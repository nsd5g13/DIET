module tm( x0,x1,x2,x3,x4,x5,x6,x7,x8,x9,x10,x11,x12,x13,x14,x15,x16,x17,x18,x19,x20,x21,x22,x23,x24,x25,x26,x27,x28,x29,x30,x31,x32,x33,x34,x35,x36,x37,x38,x39,x40,x41,x42,x43,x44,x45,x46,x47,x48,x49,x50,x51,x52,x53,x54,x55,x56,x57,x58,x59,x60,x61,x62,x63,x64,x65,x66,x67,x68,x69,x70,x71,x72,x73,x74,x75,x76,x77,x78,x79,x80,x81,x82,x83,x84,x85,x86,x87,x88,x89,x90,x91,x92,x93,x94,x95,x96,x97,x98,x99,x100,x101,x102,x103,x104,x105,x106,x107,x108,x109,x110,x111,x112,x113,x114,x115,x116,x117,x118,x119,x120,x121,x122,x123,x124,x125,x126,x127,x128,x129,x130,x131,x132,x133,x134,x135,x136,x137,x138,x139,x140,x141,x142,x143,x144,x145,x146,x147,x148,x149,x150,x151,x152,x153,x154,x155,x156,x157,x158,x159,x160,x161,x162,x163,x164,x165,x166,x167,x168,x169,x170,x171,x172,x173,x174,x175,x176,x177,x178,x179,x180,x181,x182,x183,x184,x185,x186,x187,x188,x189,x190,x191,x192,x193,x194,x195,x196,x197,x198,x199,x200,x201,x202,x203,x204,x205,x206,x207,x208,x209,x210,x211,x212,x213,x214,x215,x216,x217,x218,x219,x220,x221,x222,x223,x224,x225,x226,x227,x228,x229,x230,x231,x232,x233,x234,x235,x236,x237,x238,x239,x240,x241,x242,x243,x244,x245,x246,x247,x248,x249,x250,x251,x252,x253,x254,x255,x256,x257,x258,x259,x260,x261,x262,x263,x264,x265,x266,x267,x268,x269,x270,x271,x272,x273,x274,x275,x276,x277,x278,x279,x280,x281,x282,x283,x284,x285,x286,x287,x288,x289,x290,x291,x292,x293,x294,x295,x296,x297,x298,x299,x300,x301,x302,x303,x304,x305,x306,x307,x308,x309,x310,x311,x312,x313,x314,x315,x316,x317,x318,x319,x320,x321,x322,x323,x324,x325,x326,x327,x328,x329,x330,x331,x332,x333,x334,x335,x336,x337,x338,x339,x340,x341,x342,x343,x344,x345,x346,x347,x348,x349,x350,x351,x352,x353,x354,x355,x356,x357,x358,x359,x360,x361,x362,x363,x364,x365,x366,x367,x368,x369,x370,x371,x372,x373,x374,x375,x376,x377,x378,x379,x380,x381,x382,x383,x384,x385,x386,x387,x388,x389,x390,x391,x392,x393,x394,x395,x396,x397,x398,x399,x400,x401,x402,x403,x404,x405,x406,x407,x408,x409,x410,x411,x412,x413,x414,x415,x416,x417,x418,x419,x420,x421,x422,x423,x424,x425,x426,x427,x428,x429,x430,x431,x432,x433,x434,x435,x436,x437,x438,x439,x440,x441,x442,x443,x444,x445,x446,x447,x448,x449,x450,x451,x452,x453,x454,x455,x456,x457,x458,x459,x460,x461,x462,x463,x464,x465,x466,x467,x468,x469,x470,x471,x472,x473,x474,x475,x476,x477,x478,x479,x480,x481,x482,x483,x484,x485,x486,x487,x488,x489,x490,x491,x492,x493,x494,x495,x496,x497,x498,x499,x500,x501,x502,x503,x504,x505,x506,x507,x508,x509,x510,x511,x512,x513,x514,x515,x516,x517,x518,x519,x520,x521,x522,x523,x524,x525,x526,x527,x528,x529,x530,x531,x532,x533,x534,x535,x536,x537,x538,x539,x540,x541,x542,x543,x544,x545,x546,x547,x548,x549,x550,x551,x552,x553,x554,x555,x556,x557,x558,x559,x560,x561,x562,x563,x564,x565,x566,x567,x568,x569,x570,x571,x572,x573,x574,x575,x576,x577,x578,x579,x580,x581,x582,x583,x584,x585,x586,x587,x588,x589,x590,x591,x592,x593,x594,x595,x596,x597,x598,x599,x600,x601,x602,x603,x604,x605,x606,x607,x608,x609,x610,x611,x612,x613,x614,x615,x616,x617,x618,x619,x620,x621,x622,x623,x624,x625,x626,x627,x628,x629,x630,x631,x632,x633,x634,x635,x636,x637,x638,x639,x640,x641,x642,x643,x644,x645,x646,x647,x648,x649,x650,x651,x652,x653,x654,x655,x656,x657,x658,x659,x660,x661,x662,x663,x664,x665,x666,x667,x668,x669,x670,x671,x672,x673,x674,x675,x676,x677,x678,x679,x680,x681,x682,x683,x684,x685,x686,x687,x688,x689,x690,x691,x692,x693,x694,x695,x696,x697,x698,x699,x700,x701,x702,x703,x704,x705,x706,x707,x708,x709,x710,x711,x712,x713,x714,x715,x716,x717,x718,x719,x720,x721,x722,x723,x724,x725,x726,x727,x728,x729,x730,x731,x732,x733,x734,x735,x736,x737,x738,x739,x740,x741,x742,x743,x744,x745,x746,x747,x748,x749,x750,x751,x752,x753,x754,x755,x756,x757,x758,x759,x760,x761,x762,x763,x764,x765,x766,x767,x768,x769,x770,x771,x772,x773,x774,x775,x776,x777,x778,x779,x780,x781,x782,x783,c6228,c8114,c9123,c3431,c674,c9436,c6318,c172,c157,c2126,c6291,c7475,c8363,c5348,c051,c424,c2187,c9358,c024,c4461,c1333,c6321,c2165,c8187,c4463,c6458,c969,c1308,c6420,c9206,c4363,c918,c951,c6392,c2433,c4172,c8286,c3417,c5254,c8238,c1412,c7152,c9284,c9142,c03,c6255,c567,c416,c7125,c8369,c6441,c135,c6288,c9312,c7315,c7436,c2198,c111,c6247,c7381,c841,c0319,c2216,c3479,c0264,c0110,c7167,c1352,c7404,c6365,c22,c536,c367,c2342,c4267,c1248,c3241,c4350,c7428,c626,c5255,c3190,c537,c2145,c1360,c445,c4187,c8395,c2100,c6476,c3134,c0442,c0439,c9242,c0343,c285,c0123,c1294,c3358,c0453,c9119,c5207,c1397,c1109,c4312,c5405,c3310,c8380,c9239,c9336,c3274,c4427,c358,c947,c9191,c1379,c8139,c30,c4315,c414,c2351,c0262,c3164,c2338,c3132,c535,c062,c7180,c1256,c5171,c228,c4467,c148,c3322,c2281,c5239,c943,c133,c9155,c648,c2271,c8436,c7322,c8368,c1453,c8110,c5116,c9297,c2352,c7246,c4443,c780,c691,c3306,c3418,c295,c547,c2209,c2465,c8163,c8165,c9461,c3364,c1290,c9216,c6316,c1457,c5371,c8340,c9379,c5323,c5260,c0303,c240,c5174,c1420,c6433,c6367,c259,c7107,c188,c1262,c0426,c2200,c5480,c329,c9271,c5368,c4382,c5274,c4298,c631,c0183,c8329,c3297,c6322,c6175,c8381,c1204,c4481,c752,c066,c0108,c5411,c2252,c5271,c8401,c3143,c7266,c1179,c7429,c3126,c5242,c1380,c0178,c390,c9421,c3184,c3395,c7488,c2392,c1325,c4227,c1462,c646,c2372,c3121,c9114,c4432,c4135,c8331,c2334,c6274,c8258,c3230,c6370,c666,c4440,c2234,c874,c0357,c7396,c9225,c4434,c5182,c8151,c7358,c848,c7483,c2163,c8426,c0396,c6187,c7317,c5165,c1465,c2319,c1267,c6300,c569,c7446,c3346,c365,c359,c8105,c9230,c5412,c7355,c0417,c015,c2405,c1146,c326,c6140,c9320,c3260,c5393,c084,c0128,c12,c5406,c0189,c3379,c3137,c1466,c7173,c7103,c3426,c925,c8257,c0400,c2460,c5158,c0182,c0252,c562,c6403,c4479,c6345,c47,c039,c2263,c6385,c381,c4324,c190,c4356,c5436,c4445,c7166,c050,c3324,c891,c5431,c1284,c132,c1121,c0360,c1201,c8325,c8263,c592,c7369,c7200,c1437,c8371,c1326,c2233,c9167,c3340,c7362,c988,c1111,c297,c1175,c7150,c0298,c3456,c3138,c4352,c7468,c9373,c5367,c2361,c6327,c5347,c2404,c782,c8319,c2196,c3213,c6425,c0118,c1266,c6220,c4196,c5460,c6334,c9353,c5261,c0171,c1277,c2118,c0406,c5493,c5389,c0373,c14,c4132,c177,c893,c9209,c5491,c3487,c450,c1415,c1482,c4449,c6237,c5353,c191,c4412,c3217,c3148,c1435,c0331,c2348,c4168,c073,c8265,c252,c4188,c4270,c1142,c4224,c3160,c8162,c4292,c3116,c7473,c735,c2140,c5358,c9344,c2332,c9127,c76,c028,c8420,c8327,c3224,c0236,c9112,c9359,c210,c4208,c1239,c0391,c2250,c528,c2467,c4134,c9309,c2146,c2344,c8310,c2422,c6102,c6472,c8422,c612,c3437,c0358,c3170,c2304,c1344,c2103,c8185,c9116,c8357,c038,c8311,c4212,c0254,c5426,c3333,c5238,c0272,c4415,c4404,c8355,c7357,c5144,c3287,c5219,c235,c491,c6457,c025,c3331,c0293,c7250,c0488,c0367,c7484,c5146,c2490,c7235,c2377,c0234,c1215,c398,c1414,c5243,c8130,c7347,c7393,c7228,c964,c788,c7496,c5230,c164,c6397,c2246,c5485,c1143,c0295,c7330,c8469,c1405,c2186,c7284,c1449,c6325,c751,c6363,c5232,c5283,c0283,c7101,c5249,c747,c1145,c7236,c2458,c90,c885,c3171,c0190,c2331,c463,c534,c7132,c7297,c3149,c733,c711,c7426,c9453,c0458,c2437,c6234,c6266,c665,c1321,c4157,c57,c6418,c4381,c2474,c8296,c00,c4297,c781,c8176,c9362,c5355,c1172,c8283,c645,c8148,c0380,c2475,c0144,c7176,c9177,c336,c7239,c1167,c0411,c4102,c8215,c1370,c3470,c4181,c8440,c2341,c2318,c0258,c862,c5161,c3493,c27,c8378,c6486,c7440,c4317,c9169,c1406,c7366,c5397,c762,c6395,c6324,c911,c5398,c4314,c0223,c7211,c7187,c54,c8222,c1301,c0481,c8279,c0227,c50,c2273,c4328,c8159,c7192,c6263,c9348,c0199,c313,c2360,c3187,c5320,c9364,c5175,c963,c1305,c5432,c659,c4383,c8122,c0433,c1122,c5157,c6173,c1178,c984,c4425,c0263,c0151,c3485,c8342,c7331,c5270,c0122,c3328,c9276,c896,c4289,c5424,c790,c2430,c5107,c0469,c2413,c1350,c727,c1432,c3375,c7225,c4178,c0356,c967,c7238,c3202,c5269,c1258,c0274,c8276,c1323,c5288,c6352,c7466,c110,c7204,c1190,c0461,c4263,c1400,c6109,c9408,c4291,c5361,c5176,c5251,c9458,c8180,c7439,c5391,c493,c2419,c5478,c9473,c9341,c6482,c3407,c9361,c176,c7257,c7181,c7227,c6146,c2115,c255,c069,c0459,c6259,c3409,c865,c8367,c0164,c1383,c6319,c3102,c6139,c9143,c8494,c7442,c7435,c7291,c9433,c7373,c87,c9219,c2171,c2229,c778,c8460,c3434,c2427,c3354,c5258,c5287,c5308,c1234,c7155,c312,c1273,c2386,c4392,c7114,c8214,c6271,c1297,c9220,c2157,c2347,c3139,c554,c3243,c4269,c6353,c5240,c7280,c1320,c4332,c1300,c3350,c4290,c1282,c6130,c2366,c513,c9185,c5435,c2446,c525,c4388,c4407,c6496,c6465,c728,c0120,c6177,c0176,c597,c8271,c6176,c4229,c1193,c8421,c677,c3317,c9371,c0181,c9252,c431,c8470,c5164,c9111,c8345,c2168,c7432,c0434,c1477,c5311,c7149,c0107,c3229,c7441,c490,c6375,c7191,c8284,c0261,c0139,c638,c5233,c5417,c9422,c9391,c343,c791,c912,c7351,c9497,c4361,c640,c653,c4154,c3144,c7224,c1495,c8415,c5450,c2328,c6180,c8307,c262,c974,c121,c8416,c7161,c089,c3329,c4372,c8193,c340,c9486,c0211,c3211,c9303,c1137,c1185,c5148,c0399,c1361,c8356,c1468,c7361,c012,c2104,c8493,c7146,c0114,c4186,c366,c5145,c0218,c7324,c9465,c3394,c1268,c3474,c377,c0260,c4307,c3460,c519,c1159,c6158,c0106,c8383,c3469,c9235,c2112,c0214,c7202,c8475,c3279,c474,c729,c5322,c3408,c681,c1304,c5252,c6195,c3422,c4180,c1328,c591,c775,c35,c38,c4226,c9467,c9313,c0289,c8155,c3196,c6454,c839,c3200,c7163,c6153,c2367,c628,c9492,c8496,c4129,c80,c9176,c0207,c4391,c7140,c98,c3197,c2393,c4330,c5313,c7118,c2375,c2335,c6161,c9468,c2486,c279,c4145,c5130,c4451,c7417,c8244,c6396,c480,c1396,c5185,c6432,c4191,c45,c9446,c6142,c7186,c2236,c2218,c174,c5463,c5102,c20,c139,c0273,c9419,c2248,c8133,c6215,c8365,c1483,c7332,c9207,c0354,c4389,c4149,c8247,c134,c4378,c9187,c8134,c8390,c6218,c0378,c058,c1395,c6438,c2109,c4301,c0221,c0310,c6276,c7264,c196,c4397,c7216,c085,c3466,c9447,c6204,c819,c5290,c3244,c6303,c8439,c5235,c231,c2454,c063,c9460,c69,c1441,c161,c0268,c7499,c2150,c4336,c3482,c1331,c3406,c2483,c1182,c064,c1136,c6193,c2137,c027,c7198,c5213,c1155,c8111,c1281,c6222,c4344,c189,c2279,c8321,c4216,c7427,c9456,c5420,c7407,c5442,c1339,c0165,c1251,c6413,c9369,c1398,c5132,c2285,c394,c5197,c9200,c0168,c3351,c5481,c876,c292,c0256,c0312,c155,c0194,c2325,c5327,c5345,c3427,c3383,c1214,c01,c6243,c1438,c266,c6152,c393,c0192,c8154,c138,c7207,c7269,c2440,c9132,c6261,c1430,c1452,c1474,c7217,c8414,c5392,c9180,c153,c9316,c0487,c7212,c4244,c5256,c9228,c5241,c1424,c2388,c8211,c6148,c5275,c4170,c2181,c0389,c9168,c1358,c5246,c816,c047,c2491,c6497,c6210,c1357,c9481,c3494,c6401,c6114,c2134,c5237,c5324,c8431,c1225,c1332,c2212,c682,c8339,c1366,c4474,c8233,c686,c3262,c5369,c6308,c8452,c5133,c4232,c5396,c371,c6168,c4167,c9471,c683,c418,c6233,c5121,c581,c0270,c0322,c3313,c6178,c748,c5160,c2166,c647,c3123,c8349,c2380,c4371,c1206,c5122,c2376,c668,c7286,c6483,c3203,c9406,c5386,c9149,c1154,c4496,c6329,c2323,c737,c3491,c9282,c9337,c472,c6108,c9135,c994,c0416,c5452,c9179,c89,c8101,c6309,c8150,c6201,c042,c3468,c1244,c3207,c1355,c0478,c0425,c215,c4194,c933,c6154,c0381,c3135,c485,c6199,c7372,c6267,c0141,c7327,c126,c753,c8113,c2495,c417,c670,c234,c041,c5143,c92,c5315,c2395,c616,c9255,c3114,c4464,c6424,c4123,c3179,c044,c3236,c5490,c5217,c5404,c8246,c3248,c7348,c3338,c8240,c3352,c774,c2107,c3376,c946,c0259,c181,c8181,c6145,c8109,c1334,c2410,c5376,c9372,c0210,c4450,c8225,c4318,c898,c0448,c8387,c2400,c9248,c1115,c6227,c5263,c4251,c08,c7354,c7283,c9233,c1388,c9263,c446,c8145,c2228,c1302,c3188,c0347,c2265,c3186,c8131,c7177,c8256,c0456,c934,c9305,c043,c4271,c6171,c3218,c553,c5193,c6211,c5438,c49,c0232,c9218,c8285,c071,c694,c1410,c2421,c4437,c0444,c1375,c254,c9154,c6405,c9108,c6339,c3357,c0251,c7319,c0492,c8312,c319,c3122,c8338,c9365,c9479,c1228,c8213,c6293,c2457,c5477,c3258,c3393,c8481,c777,c9420,c9294,c5299,c3182,c9274,c1351,c9444,c769,c0484,c8178,c4494,c7292,c927,c6310,c538,c928,c3100,c8461,c741,c6400,c0250,c9355,c1336,c8202,c4230,c835,c3488,c2468,c3286,c3289,c1177,c937,c9298,c920,c7371,c2283,c166,c561,c1429,c278,c3146,c3459,c0285,c2183,c5196,c0404,c6383,c2277,c5318,c8495,c2149,c4177,c8297,c2292,c7148,c2333,c2498,c6402,c5425,c033,c4228,c0480,c1205,c9351,c5441,c6443,c5209,c9251,c4219,c7356,c272,c056,c5224,c1263,c017,c7388,c6282,c0153,c5153,c5461,c460,c5335,c936,c2471,c9134,c2299,c3360,c4320,c4109,c2113,c4438,c0422,c588,c3391,c3454,c6311,c6150,c642,c3413,c9360,c0173,c2257,c3150,c8189,c4125,c8372,c7449,c0339,c032,c4390,c281,c3298,c2431,c4242,c0371,c9477,c1106,c2215,c3129,c6284,c4343,c3425,c4419,c9430,c9171,c5325,c0238,c7410,c761,c1425,c529,c6349,c4128,c081,c29,c4176,c1488,c5104,c7433,c7376,c1257,c1158,c1218,c678,c9221,c6164,c8206,c7234,c320,c8303,c3173,c9349,c0419,c9319,c9162,c140,c6226,c3455,c9366,c5380,c7142,c4274,c2456,c7143,c734,c074,c9476,c5181,c4306,c5112,c4367,c0209,c6240,c4452,c5416,c6273,c5282,c7313,c8393,c6238,c1472,c61,c9300,c796,c1260,c2116,c7480,c8308,c3496,c973,c0338,c4160,c0241,c9270,c8465,c83,c6229,c997,c4262,c5317,c2477,c9399,c9450,c323,c5497,c3189,c1356,c8468,c5403,c91,c020,c4446,c6245,c3301,c5365,c1120,c1129,c3314,c6197,c6250,c0477,c9189,c1411,c7392,c1247,c3118,c4385,c742,c5401,c82,c7124,c9104,c1431,c325,c6407,c1377,c2173,c7308,c9402,c5387,c8216,c6217,c7231,c8212,c4200,c1107,c1157,c7300,c1455,c116,c9292,c437,c6398,c4152,c3450,c2379,c4490,c8483,c853,c1187,c1135,c4447,c9435,c4468,c855,c1209,c3294,c3227,c3133,c4342,c9172,c2359,c837,c7121,c076,c3337,c982,c0301,c861,c4300,c128,c4264,c7398,c0271,c2220,c342,c4201,c975,c9334,c459,c2309,c3449,c3288,c7482,c7312,c8434,c3446,c016,c3204,c7119,c2424,c5225,c8277,c337,c0111,c671,c866,c840,c0413,c4250,c335,c9449,c8245,c8300,c3467,c990,c6358,c7271,c0397,c4472,c2462,c5203,c061,c0246,c9363,c7259,c643,c1163,c7465,c4115,c870,c8249,c034,c8457,c249,c4430,c1387,c486,c9105,c379,c3208,c8294,c8264,c6434,c5278,c4210,c0196,c8104,c1443,c673,c1108,c6181,c3119,c2358,c851,c2194,c380,c9266,c5150,c3445,c976,c4414,c3442,c2355,c4294,c883,c0309,c355,c9144,c2232,c3181,c0208,c433,c7287,c7136,c5247,c881,c0318,c0320,c0133,c1133,c622,c4153,c4100,c6467,c3273,c4101,c784,c4235,c4260,c8194,c362,c1296,c6242,c4222,c4423,c8118,c699,c4357,c2364,c0226,c1403,c6131,c7333,c013,c1364,c593,c797,c2432,c4364,c36,c744,c2385,c5201,c9434,c6491,c842,c9247,c8322,c7273,c5192,c7249,c0186,c51,c579,c8313,c6448,c3414,c4454,c059,c28,c299,c4249,c9464,c724,c4202,c6409,c710,c8444,c3219,c257,c5245,c4106,c9498,c5292,c0436,c6290,c0355,c0286,c1197,c481,c7405,c6464,c24,c6384,c9438,c8455,c4341,c949,c3464,c026,c2139,c6185,c9193,c0311,c0281,c7141,c2230,c9317,c8441,c7452,c772,c8438,c726,c167,c9385,c1434,c7457,c018,c4253,c8499,c63,c091,c521,c324,c9454,c3268,c8250,c0342,c1354,c7203,c6213,c0253,c5453,c766,c387,c8100,c1433,c598,c9152,c1275,c3107,c7215,c2258,c4205,c1419,c7294,c466,c9389,c6184,c6307,c8405,c3278,c542,c4238,c7251,c3371,c1480,c6147,c5366,c5340,c5162,c5421,c9326,c9472,c9140,c7343,c9126,c0465,c3277,c269,c7290,c2175,c6451,c9368,c4359,c5306,c05,c4442,c080,c6393,c635,c4127,c4141,c3257,c9384,c6332,c6183,c5456,c867,c487,c9401,c4116,c6380,c6455,c5328,c2420,c4418,c6492,c9329,c1186,c8409,c467,c5468,c1324,c684,c1211,c7174,c625,c7178,c5291,c0288,c8209,c2156,c7316,c779,c0490,c552,c0160,c494,c2288,c6326,c2287,c0294,c7477,c220,c5152,c9459,c3388,c0155,c5128,c88,c1440,c1110,c159,c341,c9416,c8182,c9211,c0138,c5140,c0179,c2193,c6360,c8124,c3315,c0102,c224,c4111,c0430,c6337,c6192,c9466,c0146,c3372,c545,c2448,c945,c7419,c75,c7494,c55,c1184,c8161,c7345,c2415,c3478,c8289,c9295,c2345,c7460,c0486,c9146,c8464,c9310,c0170,c2481,c617,c5314,c9491,c9345,c2214,c6470,c7123,c1224,c8183,c6423,c833,c8323,c5208,c6138,c64,c1363,c1487,c2151,c5331,c7253,c0121,c3448,c8385,c1390,c764,c8391,c584,c844,c627,c5429,c798,c356,c636,c875,c4273,c6125,c9396,c85,c5142,c4406,c2106,c169,c0224,c3327,c1313,c9136,c9288,c2174,c773,c3498,c9262,c610,c7413,c0427,c1232,c6372,c8230,c2199,c3240,c8449,c5105,c2164,c9121,c634,c6236,c7382,c4497,c8166,c3339,c1311,c2224,c2423,c2256,c8291,c0388,c2301,c892,c4422,c8482,c094,c2136,c7350,c745,c2321,c3403,c4174,c451,c1348,c1295,c8208,c090,c1494,c2203,c369,c859,c6331,c2225,c274,c125,c5344,c4433,c4183,c971,c060,c9208,c4351,c6453,c6468,c1243,c5336,c4482,c2221,c1322,c5390,c311,c9101,c6422,c7138,c8266,c8471,c163,c3433,c2414,c623,c2298,c07,c2213,c0491,c3225,c6298,c6350,c749,c498,c9400,c1342,c2195,c9267,c4223,c9124,c7258,c669,c9327,c1490,c4248,c4444,c5149,c2390,c1194,c1309,c482,c3400,c8108,c6117,c6335,c716,c2231,c0368,c576,c4254,c5114,c9426,c6182,c154,c821,c1303,c9286,c655,c9299,c6160,c2499,c792,c84,c7193,c0372,c1404,c4287,c7171,c0150,c0277,c3261,c5302,c7218,c965,c8195,c2311,c695,c8253,c9229,c149,c0324,c0316,c1338,c3444,c1134,c5451,c0455,c4466,c495,c1448,c4215,c8190,c9291,c873,c7377,c2397,c1207,c8232,c0359,c4347,c1255,c578,c675,c2177,c2492,c9390,c1409,c6368,c3155,c7285,c4398,c8354,c310,c232,c688,c1407,c7311,c1235,c8462,c3152,c8324,c443,c2312,c2238,c9490,c4150,c5499,c6436,c7260,c1114,c8374,c4151,c568,c6260,c7220,c8361,c8419,c144,c680,c395,c2317,c5212,c5188,c1213,c7490,c375,c3304,c6444,c7303,c0112,c0364,c5298,c8358,c7233,c6404,c7370,c541,c6264,c1233,c5297,c3463,c233,c9393,c512,c7455,c321,c9495,c551,c8411,c421,c7214,c5400,c813,c6437,c2494,c2396,c9383,c5250,c2211,c8293,c271,c879,c353,c1270,c6488,c2455,c9480,c3252,c1253,c3141,c721,c399,c8382,c6354,c651,c2223,c7219,c0497,c4107,c4354,c2293,c0228,c317,c2417,c9437,c4217,c8337,c2429,c6330,c882,c1471,c7338,c1436,c1470,c057,c488,c0229,c7244,c5115,c5309,c373,c9203,c1408,c5177,c0161,c894,c0332,c9272,c0105,c4221,c3125,c983,c2276,c924,c10,c3157,c4280,c282,c3348,c62,c6257,c1450,c2408,c9264,c978,c010,c2192,c253,c1164,c2435,c7352,c198,c4182,c621,c550,c7461,c9215,c0222,c1489,c3282,c5356,c229,c0370,c6151,c0405,c088,c6373,c7272,c5330,c2451,c3386,c60,c5119,c4345,c152,c7448,c1393,c0424,c5155,c1269,c6133,c3457,c065,c9380,c6427,c8174,c5190,c3145,c868,c1138,c316,c383,c5284,c6129,c558,c6299,c4105,c419,c5377,c7487,c1166,c7105,c8295,c1212,c150,c429,c2470,c9201,c1337,c6202,c6254,c663,c123,c595,c3490,c817,c3336,c2204,c2154,c4218,c2217,c757,c1285,c4448,c6328,c594,c9170,c7464,c7438,c9487,c0390,c4321,c5312,c2227,c5489,c2268,c428,c4118,c845,c2152,c7275,c5388,c4487,c298,c2306,c2120,c8201,c6265,c1287,c836,c0245,c014,c7342,c5257,c8418,c4256,c3345,c880,c0374,c1230,c4485,c9424,c42,c171,c9387,c0284,c331,c7172,c4272,c6301,c6498,c5352,c1189,c4376,c856,c265,c7380,c4309,c8404,c8445,c5455,c9181,c9249,c9174,c5221,c0149,c1341,c5462,c9130,c6388,c8343,c368,c0197,c6110,c96,c4455,c1418,c6305,c5191,c7276,c0350,c3390,c4386,c425,c570,c5482,c114,c226,c193,c583,c0414,c6246,c0363,c2439,c6118,c6351,c812,c5458,c040,c8466,c3447,c0129,c0101,c5214,c3458,c8346,c0115,c3384,c9175,c2478,c2484,c6382,c6297,c1156,c6295,c2260,c79,c864,c9241,c0131,c7184,c9443,c7168,c6359,c8486,c7100,c2123,c396,c7254,c2340,c629,c0384,c1274,c2142,c330,c9245,c8158,c8477,c2450,c7113,c8226,c1279,c1219,c7395,c1132,c8373,c0117,c5343,c9137,c8453,c5100,c8443,c9273,c1381,c1496,c1116,c644,c16,c0454,c9159,c7188,c6107,c4304,c8137,c7112,c2329,c430,c1319,c4288,c7375,c8146,c8478,c5362,c5423,c9244,c9269,c4198,c7221,c243,c8184,c3486,c77,c3370,c1139,c2247,c4353,c3285,c7199,c7262,c8171,c6156,c284,c2438,c230,c2434,c6104,c566,c2416,c0449,c1130,c7296,c248,c3318,c5248,c793,c0483,c8447,c2270,c5117,c0437,c3497,c0315,c6466,c4410,c5360,c5349,c2180,c4373,c794,c1176,c5449,c713,c939,c2286,c3130,c9342,c3162,c0267,c8309,c4126,c0348,c818,c7344,c4133,c0201,c6341,c349,c3106,c9413,c8251,c7222,c7242,c3265,c453,c4234,c979,c3205,c1464,c7110,c3233,c820,c4394,c814,c574,c048,c5498,c5163,c944,c0498,c0475,c3451,c8410,c5409,c850,c7456,c4137,c5183,c6231,c5494,c4339,c977,c9165,c9439,c2473,c7368,c9107,c2373,c8364,c0452,c0466,c2464,c5151,c8129,c4147,c637,c9315,c449,c8379,c1202,c9147,c115,c6203,c0290,c0443,c2108,c286,c0330,c3246,c9452,c889,c0365,c4284,c8254,c8141,c4247,c2482,c075,c9258,c9217,c8304,c74,c8204,c6387,c6230,c4282,c543,c895,c4473,c3436,c0145,c9339,c3271,c872,c7412,c2313,c6333,c7116,c3397,c0328,c9287,c0314,c6191,c4416,c5483,c9431,c7443,c7423,c8456,c9198,c3234,c2222,c687,c3465,c9346,c098,c9445,c046,c6285,c218,c3153,c9182,c5173,c6374,c082,c5342,c0313,c0403,c9268,c5228,c2280,c650,c093,c654,c810,c966,c6221,c473,c1291,c6188,c2244,c4265,c0167,c5445,c5200,c0195,c478,c6281,c5427,c7205,c0156,c7241,c926,c9280,c0193,c6120,c9103,c8128,c3326,c0428,c6278,c4243,c095,c65,c2330,c2350,c2479,c0126,c3283,c6313,c0474,c357,c8442,c799,c1173,c0216,c1148,c4483,c2307,c8392,c0407,c5448,c630,c439,c7156,c3180,c3411,c1386,c7120,c26,c3499,c3323,c696,c6394,c2487,c1151,c6214,c9214,c492,c0386,c7268,c192,c2445,c8107,c333,c991,c8458,c160,c831,c1174,c1373,c4338,c913,c9238,c3172,c4316,c6296,c4486,c5180,c2133,c1497,c8402,c5296,c5307,c7209,c130,c5134,c4495,c1298,c8472,c2409,c0296,c4213,c4268,c9441,c6244,c1413,c5469,c5495,c338,c4156,c0113,c0127,c021,c1499,c6100,c0327,c2346,c9102,c2255,c7397,c5187,c3423,c7365,c8341,c9236,c7109,c9304,c2153,c921,c3161,c2442,c3303,c6223,c0282,c7261,c7389,c464,c613,c5373,c6495,c3292,c5439,c693,c442,c2128,c0334,c9223,c6406,c3489,c0206,c9378,c7318,c722,c3359,c8328,c4322,c8248,c531,c712,c7196,c9493,c522,c8123,c0134,c6141,c3247,c1238,c910,c3183,c413,c6447,c0352,c136,c4275,c0174,c6442,c2466,c2406,c3284,c0418,c932,c9139,c5472,c2132,c998,c8359,c7485,c5156,c6165,c1369,c5231,c1402,c7479,c9307,c5210,c877,c5382,c3201,c096,c3169,c4402,c2208,c4491,c0412,c070,c4240,c4112,c1126,c59,c941,c1426,c9110,c0103,c1153,c2274,c1371,c5341,c0239,c156,c2111,c241,c376,c8168,c270,c6489,c8430,c4368,c34,c9333,c238,c6209,c4457,c7245,c6386,c2162,c4384,c9183,c0220,c8102,c9409,c4492,c345,c9425,c9194,c4370,c0485,c4146,c389,c354,c4334,c572,c0462,c6484,c6494,c4175,c948,c247,c1299,c826,c556,c3415,c7147,c4225,c7425,c7411,c0317,c5211,c1327,c660,c4326,c9397,c4380,c5466,c6348,c496,c6371,c3254,c5338,c7248,c2249,c6304,c2489,c1374,c5354,c6159,c0409,c5364,c1368,c2262,c4236,c410,c3378,c147,c162,c9415,c43,c8492,c771,c8432,c378,c8425,c7495,c9178,c2296,c9128,c239,c0337,c3341,c0304,c6411,c8223,c4358,c9482,c6338,c5476,c322,c0445,c0175,c9250,c2259,c7498,c1198,c6128,c564,c1168,c3483,c3101,c5384,c972,c438,c1261,c6206,c8398,c0269,c6251,c596,c9311,c458,c2387,c2371,c7445,c3275,c3305,c6163,c587,c9293,c350,c9164,c2202,c7164,c8116,c4211,c4325,c5206,c0476,c2117,c9308,c1180,c2122,c7384,c3264,c4179,c8488,c656,c99,c8126,c1312,c2444,c0300,c573,c3342,c0217,c5418,c6121,c3267,c755,c672,c641,c7129,c3251,c1118,c5170,c4163,c4360,c7309,c6170,c6112,c1389,c9318,c3389,c9279,c0140,c6174,c277,c2197,c540,c7165,c915,c539,c4498,c5279,c6355,c619,c5118,c4148,c9347,c8149,c1445,c0432,c4499,c8491,c0159,c5124,c441,c3280,c9350,c9412,c6449,c7267,c4299,c1278,c786,c2169,c9278,c7162,c15,c011,c3361,c9370,c9405,c9145,c3178,c3471,c4237,c577,c4375,c2160,c0429,c225,c7158,c8484,c1103,c731,c7401,c8451,c0470,c0333,c9381,c3396,c9129,c5444,c8450,c2353,c2357,c4185,c117,c9256,c9474,c8336,c5381,c2412,c372,c1223,c9117,c0460,c6224,c863,c1196,c151,c5474,c415,c9234,c7335,c3212,c5285,c3419,c1252,c9374,c95,c785,c1112,c173,c4117,c2303,c6408,c3402,c6487,c1192,c477,c5159,c4458,c5329,c6399,c8186,c146,c9163,c8205,c7307,c9325,c6306,c1127,c633,c0495,c9260,c1199,c0148,c5262,c2125,c48,c849,c1427,c5138,c1498,c6478,c6115,c9489,c0266,c0125,c0450,c3309,c5113,c8423,c078,c092,c7106,c0440,c3195,c7133,c0335,c3362,c6126,c6480,c3440,c0177,c3363,c4131,c2121,c763,c3477,c4104,c559,c142,c8317,c3109,c1330,c0130,c3473,c9306,c184,c219,c1479,c9224,c1444,c3302,c7390,c3245,c7444,c072,c120,c3321,c931,c4124,c9485,c7418,c1399,c183,c411,c3462,c3216,c0472,c530,c9328,c6473,c6429,c0198,c0275,c0415,c714,c7201,c099,c7135,c9418,c5321,c8489,c351,c8192,c7194,c25,c8261,c8127,c7470,c4305,c4246,c8302,c1451,c7127,c1171,c0242,c1131,c9494,c8229,c7471,c823,c4417,c4209,c273,c8260,c8282,c127,c7408,c3476,c4308,c9283,c2272,c5437,c2327,c8164,c8389,c461,c5265,c1378,c7422,c8200,c740,c41,c560,c5276,c447,c4319,c5281,c811,c5410,c954,c2267,c7493,c3250,c420,c2300,c4293,c5370,c4428,c131,c2239,c1485,c6459,c1101,c8210,c2110,c386,c9411,c5399,c9354,c8288,c9141,c765,c6315,c9115,c4144,c3399,c6122,c1307,c7229,c1439,c1125,c8239,c9398,c6232,c3296,c0243,c296,c3308,c6456,c8386,c720,c7263,c237,c3110,c7336,c4302,c391,c599,c5433,c2219,c334,c3412,c5103,c3113,c5186,c0464,c9243,c9184,c533,c5111,c7450,c81,c3255,c2389,c4426,c4436,c5407,c4335,c6317,c31,c8221,c532,c3192,c4257,c689,c7131,c455,c956,c4255,c211,c6194,c514,c9407,c7489,c555,c5205,c7145,c9392,c7183,c118,c1124,c8463,c1227,c8314,c6190,c658,c8400,c7421,c2411,c999,c5272,c5459,c9289,c9153,c0375,c412,c7491,c6155,c3270,c3165,c3381,c3168,c8474,c3349,c6471,c9240,c5169,c212,c1385,c036,c8394,c0369,c53,c4245,c7364,c9151,c4329,c4489,c0353,c9296,c5227,c7139,c0237,c0280,c4161,c3366,c213,c1421,c8448,c1183,c986,c6378,c3405,c3325,c6343,c5167,c5216,c3356,c2241,c5402,c6249,c6103,c71,c2322,c7387,c5277,c3295,c922,c5428,c8428,c347,c214,c828,c2391,c5351,c5357,c483,c8117,c4108,c8236,c3198,c0279,c0383,c8231,c9156,c2291,c9138,c0431,c8219,c6113,c0257,c2243,c7329,c4261,c2189,c9195,c4214,c4171,c476,c3147,c0341,c1140,c4259,c216,c384,c2441,c223,c2266,c8417,c2131,c1246,c1493,c5204,c6361,c7301,c3334,c2235,c5289,c5229,c9161,c32,c5496,c3185,c4424,c9386,c1365,c388,c6474,c6435,c7255,c434,c067,c3404,c5136,c8156,c3151,c586,c1473,c4475,c3175,c9457,c0408,c2428,c0394,c5473,c2399,c4122,c2354,c2349,c7126,c3269,c8121,c4195,c2297,c5363,c6414,c0233,c5101,c6416,c1229,c0244,c897,c3166,c3108,c5198,c3416,c6270,c9113,c3253,c9133,c8115,c987,c8287,c9222,c119,c7406,c1484,c7274,c834,c6101,c1102,c7117,c8326,c4296,c9483,c815,c9427,c959,c4142,c9192,c5359,c4190,c9428,c9338,c3140,c1492,c145,c1264,c465,c1236,c1428,c8454,c961,c9440,c923,c6280,c8273,c516,c4480,c5131,c611,c698,c5172,c0249,c2310,c8172,c2182,c0152,c8320,c0326,c3276,c8384,c0421,c649,c0143,c4279,c185,c5178,c6248,c0299,c471,c2402,c3194,c5374,c6149,c5375,c4239,c4233,c6336,c2449,c426,c4377,c6428,c0395,c457,c250,c1220,c2370,c7323,c7295,c267,c168,c73,c9210,c217,c5109,c886,c5430,c8353,c180,c5434,c3163,c7282,c952,c8177,c5259,c878,c8375,c8435,c575,c7374,c8267,c4493,c4348,c7467,c5454,c1353,c2148,c0116,c58,c9404,c7434,c423,c970,c940,c6450,c3256,c2205,c314,c8135,c9277,c523,c9188,c288,c4469,c9432,c1416,c1271,c8199,c2210,c995,c33,c9356,c957,c5446,c5415,c6493,c7208,c758,c186,c5223,c1149,c6485,c370,c294,c3104,c2382,c7481,c11,c1265,c4413,c9322,c5184,c8479,c141,c4403,c0336,c0387,c2493,c2284,c2158,c275,c6460,c5218,c950,c4189,c4399,c719,c8301,c263,c515,c8143,c0276,c3158,c517,c3176,c9463,c1423,c3249,c268,c759,c0204,c3210,c7325,c1442,c7403,c4158,c7210,c7320,c8348,c9265,c5379,c8170,c019,c5475,c4155,c0438,c1372,c871,c993,c5457,c4387,c3136,c0137,c7476,c2426,c9324,c6269,c4393,c030,c8480,c589,c9499,c8147,c5487,c6169,c385,c4281,c0215,c94,c053,c260,c9462,c738,c6412,c1141,c6462,c9302,c6134,c1289,c0172,c9125,c8412,c7170,c2159,c9377,c7424,c7169,c7189,c3435,c361,c4285,c1345,c462,c756,c9376,c0401,c9301,c2245,c2305,c049,c3120,c037,c2170,c1283,c5484,c3438,c8362,c7302,c469,c1161,c8169,c8106,c5333,c3424,c1458,c8227,c916,c884,c9475,c6189,c2343,c1237,c4197,c664,c4355,c452,c8298,c1276,c055,c4173,c7334,c2485,c4139,c2362,c427,c8335,c1123,c7281,c283,c7337,c9340,c8173,c3263,c78,c4313,c6440,c8280,c5141,c917,c7363,c795,c887,c2383,c4456,c685,c0349,c112,c930,c9357,c5422,c4206,c914,c6379,c9205,c195,c6143,c5266,c67,c06,c8408,c6314,c222,c2326,c5300,c5339,c4311,c9367,c770,c0169,c725,c1314,c4462,c7197,c7472,c7122,c7328,c0157,c4374,c3385,c6431,c8388,c364,c3387,c776,c1335,c5319,c8196,c5139,c5179,c8262,c2179,c6286,c5326,c6294,c352,c1343,c9157,c7289,c3420,c4140,c717,c6256,c0265,c0292,c1165,c397,c290,c0180,c3127,c287,c8397,c6235,c1286,c4362,c3432,c0321,c7339,c293,c2295,c0457,c639,c7195,c6390,c236,c0435,c0135,c251,c2339,c2124,c4231,c5470,c5135,c0212,c9118,c624,c1152,c4165,c829,c0119,c9451,c5372,c3221,c548,c942,c8237,c3307,c7279,c9254,c276,c9442,c8476,c0231,c077,c962,c3443,c0100,c8198,c9173,c5147,c5395,c8473,c2302,c2401,c5126,c4303,c8347,c3124,c175,c087,c9388,c1475,c6347,c2167,c860,c0142,c3105,c520,c8281,c245,c0191,c0467,c3222,c4295,c1280,c8278,c1117,c888,c5253,c8485,c346,c7230,c2384,c2315,c8407,c7277,c3332,c843,c6106,c2242,c1100,c5316,c0420,c0225,c6312,c767,c8437,c256,c9150,c4346,c8370,c04,c1310,c5440,c199,c2155,c3177,c113,c2425,c197,c6258,c5486,c9455,c21,c4278,c2251,c8217,c18,c8224,c6356,c09,c0185,c4331,c3429,c8228,c2201,c5394,c8272,c7102,c657,c4477,c37,c3480,c1316,c7431,c484,c4114,c4366,c9131,c9417,c0377,c3430,c4277,c955,c9281,c7453,c825,c475,c444,c8274,c5154,c46,c2190,c6481,c3228,c5334,c6479,c7265,c7367,c8487,c2407,c6262,c690,c70,c929,c4162,c1293,c0323,c6376,c5108,c5215,c1417,c6346,c9197,c0393,c3259,c838,c079,c8433,c847,c0109,c2119,c3232,c7226,c2207,c632,c6123,c960,c5294,c1469,c2316,c7153,c6116,c3320,c1401,c66,c3193,c39,c6417,c8241,c0473,c7232,c6225,c4113,c2394,c3380,c5137,c1478,c7378,c518,c3111,c4337,c0278,c4207,c938,c9213,c7151,c031,c3131,c8235,c6137,c5264,c6369,c2114,c715,c730,c8406,c8153,c2459,c4435,c5195,c2356,c852,c1491,c3441,c6289,c3421,c2453,c7399,c9448,c0306,c5236,c1249,c2290,c3472,c7486,c122,c6205,c3319,c6186,c4203,c4453,c0493,c7104,c3242,c546,c2237,c1318,c3347,c7154,c8234,c5189,c2447,c0247,c5488,c0361,c7379,c9109,c8366,c6364,c746,c9237,c5346,c470,c5222,c6268,c827,c6463,c8330,c0392,c3365,c5295,c1104,c8427,c9394,c6357,c93,c3484,c3215,c620,c5337,c2469,c8290,c0205,c3103,c7341,c8197,c1231,c8351,c9429,c6499,c2172,c3266,c527,c1240,c0305,c9246,c029,c1162,c0496,c2443,c4400,c194,c6302,c2185,c5194,c3281,c6272,c1245,c6241,c2176,c9331,c178,c2282,c2476,c6323,c0482,c1242,c9330,c2496,c1170,c3439,c3300,c0446,c3154,c2381,c9285,c1272,c4401,c0297,c2147,c557,c2264,c0494,c2480,c3316,c5414,c4169,c9469,c6212,c360,c9335,c6124,c0235,c8138,c3398,c3335,c2289,c02,c989,c1222,c8175,c9120,c526,c8360,c7185,c919,c3167,c2374,c3368,c291,c7454,c3237,c4121,c4409,c8269,c0163,c996,c332,c8125,c9106,c0188,c022,c676,c1317,c5273,c1226,c9232,c511,c0308,c9410,c9259,c7414,c9290,c382,c2101,c1200,c1188,c2363,c0451,c280,c6219,c8218,c3226,c4103,c5123,c5443,c7306,c8413,c4441,c0213,c2365,c723,c958,c5310,c182,c7451,c7353,c4258,c8424,c9257,c2278,c9321,c227,c510,c4470,c6381,c4395,c1315,c1359,c2143,c318,c4488,c7137,c2452,c0346,c2184,c8179,c7416,c1367,c8207,c8120,c2436,c4136,c1447,c0124,c0489,c3312,c0447,c1347,c8429,c0132,c8332,c8446,c289,c1376,c4286,c1181,c9212,c858,c392,c9253,c0154,c8490,c3238,c6475,c6340,c822,c4310,c5244,c5125,c499,c0441,c5492,c8396,c8203,c7478,c0187,c435,c436,c2144,c6366,c8352,c187,c0329,c7278,c0479,c2261,c221,c5110,c7298,c9202,c9470,c9166,c035,c2188,c4429,c5304,c7463,c824,c7223,c8350,c5408,c327,c0104,c9375,c5305,c5447,c9488,c2314,c8140,c8315,c2178,c045,c5419,c6342,c4349,c6389,c4266,c1456,c2488,c4138,c6279,c7310,c1119,c6445,c5464,c8259,c2324,c5129,c3392,c9484,c732,c1446,c468,c7115,c0471,c6415,c0184,c935,c17,c9275,c3290,c3367,c6132,c315,c9190,c083,c5268,c8255,c8299,c1203,c7409,c2253,c4166,c1195,c1250,c8119,c6446,c1217,c56,c489,c3220,c6200,c0200,c6166,c8167,c9352,c0423,c086,c3199,c4333,c8112,c2336,c9100,c258,c7243,c2369,c9261,c1467,c422,c1216,c456,c9323,c7469,c739,c5280,c3410,c6391,c170,c692,c0366,c3117,c8306,c5350,c448,c7293,c8188,c1394,c585,c9148,c9204,c563,c4411,c3344,c2378,c2105,c9196,c1221,c0385,c0410,c5127,c7385,c054,c1391,c652,c667,c7447,c44,c750,c9227,c052,c6196,c614,c3156,c899,c8132,c143,c6136,c6157,c4369,c7462,c4484,c8144,c4431,c3209,c830,c618,c571,c1340,c6430,c0248,c3353,c7394,c4204,c832,c565,c5303,c2141,c544,c6469,c0345,c582,c7157,c6362,c4420,c1384,c5413,c5199,c736,c3235,c7420,c4379,c0307,c4252,c7314,c7159,c846,c4460,c0219,c8459,c7458,c3293,c7134,c5471,c0255,c615,c3369,c7346,c7179,c8334,c9332,c3159,c0325,c754,c5293,c4241,c9382,c7326,c0202,c0382,c1349,c1169,c7415,c339,c8152,c52,c9423,c1241,c7270,c985,c3355,c789,c2472,c7182,c3206,c165,c3115,c3377,c3174,c3311,c7237,c3481,c2308,c1128,c7321,c6377,c2161,c1160,c6105,c2206,c1147,c7359,c7144,c6208,c854,c3223,c7430,c0240,c2368,c1254,c3299,c6239,c2463,c2191,c8399,c2461,c857,c440,c2127,c1461,c86,c8333,c3191,c1329,c5479,c2226,c1144,c8498,c992,c4283,c0351,c9122,c1459,c4439,c9403,c2337,c0499,c1460,c0291,c4193,c1382,c768,c3495,c1486,c40,c7288,c7256,c8243,c0468,c8275,c1362,c4164,c242,c8403,c6490,c137,c760,c129,c2269,c3231,c8191,c1476,c7386,c023,c9395,c5332,c7130,c124,c7190,c7402,c6252,c1392,c7252,c7304,c6439,c0162,c479,c6111,c2403,c6216,c5106,c2129,c432,c9199,c1113,c497,c5286,c0402,c981,c8103,c2130,c524,c4365,c7474,c5234,c783,c3401,c6144,c679,c1259,c6127,c1306,c4130,c1105,c3461,c4119,c5383,c6179,c2254,c5467,c1191,c9186,c743,c7240,c0158,c4459,c2275,c8270,c5385,c0302,c6162,c6426,c5168,c3214,c2398,c7305,c1288,c8142,c6135,c1208,c6172,c0362,c662,c179,c6207,c4465,c7459,c7206,c580,c2138,c261,c9478,c97,c9160,c454,c7247,c8220,c4323,c6198,c6320,c9226,c0340,c6167,c0379,c6119,c4184,c3382,c068,c328,c3428,c3239,c4192,c2240,c3330,c6275,c2102,c6277,c9496,c3291,c3475,c8242,c661,c158,c7349,c4120,c3492,c0203,c8157,c72,c7128,c3112,c6283,c1346,c7492,c4421,c5465,c8318,c363,c2497,c7360,c980,c3453,c5226,c0376,c9231,c4159,c68,c6452,c9414,c968,c4220,c6253,c8292,c244,c1481,c3128,c0287,c8467,c097,c7175,c9158,c718,c0136,c0166,c8377,c787,c6287,c7108,c1422,c19,c7497,c549,c8252,c2294,c8376,c7391,c5378,c7111,c590,c6419,c953,c7213,c4110,c4408,c5120,c9314,c1210,c4405,c7437,c23,c374,c869,c4476,c3142,c7299,c4478,c0463,c7160,c7400,c3272,c9343,c2135,c6344,c5267,c6477,c344,c3343,c4471,c1292,c6461,c8497,c5202,c5166,c4396,c1150,c0147,c8316,c7340,c6421,c2418,c6292,c5220,c1463,c4340,c4199,c3374,c0344,c264,c3452,c3373,c8136,c8344,c8305,c1454,c8268,c13,c348,c4327,c4276,c2320,c5301,c6410,c0230,c0398,c697,c890,c8160,c246,c4143,c7383 );

input x0;
input x1;
input x2;
input x3;
input x4;
input x5;
input x6;
input x7;
input x8;
input x9;
input x10;
input x11;
input x12;
input x13;
input x14;
input x15;
input x16;
input x17;
input x18;
input x19;
input x20;
input x21;
input x22;
input x23;
input x24;
input x25;
input x26;
input x27;
input x28;
input x29;
input x30;
input x31;
input x32;
input x33;
input x34;
input x35;
input x36;
input x37;
input x38;
input x39;
input x40;
input x41;
input x42;
input x43;
input x44;
input x45;
input x46;
input x47;
input x48;
input x49;
input x50;
input x51;
input x52;
input x53;
input x54;
input x55;
input x56;
input x57;
input x58;
input x59;
input x60;
input x61;
input x62;
input x63;
input x64;
input x65;
input x66;
input x67;
input x68;
input x69;
input x70;
input x71;
input x72;
input x73;
input x74;
input x75;
input x76;
input x77;
input x78;
input x79;
input x80;
input x81;
input x82;
input x83;
input x84;
input x85;
input x86;
input x87;
input x88;
input x89;
input x90;
input x91;
input x92;
input x93;
input x94;
input x95;
input x96;
input x97;
input x98;
input x99;
input x100;
input x101;
input x102;
input x103;
input x104;
input x105;
input x106;
input x107;
input x108;
input x109;
input x110;
input x111;
input x112;
input x113;
input x114;
input x115;
input x116;
input x117;
input x118;
input x119;
input x120;
input x121;
input x122;
input x123;
input x124;
input x125;
input x126;
input x127;
input x128;
input x129;
input x130;
input x131;
input x132;
input x133;
input x134;
input x135;
input x136;
input x137;
input x138;
input x139;
input x140;
input x141;
input x142;
input x143;
input x144;
input x145;
input x146;
input x147;
input x148;
input x149;
input x150;
input x151;
input x152;
input x153;
input x154;
input x155;
input x156;
input x157;
input x158;
input x159;
input x160;
input x161;
input x162;
input x163;
input x164;
input x165;
input x166;
input x167;
input x168;
input x169;
input x170;
input x171;
input x172;
input x173;
input x174;
input x175;
input x176;
input x177;
input x178;
input x179;
input x180;
input x181;
input x182;
input x183;
input x184;
input x185;
input x186;
input x187;
input x188;
input x189;
input x190;
input x191;
input x192;
input x193;
input x194;
input x195;
input x196;
input x197;
input x198;
input x199;
input x200;
input x201;
input x202;
input x203;
input x204;
input x205;
input x206;
input x207;
input x208;
input x209;
input x210;
input x211;
input x212;
input x213;
input x214;
input x215;
input x216;
input x217;
input x218;
input x219;
input x220;
input x221;
input x222;
input x223;
input x224;
input x225;
input x226;
input x227;
input x228;
input x229;
input x230;
input x231;
input x232;
input x233;
input x234;
input x235;
input x236;
input x237;
input x238;
input x239;
input x240;
input x241;
input x242;
input x243;
input x244;
input x245;
input x246;
input x247;
input x248;
input x249;
input x250;
input x251;
input x252;
input x253;
input x254;
input x255;
input x256;
input x257;
input x258;
input x259;
input x260;
input x261;
input x262;
input x263;
input x264;
input x265;
input x266;
input x267;
input x268;
input x269;
input x270;
input x271;
input x272;
input x273;
input x274;
input x275;
input x276;
input x277;
input x278;
input x279;
input x280;
input x281;
input x282;
input x283;
input x284;
input x285;
input x286;
input x287;
input x288;
input x289;
input x290;
input x291;
input x292;
input x293;
input x294;
input x295;
input x296;
input x297;
input x298;
input x299;
input x300;
input x301;
input x302;
input x303;
input x304;
input x305;
input x306;
input x307;
input x308;
input x309;
input x310;
input x311;
input x312;
input x313;
input x314;
input x315;
input x316;
input x317;
input x318;
input x319;
input x320;
input x321;
input x322;
input x323;
input x324;
input x325;
input x326;
input x327;
input x328;
input x329;
input x330;
input x331;
input x332;
input x333;
input x334;
input x335;
input x336;
input x337;
input x338;
input x339;
input x340;
input x341;
input x342;
input x343;
input x344;
input x345;
input x346;
input x347;
input x348;
input x349;
input x350;
input x351;
input x352;
input x353;
input x354;
input x355;
input x356;
input x357;
input x358;
input x359;
input x360;
input x361;
input x362;
input x363;
input x364;
input x365;
input x366;
input x367;
input x368;
input x369;
input x370;
input x371;
input x372;
input x373;
input x374;
input x375;
input x376;
input x377;
input x378;
input x379;
input x380;
input x381;
input x382;
input x383;
input x384;
input x385;
input x386;
input x387;
input x388;
input x389;
input x390;
input x391;
input x392;
input x393;
input x394;
input x395;
input x396;
input x397;
input x398;
input x399;
input x400;
input x401;
input x402;
input x403;
input x404;
input x405;
input x406;
input x407;
input x408;
input x409;
input x410;
input x411;
input x412;
input x413;
input x414;
input x415;
input x416;
input x417;
input x418;
input x419;
input x420;
input x421;
input x422;
input x423;
input x424;
input x425;
input x426;
input x427;
input x428;
input x429;
input x430;
input x431;
input x432;
input x433;
input x434;
input x435;
input x436;
input x437;
input x438;
input x439;
input x440;
input x441;
input x442;
input x443;
input x444;
input x445;
input x446;
input x447;
input x448;
input x449;
input x450;
input x451;
input x452;
input x453;
input x454;
input x455;
input x456;
input x457;
input x458;
input x459;
input x460;
input x461;
input x462;
input x463;
input x464;
input x465;
input x466;
input x467;
input x468;
input x469;
input x470;
input x471;
input x472;
input x473;
input x474;
input x475;
input x476;
input x477;
input x478;
input x479;
input x480;
input x481;
input x482;
input x483;
input x484;
input x485;
input x486;
input x487;
input x488;
input x489;
input x490;
input x491;
input x492;
input x493;
input x494;
input x495;
input x496;
input x497;
input x498;
input x499;
input x500;
input x501;
input x502;
input x503;
input x504;
input x505;
input x506;
input x507;
input x508;
input x509;
input x510;
input x511;
input x512;
input x513;
input x514;
input x515;
input x516;
input x517;
input x518;
input x519;
input x520;
input x521;
input x522;
input x523;
input x524;
input x525;
input x526;
input x527;
input x528;
input x529;
input x530;
input x531;
input x532;
input x533;
input x534;
input x535;
input x536;
input x537;
input x538;
input x539;
input x540;
input x541;
input x542;
input x543;
input x544;
input x545;
input x546;
input x547;
input x548;
input x549;
input x550;
input x551;
input x552;
input x553;
input x554;
input x555;
input x556;
input x557;
input x558;
input x559;
input x560;
input x561;
input x562;
input x563;
input x564;
input x565;
input x566;
input x567;
input x568;
input x569;
input x570;
input x571;
input x572;
input x573;
input x574;
input x575;
input x576;
input x577;
input x578;
input x579;
input x580;
input x581;
input x582;
input x583;
input x584;
input x585;
input x586;
input x587;
input x588;
input x589;
input x590;
input x591;
input x592;
input x593;
input x594;
input x595;
input x596;
input x597;
input x598;
input x599;
input x600;
input x601;
input x602;
input x603;
input x604;
input x605;
input x606;
input x607;
input x608;
input x609;
input x610;
input x611;
input x612;
input x613;
input x614;
input x615;
input x616;
input x617;
input x618;
input x619;
input x620;
input x621;
input x622;
input x623;
input x624;
input x625;
input x626;
input x627;
input x628;
input x629;
input x630;
input x631;
input x632;
input x633;
input x634;
input x635;
input x636;
input x637;
input x638;
input x639;
input x640;
input x641;
input x642;
input x643;
input x644;
input x645;
input x646;
input x647;
input x648;
input x649;
input x650;
input x651;
input x652;
input x653;
input x654;
input x655;
input x656;
input x657;
input x658;
input x659;
input x660;
input x661;
input x662;
input x663;
input x664;
input x665;
input x666;
input x667;
input x668;
input x669;
input x670;
input x671;
input x672;
input x673;
input x674;
input x675;
input x676;
input x677;
input x678;
input x679;
input x680;
input x681;
input x682;
input x683;
input x684;
input x685;
input x686;
input x687;
input x688;
input x689;
input x690;
input x691;
input x692;
input x693;
input x694;
input x695;
input x696;
input x697;
input x698;
input x699;
input x700;
input x701;
input x702;
input x703;
input x704;
input x705;
input x706;
input x707;
input x708;
input x709;
input x710;
input x711;
input x712;
input x713;
input x714;
input x715;
input x716;
input x717;
input x718;
input x719;
input x720;
input x721;
input x722;
input x723;
input x724;
input x725;
input x726;
input x727;
input x728;
input x729;
input x730;
input x731;
input x732;
input x733;
input x734;
input x735;
input x736;
input x737;
input x738;
input x739;
input x740;
input x741;
input x742;
input x743;
input x744;
input x745;
input x746;
input x747;
input x748;
input x749;
input x750;
input x751;
input x752;
input x753;
input x754;
input x755;
input x756;
input x757;
input x758;
input x759;
input x760;
input x761;
input x762;
input x763;
input x764;
input x765;
input x766;
input x767;
input x768;
input x769;
input x770;
input x771;
input x772;
input x773;
input x774;
input x775;
input x776;
input x777;
input x778;
input x779;
input x780;
input x781;
input x782;
input x783;
output c6228;
output c8114;
output c9123;
output c3431;
output c674;
output c9436;
output c6318;
output c172;
output c157;
output c2126;
output c6291;
output c7475;
output c8363;
output c5348;
output c051;
output c424;
output c2187;
output c9358;
output c024;
output c4461;
output c1333;
output c6321;
output c2165;
output c8187;
output c4463;
output c6458;
output c969;
output c1308;
output c6420;
output c9206;
output c4363;
output c918;
output c951;
output c6392;
output c2433;
output c4172;
output c8286;
output c3417;
output c5254;
output c8238;
output c1412;
output c7152;
output c9284;
output c9142;
output c03;
output c6255;
output c567;
output c416;
output c7125;
output c8369;
output c6441;
output c135;
output c6288;
output c9312;
output c7315;
output c7436;
output c2198;
output c111;
output c6247;
output c7381;
output c841;
output c0319;
output c2216;
output c3479;
output c0264;
output c0110;
output c7167;
output c1352;
output c7404;
output c6365;
output c22;
output c536;
output c367;
output c2342;
output c4267;
output c1248;
output c3241;
output c4350;
output c7428;
output c626;
output c5255;
output c3190;
output c537;
output c2145;
output c1360;
output c445;
output c4187;
output c8395;
output c2100;
output c6476;
output c3134;
output c0442;
output c0439;
output c9242;
output c0343;
output c285;
output c0123;
output c1294;
output c3358;
output c0453;
output c9119;
output c5207;
output c1397;
output c1109;
output c4312;
output c5405;
output c3310;
output c8380;
output c9239;
output c9336;
output c3274;
output c4427;
output c358;
output c947;
output c9191;
output c1379;
output c8139;
output c30;
output c4315;
output c414;
output c2351;
output c0262;
output c3164;
output c2338;
output c3132;
output c535;
output c062;
output c7180;
output c1256;
output c5171;
output c228;
output c4467;
output c148;
output c3322;
output c2281;
output c5239;
output c943;
output c133;
output c9155;
output c648;
output c2271;
output c8436;
output c7322;
output c8368;
output c1453;
output c8110;
output c5116;
output c9297;
output c2352;
output c7246;
output c4443;
output c780;
output c691;
output c3306;
output c3418;
output c295;
output c547;
output c2209;
output c2465;
output c8163;
output c8165;
output c9461;
output c3364;
output c1290;
output c9216;
output c6316;
output c1457;
output c5371;
output c8340;
output c9379;
output c5323;
output c5260;
output c0303;
output c240;
output c5174;
output c1420;
output c6433;
output c6367;
output c259;
output c7107;
output c188;
output c1262;
output c0426;
output c2200;
output c5480;
output c329;
output c9271;
output c5368;
output c4382;
output c5274;
output c4298;
output c631;
output c0183;
output c8329;
output c3297;
output c6322;
output c6175;
output c8381;
output c1204;
output c4481;
output c752;
output c066;
output c0108;
output c5411;
output c2252;
output c5271;
output c8401;
output c3143;
output c7266;
output c1179;
output c7429;
output c3126;
output c5242;
output c1380;
output c0178;
output c390;
output c9421;
output c3184;
output c3395;
output c7488;
output c2392;
output c1325;
output c4227;
output c1462;
output c646;
output c2372;
output c3121;
output c9114;
output c4432;
output c4135;
output c8331;
output c2334;
output c6274;
output c8258;
output c3230;
output c6370;
output c666;
output c4440;
output c2234;
output c874;
output c0357;
output c7396;
output c9225;
output c4434;
output c5182;
output c8151;
output c7358;
output c848;
output c7483;
output c2163;
output c8426;
output c0396;
output c6187;
output c7317;
output c5165;
output c1465;
output c2319;
output c1267;
output c6300;
output c569;
output c7446;
output c3346;
output c365;
output c359;
output c8105;
output c9230;
output c5412;
output c7355;
output c0417;
output c015;
output c2405;
output c1146;
output c326;
output c6140;
output c9320;
output c3260;
output c5393;
output c084;
output c0128;
output c12;
output c5406;
output c0189;
output c3379;
output c3137;
output c1466;
output c7173;
output c7103;
output c3426;
output c925;
output c8257;
output c0400;
output c2460;
output c5158;
output c0182;
output c0252;
output c562;
output c6403;
output c4479;
output c6345;
output c47;
output c039;
output c2263;
output c6385;
output c381;
output c4324;
output c190;
output c4356;
output c5436;
output c4445;
output c7166;
output c050;
output c3324;
output c891;
output c5431;
output c1284;
output c132;
output c1121;
output c0360;
output c1201;
output c8325;
output c8263;
output c592;
output c7369;
output c7200;
output c1437;
output c8371;
output c1326;
output c2233;
output c9167;
output c3340;
output c7362;
output c988;
output c1111;
output c297;
output c1175;
output c7150;
output c0298;
output c3456;
output c3138;
output c4352;
output c7468;
output c9373;
output c5367;
output c2361;
output c6327;
output c5347;
output c2404;
output c782;
output c8319;
output c2196;
output c3213;
output c6425;
output c0118;
output c1266;
output c6220;
output c4196;
output c5460;
output c6334;
output c9353;
output c5261;
output c0171;
output c1277;
output c2118;
output c0406;
output c5493;
output c5389;
output c0373;
output c14;
output c4132;
output c177;
output c893;
output c9209;
output c5491;
output c3487;
output c450;
output c1415;
output c1482;
output c4449;
output c6237;
output c5353;
output c191;
output c4412;
output c3217;
output c3148;
output c1435;
output c0331;
output c2348;
output c4168;
output c073;
output c8265;
output c252;
output c4188;
output c4270;
output c1142;
output c4224;
output c3160;
output c8162;
output c4292;
output c3116;
output c7473;
output c735;
output c2140;
output c5358;
output c9344;
output c2332;
output c9127;
output c76;
output c028;
output c8420;
output c8327;
output c3224;
output c0236;
output c9112;
output c9359;
output c210;
output c4208;
output c1239;
output c0391;
output c2250;
output c528;
output c2467;
output c4134;
output c9309;
output c2146;
output c2344;
output c8310;
output c2422;
output c6102;
output c6472;
output c8422;
output c612;
output c3437;
output c0358;
output c3170;
output c2304;
output c1344;
output c2103;
output c8185;
output c9116;
output c8357;
output c038;
output c8311;
output c4212;
output c0254;
output c5426;
output c3333;
output c5238;
output c0272;
output c4415;
output c4404;
output c8355;
output c7357;
output c5144;
output c3287;
output c5219;
output c235;
output c491;
output c6457;
output c025;
output c3331;
output c0293;
output c7250;
output c0488;
output c0367;
output c7484;
output c5146;
output c2490;
output c7235;
output c2377;
output c0234;
output c1215;
output c398;
output c1414;
output c5243;
output c8130;
output c7347;
output c7393;
output c7228;
output c964;
output c788;
output c7496;
output c5230;
output c164;
output c6397;
output c2246;
output c5485;
output c1143;
output c0295;
output c7330;
output c8469;
output c1405;
output c2186;
output c7284;
output c1449;
output c6325;
output c751;
output c6363;
output c5232;
output c5283;
output c0283;
output c7101;
output c5249;
output c747;
output c1145;
output c7236;
output c2458;
output c90;
output c885;
output c3171;
output c0190;
output c2331;
output c463;
output c534;
output c7132;
output c7297;
output c3149;
output c733;
output c711;
output c7426;
output c9453;
output c0458;
output c2437;
output c6234;
output c6266;
output c665;
output c1321;
output c4157;
output c57;
output c6418;
output c4381;
output c2474;
output c8296;
output c00;
output c4297;
output c781;
output c8176;
output c9362;
output c5355;
output c1172;
output c8283;
output c645;
output c8148;
output c0380;
output c2475;
output c0144;
output c7176;
output c9177;
output c336;
output c7239;
output c1167;
output c0411;
output c4102;
output c8215;
output c1370;
output c3470;
output c4181;
output c8440;
output c2341;
output c2318;
output c0258;
output c862;
output c5161;
output c3493;
output c27;
output c8378;
output c6486;
output c7440;
output c4317;
output c9169;
output c1406;
output c7366;
output c5397;
output c762;
output c6395;
output c6324;
output c911;
output c5398;
output c4314;
output c0223;
output c7211;
output c7187;
output c54;
output c8222;
output c1301;
output c0481;
output c8279;
output c0227;
output c50;
output c2273;
output c4328;
output c8159;
output c7192;
output c6263;
output c9348;
output c0199;
output c313;
output c2360;
output c3187;
output c5320;
output c9364;
output c5175;
output c963;
output c1305;
output c5432;
output c659;
output c4383;
output c8122;
output c0433;
output c1122;
output c5157;
output c6173;
output c1178;
output c984;
output c4425;
output c0263;
output c0151;
output c3485;
output c8342;
output c7331;
output c5270;
output c0122;
output c3328;
output c9276;
output c896;
output c4289;
output c5424;
output c790;
output c2430;
output c5107;
output c0469;
output c2413;
output c1350;
output c727;
output c1432;
output c3375;
output c7225;
output c4178;
output c0356;
output c967;
output c7238;
output c3202;
output c5269;
output c1258;
output c0274;
output c8276;
output c1323;
output c5288;
output c6352;
output c7466;
output c110;
output c7204;
output c1190;
output c0461;
output c4263;
output c1400;
output c6109;
output c9408;
output c4291;
output c5361;
output c5176;
output c5251;
output c9458;
output c8180;
output c7439;
output c5391;
output c493;
output c2419;
output c5478;
output c9473;
output c9341;
output c6482;
output c3407;
output c9361;
output c176;
output c7257;
output c7181;
output c7227;
output c6146;
output c2115;
output c255;
output c069;
output c0459;
output c6259;
output c3409;
output c865;
output c8367;
output c0164;
output c1383;
output c6319;
output c3102;
output c6139;
output c9143;
output c8494;
output c7442;
output c7435;
output c7291;
output c9433;
output c7373;
output c87;
output c9219;
output c2171;
output c2229;
output c778;
output c8460;
output c3434;
output c2427;
output c3354;
output c5258;
output c5287;
output c5308;
output c1234;
output c7155;
output c312;
output c1273;
output c2386;
output c4392;
output c7114;
output c8214;
output c6271;
output c1297;
output c9220;
output c2157;
output c2347;
output c3139;
output c554;
output c3243;
output c4269;
output c6353;
output c5240;
output c7280;
output c1320;
output c4332;
output c1300;
output c3350;
output c4290;
output c1282;
output c6130;
output c2366;
output c513;
output c9185;
output c5435;
output c2446;
output c525;
output c4388;
output c4407;
output c6496;
output c6465;
output c728;
output c0120;
output c6177;
output c0176;
output c597;
output c8271;
output c6176;
output c4229;
output c1193;
output c8421;
output c677;
output c3317;
output c9371;
output c0181;
output c9252;
output c431;
output c8470;
output c5164;
output c9111;
output c8345;
output c2168;
output c7432;
output c0434;
output c1477;
output c5311;
output c7149;
output c0107;
output c3229;
output c7441;
output c490;
output c6375;
output c7191;
output c8284;
output c0261;
output c0139;
output c638;
output c5233;
output c5417;
output c9422;
output c9391;
output c343;
output c791;
output c912;
output c7351;
output c9497;
output c4361;
output c640;
output c653;
output c4154;
output c3144;
output c7224;
output c1495;
output c8415;
output c5450;
output c2328;
output c6180;
output c8307;
output c262;
output c974;
output c121;
output c8416;
output c7161;
output c089;
output c3329;
output c4372;
output c8193;
output c340;
output c9486;
output c0211;
output c3211;
output c9303;
output c1137;
output c1185;
output c5148;
output c0399;
output c1361;
output c8356;
output c1468;
output c7361;
output c012;
output c2104;
output c8493;
output c7146;
output c0114;
output c4186;
output c366;
output c5145;
output c0218;
output c7324;
output c9465;
output c3394;
output c1268;
output c3474;
output c377;
output c0260;
output c4307;
output c3460;
output c519;
output c1159;
output c6158;
output c0106;
output c8383;
output c3469;
output c9235;
output c2112;
output c0214;
output c7202;
output c8475;
output c3279;
output c474;
output c729;
output c5322;
output c3408;
output c681;
output c1304;
output c5252;
output c6195;
output c3422;
output c4180;
output c1328;
output c591;
output c775;
output c35;
output c38;
output c4226;
output c9467;
output c9313;
output c0289;
output c8155;
output c3196;
output c6454;
output c839;
output c3200;
output c7163;
output c6153;
output c2367;
output c628;
output c9492;
output c8496;
output c4129;
output c80;
output c9176;
output c0207;
output c4391;
output c7140;
output c98;
output c3197;
output c2393;
output c4330;
output c5313;
output c7118;
output c2375;
output c2335;
output c6161;
output c9468;
output c2486;
output c279;
output c4145;
output c5130;
output c4451;
output c7417;
output c8244;
output c6396;
output c480;
output c1396;
output c5185;
output c6432;
output c4191;
output c45;
output c9446;
output c6142;
output c7186;
output c2236;
output c2218;
output c174;
output c5463;
output c5102;
output c20;
output c139;
output c0273;
output c9419;
output c2248;
output c8133;
output c6215;
output c8365;
output c1483;
output c7332;
output c9207;
output c0354;
output c4389;
output c4149;
output c8247;
output c134;
output c4378;
output c9187;
output c8134;
output c8390;
output c6218;
output c0378;
output c058;
output c1395;
output c6438;
output c2109;
output c4301;
output c0221;
output c0310;
output c6276;
output c7264;
output c196;
output c4397;
output c7216;
output c085;
output c3466;
output c9447;
output c6204;
output c819;
output c5290;
output c3244;
output c6303;
output c8439;
output c5235;
output c231;
output c2454;
output c063;
output c9460;
output c69;
output c1441;
output c161;
output c0268;
output c7499;
output c2150;
output c4336;
output c3482;
output c1331;
output c3406;
output c2483;
output c1182;
output c064;
output c1136;
output c6193;
output c2137;
output c027;
output c7198;
output c5213;
output c1155;
output c8111;
output c1281;
output c6222;
output c4344;
output c189;
output c2279;
output c8321;
output c4216;
output c7427;
output c9456;
output c5420;
output c7407;
output c5442;
output c1339;
output c0165;
output c1251;
output c6413;
output c9369;
output c1398;
output c5132;
output c2285;
output c394;
output c5197;
output c9200;
output c0168;
output c3351;
output c5481;
output c876;
output c292;
output c0256;
output c0312;
output c155;
output c0194;
output c2325;
output c5327;
output c5345;
output c3427;
output c3383;
output c1214;
output c01;
output c6243;
output c1438;
output c266;
output c6152;
output c393;
output c0192;
output c8154;
output c138;
output c7207;
output c7269;
output c2440;
output c9132;
output c6261;
output c1430;
output c1452;
output c1474;
output c7217;
output c8414;
output c5392;
output c9180;
output c153;
output c9316;
output c0487;
output c7212;
output c4244;
output c5256;
output c9228;
output c5241;
output c1424;
output c2388;
output c8211;
output c6148;
output c5275;
output c4170;
output c2181;
output c0389;
output c9168;
output c1358;
output c5246;
output c816;
output c047;
output c2491;
output c6497;
output c6210;
output c1357;
output c9481;
output c3494;
output c6401;
output c6114;
output c2134;
output c5237;
output c5324;
output c8431;
output c1225;
output c1332;
output c2212;
output c682;
output c8339;
output c1366;
output c4474;
output c8233;
output c686;
output c3262;
output c5369;
output c6308;
output c8452;
output c5133;
output c4232;
output c5396;
output c371;
output c6168;
output c4167;
output c9471;
output c683;
output c418;
output c6233;
output c5121;
output c581;
output c0270;
output c0322;
output c3313;
output c6178;
output c748;
output c5160;
output c2166;
output c647;
output c3123;
output c8349;
output c2380;
output c4371;
output c1206;
output c5122;
output c2376;
output c668;
output c7286;
output c6483;
output c3203;
output c9406;
output c5386;
output c9149;
output c1154;
output c4496;
output c6329;
output c2323;
output c737;
output c3491;
output c9282;
output c9337;
output c472;
output c6108;
output c9135;
output c994;
output c0416;
output c5452;
output c9179;
output c89;
output c8101;
output c6309;
output c8150;
output c6201;
output c042;
output c3468;
output c1244;
output c3207;
output c1355;
output c0478;
output c0425;
output c215;
output c4194;
output c933;
output c6154;
output c0381;
output c3135;
output c485;
output c6199;
output c7372;
output c6267;
output c0141;
output c7327;
output c126;
output c753;
output c8113;
output c2495;
output c417;
output c670;
output c234;
output c041;
output c5143;
output c92;
output c5315;
output c2395;
output c616;
output c9255;
output c3114;
output c4464;
output c6424;
output c4123;
output c3179;
output c044;
output c3236;
output c5490;
output c5217;
output c5404;
output c8246;
output c3248;
output c7348;
output c3338;
output c8240;
output c3352;
output c774;
output c2107;
output c3376;
output c946;
output c0259;
output c181;
output c8181;
output c6145;
output c8109;
output c1334;
output c2410;
output c5376;
output c9372;
output c0210;
output c4450;
output c8225;
output c4318;
output c898;
output c0448;
output c8387;
output c2400;
output c9248;
output c1115;
output c6227;
output c5263;
output c4251;
output c08;
output c7354;
output c7283;
output c9233;
output c1388;
output c9263;
output c446;
output c8145;
output c2228;
output c1302;
output c3188;
output c0347;
output c2265;
output c3186;
output c8131;
output c7177;
output c8256;
output c0456;
output c934;
output c9305;
output c043;
output c4271;
output c6171;
output c3218;
output c553;
output c5193;
output c6211;
output c5438;
output c49;
output c0232;
output c9218;
output c8285;
output c071;
output c694;
output c1410;
output c2421;
output c4437;
output c0444;
output c1375;
output c254;
output c9154;
output c6405;
output c9108;
output c6339;
output c3357;
output c0251;
output c7319;
output c0492;
output c8312;
output c319;
output c3122;
output c8338;
output c9365;
output c9479;
output c1228;
output c8213;
output c6293;
output c2457;
output c5477;
output c3258;
output c3393;
output c8481;
output c777;
output c9420;
output c9294;
output c5299;
output c3182;
output c9274;
output c1351;
output c9444;
output c769;
output c0484;
output c8178;
output c4494;
output c7292;
output c927;
output c6310;
output c538;
output c928;
output c3100;
output c8461;
output c741;
output c6400;
output c0250;
output c9355;
output c1336;
output c8202;
output c4230;
output c835;
output c3488;
output c2468;
output c3286;
output c3289;
output c1177;
output c937;
output c9298;
output c920;
output c7371;
output c2283;
output c166;
output c561;
output c1429;
output c278;
output c3146;
output c3459;
output c0285;
output c2183;
output c5196;
output c0404;
output c6383;
output c2277;
output c5318;
output c8495;
output c2149;
output c4177;
output c8297;
output c2292;
output c7148;
output c2333;
output c2498;
output c6402;
output c5425;
output c033;
output c4228;
output c0480;
output c1205;
output c9351;
output c5441;
output c6443;
output c5209;
output c9251;
output c4219;
output c7356;
output c272;
output c056;
output c5224;
output c1263;
output c017;
output c7388;
output c6282;
output c0153;
output c5153;
output c5461;
output c460;
output c5335;
output c936;
output c2471;
output c9134;
output c2299;
output c3360;
output c4320;
output c4109;
output c2113;
output c4438;
output c0422;
output c588;
output c3391;
output c3454;
output c6311;
output c6150;
output c642;
output c3413;
output c9360;
output c0173;
output c2257;
output c3150;
output c8189;
output c4125;
output c8372;
output c7449;
output c0339;
output c032;
output c4390;
output c281;
output c3298;
output c2431;
output c4242;
output c0371;
output c9477;
output c1106;
output c2215;
output c3129;
output c6284;
output c4343;
output c3425;
output c4419;
output c9430;
output c9171;
output c5325;
output c0238;
output c7410;
output c761;
output c1425;
output c529;
output c6349;
output c4128;
output c081;
output c29;
output c4176;
output c1488;
output c5104;
output c7433;
output c7376;
output c1257;
output c1158;
output c1218;
output c678;
output c9221;
output c6164;
output c8206;
output c7234;
output c320;
output c8303;
output c3173;
output c9349;
output c0419;
output c9319;
output c9162;
output c140;
output c6226;
output c3455;
output c9366;
output c5380;
output c7142;
output c4274;
output c2456;
output c7143;
output c734;
output c074;
output c9476;
output c5181;
output c4306;
output c5112;
output c4367;
output c0209;
output c6240;
output c4452;
output c5416;
output c6273;
output c5282;
output c7313;
output c8393;
output c6238;
output c1472;
output c61;
output c9300;
output c796;
output c1260;
output c2116;
output c7480;
output c8308;
output c3496;
output c973;
output c0338;
output c4160;
output c0241;
output c9270;
output c8465;
output c83;
output c6229;
output c997;
output c4262;
output c5317;
output c2477;
output c9399;
output c9450;
output c323;
output c5497;
output c3189;
output c1356;
output c8468;
output c5403;
output c91;
output c020;
output c4446;
output c6245;
output c3301;
output c5365;
output c1120;
output c1129;
output c3314;
output c6197;
output c6250;
output c0477;
output c9189;
output c1411;
output c7392;
output c1247;
output c3118;
output c4385;
output c742;
output c5401;
output c82;
output c7124;
output c9104;
output c1431;
output c325;
output c6407;
output c1377;
output c2173;
output c7308;
output c9402;
output c5387;
output c8216;
output c6217;
output c7231;
output c8212;
output c4200;
output c1107;
output c1157;
output c7300;
output c1455;
output c116;
output c9292;
output c437;
output c6398;
output c4152;
output c3450;
output c2379;
output c4490;
output c8483;
output c853;
output c1187;
output c1135;
output c4447;
output c9435;
output c4468;
output c855;
output c1209;
output c3294;
output c3227;
output c3133;
output c4342;
output c9172;
output c2359;
output c837;
output c7121;
output c076;
output c3337;
output c982;
output c0301;
output c861;
output c4300;
output c128;
output c4264;
output c7398;
output c0271;
output c2220;
output c342;
output c4201;
output c975;
output c9334;
output c459;
output c2309;
output c3449;
output c3288;
output c7482;
output c7312;
output c8434;
output c3446;
output c016;
output c3204;
output c7119;
output c2424;
output c5225;
output c8277;
output c337;
output c0111;
output c671;
output c866;
output c840;
output c0413;
output c4250;
output c335;
output c9449;
output c8245;
output c8300;
output c3467;
output c990;
output c6358;
output c7271;
output c0397;
output c4472;
output c2462;
output c5203;
output c061;
output c0246;
output c9363;
output c7259;
output c643;
output c1163;
output c7465;
output c4115;
output c870;
output c8249;
output c034;
output c8457;
output c249;
output c4430;
output c1387;
output c486;
output c9105;
output c379;
output c3208;
output c8294;
output c8264;
output c6434;
output c5278;
output c4210;
output c0196;
output c8104;
output c1443;
output c673;
output c1108;
output c6181;
output c3119;
output c2358;
output c851;
output c2194;
output c380;
output c9266;
output c5150;
output c3445;
output c976;
output c4414;
output c3442;
output c2355;
output c4294;
output c883;
output c0309;
output c355;
output c9144;
output c2232;
output c3181;
output c0208;
output c433;
output c7287;
output c7136;
output c5247;
output c881;
output c0318;
output c0320;
output c0133;
output c1133;
output c622;
output c4153;
output c4100;
output c6467;
output c3273;
output c4101;
output c784;
output c4235;
output c4260;
output c8194;
output c362;
output c1296;
output c6242;
output c4222;
output c4423;
output c8118;
output c699;
output c4357;
output c2364;
output c0226;
output c1403;
output c6131;
output c7333;
output c013;
output c1364;
output c593;
output c797;
output c2432;
output c4364;
output c36;
output c744;
output c2385;
output c5201;
output c9434;
output c6491;
output c842;
output c9247;
output c8322;
output c7273;
output c5192;
output c7249;
output c0186;
output c51;
output c579;
output c8313;
output c6448;
output c3414;
output c4454;
output c059;
output c28;
output c299;
output c4249;
output c9464;
output c724;
output c4202;
output c6409;
output c710;
output c8444;
output c3219;
output c257;
output c5245;
output c4106;
output c9498;
output c5292;
output c0436;
output c6290;
output c0355;
output c0286;
output c1197;
output c481;
output c7405;
output c6464;
output c24;
output c6384;
output c9438;
output c8455;
output c4341;
output c949;
output c3464;
output c026;
output c2139;
output c6185;
output c9193;
output c0311;
output c0281;
output c7141;
output c2230;
output c9317;
output c8441;
output c7452;
output c772;
output c8438;
output c726;
output c167;
output c9385;
output c1434;
output c7457;
output c018;
output c4253;
output c8499;
output c63;
output c091;
output c521;
output c324;
output c9454;
output c3268;
output c8250;
output c0342;
output c1354;
output c7203;
output c6213;
output c0253;
output c5453;
output c766;
output c387;
output c8100;
output c1433;
output c598;
output c9152;
output c1275;
output c3107;
output c7215;
output c2258;
output c4205;
output c1419;
output c7294;
output c466;
output c9389;
output c6184;
output c6307;
output c8405;
output c3278;
output c542;
output c4238;
output c7251;
output c3371;
output c1480;
output c6147;
output c5366;
output c5340;
output c5162;
output c5421;
output c9326;
output c9472;
output c9140;
output c7343;
output c9126;
output c0465;
output c3277;
output c269;
output c7290;
output c2175;
output c6451;
output c9368;
output c4359;
output c5306;
output c05;
output c4442;
output c080;
output c6393;
output c635;
output c4127;
output c4141;
output c3257;
output c9384;
output c6332;
output c6183;
output c5456;
output c867;
output c487;
output c9401;
output c4116;
output c6380;
output c6455;
output c5328;
output c2420;
output c4418;
output c6492;
output c9329;
output c1186;
output c8409;
output c467;
output c5468;
output c1324;
output c684;
output c1211;
output c7174;
output c625;
output c7178;
output c5291;
output c0288;
output c8209;
output c2156;
output c7316;
output c779;
output c0490;
output c552;
output c0160;
output c494;
output c2288;
output c6326;
output c2287;
output c0294;
output c7477;
output c220;
output c5152;
output c9459;
output c3388;
output c0155;
output c5128;
output c88;
output c1440;
output c1110;
output c159;
output c341;
output c9416;
output c8182;
output c9211;
output c0138;
output c5140;
output c0179;
output c2193;
output c6360;
output c8124;
output c3315;
output c0102;
output c224;
output c4111;
output c0430;
output c6337;
output c6192;
output c9466;
output c0146;
output c3372;
output c545;
output c2448;
output c945;
output c7419;
output c75;
output c7494;
output c55;
output c1184;
output c8161;
output c7345;
output c2415;
output c3478;
output c8289;
output c9295;
output c2345;
output c7460;
output c0486;
output c9146;
output c8464;
output c9310;
output c0170;
output c2481;
output c617;
output c5314;
output c9491;
output c9345;
output c2214;
output c6470;
output c7123;
output c1224;
output c8183;
output c6423;
output c833;
output c8323;
output c5208;
output c6138;
output c64;
output c1363;
output c1487;
output c2151;
output c5331;
output c7253;
output c0121;
output c3448;
output c8385;
output c1390;
output c764;
output c8391;
output c584;
output c844;
output c627;
output c5429;
output c798;
output c356;
output c636;
output c875;
output c4273;
output c6125;
output c9396;
output c85;
output c5142;
output c4406;
output c2106;
output c169;
output c0224;
output c3327;
output c1313;
output c9136;
output c9288;
output c2174;
output c773;
output c3498;
output c9262;
output c610;
output c7413;
output c0427;
output c1232;
output c6372;
output c8230;
output c2199;
output c3240;
output c8449;
output c5105;
output c2164;
output c9121;
output c634;
output c6236;
output c7382;
output c4497;
output c8166;
output c3339;
output c1311;
output c2224;
output c2423;
output c2256;
output c8291;
output c0388;
output c2301;
output c892;
output c4422;
output c8482;
output c094;
output c2136;
output c7350;
output c745;
output c2321;
output c3403;
output c4174;
output c451;
output c1348;
output c1295;
output c8208;
output c090;
output c1494;
output c2203;
output c369;
output c859;
output c6331;
output c2225;
output c274;
output c125;
output c5344;
output c4433;
output c4183;
output c971;
output c060;
output c9208;
output c4351;
output c6453;
output c6468;
output c1243;
output c5336;
output c4482;
output c2221;
output c1322;
output c5390;
output c311;
output c9101;
output c6422;
output c7138;
output c8266;
output c8471;
output c163;
output c3433;
output c2414;
output c623;
output c2298;
output c07;
output c2213;
output c0491;
output c3225;
output c6298;
output c6350;
output c749;
output c498;
output c9400;
output c1342;
output c2195;
output c9267;
output c4223;
output c9124;
output c7258;
output c669;
output c9327;
output c1490;
output c4248;
output c4444;
output c5149;
output c2390;
output c1194;
output c1309;
output c482;
output c3400;
output c8108;
output c6117;
output c6335;
output c716;
output c2231;
output c0368;
output c576;
output c4254;
output c5114;
output c9426;
output c6182;
output c154;
output c821;
output c1303;
output c9286;
output c655;
output c9299;
output c6160;
output c2499;
output c792;
output c84;
output c7193;
output c0372;
output c1404;
output c4287;
output c7171;
output c0150;
output c0277;
output c3261;
output c5302;
output c7218;
output c965;
output c8195;
output c2311;
output c695;
output c8253;
output c9229;
output c149;
output c0324;
output c0316;
output c1338;
output c3444;
output c1134;
output c5451;
output c0455;
output c4466;
output c495;
output c1448;
output c4215;
output c8190;
output c9291;
output c873;
output c7377;
output c2397;
output c1207;
output c8232;
output c0359;
output c4347;
output c1255;
output c578;
output c675;
output c2177;
output c2492;
output c9390;
output c1409;
output c6368;
output c3155;
output c7285;
output c4398;
output c8354;
output c310;
output c232;
output c688;
output c1407;
output c7311;
output c1235;
output c8462;
output c3152;
output c8324;
output c443;
output c2312;
output c2238;
output c9490;
output c4150;
output c5499;
output c6436;
output c7260;
output c1114;
output c8374;
output c4151;
output c568;
output c6260;
output c7220;
output c8361;
output c8419;
output c144;
output c680;
output c395;
output c2317;
output c5212;
output c5188;
output c1213;
output c7490;
output c375;
output c3304;
output c6444;
output c7303;
output c0112;
output c0364;
output c5298;
output c8358;
output c7233;
output c6404;
output c7370;
output c541;
output c6264;
output c1233;
output c5297;
output c3463;
output c233;
output c9393;
output c512;
output c7455;
output c321;
output c9495;
output c551;
output c8411;
output c421;
output c7214;
output c5400;
output c813;
output c6437;
output c2494;
output c2396;
output c9383;
output c5250;
output c2211;
output c8293;
output c271;
output c879;
output c353;
output c1270;
output c6488;
output c2455;
output c9480;
output c3252;
output c1253;
output c3141;
output c721;
output c399;
output c8382;
output c6354;
output c651;
output c2223;
output c7219;
output c0497;
output c4107;
output c4354;
output c2293;
output c0228;
output c317;
output c2417;
output c9437;
output c4217;
output c8337;
output c2429;
output c6330;
output c882;
output c1471;
output c7338;
output c1436;
output c1470;
output c057;
output c488;
output c0229;
output c7244;
output c5115;
output c5309;
output c373;
output c9203;
output c1408;
output c5177;
output c0161;
output c894;
output c0332;
output c9272;
output c0105;
output c4221;
output c3125;
output c983;
output c2276;
output c924;
output c10;
output c3157;
output c4280;
output c282;
output c3348;
output c62;
output c6257;
output c1450;
output c2408;
output c9264;
output c978;
output c010;
output c2192;
output c253;
output c1164;
output c2435;
output c7352;
output c198;
output c4182;
output c621;
output c550;
output c7461;
output c9215;
output c0222;
output c1489;
output c3282;
output c5356;
output c229;
output c0370;
output c6151;
output c0405;
output c088;
output c6373;
output c7272;
output c5330;
output c2451;
output c3386;
output c60;
output c5119;
output c4345;
output c152;
output c7448;
output c1393;
output c0424;
output c5155;
output c1269;
output c6133;
output c3457;
output c065;
output c9380;
output c6427;
output c8174;
output c5190;
output c3145;
output c868;
output c1138;
output c316;
output c383;
output c5284;
output c6129;
output c558;
output c6299;
output c4105;
output c419;
output c5377;
output c7487;
output c1166;
output c7105;
output c8295;
output c1212;
output c150;
output c429;
output c2470;
output c9201;
output c1337;
output c6202;
output c6254;
output c663;
output c123;
output c595;
output c3490;
output c817;
output c3336;
output c2204;
output c2154;
output c4218;
output c2217;
output c757;
output c1285;
output c4448;
output c6328;
output c594;
output c9170;
output c7464;
output c7438;
output c9487;
output c0390;
output c4321;
output c5312;
output c2227;
output c5489;
output c2268;
output c428;
output c4118;
output c845;
output c2152;
output c7275;
output c5388;
output c4487;
output c298;
output c2306;
output c2120;
output c8201;
output c6265;
output c1287;
output c836;
output c0245;
output c014;
output c7342;
output c5257;
output c8418;
output c4256;
output c3345;
output c880;
output c0374;
output c1230;
output c4485;
output c9424;
output c42;
output c171;
output c9387;
output c0284;
output c331;
output c7172;
output c4272;
output c6301;
output c6498;
output c5352;
output c1189;
output c4376;
output c856;
output c265;
output c7380;
output c4309;
output c8404;
output c8445;
output c5455;
output c9181;
output c9249;
output c9174;
output c5221;
output c0149;
output c1341;
output c5462;
output c9130;
output c6388;
output c8343;
output c368;
output c0197;
output c6110;
output c96;
output c4455;
output c1418;
output c6305;
output c5191;
output c7276;
output c0350;
output c3390;
output c4386;
output c425;
output c570;
output c5482;
output c114;
output c226;
output c193;
output c583;
output c0414;
output c6246;
output c0363;
output c2439;
output c6118;
output c6351;
output c812;
output c5458;
output c040;
output c8466;
output c3447;
output c0129;
output c0101;
output c5214;
output c3458;
output c8346;
output c0115;
output c3384;
output c9175;
output c2478;
output c2484;
output c6382;
output c6297;
output c1156;
output c6295;
output c2260;
output c79;
output c864;
output c9241;
output c0131;
output c7184;
output c9443;
output c7168;
output c6359;
output c8486;
output c7100;
output c2123;
output c396;
output c7254;
output c2340;
output c629;
output c0384;
output c1274;
output c2142;
output c330;
output c9245;
output c8158;
output c8477;
output c2450;
output c7113;
output c8226;
output c1279;
output c1219;
output c7395;
output c1132;
output c8373;
output c0117;
output c5343;
output c9137;
output c8453;
output c5100;
output c8443;
output c9273;
output c1381;
output c1496;
output c1116;
output c644;
output c16;
output c0454;
output c9159;
output c7188;
output c6107;
output c4304;
output c8137;
output c7112;
output c2329;
output c430;
output c1319;
output c4288;
output c7375;
output c8146;
output c8478;
output c5362;
output c5423;
output c9244;
output c9269;
output c4198;
output c7221;
output c243;
output c8184;
output c3486;
output c77;
output c3370;
output c1139;
output c2247;
output c4353;
output c3285;
output c7199;
output c7262;
output c8171;
output c6156;
output c284;
output c2438;
output c230;
output c2434;
output c6104;
output c566;
output c2416;
output c0449;
output c1130;
output c7296;
output c248;
output c3318;
output c5248;
output c793;
output c0483;
output c8447;
output c2270;
output c5117;
output c0437;
output c3497;
output c0315;
output c6466;
output c4410;
output c5360;
output c5349;
output c2180;
output c4373;
output c794;
output c1176;
output c5449;
output c713;
output c939;
output c2286;
output c3130;
output c9342;
output c3162;
output c0267;
output c8309;
output c4126;
output c0348;
output c818;
output c7344;
output c4133;
output c0201;
output c6341;
output c349;
output c3106;
output c9413;
output c8251;
output c7222;
output c7242;
output c3265;
output c453;
output c4234;
output c979;
output c3205;
output c1464;
output c7110;
output c3233;
output c820;
output c4394;
output c814;
output c574;
output c048;
output c5498;
output c5163;
output c944;
output c0498;
output c0475;
output c3451;
output c8410;
output c5409;
output c850;
output c7456;
output c4137;
output c5183;
output c6231;
output c5494;
output c4339;
output c977;
output c9165;
output c9439;
output c2473;
output c7368;
output c9107;
output c2373;
output c8364;
output c0452;
output c0466;
output c2464;
output c5151;
output c8129;
output c4147;
output c637;
output c9315;
output c449;
output c8379;
output c1202;
output c9147;
output c115;
output c6203;
output c0290;
output c0443;
output c2108;
output c286;
output c0330;
output c3246;
output c9452;
output c889;
output c0365;
output c4284;
output c8254;
output c8141;
output c4247;
output c2482;
output c075;
output c9258;
output c9217;
output c8304;
output c74;
output c8204;
output c6387;
output c6230;
output c4282;
output c543;
output c895;
output c4473;
output c3436;
output c0145;
output c9339;
output c3271;
output c872;
output c7412;
output c2313;
output c6333;
output c7116;
output c3397;
output c0328;
output c9287;
output c0314;
output c6191;
output c4416;
output c5483;
output c9431;
output c7443;
output c7423;
output c8456;
output c9198;
output c3234;
output c2222;
output c687;
output c3465;
output c9346;
output c098;
output c9445;
output c046;
output c6285;
output c218;
output c3153;
output c9182;
output c5173;
output c6374;
output c082;
output c5342;
output c0313;
output c0403;
output c9268;
output c5228;
output c2280;
output c650;
output c093;
output c654;
output c810;
output c966;
output c6221;
output c473;
output c1291;
output c6188;
output c2244;
output c4265;
output c0167;
output c5445;
output c5200;
output c0195;
output c478;
output c6281;
output c5427;
output c7205;
output c0156;
output c7241;
output c926;
output c9280;
output c0193;
output c6120;
output c9103;
output c8128;
output c3326;
output c0428;
output c6278;
output c4243;
output c095;
output c65;
output c2330;
output c2350;
output c2479;
output c0126;
output c3283;
output c6313;
output c0474;
output c357;
output c8442;
output c799;
output c1173;
output c0216;
output c1148;
output c4483;
output c2307;
output c8392;
output c0407;
output c5448;
output c630;
output c439;
output c7156;
output c3180;
output c3411;
output c1386;
output c7120;
output c26;
output c3499;
output c3323;
output c696;
output c6394;
output c2487;
output c1151;
output c6214;
output c9214;
output c492;
output c0386;
output c7268;
output c192;
output c2445;
output c8107;
output c333;
output c991;
output c8458;
output c160;
output c831;
output c1174;
output c1373;
output c4338;
output c913;
output c9238;
output c3172;
output c4316;
output c6296;
output c4486;
output c5180;
output c2133;
output c1497;
output c8402;
output c5296;
output c5307;
output c7209;
output c130;
output c5134;
output c4495;
output c1298;
output c8472;
output c2409;
output c0296;
output c4213;
output c4268;
output c9441;
output c6244;
output c1413;
output c5469;
output c5495;
output c338;
output c4156;
output c0113;
output c0127;
output c021;
output c1499;
output c6100;
output c0327;
output c2346;
output c9102;
output c2255;
output c7397;
output c5187;
output c3423;
output c7365;
output c8341;
output c9236;
output c7109;
output c9304;
output c2153;
output c921;
output c3161;
output c2442;
output c3303;
output c6223;
output c0282;
output c7261;
output c7389;
output c464;
output c613;
output c5373;
output c6495;
output c3292;
output c5439;
output c693;
output c442;
output c2128;
output c0334;
output c9223;
output c6406;
output c3489;
output c0206;
output c9378;
output c7318;
output c722;
output c3359;
output c8328;
output c4322;
output c8248;
output c531;
output c712;
output c7196;
output c9493;
output c522;
output c8123;
output c0134;
output c6141;
output c3247;
output c1238;
output c910;
output c3183;
output c413;
output c6447;
output c0352;
output c136;
output c4275;
output c0174;
output c6442;
output c2466;
output c2406;
output c3284;
output c0418;
output c932;
output c9139;
output c5472;
output c2132;
output c998;
output c8359;
output c7485;
output c5156;
output c6165;
output c1369;
output c5231;
output c1402;
output c7479;
output c9307;
output c5210;
output c877;
output c5382;
output c3201;
output c096;
output c3169;
output c4402;
output c2208;
output c4491;
output c0412;
output c070;
output c4240;
output c4112;
output c1126;
output c59;
output c941;
output c1426;
output c9110;
output c0103;
output c1153;
output c2274;
output c1371;
output c5341;
output c0239;
output c156;
output c2111;
output c241;
output c376;
output c8168;
output c270;
output c6489;
output c8430;
output c4368;
output c34;
output c9333;
output c238;
output c6209;
output c4457;
output c7245;
output c6386;
output c2162;
output c4384;
output c9183;
output c0220;
output c8102;
output c9409;
output c4492;
output c345;
output c9425;
output c9194;
output c4370;
output c0485;
output c4146;
output c389;
output c354;
output c4334;
output c572;
output c0462;
output c6484;
output c6494;
output c4175;
output c948;
output c247;
output c1299;
output c826;
output c556;
output c3415;
output c7147;
output c4225;
output c7425;
output c7411;
output c0317;
output c5211;
output c1327;
output c660;
output c4326;
output c9397;
output c4380;
output c5466;
output c6348;
output c496;
output c6371;
output c3254;
output c5338;
output c7248;
output c2249;
output c6304;
output c2489;
output c1374;
output c5354;
output c6159;
output c0409;
output c5364;
output c1368;
output c2262;
output c4236;
output c410;
output c3378;
output c147;
output c162;
output c9415;
output c43;
output c8492;
output c771;
output c8432;
output c378;
output c8425;
output c7495;
output c9178;
output c2296;
output c9128;
output c239;
output c0337;
output c3341;
output c0304;
output c6411;
output c8223;
output c4358;
output c9482;
output c6338;
output c5476;
output c322;
output c0445;
output c0175;
output c9250;
output c2259;
output c7498;
output c1198;
output c6128;
output c564;
output c1168;
output c3483;
output c3101;
output c5384;
output c972;
output c438;
output c1261;
output c6206;
output c8398;
output c0269;
output c6251;
output c596;
output c9311;
output c458;
output c2387;
output c2371;
output c7445;
output c3275;
output c3305;
output c6163;
output c587;
output c9293;
output c350;
output c9164;
output c2202;
output c7164;
output c8116;
output c4211;
output c4325;
output c5206;
output c0476;
output c2117;
output c9308;
output c1180;
output c2122;
output c7384;
output c3264;
output c4179;
output c8488;
output c656;
output c99;
output c8126;
output c1312;
output c2444;
output c0300;
output c573;
output c3342;
output c0217;
output c5418;
output c6121;
output c3267;
output c755;
output c672;
output c641;
output c7129;
output c3251;
output c1118;
output c5170;
output c4163;
output c4360;
output c7309;
output c6170;
output c6112;
output c1389;
output c9318;
output c3389;
output c9279;
output c0140;
output c6174;
output c277;
output c2197;
output c540;
output c7165;
output c915;
output c539;
output c4498;
output c5279;
output c6355;
output c619;
output c5118;
output c4148;
output c9347;
output c8149;
output c1445;
output c0432;
output c4499;
output c8491;
output c0159;
output c5124;
output c441;
output c3280;
output c9350;
output c9412;
output c6449;
output c7267;
output c4299;
output c1278;
output c786;
output c2169;
output c9278;
output c7162;
output c15;
output c011;
output c3361;
output c9370;
output c9405;
output c9145;
output c3178;
output c3471;
output c4237;
output c577;
output c4375;
output c2160;
output c0429;
output c225;
output c7158;
output c8484;
output c1103;
output c731;
output c7401;
output c8451;
output c0470;
output c0333;
output c9381;
output c3396;
output c9129;
output c5444;
output c8450;
output c2353;
output c2357;
output c4185;
output c117;
output c9256;
output c9474;
output c8336;
output c5381;
output c2412;
output c372;
output c1223;
output c9117;
output c0460;
output c6224;
output c863;
output c1196;
output c151;
output c5474;
output c415;
output c9234;
output c7335;
output c3212;
output c5285;
output c3419;
output c1252;
output c9374;
output c95;
output c785;
output c1112;
output c173;
output c4117;
output c2303;
output c6408;
output c3402;
output c6487;
output c1192;
output c477;
output c5159;
output c4458;
output c5329;
output c6399;
output c8186;
output c146;
output c9163;
output c8205;
output c7307;
output c9325;
output c6306;
output c1127;
output c633;
output c0495;
output c9260;
output c1199;
output c0148;
output c5262;
output c2125;
output c48;
output c849;
output c1427;
output c5138;
output c1498;
output c6478;
output c6115;
output c9489;
output c0266;
output c0125;
output c0450;
output c3309;
output c5113;
output c8423;
output c078;
output c092;
output c7106;
output c0440;
output c3195;
output c7133;
output c0335;
output c3362;
output c6126;
output c6480;
output c3440;
output c0177;
output c3363;
output c4131;
output c2121;
output c763;
output c3477;
output c4104;
output c559;
output c142;
output c8317;
output c3109;
output c1330;
output c0130;
output c3473;
output c9306;
output c184;
output c219;
output c1479;
output c9224;
output c1444;
output c3302;
output c7390;
output c3245;
output c7444;
output c072;
output c120;
output c3321;
output c931;
output c4124;
output c9485;
output c7418;
output c1399;
output c183;
output c411;
output c3462;
output c3216;
output c0472;
output c530;
output c9328;
output c6473;
output c6429;
output c0198;
output c0275;
output c0415;
output c714;
output c7201;
output c099;
output c7135;
output c9418;
output c5321;
output c8489;
output c351;
output c8192;
output c7194;
output c25;
output c8261;
output c8127;
output c7470;
output c4305;
output c4246;
output c8302;
output c1451;
output c7127;
output c1171;
output c0242;
output c1131;
output c9494;
output c8229;
output c7471;
output c823;
output c4417;
output c4209;
output c273;
output c8260;
output c8282;
output c127;
output c7408;
output c3476;
output c4308;
output c9283;
output c2272;
output c5437;
output c2327;
output c8164;
output c8389;
output c461;
output c5265;
output c1378;
output c7422;
output c8200;
output c740;
output c41;
output c560;
output c5276;
output c447;
output c4319;
output c5281;
output c811;
output c5410;
output c954;
output c2267;
output c7493;
output c3250;
output c420;
output c2300;
output c4293;
output c5370;
output c4428;
output c131;
output c2239;
output c1485;
output c6459;
output c1101;
output c8210;
output c2110;
output c386;
output c9411;
output c5399;
output c9354;
output c8288;
output c9141;
output c765;
output c6315;
output c9115;
output c4144;
output c3399;
output c6122;
output c1307;
output c7229;
output c1439;
output c1125;
output c8239;
output c9398;
output c6232;
output c3296;
output c0243;
output c296;
output c3308;
output c6456;
output c8386;
output c720;
output c7263;
output c237;
output c3110;
output c7336;
output c4302;
output c391;
output c599;
output c5433;
output c2219;
output c334;
output c3412;
output c5103;
output c3113;
output c5186;
output c0464;
output c9243;
output c9184;
output c533;
output c5111;
output c7450;
output c81;
output c3255;
output c2389;
output c4426;
output c4436;
output c5407;
output c4335;
output c6317;
output c31;
output c8221;
output c532;
output c3192;
output c4257;
output c689;
output c7131;
output c455;
output c956;
output c4255;
output c211;
output c6194;
output c514;
output c9407;
output c7489;
output c555;
output c5205;
output c7145;
output c9392;
output c7183;
output c118;
output c1124;
output c8463;
output c1227;
output c8314;
output c6190;
output c658;
output c8400;
output c7421;
output c2411;
output c999;
output c5272;
output c5459;
output c9289;
output c9153;
output c0375;
output c412;
output c7491;
output c6155;
output c3270;
output c3165;
output c3381;
output c3168;
output c8474;
output c3349;
output c6471;
output c9240;
output c5169;
output c212;
output c1385;
output c036;
output c8394;
output c0369;
output c53;
output c4245;
output c7364;
output c9151;
output c4329;
output c4489;
output c0353;
output c9296;
output c5227;
output c7139;
output c0237;
output c0280;
output c4161;
output c3366;
output c213;
output c1421;
output c8448;
output c1183;
output c986;
output c6378;
output c3405;
output c3325;
output c6343;
output c5167;
output c5216;
output c3356;
output c2241;
output c5402;
output c6249;
output c6103;
output c71;
output c2322;
output c7387;
output c5277;
output c3295;
output c922;
output c5428;
output c8428;
output c347;
output c214;
output c828;
output c2391;
output c5351;
output c5357;
output c483;
output c8117;
output c4108;
output c8236;
output c3198;
output c0279;
output c0383;
output c8231;
output c9156;
output c2291;
output c9138;
output c0431;
output c8219;
output c6113;
output c0257;
output c2243;
output c7329;
output c4261;
output c2189;
output c9195;
output c4214;
output c4171;
output c476;
output c3147;
output c0341;
output c1140;
output c4259;
output c216;
output c384;
output c2441;
output c223;
output c2266;
output c8417;
output c2131;
output c1246;
output c1493;
output c5204;
output c6361;
output c7301;
output c3334;
output c2235;
output c5289;
output c5229;
output c9161;
output c32;
output c5496;
output c3185;
output c4424;
output c9386;
output c1365;
output c388;
output c6474;
output c6435;
output c7255;
output c434;
output c067;
output c3404;
output c5136;
output c8156;
output c3151;
output c586;
output c1473;
output c4475;
output c3175;
output c9457;
output c0408;
output c2428;
output c0394;
output c5473;
output c2399;
output c4122;
output c2354;
output c2349;
output c7126;
output c3269;
output c8121;
output c4195;
output c2297;
output c5363;
output c6414;
output c0233;
output c5101;
output c6416;
output c1229;
output c0244;
output c897;
output c3166;
output c3108;
output c5198;
output c3416;
output c6270;
output c9113;
output c3253;
output c9133;
output c8115;
output c987;
output c8287;
output c9222;
output c119;
output c7406;
output c1484;
output c7274;
output c834;
output c6101;
output c1102;
output c7117;
output c8326;
output c4296;
output c9483;
output c815;
output c9427;
output c959;
output c4142;
output c9192;
output c5359;
output c4190;
output c9428;
output c9338;
output c3140;
output c1492;
output c145;
output c1264;
output c465;
output c1236;
output c1428;
output c8454;
output c961;
output c9440;
output c923;
output c6280;
output c8273;
output c516;
output c4480;
output c5131;
output c611;
output c698;
output c5172;
output c0249;
output c2310;
output c8172;
output c2182;
output c0152;
output c8320;
output c0326;
output c3276;
output c8384;
output c0421;
output c649;
output c0143;
output c4279;
output c185;
output c5178;
output c6248;
output c0299;
output c471;
output c2402;
output c3194;
output c5374;
output c6149;
output c5375;
output c4239;
output c4233;
output c6336;
output c2449;
output c426;
output c4377;
output c6428;
output c0395;
output c457;
output c250;
output c1220;
output c2370;
output c7323;
output c7295;
output c267;
output c168;
output c73;
output c9210;
output c217;
output c5109;
output c886;
output c5430;
output c8353;
output c180;
output c5434;
output c3163;
output c7282;
output c952;
output c8177;
output c5259;
output c878;
output c8375;
output c8435;
output c575;
output c7374;
output c8267;
output c4493;
output c4348;
output c7467;
output c5454;
output c1353;
output c2148;
output c0116;
output c58;
output c9404;
output c7434;
output c423;
output c970;
output c940;
output c6450;
output c3256;
output c2205;
output c314;
output c8135;
output c9277;
output c523;
output c9188;
output c288;
output c4469;
output c9432;
output c1416;
output c1271;
output c8199;
output c2210;
output c995;
output c33;
output c9356;
output c957;
output c5446;
output c5415;
output c6493;
output c7208;
output c758;
output c186;
output c5223;
output c1149;
output c6485;
output c370;
output c294;
output c3104;
output c2382;
output c7481;
output c11;
output c1265;
output c4413;
output c9322;
output c5184;
output c8479;
output c141;
output c4403;
output c0336;
output c0387;
output c2493;
output c2284;
output c2158;
output c275;
output c6460;
output c5218;
output c950;
output c4189;
output c4399;
output c719;
output c8301;
output c263;
output c515;
output c8143;
output c0276;
output c3158;
output c517;
output c3176;
output c9463;
output c1423;
output c3249;
output c268;
output c759;
output c0204;
output c3210;
output c7325;
output c1442;
output c7403;
output c4158;
output c7210;
output c7320;
output c8348;
output c9265;
output c5379;
output c8170;
output c019;
output c5475;
output c4155;
output c0438;
output c1372;
output c871;
output c993;
output c5457;
output c4387;
output c3136;
output c0137;
output c7476;
output c2426;
output c9324;
output c6269;
output c4393;
output c030;
output c8480;
output c589;
output c9499;
output c8147;
output c5487;
output c6169;
output c385;
output c4281;
output c0215;
output c94;
output c053;
output c260;
output c9462;
output c738;
output c6412;
output c1141;
output c6462;
output c9302;
output c6134;
output c1289;
output c0172;
output c9125;
output c8412;
output c7170;
output c2159;
output c9377;
output c7424;
output c7169;
output c7189;
output c3435;
output c361;
output c4285;
output c1345;
output c462;
output c756;
output c9376;
output c0401;
output c9301;
output c2245;
output c2305;
output c049;
output c3120;
output c037;
output c2170;
output c1283;
output c5484;
output c3438;
output c8362;
output c7302;
output c469;
output c1161;
output c8169;
output c8106;
output c5333;
output c3424;
output c1458;
output c8227;
output c916;
output c884;
output c9475;
output c6189;
output c2343;
output c1237;
output c4197;
output c664;
output c4355;
output c452;
output c8298;
output c1276;
output c055;
output c4173;
output c7334;
output c2485;
output c4139;
output c2362;
output c427;
output c8335;
output c1123;
output c7281;
output c283;
output c7337;
output c9340;
output c8173;
output c3263;
output c78;
output c4313;
output c6440;
output c8280;
output c5141;
output c917;
output c7363;
output c795;
output c887;
output c2383;
output c4456;
output c685;
output c0349;
output c112;
output c930;
output c9357;
output c5422;
output c4206;
output c914;
output c6379;
output c9205;
output c195;
output c6143;
output c5266;
output c67;
output c06;
output c8408;
output c6314;
output c222;
output c2326;
output c5300;
output c5339;
output c4311;
output c9367;
output c770;
output c0169;
output c725;
output c1314;
output c4462;
output c7197;
output c7472;
output c7122;
output c7328;
output c0157;
output c4374;
output c3385;
output c6431;
output c8388;
output c364;
output c3387;
output c776;
output c1335;
output c5319;
output c8196;
output c5139;
output c5179;
output c8262;
output c2179;
output c6286;
output c5326;
output c6294;
output c352;
output c1343;
output c9157;
output c7289;
output c3420;
output c4140;
output c717;
output c6256;
output c0265;
output c0292;
output c1165;
output c397;
output c290;
output c0180;
output c3127;
output c287;
output c8397;
output c6235;
output c1286;
output c4362;
output c3432;
output c0321;
output c7339;
output c293;
output c2295;
output c0457;
output c639;
output c7195;
output c6390;
output c236;
output c0435;
output c0135;
output c251;
output c2339;
output c2124;
output c4231;
output c5470;
output c5135;
output c0212;
output c9118;
output c624;
output c1152;
output c4165;
output c829;
output c0119;
output c9451;
output c5372;
output c3221;
output c548;
output c942;
output c8237;
output c3307;
output c7279;
output c9254;
output c276;
output c9442;
output c8476;
output c0231;
output c077;
output c962;
output c3443;
output c0100;
output c8198;
output c9173;
output c5147;
output c5395;
output c8473;
output c2302;
output c2401;
output c5126;
output c4303;
output c8347;
output c3124;
output c175;
output c087;
output c9388;
output c1475;
output c6347;
output c2167;
output c860;
output c0142;
output c3105;
output c520;
output c8281;
output c245;
output c0191;
output c0467;
output c3222;
output c4295;
output c1280;
output c8278;
output c1117;
output c888;
output c5253;
output c8485;
output c346;
output c7230;
output c2384;
output c2315;
output c8407;
output c7277;
output c3332;
output c843;
output c6106;
output c2242;
output c1100;
output c5316;
output c0420;
output c0225;
output c6312;
output c767;
output c8437;
output c256;
output c9150;
output c4346;
output c8370;
output c04;
output c1310;
output c5440;
output c199;
output c2155;
output c3177;
output c113;
output c2425;
output c197;
output c6258;
output c5486;
output c9455;
output c21;
output c4278;
output c2251;
output c8217;
output c18;
output c8224;
output c6356;
output c09;
output c0185;
output c4331;
output c3429;
output c8228;
output c2201;
output c5394;
output c8272;
output c7102;
output c657;
output c4477;
output c37;
output c3480;
output c1316;
output c7431;
output c484;
output c4114;
output c4366;
output c9131;
output c9417;
output c0377;
output c3430;
output c4277;
output c955;
output c9281;
output c7453;
output c825;
output c475;
output c444;
output c8274;
output c5154;
output c46;
output c2190;
output c6481;
output c3228;
output c5334;
output c6479;
output c7265;
output c7367;
output c8487;
output c2407;
output c6262;
output c690;
output c70;
output c929;
output c4162;
output c1293;
output c0323;
output c6376;
output c5108;
output c5215;
output c1417;
output c6346;
output c9197;
output c0393;
output c3259;
output c838;
output c079;
output c8433;
output c847;
output c0109;
output c2119;
output c3232;
output c7226;
output c2207;
output c632;
output c6123;
output c960;
output c5294;
output c1469;
output c2316;
output c7153;
output c6116;
output c3320;
output c1401;
output c66;
output c3193;
output c39;
output c6417;
output c8241;
output c0473;
output c7232;
output c6225;
output c4113;
output c2394;
output c3380;
output c5137;
output c1478;
output c7378;
output c518;
output c3111;
output c4337;
output c0278;
output c4207;
output c938;
output c9213;
output c7151;
output c031;
output c3131;
output c8235;
output c6137;
output c5264;
output c6369;
output c2114;
output c715;
output c730;
output c8406;
output c8153;
output c2459;
output c4435;
output c5195;
output c2356;
output c852;
output c1491;
output c3441;
output c6289;
output c3421;
output c2453;
output c7399;
output c9448;
output c0306;
output c5236;
output c1249;
output c2290;
output c3472;
output c7486;
output c122;
output c6205;
output c3319;
output c6186;
output c4203;
output c4453;
output c0493;
output c7104;
output c3242;
output c546;
output c2237;
output c1318;
output c3347;
output c7154;
output c8234;
output c5189;
output c2447;
output c0247;
output c5488;
output c0361;
output c7379;
output c9109;
output c8366;
output c6364;
output c746;
output c9237;
output c5346;
output c470;
output c5222;
output c6268;
output c827;
output c6463;
output c8330;
output c0392;
output c3365;
output c5295;
output c1104;
output c8427;
output c9394;
output c6357;
output c93;
output c3484;
output c3215;
output c620;
output c5337;
output c2469;
output c8290;
output c0205;
output c3103;
output c7341;
output c8197;
output c1231;
output c8351;
output c9429;
output c6499;
output c2172;
output c3266;
output c527;
output c1240;
output c0305;
output c9246;
output c029;
output c1162;
output c0496;
output c2443;
output c4400;
output c194;
output c6302;
output c2185;
output c5194;
output c3281;
output c6272;
output c1245;
output c6241;
output c2176;
output c9331;
output c178;
output c2282;
output c2476;
output c6323;
output c0482;
output c1242;
output c9330;
output c2496;
output c1170;
output c3439;
output c3300;
output c0446;
output c3154;
output c2381;
output c9285;
output c1272;
output c4401;
output c0297;
output c2147;
output c557;
output c2264;
output c0494;
output c2480;
output c3316;
output c5414;
output c4169;
output c9469;
output c6212;
output c360;
output c9335;
output c6124;
output c0235;
output c8138;
output c3398;
output c3335;
output c2289;
output c02;
output c989;
output c1222;
output c8175;
output c9120;
output c526;
output c8360;
output c7185;
output c919;
output c3167;
output c2374;
output c3368;
output c291;
output c7454;
output c3237;
output c4121;
output c4409;
output c8269;
output c0163;
output c996;
output c332;
output c8125;
output c9106;
output c0188;
output c022;
output c676;
output c1317;
output c5273;
output c1226;
output c9232;
output c511;
output c0308;
output c9410;
output c9259;
output c7414;
output c9290;
output c382;
output c2101;
output c1200;
output c1188;
output c2363;
output c0451;
output c280;
output c6219;
output c8218;
output c3226;
output c4103;
output c5123;
output c5443;
output c7306;
output c8413;
output c4441;
output c0213;
output c2365;
output c723;
output c958;
output c5310;
output c182;
output c7451;
output c7353;
output c4258;
output c8424;
output c9257;
output c2278;
output c9321;
output c227;
output c510;
output c4470;
output c6381;
output c4395;
output c1315;
output c1359;
output c2143;
output c318;
output c4488;
output c7137;
output c2452;
output c0346;
output c2184;
output c8179;
output c7416;
output c1367;
output c8207;
output c8120;
output c2436;
output c4136;
output c1447;
output c0124;
output c0489;
output c3312;
output c0447;
output c1347;
output c8429;
output c0132;
output c8332;
output c8446;
output c289;
output c1376;
output c4286;
output c1181;
output c9212;
output c858;
output c392;
output c9253;
output c0154;
output c8490;
output c3238;
output c6475;
output c6340;
output c822;
output c4310;
output c5244;
output c5125;
output c499;
output c0441;
output c5492;
output c8396;
output c8203;
output c7478;
output c0187;
output c435;
output c436;
output c2144;
output c6366;
output c8352;
output c187;
output c0329;
output c7278;
output c0479;
output c2261;
output c221;
output c5110;
output c7298;
output c9202;
output c9470;
output c9166;
output c035;
output c2188;
output c4429;
output c5304;
output c7463;
output c824;
output c7223;
output c8350;
output c5408;
output c327;
output c0104;
output c9375;
output c5305;
output c5447;
output c9488;
output c2314;
output c8140;
output c8315;
output c2178;
output c045;
output c5419;
output c6342;
output c4349;
output c6389;
output c4266;
output c1456;
output c2488;
output c4138;
output c6279;
output c7310;
output c1119;
output c6445;
output c5464;
output c8259;
output c2324;
output c5129;
output c3392;
output c9484;
output c732;
output c1446;
output c468;
output c7115;
output c0471;
output c6415;
output c0184;
output c935;
output c17;
output c9275;
output c3290;
output c3367;
output c6132;
output c315;
output c9190;
output c083;
output c5268;
output c8255;
output c8299;
output c1203;
output c7409;
output c2253;
output c4166;
output c1195;
output c1250;
output c8119;
output c6446;
output c1217;
output c56;
output c489;
output c3220;
output c6200;
output c0200;
output c6166;
output c8167;
output c9352;
output c0423;
output c086;
output c3199;
output c4333;
output c8112;
output c2336;
output c9100;
output c258;
output c7243;
output c2369;
output c9261;
output c1467;
output c422;
output c1216;
output c456;
output c9323;
output c7469;
output c739;
output c5280;
output c3410;
output c6391;
output c170;
output c692;
output c0366;
output c3117;
output c8306;
output c5350;
output c448;
output c7293;
output c8188;
output c1394;
output c585;
output c9148;
output c9204;
output c563;
output c4411;
output c3344;
output c2378;
output c2105;
output c9196;
output c1221;
output c0385;
output c0410;
output c5127;
output c7385;
output c054;
output c1391;
output c652;
output c667;
output c7447;
output c44;
output c750;
output c9227;
output c052;
output c6196;
output c614;
output c3156;
output c899;
output c8132;
output c143;
output c6136;
output c6157;
output c4369;
output c7462;
output c4484;
output c8144;
output c4431;
output c3209;
output c830;
output c618;
output c571;
output c1340;
output c6430;
output c0248;
output c3353;
output c7394;
output c4204;
output c832;
output c565;
output c5303;
output c2141;
output c544;
output c6469;
output c0345;
output c582;
output c7157;
output c6362;
output c4420;
output c1384;
output c5413;
output c5199;
output c736;
output c3235;
output c7420;
output c4379;
output c0307;
output c4252;
output c7314;
output c7159;
output c846;
output c4460;
output c0219;
output c8459;
output c7458;
output c3293;
output c7134;
output c5471;
output c0255;
output c615;
output c3369;
output c7346;
output c7179;
output c8334;
output c9332;
output c3159;
output c0325;
output c754;
output c5293;
output c4241;
output c9382;
output c7326;
output c0202;
output c0382;
output c1349;
output c1169;
output c7415;
output c339;
output c8152;
output c52;
output c9423;
output c1241;
output c7270;
output c985;
output c3355;
output c789;
output c2472;
output c7182;
output c3206;
output c165;
output c3115;
output c3377;
output c3174;
output c3311;
output c7237;
output c3481;
output c2308;
output c1128;
output c7321;
output c6377;
output c2161;
output c1160;
output c6105;
output c2206;
output c1147;
output c7359;
output c7144;
output c6208;
output c854;
output c3223;
output c7430;
output c0240;
output c2368;
output c1254;
output c3299;
output c6239;
output c2463;
output c2191;
output c8399;
output c2461;
output c857;
output c440;
output c2127;
output c1461;
output c86;
output c8333;
output c3191;
output c1329;
output c5479;
output c2226;
output c1144;
output c8498;
output c992;
output c4283;
output c0351;
output c9122;
output c1459;
output c4439;
output c9403;
output c2337;
output c0499;
output c1460;
output c0291;
output c4193;
output c1382;
output c768;
output c3495;
output c1486;
output c40;
output c7288;
output c7256;
output c8243;
output c0468;
output c8275;
output c1362;
output c4164;
output c242;
output c8403;
output c6490;
output c137;
output c760;
output c129;
output c2269;
output c3231;
output c8191;
output c1476;
output c7386;
output c023;
output c9395;
output c5332;
output c7130;
output c124;
output c7190;
output c7402;
output c6252;
output c1392;
output c7252;
output c7304;
output c6439;
output c0162;
output c479;
output c6111;
output c2403;
output c6216;
output c5106;
output c2129;
output c432;
output c9199;
output c1113;
output c497;
output c5286;
output c0402;
output c981;
output c8103;
output c2130;
output c524;
output c4365;
output c7474;
output c5234;
output c783;
output c3401;
output c6144;
output c679;
output c1259;
output c6127;
output c1306;
output c4130;
output c1105;
output c3461;
output c4119;
output c5383;
output c6179;
output c2254;
output c5467;
output c1191;
output c9186;
output c743;
output c7240;
output c0158;
output c4459;
output c2275;
output c8270;
output c5385;
output c0302;
output c6162;
output c6426;
output c5168;
output c3214;
output c2398;
output c7305;
output c1288;
output c8142;
output c6135;
output c1208;
output c6172;
output c0362;
output c662;
output c179;
output c6207;
output c4465;
output c7459;
output c7206;
output c580;
output c2138;
output c261;
output c9478;
output c97;
output c9160;
output c454;
output c7247;
output c8220;
output c4323;
output c6198;
output c6320;
output c9226;
output c0340;
output c6167;
output c0379;
output c6119;
output c4184;
output c3382;
output c068;
output c328;
output c3428;
output c3239;
output c4192;
output c2240;
output c3330;
output c6275;
output c2102;
output c6277;
output c9496;
output c3291;
output c3475;
output c8242;
output c661;
output c158;
output c7349;
output c4120;
output c3492;
output c0203;
output c8157;
output c72;
output c7128;
output c3112;
output c6283;
output c1346;
output c7492;
output c4421;
output c5465;
output c8318;
output c363;
output c2497;
output c7360;
output c980;
output c3453;
output c5226;
output c0376;
output c9231;
output c4159;
output c68;
output c6452;
output c9414;
output c968;
output c4220;
output c6253;
output c8292;
output c244;
output c1481;
output c3128;
output c0287;
output c8467;
output c097;
output c7175;
output c9158;
output c718;
output c0136;
output c0166;
output c8377;
output c787;
output c6287;
output c7108;
output c1422;
output c19;
output c7497;
output c549;
output c8252;
output c2294;
output c8376;
output c7391;
output c5378;
output c7111;
output c590;
output c6419;
output c953;
output c7213;
output c4110;
output c4408;
output c5120;
output c9314;
output c1210;
output c4405;
output c7437;
output c23;
output c374;
output c869;
output c4476;
output c3142;
output c7299;
output c4478;
output c0463;
output c7160;
output c7400;
output c3272;
output c9343;
output c2135;
output c6344;
output c5267;
output c6477;
output c344;
output c3343;
output c4471;
output c1292;
output c6461;
output c8497;
output c5202;
output c5166;
output c4396;
output c1150;
output c0147;
output c8316;
output c7340;
output c6421;
output c2418;
output c6292;
output c5220;
output c1463;
output c4340;
output c4199;
output c3374;
output c0344;
output c264;
output c3452;
output c3373;
output c8136;
output c8344;
output c8305;
output c1454;
output c8268;
output c13;
output c348;
output c4327;
output c4276;
output c2320;
output c5301;
output c6410;
output c0230;
output c0398;
output c697;
output c890;
output c8160;
output c246;
output c4143;
output c7383;

assign c00 =  x174 &  x452 & ~x10 & ~x50 & ~x282 & ~x309 & ~x310 & ~x583 & ~x615 & ~x640 & ~x690 & ~x691 & ~x716 & ~x717 & ~x718 & ~x724 & ~x726 & ~x749 & ~x752;
assign c02 =  x229 &  x397 & ~x23 & ~x66 & ~x209 & ~x210 & ~x611 & ~x612 & ~x644 & ~x647 & ~x703 & ~x748 & ~x782;
assign c04 = ~x1 & ~x98 & ~x265 & ~x270 & ~x271 & ~x502 & ~x587 & ~x602 & ~x628 & ~x638 & ~x673 & ~x701 & ~x742 & ~x769;
assign c06 =  x93 &  x233 &  x289 &  x428 & ~x13 & ~x28 & ~x43 & ~x52 & ~x71 & ~x138 & ~x184 & ~x195 & ~x213 & ~x252 & ~x336 & ~x337 & ~x617 & ~x670 & ~x671 & ~x673 & ~x698 & ~x727 & ~x728 & ~x751 & ~x757 & ~x759;
assign c08 = ~x5 & ~x25 & ~x39 & ~x46 & ~x94 & ~x235 & ~x290 & ~x317 & ~x318 & ~x475 & ~x476 & ~x557 & ~x582 & ~x583 & ~x724 & ~x750 & ~x751 & ~x764;
assign c010 =  x585 & ~x2 & ~x55 & ~x248 & ~x251 & ~x252 & ~x303 & ~x304 & ~x307 & ~x333 & ~x338 & ~x392 & ~x728 & ~x729 & ~x738 & ~x739 & ~x758 & ~x783;
assign c012 =  x286 &  x482 &  x591 & ~x38 & ~x39 & ~x41 & ~x128 & ~x245 & ~x272 & ~x419 & ~x421 & ~x423 & ~x449 & ~x476 & ~x724 & ~x752;
assign c014 =  x174 &  x370 & ~x9 & ~x11 & ~x27 & ~x39 & ~x167 & ~x186 & ~x187 & ~x236 & ~x237 & ~x476 & ~x587 & ~x724 & ~x727 & ~x732;
assign c016 =  x509;
assign c018 =  x65 &  x93 &  x205 &  x345 & ~x14 & ~x466 & ~x649 & ~x727 & ~x759;
assign c020 =  x445 & ~x18 & ~x23 & ~x30 & ~x45 & ~x47 & ~x48 & ~x51 & ~x54 & ~x69 & ~x74 & ~x75 & ~x99 & ~x101 & ~x102 & ~x104 & ~x128 & ~x129 & ~x132 & ~x134 & ~x135 & ~x161 & ~x164 & ~x166 & ~x293 & ~x336 & ~x365 & ~x392 & ~x413 & ~x561 & ~x587 & ~x642 & ~x643 & ~x669 & ~x670 & ~x698 & ~x699 & ~x724 & ~x734 & ~x736 & ~x751 & ~x757 & ~x758 & ~x759 & ~x761;
assign c022 =  x143 &  x145 &  x147 &  x175 &  x397 & ~x12 & ~x310;
assign c024 =  x234 & ~x14 & ~x26 & ~x40 & ~x41 & ~x42 & ~x46 & ~x53 & ~x57 & ~x80 & ~x81 & ~x102 & ~x108 & ~x136 & ~x139 & ~x141 & ~x195 & ~x213 & ~x241 & ~x378 & ~x379 & ~x421 & ~x560 & ~x698 & ~x699 & ~x752 & ~x783;
assign c026 =  x229 &  x397 &  x426 & ~x12 & ~x243 & ~x365 & ~x366 & ~x392 & ~x680 & ~x695 & ~x722 & ~x723 & ~x730 & ~x758;
assign c028 =  x485 & ~x8 & ~x16 & ~x41 & ~x45 & ~x97 & ~x270 & ~x300 & ~x301 & ~x327 & ~x329 & ~x356 & ~x364 & ~x420 & ~x585 & ~x639 & ~x666 & ~x692 & ~x695 & ~x696 & ~x702 & ~x725 & ~x730 & ~x774 & ~x775 & ~x778;
assign c030 =  x175 &  x231 &  x482 & ~x52 & ~x53 & ~x54 & ~x55 & ~x83 & ~x96 & ~x125 & ~x181 & ~x236 & ~x364 & ~x681 & ~x703 & ~x729 & ~x731 & ~x755 & ~x768 & ~x782;
assign c032 = ~x1 & ~x2 & ~x8 & ~x10 & ~x67 & ~x134 & ~x364 & ~x581 & ~x585 & ~x617 & ~x620 & ~x637 & ~x643 & ~x645 & ~x646 & ~x648 & ~x654 & ~x673 & ~x681 & ~x690 & ~x697 & ~x701 & ~x732 & ~x748 & ~x750 & ~x782;
assign c034 =  x485 & ~x3 & ~x5 & ~x97 & ~x99 & ~x100 & ~x136 & ~x141 & ~x157 & ~x188 & ~x194 & ~x378 & ~x424 & ~x469 & ~x767 & ~x778 & ~x783;
assign c036 = ~x24 & ~x28 & ~x53 & ~x56 & ~x57 & ~x62 & ~x82 & ~x118 & ~x128 & ~x138 & ~x165 & ~x188 & ~x224 & ~x335 & ~x336 & ~x420 & ~x470 & ~x523 & ~x553 & ~x617 & ~x673 & ~x729 & ~x769;
assign c038 = ~x41 & ~x217 & ~x290 & ~x300 & ~x318 & ~x329 & ~x336 & ~x393 & ~x394 & ~x737 & ~x742 & ~x752 & ~x754 & ~x755 & ~x760 & ~x768 & ~x771;
assign c040 =  x528 & ~x129 & ~x183 & ~x240 & ~x277 & ~x297 & ~x350 & ~x414;
assign c042 =  x429 & ~x13 & ~x268 & ~x300 & ~x336 & ~x585 & ~x651 & ~x696 & ~x707 & ~x717 & ~x719 & ~x754 & ~x783;
assign c044 =  x314 &  x538 &  x539 &  x630 & ~x10 & ~x14 & ~x638 & ~x699 & ~x773 & ~x775;
assign c046 =  x248;
assign c048 =  x146 &  x147 &  x398 & ~x12 & ~x42 & ~x243 & ~x613 & ~x624 & ~x667 & ~x671 & ~x680 & ~x693 & ~x695 & ~x701 & ~x720 & ~x724 & ~x728 & ~x729 & ~x780;
assign c050 =  x592 &  x593 &  x594 &  x595 & ~x7 & ~x11 & ~x12 & ~x13 & ~x14 & ~x25 & ~x26 & ~x34 & ~x41 & ~x46 & ~x47 & ~x57 & ~x61 & ~x85 & ~x87 & ~x90 & ~x114 & ~x421 & ~x718 & ~x726 & ~x727 & ~x745 & ~x746 & ~x747 & ~x755 & ~x772 & ~x773 & ~x774 & ~x780 & ~x781 & ~x782;
assign c052 = ~x39 & ~x76 & ~x103 & ~x156 & ~x323 & ~x348 & ~x352 & ~x387 & ~x414 & ~x560 & ~x616;
assign c054 =  x167 & ~x125;
assign c056 =  x459 &  x549 & ~x3 & ~x7 & ~x18 & ~x19 & ~x20 & ~x22 & ~x29 & ~x30 & ~x41 & ~x43 & ~x56 & ~x72 & ~x82 & ~x106 & ~x114 & ~x134 & ~x280 & ~x307 & ~x352 & ~x669 & ~x696 & ~x699 & ~x701 & ~x703 & ~x720 & ~x723 & ~x725 & ~x726 & ~x727 & ~x729 & ~x748 & ~x757 & ~x760 & ~x761 & ~x781 & ~x782;
assign c058 =  x351 &  x360 &  x453 & ~x558 & ~x646 & ~x669 & ~x678 & ~x724 & ~x744;
assign c060 =  x83;
assign c062 =  x113 & ~x730;
assign c064 =  x174 &  x333 &  x369 &  x417 &  x444;
assign c066 = ~x54 & ~x212 & ~x364 & ~x464 & ~x590 & ~x666 & ~x704 & ~x715 & ~x732 & ~x770;
assign c068 = ~x27 & ~x29 & ~x41 & ~x43 & ~x77 & ~x83 & ~x166 & ~x170 & ~x213 & ~x240 & ~x281 & ~x296 & ~x558 & ~x560 & ~x586 & ~x590 & ~x618 & ~x645 & ~x693 & ~x699 & ~x706 & ~x754 & ~x759 & ~x774 & ~x783;
assign c070 =  x511 & ~x294 & ~x302 & ~x321 & ~x519 & ~x546 & ~x614 & ~x676 & ~x758;
assign c072 =  x398 &  x595 &  x622 & ~x322 & ~x347 & ~x403 & ~x737;
assign c074 =  x176 & ~x110 & ~x138 & ~x223 & ~x238 & ~x254 & ~x478 & ~x601 & ~x617 & ~x629 & ~x676 & ~x695 & ~x698 & ~x703 & ~x710 & ~x722 & ~x740 & ~x751 & ~x758 & ~x780;
assign c076 = ~x32 & ~x45 & ~x126 & ~x127 & ~x131 & ~x159 & ~x168 & ~x226 & ~x254 & ~x350 & ~x380 & ~x414 & ~x442 & ~x703 & ~x706 & ~x740 & ~x747 & ~x748 & ~x750 & ~x764 & ~x779 & ~x781;
assign c078 =  x135 &  x259 &  x508 & ~x215 & ~x275 & ~x365;
assign c080 = ~x3 & ~x17 & ~x45 & ~x47 & ~x104 & ~x128 & ~x129 & ~x134 & ~x140 & ~x158 & ~x168 & ~x224 & ~x280 & ~x295 & ~x296 & ~x297 & ~x352 & ~x353 & ~x365 & ~x412 & ~x440 & ~x468 & ~x561 & ~x588 & ~x695 & ~x700 & ~x727 & ~x736 & ~x748 & ~x752 & ~x764 & ~x776;
assign c082 =  x453 & ~x8 & ~x44 & ~x48 & ~x66 & ~x67 & ~x266 & ~x291 & ~x421 & ~x503 & ~x587;
assign c084 =  x176 &  x204 &  x482 &  x508 & ~x1 & ~x13 & ~x329 & ~x393 & ~x420 & ~x448 & ~x504 & ~x643 & ~x728 & ~x739 & ~x783;
assign c086 =  x262 &  x290 &  x342 & ~x11 & ~x27 & ~x41 & ~x46 & ~x97 & ~x99 & ~x127 & ~x353 & ~x476 & ~x669 & ~x723 & ~x724 & ~x780;
assign c088 =  x515 & ~x69 & ~x83 & ~x156 & ~x157 & ~x159 & ~x167 & ~x213 & ~x307 & ~x365 & ~x407 & ~x420 & ~x616 & ~x695 & ~x706 & ~x728 & ~x757 & ~x781;
assign c090 =  x485 & ~x0 & ~x3 & ~x10 & ~x22 & ~x27 & ~x32 & ~x42 & ~x116 & ~x141 & ~x155 & ~x182 & ~x198 & ~x224 & ~x238 & ~x392 & ~x420 & ~x640 & ~x641 & ~x642 & ~x668 & ~x671 & ~x693 & ~x695 & ~x722 & ~x725 & ~x728 & ~x747 & ~x754 & ~x763 & ~x768 & ~x776 & ~x782 & ~x783;
assign c092 =  x456 &  x707 & ~x322 & ~x363 & ~x365;
assign c094 =  x175 &  x231 &  x398 & ~x68 & ~x82 & ~x138 & ~x155 & ~x168 & ~x238 & ~x267 & ~x294 & ~x420 & ~x559 & ~x587 & ~x748;
assign c096 =  x501 &  x558 & ~x332 & ~x333 & ~x359 & ~x394;
assign c098 =  x514 &  x515 &  x516 &  x539 & ~x10 & ~x83 & ~x156 & ~x379 & ~x448 & ~x723 & ~x724 & ~x725 & ~x749;
assign c0100 =  x60 &  x90;
assign c0102 =  x204 &  x218 &  x470 & ~x271 & ~x611;
assign c0104 =  x94 &  x344 &  x372 &  x484 & ~x321;
assign c0106 = ~x43 & ~x61 & ~x67 & ~x74 & ~x151 & ~x179 & ~x224 & ~x243 & ~x247 & ~x252 & ~x476 & ~x503 & ~x557 & ~x584 & ~x616 & ~x640 & ~x643 & ~x644 & ~x672 & ~x678 & ~x691 & ~x694;
assign c0108 =  x148 & ~x19 & ~x42 & ~x280 & ~x282 & ~x337 & ~x338 & ~x562 & ~x591 & ~x592 & ~x613 & ~x621 & ~x624 & ~x625 & ~x639 & ~x640 & ~x666 & ~x670 & ~x676 & ~x694 & ~x698 & ~x699 & ~x720 & ~x722 & ~x781;
assign c0110 =  x261 &  x401 &  x569 & ~x3 & ~x6 & ~x11 & ~x12 & ~x13 & ~x29 & ~x30 & ~x40 & ~x43 & ~x59 & ~x140 & ~x143 & ~x392 & ~x393 & ~x420 & ~x644 & ~x673 & ~x698 & ~x729 & ~x756 & ~x759 & ~x760 & ~x762;
assign c0112 =  x254 &  x284 &  x426 &  x454 & ~x318 & ~x330 & ~x365;
assign c0114 = ~x82 & ~x127 & ~x168 & ~x187 & ~x242 & ~x266 & ~x476 & ~x584 & ~x638 & ~x653 & ~x673 & ~x696 & ~x711 & ~x734 & ~x746 & ~x748;
assign c0116 =  x595 & ~x4 & ~x10 & ~x46 & ~x47 & ~x93 & ~x133 & ~x164 & ~x249 & ~x707 & ~x708 & ~x724 & ~x730 & ~x735 & ~x738 & ~x755 & ~x765;
assign c0118 =  x257 &  x258 &  x342 &  x493 &  x520 &  x547 & ~x10 & ~x182 & ~x210;
assign c0120 =  x531 &  x547;
assign c0122 = ~x1 & ~x69 & ~x181 & ~x195 & ~x209 & ~x297 & ~x575 & ~x601 & ~x619 & ~x675 & ~x748;
assign c0124 = ~x6 & ~x7 & ~x21 & ~x26 & ~x29 & ~x31 & ~x34 & ~x37 & ~x40 & ~x41 & ~x49 & ~x63 & ~x122 & ~x152 & ~x196 & ~x347 & ~x476 & ~x556 & ~x558 & ~x584 & ~x612 & ~x613 & ~x615 & ~x639 & ~x665 & ~x666 & ~x667 & ~x670 & ~x674 & ~x692 & ~x693 & ~x700 & ~x719 & ~x720 & ~x727 & ~x734 & ~x740 & ~x744 & ~x764 & ~x766 & ~x770 & ~x772 & ~x774 & ~x775;
assign c0126 =  x539 &  x548 & ~x1 & ~x6 & ~x10 & ~x13 & ~x15 & ~x52 & ~x78 & ~x104 & ~x108 & ~x109 & ~x137 & ~x364 & ~x365 & ~x423 & ~x424 & ~x699 & ~x727 & ~x760 & ~x779 & ~x780;
assign c0128 =  x536 &  x543 & ~x152 & ~x240 & ~x717;
assign c0130 =  x446 &  x457 &  x458 & ~x3 & ~x16 & ~x32 & ~x44 & ~x48 & ~x57 & ~x79 & ~x97 & ~x98 & ~x364 & ~x392 & ~x393 & ~x394 & ~x420 & ~x701 & ~x724 & ~x727;
assign c0132 =  x305 &  x332 &  x455 & ~x39 & ~x97 & ~x98 & ~x337 & ~x366 & ~x640 & ~x763;
assign c0134 = ~x11 & ~x30 & ~x125 & ~x166 & ~x251 & ~x303 & ~x304 & ~x319 & ~x320 & ~x332 & ~x347 & ~x348 & ~x476 & ~x572 & ~x727 & ~x750 & ~x778 & ~x779;
assign c0136 =  x464 & ~x125 & ~x153 & ~x209 & ~x236 & ~x264 & ~x587 & ~x700 & ~x707 & ~x714 & ~x717 & ~x755 & ~x761 & ~x781;
assign c0138 = ~x100 & ~x126 & ~x269 & ~x293 & ~x350 & ~x377 & ~x379 & ~x404 & ~x415 & ~x417 & ~x447 & ~x755 & ~x758;
assign c0140 = ~x8 & ~x9 & ~x10 & ~x129 & ~x236 & ~x310 & ~x346 & ~x374 & ~x377 & ~x548 & ~x712 & ~x730 & ~x759 & ~x768;
assign c0142 =  x147 &  x231 &  x288 &  x399 & ~x193 & ~x239 & ~x294 & ~x295 & ~x732;
assign c0144 =  x111;
assign c0146 =  x507 & ~x14 & ~x32 & ~x41 & ~x263 & ~x290 & ~x331 & ~x337 & ~x366 & ~x759;
assign c0148 =  x201 &  x451 &  x479 & ~x11 & ~x43 & ~x309 & ~x365 & ~x366 & ~x637 & ~x701 & ~x744;
assign c0150 = ~x236 & ~x264 & ~x292 & ~x301 & ~x320 & ~x321 & ~x347 & ~x379 & ~x389 & ~x447 & ~x448 & ~x491 & ~x602 & ~x674;
assign c0152 =  x203 &  x455 & ~x26 & ~x82 & ~x84 & ~x157 & ~x168 & ~x324 & ~x740 & ~x754 & ~x757 & ~x761 & ~x779 & ~x782;
assign c0154 = ~x9 & ~x22 & ~x41 & ~x65 & ~x96 & ~x97 & ~x106 & ~x151 & ~x189 & ~x224 & ~x237 & ~x252 & ~x501 & ~x503 & ~x554 & ~x556 & ~x558 & ~x588 & ~x605 & ~x637 & ~x639 & ~x654 & ~x692 & ~x702 & ~x709 & ~x721;
assign c0156 = ~x4 & ~x15 & ~x80 & ~x100 & ~x239 & ~x531 & ~x558 & ~x559 & ~x561 & ~x573 & ~x599 & ~x617 & ~x626 & ~x641 & ~x648 & ~x671 & ~x675 & ~x703 & ~x723 & ~x724 & ~x729 & ~x751;
assign c0158 =  x480 & ~x65 & ~x296 & ~x318 & ~x344 & ~x348 & ~x434;
assign c0160 = ~x12 & ~x16 & ~x17 & ~x18 & ~x30 & ~x40 & ~x42 & ~x45 & ~x46 & ~x53 & ~x54 & ~x56 & ~x69 & ~x82 & ~x83 & ~x102 & ~x128 & ~x134 & ~x140 & ~x166 & ~x168 & ~x196 & ~x223 & ~x254 & ~x352 & ~x353 & ~x382 & ~x420 & ~x441 & ~x560 & ~x643 & ~x704 & ~x706 & ~x707 & ~x722 & ~x733 & ~x754 & ~x756 & ~x760 & ~x764 & ~x772 & ~x781;
assign c0162 =  x537 & ~x0 & ~x4 & ~x5 & ~x9 & ~x12 & ~x14 & ~x15 & ~x16 & ~x19 & ~x21 & ~x22 & ~x24 & ~x25 & ~x47 & ~x48 & ~x49 & ~x52 & ~x55 & ~x56 & ~x57 & ~x74 & ~x76 & ~x78 & ~x79 & ~x82 & ~x85 & ~x106 & ~x138 & ~x167 & ~x322 & ~x350 & ~x393 & ~x448 & ~x504 & ~x700 & ~x726 & ~x753 & ~x755 & ~x761 & ~x763 & ~x768 & ~x773 & ~x778 & ~x779 & ~x782 & ~x783;
assign c0164 =  x445 &  x460 &  x537 &  x538 &  x539 & ~x44 & ~x47 & ~x74 & ~x103 & ~x138 & ~x163 & ~x164 & ~x251 & ~x731 & ~x757 & ~x759;
assign c0166 =  x518 &  x530 &  x558 & ~x361 & ~x394;
assign c0168 =  x226 &  x230 &  x257 &  x536 & ~x309 & ~x365;
assign c0170 =  x205 & ~x14 & ~x134 & ~x144 & ~x183 & ~x266 & ~x659 & ~x723;
assign c0172 =  x460 & ~x21 & ~x23 & ~x41 & ~x82 & ~x158 & ~x327 & ~x356 & ~x380 & ~x381 & ~x384 & ~x437 & ~x588 & ~x697 & ~x731 & ~x756 & ~x757 & ~x781;
assign c0174 = ~x1 & ~x74 & ~x269 & ~x545 & ~x547 & ~x563 & ~x572 & ~x573 & ~x616 & ~x618 & ~x620 & ~x653 & ~x673 & ~x675;
assign c0176 =  x148 &  x204 &  x288 &  x372 & ~x2 & ~x10 & ~x13 & ~x42 & ~x50 & ~x51 & ~x53 & ~x72 & ~x75 & ~x85 & ~x105 & ~x110 & ~x138 & ~x139 & ~x166 & ~x194 & ~x196 & ~x589 & ~x671 & ~x673 & ~x703 & ~x719 & ~x756 & ~x758 & ~x781;
assign c0178 =  x203 &  x425 & ~x14 & ~x25 & ~x238 & ~x239 & ~x293 & ~x295 & ~x364 & ~x463 & ~x751;
assign c0180 =  x232 &  x446 & ~x12 & ~x40 & ~x99 & ~x158 & ~x193 & ~x296 & ~x321;
assign c0182 = ~x7 & ~x19 & ~x42 & ~x57 & ~x129 & ~x219 & ~x266 & ~x328 & ~x617 & ~x619 & ~x645 & ~x655 & ~x656 & ~x749;
assign c0184 =  x167 & ~x299;
assign c0186 =  x115 &  x397 & ~x208 & ~x255 & ~x702;
assign c0188 = ~x61 & ~x154 & ~x252 & ~x318 & ~x328 & ~x382 & ~x388 & ~x415 & ~x420 & ~x497 & ~x741;
assign c0190 = ~x56 & ~x69 & ~x111 & ~x129 & ~x156 & ~x157 & ~x183 & ~x188 & ~x212 & ~x213 & ~x240 & ~x241 & ~x274 & ~x337 & ~x435 & ~x476 & ~x532 & ~x616 & ~x668 & ~x700 & ~x724 & ~x728 & ~x741 & ~x756 & ~x767 & ~x779;
assign c0192 =  x206 &  x234 & ~x12 & ~x27 & ~x32 & ~x53 & ~x54 & ~x70 & ~x119 & ~x137 & ~x160 & ~x194 & ~x280 & ~x365 & ~x366 & ~x367 & ~x397 & ~x421 & ~x423 & ~x700;
assign c0194 = ~x37 & ~x94 & ~x143 & ~x218 & ~x243 & ~x501 & ~x527 & ~x641 & ~x643 & ~x663 & ~x680 & ~x774;
assign c0196 =  x521 & ~x28 & ~x45 & ~x47 & ~x49 & ~x51 & ~x60 & ~x62 & ~x69 & ~x76 & ~x88 & ~x89 & ~x109 & ~x138 & ~x166 & ~x307 & ~x393 & ~x421 & ~x424 & ~x643 & ~x696 & ~x702 & ~x724 & ~x733 & ~x752 & ~x753 & ~x763 & ~x773 & ~x782;
assign c0198 =  x122 & ~x27 & ~x40 & ~x127 & ~x155 & ~x156 & ~x168 & ~x297 & ~x325 & ~x338 & ~x657 & ~x719;
assign c0200 =  x481 & ~x209 & ~x237 & ~x294 & ~x319 & ~x331 & ~x347 & ~x349 & ~x364 & ~x374 & ~x375 & ~x391 & ~x459 & ~x547 & ~x574 & ~x632;
assign c0202 =  x402 &  x481 & ~x12 & ~x13 & ~x37 & ~x69 & ~x291 & ~x617 & ~x637 & ~x648 & ~x702;
assign c0204 = ~x180 & ~x209 & ~x251 & ~x265 & ~x302 & ~x332 & ~x334 & ~x346 & ~x348 & ~x349 & ~x374 & ~x407 & ~x433 & ~x462 & ~x487 & ~x603 & ~x767 & ~x768;
assign c0206 =  x205 &  x233 &  x262 &  x289 &  x317 & ~x2 & ~x12 & ~x13 & ~x14 & ~x26 & ~x27 & ~x29 & ~x40 & ~x58 & ~x60 & ~x70 & ~x81 & ~x82 & ~x86 & ~x110 & ~x112 & ~x113 & ~x140 & ~x164 & ~x167 & ~x168 & ~x224 & ~x251 & ~x309 & ~x338 & ~x339 & ~x669 & ~x672 & ~x701 & ~x706 & ~x746 & ~x756 & ~x773;
assign c0208 =  x502 & ~x12 & ~x40 & ~x124 & ~x183 & ~x303 & ~x332 & ~x377 & ~x393;
assign c0210 =  x437 & ~x6 & ~x22 & ~x53 & ~x140 & ~x517 & ~x622 & ~x639 & ~x644 & ~x648 & ~x715 & ~x728 & ~x734;
assign c0212 =  x121 & ~x76 & ~x98 & ~x213 & ~x325 & ~x326 & ~x462 & ~x560 & ~x745 & ~x746;
assign c0214 =  x543 & ~x2 & ~x6 & ~x12 & ~x31 & ~x34 & ~x41 & ~x47 & ~x126 & ~x144 & ~x307 & ~x394 & ~x420 & ~x449 & ~x752 & ~x754 & ~x764 & ~x767 & ~x776 & ~x780 & ~x781;
assign c0216 = ~x125 & ~x246 & ~x328 & ~x365 & ~x366 & ~x393 & ~x394 & ~x542 & ~x664 & ~x754;
assign c0218 =  x460 &  x510 & ~x268 & ~x353 & ~x770;
assign c0220 =  x202 &  x260 &  x426 & ~x135 & ~x309 & ~x579 & ~x642 & ~x728;
assign c0222 =  x203 &  x259 &  x415 & ~x12 & ~x96 & ~x609 & ~x612 & ~x640 & ~x747 & ~x748;
assign c0224 =  x481 &  x484 & ~x6 & ~x12 & ~x13 & ~x14 & ~x82 & ~x106 & ~x153 & ~x392 & ~x448 & ~x588 & ~x667 & ~x668 & ~x726 & ~x755 & ~x774;
assign c0226 = ~x0 & ~x2 & ~x25 & ~x54 & ~x55 & ~x69 & ~x98 & ~x183 & ~x309 & ~x476 & ~x501 & ~x504 & ~x523 & ~x529 & ~x530 & ~x531 & ~x550 & ~x557 & ~x587 & ~x592 & ~x603 & ~x639 & ~x657 & ~x695 & ~x701 & ~x712 & ~x760;
assign c0228 =  x547 & ~x1 & ~x11 & ~x33 & ~x44 & ~x56 & ~x70 & ~x76 & ~x99 & ~x102 & ~x106 & ~x108 & ~x140 & ~x195 & ~x420 & ~x421 & ~x424 & ~x449 & ~x450 & ~x477 & ~x697 & ~x717 & ~x724 & ~x725 & ~x735 & ~x756 & ~x760 & ~x782;
assign c0230 =  x261 &  x509 & ~x27 & ~x40 & ~x72 & ~x321 & ~x368 & ~x394 & ~x396 & ~x420 & ~x421 & ~x451 & ~x477 & ~x698 & ~x699 & ~x714 & ~x728 & ~x759;
assign c0232 =  x205 &  x233 & ~x11 & ~x40 & ~x53 & ~x63 & ~x125 & ~x126 & ~x165 & ~x210 & ~x251 & ~x336 & ~x391 & ~x420 & ~x671 & ~x753 & ~x754 & ~x760;
assign c0234 =  x313 &  x454 & ~x152 & ~x153 & ~x161 & ~x347 & ~x586 & ~x744 & ~x747 & ~x783;
assign c0236 =  x194 & ~x71 & ~x185 & ~x213 & ~x243;
assign c0238 =  x434 &  x465 &  x520 & ~x124 & ~x743;
assign c0240 =  x231 &  x259 &  x287 &  x455 & ~x4 & ~x10 & ~x11 & ~x22 & ~x41 & ~x47 & ~x49 & ~x68 & ~x124 & ~x152 & ~x180 & ~x181 & ~x208 & ~x448 & ~x691 & ~x701 & ~x719 & ~x731 & ~x732 & ~x744 & ~x754 & ~x756 & ~x770 & ~x772 & ~x776 & ~x778 & ~x781 & ~x782;
assign c0242 =  x259 &  x483 & ~x11 & ~x31 & ~x41 & ~x84 & ~x322 & ~x325 & ~x357 & ~x530 & ~x532 & ~x559 & ~x727 & ~x738 & ~x755 & ~x775;
assign c0244 = ~x13 & ~x39 & ~x47 & ~x48 & ~x97 & ~x135 & ~x168 & ~x192 & ~x207 & ~x337 & ~x587 & ~x594 & ~x617 & ~x623 & ~x626 & ~x665 & ~x675 & ~x680 & ~x692 & ~x698 & ~x719 & ~x726 & ~x729 & ~x730 & ~x737 & ~x755 & ~x760 & ~x769;
assign c0246 =  x484 &  x485 &  x487 & ~x43 & ~x242 & ~x324 & ~x380 & ~x382 & ~x666;
assign c0248 =  x592 & ~x10 & ~x122 & ~x239 & ~x294 & ~x345 & ~x346 & ~x696 & ~x744 & ~x745 & ~x781;
assign c0250 =  x575 & ~x16 & ~x29 & ~x37 & ~x49 & ~x50 & ~x61 & ~x77 & ~x133 & ~x138 & ~x164 & ~x204 & ~x226 & ~x307 & ~x421 & ~x477 & ~x698 & ~x753 & ~x760 & ~x762 & ~x780;
assign c0252 =  x92 &  x232 &  x288 &  x343 & ~x3 & ~x13 & ~x14 & ~x25 & ~x111 & ~x311 & ~x366 & ~x671 & ~x676 & ~x677;
assign c0254 = ~x3 & ~x15 & ~x28 & ~x129 & ~x211 & ~x212 & ~x223 & ~x272 & ~x332 & ~x351 & ~x643 & ~x658 & ~x675 & ~x703 & ~x711 & ~x724 & ~x750 & ~x751 & ~x756 & ~x765 & ~x778 & ~x779;
assign c0256 =  x166 & ~x37 & ~x122 & ~x245 & ~x419;
assign c0258 = ~x21 & ~x56 & ~x130 & ~x327 & ~x337 & ~x356 & ~x475 & ~x476 & ~x529 & ~x586 & ~x602 & ~x655 & ~x694 & ~x701 & ~x702 & ~x703 & ~x705 & ~x733 & ~x752 & ~x757 & ~x759 & ~x778 & ~x781 & ~x783;
assign c0260 =  x149 &  x204 &  x475 & ~x51 & ~x365 & ~x366;
assign c0262 = ~x2 & ~x10 & ~x32 & ~x48 & ~x60 & ~x63 & ~x74 & ~x77 & ~x78 & ~x85 & ~x91 & ~x116 & ~x142 & ~x273 & ~x423 & ~x427 & ~x449 & ~x451 & ~x724 & ~x729 & ~x735 & ~x780;
assign c0264 = ~x30 & ~x163 & ~x170 & ~x172 & ~x184 & ~x351 & ~x454 & ~x479 & ~x702 & ~x745 & ~x772;
assign c0266 = ~x40 & ~x124 & ~x180 & ~x208 & ~x295 & ~x322 & ~x329 & ~x346 & ~x364 & ~x391 & ~x616 & ~x700 & ~x724;
assign c0268 =  x261 & ~x4 & ~x13 & ~x30 & ~x42 & ~x161 & ~x162 & ~x163 & ~x164 & ~x166 & ~x190 & ~x195 & ~x219 & ~x324 & ~x353 & ~x410 & ~x412 & ~x437 & ~x467 & ~x673 & ~x704 & ~x727 & ~x732 & ~x783;
assign c0270 =  x168;
assign c0272 =  x373 &  x457 &  x484 & ~x0 & ~x1 & ~x8 & ~x24 & ~x30 & ~x58 & ~x84 & ~x86 & ~x321 & ~x330 & ~x392 & ~x448 & ~x449 & ~x559 & ~x587 & ~x614 & ~x669 & ~x700 & ~x701 & ~x726 & ~x727 & ~x728 & ~x762 & ~x768 & ~x780;
assign c0274 =  x35 &  x480;
assign c0276 = ~x69 & ~x70 & ~x88 & ~x107 & ~x115 & ~x117 & ~x118 & ~x128 & ~x135 & ~x140 & ~x336 & ~x367 & ~x378 & ~x394 & ~x395 & ~x396 & ~x423 & ~x442 & ~x476 & ~x696 & ~x754 & ~x760 & ~x762;
assign c0278 =  x264 & ~x50 & ~x70 & ~x197 & ~x351 & ~x366 & ~x398 & ~x422 & ~x423 & ~x480 & ~x669 & ~x750 & ~x779;
assign c0280 =  x149 &  x316 &  x345 &  x346 &  x401 & ~x167 & ~x182 & ~x561;
assign c0282 =  x120 &  x232 &  x260 &  x315 &  x399 & ~x252 & ~x281 & ~x575 & ~x587 & ~x631 & ~x641 & ~x670 & ~x672 & ~x674 & ~x684 & ~x703 & ~x712;
assign c0284 = ~x82 & ~x128 & ~x154 & ~x168 & ~x266 & ~x328 & ~x502 & ~x530 & ~x571 & ~x628 & ~x645 & ~x701 & ~x703 & ~x725 & ~x751;
assign c0286 = ~x33 & ~x154 & ~x182 & ~x213 & ~x237 & ~x281 & ~x329 & ~x375 & ~x376 & ~x377 & ~x408 & ~x492 & ~x519 & ~x697 & ~x701 & ~x729;
assign c0288 =  x288 &  x315 &  x458 & ~x39 & ~x46 & ~x52 & ~x54 & ~x184 & ~x325 & ~x420 & ~x698;
assign c0290 =  x344 &  x680 & ~x295 & ~x376 & ~x393 & ~x766;
assign c0292 =  x207 & ~x12 & ~x15 & ~x41 & ~x71 & ~x98 & ~x107 & ~x109 & ~x127 & ~x157 & ~x352 & ~x364 & ~x392 & ~x423 & ~x448 & ~x731 & ~x765;
assign c0294 =  x234 &  x262 &  x289 & ~x0 & ~x12 & ~x13 & ~x16 & ~x22 & ~x25 & ~x42 & ~x44 & ~x45 & ~x52 & ~x68 & ~x72 & ~x137 & ~x268 & ~x307 & ~x420 & ~x424 & ~x699 & ~x726 & ~x727 & ~x745 & ~x773 & ~x781;
assign c0296 =  x119 &  x147 &  x423 &  x425 & ~x208 & ~x704 & ~x722 & ~x752;
assign c0298 = ~x27 & ~x83 & ~x112 & ~x161 & ~x166 & ~x220 & ~x221 & ~x380 & ~x467 & ~x589 & ~x632 & ~x640 & ~x647 & ~x676 & ~x683 & ~x694 & ~x695 & ~x700 & ~x722 & ~x725 & ~x739;
assign c0300 = ~x124 & ~x151 & ~x179 & ~x215 & ~x240 & ~x272 & ~x336 & ~x447 & ~x476 & ~x489 & ~x502 & ~x529 & ~x588 & ~x612 & ~x646 & ~x647 & ~x670 & ~x695 & ~x707 & ~x723 & ~x724 & ~x726 & ~x730;
assign c0302 =  x256 &  x257 &  x508 & ~x25 & ~x47 & ~x70 & ~x71 & ~x295 & ~x393 & ~x724 & ~x730;
assign c0304 =  x514 & ~x4 & ~x14 & ~x15 & ~x16 & ~x41 & ~x43 & ~x48 & ~x53 & ~x76 & ~x108 & ~x128 & ~x135 & ~x325 & ~x352 & ~x384 & ~x413 & ~x639 & ~x696 & ~x756 & ~x775;
assign c0306 =  x427 & ~x336 & ~x476 & ~x486 & ~x532 & ~x585 & ~x588 & ~x615 & ~x645 & ~x653 & ~x668 & ~x691 & ~x718 & ~x719 & ~x720 & ~x742 & ~x752 & ~x756;
assign c0308 =  x431 &  x510 & ~x28 & ~x43 & ~x111 & ~x322 & ~x330 & ~x586 & ~x637 & ~x642 & ~x700 & ~x703 & ~x739;
assign c0310 = ~x4 & ~x15 & ~x16 & ~x20 & ~x22 & ~x30 & ~x41 & ~x43 & ~x44 & ~x51 & ~x55 & ~x56 & ~x57 & ~x72 & ~x73 & ~x100 & ~x102 & ~x106 & ~x113 & ~x128 & ~x136 & ~x223 & ~x246 & ~x251 & ~x279 & ~x448 & ~x504 & ~x559 & ~x614 & ~x615 & ~x644 & ~x645 & ~x646 & ~x654 & ~x655 & ~x665 & ~x667 & ~x670 & ~x675 & ~x681 & ~x699 & ~x706 & ~x716 & ~x718 & ~x721 & ~x727 & ~x730 & ~x742 & ~x745 & ~x748 & ~x753 & ~x758 & ~x760 & ~x763 & ~x771 & ~x772 & ~x774 & ~x782;
assign c0312 = ~x13 & ~x25 & ~x31 & ~x42 & ~x80 & ~x99 & ~x110 & ~x132 & ~x133 & ~x160 & ~x188 & ~x196 & ~x279 & ~x364 & ~x406 & ~x466 & ~x507 & ~x670 & ~x737 & ~x756;
assign c0314 =  x506 & ~x153 & ~x346 & ~x708 & ~x730;
assign c0316 =  x90 &  x147 &  x342 & ~x135 & ~x300 & ~x325 & ~x410;
assign c0318 =  x495 & ~x181 & ~x237 & ~x238 & ~x270 & ~x695 & ~x722 & ~x734 & ~x742 & ~x743 & ~x751 & ~x754 & ~x761;
assign c0320 =  x146 &  x174 &  x426 & ~x0 & ~x11 & ~x13 & ~x14 & ~x23 & ~x41 & ~x55 & ~x187 & ~x224 & ~x309 & ~x337 & ~x588 & ~x643 & ~x671 & ~x702 & ~x725 & ~x728 & ~x749 & ~x750 & ~x765 & ~x778;
assign c0322 =  x439 &  x510 & ~x154 & ~x181 & ~x394 & ~x708 & ~x709 & ~x741;
assign c0324 =  x434 &  x480 & ~x12 & ~x46 & ~x266 & ~x676 & ~x703 & ~x744 & ~x766;
assign c0326 = ~x32 & ~x163 & ~x195 & ~x220 & ~x392 & ~x468 & ~x579 & ~x615 & ~x646 & ~x689 & ~x693 & ~x707 & ~x708 & ~x723 & ~x728 & ~x732 & ~x736 & ~x746 & ~x770;
assign c0328 =  x261 &  x289 &  x317 &  x485 & ~x5 & ~x8 & ~x33 & ~x73 & ~x78 & ~x81 & ~x99 & ~x125 & ~x141 & ~x153 & ~x196 & ~x392 & ~x674 & ~x694 & ~x707 & ~x722 & ~x733 & ~x752 & ~x774 & ~x780;
assign c0330 =  x94 &  x233 &  x372 & ~x199 & ~x200 & ~x548 & ~x589;
assign c0332 =  x507 & ~x4 & ~x54 & ~x69 & ~x99 & ~x100 & ~x211 & ~x304 & ~x320 & ~x364 & ~x394 & ~x703 & ~x737 & ~x738 & ~x783;
assign c0334 = ~x30 & ~x52 & ~x53 & ~x77 & ~x167 & ~x194 & ~x223 & ~x269 & ~x351 & ~x356 & ~x382 & ~x436 & ~x441 & ~x492 & ~x493 & ~x494 & ~x587 & ~x643 & ~x671 & ~x696 & ~x749 & ~x760 & ~x780;
assign c0336 =  x147 &  x203 &  x426 & ~x24 & ~x27 & ~x38 & ~x69 & ~x112 & ~x139 & ~x140 & ~x154 & ~x224 & ~x294 & ~x296 & ~x421 & ~x723 & ~x729 & ~x730 & ~x752 & ~x753 & ~x757 & ~x780 & ~x781;
assign c0338 =  x145 &  x174 &  x478 &  x480 &  x481 &  x508 & ~x9 & ~x730;
assign c0340 =  x399 & ~x29 & ~x56 & ~x235 & ~x236 & ~x291 & ~x609 & ~x613 & ~x614 & ~x634 & ~x717;
assign c0342 =  x259 &  x281 &  x315 & ~x228;
assign c0344 =  x479 & ~x13 & ~x23 & ~x38 & ~x178 & ~x273 & ~x289 & ~x557 & ~x560 & ~x652 & ~x664 & ~x696 & ~x729;
assign c0346 =  x262 & ~x3 & ~x5 & ~x50 & ~x63 & ~x80 & ~x100 & ~x101 & ~x129 & ~x131 & ~x157 & ~x158 & ~x159 & ~x162 & ~x192 & ~x199 & ~x224 & ~x226 & ~x280 & ~x392 & ~x421 & ~x673 & ~x697 & ~x752 & ~x763 & ~x767 & ~x773 & ~x774;
assign c0348 =  x202 &  x230 &  x454 & ~x5 & ~x24 & ~x47 & ~x150 & ~x180 & ~x373 & ~x392 & ~x732 & ~x755 & ~x770;
assign c0350 =  x206 & ~x24 & ~x41 & ~x57 & ~x80 & ~x86 & ~x97 & ~x110 & ~x114 & ~x129 & ~x130 & ~x155 & ~x252 & ~x336 & ~x365 & ~x369 & ~x392 & ~x448 & ~x560 & ~x697 & ~x716 & ~x738;
assign c0352 =  x223;
assign c0354 =  x173 & ~x1 & ~x8 & ~x13 & ~x15 & ~x28 & ~x40 & ~x42 & ~x49 & ~x82 & ~x83 & ~x610 & ~x643 & ~x645 & ~x665 & ~x700 & ~x723 & ~x739 & ~x747 & ~x748 & ~x755 & ~x772;
assign c0356 = ~x17 & ~x36 & ~x61 & ~x83 & ~x84 & ~x110 & ~x113 & ~x121 & ~x122 & ~x246 & ~x393 & ~x477 & ~x532 & ~x560 & ~x586 & ~x665 & ~x703 & ~x722 & ~x726 & ~x737 & ~x741 & ~x746 & ~x760;
assign c0358 =  x227 & ~x1 & ~x26 & ~x29 & ~x38 & ~x39 & ~x55 & ~x57 & ~x95 & ~x159 & ~x280 & ~x338 & ~x365 & ~x702 & ~x703 & ~x730 & ~x731 & ~x759 & ~x764 & ~x766 & ~x776 & ~x780;
assign c0360 =  x111;
assign c0362 =  x229 &  x230 &  x479 &  x480 &  x508 & ~x243 & ~x643 & ~x730 & ~x753 & ~x759;
assign c0364 = ~x0 & ~x13 & ~x47 & ~x210 & ~x269 & ~x278 & ~x295 & ~x323 & ~x439 & ~x653 & ~x680 & ~x681 & ~x693 & ~x700 & ~x703 & ~x725 & ~x728 & ~x731 & ~x746 & ~x764;
assign c0366 =  x458 &  x578 &  x632 & ~x40 & ~x70 & ~x153;
assign c0368 =  x257 & ~x13 & ~x44 & ~x66 & ~x365 & ~x556 & ~x609 & ~x615 & ~x638 & ~x647 & ~x668 & ~x669 & ~x693 & ~x699 & ~x707 & ~x723 & ~x760 & ~x774 & ~x775 & ~x777 & ~x783;
assign c0370 =  x648 & ~x10 & ~x12 & ~x186 & ~x216 & ~x240 & ~x268 & ~x352 & ~x671 & ~x728 & ~x751 & ~x754 & ~x763 & ~x780;
assign c0372 =  x53;
assign c0374 = ~x12 & ~x19 & ~x21 & ~x73 & ~x213 & ~x228 & ~x350 & ~x420 & ~x435 & ~x450 & ~x723 & ~x749 & ~x777 & ~x778 & ~x782;
assign c0376 = ~x9 & ~x30 & ~x36 & ~x39 & ~x93 & ~x113 & ~x122 & ~x141 & ~x145 & ~x172 & ~x235 & ~x247 & ~x291 & ~x292 & ~x319 & ~x477 & ~x615 & ~x690 & ~x724 & ~x726 & ~x744;
assign c0378 =  x403 &  x483 & ~x1 & ~x21 & ~x43 & ~x46 & ~x308 & ~x447 & ~x559 & ~x584 & ~x587 & ~x616 & ~x639 & ~x643 & ~x665 & ~x668 & ~x692 & ~x695 & ~x696 & ~x701 & ~x744;
assign c0380 =  x342 & ~x13 & ~x21 & ~x48 & ~x247 & ~x263 & ~x393 & ~x587 & ~x616 & ~x671 & ~x694 & ~x729 & ~x737 & ~x780;
assign c0382 =  x458 & ~x16 & ~x20 & ~x30 & ~x46 & ~x55 & ~x66 & ~x73 & ~x77 & ~x97 & ~x101 & ~x141 & ~x182 & ~x349 & ~x393 & ~x641 & ~x668 & ~x692 & ~x722 & ~x729 & ~x740 & ~x746 & ~x757 & ~x782;
assign c0384 = ~x10 & ~x12 & ~x39 & ~x62 & ~x139 & ~x239 & ~x270 & ~x276 & ~x336 & ~x357 & ~x380 & ~x699 & ~x724 & ~x725 & ~x746 & ~x749 & ~x768 & ~x771 & ~x773 & ~x776;
assign c0386 =  x361 &  x389 &  x428 & ~x12 & ~x97 & ~x99 & ~x730;
assign c0388 =  x517 & ~x5 & ~x11 & ~x17 & ~x19 & ~x46 & ~x75 & ~x355 & ~x383 & ~x384 & ~x411 & ~x420 & ~x439 & ~x440 & ~x467 & ~x495 & ~x522 & ~x671 & ~x698 & ~x725 & ~x730 & ~x757 & ~x759 & ~x781 & ~x782 & ~x783;
assign c0390 =  x453 &  x601 & ~x28 & ~x605 & ~x633 & ~x659 & ~x688 & ~x715 & ~x726 & ~x766 & ~x768 & ~x770;
assign c0392 =  x591 & ~x13 & ~x15 & ~x41 & ~x44 & ~x45 & ~x46 & ~x100 & ~x102 & ~x128 & ~x129 & ~x157 & ~x321 & ~x322 & ~x348 & ~x393 & ~x420 & ~x421 & ~x448 & ~x449 & ~x476 & ~x504 & ~x643 & ~x669 & ~x724 & ~x767 & ~x771 & ~x782 & ~x783;
assign c0394 = ~x122 & ~x244 & ~x290 & ~x330 & ~x392 & ~x420 & ~x476 & ~x666 & ~x667 & ~x673 & ~x696 & ~x724 & ~x727 & ~x730 & ~x731 & ~x739 & ~x780 & ~x782;
assign c0396 =  x539 & ~x4 & ~x5 & ~x10 & ~x16 & ~x18 & ~x41 & ~x100 & ~x323 & ~x645 & ~x678 & ~x693 & ~x705 & ~x717 & ~x751 & ~x767 & ~x770;
assign c0398 =  x368 & ~x42 & ~x236 & ~x239 & ~x281 & ~x308 & ~x408 & ~x435 & ~x490 & ~x584 & ~x611 & ~x614 & ~x644 & ~x693;
assign c0400 =  x570 &  x593 &  x596 & ~x33 & ~x36 & ~x38 & ~x392 & ~x450 & ~x726 & ~x778;
assign c0402 =  x225 &  x479 &  x480;
assign c0404 =  x370 &  x433 &  x454 & ~x54 & ~x208 & ~x556 & ~x583 & ~x584 & ~x610 & ~x671 & ~x694 & ~x700 & ~x762 & ~x776;
assign c0406 =  x34 &  x508;
assign c0408 =  x319 &  x341 &  x458 & ~x184 & ~x211 & ~x268 & ~x269 & ~x500;
assign c0410 =  x313 &  x510 &  x536 & ~x6 & ~x11 & ~x21 & ~x70 & ~x108 & ~x393 & ~x423 & ~x424 & ~x742;
assign c0412 =  x231 & ~x68 & ~x127 & ~x210 & ~x266 & ~x292 & ~x656 & ~x731;
assign c0414 = ~x1 & ~x4 & ~x24 & ~x28 & ~x40 & ~x44 & ~x186 & ~x252 & ~x253 & ~x281 & ~x475 & ~x476 & ~x586 & ~x602 & ~x616 & ~x628 & ~x629 & ~x645 & ~x649 & ~x669 & ~x674 & ~x676 & ~x682 & ~x699 & ~x701 & ~x710 & ~x749 & ~x754;
assign c0416 = ~x31 & ~x52 & ~x74 & ~x219 & ~x494 & ~x531 & ~x557 & ~x560 & ~x577 & ~x587 & ~x615 & ~x639 & ~x642 & ~x655 & ~x699 & ~x709 & ~x723 & ~x762;
assign c0418 =  x428 &  x512 &  x568 &  x577 &  x625 & ~x422;
assign c0420 =  x379 &  x401 & ~x19 & ~x365 & ~x460 & ~x650 & ~x750;
assign c0422 =  x259 &  x454 &  x511 &  x546 & ~x6 & ~x20 & ~x393 & ~x670 & ~x748;
assign c0424 =  x539 &  x566 &  x567 &  x603 & ~x351 & ~x422 & ~x423 & ~x451;
assign c0426 =  x197 &  x508;
assign c0428 =  x233 &  x482 & ~x12 & ~x57 & ~x140 & ~x294 & ~x364 & ~x531 & ~x577 & ~x642 & ~x671 & ~x686 & ~x697;
assign c0430 =  x446 &  x483 &  x484 &  x547 & ~x7 & ~x12 & ~x14 & ~x693 & ~x695;
assign c0432 =  x261 &  x262 &  x263 &  x288 &  x317 &  x457 & ~x11 & ~x13 & ~x28 & ~x40 & ~x43 & ~x128 & ~x168 & ~x196 & ~x449 & ~x753 & ~x755;
assign c0434 =  x462 &  x463 &  x483 &  x511 &  x538 & ~x33 & ~x394 & ~x423 & ~x424 & ~x738 & ~x764;
assign c0436 =  x474 &  x602 &  x657 & ~x366 & ~x716;
assign c0438 = ~x40 & ~x42 & ~x98 & ~x153 & ~x243 & ~x244 & ~x245 & ~x434 & ~x472 & ~x532 & ~x607 & ~x674 & ~x686 & ~x752;
assign c0440 =  x202 & ~x16 & ~x20 & ~x28 & ~x38 & ~x46 & ~x65 & ~x74 & ~x301 & ~x309 & ~x615 & ~x644 & ~x700 & ~x703 & ~x704 & ~x731 & ~x748 & ~x757 & ~x764 & ~x765;
assign c0442 =  x205 &  x232 & ~x124 & ~x128 & ~x182 & ~x211 & ~x294 & ~x588 & ~x660;
assign c0444 =  x166 & ~x242;
assign c0446 =  x259 &  x536 & ~x26 & ~x40 & ~x41 & ~x66 & ~x94 & ~x95 & ~x98 & ~x153 & ~x586 & ~x702 & ~x767 & ~x781;
assign c0448 =  x143 &  x173 &  x174 &  x399 &  x452;
assign c0450 =  x205 & ~x12 & ~x55 & ~x294 & ~x306 & ~x308 & ~x340 & ~x393 & ~x548 & ~x603 & ~x711 & ~x729 & ~x767;
assign c0452 =  x260 & ~x3 & ~x13 & ~x57 & ~x311 & ~x321 & ~x330 & ~x476 & ~x602 & ~x685 & ~x686 & ~x704 & ~x711 & ~x739;
assign c0454 =  x148 & ~x109 & ~x136 & ~x164 & ~x208 & ~x264 & ~x364 & ~x652 & ~x653 & ~x654 & ~x694 & ~x709 & ~x730 & ~x731 & ~x751 & ~x756;
assign c0456 =  x31;
assign c0458 =  x543 &  x577 &  x605 & ~x6 & ~x9 & ~x14 & ~x42 & ~x57 & ~x196 & ~x392 & ~x451 & ~x752 & ~x753;
assign c0460 =  x230 & ~x5 & ~x21 & ~x37 & ~x42 & ~x54 & ~x126 & ~x139 & ~x237 & ~x249 & ~x614 & ~x670 & ~x673 & ~x682 & ~x703 & ~x707 & ~x727 & ~x752 & ~x762 & ~x772;
assign c0462 = ~x2 & ~x6 & ~x15 & ~x24 & ~x29 & ~x41 & ~x45 & ~x49 & ~x54 & ~x73 & ~x75 & ~x77 & ~x80 & ~x104 & ~x133 & ~x136 & ~x138 & ~x140 & ~x157 & ~x160 & ~x168 & ~x169 & ~x353 & ~x439 & ~x440 & ~x467 & ~x587 & ~x701 & ~x728 & ~x733 & ~x748 & ~x775 & ~x782;
assign c0464 =  x287 &  x315 &  x343 &  x455 &  x483 &  x511 &  x539 & ~x10 & ~x218 & ~x291 & ~x532 & ~x587 & ~x614 & ~x698 & ~x731 & ~x783;
assign c0466 =  x234 & ~x45 & ~x71 & ~x79 & ~x141 & ~x162 & ~x279 & ~x356 & ~x392 & ~x437 & ~x493 & ~x560 & ~x754 & ~x758 & ~x781;
assign c0468 =  x118 &  x333 &  x361 &  x453;
assign c0470 =  x455 & ~x25 & ~x83 & ~x209 & ~x265 & ~x308 & ~x556 & ~x660 & ~x665 & ~x708 & ~x714 & ~x736 & ~x752 & ~x760 & ~x761;
assign c0474 =  x313 &  x543 &  x566 &  x568;
assign c0476 =  x559 & ~x303;
assign c0478 =  x460 & ~x20 & ~x44 & ~x169 & ~x240 & ~x268 & ~x297 & ~x353 & ~x382 & ~x642 & ~x674 & ~x678 & ~x695 & ~x729 & ~x754;
assign c0480 =  x233 & ~x29 & ~x211 & ~x266 & ~x587 & ~x603 & ~x618 & ~x641 & ~x657 & ~x683 & ~x697 & ~x732 & ~x753;
assign c0482 = ~x8 & ~x27 & ~x40 & ~x158 & ~x191 & ~x220 & ~x224 & ~x322 & ~x376 & ~x380 & ~x409 & ~x413 & ~x464 & ~x466 & ~x496 & ~x754 & ~x755;
assign c0484 = ~x12 & ~x28 & ~x85 & ~x126 & ~x154 & ~x156 & ~x187 & ~x211 & ~x268 & ~x298 & ~x322 & ~x350 & ~x362 & ~x377 & ~x405 & ~x476 & ~x741 & ~x754 & ~x782;
assign c0486 =  x314 & ~x1 & ~x6 & ~x8 & ~x13 & ~x31 & ~x33 & ~x38 & ~x39 & ~x41 & ~x56 & ~x67 & ~x95 & ~x122 & ~x123 & ~x124 & ~x125 & ~x152 & ~x207 & ~x208 & ~x246 & ~x504 & ~x586 & ~x640 & ~x667 & ~x695 & ~x698 & ~x725 & ~x726 & ~x729 & ~x730 & ~x732 & ~x753 & ~x757 & ~x759 & ~x781 & ~x782 & ~x783;
assign c0488 =  x260 &  x345 &  x457 &  x485 &  x486 &  x625;
assign c0490 =  x593 & ~x11 & ~x21 & ~x28 & ~x45 & ~x47 & ~x213 & ~x224 & ~x280 & ~x378 & ~x379 & ~x387 & ~x450 & ~x696 & ~x775;
assign c0492 =  x229 &  x480 & ~x11 & ~x13 & ~x18 & ~x41 & ~x289 & ~x329 & ~x448 & ~x730 & ~x780;
assign c0494 = ~x140 & ~x181 & ~x210 & ~x237 & ~x263 & ~x290 & ~x294 & ~x319 & ~x348 & ~x351 & ~x374 & ~x404 & ~x419 & ~x432 & ~x475 & ~x504 & ~x604 & ~x659 & ~x728 & ~x781 & ~x782;
assign c0496 =  x147 &  x148 &  x176 & ~x1 & ~x18 & ~x27 & ~x56 & ~x181 & ~x584 & ~x623 & ~x649 & ~x691 & ~x701 & ~x703 & ~x718 & ~x727 & ~x730 & ~x756 & ~x778;
assign c0498 =  x63 &  x149 &  x261 &  x315 &  x343 & ~x394 & ~x421;
assign c01 =  x627 & ~x1 & ~x27 & ~x44 & ~x54 & ~x447 & ~x476 & ~x532 & ~x564 & ~x591 & ~x617 & ~x618 & ~x648 & ~x702 & ~x726 & ~x729 & ~x733 & ~x754 & ~x757 & ~x759 & ~x760;
assign c03 =  x241 &  x593 & ~x196 & ~x206 & ~x390;
assign c05 = ~x1 & ~x24 & ~x26 & ~x30 & ~x52 & ~x53 & ~x54 & ~x57 & ~x58 & ~x80 & ~x83 & ~x84 & ~x85 & ~x110 & ~x138 & ~x140 & ~x141 & ~x142 & ~x144 & ~x169 & ~x180 & ~x199 & ~x200 & ~x222 & ~x227 & ~x249 & ~x255 & ~x261 & ~x310 & ~x337 & ~x642 & ~x755 & ~x757 & ~x776;
assign c07 =  x572 &  x630 & ~x6 & ~x139 & ~x614 & ~x624 & ~x705 & ~x727 & ~x764;
assign c09 = ~x24 & ~x55 & ~x83 & ~x237 & ~x400 & ~x428 & ~x446 & ~x455 & ~x475 & ~x558 & ~x559 & ~x561 & ~x589 & ~x672 & ~x673 & ~x728 & ~x757 & ~x760 & ~x775;
assign c011 =  x699;
assign c013 = ~x208 & ~x398 & ~x399 & ~x453 & ~x480 & ~x535;
assign c015 =  x265 &  x266 & ~x194 & ~x597 & ~x652 & ~x664;
assign c017 =  x451 & ~x4 & ~x103 & ~x172 & ~x174 & ~x229 & ~x253 & ~x283;
assign c019 =  x405 & ~x7 & ~x417 & ~x503 & ~x522 & ~x607 & ~x730;
assign c021 = ~x155 & ~x180 & ~x341 & ~x396 & ~x474 & ~x480 & ~x497 & ~x524 & ~x525 & ~x559 & ~x590 & ~x646;
assign c023 =  x716 &  x717 & ~x258 & ~x782;
assign c025 =  x634 & ~x445 & ~x497 & ~x515 & ~x543;
assign c027 =  x211 &  x235 &  x236 & ~x529 & ~x551 & ~x607;
assign c029 =  x368 &  x423 & ~x82 & ~x142 & ~x168 & ~x197 & ~x253 & ~x509 & ~x537;
assign c031 =  x221 & ~x36 & ~x467 & ~x521 & ~x522;
assign c033 =  x118 & ~x398 & ~x643 & ~x727;
assign c035 = ~x32 & ~x58 & ~x61 & ~x88 & ~x89 & ~x113 & ~x114 & ~x144 & ~x147 & ~x174 & ~x193 & ~x228 & ~x254 & ~x255 & ~x284 & ~x312 & ~x623 & ~x705;
assign c037 =  x418 & ~x378 & ~x382 & ~x515 & ~x627;
assign c039 =  x669 & ~x531 & ~x559;
assign c041 = ~x113 & ~x177 & ~x232 & ~x376 & ~x459 & ~x515 & ~x626 & ~x655 & ~x683 & ~x710;
assign c043 =  x565 & ~x3 & ~x17 & ~x24 & ~x27 & ~x31 & ~x84 & ~x85 & ~x108 & ~x113 & ~x114 & ~x142 & ~x171 & ~x191 & ~x196 & ~x199 & ~x225 & ~x226 & ~x227 & ~x253 & ~x278 & ~x305 & ~x310 & ~x334 & ~x336 & ~x388 & ~x756;
assign c045 =  x574 &  x603 & ~x26 & ~x29 & ~x475 & ~x513 & ~x528 & ~x529 & ~x557 & ~x585 & ~x755;
assign c047 = ~x1 & ~x19 & ~x28 & ~x50 & ~x68 & ~x110 & ~x112 & ~x172 & ~x433 & ~x597 & ~x651 & ~x652 & ~x653 & ~x679 & ~x710 & ~x735;
assign c049 =  x325 &  x350 &  x486 & ~x24 & ~x78 & ~x139 & ~x140 & ~x168 & ~x615 & ~x757;
assign c051 = ~x50 & ~x78 & ~x393 & ~x421 & ~x463 & ~x489 & ~x515 & ~x544 & ~x547 & ~x601 & ~x602 & ~x631 & ~x661 & ~x716 & ~x731 & ~x772;
assign c053 = ~x18 & ~x114 & ~x118 & ~x139 & ~x141 & ~x168 & ~x197 & ~x198 & ~x378 & ~x432 & ~x487 & ~x514 & ~x542 & ~x571 & ~x599 & ~x735 & ~x736 & ~x761 & ~x777;
assign c055 =  x678 & ~x400 & ~x427;
assign c057 = ~x19 & ~x57 & ~x140 & ~x169 & ~x197 & ~x203 & ~x253 & ~x254 & ~x597 & ~x627 & ~x711 & ~x736 & ~x737 & ~x740 & ~x746 & ~x769 & ~x783;
assign c059 =  x323 &  x430 & ~x23 & ~x25 & ~x27 & ~x53 & ~x115 & ~x170 & ~x224 & ~x279 & ~x385 & ~x783;
assign c061 =  x297 &  x320 &  x402;
assign c063 =  x124 & ~x10 & ~x651 & ~x679;
assign c065 =  x125 &  x154 &  x207 & ~x2 & ~x503;
assign c067 =  x310;
assign c069 =  x453 & ~x43 & ~x107 & ~x178 & ~x349 & ~x377 & ~x393 & ~x460 & ~x487 & ~x570 & ~x710 & ~x761 & ~x770;
assign c071 =  x389 &  x416 & ~x26 & ~x61 & ~x379 & ~x380 & ~x381 & ~x434 & ~x651 & ~x682 & ~x753;
assign c073 =  x10 &  x37;
assign c075 = ~x292 & ~x294 & ~x479 & ~x483 & ~x531 & ~x534 & ~x557 & ~x558 & ~x585 & ~x612 & ~x757 & ~x761 & ~x776;
assign c077 =  x606 & ~x0 & ~x497 & ~x499 & ~x503 & ~x626;
assign c079 =  x433 & ~x26 & ~x131 & ~x184 & ~x453 & ~x502 & ~x530 & ~x531 & ~x549 & ~x559 & ~x754;
assign c081 = ~x55 & ~x151 & ~x260;
assign c083 =  x179 &  x338;
assign c085 =  x424 &  x451 & ~x0 & ~x1 & ~x3 & ~x24 & ~x26 & ~x31 & ~x33 & ~x51 & ~x52 & ~x53 & ~x54 & ~x58 & ~x61 & ~x79 & ~x82 & ~x85 & ~x89 & ~x107 & ~x109 & ~x113 & ~x137 & ~x138 & ~x139 & ~x141 & ~x143 & ~x167 & ~x168 & ~x169 & ~x170 & ~x172 & ~x197 & ~x198 & ~x252 & ~x253 & ~x281 & ~x336 & ~x672 & ~x697 & ~x726 & ~x727 & ~x751 & ~x752 & ~x781 & ~x783;
assign c087 =  x275 &  x303 &  x331 & ~x1 & ~x392 & ~x436 & ~x491 & ~x517 & ~x546 & ~x547 & ~x576 & ~x756 & ~x769;
assign c089 = ~x1 & ~x17 & ~x20 & ~x43 & ~x45 & ~x50 & ~x82 & ~x110 & ~x111 & ~x139 & ~x322 & ~x348 & ~x504 & ~x508 & ~x532 & ~x534 & ~x536 & ~x537 & ~x564 & ~x565 & ~x644 & ~x647 & ~x671 & ~x700;
assign c091 =  x658 & ~x43 & ~x56 & ~x183 & ~x302 & ~x305 & ~x419 & ~x589 & ~x615 & ~x616 & ~x701 & ~x730;
assign c093 =  x294 &  x296 &  x496;
assign c095 = ~x119 & ~x408 & ~x436 & ~x517 & ~x546 & ~x569 & ~x629 & ~x653 & ~x693;
assign c097 = ~x3 & ~x7 & ~x22 & ~x51 & ~x52 & ~x54 & ~x60 & ~x78 & ~x79 & ~x80 & ~x82 & ~x83 & ~x87 & ~x107 & ~x109 & ~x114 & ~x115 & ~x135 & ~x136 & ~x140 & ~x163 & ~x169 & ~x190 & ~x219 & ~x248 & ~x250 & ~x305 & ~x362 & ~x391 & ~x417 & ~x418 & ~x473 & ~x572 & ~x699 & ~x753 & ~x778;
assign c099 =  x675 & ~x627 & ~x628 & ~x658 & ~x659;
assign c0101 =  x546 &  x634 &  x662;
assign c0103 =  x358 &  x454 & ~x16 & ~x35 & ~x325 & ~x378 & ~x489 & ~x547;
assign c0105 = ~x7 & ~x58 & ~x90 & ~x452 & ~x508 & ~x509 & ~x564 & ~x594 & ~x621 & ~x650 & ~x733 & ~x772;
assign c0107 =  x152 &  x179 &  x312 & ~x28 & ~x223 & ~x225 & ~x252;
assign c0109 =  x67 &  x68 & ~x61 & ~x102;
assign c0111 =  x256 &  x283 &  x338 &  x339 & ~x1 & ~x26 & ~x27 & ~x83 & ~x85 & ~x280;
assign c0113 =  x243 & ~x19 & ~x380 & ~x525 & ~x526 & ~x569 & ~x654 & ~x736;
assign c0115 = ~x19 & ~x20 & ~x21 & ~x26 & ~x55 & ~x71 & ~x83 & ~x116 & ~x135 & ~x141 & ~x143 & ~x169 & ~x179 & ~x220 & ~x221 & ~x224 & ~x226 & ~x247 & ~x249 & ~x277 & ~x278 & ~x281 & ~x282 & ~x305 & ~x306 & ~x308 & ~x334 & ~x335 & ~x365 & ~x419 & ~x783;
assign c0117 =  x577 &  x580 & ~x109 & ~x279 & ~x474 & ~x502;
assign c0119 =  x154 &  x155 &  x181 & ~x54 & ~x81 & ~x112 & ~x139 & ~x166 & ~x196 & ~x642 & ~x747;
assign c0121 =  x406 & ~x98 & ~x180 & ~x295 & ~x427 & ~x482;
assign c0123 =  x212 & ~x55 & ~x260;
assign c0125 = ~x0 & ~x5 & ~x27 & ~x29 & ~x30 & ~x31 & ~x55 & ~x56 & ~x83 & ~x86 & ~x87 & ~x141 & ~x142 & ~x170 & ~x196 & ~x251 & ~x349 & ~x378 & ~x392 & ~x393 & ~x406 & ~x421 & ~x434 & ~x518 & ~x570 & ~x599 & ~x727 & ~x735 & ~x757;
assign c0127 =  x747 & ~x68;
assign c0129 = ~x24 & ~x249 & ~x274 & ~x276 & ~x302 & ~x304 & ~x331 & ~x332 & ~x334 & ~x365 & ~x388 & ~x389 & ~x392 & ~x414 & ~x441 & ~x443 & ~x611 & ~x612 & ~x614 & ~x640 & ~x671 & ~x726 & ~x761 & ~x783;
assign c0131 = ~x19 & ~x70 & ~x71 & ~x367 & ~x368 & ~x396 & ~x420 & ~x423 & ~x424 & ~x452 & ~x479 & ~x506 & ~x524 & ~x526 & ~x559 & ~x562 & ~x614 & ~x618 & ~x646 & ~x705 & ~x729 & ~x733 & ~x753;
assign c0133 =  x658 & ~x291 & ~x456 & ~x534 & ~x589 & ~x674;
assign c0135 =  x256 &  x283 &  x311 & ~x2 & ~x28 & ~x56 & ~x534 & ~x560 & ~x562 & ~x590 & ~x617 & ~x729 & ~x750 & ~x758 & ~x759;
assign c0137 =  x350 &  x594 & ~x55 & ~x473 & ~x502 & ~x533 & ~x561;
assign c0139 = ~x6 & ~x20 & ~x58 & ~x117 & ~x152 & ~x179 & ~x190 & ~x193 & ~x252 & ~x254 & ~x279 & ~x282 & ~x339 & ~x576 & ~x610 & ~x639 & ~x761;
assign c0141 =  x352 & ~x267 & ~x480 & ~x534 & ~x563 & ~x590;
assign c0143 = ~x36 & ~x60 & ~x90 & ~x114 & ~x169 & ~x197 & ~x511 & ~x542 & ~x571 & ~x655 & ~x676 & ~x685;
assign c0145 =  x208 & ~x348 & ~x374 & ~x403;
assign c0147 = ~x27 & ~x51 & ~x99 & ~x160 & ~x452 & ~x453 & ~x508 & ~x534 & ~x562 & ~x611 & ~x640 & ~x644 & ~x730 & ~x753 & ~x766 & ~x770;
assign c0149 = ~x6 & ~x35 & ~x61 & ~x91 & ~x138 & ~x173 & ~x174 & ~x351 & ~x353 & ~x406 & ~x460 & ~x544 & ~x545 & ~x665 & ~x761;
assign c0151 =  x602 & ~x1 & ~x43 & ~x44 & ~x537 & ~x591 & ~x592 & ~x702 & ~x750 & ~x769;
assign c0153 =  x11 & ~x225;
assign c0155 = ~x1 & ~x5 & ~x15 & ~x106 & ~x138 & ~x407 & ~x436 & ~x542 & ~x570 & ~x626 & ~x627 & ~x633 & ~x654 & ~x657 & ~x659 & ~x660 & ~x718 & ~x736 & ~x739 & ~x761 & ~x762 & ~x769 & ~x777;
assign c0157 = ~x28 & ~x36 & ~x64 & ~x91 & ~x194 & ~x282 & ~x411 & ~x420 & ~x438 & ~x489 & ~x516 & ~x546 & ~x631 & ~x747;
assign c0159 = ~x26 & ~x168 & ~x337 & ~x764;
assign c0161 =  x41 & ~x72 & ~x782;
assign c0163 = ~x5 & ~x28 & ~x54 & ~x79 & ~x149 & ~x366 & ~x421 & ~x518 & ~x542 & ~x544 & ~x545 & ~x546 & ~x547 & ~x549 & ~x576 & ~x735 & ~x763 & ~x764;
assign c0165 = ~x19 & ~x22 & ~x34 & ~x35 & ~x70 & ~x79 & ~x136 & ~x366 & ~x407 & ~x488 & ~x516 & ~x518 & ~x572 & ~x600 & ~x602 & ~x668 & ~x687 & ~x765 & ~x777 & ~x778;
assign c0167 =  x240 &  x367 & ~x140 & ~x196;
assign c0169 =  x91 & ~x23 & ~x51 & ~x304 & ~x444 & ~x445 & ~x471 & ~x472 & ~x501 & ~x505 & ~x506;
assign c0171 = ~x85 & ~x354 & ~x379 & ~x432 & ~x436 & ~x458 & ~x459 & ~x545 & ~x595 & ~x624 & ~x649 & ~x762;
assign c0173 = ~x260 & ~x628 & ~x656;
assign c0175 = ~x6 & ~x28 & ~x29 & ~x30 & ~x51 & ~x52 & ~x71 & ~x79 & ~x99 & ~x107 & ~x109 & ~x114 & ~x136 & ~x138 & ~x139 & ~x164 & ~x170 & ~x191 & ~x197 & ~x220 & ~x248 & ~x250 & ~x251 & ~x291 & ~x391 & ~x401 & ~x699 & ~x726 & ~x776;
assign c0177 = ~x30 & ~x34 & ~x59 & ~x86 & ~x143 & ~x144 & ~x195 & ~x596 & ~x726;
assign c0179 =  x301 &  x329 & ~x28 & ~x31 & ~x57 & ~x438 & ~x463 & ~x627 & ~x683;
assign c0181 =  x183 & ~x28 & ~x44 & ~x351 & ~x461 & ~x711;
assign c0183 =  x575 & ~x157 & ~x184 & ~x290 & ~x507 & ~x535 & ~x557 & ~x558 & ~x644 & ~x645;
assign c0185 = ~x3 & ~x8 & ~x27 & ~x29 & ~x34 & ~x39 & ~x42 & ~x50 & ~x60 & ~x81 & ~x89 & ~x105 & ~x131 & ~x145 & ~x169 & ~x226 & ~x227 & ~x254 & ~x569 & ~x597 & ~x598 & ~x626 & ~x655 & ~x707 & ~x708 & ~x744 & ~x761 & ~x766 & ~x767 & ~x773;
assign c0187 = ~x2 & ~x13 & ~x16 & ~x18 & ~x22 & ~x28 & ~x29 & ~x42 & ~x65 & ~x82 & ~x110 & ~x113 & ~x139 & ~x141 & ~x143 & ~x169 & ~x171 & ~x198 & ~x226 & ~x253 & ~x281 & ~x282 & ~x308 & ~x571 & ~x598 & ~x599 & ~x600 & ~x626 & ~x656 & ~x681 & ~x684;
assign c0189 =  x306 & ~x451 & ~x509;
assign c0191 = ~x15 & ~x247 & ~x249 & ~x274 & ~x301 & ~x307 & ~x391 & ~x419 & ~x443 & ~x472 & ~x473 & ~x498 & ~x587 & ~x668 & ~x698 & ~x731;
assign c0193 = ~x10 & ~x147 & ~x167 & ~x177 & ~x339 & ~x381 & ~x544 & ~x545 & ~x603;
assign c0195 = ~x1 & ~x7 & ~x52 & ~x55 & ~x76 & ~x89 & ~x106 & ~x117 & ~x143 & ~x144 & ~x167 & ~x511 & ~x539 & ~x565 & ~x593 & ~x594 & ~x620 & ~x621 & ~x622 & ~x652 & ~x674 & ~x675 & ~x680 & ~x681 & ~x703 & ~x712 & ~x737 & ~x738 & ~x739 & ~x760;
assign c0197 =  x207 & ~x24 & ~x49 & ~x55 & ~x107 & ~x202 & ~x503 & ~x586 & ~x722 & ~x753 & ~x782;
assign c0199 =  x399 & ~x25 & ~x47 & ~x72 & ~x104 & ~x114 & ~x135 & ~x220 & ~x279 & ~x331 & ~x446 & ~x504 & ~x698;
assign c0201 =  x455 & ~x19 & ~x28 & ~x36 & ~x55 & ~x112 & ~x407 & ~x436 & ~x464 & ~x570 & ~x599 & ~x627 & ~x655 & ~x682 & ~x710 & ~x727 & ~x765 & ~x767 & ~x783;
assign c0203 =  x454 & ~x22 & ~x31 & ~x32 & ~x82 & ~x83 & ~x86 & ~x107 & ~x164 & ~x172 & ~x192 & ~x225 & ~x248 & ~x254 & ~x276 & ~x281 & ~x388 & ~x417 & ~x419;
assign c0205 =  x268 &  x269 & ~x26 & ~x289 & ~x531 & ~x710;
assign c0207 =  x303 & ~x460 & ~x462 & ~x463 & ~x464 & ~x520 & ~x576 & ~x600 & ~x658 & ~x684;
assign c0209 =  x399 &  x454 & ~x10 & ~x82 & ~x136 & ~x433 & ~x435 & ~x462 & ~x464 & ~x516 & ~x518 & ~x705 & ~x736 & ~x771 & ~x783;
assign c0211 =  x353 & ~x16 & ~x335 & ~x361 & ~x362 & ~x413 & ~x417 & ~x441;
assign c0213 =  x648 & ~x561 & ~x570 & ~x627 & ~x736 & ~x762;
assign c0215 = ~x167 & ~x188 & ~x237 & ~x400 & ~x453 & ~x482 & ~x531 & ~x532 & ~x724;
assign c0217 = ~x0 & ~x1 & ~x47 & ~x106 & ~x180 & ~x399 & ~x426 & ~x453 & ~x454 & ~x509 & ~x729 & ~x731 & ~x755 & ~x757 & ~x778 & ~x783;
assign c0219 =  x208 &  x315 & ~x9 & ~x512 & ~x541 & ~x596 & ~x624 & ~x625 & ~x652;
assign c0221 =  x215 & ~x27 & ~x59 & ~x231 & ~x461;
assign c0223 =  x236 &  x342 & ~x625 & ~x683;
assign c0225 =  x153 &  x398 & ~x6 & ~x56 & ~x110 & ~x140 & ~x144 & ~x167 & ~x170 & ~x223 & ~x225 & ~x252 & ~x749 & ~x779;
assign c0227 =  x724;
assign c0229 =  x295 & ~x40 & ~x126 & ~x127 & ~x279 & ~x333 & ~x391 & ~x502 & ~x783;
assign c0231 =  x265 &  x292 & ~x569 & ~x597 & ~x652 & ~x654;
assign c0233 = ~x470 & ~x498 & ~x525 & ~x554;
assign c0235 = ~x27 & ~x36 & ~x79 & ~x96 & ~x110 & ~x408 & ~x491 & ~x515 & ~x517 & ~x544 & ~x546 & ~x548 & ~x571 & ~x599 & ~x602 & ~x603 & ~x630 & ~x742 & ~x756 & ~x765;
assign c0237 =  x175 & ~x27 & ~x395 & ~x396 & ~x397 & ~x425 & ~x477 & ~x479 & ~x503 & ~x505 & ~x531 & ~x536 & ~x586 & ~x588 & ~x616 & ~x618 & ~x646 & ~x647 & ~x671 & ~x700 & ~x702;
assign c0239 = ~x4 & ~x308 & ~x348 & ~x375 & ~x376 & ~x384 & ~x404 & ~x433 & ~x459 & ~x541 & ~x676 & ~x678 & ~x679 & ~x707 & ~x727;
assign c0241 = ~x26 & ~x139 & ~x324 & ~x336 & ~x379 & ~x382 & ~x383 & ~x411 & ~x433 & ~x438 & ~x439 & ~x464 & ~x466 & ~x493 & ~x516 & ~x517 & ~x518 & ~x521 & ~x522 & ~x656 & ~x727 & ~x769 & ~x776 & ~x783;
assign c0243 =  x706 & ~x53 & ~x135 & ~x142 & ~x160 & ~x227 & ~x418 & ~x446;
assign c0245 = ~x0 & ~x21 & ~x75 & ~x84 & ~x134 & ~x136 & ~x191 & ~x211 & ~x250 & ~x277 & ~x306 & ~x402 & ~x419 & ~x446 & ~x591 & ~x646 & ~x701 & ~x730;
assign c0247 =  x365 &  x393 &  x394;
assign c0249 =  x65 & ~x30 & ~x123;
assign c0251 =  x70 & ~x734;
assign c0253 = ~x52 & ~x84 & ~x111 & ~x112 & ~x182 & ~x280 & ~x304 & ~x305 & ~x306 & ~x307 & ~x359 & ~x360 & ~x362 & ~x384 & ~x388 & ~x416 & ~x417 & ~x418 & ~x439 & ~x502 & ~x556 & ~x587 & ~x613 & ~x643;
assign c0255 =  x633 & ~x496 & ~x502 & ~x715;
assign c0257 =  x687 & ~x447 & ~x500 & ~x523 & ~x525 & ~x526 & ~x581 & ~x607 & ~x611;
assign c0259 =  x398 &  x452 & ~x44 & ~x166 & ~x414 & ~x460 & ~x469;
assign c0261 = ~x0 & ~x17 & ~x19 & ~x44 & ~x55 & ~x59 & ~x60 & ~x71 & ~x86 & ~x111 & ~x113 & ~x140 & ~x168 & ~x169 & ~x435 & ~x470 & ~x489 & ~x710 & ~x783;
assign c0263 =  x211 & ~x26 & ~x407 & ~x684 & ~x745 & ~x763;
assign c0265 = ~x6 & ~x18 & ~x36 & ~x91 & ~x381 & ~x407 & ~x409 & ~x460 & ~x487 & ~x571 & ~x573 & ~x598 & ~x626 & ~x655 & ~x683 & ~x711 & ~x713 & ~x715;
assign c0267 = ~x325 & ~x380 & ~x403 & ~x459 & ~x517;
assign c0269 = ~x0 & ~x68 & ~x112 & ~x113 & ~x252 & ~x275 & ~x388 & ~x389 & ~x417 & ~x487 & ~x624 & ~x734 & ~x753;
assign c0271 =  x480 & ~x0 & ~x5 & ~x21 & ~x24 & ~x26 & ~x31 & ~x32 & ~x35 & ~x51 & ~x56 & ~x80 & ~x83 & ~x90 & ~x107 & ~x115 & ~x137 & ~x139 & ~x142 & ~x167 & ~x172 & ~x196 & ~x197 & ~x227 & ~x281 & ~x283 & ~x337 & ~x392 & ~x676 & ~x777 & ~x783;
assign c0273 =  x270 &  x313 &  x340 & ~x55 & ~x59 & ~x82 & ~x83 & ~x140 & ~x141 & ~x308;
assign c0275 =  x426 &  x480 & ~x21 & ~x108 & ~x114 & ~x135 & ~x193 & ~x281 & ~x282 & ~x484 & ~x670 & ~x783;
assign c0277 = ~x348 & ~x403 & ~x433 & ~x458 & ~x490 & ~x515 & ~x542 & ~x568 & ~x651 & ~x705 & ~x734 & ~x760;
assign c0279 = ~x48 & ~x56 & ~x65 & ~x93 & ~x109 & ~x111 & ~x148 & ~x202 & ~x224 & ~x227 & ~x229 & ~x252 & ~x254 & ~x255 & ~x257 & ~x283 & ~x284 & ~x706 & ~x778;
assign c0281 =  x182 & ~x322 & ~x377 & ~x591;
assign c0283 =  x241 &  x242 &  x269 & ~x23 & ~x24 & ~x336 & ~x364 & ~x391 & ~x392 & ~x419 & ~x700 & ~x767;
assign c0285 = ~x53 & ~x54 & ~x111 & ~x344 & ~x372 & ~x373 & ~x400 & ~x454 & ~x588 & ~x589 & ~x617 & ~x644 & ~x699 & ~x772;
assign c0287 =  x719 &  x749;
assign c0289 =  x379 &  x656 &  x657 & ~x1 & ~x222 & ~x756 & ~x780;
assign c0291 =  x400 &  x510 & ~x10 & ~x19 & ~x28 & ~x56 & ~x111 & ~x489 & ~x545 & ~x573 & ~x603 & ~x775;
assign c0293 =  x255 &  x310 &  x366 & ~x57 & ~x779;
assign c0295 =  x397 &  x425 & ~x0 & ~x1 & ~x17 & ~x30 & ~x48 & ~x61 & ~x62 & ~x85 & ~x90 & ~x191 & ~x228 & ~x252 & ~x254 & ~x282 & ~x758 & ~x778;
assign c0297 =  x482 & ~x145 & ~x436 & ~x463 & ~x544 & ~x597 & ~x707;
assign c0299 =  x717 & ~x555;
assign c0301 =  x246 & ~x1 & ~x7 & ~x21 & ~x25 & ~x33 & ~x51 & ~x84 & ~x111 & ~x232 & ~x596 & ~x699 & ~x755;
assign c0303 =  x667 & ~x528 & ~x557;
assign c0305 = ~x0 & ~x17 & ~x71 & ~x73 & ~x132 & ~x167 & ~x194 & ~x251 & ~x273 & ~x281 & ~x284 & ~x302 & ~x304 & ~x329 & ~x330 & ~x331 & ~x332 & ~x333 & ~x359 & ~x360 & ~x363 & ~x388 & ~x391 & ~x638 & ~x724 & ~x783;
assign c0307 = ~x2 & ~x53 & ~x179 & ~x221 & ~x316 & ~x361 & ~x363 & ~x389 & ~x417 & ~x531 & ~x783;
assign c0309 =  x151 & ~x540 & ~x649 & ~x705;
assign c0311 = ~x20 & ~x104 & ~x311 & ~x423 & ~x498 & ~x499 & ~x525 & ~x528 & ~x552 & ~x554 & ~x641 & ~x643 & ~x645 & ~x696 & ~x763;
assign c0313 = ~x21 & ~x109 & ~x112 & ~x336 & ~x377 & ~x404 & ~x433 & ~x488 & ~x490 & ~x515 & ~x576 & ~x601 & ~x603 & ~x629 & ~x678 & ~x679 & ~x707 & ~x733;
assign c0315 =  x237 &  x238 &  x296 & ~x55;
assign c0317 =  x296 & ~x98 & ~x316 & ~x777;
assign c0319 =  x256 &  x283 &  x338 &  x366 & ~x30 & ~x763;
assign c0321 = ~x126 & ~x160 & ~x241 & ~x265 & ~x367 & ~x396 & ~x452 & ~x562 & ~x587 & ~x613 & ~x619 & ~x672 & ~x673 & ~x731;
assign c0323 =  x426 & ~x8 & ~x21 & ~x23 & ~x24 & ~x25 & ~x26 & ~x51 & ~x61 & ~x77 & ~x140 & ~x144 & ~x169 & ~x172 & ~x196 & ~x197 & ~x199 & ~x223 & ~x231 & ~x251 & ~x282 & ~x643 & ~x670 & ~x729;
assign c0325 = ~x5 & ~x31 & ~x60 & ~x115 & ~x224 & ~x503 & ~x652;
assign c0327 =  x343 &  x344 &  x370 &  x371 & ~x84 & ~x433 & ~x575 & ~x608 & ~x632 & ~x691 & ~x736 & ~x763 & ~x766;
assign c0329 =  x163 & ~x506 & ~x534 & ~x543;
assign c0331 =  x240 &  x266 &  x267 &  x293 & ~x63 & ~x750 & ~x772;
assign c0333 =  x660 &  x661 & ~x528 & ~x652;
assign c0335 =  x266 &  x565 & ~x221 & ~x226 & ~x282 & ~x390 & ~x391 & ~x473 & ~x502;
assign c0337 = ~x0 & ~x3 & ~x29 & ~x43 & ~x83 & ~x235 & ~x236 & ~x395 & ~x397 & ~x420 & ~x423 & ~x424 & ~x452 & ~x476 & ~x525 & ~x526 & ~x531 & ~x645 & ~x673 & ~x728 & ~x750 & ~x763;
assign c0339 =  x328 &  x356 & ~x51 & ~x55 & ~x475 & ~x501 & ~x503 & ~x558 & ~x764;
assign c0341 =  x404 & ~x19 & ~x111 & ~x236 & ~x426 & ~x452 & ~x472 & ~x500;
assign c0343 = ~x15 & ~x83 & ~x238 & ~x239 & ~x250 & ~x396 & ~x422 & ~x451 & ~x497 & ~x500 & ~x501 & ~x524 & ~x526 & ~x527 & ~x529 & ~x557 & ~x580 & ~x582 & ~x672 & ~x761 & ~x782;
assign c0345 = ~x168 & ~x219 & ~x247 & ~x248 & ~x251 & ~x274 & ~x331 & ~x364 & ~x389 & ~x441 & ~x442 & ~x445 & ~x471 & ~x620;
assign c0347 = ~x297 & ~x374 & ~x401 & ~x429 & ~x458 & ~x484 & ~x512 & ~x540 & ~x567 & ~x593 & ~x594 & ~x621;
assign c0349 =  x481 &  x537 &  x564 & ~x29 & ~x406 & ~x515 & ~x517 & ~x571 & ~x572 & ~x599 & ~x706 & ~x736 & ~x739;
assign c0351 = ~x2 & ~x86 & ~x135 & ~x190 & ~x191 & ~x219 & ~x253 & ~x280 & ~x309 & ~x335 & ~x387 & ~x418 & ~x419 & ~x471 & ~x601 & ~x661 & ~x719;
assign c0353 = ~x15 & ~x265 & ~x397 & ~x454 & ~x480 & ~x537 & ~x590 & ~x614 & ~x699 & ~x761;
assign c0355 = ~x18 & ~x40 & ~x421 & ~x422 & ~x425 & ~x525 & ~x526 & ~x534 & ~x564 & ~x620 & ~x730;
assign c0357 = ~x18 & ~x29 & ~x44 & ~x45 & ~x74 & ~x75 & ~x83 & ~x103 & ~x218 & ~x219 & ~x250 & ~x277 & ~x305 & ~x331 & ~x333 & ~x335 & ~x360 & ~x361 & ~x388 & ~x389 & ~x420 & ~x444 & ~x445 & ~x446 & ~x447 & ~x527 & ~x529 & ~x530 & ~x747;
assign c0359 =  x416 &  x417 & ~x91 & ~x141 & ~x511 & ~x538 & ~x565 & ~x566 & ~x781;
assign c0361 = ~x7 & ~x8 & ~x18 & ~x25 & ~x29 & ~x32 & ~x33 & ~x42 & ~x58 & ~x59 & ~x60 & ~x71 & ~x83 & ~x85 & ~x86 & ~x87 & ~x96 & ~x114 & ~x115 & ~x141 & ~x142 & ~x143 & ~x144 & ~x169 & ~x170 & ~x196 & ~x392 & ~x460 & ~x487 & ~x515 & ~x516 & ~x544 & ~x545 & ~x571 & ~x573 & ~x601 & ~x603 & ~x627 & ~x629 & ~x630 & ~x643 & ~x656 & ~x683 & ~x710 & ~x711 & ~x714 & ~x764 & ~x767;
assign c0363 =  x742 & ~x331 & ~x637 & ~x645;
assign c0365 = ~x127 & ~x131 & ~x132 & ~x397 & ~x422 & ~x425 & ~x454 & ~x478 & ~x563 & ~x620 & ~x646 & ~x674 & ~x702 & ~x703 & ~x783;
assign c0367 = ~x27 & ~x54 & ~x82 & ~x373 & ~x401 & ~x427 & ~x533 & ~x560 & ~x562 & ~x588 & ~x589 & ~x616 & ~x645 & ~x672 & ~x729 & ~x745 & ~x746 & ~x773 & ~x782;
assign c0369 = ~x3 & ~x12 & ~x49 & ~x61 & ~x107 & ~x110 & ~x117 & ~x199 & ~x224 & ~x226 & ~x254 & ~x568 & ~x570 & ~x626 & ~x710 & ~x739 & ~x742 & ~x749 & ~x765 & ~x776;
assign c0371 = ~x28 & ~x84 & ~x347 & ~x374 & ~x375 & ~x402 & ~x431 & ~x432 & ~x441 & ~x448 & ~x485 & ~x512 & ~x623 & ~x650 & ~x678 & ~x729 & ~x760 & ~x762;
assign c0373 = ~x26 & ~x54 & ~x55 & ~x179 & ~x197 & ~x199 & ~x206 & ~x234 & ~x282 & ~x338 & ~x367 & ~x571 & ~x683;
assign c0375 =  x409 & ~x43 & ~x138 & ~x273 & ~x429;
assign c0377 =  x550 & ~x194 & ~x331 & ~x459 & ~x611 & ~x670;
assign c0379 = ~x57 & ~x150 & ~x177 & ~x205 & ~x223 & ~x286 & ~x313 & ~x763 & ~x771;
assign c0381 = ~x1 & ~x54 & ~x78 & ~x79 & ~x83 & ~x108 & ~x136 & ~x138 & ~x151 & ~x366 & ~x379 & ~x464 & ~x489 & ~x519 & ~x546 & ~x547 & ~x548 & ~x574 & ~x656 & ~x683 & ~x684 & ~x755 & ~x762 & ~x764 & ~x769 & ~x780;
assign c0383 =  x129 &  x156 & ~x15 & ~x67 & ~x603;
assign c0385 = ~x48 & ~x67 & ~x82 & ~x111 & ~x136 & ~x142 & ~x146 & ~x195 & ~x200 & ~x201 & ~x282 & ~x336 & ~x647 & ~x653 & ~x684 & ~x698 & ~x710 & ~x738 & ~x740 & ~x746 & ~x772 & ~x779;
assign c0387 =  x374 & ~x1 & ~x19 & ~x28 & ~x65 & ~x93 & ~x145 & ~x147 & ~x175 & ~x201 & ~x202 & ~x717 & ~x767;
assign c0389 =  x398 & ~x0 & ~x1 & ~x4 & ~x20 & ~x22 & ~x24 & ~x25 & ~x26 & ~x27 & ~x28 & ~x29 & ~x30 & ~x31 & ~x32 & ~x41 & ~x43 & ~x51 & ~x52 & ~x55 & ~x56 & ~x57 & ~x58 & ~x60 & ~x81 & ~x83 & ~x84 & ~x85 & ~x86 & ~x88 & ~x89 & ~x108 & ~x109 & ~x111 & ~x112 & ~x113 & ~x114 & ~x115 & ~x136 & ~x137 & ~x140 & ~x142 & ~x143 & ~x144 & ~x165 & ~x166 & ~x167 & ~x168 & ~x169 & ~x170 & ~x171 & ~x194 & ~x195 & ~x196 & ~x197 & ~x198 & ~x199 & ~x224 & ~x225 & ~x226 & ~x227 & ~x252 & ~x253 & ~x280 & ~x281 & ~x282 & ~x308 & ~x309 & ~x310 & ~x336 & ~x337 & ~x364 & ~x615 & ~x644 & ~x669 & ~x697 & ~x699 & ~x725 & ~x726 & ~x727 & ~x729 & ~x749 & ~x757 & ~x758 & ~x764 & ~x765 & ~x767 & ~x776 & ~x781 & ~x782 & ~x783;
assign c0391 =  x435 & ~x53 & ~x107 & ~x131 & ~x184 & ~x185 & ~x191 & ~x221 & ~x276 & ~x392 & ~x447;
assign c0393 =  x183 &  x210 & ~x463 & ~x782;
assign c0395 =  x641 & ~x170 & ~x225;
assign c0397 = ~x26 & ~x111 & ~x180 & ~x342 & ~x343 & ~x369 & ~x370 & ~x398 & ~x453 & ~x480 & ~x779;
assign c0399 = ~x20 & ~x44 & ~x68 & ~x72 & ~x75 & ~x481 & ~x508 & ~x509 & ~x533 & ~x535 & ~x537 & ~x560 & ~x561 & ~x563 & ~x590 & ~x616 & ~x617 & ~x619 & ~x620 & ~x674 & ~x727 & ~x753 & ~x756 & ~x763 & ~x764 & ~x768 & ~x769 & ~x778 & ~x779;
assign c0401 =  x269 & ~x86 & ~x113 & ~x115 & ~x625 & ~x682;
assign c0403 = ~x352 & ~x433 & ~x434 & ~x460 & ~x518 & ~x546 & ~x597 & ~x652 & ~x687 & ~x688 & ~x736 & ~x744 & ~x762;
assign c0405 =  x277 & ~x120 & ~x377 & ~x378 & ~x513 & ~x542 & ~x569 & ~x600;
assign c0407 =  x215 & ~x417 & ~x443 & ~x444 & ~x616;
assign c0409 =  x378 &  x653 &  x682 & ~x26 & ~x112 & ~x280;
assign c0411 = ~x0 & ~x24 & ~x43 & ~x71 & ~x291 & ~x395 & ~x424 & ~x449 & ~x452 & ~x479 & ~x480 & ~x508 & ~x564 & ~x614 & ~x699 & ~x764 & ~x766;
assign c0413 =  x382 & ~x83 & ~x470 & ~x528 & ~x529 & ~x530;
assign c0415 = ~x82 & ~x108 & ~x164 & ~x167 & ~x176 & ~x202 & ~x203 & ~x231 & ~x285 & ~x287;
assign c0417 = ~x25 & ~x374 & ~x402 & ~x430 & ~x431 & ~x432 & ~x460 & ~x486 & ~x488 & ~x621 & ~x648 & ~x650 & ~x651 & ~x678 & ~x707 & ~x732 & ~x734 & ~x761 & ~x762;
assign c0419 = ~x1 & ~x14 & ~x30 & ~x54 & ~x57 & ~x84 & ~x112 & ~x293 & ~x401 & ~x402 & ~x429 & ~x457 & ~x511 & ~x539 & ~x566 & ~x593 & ~x642 & ~x643 & ~x775;
assign c0421 =  x629 & ~x32 & ~x59 & ~x195 & ~x536 & ~x559 & ~x564 & ~x619 & ~x648 & ~x677 & ~x722 & ~x723 & ~x750 & ~x782;
assign c0423 = ~x17 & ~x23 & ~x25 & ~x30 & ~x31 & ~x44 & ~x51 & ~x60 & ~x79 & ~x115 & ~x117 & ~x144 & ~x168 & ~x169 & ~x172 & ~x173 & ~x180 & ~x197 & ~x201 & ~x207 & ~x228 & ~x282 & ~x283 & ~x338 & ~x339 & ~x643 & ~x729 & ~x783;
assign c0425 =  x179 &  x314 & ~x63 & ~x679;
assign c0427 =  x610 & ~x400 & ~x447 & ~x557 & ~x585;
assign c0429 = ~x2 & ~x9 & ~x18 & ~x19 & ~x23 & ~x24 & ~x30 & ~x31 & ~x32 & ~x33 & ~x51 & ~x56 & ~x61 & ~x82 & ~x84 & ~x87 & ~x108 & ~x109 & ~x113 & ~x114 & ~x137 & ~x138 & ~x139 & ~x141 & ~x142 & ~x165 & ~x169 & ~x172 & ~x193 & ~x196 & ~x198 & ~x221 & ~x224 & ~x227 & ~x228 & ~x253 & ~x255 & ~x280 & ~x281 & ~x307 & ~x309 & ~x310 & ~x336 & ~x337 & ~x363 & ~x365 & ~x391 & ~x448 & ~x577 & ~x726 & ~x728 & ~x730 & ~x781 & ~x782;
assign c0431 =  x183 &  x209 & ~x196 & ~x434 & ~x783;
assign c0433 = ~x54 & ~x261 & ~x313 & ~x314 & ~x340 & ~x341 & ~x368 & ~x396 & ~x420 & ~x587;
assign c0435 =  x158 & ~x83 & ~x140 & ~x231;
assign c0437 =  x13;
assign c0439 =  x426 & ~x31 & ~x41 & ~x50 & ~x80 & ~x108 & ~x137 & ~x379 & ~x433 & ~x570 & ~x599 & ~x629 & ~x630 & ~x762;
assign c0441 = ~x79 & ~x132 & ~x139 & ~x159 & ~x184 & ~x275 & ~x305 & ~x448 & ~x478 & ~x527 & ~x530 & ~x555 & ~x556 & ~x558 & ~x559 & ~x747 & ~x778;
assign c0443 = ~x23 & ~x56 & ~x78 & ~x348 & ~x507 & ~x510 & ~x702 & ~x769 & ~x781;
assign c0445 = ~x91 & ~x147 & ~x282 & ~x382 & ~x383 & ~x438 & ~x462 & ~x595 & ~x621 & ~x677 & ~x703;
assign c0447 =  x126 &  x153 &  x180 & ~x27 & ~x56 & ~x140 & ~x503 & ~x747 & ~x749 & ~x763;
assign c0449 =  x462 & ~x103 & ~x106 & ~x130 & ~x131 & ~x238 & ~x267 & ~x482 & ~x503 & ~x510;
assign c0451 =  x394 & ~x3 & ~x31 & ~x57 & ~x83 & ~x85 & ~x86 & ~x87 & ~x111 & ~x113 & ~x140 & ~x142 & ~x754 & ~x762 & ~x765 & ~x774;
assign c0453 =  x292 & ~x37 & ~x653;
assign c0455 = ~x50 & ~x51 & ~x136 & ~x379 & ~x460 & ~x462 & ~x518 & ~x570 & ~x573 & ~x598 & ~x629 & ~x631 & ~x632 & ~x660 & ~x661 & ~x707;
assign c0457 =  x674 & ~x56 & ~x281 & ~x308 & ~x736;
assign c0459 = ~x1 & ~x8 & ~x9 & ~x21 & ~x26 & ~x28 & ~x35 & ~x54 & ~x56 & ~x57 & ~x63 & ~x84 & ~x85 & ~x110 & ~x111 & ~x112 & ~x140 & ~x143 & ~x144 & ~x168 & ~x169 & ~x170 & ~x171 & ~x280 & ~x518 & ~x520 & ~x546 & ~x547 & ~x549 & ~x576 & ~x577 & ~x605 & ~x606 & ~x634 & ~x636 & ~x664 & ~x692 & ~x718 & ~x743 & ~x744 & ~x747 & ~x757 & ~x761 & ~x763 & ~x764 & ~x768 & ~x771;
assign c0461 = ~x10 & ~x25 & ~x45 & ~x147 & ~x181 & ~x255 & ~x393 & ~x408 & ~x550 & ~x719;
assign c0463 = ~x1 & ~x2 & ~x6 & ~x7 & ~x19 & ~x27 & ~x28 & ~x29 & ~x38 & ~x53 & ~x82 & ~x88 & ~x92 & ~x109 & ~x111 & ~x112 & ~x113 & ~x120 & ~x139 & ~x174 & ~x175 & ~x200 & ~x202 & ~x227 & ~x229 & ~x230 & ~x255 & ~x257 & ~x283 & ~x284 & ~x729 & ~x746 & ~x747 & ~x755 & ~x756 & ~x762 & ~x775;
assign c0465 =  x683 & ~x274 & ~x276 & ~x306 & ~x620;
assign c0467 = ~x113 & ~x265 & ~x319 & ~x399 & ~x426 & ~x503 & ~x532 & ~x589;
assign c0469 = ~x15 & ~x28 & ~x44 & ~x47 & ~x71 & ~x99 & ~x139 & ~x348 & ~x448 & ~x449 & ~x450 & ~x451 & ~x478 & ~x479 & ~x480 & ~x557 & ~x562 & ~x588 & ~x612 & ~x615 & ~x619 & ~x640 & ~x641 & ~x643 & ~x667 & ~x695 & ~x703 & ~x722 & ~x727 & ~x732 & ~x751 & ~x752 & ~x758 & ~x759 & ~x761 & ~x776;
assign c0471 = ~x29 & ~x32 & ~x195 & ~x197 & ~x247 & ~x274 & ~x275 & ~x302 & ~x304 & ~x331 & ~x391 & ~x418 & ~x445 & ~x446 & ~x497 & ~x558 & ~x584 & ~x611 & ~x642;
assign c0473 =  x327 & ~x25 & ~x389 & ~x390 & ~x443 & ~x471 & ~x764;
assign c0475 =  x648 & ~x335 & ~x543 & ~x627 & ~x658 & ~x682;
assign c0477 = ~x7 & ~x68 & ~x89 & ~x95 & ~x201 & ~x228 & ~x256 & ~x283 & ~x284 & ~x543 & ~x746;
assign c0479 =  x240 &  x515 & ~x567 & ~x650;
assign c0481 =  x416 & ~x5 & ~x62 & ~x353 & ~x405 & ~x406 & ~x623 & ~x652 & ~x677 & ~x678 & ~x761;
assign c0483 =  x239 & ~x1 & ~x23 & ~x53 & ~x81 & ~x84 & ~x139 & ~x142 & ~x196 & ~x199 & ~x224 & ~x225 & ~x227 & ~x253 & ~x475 & ~x503 & ~x753 & ~x754 & ~x755 & ~x759 & ~x770;
assign c0485 =  x398 & ~x54 & ~x107 & ~x151 & ~x296 & ~x352 & ~x486 & ~x624 & ~x683 & ~x722;
assign c0487 =  x718 & ~x277 & ~x308 & ~x553 & ~x582 & ~x671;
assign c0489 =  x228 & ~x441 & ~x473 & ~x474 & ~x479 & ~x498 & ~x501 & ~x588;
assign c0491 =  x90 & ~x304 & ~x305 & ~x362 & ~x391 & ~x445 & ~x446 & ~x447 & ~x474 & ~x503 & ~x561 & ~x616;
assign c0493 = ~x37 & ~x92 & ~x94 & ~x380 & ~x407 & ~x542 & ~x569 & ~x570 & ~x597 & ~x599 & ~x629 & ~x656 & ~x657 & ~x683 & ~x684 & ~x705;
assign c0495 =  x572 & ~x43 & ~x346 & ~x347 & ~x564 & ~x592 & ~x704 & ~x757;
assign c0497 =  x710 &  x712 & ~x475 & ~x562 & ~x589 & ~x590 & ~x617 & ~x619 & ~x670 & ~x753;
assign c0499 = ~x84 & ~x362 & ~x413 & ~x440 & ~x475 & ~x495 & ~x496;
assign c10 = ~x154 & ~x324 & ~x680;
assign c14 =  x231 &  x401 & ~x419 & ~x481 & ~x656;
assign c16 = ~x1 & ~x4 & ~x16 & ~x21 & ~x22 & ~x23 & ~x24 & ~x27 & ~x29 & ~x30 & ~x53 & ~x56 & ~x60 & ~x79 & ~x81 & ~x86 & ~x88 & ~x107 & ~x108 & ~x109 & ~x110 & ~x112 & ~x140 & ~x143 & ~x144 & ~x164 & ~x165 & ~x166 & ~x167 & ~x168 & ~x193 & ~x194 & ~x195 & ~x196 & ~x199 & ~x221 & ~x223 & ~x224 & ~x225 & ~x251 & ~x278 & ~x280 & ~x281 & ~x283 & ~x304 & ~x306 & ~x307 & ~x309 & ~x333 & ~x337 & ~x361 & ~x362 & ~x367 & ~x390 & ~x391 & ~x392 & ~x394 & ~x395 & ~x396 & ~x418 & ~x420 & ~x421 & ~x423 & ~x424 & ~x448 & ~x450 & ~x451 & ~x452 & ~x453 & ~x459 & ~x460 & ~x474 & ~x475 & ~x476 & ~x477 & ~x479 & ~x480 & ~x481 & ~x503 & ~x505 & ~x507 & ~x508 & ~x531 & ~x532 & ~x533 & ~x534 & ~x559 & ~x560 & ~x561 & ~x562 & ~x586 & ~x588 & ~x589 & ~x590 & ~x600 & ~x601 & ~x616 & ~x617 & ~x629 & ~x630 & ~x631 & ~x644 & ~x645 & ~x669 & ~x672 & ~x724 & ~x726 & ~x752 & ~x755 & ~x756 & ~x757 & ~x780 & ~x781;
assign c18 =  x711 & ~x28 & ~x81 & ~x118 & ~x144 & ~x146 & ~x172 & ~x203 & ~x229 & ~x230 & ~x287 & ~x313 & ~x314 & ~x338 & ~x341 & ~x342 & ~x343 & ~x419 & ~x423 & ~x477 & ~x643 & ~x646 & ~x671 & ~x686 & ~x717 & ~x719 & ~x728 & ~x747 & ~x774;
assign c110 =  x351 &  x521 & ~x0 & ~x62 & ~x85 & ~x89 & ~x119 & ~x131 & ~x158 & ~x161 & ~x165 & ~x168 & ~x173 & ~x174 & ~x185 & ~x188 & ~x189 & ~x194 & ~x202 & ~x214 & ~x225 & ~x230 & ~x244 & ~x246 & ~x252 & ~x256 & ~x284 & ~x303 & ~x306 & ~x307 & ~x330 & ~x335 & ~x336 & ~x338 & ~x357 & ~x358 & ~x361 & ~x368 & ~x369 & ~x370 & ~x416 & ~x423 & ~x425 & ~x445 & ~x470 & ~x472 & ~x473 & ~x475 & ~x483 & ~x527 & ~x533 & ~x557 & ~x558 & ~x618 & ~x620 & ~x639 & ~x666 & ~x671 & ~x676 & ~x677 & ~x697 & ~x705 & ~x721 & ~x724 & ~x736 & ~x759;
assign c112 =  x704 & ~x424 & ~x446 & ~x475 & ~x544 & ~x561 & ~x563 & ~x600 & ~x617 & ~x618 & ~x628 & ~x645 & ~x709 & ~x735 & ~x737;
assign c114 =  x326 &  x552 & ~x1 & ~x58 & ~x82 & ~x86 & ~x134 & ~x165 & ~x221 & ~x249 & ~x250 & ~x252 & ~x283 & ~x311 & ~x312 & ~x313 & ~x342 & ~x361 & ~x369 & ~x393 & ~x418 & ~x422 & ~x450 & ~x477 & ~x478 & ~x502 & ~x530 & ~x533 & ~x560 & ~x587 & ~x615 & ~x641 & ~x644 & ~x669 & ~x671 & ~x700 & ~x725 & ~x728 & ~x730 & ~x752 & ~x754 & ~x782;
assign c116 = ~x43 & ~x194 & ~x416 & ~x442 & ~x467 & ~x500 & ~x503 & ~x598 & ~x630 & ~x686 & ~x749;
assign c118 = ~x3 & ~x5 & ~x22 & ~x45 & ~x57 & ~x74 & ~x87 & ~x98 & ~x100 & ~x135 & ~x143 & ~x194 & ~x199 & ~x240 & ~x257 & ~x286 & ~x287 & ~x309 & ~x326 & ~x366 & ~x445 & ~x447 & ~x451 & ~x452 & ~x453 & ~x482 & ~x498 & ~x500 & ~x502 & ~x503 & ~x527 & ~x528 & ~x529 & ~x530 & ~x555 & ~x563 & ~x564 & ~x585 & ~x727 & ~x728 & ~x748 & ~x751 & ~x755;
assign c120 =  x678 & ~x0 & ~x24 & ~x26 & ~x54 & ~x100 & ~x111 & ~x223 & ~x251 & ~x254 & ~x280 & ~x307 & ~x390 & ~x391 & ~x392 & ~x393 & ~x475 & ~x506 & ~x517 & ~x545 & ~x563 & ~x572 & ~x656 & ~x729;
assign c122 =  x202 &  x428 & ~x180 & ~x627;
assign c124 =  x180 &  x322 &  x379 &  x407 & ~x42 & ~x276 & ~x442 & ~x609 & ~x722;
assign c126 =  x351 &  x379 & ~x21 & ~x107 & ~x133 & ~x138 & ~x145 & ~x146 & ~x185 & ~x211 & ~x212 & ~x222 & ~x241 & ~x280 & ~x299 & ~x304 & ~x327 & ~x357 & ~x368 & ~x482 & ~x483 & ~x510 & ~x528 & ~x555 & ~x583 & ~x614 & ~x619 & ~x621 & ~x647 & ~x701 & ~x727;
assign c128 = ~x0 & ~x5 & ~x32 & ~x46 & ~x83 & ~x87 & ~x105 & ~x141 & ~x166 & ~x173 & ~x189 & ~x248 & ~x276 & ~x277 & ~x303 & ~x305 & ~x308 & ~x309 & ~x334 & ~x335 & ~x336 & ~x367 & ~x369 & ~x373 & ~x374 & ~x375 & ~x376 & ~x394 & ~x396 & ~x419 & ~x422 & ~x423 & ~x446 & ~x527 & ~x545 & ~x546 & ~x556 & ~x557 & ~x562 & ~x575 & ~x586 & ~x589 & ~x643 & ~x671 & ~x729 & ~x731 & ~x749;
assign c130 =  x485 & ~x152 & ~x417 & ~x488 & ~x563 & ~x598 & ~x654 & ~x708;
assign c132 = ~x1 & ~x3 & ~x4 & ~x20 & ~x23 & ~x30 & ~x45 & ~x46 & ~x50 & ~x53 & ~x56 & ~x57 & ~x58 & ~x59 & ~x71 & ~x72 & ~x74 & ~x76 & ~x81 & ~x82 & ~x86 & ~x98 & ~x102 & ~x103 & ~x104 & ~x105 & ~x108 & ~x110 & ~x112 & ~x128 & ~x129 & ~x137 & ~x138 & ~x143 & ~x156 & ~x166 & ~x167 & ~x183 & ~x221 & ~x223 & ~x224 & ~x249 & ~x277 & ~x298 & ~x307 & ~x333 & ~x336 & ~x337 & ~x353 & ~x363 & ~x391 & ~x418 & ~x419 & ~x421 & ~x444 & ~x445 & ~x449 & ~x479 & ~x499 & ~x524 & ~x525 & ~x526 & ~x529 & ~x533 & ~x534 & ~x552 & ~x555 & ~x559 & ~x588 & ~x756 & ~x782;
assign c134 = ~x0 & ~x1 & ~x2 & ~x6 & ~x7 & ~x18 & ~x20 & ~x22 & ~x23 & ~x25 & ~x27 & ~x28 & ~x29 & ~x30 & ~x32 & ~x33 & ~x35 & ~x49 & ~x50 & ~x53 & ~x54 & ~x55 & ~x56 & ~x57 & ~x59 & ~x60 & ~x61 & ~x63 & ~x73 & ~x76 & ~x78 & ~x79 & ~x80 & ~x83 & ~x84 & ~x86 & ~x87 & ~x89 & ~x90 & ~x103 & ~x108 & ~x109 & ~x110 & ~x112 & ~x113 & ~x114 & ~x115 & ~x118 & ~x120 & ~x131 & ~x132 & ~x133 & ~x134 & ~x135 & ~x136 & ~x138 & ~x139 & ~x142 & ~x143 & ~x146 & ~x166 & ~x167 & ~x170 & ~x171 & ~x172 & ~x175 & ~x177 & ~x188 & ~x190 & ~x191 & ~x192 & ~x196 & ~x198 & ~x199 & ~x201 & ~x203 & ~x205 & ~x215 & ~x216 & ~x218 & ~x224 & ~x225 & ~x226 & ~x227 & ~x229 & ~x230 & ~x232 & ~x233 & ~x244 & ~x245 & ~x246 & ~x249 & ~x250 & ~x252 & ~x259 & ~x260 & ~x273 & ~x275 & ~x276 & ~x280 & ~x282 & ~x287 & ~x301 & ~x303 & ~x304 & ~x305 & ~x306 & ~x308 & ~x309 & ~x310 & ~x311 & ~x313 & ~x314 & ~x315 & ~x316 & ~x327 & ~x328 & ~x330 & ~x332 & ~x334 & ~x335 & ~x337 & ~x339 & ~x340 & ~x343 & ~x344 & ~x357 & ~x362 & ~x364 & ~x365 & ~x366 & ~x367 & ~x369 & ~x370 & ~x371 & ~x387 & ~x391 & ~x393 & ~x394 & ~x396 & ~x399 & ~x400 & ~x415 & ~x416 & ~x417 & ~x419 & ~x421 & ~x423 & ~x424 & ~x425 & ~x426 & ~x442 & ~x443 & ~x445 & ~x449 & ~x450 & ~x471 & ~x473 & ~x474 & ~x475 & ~x478 & ~x479 & ~x480 & ~x481 & ~x500 & ~x501 & ~x502 & ~x503 & ~x504 & ~x505 & ~x506 & ~x507 & ~x508 & ~x528 & ~x529 & ~x532 & ~x533 & ~x534 & ~x535 & ~x536 & ~x540 & ~x555 & ~x557 & ~x558 & ~x559 & ~x560 & ~x561 & ~x563 & ~x564 & ~x565 & ~x581 & ~x584 & ~x587 & ~x588 & ~x590 & ~x591 & ~x608 & ~x612 & ~x614 & ~x616 & ~x617 & ~x618 & ~x619 & ~x620 & ~x636 & ~x637 & ~x642 & ~x643 & ~x645 & ~x647 & ~x663 & ~x664 & ~x665 & ~x667 & ~x668 & ~x669 & ~x670 & ~x671 & ~x672 & ~x674 & ~x675 & ~x676 & ~x691 & ~x693 & ~x694 & ~x696 & ~x698 & ~x700 & ~x701 & ~x704 & ~x705 & ~x720 & ~x721 & ~x724 & ~x725 & ~x726 & ~x730 & ~x732 & ~x733 & ~x747 & ~x750 & ~x751 & ~x752 & ~x754 & ~x756 & ~x759 & ~x774 & ~x776 & ~x778 & ~x780;
assign c136 =  x297 &  x524 & ~x0 & ~x24 & ~x26 & ~x54 & ~x58 & ~x86 & ~x87 & ~x107 & ~x135 & ~x136 & ~x139 & ~x165 & ~x168 & ~x193 & ~x194 & ~x197 & ~x224 & ~x249 & ~x250 & ~x251 & ~x275 & ~x278 & ~x303 & ~x309 & ~x333 & ~x342 & ~x362 & ~x368 & ~x369 & ~x391 & ~x394 & ~x395 & ~x418 & ~x450 & ~x477 & ~x504 & ~x532 & ~x585 & ~x613 & ~x641 & ~x644 & ~x672 & ~x673 & ~x698 & ~x732 & ~x752 & ~x754 & ~x755 & ~x757;
assign c138 =  x89 &  x593;
assign c140 =  x407 &  x464 &  x656 & ~x412 & ~x439 & ~x603 & ~x649;
assign c142 =  x494 & ~x109 & ~x115 & ~x146 & ~x247 & ~x256 & ~x283 & ~x313 & ~x335 & ~x342 & ~x397 & ~x398 & ~x399 & ~x428 & ~x457 & ~x459 & ~x609 & ~x733 & ~x747;
assign c144 =  x246 &  x646;
assign c146 =  x675 & ~x97 & ~x597;
assign c148 = ~x471 & ~x496 & ~x498 & ~x502 & ~x505 & ~x627 & ~x629 & ~x723 & ~x724;
assign c150 =  x326 &  x469 & ~x27 & ~x53 & ~x56 & ~x57 & ~x58 & ~x80 & ~x81 & ~x111 & ~x113 & ~x136 & ~x139 & ~x197 & ~x253 & ~x254 & ~x283 & ~x311 & ~x333 & ~x340 & ~x361 & ~x362 & ~x367 & ~x369 & ~x418 & ~x419 & ~x447 & ~x561 & ~x587 & ~x614 & ~x643 & ~x669 & ~x696 & ~x755 & ~x782;
assign c152 =  x147 &  x566 &  x703;
assign c154 = ~x17 & ~x139 & ~x224 & ~x253 & ~x336 & ~x446 & ~x490 & ~x506 & ~x508 & ~x517 & ~x533 & ~x535 & ~x536 & ~x544 & ~x545 & ~x563 & ~x599 & ~x600 & ~x617 & ~x618 & ~x642 & ~x645 & ~x708 & ~x736;
assign c156 =  x662 & ~x71 & ~x166 & ~x251 & ~x279 & ~x364 & ~x533 & ~x552 & ~x557 & ~x616 & ~x656 & ~x715;
assign c158 =  x352 &  x550 & ~x60 & ~x102 & ~x135 & ~x172 & ~x187 & ~x190 & ~x191 & ~x271 & ~x275 & ~x276 & ~x314 & ~x342 & ~x392 & ~x395 & ~x396 & ~x480 & ~x529 & ~x537 & ~x584 & ~x620 & ~x621 & ~x732 & ~x777;
assign c160 =  x354 &  x524 &  x743 & ~x81 & ~x249 & ~x423 & ~x668 & ~x724;
assign c162 =  x68 &  x323 &  x436 &  x493 & ~x4 & ~x115 & ~x258 & ~x314 & ~x419 & ~x426 & ~x444 & ~x471 & ~x555 & ~x619 & ~x643 & ~x672 & ~x674 & ~x676 & ~x752 & ~x760 & ~x780;
assign c164 =  x709 &  x739 & ~x142 & ~x369 & ~x686 & ~x688;
assign c166 =  x551 &  x555 & ~x415 & ~x632;
assign c168 =  x240 &  x267 & ~x192 & ~x394 & ~x422 & ~x450 & ~x500 & ~x575 & ~x576 & ~x589 & ~x605 & ~x638 & ~x749 & ~x780;
assign c170 =  x323 &  x437 &  x465 &  x494 & ~x107 & ~x116 & ~x117 & ~x193 & ~x223 & ~x229 & ~x230 & ~x254 & ~x257 & ~x277 & ~x304 & ~x308 & ~x309 & ~x330 & ~x367 & ~x370 & ~x389 & ~x396 & ~x397 & ~x426 & ~x427 & ~x474 & ~x560 & ~x669 & ~x670 & ~x674 & ~x675 & ~x693 & ~x695 & ~x703 & ~x705 & ~x721 & ~x733 & ~x749 & ~x759 & ~x761;
assign c172 =  x705 & ~x56 & ~x111 & ~x195 & ~x335 & ~x392 & ~x451 & ~x474 & ~x475 & ~x478 & ~x479 & ~x504 & ~x509 & ~x562 & ~x616;
assign c174 = ~x58 & ~x103 & ~x109 & ~x141 & ~x164 & ~x222 & ~x229 & ~x253 & ~x283 & ~x315 & ~x316 & ~x317 & ~x334 & ~x336 & ~x342 & ~x343 & ~x344 & ~x346 & ~x347 & ~x391 & ~x396 & ~x490 & ~x492 & ~x504 & ~x530 & ~x549 & ~x697 & ~x700 & ~x752 & ~x779;
assign c176 =  x326 &  x441 &  x744 & ~x108 & ~x135 & ~x192 & ~x221 & ~x283 & ~x561 & ~x669;
assign c178 =  x552 &  x553 & ~x53 & ~x360 & ~x389 & ~x449 & ~x639 & ~x641 & ~x665 & ~x669 & ~x724;
assign c180 =  x684 & ~x147 & ~x205 & ~x240 & ~x315 & ~x495 & ~x768;
assign c182 =  x352 & ~x24 & ~x27 & ~x29 & ~x51 & ~x79 & ~x136 & ~x195 & ~x276 & ~x280 & ~x306 & ~x309 & ~x332 & ~x333 & ~x334 & ~x337 & ~x389 & ~x418 & ~x449 & ~x460 & ~x461 & ~x462 & ~x476 & ~x505 & ~x588 & ~x604 & ~x608 & ~x643 & ~x669 & ~x722 & ~x723 & ~x752 & ~x753 & ~x781;
assign c184 = ~x23 & ~x29 & ~x55 & ~x57 & ~x107 & ~x109 & ~x114 & ~x117 & ~x144 & ~x166 & ~x195 & ~x197 & ~x223 & ~x230 & ~x255 & ~x256 & ~x277 & ~x281 & ~x287 & ~x313 & ~x334 & ~x366 & ~x397 & ~x406 & ~x422 & ~x428 & ~x429 & ~x431 & ~x432 & ~x433 & ~x435 & ~x449 & ~x473 & ~x479 & ~x504 & ~x507 & ~x529 & ~x530 & ~x587 & ~x588 & ~x589 & ~x614 & ~x644 & ~x667 & ~x673 & ~x674 & ~x694 & ~x697 & ~x698 & ~x700 & ~x728 & ~x756 & ~x757;
assign c186 =  x90 & ~x96 & ~x506;
assign c188 = ~x27 & ~x80 & ~x81 & ~x82 & ~x109 & ~x111 & ~x114 & ~x196 & ~x306 & ~x391 & ~x418 & ~x449 & ~x462 & ~x503 & ~x600 & ~x601 & ~x602 & ~x631 & ~x660 & ~x661 & ~x692 & ~x695 & ~x721 & ~x722 & ~x725 & ~x756 & ~x776 & ~x777 & ~x779 & ~x782;
assign c190 =  x379 &  x578 & ~x28 & ~x31 & ~x58 & ~x79 & ~x106 & ~x140 & ~x141 & ~x142 & ~x163 & ~x164 & ~x224 & ~x246 & ~x254 & ~x285 & ~x302 & ~x304 & ~x306 & ~x311 & ~x313 & ~x334 & ~x338 & ~x422 & ~x443 & ~x477 & ~x481 & ~x483 & ~x502 & ~x505 & ~x506 & ~x507 & ~x512 & ~x563 & ~x674 & ~x702;
assign c192 = ~x96 & ~x97 & ~x181 & ~x296 & ~x362 & ~x417 & ~x545 & ~x572 & ~x708;
assign c194 = ~x4 & ~x21 & ~x22 & ~x24 & ~x27 & ~x28 & ~x29 & ~x53 & ~x54 & ~x58 & ~x62 & ~x78 & ~x80 & ~x84 & ~x85 & ~x89 & ~x90 & ~x105 & ~x109 & ~x119 & ~x134 & ~x137 & ~x139 & ~x141 & ~x142 & ~x145 & ~x165 & ~x171 & ~x172 & ~x190 & ~x194 & ~x195 & ~x198 & ~x202 & ~x220 & ~x222 & ~x224 & ~x230 & ~x248 & ~x276 & ~x281 & ~x283 & ~x305 & ~x313 & ~x314 & ~x338 & ~x339 & ~x340 & ~x341 & ~x342 & ~x343 & ~x344 & ~x345 & ~x346 & ~x347 & ~x348 & ~x349 & ~x350 & ~x360 & ~x373 & ~x388 & ~x392 & ~x418 & ~x419 & ~x420 & ~x421 & ~x445 & ~x448 & ~x473 & ~x475 & ~x504 & ~x529 & ~x530 & ~x586 & ~x612 & ~x615 & ~x617 & ~x668 & ~x669 & ~x671 & ~x673 & ~x674 & ~x699 & ~x700 & ~x723 & ~x724 & ~x753;
assign c196 = ~x66 & ~x97 & ~x167 & ~x363 & ~x388 & ~x412 & ~x414 & ~x443 & ~x487 & ~x679 & ~x706 & ~x707 & ~x734;
assign c198 = ~x98 & ~x126 & ~x270 & ~x324 & ~x335 & ~x352 & ~x469 & ~x471 & ~x475 & ~x504 & ~x516 & ~x711 & ~x763 & ~x768;
assign c1100 =  x654 &  x741 & ~x271 & ~x331 & ~x340 & ~x471 & ~x515 & ~x759;
assign c1102 =  x330 & ~x525;
assign c1104 =  x620 & ~x24 & ~x152 & ~x234 & ~x441 & ~x598 & ~x679 & ~x733;
assign c1106 = ~x18 & ~x51 & ~x77 & ~x81 & ~x85 & ~x87 & ~x165 & ~x195 & ~x251 & ~x255 & ~x281 & ~x338 & ~x397 & ~x400 & ~x404 & ~x419 & ~x421 & ~x478 & ~x544 & ~x545 & ~x602 & ~x603 & ~x605 & ~x724 & ~x778;
assign c1108 =  x664 & ~x16 & ~x17 & ~x71 & ~x73 & ~x79 & ~x501 & ~x525 & ~x553 & ~x629 & ~x710;
assign c1110 =  x642;
assign c1112 =  x627 & ~x114 & ~x145 & ~x175 & ~x254 & ~x306 & ~x338 & ~x341 & ~x477 & ~x515 & ~x517 & ~x518 & ~x544 & ~x643 & ~x723 & ~x755 & ~x778;
assign c1114 =  x239 & ~x4 & ~x19 & ~x24 & ~x108 & ~x115 & ~x141 & ~x172 & ~x194 & ~x197 & ~x227 & ~x251 & ~x254 & ~x276 & ~x279 & ~x305 & ~x312 & ~x335 & ~x337 & ~x338 & ~x339 & ~x340 & ~x341 & ~x360 & ~x364 & ~x393 & ~x420 & ~x421 & ~x424 & ~x452 & ~x475 & ~x477 & ~x479 & ~x480 & ~x490 & ~x491 & ~x503 & ~x510 & ~x511 & ~x530 & ~x559 & ~x565 & ~x585 & ~x589 & ~x618 & ~x673 & ~x675 & ~x698 & ~x702 & ~x723 & ~x726 & ~x731 & ~x749 & ~x750 & ~x751 & ~x754 & ~x761 & ~x776;
assign c1116 = ~x185 & ~x240 & ~x241 & ~x287 & ~x298 & ~x353 & ~x369 & ~x383 & ~x438 & ~x596 & ~x706;
assign c1118 =  x1;
assign c1120 = ~x28 & ~x59 & ~x104 & ~x129 & ~x143 & ~x173 & ~x198 & ~x199 & ~x241 & ~x255 & ~x269 & ~x286 & ~x298 & ~x299 & ~x312 & ~x314 & ~x327 & ~x328 & ~x354 & ~x385 & ~x413 & ~x425 & ~x451 & ~x480 & ~x538 & ~x539 & ~x544 & ~x642 & ~x671 & ~x721 & ~x752 & ~x754;
assign c1122 =  x609;
assign c1124 =  x634 & ~x448 & ~x497 & ~x534 & ~x572 & ~x582 & ~x746 & ~x773;
assign c1126 = ~x4 & ~x17 & ~x20 & ~x23 & ~x24 & ~x27 & ~x29 & ~x30 & ~x32 & ~x44 & ~x52 & ~x53 & ~x54 & ~x58 & ~x81 & ~x84 & ~x85 & ~x107 & ~x110 & ~x111 & ~x113 & ~x114 & ~x115 & ~x137 & ~x143 & ~x144 & ~x164 & ~x168 & ~x169 & ~x171 & ~x200 & ~x220 & ~x221 & ~x222 & ~x225 & ~x227 & ~x249 & ~x251 & ~x275 & ~x278 & ~x281 & ~x283 & ~x308 & ~x312 & ~x313 & ~x335 & ~x336 & ~x337 & ~x361 & ~x362 & ~x365 & ~x392 & ~x417 & ~x419 & ~x420 & ~x421 & ~x423 & ~x424 & ~x447 & ~x448 & ~x449 & ~x454 & ~x472 & ~x474 & ~x481 & ~x505 & ~x506 & ~x508 & ~x509 & ~x516 & ~x534 & ~x537 & ~x544 & ~x545 & ~x546 & ~x558 & ~x559 & ~x563 & ~x564 & ~x575 & ~x590 & ~x613 & ~x616 & ~x642 & ~x643 & ~x644 & ~x646 & ~x670 & ~x672 & ~x674 & ~x697 & ~x698 & ~x699 & ~x725 & ~x726 & ~x727 & ~x728 & ~x729 & ~x752 & ~x754 & ~x755 & ~x757;
assign c1128 = ~x24 & ~x29 & ~x75 & ~x77 & ~x79 & ~x81 & ~x85 & ~x103 & ~x104 & ~x110 & ~x138 & ~x144 & ~x145 & ~x160 & ~x161 & ~x162 & ~x199 & ~x222 & ~x224 & ~x225 & ~x277 & ~x281 & ~x282 & ~x285 & ~x311 & ~x340 & ~x341 & ~x391 & ~x392 & ~x395 & ~x396 & ~x397 & ~x399 & ~x400 & ~x401 & ~x402 & ~x403 & ~x404 & ~x426 & ~x447 & ~x474 & ~x529 & ~x546 & ~x547 & ~x548 & ~x549 & ~x615 & ~x645 & ~x668 & ~x671 & ~x702;
assign c1130 =  x711 & ~x0 & ~x27 & ~x29 & ~x32 & ~x54 & ~x85 & ~x113 & ~x137 & ~x170 & ~x229 & ~x255 & ~x277 & ~x281 & ~x283 & ~x306 & ~x390 & ~x397 & ~x424 & ~x451 & ~x476 & ~x507 & ~x533 & ~x589 & ~x628 & ~x658 & ~x669 & ~x718 & ~x724 & ~x729 & ~x731 & ~x747 & ~x780;
assign c1132 =  x348 & ~x33 & ~x116 & ~x118 & ~x202 & ~x212 & ~x270 & ~x314 & ~x354 & ~x399 & ~x426 & ~x456 & ~x457 & ~x553 & ~x566 & ~x582 & ~x587;
assign c1134 =  x38 &  x322 &  x351 & ~x62 & ~x109 & ~x148 & ~x312 & ~x337 & ~x367 & ~x423 & ~x481 & ~x590 & ~x781;
assign c1136 = ~x17 & ~x26 & ~x28 & ~x32 & ~x86 & ~x142 & ~x169 & ~x195 & ~x196 & ~x250 & ~x306 & ~x311 & ~x363 & ~x367 & ~x389 & ~x393 & ~x394 & ~x418 & ~x419 & ~x422 & ~x433 & ~x447 & ~x450 & ~x452 & ~x476 & ~x520 & ~x584 & ~x589 & ~x633 & ~x634 & ~x638 & ~x639 & ~x644 & ~x662 & ~x666 & ~x667 & ~x668 & ~x669 & ~x671 & ~x721 & ~x750 & ~x752;
assign c1138 =  x684 & ~x62 & ~x90 & ~x101 & ~x147 & ~x241 & ~x269 & ~x283 & ~x326 & ~x424 & ~x426 & ~x438 & ~x447 & ~x505;
assign c1140 =  x153 &  x295 &  x324 & ~x14 & ~x117 & ~x364 & ~x547 & ~x548 & ~x591 & ~x749;
assign c1142 = ~x27 & ~x139 & ~x143 & ~x166 & ~x199 & ~x222 & ~x253 & ~x308 & ~x363 & ~x367 & ~x368 & ~x377 & ~x398 & ~x403 & ~x422 & ~x448 & ~x477 & ~x478 & ~x506 & ~x546 & ~x561 & ~x576 & ~x577 & ~x585 & ~x668 & ~x671 & ~x697 & ~x748 & ~x755 & ~x783;
assign c1144 =  x436 & ~x91 & ~x100 & ~x143 & ~x146 & ~x165 & ~x170 & ~x221 & ~x233 & ~x317 & ~x328 & ~x341 & ~x420 & ~x566 & ~x674 & ~x747;
assign c1146 =  x594 & ~x452 & ~x480 & ~x561 & ~x601 & ~x631;
assign c1148 =  x407 &  x548 &  x577 & ~x145 & ~x268 & ~x269;
assign c1150 =  x330 &  x356 & ~x16 & ~x445 & ~x446;
assign c1152 = ~x146 & ~x249 & ~x298 & ~x328 & ~x355 & ~x384 & ~x415 & ~x483 & ~x545 & ~x547 & ~x549 & ~x594 & ~x631;
assign c1154 =  x128 &  x217 & ~x249 & ~x304 & ~x305 & ~x390;
assign c1156 =  x97 &  x239 &  x267 &  x296 & ~x5 & ~x14 & ~x49 & ~x54 & ~x77 & ~x110 & ~x228 & ~x229 & ~x308 & ~x309 & ~x365 & ~x366 & ~x393 & ~x422 & ~x444 & ~x449 & ~x477 & ~x505 & ~x529 & ~x637 & ~x639 & ~x640 & ~x645 & ~x666 & ~x668 & ~x677 & ~x703 & ~x722 & ~x723 & ~x783;
assign c1158 =  x211 &  x296 & ~x15 & ~x58 & ~x109 & ~x113 & ~x164 & ~x166 & ~x168 & ~x192 & ~x221 & ~x251 & ~x277 & ~x310 & ~x337 & ~x361 & ~x396 & ~x481 & ~x504 & ~x507 & ~x511 & ~x520 & ~x538 & ~x751;
assign c1160 =  x634 &  x663 &  x666 & ~x657;
assign c1162 = ~x30 & ~x53 & ~x54 & ~x58 & ~x87 & ~x109 & ~x112 & ~x115 & ~x117 & ~x136 & ~x145 & ~x146 & ~x147 & ~x166 & ~x167 & ~x169 & ~x170 & ~x172 & ~x176 & ~x177 & ~x189 & ~x193 & ~x194 & ~x199 & ~x201 & ~x229 & ~x249 & ~x258 & ~x277 & ~x279 & ~x286 & ~x306 & ~x315 & ~x331 & ~x337 & ~x342 & ~x364 & ~x365 & ~x389 & ~x390 & ~x393 & ~x395 & ~x398 & ~x418 & ~x420 & ~x447 & ~x448 & ~x450 & ~x452 & ~x454 & ~x455 & ~x475 & ~x484 & ~x485 & ~x486 & ~x488 & ~x489 & ~x490 & ~x506 & ~x534 & ~x561 & ~x589 & ~x619 & ~x642 & ~x645 & ~x676 & ~x696 & ~x698 & ~x752 & ~x753 & ~x760 & ~x761;
assign c1164 =  x39 &  x96 &  x239 &  x267 &  x295 & ~x192 & ~x253 & ~x254 & ~x282 & ~x304 & ~x306 & ~x450 & ~x479 & ~x498 & ~x583 & ~x619 & ~x621 & ~x665 & ~x704 & ~x782;
assign c1166 =  x436 & ~x193 & ~x211 & ~x304 & ~x382 & ~x414 & ~x444 & ~x474 & ~x516 & ~x722;
assign c1168 =  x684 & ~x147 & ~x171 & ~x212 & ~x313 & ~x325 & ~x355 & ~x381 & ~x411 & ~x438 & ~x466 & ~x495 & ~x594 & ~x622 & ~x648 & ~x705;
assign c1170 =  x524 & ~x30 & ~x54 & ~x56 & ~x86 & ~x112 & ~x137 & ~x139 & ~x165 & ~x167 & ~x169 & ~x193 & ~x194 & ~x196 & ~x197 & ~x221 & ~x224 & ~x248 & ~x249 & ~x251 & ~x252 & ~x254 & ~x277 & ~x278 & ~x279 & ~x281 & ~x333 & ~x362 & ~x389 & ~x391 & ~x393 & ~x394 & ~x418 & ~x419 & ~x422 & ~x423 & ~x448 & ~x450 & ~x475 & ~x477 & ~x533 & ~x633 & ~x634 & ~x638 & ~x641 & ~x642 & ~x663 & ~x664 & ~x665 & ~x666 & ~x667 & ~x668 & ~x671 & ~x694 & ~x697 & ~x699 & ~x722 & ~x723 & ~x725 & ~x727 & ~x728 & ~x751 & ~x753 & ~x754 & ~x780 & ~x781;
assign c1172 =  x433 & ~x71 & ~x268 & ~x269 & ~x285 & ~x326 & ~x426 & ~x484 & ~x512 & ~x539 & ~x581 & ~x672 & ~x723 & ~x747;
assign c1174 =  x435 & ~x100 & ~x128 & ~x130 & ~x174 & ~x193 & ~x272 & ~x313 & ~x340 & ~x381 & ~x438 & ~x442 & ~x479 & ~x566 & ~x754 & ~x776;
assign c1176 =  x303 &  x579 & ~x470;
assign c1178 =  x407 &  x436 & ~x84 & ~x137 & ~x141 & ~x184 & ~x222 & ~x304 & ~x328 & ~x381 & ~x410 & ~x411 & ~x442 & ~x616 & ~x624 & ~x706 & ~x735;
assign c1180 = ~x50 & ~x52 & ~x55 & ~x56 & ~x58 & ~x79 & ~x80 & ~x85 & ~x112 & ~x114 & ~x115 & ~x136 & ~x167 & ~x168 & ~x169 & ~x195 & ~x196 & ~x221 & ~x223 & ~x226 & ~x252 & ~x279 & ~x282 & ~x306 & ~x309 & ~x310 & ~x311 & ~x312 & ~x333 & ~x338 & ~x342 & ~x361 & ~x364 & ~x365 & ~x391 & ~x396 & ~x397 & ~x418 & ~x419 & ~x420 & ~x422 & ~x427 & ~x429 & ~x431 & ~x432 & ~x433 & ~x435 & ~x436 & ~x449 & ~x450 & ~x452 & ~x475 & ~x476 & ~x478 & ~x504 & ~x505 & ~x586 & ~x587 & ~x588 & ~x614 & ~x670 & ~x725 & ~x728 & ~x753 & ~x759;
assign c1182 = ~x0 & ~x1 & ~x2 & ~x5 & ~x23 & ~x27 & ~x28 & ~x31 & ~x55 & ~x59 & ~x72 & ~x82 & ~x84 & ~x86 & ~x112 & ~x113 & ~x115 & ~x130 & ~x158 & ~x166 & ~x169 & ~x170 & ~x192 & ~x193 & ~x194 & ~x195 & ~x199 & ~x200 & ~x221 & ~x223 & ~x277 & ~x279 & ~x283 & ~x305 & ~x307 & ~x311 & ~x336 & ~x337 & ~x339 & ~x361 & ~x362 & ~x365 & ~x366 & ~x368 & ~x369 & ~x390 & ~x391 & ~x395 & ~x396 & ~x417 & ~x423 & ~x446 & ~x450 & ~x476 & ~x477 & ~x481 & ~x501 & ~x504 & ~x506 & ~x509 & ~x529 & ~x536 & ~x557 & ~x558 & ~x560 & ~x564 & ~x590 & ~x646 & ~x656 & ~x658 & ~x659 & ~x669 & ~x670 & ~x686 & ~x700 & ~x702 & ~x726 & ~x727 & ~x752 & ~x753 & ~x755 & ~x756 & ~x758 & ~x763;
assign c1184 =  x268 &  x411 & ~x105 & ~x194 & ~x197 & ~x229 & ~x248 & ~x282 & ~x283 & ~x312 & ~x340 & ~x397 & ~x399 & ~x533 & ~x585 & ~x641 & ~x672 & ~x675 & ~x698 & ~x783;
assign c1186 =  x174 & ~x44 & ~x406 & ~x654;
assign c1188 =  x730 & ~x562;
assign c1190 = ~x21 & ~x24 & ~x25 & ~x74 & ~x82 & ~x86 & ~x88 & ~x108 & ~x109 & ~x129 & ~x137 & ~x140 & ~x144 & ~x146 & ~x147 & ~x168 & ~x175 & ~x194 & ~x216 & ~x226 & ~x245 & ~x250 & ~x254 & ~x269 & ~x270 & ~x278 & ~x298 & ~x310 & ~x312 & ~x314 & ~x326 & ~x329 & ~x333 & ~x334 & ~x335 & ~x354 & ~x360 & ~x361 & ~x362 & ~x364 & ~x368 & ~x369 & ~x386 & ~x415 & ~x454 & ~x481 & ~x482 & ~x483 & ~x502 & ~x506 & ~x508 & ~x511 & ~x526 & ~x528 & ~x539 & ~x540 & ~x544 & ~x555 & ~x560 & ~x593 & ~x594 & ~x614 & ~x645 & ~x724 & ~x726 & ~x728 & ~x776 & ~x780;
assign c1192 =  x557;
assign c1194 =  x326 &  x497 & ~x283 & ~x368 & ~x369 & ~x395 & ~x398 & ~x476 & ~x641 & ~x668 & ~x725;
assign c1196 = ~x18 & ~x19 & ~x48 & ~x51 & ~x88 & ~x106 & ~x110 & ~x163 & ~x165 & ~x193 & ~x248 & ~x254 & ~x278 & ~x361 & ~x394 & ~x399 & ~x400 & ~x401 & ~x402 & ~x403 & ~x421 & ~x479 & ~x573 & ~x574 & ~x602 & ~x603 & ~x605 & ~x671 & ~x702 & ~x722 & ~x729 & ~x762;
assign c1198 =  x298 &  x440 & ~x56 & ~x84 & ~x113 & ~x198 & ~x251 & ~x254 & ~x283 & ~x305 & ~x334 & ~x340 & ~x341 & ~x361 & ~x368 & ~x369 & ~x370 & ~x391 & ~x392 & ~x396 & ~x423 & ~x449 & ~x450 & ~x475 & ~x478 & ~x532 & ~x561 & ~x562 & ~x586 & ~x617 & ~x643 & ~x645 & ~x670 & ~x725 & ~x726 & ~x755 & ~x782;
assign c1200 = ~x1 & ~x16 & ~x17 & ~x23 & ~x29 & ~x43 & ~x44 & ~x45 & ~x50 & ~x54 & ~x56 & ~x82 & ~x97 & ~x106 & ~x137 & ~x139 & ~x140 & ~x165 & ~x168 & ~x195 & ~x223 & ~x249 & ~x251 & ~x278 & ~x280 & ~x306 & ~x308 & ~x363 & ~x390 & ~x391 & ~x445 & ~x447 & ~x474 & ~x475 & ~x495 & ~x496 & ~x497 & ~x498 & ~x499 & ~x528 & ~x529 & ~x530 & ~x531 & ~x654 & ~x681 & ~x709 & ~x710 & ~x740 & ~x756;
assign c1202 = ~x5 & ~x24 & ~x25 & ~x28 & ~x29 & ~x30 & ~x58 & ~x60 & ~x76 & ~x78 & ~x79 & ~x82 & ~x84 & ~x86 & ~x91 & ~x107 & ~x108 & ~x114 & ~x115 & ~x117 & ~x135 & ~x138 & ~x143 & ~x165 & ~x199 & ~x222 & ~x226 & ~x227 & ~x254 & ~x255 & ~x256 & ~x279 & ~x312 & ~x313 & ~x337 & ~x338 & ~x344 & ~x346 & ~x347 & ~x348 & ~x366 & ~x368 & ~x373 & ~x391 & ~x397 & ~x422 & ~x424 & ~x451 & ~x517 & ~x532 & ~x546 & ~x558 & ~x613 & ~x616 & ~x617 & ~x698 & ~x754 & ~x755 & ~x757 & ~x763;
assign c1204 =  x124 & ~x43 & ~x174 & ~x215 & ~x279 & ~x340 & ~x383 & ~x394 & ~x482 & ~x530 & ~x723 & ~x730 & ~x744 & ~x749;
assign c1206 =  x70 & ~x5 & ~x36 & ~x54 & ~x59 & ~x74 & ~x77 & ~x81 & ~x82 & ~x85 & ~x102 & ~x111 & ~x112 & ~x132 & ~x133 & ~x139 & ~x140 & ~x141 & ~x142 & ~x143 & ~x146 & ~x162 & ~x164 & ~x171 & ~x172 & ~x173 & ~x192 & ~x197 & ~x198 & ~x201 & ~x224 & ~x225 & ~x228 & ~x231 & ~x244 & ~x245 & ~x248 & ~x250 & ~x255 & ~x258 & ~x277 & ~x279 & ~x312 & ~x313 & ~x336 & ~x338 & ~x341 & ~x342 & ~x366 & ~x370 & ~x371 & ~x392 & ~x396 & ~x400 & ~x401 & ~x421 & ~x423 & ~x429 & ~x431 & ~x443 & ~x444 & ~x448 & ~x454 & ~x472 & ~x477 & ~x479 & ~x500 & ~x504 & ~x507 & ~x530 & ~x533 & ~x534 & ~x535 & ~x559 & ~x586 & ~x591 & ~x608 & ~x610 & ~x614 & ~x615 & ~x616 & ~x644 & ~x663 & ~x668 & ~x669 & ~x671 & ~x672 & ~x673 & ~x692 & ~x693 & ~x696 & ~x703 & ~x721 & ~x722 & ~x727 & ~x728 & ~x749 & ~x755 & ~x756 & ~x777 & ~x783;
assign c1208 =  x301 & ~x0 & ~x15 & ~x16 & ~x23 & ~x45 & ~x47 & ~x49 & ~x305 & ~x332 & ~x360 & ~x391 & ~x417;
assign c1210 = ~x0 & ~x1 & ~x20 & ~x24 & ~x27 & ~x28 & ~x43 & ~x51 & ~x53 & ~x72 & ~x80 & ~x81 & ~x82 & ~x84 & ~x109 & ~x110 & ~x112 & ~x139 & ~x165 & ~x167 & ~x168 & ~x169 & ~x170 & ~x192 & ~x193 & ~x195 & ~x249 & ~x250 & ~x251 & ~x278 & ~x279 & ~x305 & ~x306 & ~x361 & ~x363 & ~x390 & ~x393 & ~x418 & ~x420 & ~x444 & ~x446 & ~x447 & ~x473 & ~x476 & ~x498 & ~x499 & ~x500 & ~x505 & ~x523 & ~x528 & ~x529 & ~x532 & ~x533 & ~x534 & ~x560 & ~x686 & ~x715 & ~x743 & ~x772 & ~x773 & ~x774 & ~x776 & ~x778 & ~x781 & ~x782;
assign c1212 =  x127 &  x297 &  x354 &  x411 & ~x83 & ~x193 & ~x283 & ~x310 & ~x338 & ~x365 & ~x562 & ~x589 & ~x696;
assign c1214 = ~x508 & ~x509 & ~x563 & ~x575 & ~x636 & ~x768;
assign c1216 = ~x24 & ~x27 & ~x28 & ~x29 & ~x51 & ~x58 & ~x81 & ~x82 & ~x83 & ~x84 & ~x113 & ~x114 & ~x138 & ~x140 & ~x142 & ~x143 & ~x171 & ~x198 & ~x223 & ~x226 & ~x227 & ~x254 & ~x279 & ~x283 & ~x306 & ~x307 & ~x309 & ~x333 & ~x334 & ~x336 & ~x362 & ~x363 & ~x364 & ~x366 & ~x367 & ~x388 & ~x389 & ~x394 & ~x396 & ~x418 & ~x422 & ~x423 & ~x424 & ~x425 & ~x448 & ~x450 & ~x451 & ~x452 & ~x454 & ~x475 & ~x476 & ~x479 & ~x490 & ~x491 & ~x509 & ~x531 & ~x560 & ~x562 & ~x618 & ~x643 & ~x645 & ~x668 & ~x669 & ~x672 & ~x674 & ~x694 & ~x722 & ~x725 & ~x729 & ~x752 & ~x754 & ~x758;
assign c1218 = ~x0 & ~x1 & ~x4 & ~x5 & ~x22 & ~x23 & ~x25 & ~x26 & ~x27 & ~x28 & ~x29 & ~x31 & ~x32 & ~x50 & ~x52 & ~x53 & ~x54 & ~x55 & ~x56 & ~x57 & ~x58 & ~x79 & ~x80 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x86 & ~x91 & ~x103 & ~x107 & ~x108 & ~x109 & ~x110 & ~x111 & ~x112 & ~x113 & ~x115 & ~x136 & ~x137 & ~x140 & ~x141 & ~x142 & ~x143 & ~x164 & ~x165 & ~x166 & ~x167 & ~x168 & ~x169 & ~x170 & ~x191 & ~x193 & ~x194 & ~x195 & ~x196 & ~x197 & ~x200 & ~x219 & ~x221 & ~x222 & ~x223 & ~x224 & ~x225 & ~x246 & ~x249 & ~x251 & ~x276 & ~x277 & ~x278 & ~x279 & ~x280 & ~x281 & ~x282 & ~x283 & ~x302 & ~x304 & ~x305 & ~x307 & ~x308 & ~x309 & ~x311 & ~x331 & ~x333 & ~x335 & ~x336 & ~x337 & ~x339 & ~x342 & ~x343 & ~x360 & ~x361 & ~x362 & ~x363 & ~x364 & ~x365 & ~x366 & ~x367 & ~x368 & ~x373 & ~x387 & ~x388 & ~x389 & ~x390 & ~x391 & ~x392 & ~x393 & ~x394 & ~x403 & ~x416 & ~x417 & ~x418 & ~x419 & ~x420 & ~x421 & ~x422 & ~x423 & ~x424 & ~x428 & ~x445 & ~x446 & ~x447 & ~x448 & ~x449 & ~x450 & ~x451 & ~x471 & ~x472 & ~x474 & ~x475 & ~x476 & ~x477 & ~x478 & ~x479 & ~x500 & ~x502 & ~x504 & ~x505 & ~x506 & ~x529 & ~x532 & ~x533 & ~x534 & ~x556 & ~x557 & ~x559 & ~x560 & ~x561 & ~x563 & ~x583 & ~x585 & ~x587 & ~x588 & ~x589 & ~x590 & ~x608 & ~x609 & ~x611 & ~x614 & ~x615 & ~x616 & ~x619 & ~x632 & ~x633 & ~x634 & ~x635 & ~x636 & ~x637 & ~x638 & ~x639 & ~x640 & ~x641 & ~x642 & ~x643 & ~x644 & ~x661 & ~x662 & ~x663 & ~x664 & ~x665 & ~x666 & ~x667 & ~x668 & ~x669 & ~x670 & ~x671 & ~x690 & ~x691 & ~x692 & ~x693 & ~x694 & ~x695 & ~x696 & ~x697 & ~x698 & ~x699 & ~x700 & ~x701 & ~x718 & ~x720 & ~x721 & ~x722 & ~x723 & ~x724 & ~x725 & ~x726 & ~x727 & ~x728 & ~x729 & ~x731 & ~x748 & ~x749 & ~x751 & ~x752 & ~x754 & ~x755 & ~x756 & ~x757 & ~x758 & ~x761 & ~x762 & ~x763 & ~x776 & ~x777 & ~x778 & ~x779 & ~x780 & ~x781 & ~x782 & ~x783;
assign c1220 = ~x107 & ~x208 & ~x279 & ~x366 & ~x394 & ~x420 & ~x422 & ~x505 & ~x535 & ~x537 & ~x564 & ~x628 & ~x646 & ~x656 & ~x658 & ~x685 & ~x755;
assign c1222 =  x239 &  x352 &  x409 & ~x28 & ~x43 & ~x72 & ~x108 & ~x138 & ~x169 & ~x192 & ~x197 & ~x250 & ~x422 & ~x442 & ~x665 & ~x667;
assign c1224 =  x703 & ~x125 & ~x489 & ~x708;
assign c1226 =  x324 & ~x21 & ~x28 & ~x32 & ~x54 & ~x59 & ~x136 & ~x137 & ~x221 & ~x280 & ~x305 & ~x306 & ~x388 & ~x389 & ~x393 & ~x431 & ~x433 & ~x446 & ~x449 & ~x475 & ~x478 & ~x503 & ~x617 & ~x631 & ~x632 & ~x661 & ~x664 & ~x665 & ~x672 & ~x695 & ~x726 & ~x752 & ~x754;
assign c1228 = ~x20 & ~x26 & ~x32 & ~x53 & ~x108 & ~x136 & ~x140 & ~x160 & ~x165 & ~x250 & ~x276 & ~x341 & ~x393 & ~x396 & ~x399 & ~x401 & ~x402 & ~x405 & ~x449 & ~x455 & ~x477 & ~x530 & ~x546 & ~x547 & ~x557 & ~x559 & ~x576 & ~x577 & ~x585 & ~x668 & ~x674 & ~x696 & ~x728 & ~x759;
assign c1230 =  x713 &  x714 & ~x0 & ~x2 & ~x21 & ~x26 & ~x28 & ~x86 & ~x91 & ~x108 & ~x114 & ~x118 & ~x137 & ~x140 & ~x142 & ~x143 & ~x169 & ~x170 & ~x171 & ~x199 & ~x222 & ~x224 & ~x225 & ~x226 & ~x250 & ~x251 & ~x253 & ~x277 & ~x282 & ~x283 & ~x305 & ~x308 & ~x309 & ~x310 & ~x311 & ~x333 & ~x336 & ~x337 & ~x339 & ~x363 & ~x369 & ~x389 & ~x391 & ~x392 & ~x418 & ~x420 & ~x421 & ~x422 & ~x448 & ~x451 & ~x476 & ~x479 & ~x504 & ~x506 & ~x507 & ~x512 & ~x532 & ~x558 & ~x560 & ~x588 & ~x613 & ~x641 & ~x642 & ~x643 & ~x644 & ~x659 & ~x660 & ~x661 & ~x662 & ~x663 & ~x665 & ~x667 & ~x668 & ~x669 & ~x670 & ~x671 & ~x691 & ~x692 & ~x693 & ~x694 & ~x695 & ~x696 & ~x699 & ~x700 & ~x701 & ~x702 & ~x722 & ~x723 & ~x724 & ~x751 & ~x752 & ~x755 & ~x780 & ~x782 & ~x783;
assign c1232 = ~x46 & ~x67 & ~x96 & ~x234 & ~x262 & ~x351 & ~x362 & ~x417 & ~x468 & ~x476 & ~x543 & ~x571 & ~x598;
assign c1234 =  x67 &  x124 &  x266 &  x351 & ~x0 & ~x109 & ~x144 & ~x368 & ~x389 & ~x394 & ~x481 & ~x533 & ~x618 & ~x669 & ~x693 & ~x694 & ~x696 & ~x721;
assign c1236 =  x711 & ~x2 & ~x6 & ~x53 & ~x55 & ~x59 & ~x77 & ~x79 & ~x88 & ~x89 & ~x117 & ~x118 & ~x138 & ~x144 & ~x164 & ~x165 & ~x166 & ~x167 & ~x169 & ~x172 & ~x173 & ~x195 & ~x196 & ~x200 & ~x201 & ~x223 & ~x224 & ~x226 & ~x228 & ~x229 & ~x247 & ~x251 & ~x277 & ~x278 & ~x279 & ~x280 & ~x282 & ~x283 & ~x304 & ~x311 & ~x312 & ~x332 & ~x333 & ~x334 & ~x336 & ~x337 & ~x339 & ~x340 & ~x341 & ~x342 & ~x361 & ~x364 & ~x365 & ~x366 & ~x367 & ~x369 & ~x393 & ~x394 & ~x395 & ~x419 & ~x421 & ~x422 & ~x424 & ~x447 & ~x448 & ~x449 & ~x450 & ~x451 & ~x452 & ~x477 & ~x478 & ~x479 & ~x501 & ~x503 & ~x534 & ~x535 & ~x559 & ~x586 & ~x589 & ~x611 & ~x612 & ~x613 & ~x614 & ~x615 & ~x616 & ~x639 & ~x640 & ~x669 & ~x670 & ~x673 & ~x674 & ~x687 & ~x688 & ~x699 & ~x700 & ~x718 & ~x722 & ~x723 & ~x725 & ~x727 & ~x728 & ~x729 & ~x748 & ~x749 & ~x750 & ~x759 & ~x761 & ~x762 & ~x763 & ~x774 & ~x776 & ~x778 & ~x780 & ~x782;
assign c1238 = ~x28 & ~x97 & ~x140 & ~x166 & ~x179 & ~x194 & ~x250 & ~x334 & ~x419 & ~x449 & ~x467 & ~x468 & ~x473 & ~x475 & ~x477 & ~x478 & ~x498 & ~x499 & ~x501 & ~x544 & ~x561 & ~x654 & ~x655 & ~x682 & ~x764;
assign c1240 =  x408 & ~x79 & ~x192 & ~x278 & ~x315 & ~x422 & ~x423 & ~x486 & ~x489 & ~x490 & ~x491 & ~x721;
assign c1242 = ~x69 & ~x97 & ~x418 & ~x451 & ~x488 & ~x561 & ~x571 & ~x588 & ~x644 & ~x680 & ~x708 & ~x709;
assign c1244 =  x729 & ~x42;
assign c1246 =  x39 &  x68 &  x96 &  x153 &  x295 &  x296 &  x323 & ~x31 & ~x193 & ~x254 & ~x395 & ~x779;
assign c1248 = ~x0 & ~x2 & ~x23 & ~x26 & ~x27 & ~x28 & ~x30 & ~x31 & ~x47 & ~x53 & ~x56 & ~x57 & ~x58 & ~x78 & ~x83 & ~x85 & ~x110 & ~x112 & ~x133 & ~x140 & ~x143 & ~x166 & ~x167 & ~x168 & ~x170 & ~x172 & ~x190 & ~x193 & ~x194 & ~x199 & ~x222 & ~x223 & ~x228 & ~x249 & ~x250 & ~x251 & ~x252 & ~x254 & ~x255 & ~x273 & ~x279 & ~x284 & ~x285 & ~x308 & ~x309 & ~x312 & ~x313 & ~x334 & ~x335 & ~x341 & ~x363 & ~x364 & ~x366 & ~x367 & ~x396 & ~x397 & ~x421 & ~x425 & ~x426 & ~x447 & ~x448 & ~x450 & ~x451 & ~x453 & ~x454 & ~x455 & ~x474 & ~x475 & ~x477 & ~x479 & ~x481 & ~x482 & ~x483 & ~x488 & ~x490 & ~x501 & ~x508 & ~x511 & ~x528 & ~x529 & ~x530 & ~x531 & ~x534 & ~x536 & ~x557 & ~x560 & ~x562 & ~x564 & ~x584 & ~x585 & ~x587 & ~x588 & ~x590 & ~x591 & ~x616 & ~x617 & ~x619 & ~x631 & ~x643 & ~x673 & ~x674 & ~x698 & ~x699 & ~x700 & ~x725 & ~x726 & ~x728 & ~x750 & ~x752 & ~x753 & ~x754 & ~x755 & ~x779 & ~x780 & ~x781 & ~x782;
assign c1250 =  x9 &  x428 & ~x562 & ~x645;
assign c1252 =  x552 &  x555 & ~x439 & ~x640 & ~x724;
assign c1254 =  x579 &  x581 & ~x445 & ~x599;
assign c1256 =  x409 & ~x0 & ~x5 & ~x26 & ~x53 & ~x54 & ~x58 & ~x60 & ~x82 & ~x110 & ~x115 & ~x138 & ~x141 & ~x142 & ~x194 & ~x196 & ~x197 & ~x225 & ~x249 & ~x253 & ~x278 & ~x308 & ~x339 & ~x361 & ~x365 & ~x389 & ~x391 & ~x394 & ~x396 & ~x397 & ~x417 & ~x420 & ~x421 & ~x424 & ~x425 & ~x426 & ~x427 & ~x449 & ~x450 & ~x453 & ~x454 & ~x478 & ~x490 & ~x506 & ~x508 & ~x520 & ~x536 & ~x589 & ~x590 & ~x617 & ~x695 & ~x696 & ~x751 & ~x752 & ~x757 & ~x782;
assign c1258 =  x760;
assign c1260 =  x680 & ~x144 & ~x198 & ~x200 & ~x201 & ~x256 & ~x287 & ~x456 & ~x646 & ~x689 & ~x720 & ~x728;
assign c1262 =  x607 &  x608 &  x609 & ~x472 & ~x473 & ~x659 & ~x724;
assign c1264 =  x577 &  x742 & ~x190 & ~x254 & ~x449 & ~x562 & ~x660 & ~x689 & ~x695 & ~x726;
assign c1266 =  x406 &  x491 & ~x32 & ~x86 & ~x118 & ~x119 & ~x139 & ~x146 & ~x147 & ~x148 & ~x174 & ~x175 & ~x203 & ~x213 & ~x240 & ~x241 & ~x242 & ~x245 & ~x246 & ~x277 & ~x311 & ~x313 & ~x333 & ~x356 & ~x362 & ~x368 & ~x384 & ~x389 & ~x411 & ~x423 & ~x440 & ~x442 & ~x445 & ~x455 & ~x468 & ~x469 & ~x470 & ~x471 & ~x473 & ~x483 & ~x496 & ~x497 & ~x509 & ~x512 & ~x532 & ~x534 & ~x536 & ~x539 & ~x591 & ~x640 & ~x694 & ~x705 & ~x722;
assign c1268 =  x374 &  x376 &  x380 &  x551 & ~x192 & ~x222 & ~x395 & ~x423 & ~x479 & ~x752;
assign c1270 = ~x0 & ~x24 & ~x52 & ~x55 & ~x58 & ~x59 & ~x81 & ~x85 & ~x108 & ~x136 & ~x139 & ~x140 & ~x143 & ~x146 & ~x164 & ~x166 & ~x168 & ~x170 & ~x171 & ~x203 & ~x223 & ~x225 & ~x229 & ~x249 & ~x253 & ~x254 & ~x311 & ~x313 & ~x339 & ~x342 & ~x368 & ~x388 & ~x394 & ~x396 & ~x398 & ~x399 & ~x417 & ~x419 & ~x428 & ~x447 & ~x487 & ~x489 & ~x502 & ~x505 & ~x531 & ~x532 & ~x560 & ~x563 & ~x585 & ~x614 & ~x671 & ~x689 & ~x690 & ~x691 & ~x698 & ~x719 & ~x746 & ~x747 & ~x749 & ~x750 & ~x751 & ~x756 & ~x775 & ~x777 & ~x779 & ~x781 & ~x783;
assign c1272 =  x687 & ~x56 & ~x78 & ~x79 & ~x107 & ~x142 & ~x251 & ~x253 & ~x331 & ~x372 & ~x389 & ~x400 & ~x423 & ~x471 & ~x605 & ~x633 & ~x664 & ~x710 & ~x722 & ~x723 & ~x739 & ~x754;
assign c1274 = ~x5 & ~x6 & ~x21 & ~x24 & ~x69 & ~x84 & ~x166 & ~x193 & ~x250 & ~x306 & ~x308 & ~x335 & ~x336 & ~x352 & ~x361 & ~x362 & ~x391 & ~x417 & ~x419 & ~x448 & ~x472 & ~x474 & ~x504 & ~x523 & ~x528 & ~x532 & ~x534 & ~x551 & ~x553 & ~x738 & ~x780;
assign c1276 = ~x1 & ~x3 & ~x4 & ~x18 & ~x20 & ~x22 & ~x25 & ~x26 & ~x28 & ~x29 & ~x32 & ~x33 & ~x47 & ~x49 & ~x51 & ~x53 & ~x59 & ~x71 & ~x74 & ~x76 & ~x79 & ~x80 & ~x84 & ~x87 & ~x94 & ~x104 & ~x106 & ~x107 & ~x110 & ~x112 & ~x130 & ~x132 & ~x133 & ~x134 & ~x135 & ~x136 & ~x137 & ~x139 & ~x140 & ~x142 & ~x143 & ~x160 & ~x165 & ~x168 & ~x169 & ~x170 & ~x191 & ~x199 & ~x218 & ~x220 & ~x221 & ~x222 & ~x224 & ~x226 & ~x227 & ~x245 & ~x250 & ~x251 & ~x253 & ~x282 & ~x307 & ~x309 & ~x310 & ~x311 & ~x320 & ~x333 & ~x336 & ~x339 & ~x341 & ~x360 & ~x363 & ~x365 & ~x366 & ~x391 & ~x392 & ~x396 & ~x418 & ~x419 & ~x423 & ~x446 & ~x448 & ~x476 & ~x478 & ~x479 & ~x499 & ~x500 & ~x504 & ~x505 & ~x507 & ~x509 & ~x510 & ~x529 & ~x530 & ~x531 & ~x532 & ~x533 & ~x537 & ~x565 & ~x587 & ~x591 & ~x613 & ~x620 & ~x698 & ~x700 & ~x701 & ~x726 & ~x730 & ~x756 & ~x759 & ~x781;
assign c1278 =  x569 & ~x110 & ~x225 & ~x237 & ~x435 & ~x479 & ~x533 & ~x564 & ~x615 & ~x682 & ~x709;
assign c1280 =  x70 &  x269 &  x383 & ~x55 & ~x142 & ~x170 & ~x277 & ~x283 & ~x309 & ~x335 & ~x341 & ~x365 & ~x389 & ~x502 & ~x535 & ~x564 & ~x585 & ~x586 & ~x614 & ~x729;
assign c1282 =  x409 & ~x1 & ~x60 & ~x80 & ~x87 & ~x105 & ~x106 & ~x114 & ~x115 & ~x133 & ~x135 & ~x190 & ~x194 & ~x222 & ~x226 & ~x253 & ~x278 & ~x305 & ~x310 & ~x336 & ~x337 & ~x340 & ~x366 & ~x367 & ~x394 & ~x416 & ~x421 & ~x447 & ~x454 & ~x487 & ~x489 & ~x492 & ~x509 & ~x563 & ~x586 & ~x644 & ~x669 & ~x672 & ~x674 & ~x702 & ~x723 & ~x783;
assign c1284 =  x713 & ~x9 & ~x176 & ~x193 & ~x194 & ~x196 & ~x199 & ~x202 & ~x204 & ~x279 & ~x306 & ~x337 & ~x391 & ~x422 & ~x544 & ~x586 & ~x659 & ~x691 & ~x724;
assign c1286 = ~x21 & ~x45 & ~x84 & ~x115 & ~x119 & ~x131 & ~x143 & ~x159 & ~x172 & ~x185 & ~x190 & ~x197 & ~x212 & ~x213 & ~x225 & ~x229 & ~x239 & ~x240 & ~x250 & ~x269 & ~x271 & ~x277 & ~x284 & ~x285 & ~x336 & ~x339 & ~x341 & ~x342 & ~x360 & ~x369 & ~x381 & ~x392 & ~x410 & ~x417 & ~x421 & ~x426 & ~x438 & ~x451 & ~x454 & ~x455 & ~x466 & ~x467 & ~x474 & ~x495 & ~x525 & ~x552 & ~x562 & ~x584 & ~x611 & ~x618 & ~x665 & ~x672 & ~x702 & ~x728 & ~x749 & ~x751 & ~x777;
assign c1288 =  x99 &  x127 &  x269 &  x297 & ~x32 & ~x134 & ~x161 & ~x166 & ~x193 & ~x194 & ~x306 & ~x341 & ~x363 & ~x369 & ~x450 & ~x451 & ~x533 & ~x669 & ~x702 & ~x720 & ~x724 & ~x760 & ~x764 & ~x782;
assign c1290 =  x739 & ~x94 & ~x109 & ~x115 & ~x117 & ~x171 & ~x250 & ~x258 & ~x314 & ~x330 & ~x363 & ~x506 & ~x694 & ~x698 & ~x701 & ~x717 & ~x720 & ~x728 & ~x774 & ~x775;
assign c1292 =  x712 & ~x24 & ~x28 & ~x79 & ~x84 & ~x87 & ~x103 & ~x115 & ~x140 & ~x143 & ~x169 & ~x171 & ~x251 & ~x277 & ~x278 & ~x305 & ~x307 & ~x332 & ~x333 & ~x334 & ~x361 & ~x363 & ~x389 & ~x419 & ~x423 & ~x450 & ~x474 & ~x477 & ~x501 & ~x506 & ~x507 & ~x534 & ~x558 & ~x562 & ~x599 & ~x600 & ~x629 & ~x630 & ~x658 & ~x659 & ~x660 & ~x670 & ~x692 & ~x695 & ~x756 & ~x782;
assign c1294 =  x295 &  x352 & ~x4 & ~x5 & ~x25 & ~x30 & ~x81 & ~x109 & ~x112 & ~x165 & ~x198 & ~x222 & ~x250 & ~x305 & ~x309 & ~x311 & ~x328 & ~x332 & ~x337 & ~x358 & ~x364 & ~x367 & ~x387 & ~x389 & ~x390 & ~x394 & ~x425 & ~x449 & ~x450 & ~x474 & ~x525 & ~x563 & ~x590 & ~x591 & ~x612 & ~x638 & ~x666 & ~x667 & ~x669 & ~x675 & ~x690 & ~x693 & ~x694 & ~x719 & ~x722 & ~x749 & ~x752 & ~x780;
assign c1296 = ~x21 & ~x25 & ~x27 & ~x57 & ~x81 & ~x82 & ~x83 & ~x84 & ~x109 & ~x110 & ~x111 & ~x137 & ~x138 & ~x166 & ~x222 & ~x223 & ~x225 & ~x250 & ~x281 & ~x307 & ~x325 & ~x335 & ~x363 & ~x390 & ~x446 & ~x448 & ~x449 & ~x468 & ~x472 & ~x474 & ~x477 & ~x495 & ~x499 & ~x502 & ~x505 & ~x506 & ~x517 & ~x524 & ~x525 & ~x526 & ~x528 & ~x533 & ~x559 & ~x781;
assign c1298 = ~x2 & ~x4 & ~x22 & ~x28 & ~x32 & ~x51 & ~x52 & ~x54 & ~x58 & ~x60 & ~x79 & ~x80 & ~x83 & ~x84 & ~x86 & ~x107 & ~x108 & ~x110 & ~x112 & ~x114 & ~x136 & ~x137 & ~x138 & ~x139 & ~x142 & ~x165 & ~x167 & ~x168 & ~x198 & ~x224 & ~x226 & ~x252 & ~x254 & ~x278 & ~x304 & ~x308 & ~x309 & ~x333 & ~x335 & ~x336 & ~x337 & ~x362 & ~x365 & ~x366 & ~x389 & ~x391 & ~x392 & ~x394 & ~x420 & ~x421 & ~x445 & ~x446 & ~x447 & ~x448 & ~x476 & ~x501 & ~x503 & ~x504 & ~x515 & ~x530 & ~x586 & ~x589 & ~x617 & ~x629 & ~x630 & ~x632 & ~x633 & ~x640 & ~x641 & ~x642 & ~x658 & ~x661 & ~x662 & ~x665 & ~x666 & ~x668 & ~x673 & ~x693 & ~x694 & ~x695 & ~x697 & ~x700 & ~x701 & ~x722 & ~x725 & ~x726 & ~x752 & ~x753 & ~x754 & ~x779;
assign c1300 =  x663 &  x695 & ~x183;
assign c1302 =  x677 & ~x324 & ~x563 & ~x588 & ~x590 & ~x591;
assign c1304 =  x96 &  x319 &  x321 & ~x48 & ~x106 & ~x109 & ~x111 & ~x114 & ~x143 & ~x222 & ~x223 & ~x251 & ~x280 & ~x366 & ~x368 & ~x400 & ~x426 & ~x429 & ~x430 & ~x475 & ~x477 & ~x506 & ~x533 & ~x617 & ~x730 & ~x780 & ~x782;
assign c1306 =  x483 & ~x16 & ~x38 & ~x39 & ~x110 & ~x137 & ~x166 & ~x222 & ~x251 & ~x416 & ~x417 & ~x444 & ~x445 & ~x446 & ~x467 & ~x468 & ~x469 & ~x514 & ~x652 & ~x679 & ~x734;
assign c1308 = ~x16 & ~x20 & ~x23 & ~x24 & ~x28 & ~x47 & ~x54 & ~x55 & ~x56 & ~x57 & ~x71 & ~x74 & ~x77 & ~x80 & ~x83 & ~x102 & ~x104 & ~x106 & ~x128 & ~x137 & ~x142 & ~x143 & ~x164 & ~x165 & ~x167 & ~x168 & ~x192 & ~x197 & ~x224 & ~x249 & ~x280 & ~x281 & ~x305 & ~x307 & ~x335 & ~x337 & ~x364 & ~x416 & ~x421 & ~x444 & ~x445 & ~x469 & ~x477 & ~x504 & ~x505 & ~x532 & ~x652 & ~x688 & ~x706 & ~x718 & ~x724 & ~x725 & ~x726 & ~x727 & ~x735 & ~x746 & ~x750 & ~x751 & ~x752 & ~x763 & ~x780 & ~x783;
assign c1310 =  x183 &  x325 & ~x16 & ~x27 & ~x28 & ~x44 & ~x83 & ~x105 & ~x107 & ~x142 & ~x171 & ~x172 & ~x224 & ~x277 & ~x278 & ~x281 & ~x305 & ~x307 & ~x312 & ~x394 & ~x396 & ~x418 & ~x427 & ~x451 & ~x480 & ~x501 & ~x504 & ~x646 & ~x666 & ~x672 & ~x693 & ~x697 & ~x698 & ~x702 & ~x730 & ~x733 & ~x753 & ~x781 & ~x783;
assign c1312 =  x607 &  x610 & ~x72 & ~x723;
assign c1314 =  x375 & ~x0 & ~x19 & ~x20 & ~x21 & ~x24 & ~x25 & ~x26 & ~x27 & ~x29 & ~x30 & ~x47 & ~x51 & ~x53 & ~x54 & ~x56 & ~x57 & ~x77 & ~x78 & ~x79 & ~x80 & ~x83 & ~x84 & ~x106 & ~x108 & ~x110 & ~x111 & ~x115 & ~x119 & ~x133 & ~x135 & ~x137 & ~x138 & ~x140 & ~x141 & ~x143 & ~x162 & ~x165 & ~x166 & ~x167 & ~x188 & ~x193 & ~x194 & ~x196 & ~x199 & ~x200 & ~x201 & ~x222 & ~x223 & ~x224 & ~x226 & ~x228 & ~x247 & ~x249 & ~x251 & ~x252 & ~x253 & ~x254 & ~x255 & ~x256 & ~x278 & ~x279 & ~x280 & ~x281 & ~x282 & ~x283 & ~x284 & ~x305 & ~x306 & ~x307 & ~x308 & ~x310 & ~x332 & ~x333 & ~x338 & ~x363 & ~x364 & ~x367 & ~x391 & ~x393 & ~x394 & ~x418 & ~x420 & ~x421 & ~x422 & ~x426 & ~x444 & ~x449 & ~x450 & ~x452 & ~x454 & ~x455 & ~x456 & ~x457 & ~x473 & ~x477 & ~x482 & ~x483 & ~x484 & ~x485 & ~x486 & ~x487 & ~x502 & ~x503 & ~x504 & ~x505 & ~x506 & ~x507 & ~x528 & ~x529 & ~x530 & ~x533 & ~x558 & ~x561 & ~x589 & ~x614 & ~x641 & ~x642 & ~x643 & ~x646 & ~x669 & ~x673 & ~x674 & ~x698 & ~x699 & ~x700 & ~x724 & ~x726 & ~x727 & ~x730 & ~x752 & ~x753 & ~x754 & ~x761 & ~x780 & ~x781 & ~x782 & ~x783;
assign c1316 =  x238 & ~x53 & ~x116 & ~x168 & ~x171 & ~x192 & ~x222 & ~x224 & ~x228 & ~x249 & ~x306 & ~x310 & ~x331 & ~x335 & ~x338 & ~x341 & ~x342 & ~x364 & ~x371 & ~x392 & ~x420 & ~x422 & ~x423 & ~x445 & ~x448 & ~x449 & ~x473 & ~x478 & ~x501 & ~x560 & ~x561 & ~x562 & ~x586 & ~x616 & ~x629 & ~x659 & ~x669 & ~x673 & ~x690 & ~x694 & ~x696 & ~x703 & ~x726 & ~x754 & ~x777;
assign c1318 =  x655 & ~x5 & ~x141 & ~x174 & ~x189 & ~x193 & ~x212 & ~x214 & ~x338 & ~x381 & ~x417 & ~x425 & ~x438 & ~x479 & ~x503 & ~x528 & ~x554 & ~x562 & ~x609 & ~x752 & ~x777;
assign c1320 =  x295 &  x352 &  x465 & ~x29 & ~x34 & ~x48 & ~x59 & ~x76 & ~x168 & ~x202 & ~x220 & ~x230 & ~x285 & ~x360 & ~x367 & ~x384 & ~x481 & ~x499 & ~x510 & ~x581 & ~x619 & ~x621 & ~x639 & ~x674 & ~x678 & ~x693 & ~x700 & ~x719 & ~x733 & ~x734 & ~x758;
assign c1322 =  x674 & ~x40 & ~x417 & ~x442 & ~x444 & ~x571 & ~x706;
assign c1324 =  x211 &  x353 & ~x1 & ~x15 & ~x16 & ~x17 & ~x24 & ~x25 & ~x28 & ~x43 & ~x44 & ~x81 & ~x111 & ~x113 & ~x137 & ~x138 & ~x141 & ~x164 & ~x165 & ~x166 & ~x168 & ~x192 & ~x193 & ~x195 & ~x221 & ~x222 & ~x223 & ~x224 & ~x249 & ~x250 & ~x277 & ~x278 & ~x280 & ~x281 & ~x305 & ~x306 & ~x307 & ~x308 & ~x309 & ~x332 & ~x360 & ~x361 & ~x362 & ~x364 & ~x390 & ~x418 & ~x420 & ~x421 & ~x448 & ~x450 & ~x473 & ~x475 & ~x477 & ~x506 & ~x588 & ~x664 & ~x668 & ~x670 & ~x692 & ~x694 & ~x696 & ~x697 & ~x698 & ~x699 & ~x723 & ~x724 & ~x725 & ~x726 & ~x729 & ~x751 & ~x753 & ~x763 & ~x764 & ~x777 & ~x780;
assign c1326 =  x146 &  x580;
assign c1328 = ~x12 & ~x14 & ~x22 & ~x54 & ~x56 & ~x69 & ~x96 & ~x97 & ~x418 & ~x449 & ~x476 & ~x515 & ~x541 & ~x542 & ~x678 & ~x705 & ~x760;
assign c1330 = ~x2 & ~x8 & ~x19 & ~x28 & ~x36 & ~x48 & ~x49 & ~x54 & ~x75 & ~x76 & ~x77 & ~x83 & ~x86 & ~x89 & ~x109 & ~x111 & ~x115 & ~x140 & ~x167 & ~x278 & ~x290 & ~x333 & ~x335 & ~x389 & ~x393 & ~x419 & ~x420 & ~x433 & ~x448 & ~x476 & ~x600 & ~x690 & ~x699 & ~x700 & ~x702 & ~x722 & ~x725 & ~x747 & ~x753 & ~x763 & ~x775;
assign c1332 =  x322 &  x436 & ~x53 & ~x59 & ~x81 & ~x143 & ~x175 & ~x186 & ~x201 & ~x211 & ~x213 & ~x214 & ~x243 & ~x253 & ~x270 & ~x272 & ~x276 & ~x286 & ~x314 & ~x332 & ~x343 & ~x356 & ~x357 & ~x384 & ~x427 & ~x444 & ~x448 & ~x503 & ~x526 & ~x583 & ~x586 & ~x639 & ~x648;
assign c1334 = ~x106 & ~x115 & ~x192 & ~x273 & ~x286 & ~x327 & ~x388 & ~x424 & ~x428 & ~x446 & ~x509 & ~x512 & ~x517 & ~x532 & ~x538 & ~x575 & ~x691 & ~x697 & ~x719 & ~x776;
assign c1336 =  x145 &  x748;
assign c1338 = ~x18 & ~x78 & ~x83 & ~x109 & ~x172 & ~x194 & ~x305 & ~x311 & ~x349 & ~x367 & ~x368 & ~x373 & ~x374 & ~x375 & ~x391 & ~x423 & ~x424 & ~x507 & ~x576 & ~x577 & ~x584 & ~x605 & ~x608 & ~x641 & ~x724;
assign c1340 = ~x0 & ~x17 & ~x53 & ~x55 & ~x96 & ~x124 & ~x138 & ~x139 & ~x195 & ~x196 & ~x197 & ~x198 & ~x212 & ~x222 & ~x223 & ~x251 & ~x278 & ~x306 & ~x334 & ~x391 & ~x417 & ~x418 & ~x446 & ~x447 & ~x474 & ~x478 & ~x479 & ~x507 & ~x517 & ~x532 & ~x561 & ~x599 & ~x736 & ~x756 & ~x763;
assign c1342 = ~x17 & ~x21 & ~x97 & ~x233 & ~x307 & ~x468 & ~x569 & ~x678 & ~x681 & ~x706 & ~x733 & ~x763;
assign c1344 = ~x5 & ~x25 & ~x31 & ~x34 & ~x56 & ~x84 & ~x106 & ~x107 & ~x134 & ~x136 & ~x143 & ~x168 & ~x170 & ~x199 & ~x221 & ~x226 & ~x228 & ~x255 & ~x275 & ~x334 & ~x338 & ~x340 & ~x374 & ~x391 & ~x392 & ~x393 & ~x400 & ~x401 & ~x402 & ~x403 & ~x406 & ~x422 & ~x423 & ~x444 & ~x530 & ~x558 & ~x605 & ~x614 & ~x615 & ~x634 & ~x636 & ~x641 & ~x645 & ~x662 & ~x670 & ~x694 & ~x725 & ~x760;
assign c1346 =  x380 &  x551 & ~x0 & ~x1 & ~x2 & ~x24 & ~x27 & ~x30 & ~x53 & ~x56 & ~x57 & ~x79 & ~x80 & ~x81 & ~x82 & ~x85 & ~x107 & ~x108 & ~x109 & ~x112 & ~x136 & ~x137 & ~x138 & ~x139 & ~x163 & ~x164 & ~x167 & ~x193 & ~x195 & ~x196 & ~x220 & ~x221 & ~x223 & ~x224 & ~x225 & ~x226 & ~x249 & ~x250 & ~x253 & ~x277 & ~x281 & ~x306 & ~x307 & ~x334 & ~x335 & ~x361 & ~x362 & ~x389 & ~x391 & ~x392 & ~x394 & ~x416 & ~x417 & ~x419 & ~x421 & ~x422 & ~x423 & ~x424 & ~x425 & ~x443 & ~x444 & ~x445 & ~x448 & ~x449 & ~x477 & ~x479 & ~x503 & ~x504 & ~x532 & ~x533 & ~x534 & ~x588 & ~x640 & ~x642 & ~x667 & ~x668 & ~x669 & ~x670 & ~x671 & ~x694 & ~x695 & ~x696 & ~x699 & ~x700 & ~x721 & ~x722 & ~x723 & ~x724 & ~x727 & ~x728 & ~x729 & ~x731 & ~x751 & ~x752 & ~x756 & ~x778 & ~x780 & ~x781 & ~x782 & ~x783;
assign c1348 =  x217 &  x537;
assign c1350 =  x241 &  x269 &  x411 & ~x24 & ~x53 & ~x87 & ~x250 & ~x284 & ~x311 & ~x367 & ~x398 & ~x399 & ~x477 & ~x502 & ~x589 & ~x722 & ~x755;
assign c1352 =  x713 &  x742 & ~x79 & ~x91 & ~x147 & ~x203 & ~x204 & ~x231 & ~x344 & ~x372 & ~x373 & ~x391 & ~x709 & ~x738 & ~x767 & ~x776;
assign c1354 =  x268 & ~x22 & ~x51 & ~x56 & ~x57 & ~x119 & ~x137 & ~x164 & ~x165 & ~x222 & ~x225 & ~x227 & ~x275 & ~x282 & ~x362 & ~x391 & ~x404 & ~x406 & ~x445 & ~x447 & ~x476 & ~x502 & ~x531 & ~x548 & ~x557 & ~x560 & ~x616 & ~x665 & ~x669 & ~x694 & ~x697 & ~x699 & ~x701 & ~x735 & ~x749 & ~x755 & ~x761;
assign c1356 = ~x6 & ~x89 & ~x90 & ~x105 & ~x142 & ~x155 & ~x184 & ~x226 & ~x270 & ~x288 & ~x298 & ~x316 & ~x342 & ~x355 & ~x369 & ~x370 & ~x400 & ~x478 & ~x497 & ~x524 & ~x525 & ~x526 & ~x538 & ~x554 & ~x723 & ~x754;
assign c1358 =  x349 &  x350 & ~x52 & ~x84 & ~x137 & ~x167 & ~x195 & ~x221 & ~x250 & ~x276 & ~x282 & ~x305 & ~x311 & ~x333 & ~x338 & ~x420 & ~x451 & ~x457 & ~x458 & ~x459 & ~x460 & ~x461 & ~x481 & ~x484 & ~x644 & ~x663 & ~x664 & ~x668 & ~x693 & ~x694 & ~x697 & ~x699 & ~x724 & ~x751 & ~x765 & ~x779;
assign c1360 = ~x25 & ~x53 & ~x58 & ~x81 & ~x82 & ~x85 & ~x86 & ~x104 & ~x106 & ~x110 & ~x115 & ~x137 & ~x138 & ~x139 & ~x143 & ~x144 & ~x165 & ~x170 & ~x171 & ~x172 & ~x195 & ~x199 & ~x200 & ~x226 & ~x228 & ~x250 & ~x254 & ~x280 & ~x307 & ~x338 & ~x362 & ~x364 & ~x367 & ~x391 & ~x395 & ~x397 & ~x398 & ~x420 & ~x422 & ~x423 & ~x427 & ~x428 & ~x429 & ~x430 & ~x431 & ~x433 & ~x451 & ~x479 & ~x505 & ~x506 & ~x560 & ~x574 & ~x575 & ~x576 & ~x588 & ~x606 & ~x617 & ~x670 & ~x674 & ~x696 & ~x699 & ~x701 & ~x724 & ~x728 & ~x751 & ~x752 & ~x757;
assign c1362 = ~x31 & ~x116 & ~x128 & ~x139 & ~x142 & ~x145 & ~x147 & ~x162 & ~x168 & ~x173 & ~x174 & ~x200 & ~x218 & ~x229 & ~x242 & ~x243 & ~x250 & ~x270 & ~x271 & ~x277 & ~x286 & ~x299 & ~x310 & ~x340 & ~x341 & ~x342 & ~x365 & ~x366 & ~x368 & ~x390 & ~x391 & ~x398 & ~x400 & ~x423 & ~x426 & ~x448 & ~x450 & ~x454 & ~x455 & ~x482 & ~x484 & ~x485 & ~x486 & ~x487 & ~x488 & ~x500 & ~x502 & ~x529 & ~x563 & ~x611 & ~x614 & ~x617 & ~x618 & ~x619 & ~x645 & ~x674 & ~x675 & ~x702 & ~x724 & ~x731 & ~x753 & ~x755 & ~x757;
assign c1364 = ~x4 & ~x23 & ~x28 & ~x84 & ~x107 & ~x115 & ~x131 & ~x143 & ~x165 & ~x172 & ~x201 & ~x222 & ~x225 & ~x252 & ~x256 & ~x306 & ~x310 & ~x311 & ~x336 & ~x338 & ~x364 & ~x368 & ~x394 & ~x397 & ~x399 & ~x419 & ~x422 & ~x425 & ~x426 & ~x447 & ~x476 & ~x530 & ~x535 & ~x588 & ~x613 & ~x657 & ~x658 & ~x671 & ~x686 & ~x687 & ~x688 & ~x717 & ~x723 & ~x745 & ~x761 & ~x779;
assign c1366 =  x96 & ~x0 & ~x43 & ~x72 & ~x105 & ~x132 & ~x241 & ~x242 & ~x243 & ~x271 & ~x298 & ~x364 & ~x382 & ~x383 & ~x399 & ~x439 & ~x441 & ~x447 & ~x503 & ~x527 & ~x559 & ~x763 & ~x782;
assign c1368 = ~x31 & ~x33 & ~x76 & ~x78 & ~x83 & ~x85 & ~x88 & ~x104 & ~x105 & ~x113 & ~x114 & ~x116 & ~x139 & ~x140 & ~x143 & ~x144 & ~x168 & ~x170 & ~x197 & ~x198 & ~x199 & ~x227 & ~x252 & ~x255 & ~x280 & ~x281 & ~x306 & ~x311 & ~x312 & ~x314 & ~x341 & ~x360 & ~x363 & ~x369 & ~x388 & ~x397 & ~x399 & ~x427 & ~x428 & ~x429 & ~x430 & ~x431 & ~x432 & ~x433 & ~x449 & ~x450 & ~x531 & ~x532 & ~x559 & ~x589 & ~x604 & ~x605 & ~x663 & ~x670 & ~x695 & ~x696 & ~x700 & ~x701 & ~x722 & ~x729 & ~x733 & ~x735 & ~x753 & ~x754 & ~x756;
assign c1370 =  x407 &  x492 &  x548 & ~x31 & ~x55 & ~x75 & ~x88 & ~x108 & ~x109 & ~x115 & ~x137 & ~x138 & ~x147 & ~x163 & ~x175 & ~x248 & ~x249 & ~x270 & ~x327 & ~x330 & ~x331 & ~x355 & ~x383 & ~x385 & ~x393 & ~x395 & ~x417 & ~x445 & ~x479 & ~x505 & ~x510 & ~x553 & ~x554 & ~x558 & ~x586 & ~x614 & ~x619 & ~x642 & ~x645 & ~x649 & ~x650 & ~x692 & ~x695 & ~x701 & ~x719 & ~x777 & ~x778 & ~x783;
assign c1372 = ~x0 & ~x53 & ~x56 & ~x75 & ~x81 & ~x82 & ~x87 & ~x90 & ~x105 & ~x111 & ~x112 & ~x113 & ~x115 & ~x116 & ~x135 & ~x144 & ~x167 & ~x194 & ~x198 & ~x202 & ~x222 & ~x224 & ~x227 & ~x229 & ~x230 & ~x254 & ~x255 & ~x258 & ~x278 & ~x283 & ~x287 & ~x305 & ~x310 & ~x311 & ~x312 & ~x341 & ~x342 & ~x348 & ~x367 & ~x369 & ~x371 & ~x372 & ~x373 & ~x374 & ~x375 & ~x396 & ~x445 & ~x446 & ~x473 & ~x474 & ~x477 & ~x478 & ~x504 & ~x505 & ~x507 & ~x534 & ~x557 & ~x560 & ~x587 & ~x611 & ~x614 & ~x615 & ~x642 & ~x661 & ~x670 & ~x671 & ~x672 & ~x697 & ~x698 & ~x700 & ~x701 & ~x720 & ~x730 & ~x750 & ~x777;
assign c1374 =  x672;
assign c1376 =  x354 &  x524 &  x553 & ~x137 & ~x139 & ~x168 & ~x169 & ~x280 & ~x281 & ~x306 & ~x366 & ~x392 & ~x393 & ~x395 & ~x417 & ~x425 & ~x446 & ~x451 & ~x477 & ~x478 & ~x502 & ~x504 & ~x505 & ~x669 & ~x752;
assign c1378 = ~x19 & ~x72 & ~x85 & ~x89 & ~x91 & ~x107 & ~x115 & ~x120 & ~x132 & ~x172 & ~x176 & ~x187 & ~x203 & ~x232 & ~x275 & ~x304 & ~x316 & ~x339 & ~x367 & ~x373 & ~x374 & ~x391 & ~x450 & ~x557 & ~x564 & ~x589 & ~x614 & ~x648 & ~x649 & ~x690 & ~x694 & ~x732 & ~x747 & ~x754;
assign c1380 =  x593 & ~x24 & ~x52 & ~x79 & ~x108 & ~x136 & ~x166 & ~x195 & ~x222 & ~x362 & ~x363 & ~x418 & ~x419 & ~x505 & ~x625 & ~x651 & ~x652 & ~x707 & ~x708 & ~x733 & ~x748 & ~x779 & ~x780 & ~x782;
assign c1382 = ~x1 & ~x25 & ~x28 & ~x30 & ~x53 & ~x54 & ~x55 & ~x57 & ~x60 & ~x78 & ~x79 & ~x80 & ~x85 & ~x86 & ~x87 & ~x88 & ~x106 & ~x107 & ~x110 & ~x111 & ~x112 & ~x114 & ~x116 & ~x137 & ~x138 & ~x168 & ~x169 & ~x170 & ~x171 & ~x172 & ~x189 & ~x193 & ~x197 & ~x198 & ~x200 & ~x217 & ~x224 & ~x225 & ~x249 & ~x251 & ~x253 & ~x254 & ~x256 & ~x278 & ~x282 & ~x284 & ~x287 & ~x311 & ~x312 & ~x337 & ~x341 & ~x360 & ~x361 & ~x363 & ~x364 & ~x365 & ~x367 & ~x368 & ~x369 & ~x390 & ~x391 & ~x393 & ~x395 & ~x396 & ~x419 & ~x420 & ~x423 & ~x424 & ~x425 & ~x426 & ~x445 & ~x449 & ~x451 & ~x452 & ~x453 & ~x454 & ~x475 & ~x476 & ~x477 & ~x480 & ~x482 & ~x483 & ~x485 & ~x491 & ~x504 & ~x505 & ~x509 & ~x511 & ~x514 & ~x515 & ~x519 & ~x533 & ~x559 & ~x560 & ~x586 & ~x587 & ~x588 & ~x617 & ~x643 & ~x669 & ~x697 & ~x699 & ~x725 & ~x726 & ~x728 & ~x730 & ~x747 & ~x749 & ~x752 & ~x755 & ~x757 & ~x758 & ~x759;
assign c1384 =  x759 & ~x152 & ~x393 & ~x489 & ~x517 & ~x590 & ~x614;
assign c1386 =  x41 & ~x27 & ~x29 & ~x79 & ~x164 & ~x167 & ~x173 & ~x202 & ~x225 & ~x226 & ~x228 & ~x247 & ~x281 & ~x283 & ~x335 & ~x343 & ~x369 & ~x372 & ~x374 & ~x377 & ~x395 & ~x402 & ~x449 & ~x617 & ~x635 & ~x668 & ~x674 & ~x702 & ~x726 & ~x729 & ~x763;
assign c1388 =  x90 &  x702;
assign c1390 =  x577 & ~x3 & ~x53 & ~x60 & ~x81 & ~x87 & ~x109 & ~x111 & ~x137 & ~x142 & ~x166 & ~x172 & ~x173 & ~x193 & ~x195 & ~x199 & ~x200 & ~x202 & ~x222 & ~x246 & ~x251 & ~x252 & ~x256 & ~x276 & ~x280 & ~x281 & ~x282 & ~x283 & ~x303 & ~x306 & ~x310 & ~x311 & ~x338 & ~x339 & ~x362 & ~x367 & ~x394 & ~x417 & ~x421 & ~x449 & ~x451 & ~x452 & ~x475 & ~x501 & ~x558 & ~x561 & ~x588 & ~x591 & ~x614 & ~x617 & ~x645 & ~x646 & ~x647 & ~x660 & ~x663 & ~x669 & ~x676 & ~x691 & ~x692 & ~x693 & ~x695 & ~x699 & ~x701 & ~x722 & ~x723 & ~x724 & ~x725 & ~x727 & ~x751 & ~x752 & ~x764 & ~x782;
assign c1392 =  x350 &  x378 &  x407 &  x436 &  x464 &  x521 & ~x118 & ~x147 & ~x176 & ~x193 & ~x330 & ~x341 & ~x361 & ~x440 & ~x478 & ~x479 & ~x511 & ~x621 & ~x694;
assign c1394 =  x239 & ~x29 & ~x172 & ~x314 & ~x361 & ~x420 & ~x506 & ~x518 & ~x576 & ~x646 & ~x720 & ~x752;
assign c1396 =  x272 &  x409 & ~x43 & ~x44 & ~x194 & ~x249 & ~x250 & ~x725;
assign c1398 =  x68 &  x210 &  x295 & ~x59 & ~x71 & ~x85 & ~x105 & ~x136 & ~x224 & ~x248 & ~x277 & ~x333 & ~x501 & ~x666 & ~x723 & ~x724 & ~x730 & ~x749;
assign c1400 =  x581 &  x584 & ~x417 & ~x696;
assign c1402 = ~x5 & ~x17 & ~x18 & ~x26 & ~x27 & ~x44 & ~x56 & ~x72 & ~x73 & ~x75 & ~x81 & ~x82 & ~x85 & ~x110 & ~x113 & ~x138 & ~x141 & ~x167 & ~x168 & ~x169 & ~x197 & ~x224 & ~x249 & ~x253 & ~x254 & ~x276 & ~x279 & ~x281 & ~x308 & ~x333 & ~x335 & ~x363 & ~x390 & ~x391 & ~x393 & ~x417 & ~x418 & ~x419 & ~x446 & ~x448 & ~x449 & ~x450 & ~x475 & ~x478 & ~x499 & ~x501 & ~x502 & ~x503 & ~x504 & ~x505 & ~x506 & ~x507 & ~x524 & ~x527 & ~x529 & ~x531 & ~x532 & ~x534 & ~x551 & ~x552 & ~x553 & ~x554 & ~x555 & ~x556 & ~x557 & ~x558 & ~x559 & ~x561 & ~x562 & ~x563 & ~x583 & ~x584 & ~x585 & ~x586 & ~x600 & ~x617 & ~x618 & ~x682 & ~x709 & ~x710 & ~x727 & ~x736 & ~x738 & ~x763;
assign c1404 = ~x16 & ~x21 & ~x26 & ~x28 & ~x31 & ~x54 & ~x55 & ~x57 & ~x83 & ~x85 & ~x110 & ~x112 & ~x114 & ~x115 & ~x137 & ~x138 & ~x141 & ~x142 & ~x144 & ~x166 & ~x167 & ~x168 & ~x170 & ~x171 & ~x198 & ~x221 & ~x222 & ~x224 & ~x225 & ~x226 & ~x250 & ~x253 & ~x254 & ~x278 & ~x279 & ~x306 & ~x307 & ~x310 & ~x333 & ~x334 & ~x362 & ~x365 & ~x390 & ~x392 & ~x393 & ~x417 & ~x419 & ~x420 & ~x422 & ~x423 & ~x446 & ~x447 & ~x450 & ~x451 & ~x452 & ~x473 & ~x474 & ~x475 & ~x479 & ~x502 & ~x503 & ~x504 & ~x507 & ~x508 & ~x528 & ~x529 & ~x530 & ~x533 & ~x534 & ~x535 & ~x536 & ~x551 & ~x552 & ~x553 & ~x554 & ~x555 & ~x556 & ~x558 & ~x559 & ~x560 & ~x562 & ~x563 & ~x564 & ~x580 & ~x581 & ~x582 & ~x583 & ~x584 & ~x585 & ~x586 & ~x590 & ~x591 & ~x618 & ~x643 & ~x670 & ~x671 & ~x673 & ~x698 & ~x709 & ~x710 & ~x711 & ~x725 & ~x726 & ~x727 & ~x728 & ~x736 & ~x737 & ~x738 & ~x752 & ~x755 & ~x756 & ~x763 & ~x764 & ~x765 & ~x766 & ~x774;
assign c1406 =  x181 &  x323 &  x436 & ~x43 & ~x44 & ~x72 & ~x194 & ~x220 & ~x229 & ~x230 & ~x389 & ~x398 & ~x611 & ~x646 & ~x723;
assign c1408 =  x212 &  x354 &  x411 & ~x22 & ~x30 & ~x51 & ~x54 & ~x55 & ~x76 & ~x77 & ~x78 & ~x79 & ~x82 & ~x87 & ~x105 & ~x107 & ~x111 & ~x115 & ~x194 & ~x222 & ~x252 & ~x254 & ~x276 & ~x279 & ~x280 & ~x281 & ~x282 & ~x308 & ~x310 & ~x335 & ~x336 & ~x337 & ~x362 & ~x366 & ~x368 & ~x390 & ~x391 & ~x394 & ~x395 & ~x397 & ~x422 & ~x423 & ~x448 & ~x450 & ~x478 & ~x504 & ~x532 & ~x645 & ~x669 & ~x697 & ~x698 & ~x699 & ~x725 & ~x729 & ~x753 & ~x755 & ~x780;
assign c1410 = ~x25 & ~x115 & ~x168 & ~x304 & ~x337 & ~x371 & ~x374 & ~x375 & ~x377 & ~x576 & ~x633 & ~x639 & ~x663 & ~x664 & ~x692 & ~x724;
assign c1412 =  x352 &  x437 & ~x91 & ~x144 & ~x145 & ~x156 & ~x202 & ~x257 & ~x315 & ~x367 & ~x425 & ~x510 & ~x666;
assign c1414 =  x485 & ~x30 & ~x44 & ~x125 & ~x196 & ~x223 & ~x252 & ~x280 & ~x338 & ~x364 & ~x418 & ~x509 & ~x536 & ~x544 & ~x571 & ~x599;
assign c1416 =  x732 & ~x545 & ~x564;
assign c1418 =  x356 & ~x25 & ~x45 & ~x124 & ~x226 & ~x477 & ~x496 & ~x499 & ~x502 & ~x654;
assign c1420 = ~x26 & ~x27 & ~x32 & ~x51 & ~x53 & ~x55 & ~x56 & ~x81 & ~x87 & ~x88 & ~x110 & ~x111 & ~x113 & ~x134 & ~x142 & ~x144 & ~x171 & ~x222 & ~x223 & ~x224 & ~x227 & ~x249 & ~x250 & ~x254 & ~x282 & ~x334 & ~x337 & ~x339 & ~x341 & ~x368 & ~x388 & ~x389 & ~x445 & ~x446 & ~x448 & ~x452 & ~x459 & ~x460 & ~x475 & ~x477 & ~x480 & ~x503 & ~x504 & ~x506 & ~x531 & ~x560 & ~x562 & ~x591 & ~x601 & ~x617 & ~x618 & ~x632 & ~x634 & ~x640 & ~x664 & ~x665 & ~x667 & ~x692 & ~x698 & ~x702 & ~x748 & ~x754 & ~x756 & ~x761 & ~x766;
assign c1422 =  x654 & ~x201 & ~x203 & ~x341 & ~x382 & ~x482 & ~x665 & ~x738;
assign c1424 =  x156 &  x298 & ~x81 & ~x226 & ~x253 & ~x283 & ~x419 & ~x452 & ~x478 & ~x585 & ~x605 & ~x643 & ~x664 & ~x673 & ~x693 & ~x696 & ~x725 & ~x749;
assign c1426 =  x733 & ~x87 & ~x153 & ~x339 & ~x477 & ~x506 & ~x564 & ~x591;
assign c1428 = ~x20 & ~x85 & ~x167 & ~x239 & ~x240 & ~x249 & ~x250 & ~x260 & ~x268 & ~x269 & ~x288 & ~x304 & ~x333 & ~x381 & ~x395 & ~x410 & ~x448 & ~x455 & ~x479 & ~x495 & ~x530 & ~x665 & ~x724 & ~x758 & ~x763;
assign c1430 =  x154 &  x296 & ~x52 & ~x108 & ~x112 & ~x114 & ~x164 & ~x166 & ~x193 & ~x195 & ~x198 & ~x249 & ~x334 & ~x360 & ~x364 & ~x368 & ~x395 & ~x446 & ~x450 & ~x506 & ~x574 & ~x603 & ~x604 & ~x645 & ~x671 & ~x695 & ~x696 & ~x697 & ~x722 & ~x723;
assign c1432 =  x211 &  x240 &  x353 & ~x91 & ~x165 & ~x398 & ~x423 & ~x605 & ~x722;
assign c1434 =  x324 &  x353 &  x381 &  x438 & ~x22 & ~x51 & ~x59 & ~x75 & ~x85 & ~x129 & ~x165 & ~x199 & ~x249 & ~x276 & ~x277 & ~x280 & ~x308 & ~x329 & ~x339 & ~x415 & ~x447 & ~x477 & ~x500 & ~x535 & ~x611 & ~x616 & ~x751 & ~x753;
assign c1436 =  x70 &  x296 & ~x25 & ~x32 & ~x60 & ~x109 & ~x169 & ~x192 & ~x253 & ~x304 & ~x306 & ~x399 & ~x416 & ~x423 & ~x426 & ~x428 & ~x430 & ~x431 & ~x449 & ~x588 & ~x640 & ~x645 & ~x667 & ~x735;
assign c1440 =  x651 & ~x84 & ~x137 & ~x226 & ~x254 & ~x309 & ~x363 & ~x391 & ~x474 & ~x475 & ~x502 & ~x533 & ~x536 & ~x562 & ~x563 & ~x565 & ~x573 & ~x588 & ~x590 & ~x592 & ~x618 & ~x646 & ~x657 & ~x673 & ~x674 & ~x685 & ~x713 & ~x754 & ~x756;
assign c1442 =  x371 &  x679;
assign c1444 =  x353 &  x523 & ~x53 & ~x102 & ~x111 & ~x113 & ~x144 & ~x161 & ~x170 & ~x192 & ~x226 & ~x246 & ~x276 & ~x277 & ~x309 & ~x311 & ~x333 & ~x390 & ~x392 & ~x424 & ~x445 & ~x447 & ~x449 & ~x476 & ~x564 & ~x615 & ~x668 & ~x696 & ~x697 & ~x698 & ~x699 & ~x723 & ~x728 & ~x730 & ~x749 & ~x755 & ~x782;
assign c1446 =  x273 &  x370 &  x401 & ~x363 & ~x445;
assign c1448 =  x129 &  x271 & ~x78 & ~x395 & ~x605 & ~x606;
assign c1450 = ~x0 & ~x2 & ~x24 & ~x31 & ~x51 & ~x58 & ~x78 & ~x112 & ~x132 & ~x144 & ~x161 & ~x162 & ~x222 & ~x254 & ~x278 & ~x282 & ~x283 & ~x309 & ~x362 & ~x446 & ~x508 & ~x510 & ~x511 & ~x515 & ~x516 & ~x517 & ~x518 & ~x535 & ~x536 & ~x630 & ~x646 & ~x659 & ~x660 & ~x671;
assign c1452 = ~x23 & ~x43 & ~x44 & ~x79 & ~x81 & ~x102 & ~x119 & ~x131 & ~x139 & ~x167 & ~x171 & ~x185 & ~x200 & ~x201 & ~x212 & ~x214 & ~x216 & ~x226 & ~x242 & ~x244 & ~x245 & ~x257 & ~x269 & ~x278 & ~x303 & ~x312 & ~x313 & ~x370 & ~x382 & ~x389 & ~x391 & ~x424 & ~x426 & ~x438 & ~x439 & ~x451 & ~x453 & ~x454 & ~x480 & ~x483 & ~x484 & ~x503 & ~x526 & ~x530 & ~x537 & ~x539 & ~x553 & ~x565 & ~x585 & ~x594 & ~x610 & ~x611 & ~x613 & ~x643 & ~x675 & ~x694 & ~x702;
assign c1454 = ~x0 & ~x1 & ~x3 & ~x4 & ~x16 & ~x20 & ~x22 & ~x23 & ~x24 & ~x25 & ~x27 & ~x30 & ~x44 & ~x51 & ~x52 & ~x53 & ~x55 & ~x57 & ~x59 & ~x60 & ~x71 & ~x80 & ~x81 & ~x85 & ~x86 & ~x109 & ~x110 & ~x113 & ~x114 & ~x136 & ~x137 & ~x138 & ~x165 & ~x167 & ~x168 & ~x192 & ~x193 & ~x196 & ~x213 & ~x220 & ~x221 & ~x224 & ~x225 & ~x226 & ~x248 & ~x250 & ~x251 & ~x252 & ~x254 & ~x261 & ~x275 & ~x277 & ~x279 & ~x280 & ~x281 & ~x304 & ~x307 & ~x308 & ~x309 & ~x332 & ~x333 & ~x334 & ~x336 & ~x360 & ~x361 & ~x363 & ~x364 & ~x365 & ~x366 & ~x389 & ~x390 & ~x391 & ~x392 & ~x412 & ~x413 & ~x414 & ~x415 & ~x416 & ~x417 & ~x418 & ~x419 & ~x420 & ~x422 & ~x423 & ~x424 & ~x425 & ~x439 & ~x440 & ~x441 & ~x442 & ~x444 & ~x445 & ~x446 & ~x447 & ~x449 & ~x450 & ~x451 & ~x452 & ~x469 & ~x470 & ~x471 & ~x473 & ~x474 & ~x475 & ~x477 & ~x478 & ~x479 & ~x482 & ~x502 & ~x503 & ~x504 & ~x505 & ~x506 & ~x532 & ~x533 & ~x534 & ~x559 & ~x587 & ~x588 & ~x615 & ~x616 & ~x643 & ~x647 & ~x671 & ~x698 & ~x699 & ~x721 & ~x723 & ~x724 & ~x725 & ~x726 & ~x727 & ~x749 & ~x750 & ~x751 & ~x752 & ~x754 & ~x755 & ~x756 & ~x774 & ~x775 & ~x777 & ~x778 & ~x779 & ~x781 & ~x783;
assign c1456 =  x381 & ~x226 & ~x389 & ~x395 & ~x420 & ~x432 & ~x434 & ~x449 & ~x454 & ~x605 & ~x641 & ~x664 & ~x665 & ~x725 & ~x726;
assign c1458 =  x408 & ~x14 & ~x49 & ~x81 & ~x93 & ~x120 & ~x196 & ~x278 & ~x313 & ~x314 & ~x390 & ~x519 & ~x547 & ~x589 & ~x594 & ~x696 & ~x781;
assign c1460 = ~x0 & ~x1 & ~x4 & ~x28 & ~x29 & ~x48 & ~x51 & ~x53 & ~x75 & ~x76 & ~x78 & ~x86 & ~x111 & ~x112 & ~x168 & ~x225 & ~x252 & ~x264 & ~x309 & ~x310 & ~x339 & ~x390 & ~x393 & ~x422 & ~x444 & ~x445 & ~x446 & ~x447 & ~x448 & ~x449 & ~x475 & ~x481 & ~x482 & ~x508 & ~x599 & ~x600 & ~x729 & ~x736 & ~x737 & ~x757 & ~x783;
assign c1462 =  x82;
assign c1464 = ~x0 & ~x3 & ~x26 & ~x47 & ~x87 & ~x106 & ~x114 & ~x115 & ~x135 & ~x139 & ~x145 & ~x160 & ~x164 & ~x170 & ~x173 & ~x194 & ~x197 & ~x199 & ~x200 & ~x224 & ~x225 & ~x229 & ~x251 & ~x255 & ~x314 & ~x334 & ~x337 & ~x338 & ~x339 & ~x341 & ~x342 & ~x343 & ~x364 & ~x367 & ~x369 & ~x374 & ~x387 & ~x400 & ~x401 & ~x403 & ~x415 & ~x418 & ~x420 & ~x423 & ~x430 & ~x432 & ~x433 & ~x434 & ~x449 & ~x451 & ~x533 & ~x558 & ~x585 & ~x588 & ~x641 & ~x643 & ~x647 & ~x668 & ~x671 & ~x676 & ~x728 & ~x753 & ~x762;
assign c1466 =  x126 &  x212 &  x268 &  x326 & ~x47 & ~x55 & ~x80 & ~x83 & ~x107 & ~x136 & ~x162 & ~x163 & ~x198 & ~x199 & ~x282 & ~x306 & ~x308 & ~x310 & ~x364 & ~x366 & ~x367 & ~x389 & ~x394 & ~x395 & ~x418 & ~x419 & ~x448 & ~x452 & ~x478 & ~x587 & ~x616 & ~x641 & ~x644 & ~x669 & ~x670 & ~x696 & ~x700 & ~x726 & ~x732 & ~x759 & ~x780 & ~x782;
assign c1468 = ~x25 & ~x54 & ~x56 & ~x69 & ~x97 & ~x223 & ~x224 & ~x225 & ~x363 & ~x447 & ~x450 & ~x480 & ~x507 & ~x535 & ~x545 & ~x563 & ~x572 & ~x573 & ~x589 & ~x600 & ~x629 & ~x658 & ~x686 & ~x709;
assign c1470 =  x377 &  x520 & ~x1 & ~x5 & ~x24 & ~x27 & ~x31 & ~x73 & ~x82 & ~x88 & ~x117 & ~x136 & ~x137 & ~x148 & ~x169 & ~x174 & ~x195 & ~x218 & ~x219 & ~x227 & ~x252 & ~x269 & ~x278 & ~x279 & ~x304 & ~x306 & ~x307 & ~x309 & ~x313 & ~x337 & ~x360 & ~x363 & ~x367 & ~x387 & ~x390 & ~x392 & ~x395 & ~x445 & ~x468 & ~x470 & ~x473 & ~x482 & ~x496 & ~x525 & ~x527 & ~x535 & ~x592 & ~x593 & ~x619 & ~x669 & ~x692 & ~x694 & ~x696 & ~x722 & ~x764;
assign c1472 =  x701;
assign c1474 = ~x16 & ~x18 & ~x44 & ~x83 & ~x97 & ~x125 & ~x208 & ~x390 & ~x406 & ~x415 & ~x433 & ~x449 & ~x544 & ~x653 & ~x764;
assign c1476 =  x294 & ~x25 & ~x87 & ~x102 & ~x119 & ~x136 & ~x147 & ~x171 & ~x182 & ~x183 & ~x184 & ~x230 & ~x277 & ~x387 & ~x414 & ~x452 & ~x479 & ~x526 & ~x618 & ~x667;
assign c1478 = ~x60 & ~x91 & ~x104 & ~x107 & ~x166 & ~x193 & ~x224 & ~x275 & ~x305 & ~x339 & ~x394 & ~x395 & ~x397 & ~x399 & ~x400 & ~x402 & ~x403 & ~x406 & ~x418 & ~x421 & ~x428 & ~x447 & ~x454 & ~x505 & ~x562 & ~x575 & ~x576 & ~x608 & ~x670 & ~x699 & ~x703 & ~x730 & ~x755 & ~x762 & ~x781;
assign c1480 =  x401 & ~x151 & ~x305 & ~x360 & ~x412 & ~x440 & ~x542 & ~x597;
assign c1482 =  x619 & ~x42 & ~x51 & ~x97 & ~x111 & ~x391 & ~x487 & ~x596 & ~x677;
assign c1484 = ~x0 & ~x3 & ~x24 & ~x28 & ~x51 & ~x53 & ~x58 & ~x59 & ~x79 & ~x83 & ~x84 & ~x108 & ~x109 & ~x111 & ~x135 & ~x136 & ~x140 & ~x141 & ~x142 & ~x164 & ~x167 & ~x169 & ~x191 & ~x193 & ~x194 & ~x195 & ~x196 & ~x198 & ~x221 & ~x222 & ~x226 & ~x247 & ~x248 & ~x249 & ~x251 & ~x252 & ~x276 & ~x277 & ~x278 & ~x279 & ~x280 & ~x281 & ~x304 & ~x305 & ~x307 & ~x309 & ~x333 & ~x336 & ~x362 & ~x363 & ~x364 & ~x366 & ~x389 & ~x392 & ~x394 & ~x418 & ~x419 & ~x420 & ~x421 & ~x422 & ~x446 & ~x447 & ~x448 & ~x449 & ~x450 & ~x477 & ~x478 & ~x479 & ~x506 & ~x512 & ~x513 & ~x514 & ~x515 & ~x516 & ~x517 & ~x534 & ~x630 & ~x631 & ~x643 & ~x660 & ~x661 & ~x666 & ~x667 & ~x669 & ~x693 & ~x694 & ~x695 & ~x696 & ~x697 & ~x722 & ~x723 & ~x724 & ~x751 & ~x752 & ~x753 & ~x757 & ~x761 & ~x781 & ~x783;
assign c1486 =  x439 & ~x5 & ~x24 & ~x26 & ~x28 & ~x29 & ~x51 & ~x77 & ~x81 & ~x83 & ~x87 & ~x104 & ~x105 & ~x113 & ~x172 & ~x189 & ~x195 & ~x199 & ~x249 & ~x253 & ~x278 & ~x280 & ~x286 & ~x307 & ~x312 & ~x314 & ~x336 & ~x337 & ~x342 & ~x361 & ~x368 & ~x387 & ~x418 & ~x423 & ~x445 & ~x448 & ~x451 & ~x452 & ~x472 & ~x475 & ~x478 & ~x480 & ~x501 & ~x559 & ~x585 & ~x588 & ~x590 & ~x615 & ~x644 & ~x645 & ~x647 & ~x670 & ~x672 & ~x674 & ~x698 & ~x699 & ~x719 & ~x728 & ~x752 & ~x775 & ~x781;
assign c1488 = ~x48 & ~x106 & ~x144 & ~x167 & ~x199 & ~x335 & ~x398 & ~x426 & ~x427 & ~x429 & ~x430 & ~x431 & ~x455 & ~x456 & ~x475 & ~x534 & ~x562 & ~x587 & ~x589 & ~x602 & ~x617 & ~x631 & ~x632 & ~x633 & ~x634 & ~x663 & ~x694 & ~x695 & ~x701 & ~x722 & ~x755 & ~x783;
assign c1490 =  x66 & ~x2 & ~x12 & ~x23 & ~x75 & ~x77 & ~x79 & ~x106 & ~x119 & ~x120 & ~x134 & ~x137 & ~x146 & ~x147 & ~x164 & ~x168 & ~x169 & ~x192 & ~x198 & ~x222 & ~x229 & ~x230 & ~x251 & ~x285 & ~x310 & ~x311 & ~x363 & ~x365 & ~x368 & ~x369 & ~x390 & ~x392 & ~x423 & ~x445 & ~x449 & ~x506 & ~x511 & ~x536 & ~x557 & ~x561 & ~x562 & ~x586 & ~x618 & ~x644 & ~x645 & ~x675 & ~x725 & ~x752 & ~x758 & ~x778 & ~x779;
assign c1492 =  x35 & ~x30 & ~x85 & ~x87 & ~x170 & ~x225 & ~x309 & ~x337 & ~x478 & ~x505 & ~x560 & ~x561 & ~x575 & ~x590;
assign c1494 =  x299 & ~x3 & ~x18 & ~x20 & ~x25 & ~x28 & ~x46 & ~x49 & ~x51 & ~x55 & ~x80 & ~x86 & ~x96 & ~x108 & ~x137 & ~x138 & ~x139 & ~x168 & ~x193 & ~x194 & ~x223 & ~x225 & ~x250 & ~x251 & ~x275 & ~x276 & ~x277 & ~x304 & ~x305 & ~x306 & ~x307 & ~x308 & ~x310 & ~x332 & ~x334 & ~x336 & ~x363 & ~x390 & ~x420 & ~x444 & ~x448 & ~x449 & ~x451 & ~x476 & ~x479 & ~x502 & ~x506 & ~x507 & ~x531 & ~x532 & ~x560 & ~x587 & ~x588 & ~x589 & ~x615 & ~x616 & ~x698 & ~x764 & ~x765 & ~x782 & ~x783;
assign c1496 =  x320 & ~x12 & ~x16 & ~x20 & ~x52 & ~x82 & ~x223 & ~x262 & ~x389 & ~x404 & ~x418 & ~x419 & ~x432 & ~x447 & ~x532;
assign c1498 =  x757;
assign c11 =  x390;
assign c13 =  x240 &  x405 & ~x316 & ~x358 & ~x477 & ~x503 & ~x559 & ~x587;
assign c15 = ~x26 & ~x59 & ~x167 & ~x243 & ~x247 & ~x357 & ~x384 & ~x441 & ~x445 & ~x468 & ~x631 & ~x655 & ~x656 & ~x658 & ~x684 & ~x759;
assign c17 =  x520 &  x547 &  x602 & ~x0 & ~x20 & ~x30 & ~x50 & ~x83 & ~x140 & ~x169 & ~x194 & ~x280 & ~x336 & ~x364 & ~x394 & ~x419 & ~x420 & ~x449 & ~x506 & ~x532 & ~x561 & ~x614 & ~x616 & ~x669 & ~x671 & ~x672 & ~x700 & ~x725 & ~x731 & ~x753 & ~x754 & ~x761 & ~x780;
assign c19 =  x547 &  x602 &  x656 & ~x53 & ~x197 & ~x448 & ~x503 & ~x504 & ~x563 & ~x588 & ~x589 & ~x671 & ~x727;
assign c111 =  x183 &  x267 & ~x68 & ~x559 & ~x587 & ~x615 & ~x623 & ~x778;
assign c113 =  x517 & ~x272 & ~x299 & ~x520;
assign c115 =  x96 & ~x0 & ~x2 & ~x4 & ~x6 & ~x25 & ~x29 & ~x30 & ~x53 & ~x55 & ~x112 & ~x113 & ~x141 & ~x168 & ~x169 & ~x195 & ~x225 & ~x249 & ~x280 & ~x351 & ~x359 & ~x360 & ~x389 & ~x419 & ~x441 & ~x444 & ~x448 & ~x471 & ~x472 & ~x499 & ~x501 & ~x502 & ~x531 & ~x782 & ~x783;
assign c117 =  x323 &  x435 &  x463 & ~x68 & ~x124 & ~x674 & ~x731;
assign c119 =  x485 & ~x551 & ~x606 & ~x659 & ~x660 & ~x756;
assign c121 =  x399 &  x623 & ~x404 & ~x406 & ~x431 & ~x459;
assign c123 = ~x19 & ~x54 & ~x71 & ~x109 & ~x266 & ~x478 & ~x495 & ~x550 & ~x633 & ~x660 & ~x782;
assign c125 =  x611 & ~x580 & ~x609;
assign c127 =  x312 & ~x371 & ~x398 & ~x399 & ~x454;
assign c129 =  x257 & ~x0 & ~x110 & ~x336 & ~x343 & ~x399 & ~x779;
assign c131 = ~x0 & ~x1 & ~x2 & ~x3 & ~x5 & ~x19 & ~x25 & ~x27 & ~x29 & ~x30 & ~x31 & ~x32 & ~x34 & ~x35 & ~x40 & ~x54 & ~x57 & ~x58 & ~x86 & ~x87 & ~x96 & ~x111 & ~x113 & ~x117 & ~x118 & ~x140 & ~x141 & ~x142 & ~x169 & ~x170 & ~x195 & ~x224 & ~x225 & ~x250 & ~x251 & ~x253 & ~x279 & ~x282 & ~x308 & ~x336 & ~x379 & ~x683 & ~x727 & ~x737 & ~x756 & ~x764 & ~x780 & ~x783;
assign c133 = ~x69 & ~x84 & ~x447 & ~x485 & ~x527 & ~x569 & ~x584 & ~x644 & ~x673 & ~x700 & ~x728 & ~x731 & ~x757 & ~x766 & ~x767 & ~x783;
assign c135 =  x170;
assign c137 =  x460 & ~x24 & ~x257 & ~x308 & ~x364 & ~x476 & ~x577 & ~x630 & ~x732;
assign c139 =  x390;
assign c141 =  x416 & ~x440;
assign c143 = ~x213 & ~x339 & ~x340 & ~x439 & ~x466 & ~x521 & ~x666 & ~x704 & ~x755;
assign c145 =  x659 &  x686 &  x713 &  x739 & ~x1 & ~x3 & ~x225 & ~x532 & ~x642 & ~x729 & ~x755 & ~x758;
assign c147 =  x462 &  x488 &  x541 & ~x54 & ~x56 & ~x756 & ~x781;
assign c149 =  x515 &  x571 &  x739 & ~x22 & ~x364;
assign c151 = ~x83 & ~x411 & ~x436 & ~x465 & ~x492 & ~x494 & ~x549 & ~x603 & ~x773;
assign c153 = ~x24 & ~x30 & ~x39 & ~x158 & ~x428 & ~x526 & ~x565 & ~x594 & ~x674 & ~x679 & ~x764 & ~x771;
assign c155 = ~x8 & ~x12 & ~x34 & ~x37 & ~x39 & ~x55 & ~x65 & ~x87 & ~x111 & ~x114 & ~x139 & ~x140 & ~x419 & ~x617 & ~x647 & ~x654 & ~x673 & ~x682 & ~x697 & ~x701 & ~x730 & ~x738 & ~x739 & ~x753 & ~x765 & ~x783;
assign c157 =  x533;
assign c159 = ~x27 & ~x105 & ~x134 & ~x186 & ~x452 & ~x467 & ~x493 & ~x496 & ~x548 & ~x774;
assign c161 =  x291 &  x319 & ~x27 & ~x80 & ~x204 & ~x205 & ~x259 & ~x284 & ~x501;
assign c163 =  x367 & ~x400 & ~x401;
assign c165 =  x348 & ~x109 & ~x630 & ~x655 & ~x657;
assign c167 =  x490 &  x517 &  x545 & ~x83 & ~x254 & ~x300 & ~x442 & ~x783;
assign c169 =  x508 & ~x1 & ~x26 & ~x31 & ~x58 & ~x89 & ~x116 & ~x304 & ~x547 & ~x574 & ~x601 & ~x602;
assign c171 =  x741 & ~x0 & ~x390 & ~x422 & ~x450 & ~x479 & ~x502 & ~x523 & ~x605 & ~x645 & ~x728;
assign c173 =  x183 &  x211 &  x267 & ~x243 & ~x467 & ~x701;
assign c175 = ~x22 & ~x26 & ~x29 & ~x30 & ~x49 & ~x50 & ~x52 & ~x56 & ~x78 & ~x83 & ~x86 & ~x106 & ~x109 & ~x111 & ~x112 & ~x134 & ~x135 & ~x136 & ~x139 & ~x164 & ~x191 & ~x192 & ~x194 & ~x218 & ~x224 & ~x248 & ~x251 & ~x278 & ~x279 & ~x306 & ~x335 & ~x336 & ~x360 & ~x387 & ~x414 & ~x415 & ~x437 & ~x444 & ~x446 & ~x464 & ~x493 & ~x502 & ~x548 & ~x560 & ~x756 & ~x758;
assign c177 =  x397 & ~x56 & ~x60 & ~x82 & ~x86 & ~x87 & ~x110 & ~x111 & ~x114 & ~x142 & ~x166 & ~x167 & ~x198 & ~x199 & ~x224 & ~x225 & ~x253 & ~x281 & ~x283 & ~x311 & ~x376 & ~x559 & ~x589 & ~x671 & ~x672 & ~x700 & ~x755;
assign c179 =  x545 & ~x1 & ~x2 & ~x66 & ~x109 & ~x195 & ~x355 & ~x383 & ~x419 & ~x757 & ~x782;
assign c181 =  x42 &  x155 &  x239 &  x351;
assign c183 =  x459 &  x543 & ~x2 & ~x36 & ~x90 & ~x112 & ~x136 & ~x145 & ~x168 & ~x419 & ~x449 & ~x783;
assign c185 = ~x84 & ~x110 & ~x111 & ~x112 & ~x225 & ~x274 & ~x281 & ~x303 & ~x332 & ~x335 & ~x363 & ~x445 & ~x447 & ~x531 & ~x557 & ~x558 & ~x633 & ~x662 & ~x688 & ~x689 & ~x709 & ~x713 & ~x714 & ~x716 & ~x737 & ~x740 & ~x742 & ~x755 & ~x756 & ~x778;
assign c187 = ~x110 & ~x419 & ~x447 & ~x487 & ~x503 & ~x530 & ~x542 & ~x565 & ~x571 & ~x572 & ~x584 & ~x617 & ~x620 & ~x626 & ~x651 & ~x678 & ~x680 & ~x699 & ~x700 & ~x728 & ~x755 & ~x765;
assign c189 =  x575 &  x630 & ~x660 & ~x779;
assign c191 =  x75 & ~x22 & ~x317 & ~x682;
assign c193 =  x662 & ~x68 & ~x168 & ~x556 & ~x665 & ~x751;
assign c195 = ~x327 & ~x380 & ~x381 & ~x383 & ~x408 & ~x409 & ~x435 & ~x638 & ~x671 & ~x704;
assign c197 =  x179 & ~x4 & ~x141 & ~x377 & ~x404 & ~x405 & ~x459;
assign c199 = ~x27 & ~x82 & ~x137 & ~x309 & ~x447 & ~x526 & ~x572 & ~x581 & ~x598 & ~x642 & ~x645 & ~x647 & ~x669 & ~x705 & ~x712 & ~x739 & ~x761 & ~x764;
assign c1101 =  x632 &  x659 &  x685 & ~x25 & ~x196 & ~x508 & ~x561 & ~x562 & ~x563 & ~x590 & ~x618 & ~x696 & ~x697 & ~x702 & ~x754 & ~x781;
assign c1103 = ~x21 & ~x50 & ~x51 & ~x85 & ~x336 & ~x351 & ~x420 & ~x492 & ~x547 & ~x574 & ~x598 & ~x602 & ~x626 & ~x654 & ~x759 & ~x760;
assign c1105 =  x203 & ~x345 & ~x346 & ~x372 & ~x373 & ~x450 & ~x455 & ~x533 & ~x587 & ~x617 & ~x644 & ~x672 & ~x754 & ~x757 & ~x760;
assign c1107 =  x524 &  x610 & ~x278 & ~x332 & ~x529 & ~x739;
assign c1109 =  x411 &  x439 &  x467 & ~x276 & ~x659 & ~x713 & ~x741;
assign c1111 =  x401 & ~x9 & ~x36 & ~x494 & ~x578 & ~x605;
assign c1113 =  x488 & ~x185 & ~x576 & ~x760;
assign c1115 =  x423 & ~x27 & ~x30 & ~x87 & ~x170 & ~x197 & ~x223 & ~x274 & ~x757;
assign c1117 = ~x3 & ~x25 & ~x110 & ~x394 & ~x466 & ~x493 & ~x521 & ~x533 & ~x615 & ~x760;
assign c1119 =  x166;
assign c1121 =  x349 &  x405 &  x460 & ~x259 & ~x577;
assign c1123 =  x632 &  x659 &  x686 & ~x56 & ~x140 & ~x422 & ~x450 & ~x477 & ~x479 & ~x535 & ~x565 & ~x589 & ~x590 & ~x616 & ~x619 & ~x644 & ~x675 & ~x703;
assign c1125 = ~x242 & ~x284 & ~x370 & ~x495 & ~x521 & ~x522 & ~x548 & ~x638 & ~x648 & ~x760;
assign c1127 = ~x10 & ~x124 & ~x483 & ~x623 & ~x681 & ~x709;
assign c1129 = ~x126 & ~x154 & ~x192 & ~x250 & ~x392 & ~x493 & ~x521 & ~x578 & ~x603 & ~x630;
assign c1131 =  x603 &  x658 &  x684 & ~x0 & ~x21 & ~x23 & ~x30 & ~x50 & ~x53 & ~x56 & ~x59 & ~x84 & ~x112 & ~x192 & ~x197 & ~x224 & ~x421 & ~x508 & ~x697 & ~x699 & ~x724 & ~x727;
assign c1133 =  x231 & ~x319 & ~x400 & ~x428 & ~x624 & ~x680;
assign c1135 =  x491 &  x517 &  x544 &  x571 & ~x216 & ~x280;
assign c1137 =  x154 &  x210 &  x238 & ~x25 & ~x27 & ~x30 & ~x32 & ~x83 & ~x110 & ~x114 & ~x138 & ~x223 & ~x279 & ~x380 & ~x447 & ~x502 & ~x504 & ~x728;
assign c1139 =  x536 & ~x26 & ~x69 & ~x82 & ~x113 & ~x115 & ~x143 & ~x144 & ~x172 & ~x252 & ~x282 & ~x502 & ~x701;
assign c1141 =  x150 & ~x8 & ~x23 & ~x389 & ~x390 & ~x405 & ~x415 & ~x470 & ~x499 & ~x542 & ~x760;
assign c1143 =  x164 & ~x247 & ~x303 & ~x392;
assign c1145 = ~x24 & ~x84 & ~x87 & ~x90 & ~x115 & ~x142 & ~x145 & ~x173 & ~x331 & ~x392 & ~x421 & ~x474 & ~x515 & ~x529 & ~x542 & ~x571 & ~x599 & ~x612 & ~x615 & ~x627 & ~x653 & ~x710 & ~x736 & ~x756 & ~x764;
assign c1147 =  x398 &  x426 &  x482 &  x510 & ~x283 & ~x284 & ~x340 & ~x367 & ~x392 & ~x420 & ~x671 & ~x759;
assign c1149 =  x155 &  x267 & ~x30 & ~x275 & ~x470 & ~x495 & ~x496;
assign c1151 = ~x2 & ~x31 & ~x81 & ~x85 & ~x140 & ~x392 & ~x475 & ~x503 & ~x515 & ~x527 & ~x543 & ~x569 & ~x571 & ~x588 & ~x596 & ~x597 & ~x618 & ~x625 & ~x643 & ~x644 & ~x646 & ~x653 & ~x675 & ~x682 & ~x697 & ~x698 & ~x699 & ~x708 & ~x727 & ~x728 & ~x737 & ~x755 & ~x764;
assign c1153 =  x490 & ~x404 & ~x614;
assign c1155 =  x293 &  x370 & ~x272 & ~x301;
assign c1157 =  x738 & ~x85 & ~x552 & ~x578 & ~x579 & ~x605;
assign c1159 =  x129 & ~x4 & ~x60 & ~x281 & ~x310 & ~x332 & ~x359 & ~x414 & ~x472 & ~x501 & ~x528 & ~x531 & ~x555 & ~x597 & ~x728 & ~x729;
assign c1161 = ~x1 & ~x2 & ~x3 & ~x27 & ~x28 & ~x29 & ~x55 & ~x56 & ~x57 & ~x58 & ~x59 & ~x83 & ~x85 & ~x86 & ~x89 & ~x104 & ~x106 & ~x111 & ~x113 & ~x114 & ~x115 & ~x140 & ~x141 & ~x142 & ~x143 & ~x161 & ~x168 & ~x169 & ~x170 & ~x171 & ~x174 & ~x189 & ~x196 & ~x197 & ~x217 & ~x218 & ~x219 & ~x220 & ~x224 & ~x227 & ~x228 & ~x245 & ~x246 & ~x247 & ~x248 & ~x249 & ~x252 & ~x273 & ~x274 & ~x275 & ~x280 & ~x304 & ~x306 & ~x309 & ~x333 & ~x362 & ~x366 & ~x393 & ~x414 & ~x417 & ~x418 & ~x420 & ~x444 & ~x473 & ~x475 & ~x575 & ~x603 & ~x629 & ~x630 & ~x643 & ~x656 & ~x657 & ~x671 & ~x756 & ~x759 & ~x783;
assign c1163 =  x458 & ~x58 & ~x82 & ~x551 & ~x578 & ~x579 & ~x605 & ~x659 & ~x755;
assign c1165 =  x574 & ~x18 & ~x394 & ~x414 & ~x478 & ~x513 & ~x671;
assign c1167 = ~x3 & ~x27 & ~x86 & ~x115 & ~x141 & ~x274 & ~x334 & ~x432 & ~x445 & ~x448 & ~x472 & ~x473 & ~x487 & ~x526 & ~x529 & ~x532 & ~x541 & ~x543 & ~x625 & ~x651 & ~x680 & ~x756;
assign c1169 =  x554 &  x582 & ~x323 & ~x408;
assign c1171 =  x519 &  x546 &  x572 &  x573 & ~x87 & ~x537 & ~x560;
assign c1173 = ~x32 & ~x112 & ~x141 & ~x169 & ~x251 & ~x513 & ~x543 & ~x562 & ~x568 & ~x571 & ~x591 & ~x596 & ~x625 & ~x643 & ~x653 & ~x681 & ~x695 & ~x736 & ~x766 & ~x767 & ~x780;
assign c1175 =  x314 & ~x215 & ~x224 & ~x272 & ~x277 & ~x305 & ~x755 & ~x772 & ~x782;
assign c1177 =  x313 & ~x30 & ~x82 & ~x141 & ~x188 & ~x226 & ~x421 & ~x475 & ~x531 & ~x557 & ~x561 & ~x587 & ~x613 & ~x614 & ~x616 & ~x670 & ~x672 & ~x777;
assign c1179 = ~x1 & ~x3 & ~x4 & ~x5 & ~x29 & ~x32 & ~x52 & ~x57 & ~x82 & ~x136 & ~x279 & ~x336 & ~x382 & ~x392 & ~x408 & ~x410 & ~x437 & ~x438 & ~x464 & ~x466 & ~x494 & ~x520 & ~x522 & ~x547 & ~x550 & ~x576 & ~x757 & ~x783;
assign c1181 = ~x82 & ~x128 & ~x135 & ~x138 & ~x225 & ~x364 & ~x394 & ~x450 & ~x466 & ~x521 & ~x522 & ~x576 & ~x631 & ~x669 & ~x731;
assign c1183 =  x468 &  x496 &  x552 & ~x277 & ~x305 & ~x332 & ~x336 & ~x473 & ~x500 & ~x772 & ~x778;
assign c1185 = ~x2 & ~x22 & ~x45 & ~x84 & ~x110 & ~x112 & ~x140 & ~x166 & ~x168 & ~x224 & ~x270 & ~x271 & ~x297 & ~x523 & ~x577 & ~x604 & ~x605 & ~x631;
assign c1187 = ~x15 & ~x53 & ~x57 & ~x76 & ~x80 & ~x134 & ~x145 & ~x223 & ~x226 & ~x246 & ~x324 & ~x587 & ~x604 & ~x674 & ~x679 & ~x698 & ~x727 & ~x731 & ~x778 & ~x782;
assign c1189 = ~x8 & ~x11 & ~x13 & ~x14 & ~x19 & ~x26 & ~x609 & ~x645 & ~x672 & ~x676 & ~x702 & ~x705 & ~x732 & ~x733 & ~x735 & ~x740 & ~x751 & ~x753 & ~x754 & ~x762 & ~x769 & ~x773 & ~x774;
assign c1191 = ~x0 & ~x1 & ~x2 & ~x29 & ~x83 & ~x96 & ~x123 & ~x151 & ~x364 & ~x410 & ~x438 & ~x448 & ~x466 & ~x521 & ~x522 & ~x549 & ~x577 & ~x605 & ~x634 & ~x671 & ~x728 & ~x756 & ~x783;
assign c1193 =  x228 & ~x2 & ~x86 & ~x343 & ~x364 & ~x371 & ~x699 & ~x755;
assign c1195 =  x276 & ~x612 & ~x616 & ~x648 & ~x676 & ~x677;
assign c1197 =  x254 & ~x757 & ~x778;
assign c1199 = ~x4 & ~x19 & ~x48 & ~x85 & ~x90 & ~x146 & ~x168 & ~x170 & ~x267 & ~x323 & ~x405 & ~x406 & ~x444 & ~x669;
assign c1201 =  x606 &  x633 &  x634 &  x661 &  x688 & ~x84 & ~x110 & ~x140 & ~x645 & ~x672;
assign c1203 =  x509 & ~x0 & ~x4 & ~x23 & ~x29 & ~x56 & ~x58 & ~x59 & ~x82 & ~x84 & ~x86 & ~x87 & ~x336 & ~x503 & ~x529 & ~x614 & ~x615 & ~x671 & ~x672 & ~x699 & ~x701 & ~x727 & ~x738 & ~x739 & ~x766 & ~x781;
assign c1205 =  x533;
assign c1207 = ~x17 & ~x50 & ~x84 & ~x87 & ~x112 & ~x114 & ~x116 & ~x138 & ~x218 & ~x247 & ~x248 & ~x252 & ~x305 & ~x306 & ~x333 & ~x386 & ~x414 & ~x415 & ~x436 & ~x464 & ~x490 & ~x498 & ~x547 & ~x574 & ~x758;
assign c1209 =  x446;
assign c1211 =  x208 &  x402 &  x485 & ~x84 & ~x417 & ~x560;
assign c1213 = ~x23 & ~x28 & ~x32 & ~x51 & ~x54 & ~x80 & ~x135 & ~x163 & ~x504 & ~x521 & ~x548 & ~x560 & ~x644 & ~x706 & ~x735;
assign c1215 =  x166;
assign c1217 =  x371 &  x427 &  x455 & ~x5 & ~x85 & ~x640 & ~x697 & ~x704 & ~x725 & ~x733 & ~x758;
assign c1219 = ~x9 & ~x84 & ~x87 & ~x139 & ~x167 & ~x416 & ~x551 & ~x552 & ~x560 & ~x577 & ~x604 & ~x606 & ~x615 & ~x632 & ~x633 & ~x659 & ~x661 & ~x687;
assign c1221 =  x259 &  x287 & ~x690 & ~x701 & ~x718 & ~x730 & ~x747 & ~x756 & ~x773;
assign c1223 = ~x20 & ~x243 & ~x495 & ~x521 & ~x528 & ~x540 & ~x550 & ~x576 & ~x595 & ~x642;
assign c1225 =  x194;
assign c1227 =  x238 &  x294 & ~x9 & ~x36 & ~x497;
assign c1229 = ~x1 & ~x2 & ~x3 & ~x26 & ~x31 & ~x35 & ~x58 & ~x83 & ~x88 & ~x89 & ~x114 & ~x117 & ~x141 & ~x142 & ~x191 & ~x304 & ~x330 & ~x602 & ~x630 & ~x656 & ~x657 & ~x682 & ~x683 & ~x684 & ~x690 & ~x718 & ~x737;
assign c1231 =  x258 & ~x2 & ~x24 & ~x53 & ~x54 & ~x84 & ~x85 & ~x87 & ~x111 & ~x137 & ~x139 & ~x196 & ~x224 & ~x373 & ~x391 & ~x401 & ~x417 & ~x420 & ~x428 & ~x445 & ~x455 & ~x456 & ~x473 & ~x474 & ~x483 & ~x484 & ~x503 & ~x505 & ~x511 & ~x531 & ~x533 & ~x560 & ~x561 & ~x588 & ~x589 & ~x616 & ~x644 & ~x672 & ~x673 & ~x698 & ~x700 & ~x701 & ~x756 & ~x758 & ~x783;
assign c1233 = ~x162 & ~x168 & ~x284 & ~x469 & ~x473 & ~x501 & ~x522 & ~x529 & ~x548 & ~x658;
assign c1235 = ~x1 & ~x3 & ~x4 & ~x160 & ~x166 & ~x415 & ~x420 & ~x438 & ~x465 & ~x467 & ~x495 & ~x548 & ~x702 & ~x763;
assign c1237 =  x361 & ~x643 & ~x696;
assign c1239 =  x745 & ~x29 & ~x133 & ~x190 & ~x558 & ~x617 & ~x641 & ~x643 & ~x686;
assign c1241 =  x401 &  x456 &  x484 & ~x0 & ~x32 & ~x170 & ~x171 & ~x244 & ~x304 & ~x336 & ~x761;
assign c1243 =  x540 &  x708 &  x736;
assign c1245 =  x509 &  x621 & ~x284;
assign c1247 =  x435 & ~x27 & ~x346 & ~x402 & ~x455 & ~x589 & ~x761;
assign c1249 =  x128 &  x156 &  x212 &  x240 & ~x59 & ~x168 & ~x270 & ~x781 & ~x783;
assign c1251 = ~x18 & ~x31 & ~x320 & ~x363 & ~x454 & ~x482 & ~x509 & ~x510 & ~x527 & ~x533 & ~x536 & ~x539 & ~x559 & ~x561 & ~x567 & ~x593 & ~x617 & ~x620 & ~x623 & ~x641 & ~x642 & ~x645 & ~x648 & ~x650 & ~x651 & ~x677 & ~x706 & ~x707 & ~x713 & ~x756;
assign c1253 =  x239 &  x267 &  x406 &  x434 &  x490 & ~x29 & ~x31 & ~x56 & ~x614;
assign c1255 =  x506 & ~x249 & ~x280 & ~x336;
assign c1257 =  x96 & ~x139 & ~x238 & ~x294 & ~x322 & ~x336 & ~x419 & ~x585 & ~x706;
assign c1259 =  x148 & ~x24 & ~x55 & ~x57 & ~x140 & ~x168 & ~x502 & ~x504 & ~x506 & ~x507 & ~x509 & ~x510 & ~x532 & ~x533 & ~x538 & ~x562 & ~x566 & ~x588 & ~x589 & ~x592 & ~x594 & ~x614 & ~x617 & ~x619 & ~x620 & ~x621 & ~x622 & ~x623 & ~x645 & ~x647 & ~x649 & ~x650 & ~x651 & ~x675 & ~x676 & ~x677 & ~x678 & ~x679 & ~x698 & ~x701 & ~x702 & ~x705 & ~x707 & ~x726 & ~x732 & ~x735 & ~x760 & ~x761 & ~x763 & ~x780;
assign c1261 =  x406 &  x434 & ~x187 & ~x215 & ~x549;
assign c1263 =  x331 & ~x392 & ~x440;
assign c1265 = ~x266 & ~x595 & ~x618 & ~x650 & ~x674 & ~x680 & ~x712 & ~x728 & ~x730 & ~x737 & ~x780;
assign c1267 =  x605 &  x631 &  x658 & ~x25 & ~x55 & ~x57 & ~x110 & ~x139 & ~x223 & ~x251 & ~x536 & ~x560 & ~x588 & ~x616 & ~x642 & ~x643 & ~x672 & ~x756 & ~x758 & ~x783;
assign c1269 =  x417 &  x445;
assign c1271 =  x185 &  x213 &  x241 & ~x2 & ~x3 & ~x70 & ~x82 & ~x97 & ~x114 & ~x392 & ~x419 & ~x447 & ~x471 & ~x472 & ~x501 & ~x528 & ~x530 & ~x559 & ~x615;
assign c1273 =  x382 & ~x5 & ~x25 & ~x29 & ~x32 & ~x54 & ~x56 & ~x83 & ~x86 & ~x197 & ~x530 & ~x541 & ~x557 & ~x569 & ~x626 & ~x643 & ~x654 & ~x709 & ~x765;
assign c1275 =  x202 & ~x343 & ~x371 & ~x421 & ~x556 & ~x671 & ~x673 & ~x730 & ~x753 & ~x754 & ~x778;
assign c1277 =  x234 &  x289 & ~x169 & ~x405 & ~x460 & ~x725;
assign c1279 =  x378 & ~x68 & ~x208 & ~x345 & ~x624 & ~x644;
assign c1281 =  x268 & ~x64 & ~x69 & ~x70 & ~x97 & ~x196 & ~x500 & ~x559 & ~x584 & ~x587 & ~x615 & ~x645 & ~x731 & ~x757 & ~x760;
assign c1283 =  x517 &  x544 &  x572 & ~x23 & ~x281 & ~x356 & ~x533;
assign c1285 =  x535 & ~x31 & ~x87 & ~x301 & ~x329 & ~x615;
assign c1287 =  x322 &  x377 & ~x285 & ~x370 & ~x371 & ~x495 & ~x522;
assign c1289 =  x162 & ~x417 & ~x528 & ~x529 & ~x555 & ~x584 & ~x701 & ~x754 & ~x760;
assign c1291 = ~x4 & ~x12 & ~x36 & ~x39 & ~x56 & ~x66 & ~x93 & ~x104 & ~x329 & ~x331 & ~x364 & ~x391 & ~x445 & ~x471 & ~x472 & ~x501 & ~x515 & ~x527 & ~x530 & ~x556 & ~x728;
assign c1293 = ~x4 & ~x197 & ~x221 & ~x246 & ~x274 & ~x303 & ~x330 & ~x351 & ~x379 & ~x435 & ~x462 & ~x626 & ~x689;
assign c1295 =  x466 &  x494 &  x549 & ~x84 & ~x274 & ~x336 & ~x359 & ~x531 & ~x587 & ~x672 & ~x769 & ~x770;
assign c1297 =  x445;
assign c1299 =  x459 &  x515 & ~x366 & ~x450 & ~x531;
assign c1301 = ~x10 & ~x12 & ~x24 & ~x28 & ~x41 & ~x67 & ~x106 & ~x164 & ~x264 & ~x413 & ~x469 & ~x558 & ~x585 & ~x613 & ~x615 & ~x670;
assign c1303 =  x154 &  x182 & ~x32 & ~x84 & ~x104 & ~x195 & ~x325 & ~x352 & ~x783;
assign c1305 =  x100 & ~x469 & ~x551;
assign c1307 = ~x21 & ~x122 & ~x123 & ~x151 & ~x337 & ~x392 & ~x440 & ~x467 & ~x468 & ~x497 & ~x524 & ~x531 & ~x551 & ~x558 & ~x612 & ~x643 & ~x667 & ~x705 & ~x722 & ~x733 & ~x753 & ~x762 & ~x763;
assign c1309 =  x547 &  x573 & ~x114 & ~x144 & ~x394 & ~x405 & ~x432 & ~x541;
assign c1311 =  x463 &  x490 & ~x54 & ~x169 & ~x227 & ~x364 & ~x449 & ~x561 & ~x616 & ~x639;
assign c1313 =  x367 & ~x83 & ~x112 & ~x225 & ~x454 & ~x783;
assign c1315 =  x150 &  x178 &  x261 & ~x2 & ~x44 & ~x100 & ~x476 & ~x477 & ~x732;
assign c1317 =  x440 &  x582 & ~x276 & ~x743;
assign c1319 = ~x80 & ~x134 & ~x163 & ~x165 & ~x191 & ~x192 & ~x248 & ~x249 & ~x305 & ~x336 & ~x488 & ~x492 & ~x548 & ~x576 & ~x603 & ~x630 & ~x658 & ~x760 & ~x778;
assign c1321 =  x305 & ~x552 & ~x581 & ~x694 & ~x698 & ~x724 & ~x755;
assign c1323 =  x515 & ~x18 & ~x240 & ~x548 & ~x647;
assign c1325 =  x507 & ~x221 & ~x250 & ~x547;
assign c1327 =  x150 & ~x56 & ~x139 & ~x265 & ~x294 & ~x703 & ~x729;
assign c1329 = ~x8 & ~x12 & ~x38 & ~x40 & ~x65 & ~x111 & ~x167 & ~x171 & ~x226 & ~x417 & ~x471 & ~x472 & ~x498 & ~x526 & ~x528;
assign c1331 =  x377 & ~x308 & ~x616 & ~x655 & ~x705 & ~x783;
assign c1333 = ~x27 & ~x140 & ~x208 & ~x424 & ~x467 & ~x550 & ~x578 & ~x605 & ~x634 & ~x648 & ~x661 & ~x732;
assign c1335 =  x179 & ~x323 & ~x351 & ~x432 & ~x449 & ~x640 & ~x755;
assign c1337 = ~x4 & ~x139 & ~x357 & ~x433 & ~x434 & ~x458 & ~x514 & ~x542 & ~x569 & ~x613 & ~x615 & ~x704 & ~x781;
assign c1339 = ~x16 & ~x54 & ~x72 & ~x112 & ~x238 & ~x239 & ~x266 & ~x294 & ~x364 & ~x420 & ~x702 & ~x705 & ~x729 & ~x730 & ~x732;
assign c1341 =  x394 & ~x27 & ~x750;
assign c1343 =  x254 & ~x4 & ~x728 & ~x760;
assign c1345 =  x520 &  x548 &  x574 &  x600 & ~x614 & ~x753;
assign c1347 =  x100 & ~x187 & ~x338 & ~x362 & ~x513 & ~x541 & ~x624 & ~x652;
assign c1349 =  x424 &  x508 & ~x226 & ~x255 & ~x458 & ~x689;
assign c1351 =  x375 & ~x107 & ~x468 & ~x523;
assign c1353 = ~x52 & ~x71 & ~x211 & ~x266 & ~x267 & ~x668 & ~x675 & ~x705 & ~x732 & ~x761 & ~x776;
assign c1355 =  x317 &  x400 & ~x8 & ~x139 & ~x393 & ~x420 & ~x614 & ~x645 & ~x648 & ~x675 & ~x676 & ~x705 & ~x730 & ~x758;
assign c1357 = ~x140 & ~x245 & ~x248 & ~x273 & ~x276 & ~x349 & ~x378 & ~x406 & ~x433 & ~x461 & ~x462 & ~x489 & ~x683 & ~x754;
assign c1359 = ~x23 & ~x84 & ~x140 & ~x251 & ~x336 & ~x337 & ~x374 & ~x376 & ~x402 & ~x403 & ~x404 & ~x420 & ~x430 & ~x486 & ~x543 & ~x587 & ~x626 & ~x644 & ~x709 & ~x729 & ~x730 & ~x766;
assign c1361 = ~x31 & ~x73 & ~x136 & ~x156 & ~x211 & ~x239 & ~x310 & ~x365 & ~x448 & ~x504 & ~x522 & ~x550 & ~x577 & ~x604 & ~x672;
assign c1363 = ~x3 & ~x6 & ~x9 & ~x34 & ~x55 & ~x82 & ~x276 & ~x578 & ~x662 & ~x688 & ~x713 & ~x717 & ~x718 & ~x768;
assign c1365 =  x377 &  x458 &  x513 & ~x8 & ~x54 & ~x80 & ~x109 & ~x223 & ~x332 & ~x388 & ~x783;
assign c1367 =  x350 & ~x68 & ~x76 & ~x123 & ~x439 & ~x441 & ~x535 & ~x590 & ~x669 & ~x730;
assign c1369 =  x185 & ~x36 & ~x98 & ~x196 & ~x224 & ~x469 & ~x472 & ~x475 & ~x585 & ~x616 & ~x640 & ~x643 & ~x753 & ~x761;
assign c1371 = ~x4 & ~x43 & ~x71 & ~x99 & ~x112 & ~x140 & ~x162 & ~x217 & ~x248 & ~x307 & ~x434 & ~x634 & ~x691 & ~x749 & ~x773 & ~x783;
assign c1373 = ~x51 & ~x86 & ~x190 & ~x202 & ~x386 & ~x438 & ~x465 & ~x467 & ~x521 & ~x549 & ~x611 & ~x773;
assign c1375 =  x375 & ~x0 & ~x80 & ~x133 & ~x137 & ~x556 & ~x605 & ~x756 & ~x758;
assign c1377 =  x371 & ~x202 & ~x332 & ~x732;
assign c1379 =  x676 & ~x5 & ~x7 & ~x62 & ~x177 & ~x260 & ~x278 & ~x757;
assign c1381 =  x547 &  x600 &  x601 & ~x1 & ~x26 & ~x29 & ~x32 & ~x80 & ~x87 & ~x141 & ~x309 & ~x336 & ~x364 & ~x365 & ~x474 & ~x501 & ~x502 & ~x531 & ~x532 & ~x560 & ~x617 & ~x644 & ~x700 & ~x755 & ~x777;
assign c1383 =  x316 &  x344 &  x371 & ~x6 & ~x28 & ~x31 & ~x49 & ~x84 & ~x85 & ~x138 & ~x201 & ~x224 & ~x448 & ~x731 & ~x732 & ~x782;
assign c1385 =  x312 &  x467 & ~x331 & ~x388 & ~x771 & ~x773 & ~x777;
assign c1387 = ~x0 & ~x4 & ~x29 & ~x55 & ~x58 & ~x59 & ~x134 & ~x140 & ~x141 & ~x142 & ~x220 & ~x224 & ~x250 & ~x487 & ~x488 & ~x515 & ~x543 & ~x547 & ~x572 & ~x599 & ~x627 & ~x655 & ~x657 & ~x711 & ~x738 & ~x753;
assign c1389 =  x315 & ~x33 & ~x51 & ~x90 & ~x117 & ~x142 & ~x143 & ~x144 & ~x146 & ~x201 & ~x252 & ~x302 & ~x303 & ~x308 & ~x330 & ~x331 & ~x358 & ~x445 & ~x759 & ~x760 & ~x761;
assign c1391 =  x612 & ~x0 & ~x3 & ~x17 & ~x26 & ~x31 & ~x46 & ~x54 & ~x56 & ~x82 & ~x168 & ~x224 & ~x335 & ~x336 & ~x393 & ~x579 & ~x580 & ~x606 & ~x607 & ~x608 & ~x633 & ~x634 & ~x635 & ~x636 & ~x661 & ~x662 & ~x663 & ~x687;
assign c1393 =  x664 & ~x8 & ~x52 & ~x85 & ~x87 & ~x614 & ~x695 & ~x726 & ~x760 & ~x762 & ~x766;
assign c1395 =  x718 & ~x37 & ~x52 & ~x77 & ~x413 & ~x553 & ~x589 & ~x619 & ~x644 & ~x699;
assign c1397 =  x520 &  x576 & ~x83 & ~x169 & ~x254 & ~x374 & ~x401 & ~x429 & ~x457 & ~x476 & ~x559 & ~x615 & ~x643 & ~x645 & ~x701 & ~x755;
assign c1399 =  x469 & ~x45 & ~x474 & ~x664 & ~x692 & ~x717 & ~x719 & ~x721 & ~x747 & ~x772 & ~x778;
assign c1401 =  x318 & ~x257 & ~x312 & ~x730 & ~x731;
assign c1403 =  x389;
assign c1405 =  x433 & ~x10 & ~x12 & ~x25 & ~x38 & ~x39 & ~x53 & ~x66 & ~x447 & ~x732 & ~x734 & ~x758;
assign c1407 =  x523 & ~x52 & ~x56 & ~x107 & ~x135 & ~x166 & ~x167 & ~x193 & ~x197 & ~x224 & ~x226 & ~x274 & ~x296 & ~x303 & ~x352 & ~x379 & ~x392 & ~x779;
assign c1409 =  x208 &  x632 &  x659 &  x686;
assign c1411 =  x632 &  x659 &  x687 & ~x513 & ~x648 & ~x701;
assign c1413 =  x164 &  x323;
assign c1415 =  x295 & ~x11 & ~x12 & ~x13 & ~x23 & ~x24 & ~x37 & ~x38 & ~x39 & ~x40 & ~x58 & ~x64 & ~x65 & ~x86 & ~x93 & ~x198 & ~x227 & ~x252 & ~x280 & ~x282 & ~x499 & ~x500 & ~x559 & ~x699 & ~x729 & ~x755;
assign c1417 = ~x12 & ~x33 & ~x224 & ~x247 & ~x441 & ~x487 & ~x503 & ~x551 & ~x554 & ~x592;
assign c1419 = ~x141 & ~x196 & ~x198 & ~x215 & ~x442 & ~x468 & ~x502 & ~x522 & ~x549 & ~x632 & ~x641 & ~x761 & ~x781;
assign c1421 = ~x0 & ~x26 & ~x196 & ~x280 & ~x577 & ~x597 & ~x605 & ~x606 & ~x635 & ~x659 & ~x662 & ~x680 & ~x689 & ~x690 & ~x708 & ~x714 & ~x715 & ~x765 & ~x771 & ~x775;
assign c1423 = ~x6 & ~x33 & ~x55 & ~x59 & ~x60 & ~x61 & ~x62 & ~x83 & ~x84 & ~x85 & ~x114 & ~x116 & ~x196 & ~x274 & ~x302 & ~x304 & ~x307 & ~x333 & ~x358 & ~x359 & ~x387 & ~x389 & ~x416 & ~x420 & ~x660 & ~x715 & ~x740 & ~x742 & ~x744 & ~x765 & ~x767 & ~x768 & ~x769 & ~x770;
assign c1425 =  x73 & ~x28 & ~x114 & ~x345 & ~x472 & ~x473 & ~x656;
assign c1427 =  x260 & ~x12 & ~x37 & ~x771;
assign c1429 =  x549 &  x603 & ~x25 & ~x322 & ~x757 & ~x778;
assign c1431 =  x80 & ~x219;
assign c1433 = ~x2 & ~x10 & ~x218 & ~x279 & ~x432 & ~x516 & ~x600 & ~x615 & ~x616 & ~x659 & ~x687 & ~x713;
assign c1435 =  x389 & ~x700;
assign c1437 =  x576 &  x603 &  x630 &  x657 & ~x0 & ~x27 & ~x51 & ~x52 & ~x55 & ~x168 & ~x252 & ~x335 & ~x336 & ~x477 & ~x479 & ~x503 & ~x504 & ~x529 & ~x530 & ~x534 & ~x561 & ~x562 & ~x585 & ~x586 & ~x588 & ~x590 & ~x615 & ~x673 & ~x700 & ~x701 & ~x730 & ~x754 & ~x755 & ~x781 & ~x783;
assign c1439 =  x165 & ~x274;
assign c1441 =  x634 &  x661 &  x687 &  x714 & ~x28 & ~x278 & ~x558 & ~x700 & ~x726;
assign c1443 =  x126 &  x182 & ~x162 & ~x241 & ~x533;
assign c1445 =  x397 &  x425 & ~x0 & ~x26 & ~x28 & ~x88 & ~x115 & ~x282 & ~x330 & ~x700;
assign c1447 = ~x1 & ~x56 & ~x82 & ~x114 & ~x139 & ~x223 & ~x247 & ~x362 & ~x436 & ~x547 & ~x604 & ~x605 & ~x631 & ~x686 & ~x766 & ~x767;
assign c1449 =  x517 &  x545 & ~x320 & ~x642 & ~x678 & ~x706;
assign c1451 = ~x97 & ~x456 & ~x543 & ~x616 & ~x624 & ~x639 & ~x652 & ~x766;
assign c1453 =  x491 &  x518 &  x545 & ~x29 & ~x31 & ~x81 & ~x109 & ~x167 & ~x188 & ~x218 & ~x222 & ~x223 & ~x244 & ~x245 & ~x250 & ~x254 & ~x273 & ~x274 & ~x275 & ~x280 & ~x283 & ~x301 & ~x337 & ~x391 & ~x448 & ~x532 & ~x559 & ~x588 & ~x614 & ~x642 & ~x754 & ~x757;
assign c1455 =  x462 &  x516 & ~x140 & ~x217 & ~x273 & ~x301 & ~x336 & ~x502 & ~x504 & ~x605;
assign c1457 =  x527 & ~x82 & ~x195 & ~x496 & ~x523;
assign c1459 =  x403 & ~x32 & ~x59 & ~x166 & ~x418 & ~x475 & ~x477 & ~x532 & ~x577 & ~x607 & ~x633 & ~x635 & ~x654 & ~x672;
assign c1461 =  x356 & ~x5 & ~x240 & ~x708 & ~x733;
assign c1463 = ~x197 & ~x440 & ~x443 & ~x459 & ~x487 & ~x496 & ~x514 & ~x515 & ~x523 & ~x541 & ~x569 & ~x580 & ~x596 & ~x597 & ~x616 & ~x625;
assign c1465 =  x487 &  x542 & ~x186 & ~x213 & ~x734;
assign c1467 = ~x1 & ~x2 & ~x30 & ~x54 & ~x56 & ~x81 & ~x82 & ~x87 & ~x112 & ~x116 & ~x139 & ~x144 & ~x190 & ~x198 & ~x218 & ~x219 & ~x221 & ~x223 & ~x246 & ~x247 & ~x253 & ~x278 & ~x279 & ~x307 & ~x309 & ~x335 & ~x336 & ~x361 & ~x418 & ~x419 & ~x447 & ~x503 & ~x576 & ~x603 & ~x628 & ~x629 & ~x656 & ~x657 & ~x671 & ~x711 & ~x729 & ~x755;
assign c1469 = ~x2 & ~x221 & ~x226 & ~x246 & ~x275 & ~x276 & ~x390 & ~x433 & ~x517 & ~x544 & ~x631 & ~x658 & ~x659 & ~x711 & ~x713 & ~x714 & ~x767 & ~x783;
assign c1471 =  x406 &  x486 & ~x344 & ~x372 & ~x400 & ~x781;
assign c1473 = ~x39 & ~x179 & ~x452 & ~x476 & ~x542 & ~x623 & ~x637 & ~x647 & ~x652 & ~x675 & ~x773 & ~x782;
assign c1475 =  x269 & ~x55 & ~x252 & ~x366 & ~x440 & ~x468 & ~x475 & ~x514 & ~x515 & ~x531 & ~x554 & ~x612 & ~x641 & ~x642 & ~x673 & ~x701;
assign c1477 =  x155 &  x211 &  x351 & ~x48 & ~x89 & ~x525 & ~x783;
assign c1479 =  x67 &  x93 &  x121 & ~x421 & ~x614 & ~x622 & ~x642 & ~x650;
assign c1481 =  x575 &  x629 &  x630 & ~x26 & ~x58 & ~x61 & ~x117 & ~x164 & ~x196 & ~x531 & ~x585 & ~x641 & ~x725 & ~x731 & ~x751;
assign c1483 =  x740 & ~x300 & ~x326 & ~x605;
assign c1485 =  x229 & ~x23 & ~x344 & ~x371 & ~x399 & ~x427 & ~x477 & ~x532 & ~x587 & ~x588 & ~x616 & ~x643 & ~x644 & ~x757;
assign c1487 = ~x5 & ~x27 & ~x85 & ~x139 & ~x356 & ~x412 & ~x440 & ~x468 & ~x495 & ~x542 & ~x570 & ~x582 & ~x762;
assign c1489 =  x423 & ~x5 & ~x27 & ~x55 & ~x83 & ~x84 & ~x111 & ~x112 & ~x166 & ~x168 & ~x170 & ~x196 & ~x197 & ~x224 & ~x252 & ~x274 & ~x642 & ~x728 & ~x755 & ~x773 & ~x783;
assign c1491 =  x241 &  x339 &  x367;
assign c1493 =  x184 &  x492 &  x548 & ~x511 & ~x542;
assign c1495 =  x603 &  x631 &  x657 & ~x280 & ~x609;
assign c1497 =  x129 &  x241 & ~x1 & ~x29 & ~x272 & ~x336 & ~x557 & ~x559 & ~x585;
assign c1499 =  x366 & ~x401;
assign c20 =  x161 & ~x262 & ~x399 & ~x426 & ~x545 & ~x546 & ~x573 & ~x629 & ~x683 & ~x711 & ~x740 & ~x776;
assign c22 =  x153 &  x181 &  x542 & ~x218 & ~x245 & ~x250 & ~x251 & ~x269 & ~x392 & ~x552 & ~x557 & ~x560 & ~x605 & ~x611 & ~x678 & ~x736 & ~x760 & ~x764;
assign c24 = ~x17 & ~x28 & ~x46 & ~x76 & ~x77 & ~x84 & ~x87 & ~x102 & ~x105 & ~x109 & ~x110 & ~x132 & ~x134 & ~x138 & ~x163 & ~x170 & ~x171 & ~x184 & ~x189 & ~x190 & ~x193 & ~x199 & ~x212 & ~x220 & ~x222 & ~x225 & ~x248 & ~x277 & ~x281 & ~x303 & ~x306 & ~x309 & ~x310 & ~x333 & ~x336 & ~x339 & ~x361 & ~x362 & ~x365 & ~x366 & ~x386 & ~x395 & ~x413 & ~x417 & ~x420 & ~x421 & ~x422 & ~x423 & ~x440 & ~x443 & ~x477 & ~x480 & ~x494 & ~x502 & ~x503 & ~x505 & ~x506 & ~x520 & ~x521 & ~x526 & ~x531 & ~x532 & ~x536 & ~x556 & ~x564 & ~x566 & ~x567 & ~x580 & ~x583 & ~x590 & ~x591 & ~x594 & ~x595 & ~x608 & ~x616 & ~x618 & ~x622 & ~x637 & ~x638 & ~x647 & ~x665 & ~x668 & ~x671 & ~x676 & ~x693 & ~x696 & ~x697 & ~x701 & ~x703 & ~x706 & ~x725 & ~x751 & ~x758 & ~x759;
assign c26 =  x371 & ~x0 & ~x2 & ~x3 & ~x4 & ~x18 & ~x20 & ~x21 & ~x23 & ~x24 & ~x25 & ~x26 & ~x27 & ~x28 & ~x29 & ~x30 & ~x31 & ~x32 & ~x49 & ~x51 & ~x52 & ~x53 & ~x54 & ~x55 & ~x56 & ~x58 & ~x60 & ~x61 & ~x78 & ~x79 & ~x80 & ~x82 & ~x83 & ~x84 & ~x85 & ~x86 & ~x87 & ~x88 & ~x107 & ~x108 & ~x109 & ~x112 & ~x113 & ~x114 & ~x115 & ~x116 & ~x136 & ~x138 & ~x139 & ~x140 & ~x141 & ~x142 & ~x143 & ~x163 & ~x164 & ~x165 & ~x168 & ~x169 & ~x170 & ~x171 & ~x172 & ~x191 & ~x192 & ~x193 & ~x194 & ~x196 & ~x197 & ~x198 & ~x220 & ~x221 & ~x223 & ~x224 & ~x225 & ~x226 & ~x227 & ~x247 & ~x248 & ~x249 & ~x251 & ~x254 & ~x255 & ~x275 & ~x277 & ~x278 & ~x279 & ~x280 & ~x304 & ~x305 & ~x306 & ~x309 & ~x310 & ~x311 & ~x332 & ~x333 & ~x334 & ~x338 & ~x360 & ~x361 & ~x362 & ~x363 & ~x365 & ~x366 & ~x367 & ~x388 & ~x390 & ~x391 & ~x392 & ~x394 & ~x416 & ~x417 & ~x419 & ~x420 & ~x421 & ~x422 & ~x444 & ~x446 & ~x447 & ~x448 & ~x450 & ~x471 & ~x472 & ~x473 & ~x476 & ~x477 & ~x478 & ~x498 & ~x499 & ~x500 & ~x501 & ~x503 & ~x506 & ~x519 & ~x527 & ~x528 & ~x529 & ~x530 & ~x531 & ~x532 & ~x546 & ~x547 & ~x555 & ~x556 & ~x557 & ~x558 & ~x560 & ~x561 & ~x562 & ~x573 & ~x574 & ~x575 & ~x584 & ~x585 & ~x586 & ~x587 & ~x589 & ~x601 & ~x602 & ~x613 & ~x614 & ~x615 & ~x616 & ~x617 & ~x641 & ~x642 & ~x644 & ~x645 & ~x669 & ~x670 & ~x671 & ~x672 & ~x673 & ~x674 & ~x697 & ~x698 & ~x699 & ~x700 & ~x725 & ~x726 & ~x727 & ~x728 & ~x729 & ~x730 & ~x731 & ~x752 & ~x754 & ~x755 & ~x756 & ~x757 & ~x758 & ~x780 & ~x781 & ~x782 & ~x783;
assign c28 = ~x0 & ~x2 & ~x3 & ~x22 & ~x26 & ~x27 & ~x32 & ~x33 & ~x51 & ~x52 & ~x55 & ~x58 & ~x72 & ~x78 & ~x84 & ~x86 & ~x88 & ~x107 & ~x108 & ~x109 & ~x110 & ~x115 & ~x116 & ~x135 & ~x137 & ~x138 & ~x139 & ~x140 & ~x143 & ~x144 & ~x161 & ~x162 & ~x163 & ~x164 & ~x168 & ~x170 & ~x171 & ~x190 & ~x191 & ~x193 & ~x195 & ~x198 & ~x199 & ~x200 & ~x219 & ~x224 & ~x225 & ~x227 & ~x244 & ~x245 & ~x247 & ~x248 & ~x250 & ~x280 & ~x285 & ~x303 & ~x305 & ~x324 & ~x333 & ~x334 & ~x335 & ~x351 & ~x360 & ~x361 & ~x363 & ~x364 & ~x379 & ~x391 & ~x407 & ~x422 & ~x446 & ~x447 & ~x474 & ~x505 & ~x531 & ~x559 & ~x561 & ~x562 & ~x587 & ~x588 & ~x614 & ~x617 & ~x640 & ~x646 & ~x668 & ~x670 & ~x672 & ~x690 & ~x695 & ~x698 & ~x700 & ~x726 & ~x728 & ~x754 & ~x755 & ~x756 & ~x782 & ~x783;
assign c210 = ~x3 & ~x5 & ~x6 & ~x27 & ~x55 & ~x168 & ~x305 & ~x306 & ~x360 & ~x362 & ~x365 & ~x370 & ~x371 & ~x372 & ~x387 & ~x389 & ~x391 & ~x393 & ~x398 & ~x399 & ~x415 & ~x416 & ~x419 & ~x445 & ~x447 & ~x450 & ~x454 & ~x456 & ~x472 & ~x474 & ~x480 & ~x482 & ~x484 & ~x500 & ~x503 & ~x506 & ~x507 & ~x509 & ~x511 & ~x512 & ~x528 & ~x531 & ~x536 & ~x556 & ~x560 & ~x562 & ~x564 & ~x565 & ~x566 & ~x571 & ~x589 & ~x591 & ~x594 & ~x597 & ~x598 & ~x599 & ~x615 & ~x616 & ~x618 & ~x620 & ~x622 & ~x623 & ~x624 & ~x626 & ~x627 & ~x643 & ~x653 & ~x670 & ~x674 & ~x676 & ~x678 & ~x698 & ~x701 & ~x713 & ~x729 & ~x730 & ~x755 & ~x783;
assign c212 =  x131 & ~x27 & ~x30 & ~x56 & ~x57 & ~x70 & ~x96 & ~x195 & ~x317 & ~x335 & ~x362 & ~x387 & ~x391 & ~x415 & ~x427 & ~x697 & ~x755 & ~x782;
assign c214 = ~x16 & ~x71 & ~x98 & ~x125 & ~x165 & ~x193 & ~x250 & ~x289 & ~x399 & ~x416 & ~x426 & ~x600 & ~x627 & ~x710 & ~x737;
assign c216 =  x133 & ~x2 & ~x55 & ~x168 & ~x196 & ~x247 & ~x249 & ~x251 & ~x278 & ~x279 & ~x304 & ~x307 & ~x345 & ~x361 & ~x363 & ~x371 & ~x398 & ~x399 & ~x419 & ~x454 & ~x510 & ~x700 & ~x756;
assign c218 = ~x3 & ~x5 & ~x24 & ~x26 & ~x30 & ~x59 & ~x60 & ~x125 & ~x139 & ~x166 & ~x169 & ~x223 & ~x279 & ~x281 & ~x291 & ~x346 & ~x361 & ~x363 & ~x373 & ~x400 & ~x456 & ~x484 & ~x539 & ~x712 & ~x740 & ~x742 & ~x768;
assign c220 =  x97 &  x125 &  x181 &  x209 &  x237 & ~x2 & ~x22 & ~x31 & ~x79 & ~x135 & ~x137 & ~x138 & ~x167 & ~x169 & ~x221 & ~x251 & ~x268 & ~x304 & ~x307 & ~x308 & ~x309 & ~x335 & ~x337 & ~x475 & ~x555 & ~x558 & ~x579 & ~x587 & ~x603 & ~x605 & ~x607 & ~x608 & ~x611 & ~x614 & ~x637 & ~x670 & ~x704 & ~x705 & ~x724 & ~x729 & ~x757 & ~x783;
assign c222 = ~x7 & ~x24 & ~x34 & ~x61 & ~x84 & ~x86 & ~x89 & ~x91 & ~x114 & ~x116 & ~x142 & ~x144 & ~x145 & ~x147 & ~x152 & ~x170 & ~x172 & ~x173 & ~x174 & ~x175 & ~x180 & ~x419 & ~x443 & ~x445 & ~x446 & ~x473 & ~x482 & ~x500 & ~x502 & ~x508 & ~x509 & ~x528 & ~x529 & ~x530 & ~x531 & ~x535 & ~x536 & ~x537 & ~x559 & ~x560 & ~x562 & ~x565 & ~x566 & ~x586 & ~x592 & ~x619 & ~x626 & ~x627 & ~x642 & ~x643 & ~x644 & ~x651 & ~x653 & ~x654 & ~x655 & ~x668 & ~x674 & ~x675 & ~x677 & ~x678 & ~x681 & ~x682 & ~x697 & ~x699 & ~x700 & ~x701 & ~x703 & ~x705 & ~x706 & ~x707 & ~x708 & ~x709 & ~x728 & ~x730 & ~x752 & ~x756 & ~x757 & ~x758 & ~x759 & ~x762 & ~x778 & ~x779 & ~x783;
assign c224 =  x597 & ~x3 & ~x27 & ~x28 & ~x50 & ~x57 & ~x59 & ~x80 & ~x84 & ~x86 & ~x107 & ~x108 & ~x109 & ~x114 & ~x134 & ~x141 & ~x164 & ~x166 & ~x167 & ~x169 & ~x171 & ~x172 & ~x199 & ~x219 & ~x221 & ~x222 & ~x224 & ~x226 & ~x227 & ~x247 & ~x252 & ~x278 & ~x305 & ~x309 & ~x334 & ~x361 & ~x362 & ~x393 & ~x420 & ~x446 & ~x448 & ~x475 & ~x477 & ~x505 & ~x547 & ~x559 & ~x573 & ~x575 & ~x587 & ~x613 & ~x614 & ~x629 & ~x645 & ~x671 & ~x698 & ~x729 & ~x755 & ~x782;
assign c226 =  x436 & ~x49 & ~x53 & ~x79 & ~x81 & ~x88 & ~x106 & ~x115 & ~x132 & ~x160 & ~x163 & ~x164 & ~x172 & ~x195 & ~x198 & ~x200 & ~x221 & ~x242 & ~x243 & ~x246 & ~x247 & ~x254 & ~x269 & ~x297 & ~x311 & ~x351 & ~x394 & ~x448 & ~x471 & ~x499 & ~x506 & ~x522 & ~x524 & ~x525 & ~x526 & ~x532 & ~x558 & ~x584 & ~x587 & ~x615 & ~x616 & ~x639 & ~x675 & ~x702 & ~x703 & ~x728 & ~x757 & ~x761;
assign c228 =  x73 &  x127 & ~x54 & ~x56 & ~x111 & ~x218 & ~x252 & ~x253 & ~x280 & ~x309 & ~x337 & ~x389 & ~x390 & ~x419 & ~x447 & ~x502 & ~x700 & ~x720 & ~x729 & ~x755 & ~x766 & ~x774 & ~x782;
assign c230 =  x322 &  x323 &  x630 & ~x3 & ~x59 & ~x87 & ~x194 & ~x208 & ~x473 & ~x611 & ~x637 & ~x639 & ~x750 & ~x783;
assign c232 = ~x1 & ~x3 & ~x140 & ~x222 & ~x224 & ~x251 & ~x280 & ~x307 & ~x334 & ~x360 & ~x361 & ~x390 & ~x399 & ~x415 & ~x417 & ~x425 & ~x427 & ~x454 & ~x473 & ~x499 & ~x500 & ~x501 & ~x503 & ~x506 & ~x507 & ~x511 & ~x527 & ~x528 & ~x531 & ~x542 & ~x557 & ~x558 & ~x566 & ~x568 & ~x587 & ~x593 & ~x595 & ~x596 & ~x598 & ~x611 & ~x616 & ~x619 & ~x626 & ~x627 & ~x639 & ~x641 & ~x653 & ~x668 & ~x674 & ~x675 & ~x677 & ~x701 & ~x702 & ~x706 & ~x707 & ~x708 & ~x725 & ~x732 & ~x733 & ~x742 & ~x757 & ~x760 & ~x761 & ~x768 & ~x780 & ~x781;
assign c234 =  x464 & ~x32 & ~x132 & ~x243 & ~x325 & ~x379 & ~x405;
assign c236 = ~x1 & ~x26 & ~x45 & ~x73 & ~x83 & ~x87 & ~x135 & ~x157 & ~x174 & ~x185 & ~x188 & ~x194 & ~x212 & ~x240 & ~x268 & ~x279 & ~x281 & ~x295 & ~x303 & ~x312 & ~x335 & ~x362 & ~x421 & ~x443 & ~x447 & ~x449 & ~x450 & ~x470 & ~x478 & ~x499 & ~x505 & ~x528 & ~x529 & ~x535 & ~x551 & ~x558 & ~x562 & ~x582 & ~x587 & ~x590 & ~x591 & ~x645 & ~x647 & ~x652 & ~x679 & ~x703 & ~x748 & ~x752 & ~x756 & ~x776;
assign c238 =  x189 & ~x346 & ~x388 & ~x454 & ~x538 & ~x714;
assign c240 = ~x140 & ~x319 & ~x320 & ~x334 & ~x359 & ~x363 & ~x389 & ~x398 & ~x399 & ~x416 & ~x421 & ~x445 & ~x447 & ~x460 & ~x473 & ~x506 & ~x511 & ~x532 & ~x539 & ~x586 & ~x589 & ~x592 & ~x593 & ~x595 & ~x614 & ~x627 & ~x642 & ~x646 & ~x651 & ~x681 & ~x704 & ~x707;
assign c242 = ~x3 & ~x29 & ~x51 & ~x52 & ~x53 & ~x55 & ~x78 & ~x82 & ~x84 & ~x110 & ~x137 & ~x140 & ~x143 & ~x156 & ~x168 & ~x199 & ~x246 & ~x275 & ~x278 & ~x304 & ~x305 & ~x308 & ~x335 & ~x385 & ~x387 & ~x392 & ~x413 & ~x419 & ~x426 & ~x439 & ~x443 & ~x448 & ~x455 & ~x466 & ~x470 & ~x483 & ~x493 & ~x501 & ~x502 & ~x510 & ~x520 & ~x521 & ~x531 & ~x535 & ~x551 & ~x556 & ~x560 & ~x582 & ~x589 & ~x596 & ~x597 & ~x620 & ~x621 & ~x641 & ~x645 & ~x663 & ~x664 & ~x681 & ~x695 & ~x701 & ~x755 & ~x762;
assign c244 =  x369 & ~x26 & ~x28 & ~x29 & ~x31 & ~x84 & ~x86 & ~x108 & ~x109 & ~x114 & ~x115 & ~x137 & ~x138 & ~x141 & ~x142 & ~x164 & ~x165 & ~x166 & ~x169 & ~x170 & ~x196 & ~x197 & ~x220 & ~x221 & ~x222 & ~x223 & ~x224 & ~x225 & ~x226 & ~x247 & ~x248 & ~x249 & ~x250 & ~x251 & ~x253 & ~x277 & ~x280 & ~x282 & ~x305 & ~x306 & ~x310 & ~x335 & ~x337 & ~x363 & ~x365 & ~x366 & ~x391 & ~x419 & ~x421 & ~x445 & ~x446 & ~x448 & ~x472 & ~x474 & ~x475 & ~x501 & ~x504 & ~x519 & ~x520 & ~x532 & ~x546 & ~x547 & ~x559 & ~x560 & ~x573 & ~x574 & ~x700 & ~x753 & ~x754 & ~x781;
assign c246 =  x464 & ~x0 & ~x30 & ~x55 & ~x79 & ~x107 & ~x109 & ~x112 & ~x136 & ~x142 & ~x199 & ~x221 & ~x245 & ~x250 & ~x254 & ~x269 & ~x270 & ~x324 & ~x351 & ~x420 & ~x504 & ~x526 & ~x551 & ~x557 & ~x583 & ~x608 & ~x609 & ~x610 & ~x611 & ~x613 & ~x615 & ~x639 & ~x669 & ~x671 & ~x700 & ~x726 & ~x730 & ~x731 & ~x734 & ~x760;
assign c248 =  x321 &  x345 & ~x1 & ~x2 & ~x3 & ~x23 & ~x24 & ~x27 & ~x32 & ~x52 & ~x54 & ~x56 & ~x57 & ~x58 & ~x59 & ~x60 & ~x80 & ~x82 & ~x87 & ~x88 & ~x107 & ~x108 & ~x111 & ~x133 & ~x134 & ~x139 & ~x141 & ~x142 & ~x144 & ~x145 & ~x161 & ~x167 & ~x168 & ~x169 & ~x172 & ~x192 & ~x194 & ~x196 & ~x220 & ~x221 & ~x222 & ~x225 & ~x277 & ~x278 & ~x336 & ~x364 & ~x390 & ~x392 & ~x417 & ~x419 & ~x445 & ~x446 & ~x448 & ~x471 & ~x472 & ~x476 & ~x477 & ~x498 & ~x501 & ~x503 & ~x504 & ~x505 & ~x524 & ~x527 & ~x530 & ~x532 & ~x550 & ~x551 & ~x555 & ~x558 & ~x587 & ~x610 & ~x611 & ~x636 & ~x638 & ~x639 & ~x640 & ~x641 & ~x642 & ~x646 & ~x648 & ~x649 & ~x669 & ~x677 & ~x678 & ~x679 & ~x680 & ~x703 & ~x705 & ~x707 & ~x708 & ~x725 & ~x729 & ~x732 & ~x733 & ~x754 & ~x780;
assign c250 =  x83;
assign c252 =  x427 &  x542 & ~x80 & ~x85 & ~x86 & ~x132 & ~x136 & ~x193 & ~x197 & ~x226 & ~x305 & ~x338 & ~x390 & ~x392 & ~x447 & ~x448 & ~x475 & ~x531 & ~x534 & ~x556 & ~x559 & ~x561 & ~x582 & ~x589 & ~x611 & ~x615 & ~x640 & ~x670 & ~x695 & ~x704 & ~x730 & ~x731;
assign c254 =  x157 &  x240 &  x296 & ~x301 & ~x318 & ~x361 & ~x367 & ~x385 & ~x412 & ~x414 & ~x416 & ~x425 & ~x469 & ~x471 & ~x473 & ~x474 & ~x500 & ~x528 & ~x561 & ~x563 & ~x585 & ~x588 & ~x590 & ~x591 & ~x637 & ~x649;
assign c256 =  x678 &  x732 & ~x491;
assign c258 = ~x1 & ~x112 & ~x276 & ~x305 & ~x390 & ~x400 & ~x418 & ~x426 & ~x453 & ~x455 & ~x509 & ~x544 & ~x626 & ~x627 & ~x629 & ~x652 & ~x654 & ~x657 & ~x680 & ~x700 & ~x707 & ~x735 & ~x740 & ~x757 & ~x760;
assign c260 = ~x0 & ~x26 & ~x166 & ~x193 & ~x221 & ~x240 & ~x248 & ~x274 & ~x275 & ~x276 & ~x289 & ~x302 & ~x324 & ~x352 & ~x361 & ~x380 & ~x408 & ~x409 & ~x436 & ~x463;
assign c262 =  x492 & ~x50 & ~x134 & ~x137 & ~x221 & ~x224 & ~x227 & ~x247 & ~x252 & ~x254 & ~x351 & ~x379 & ~x604;
assign c264 =  x310 & ~x152 & ~x179 & ~x453;
assign c266 =  x354 & ~x25 & ~x48 & ~x61 & ~x82 & ~x87 & ~x88 & ~x90 & ~x107 & ~x136 & ~x137 & ~x166 & ~x190 & ~x213 & ~x214 & ~x222 & ~x240 & ~x280 & ~x282 & ~x310 & ~x386 & ~x387 & ~x422 & ~x441 & ~x445 & ~x475 & ~x497 & ~x499 & ~x534 & ~x557 & ~x585 & ~x586 & ~x617 & ~x639 & ~x641 & ~x701 & ~x702 & ~x754 & ~x759;
assign c268 = ~x0 & ~x34 & ~x53 & ~x89 & ~x106 & ~x113 & ~x114 & ~x115 & ~x147 & ~x159 & ~x164 & ~x196 & ~x216 & ~x217 & ~x226 & ~x255 & ~x279 & ~x417 & ~x439 & ~x440 & ~x467 & ~x470 & ~x477 & ~x479 & ~x506 & ~x507 & ~x520 & ~x522 & ~x524 & ~x528 & ~x536 & ~x548 & ~x551 & ~x552 & ~x553 & ~x554 & ~x562 & ~x591 & ~x608 & ~x625 & ~x642 & ~x644 & ~x646 & ~x648 & ~x653 & ~x664 & ~x680 & ~x681 & ~x721 & ~x728 & ~x758 & ~x774 & ~x777 & ~x779;
assign c270 = ~x1 & ~x7 & ~x15 & ~x19 & ~x25 & ~x26 & ~x34 & ~x51 & ~x58 & ~x60 & ~x88 & ~x116 & ~x129 & ~x196 & ~x219 & ~x220 & ~x278 & ~x303 & ~x305 & ~x310 & ~x326 & ~x330 & ~x337 & ~x353 & ~x361 & ~x380 & ~x445 & ~x500 & ~x505 & ~x531 & ~x534 & ~x557 & ~x577 & ~x579 & ~x580 & ~x617 & ~x618 & ~x641 & ~x645 & ~x663 & ~x665 & ~x671 & ~x672 & ~x679 & ~x696 & ~x698 & ~x705 & ~x724 & ~x727 & ~x735 & ~x762;
assign c272 = ~x2 & ~x5 & ~x23 & ~x27 & ~x30 & ~x51 & ~x52 & ~x58 & ~x59 & ~x60 & ~x81 & ~x85 & ~x112 & ~x113 & ~x114 & ~x136 & ~x165 & ~x167 & ~x193 & ~x198 & ~x199 & ~x217 & ~x224 & ~x226 & ~x235 & ~x253 & ~x278 & ~x279 & ~x281 & ~x308 & ~x333 & ~x334 & ~x338 & ~x361 & ~x363 & ~x387 & ~x391 & ~x441 & ~x447 & ~x477 & ~x483 & ~x499 & ~x501 & ~x511 & ~x529 & ~x539 & ~x557 & ~x560 & ~x585 & ~x613 & ~x614 & ~x642 & ~x643 & ~x655 & ~x670 & ~x683 & ~x690 & ~x692 & ~x698 & ~x699 & ~x700 & ~x710 & ~x729 & ~x739;
assign c274 = ~x54 & ~x55 & ~x222 & ~x300 & ~x363 & ~x368 & ~x385 & ~x401 & ~x412 & ~x413 & ~x420 & ~x441 & ~x473 & ~x478 & ~x479 & ~x503 & ~x514 & ~x527 & ~x581 & ~x586 & ~x598 & ~x625 & ~x628 & ~x642 & ~x653 & ~x663 & ~x665 & ~x674 & ~x682 & ~x698 & ~x707 & ~x710 & ~x727 & ~x728 & ~x748 & ~x749 & ~x758 & ~x777;
assign c276 =  x426 & ~x25 & ~x27 & ~x29 & ~x31 & ~x55 & ~x57 & ~x61 & ~x81 & ~x87 & ~x109 & ~x110 & ~x113 & ~x116 & ~x136 & ~x137 & ~x142 & ~x143 & ~x145 & ~x162 & ~x165 & ~x168 & ~x188 & ~x192 & ~x196 & ~x197 & ~x198 & ~x199 & ~x218 & ~x219 & ~x227 & ~x244 & ~x248 & ~x252 & ~x253 & ~x270 & ~x278 & ~x281 & ~x307 & ~x310 & ~x335 & ~x336 & ~x391 & ~x419 & ~x422 & ~x446 & ~x450 & ~x502 & ~x503 & ~x505 & ~x506 & ~x533 & ~x559 & ~x561 & ~x582 & ~x584 & ~x586 & ~x587 & ~x589 & ~x610 & ~x611 & ~x612 & ~x613 & ~x616 & ~x617 & ~x640 & ~x641 & ~x643 & ~x644 & ~x672 & ~x695 & ~x696 & ~x698 & ~x702 & ~x725 & ~x729 & ~x757 & ~x758;
assign c278 = ~x40 & ~x68 & ~x82 & ~x84 & ~x94 & ~x95 & ~x389 & ~x390 & ~x444 & ~x452 & ~x460 & ~x473 & ~x506 & ~x507 & ~x591 & ~x619 & ~x648 & ~x649 & ~x655 & ~x676 & ~x681 & ~x700 & ~x708 & ~x710;
assign c280 =  x236 &  x435 &  x462 &  x489 &  x516 & ~x57 & ~x113 & ~x135 & ~x323 & ~x364 & ~x524 & ~x528 & ~x559 & ~x582 & ~x583 & ~x584 & ~x588 & ~x612 & ~x613 & ~x641 & ~x726 & ~x730 & ~x734 & ~x755;
assign c282 =  x102 &  x184 &  x464 & ~x28 & ~x82 & ~x85 & ~x362 & ~x386 & ~x417 & ~x499 & ~x609 & ~x620 & ~x665 & ~x701 & ~x758;
assign c284 = ~x29 & ~x32 & ~x52 & ~x56 & ~x115 & ~x143 & ~x157 & ~x166 & ~x184 & ~x197 & ~x249 & ~x253 & ~x276 & ~x277 & ~x278 & ~x279 & ~x307 & ~x309 & ~x362 & ~x416 & ~x418 & ~x439 & ~x465 & ~x472 & ~x491 & ~x493 & ~x494 & ~x503 & ~x518 & ~x520 & ~x547 & ~x549 & ~x553 & ~x565 & ~x577 & ~x578 & ~x593 & ~x755;
assign c286 = ~x31 & ~x55 & ~x57 & ~x192 & ~x246 & ~x247 & ~x250 & ~x274 & ~x305 & ~x306 & ~x334 & ~x344 & ~x372 & ~x389 & ~x400 & ~x407 & ~x434 & ~x462 & ~x503 & ~x517 & ~x518 & ~x573 & ~x574 & ~x748 & ~x756;
assign c288 =  x367 & ~x234 & ~x406 & ~x473;
assign c290 = ~x2 & ~x25 & ~x125 & ~x153 & ~x361 & ~x391 & ~x455 & ~x484 & ~x500 & ~x507 & ~x528 & ~x530 & ~x558 & ~x586 & ~x627 & ~x654 & ~x655 & ~x673 & ~x700 & ~x709 & ~x713 & ~x729 & ~x730 & ~x736 & ~x737 & ~x739 & ~x741 & ~x755 & ~x757 & ~x768 & ~x782;
assign c292 =  x102 & ~x194 & ~x252 & ~x385 & ~x488 & ~x503 & ~x532 & ~x557 & ~x558 & ~x588 & ~x613 & ~x618 & ~x619 & ~x664 & ~x666 & ~x700 & ~x730 & ~x731 & ~x752;
assign c294 =  x296 & ~x22 & ~x54 & ~x132 & ~x138 & ~x167 & ~x195 & ~x196 & ~x356 & ~x384 & ~x412 & ~x413 & ~x424 & ~x441 & ~x443 & ~x451 & ~x452 & ~x469 & ~x470 & ~x474 & ~x482 & ~x484 & ~x498 & ~x501 & ~x502 & ~x524 & ~x525 & ~x526 & ~x533 & ~x540 & ~x559 & ~x560 & ~x561 & ~x569 & ~x584 & ~x596 & ~x613 & ~x618 & ~x623 & ~x626 & ~x637 & ~x647 & ~x650 & ~x653 & ~x699 & ~x701 & ~x705 & ~x706 & ~x726 & ~x727 & ~x729 & ~x735 & ~x750 & ~x779 & ~x781;
assign c296 =  x733 & ~x16 & ~x218 & ~x518 & ~x747;
assign c298 =  x506 & ~x426 & ~x548;
assign c2100 =  x518 & ~x26 & ~x29 & ~x55 & ~x111 & ~x115 & ~x139 & ~x142 & ~x165 & ~x225 & ~x249 & ~x252 & ~x297 & ~x298 & ~x300 & ~x309 & ~x352 & ~x353 & ~x380 & ~x419 & ~x552 & ~x559 & ~x577 & ~x578 & ~x580 & ~x588 & ~x603 & ~x608 & ~x631 & ~x633 & ~x637 & ~x661 & ~x696 & ~x725 & ~x729 & ~x734;
assign c2102 = ~x16 & ~x25 & ~x53 & ~x58 & ~x81 & ~x82 & ~x84 & ~x85 & ~x86 & ~x87 & ~x141 & ~x166 & ~x168 & ~x223 & ~x248 & ~x275 & ~x277 & ~x289 & ~x306 & ~x307 & ~x332 & ~x344 & ~x361 & ~x372 & ~x417 & ~x435 & ~x446 & ~x503 & ~x602 & ~x629 & ~x655 & ~x682 & ~x728 & ~x776;
assign c2104 =  x156 &  x159 & ~x27 & ~x55 & ~x58 & ~x85 & ~x96 & ~x139 & ~x251 & ~x272 & ~x274 & ~x277 & ~x278 & ~x280 & ~x302 & ~x303 & ~x305 & ~x307 & ~x330 & ~x331 & ~x334 & ~x335 & ~x359 & ~x363 & ~x388 & ~x391 & ~x415 & ~x416 & ~x417 & ~x420 & ~x445 & ~x531 & ~x588 & ~x673 & ~x701 & ~x778;
assign c2106 =  x674;
assign c2108 = ~x4 & ~x85 & ~x306 & ~x310 & ~x338 & ~x356 & ~x385 & ~x387 & ~x396 & ~x418 & ~x420 & ~x421 & ~x438 & ~x449 & ~x451 & ~x473 & ~x485 & ~x499 & ~x503 & ~x508 & ~x531 & ~x535 & ~x540 & ~x550 & ~x579 & ~x584 & ~x591 & ~x592 & ~x597 & ~x598 & ~x599 & ~x621 & ~x626 & ~x627 & ~x638 & ~x670 & ~x690 & ~x704 & ~x718 & ~x723 & ~x782;
assign c2110 =  x411 & ~x28 & ~x51 & ~x54 & ~x191 & ~x192 & ~x193 & ~x219 & ~x245 & ~x261 & ~x303 & ~x548 & ~x575 & ~x665;
assign c2112 = ~x0 & ~x4 & ~x27 & ~x34 & ~x37 & ~x61 & ~x107 & ~x109 & ~x112 & ~x140 & ~x252 & ~x300 & ~x301 & ~x306 & ~x329 & ~x357 & ~x358 & ~x363 & ~x385 & ~x388 & ~x396 & ~x398 & ~x399 & ~x429 & ~x453 & ~x455 & ~x457 & ~x479 & ~x481 & ~x482 & ~x497 & ~x501 & ~x502 & ~x510 & ~x512 & ~x513 & ~x527 & ~x537 & ~x541 & ~x557 & ~x559 & ~x563 & ~x565 & ~x579 & ~x584 & ~x615 & ~x616 & ~x620 & ~x621 & ~x624 & ~x626 & ~x635 & ~x649 & ~x652 & ~x654 & ~x666 & ~x672 & ~x677 & ~x678 & ~x681 & ~x691 & ~x704 & ~x706 & ~x707 & ~x710 & ~x727 & ~x729 & ~x734 & ~x758 & ~x763 & ~x778;
assign c2114 =  x412 & ~x234 & ~x247 & ~x316 & ~x407 & ~x463;
assign c2116 =  x187 & ~x4 & ~x23 & ~x25 & ~x26 & ~x84 & ~x307 & ~x318 & ~x319 & ~x332 & ~x333 & ~x335 & ~x344 & ~x345 & ~x361 & ~x372 & ~x389 & ~x391 & ~x392 & ~x401 & ~x419 & ~x427 & ~x443 & ~x444 & ~x445 & ~x446 & ~x448 & ~x455 & ~x456 & ~x472 & ~x473 & ~x474 & ~x483 & ~x502 & ~x503 & ~x505 & ~x539 & ~x559 & ~x588 & ~x644 & ~x673 & ~x700 & ~x729 & ~x759;
assign c2118 =  x344 &  x372 & ~x0 & ~x6 & ~x7 & ~x22 & ~x56 & ~x57 & ~x80 & ~x81 & ~x86 & ~x89 & ~x90 & ~x107 & ~x111 & ~x112 & ~x113 & ~x114 & ~x116 & ~x117 & ~x135 & ~x138 & ~x142 & ~x143 & ~x144 & ~x145 & ~x160 & ~x162 & ~x164 & ~x165 & ~x168 & ~x174 & ~x193 & ~x194 & ~x201 & ~x219 & ~x222 & ~x227 & ~x229 & ~x253 & ~x254 & ~x281 & ~x283 & ~x359 & ~x363 & ~x364 & ~x390 & ~x414 & ~x416 & ~x417 & ~x418 & ~x445 & ~x447 & ~x448 & ~x450 & ~x452 & ~x453 & ~x472 & ~x473 & ~x475 & ~x477 & ~x480 & ~x499 & ~x502 & ~x506 & ~x508 & ~x533 & ~x556 & ~x557 & ~x560 & ~x563 & ~x564 & ~x583 & ~x588 & ~x610 & ~x611 & ~x614 & ~x615 & ~x616 & ~x618 & ~x620 & ~x621 & ~x637 & ~x643 & ~x644 & ~x645 & ~x648 & ~x649 & ~x665 & ~x667 & ~x670 & ~x672 & ~x677 & ~x694 & ~x695 & ~x701 & ~x702 & ~x703 & ~x705 & ~x728 & ~x732 & ~x733 & ~x751 & ~x756 & ~x759 & ~x761 & ~x762 & ~x779 & ~x783;
assign c2120 =  x438 & ~x4 & ~x24 & ~x27 & ~x28 & ~x29 & ~x32 & ~x47 & ~x57 & ~x58 & ~x59 & ~x60 & ~x78 & ~x79 & ~x82 & ~x83 & ~x86 & ~x104 & ~x106 & ~x107 & ~x111 & ~x112 & ~x138 & ~x139 & ~x140 & ~x162 & ~x165 & ~x166 & ~x167 & ~x169 & ~x190 & ~x192 & ~x194 & ~x195 & ~x200 & ~x220 & ~x221 & ~x225 & ~x227 & ~x246 & ~x249 & ~x250 & ~x253 & ~x269 & ~x271 & ~x273 & ~x274 & ~x279 & ~x280 & ~x297 & ~x308 & ~x325 & ~x327 & ~x334 & ~x335 & ~x352 & ~x364 & ~x391 & ~x419 & ~x448 & ~x475 & ~x476 & ~x503 & ~x530 & ~x531 & ~x532 & ~x533 & ~x550 & ~x559 & ~x561 & ~x578 & ~x579 & ~x580 & ~x581 & ~x582 & ~x588 & ~x608 & ~x610 & ~x611 & ~x614 & ~x637 & ~x641 & ~x669 & ~x697 & ~x700 & ~x701 & ~x706 & ~x727 & ~x729 & ~x758 & ~x759 & ~x762;
assign c2122 =  x427 & ~x3 & ~x4 & ~x24 & ~x28 & ~x32 & ~x52 & ~x54 & ~x56 & ~x79 & ~x89 & ~x105 & ~x112 & ~x113 & ~x116 & ~x132 & ~x136 & ~x137 & ~x140 & ~x161 & ~x171 & ~x172 & ~x191 & ~x192 & ~x193 & ~x194 & ~x220 & ~x223 & ~x250 & ~x254 & ~x276 & ~x278 & ~x283 & ~x308 & ~x332 & ~x335 & ~x339 & ~x366 & ~x394 & ~x418 & ~x420 & ~x445 & ~x473 & ~x474 & ~x478 & ~x531 & ~x534 & ~x556 & ~x558 & ~x584 & ~x587 & ~x590 & ~x606 & ~x607 & ~x617 & ~x635 & ~x637 & ~x639 & ~x640 & ~x643 & ~x644 & ~x665 & ~x670 & ~x671 & ~x674 & ~x694 & ~x729 & ~x757 & ~x758 & ~x783;
assign c2124 =  x129 &  x156 & ~x0 & ~x29 & ~x57 & ~x97 & ~x222 & ~x244 & ~x248 & ~x249 & ~x250 & ~x252 & ~x274 & ~x275 & ~x277 & ~x289 & ~x331 & ~x332 & ~x390 & ~x391 & ~x418 & ~x469 & ~x472 & ~x644 & ~x746 & ~x752 & ~x780 & ~x781;
assign c2126 =  x506 &  x618 &  x674;
assign c2128 =  x298 & ~x1 & ~x2 & ~x23 & ~x27 & ~x30 & ~x32 & ~x33 & ~x83 & ~x84 & ~x141 & ~x143 & ~x156 & ~x165 & ~x166 & ~x170 & ~x171 & ~x185 & ~x196 & ~x197 & ~x211 & ~x224 & ~x253 & ~x335 & ~x358 & ~x359 & ~x360 & ~x361 & ~x363 & ~x444 & ~x473 & ~x475 & ~x500 & ~x519 & ~x530 & ~x531 & ~x559 & ~x729;
assign c2130 =  x216 & ~x5 & ~x152 & ~x179 & ~x374 & ~x388 & ~x389 & ~x391 & ~x472 & ~x477 & ~x483 & ~x511 & ~x528 & ~x530 & ~x539 & ~x567 & ~x591 & ~x595 & ~x669 & ~x697;
assign c2132 =  x678 & ~x16 & ~x31 & ~x82 & ~x110 & ~x193 & ~x195 & ~x248 & ~x278 & ~x308 & ~x364 & ~x390 & ~x416 & ~x463 & ~x490 & ~x545 & ~x573 & ~x600 & ~x755 & ~x757;
assign c2134 =  x95 & ~x134 & ~x146 & ~x174 & ~x184 & ~x224 & ~x247 & ~x279 & ~x336 & ~x441 & ~x466 & ~x493 & ~x499 & ~x529 & ~x536 & ~x538 & ~x578 & ~x594 & ~x651 & ~x666;
assign c2136 =  x560;
assign c2138 =  x455 &  x483 & ~x0 & ~x1 & ~x6 & ~x26 & ~x27 & ~x31 & ~x47 & ~x54 & ~x55 & ~x78 & ~x79 & ~x80 & ~x82 & ~x84 & ~x88 & ~x106 & ~x109 & ~x111 & ~x134 & ~x140 & ~x142 & ~x160 & ~x162 & ~x164 & ~x165 & ~x166 & ~x167 & ~x168 & ~x193 & ~x197 & ~x220 & ~x221 & ~x248 & ~x253 & ~x254 & ~x255 & ~x278 & ~x279 & ~x280 & ~x304 & ~x309 & ~x335 & ~x336 & ~x337 & ~x366 & ~x391 & ~x393 & ~x416 & ~x417 & ~x445 & ~x446 & ~x449 & ~x474 & ~x475 & ~x500 & ~x503 & ~x505 & ~x529 & ~x530 & ~x533 & ~x535 & ~x536 & ~x560 & ~x582 & ~x584 & ~x586 & ~x587 & ~x588 & ~x615 & ~x616 & ~x619 & ~x620 & ~x640 & ~x642 & ~x644 & ~x667 & ~x670 & ~x672 & ~x674 & ~x675 & ~x676 & ~x695 & ~x700 & ~x701 & ~x702 & ~x723 & ~x724 & ~x731 & ~x751 & ~x755 & ~x759 & ~x760 & ~x781;
assign c2140 =  x492 & ~x7 & ~x112 & ~x140 & ~x335 & ~x389 & ~x427 & ~x447 & ~x455 & ~x476 & ~x479 & ~x483 & ~x537 & ~x538 & ~x539 & ~x540 & ~x566 & ~x569 & ~x588 & ~x596 & ~x599 & ~x625 & ~x642 & ~x646 & ~x673 & ~x704 & ~x741;
assign c2142 =  x183 & ~x1 & ~x4 & ~x26 & ~x55 & ~x58 & ~x85 & ~x108 & ~x110 & ~x140 & ~x271 & ~x299 & ~x320 & ~x327 & ~x328 & ~x330 & ~x335 & ~x344 & ~x355 & ~x356 & ~x359 & ~x364 & ~x384 & ~x394 & ~x395 & ~x411 & ~x415 & ~x417 & ~x419 & ~x422 & ~x442 & ~x444 & ~x451 & ~x453 & ~x473 & ~x474 & ~x478 & ~x499 & ~x501 & ~x502 & ~x504 & ~x530 & ~x531 & ~x535 & ~x555 & ~x563 & ~x582 & ~x586 & ~x592 & ~x610 & ~x615 & ~x618 & ~x619 & ~x620 & ~x647 & ~x670 & ~x672 & ~x673 & ~x678 & ~x699 & ~x702 & ~x704 & ~x705 & ~x706 & ~x731 & ~x732 & ~x733 & ~x757;
assign c2144 =  x380 &  x460 & ~x88 & ~x133 & ~x139 & ~x142 & ~x170 & ~x191 & ~x194 & ~x212 & ~x213 & ~x218 & ~x224 & ~x248 & ~x278 & ~x442 & ~x466 & ~x469 & ~x471 & ~x492 & ~x522 & ~x530 & ~x549 & ~x550 & ~x647 & ~x671 & ~x674 & ~x676 & ~x699 & ~x703 & ~x733 & ~x759;
assign c2146 =  x477 & ~x425;
assign c2148 = ~x1 & ~x27 & ~x31 & ~x32 & ~x96 & ~x112 & ~x152 & ~x391 & ~x404 & ~x425 & ~x431 & ~x513 & ~x514 & ~x596 & ~x768 & ~x769 & ~x778;
assign c2150 =  x315 & ~x27 & ~x52 & ~x56 & ~x81 & ~x112 & ~x117 & ~x170 & ~x195 & ~x360 & ~x385 & ~x442 & ~x449 & ~x470 & ~x500 & ~x501 & ~x503 & ~x507 & ~x524 & ~x528 & ~x563 & ~x580 & ~x590 & ~x607 & ~x608 & ~x611 & ~x613 & ~x620 & ~x670 & ~x674 & ~x694 & ~x705 & ~x729 & ~x732 & ~x736 & ~x754 & ~x757 & ~x761 & ~x762 & ~x781;
assign c2152 =  x349 & ~x1 & ~x3 & ~x28 & ~x31 & ~x80 & ~x90 & ~x111 & ~x136 & ~x138 & ~x140 & ~x164 & ~x190 & ~x201 & ~x218 & ~x223 & ~x243 & ~x250 & ~x252 & ~x262 & ~x291 & ~x306 & ~x334 & ~x363 & ~x393 & ~x417 & ~x420 & ~x503 & ~x530 & ~x563 & ~x606 & ~x607 & ~x615 & ~x637 & ~x639 & ~x666 & ~x696 & ~x758 & ~x779 & ~x780;
assign c2154 = ~x1 & ~x2 & ~x22 & ~x23 & ~x31 & ~x52 & ~x54 & ~x78 & ~x82 & ~x86 & ~x88 & ~x89 & ~x108 & ~x137 & ~x190 & ~x192 & ~x194 & ~x196 & ~x199 & ~x214 & ~x218 & ~x219 & ~x222 & ~x229 & ~x240 & ~x241 & ~x243 & ~x248 & ~x249 & ~x251 & ~x256 & ~x257 & ~x268 & ~x275 & ~x332 & ~x333 & ~x334 & ~x337 & ~x338 & ~x339 & ~x357 & ~x366 & ~x367 & ~x388 & ~x391 & ~x395 & ~x413 & ~x418 & ~x442 & ~x445 & ~x447 & ~x467 & ~x470 & ~x494 & ~x495 & ~x500 & ~x505 & ~x521 & ~x524 & ~x525 & ~x530 & ~x531 & ~x533 & ~x536 & ~x552 & ~x553 & ~x558 & ~x564 & ~x582 & ~x583 & ~x586 & ~x608 & ~x611 & ~x615 & ~x641 & ~x643 & ~x645 & ~x647 & ~x649 & ~x669 & ~x673 & ~x676 & ~x690 & ~x698 & ~x700 & ~x702 & ~x704 & ~x705 & ~x706 & ~x722 & ~x735 & ~x748 & ~x749 & ~x755 & ~x757 & ~x760 & ~x761 & ~x762 & ~x763 & ~x776 & ~x780;
assign c2156 =  x408 &  x435 &  x462 &  x463 & ~x32 & ~x84 & ~x114 & ~x118 & ~x165 & ~x192 & ~x193 & ~x194 & ~x361 & ~x387 & ~x390 & ~x392 & ~x416 & ~x417 & ~x418 & ~x419 & ~x439 & ~x440 & ~x444 & ~x446 & ~x466 & ~x475 & ~x479 & ~x494 & ~x498 & ~x523 & ~x524 & ~x533 & ~x562 & ~x569 & ~x586 & ~x589 & ~x607 & ~x611 & ~x615 & ~x618 & ~x650 & ~x651 & ~x670 & ~x696 & ~x697 & ~x702 & ~x729 & ~x755 & ~x757 & ~x781;
assign c2158 =  x453 &  x481 &  x509 &  x537 & ~x4 & ~x28 & ~x29 & ~x30 & ~x81 & ~x84 & ~x106 & ~x108 & ~x109 & ~x111 & ~x136 & ~x137 & ~x138 & ~x141 & ~x142 & ~x162 & ~x163 & ~x168 & ~x190 & ~x194 & ~x195 & ~x219 & ~x220 & ~x222 & ~x250 & ~x251 & ~x252 & ~x254 & ~x276 & ~x277 & ~x281 & ~x282 & ~x307 & ~x310 & ~x336 & ~x338 & ~x363 & ~x393 & ~x419 & ~x446 & ~x474 & ~x501 & ~x502 & ~x504 & ~x558 & ~x559 & ~x562 & ~x587 & ~x588 & ~x589 & ~x616 & ~x617 & ~x641 & ~x645 & ~x672 & ~x673 & ~x701 & ~x727 & ~x755 & ~x758 & ~x782;
assign c2160 = ~x0 & ~x3 & ~x29 & ~x86 & ~x101 & ~x102 & ~x129 & ~x131 & ~x137 & ~x163 & ~x169 & ~x170 & ~x183 & ~x185 & ~x200 & ~x212 & ~x227 & ~x239 & ~x255 & ~x303 & ~x305 & ~x309 & ~x337 & ~x363 & ~x385 & ~x388 & ~x389 & ~x391 & ~x415 & ~x416 & ~x442 & ~x443 & ~x467 & ~x494 & ~x495 & ~x520 & ~x521 & ~x525 & ~x526 & ~x549 & ~x578 & ~x579 & ~x589 & ~x595 & ~x608 & ~x623 & ~x650 & ~x651 & ~x652 & ~x726;
assign c2162 =  x518 & ~x64 & ~x146 & ~x349 & ~x370 & ~x389 & ~x391 & ~x399 & ~x427 & ~x511 & ~x619 & ~x668 & ~x680 & ~x705 & ~x731 & ~x733 & ~x756 & ~x758 & ~x782;
assign c2164 = ~x6 & ~x26 & ~x27 & ~x28 & ~x35 & ~x53 & ~x59 & ~x79 & ~x80 & ~x86 & ~x91 & ~x101 & ~x106 & ~x116 & ~x159 & ~x162 & ~x170 & ~x184 & ~x212 & ~x219 & ~x329 & ~x330 & ~x337 & ~x358 & ~x364 & ~x387 & ~x391 & ~x393 & ~x418 & ~x422 & ~x440 & ~x448 & ~x449 & ~x450 & ~x467 & ~x477 & ~x498 & ~x502 & ~x508 & ~x524 & ~x530 & ~x548 & ~x579 & ~x591 & ~x622 & ~x637 & ~x643 & ~x646 & ~x648 & ~x650 & ~x653 & ~x670 & ~x673 & ~x679 & ~x694 & ~x697 & ~x700 & ~x701 & ~x706 & ~x726 & ~x733 & ~x752 & ~x761;
assign c2166 = ~x55 & ~x69 & ~x70 & ~x84 & ~x221 & ~x224 & ~x246 & ~x247 & ~x251 & ~x263 & ~x284 & ~x289 & ~x305 & ~x310 & ~x312 & ~x316 & ~x336 & ~x340 & ~x389 & ~x390 & ~x391 & ~x392 & ~x415 & ~x418 & ~x420 & ~x442 & ~x448 & ~x510 & ~x566 & ~x668 & ~x693 & ~x728 & ~x781;
assign c2168 =  x96 &  x462 &  x489 &  x516 & ~x23 & ~x51 & ~x52 & ~x103 & ~x104 & ~x107 & ~x165 & ~x171 & ~x188 & ~x189 & ~x221 & ~x224 & ~x243 & ~x310 & ~x504 & ~x527 & ~x553 & ~x557 & ~x578 & ~x583 & ~x584 & ~x638 & ~x645 & ~x678 & ~x705 & ~x706;
assign c2170 = ~x1 & ~x62 & ~x85 & ~x198 & ~x223 & ~x227 & ~x335 & ~x358 & ~x359 & ~x362 & ~x371 & ~x388 & ~x389 & ~x394 & ~x421 & ~x424 & ~x429 & ~x446 & ~x476 & ~x486 & ~x499 & ~x503 & ~x514 & ~x525 & ~x529 & ~x533 & ~x534 & ~x538 & ~x542 & ~x555 & ~x562 & ~x564 & ~x569 & ~x588 & ~x598 & ~x599 & ~x600 & ~x617 & ~x624 & ~x625 & ~x642 & ~x655 & ~x665 & ~x668 & ~x673 & ~x692 & ~x719 & ~x732 & ~x753 & ~x757 & ~x758 & ~x761 & ~x780;
assign c2172 =  x431 & ~x32 & ~x58 & ~x59 & ~x85 & ~x87 & ~x111 & ~x128 & ~x137 & ~x138 & ~x141 & ~x142 & ~x155 & ~x166 & ~x167 & ~x195 & ~x254 & ~x279 & ~x281 & ~x334 & ~x359 & ~x363 & ~x384 & ~x385 & ~x417 & ~x440 & ~x447 & ~x448 & ~x465 & ~x477 & ~x525 & ~x526 & ~x555 & ~x560 & ~x611 & ~x613 & ~x642 & ~x759;
assign c2174 =  x312 & ~x204 & ~x617 & ~x620 & ~x758;
assign c2176 =  x342 & ~x1 & ~x3 & ~x28 & ~x29 & ~x30 & ~x31 & ~x56 & ~x58 & ~x60 & ~x61 & ~x76 & ~x80 & ~x86 & ~x89 & ~x104 & ~x105 & ~x107 & ~x116 & ~x132 & ~x133 & ~x135 & ~x137 & ~x138 & ~x139 & ~x141 & ~x142 & ~x143 & ~x145 & ~x161 & ~x162 & ~x164 & ~x166 & ~x167 & ~x169 & ~x170 & ~x171 & ~x192 & ~x194 & ~x196 & ~x198 & ~x223 & ~x225 & ~x226 & ~x250 & ~x251 & ~x307 & ~x309 & ~x364 & ~x391 & ~x392 & ~x393 & ~x418 & ~x421 & ~x422 & ~x447 & ~x449 & ~x450 & ~x473 & ~x475 & ~x476 & ~x478 & ~x497 & ~x499 & ~x500 & ~x502 & ~x503 & ~x506 & ~x530 & ~x531 & ~x533 & ~x551 & ~x552 & ~x555 & ~x556 & ~x557 & ~x581 & ~x582 & ~x583 & ~x585 & ~x611 & ~x612 & ~x613 & ~x614 & ~x616 & ~x637 & ~x639 & ~x641 & ~x643 & ~x644 & ~x645 & ~x647 & ~x648 & ~x666 & ~x669 & ~x670 & ~x671 & ~x678 & ~x696 & ~x697 & ~x700 & ~x701 & ~x702 & ~x703 & ~x704 & ~x705 & ~x707 & ~x728 & ~x729 & ~x731 & ~x733 & ~x753 & ~x756 & ~x757 & ~x758 & ~x760 & ~x761 & ~x766 & ~x783;
assign c2178 =  x155 &  x156 & ~x24 & ~x25 & ~x29 & ~x31 & ~x52 & ~x53 & ~x59 & ~x84 & ~x111 & ~x113 & ~x197 & ~x216 & ~x218 & ~x221 & ~x222 & ~x227 & ~x235 & ~x236 & ~x242 & ~x243 & ~x245 & ~x253 & ~x254 & ~x259 & ~x270 & ~x272 & ~x298 & ~x306 & ~x308 & ~x310 & ~x336 & ~x338 & ~x362 & ~x363 & ~x394 & ~x446 & ~x447 & ~x449 & ~x502 & ~x534 & ~x582 & ~x585 & ~x613 & ~x637 & ~x669 & ~x671 & ~x697 & ~x730 & ~x760;
assign c2180 = ~x12 & ~x38 & ~x83 & ~x93 & ~x109 & ~x140 & ~x359 & ~x375 & ~x386 & ~x390 & ~x411 & ~x412 & ~x417 & ~x427 & ~x454 & ~x473 & ~x501 & ~x502 & ~x529 & ~x535 & ~x662 & ~x671 & ~x690 & ~x719 & ~x722 & ~x753;
assign c2182 =  x412 & ~x24 & ~x26 & ~x55 & ~x58 & ~x84 & ~x85 & ~x113 & ~x138 & ~x168 & ~x196 & ~x224 & ~x305 & ~x323 & ~x363 & ~x419 & ~x447 & ~x575 & ~x576 & ~x601 & ~x602 & ~x603 & ~x631 & ~x632 & ~x750 & ~x780;
assign c2184 =  x213 &  x214 & ~x140 & ~x152 & ~x374 & ~x375 & ~x447 & ~x481 & ~x482 & ~x505 & ~x531 & ~x532 & ~x535 & ~x562 & ~x585 & ~x613 & ~x622 & ~x643 & ~x649 & ~x699 & ~x724 & ~x731 & ~x734 & ~x756 & ~x761;
assign c2186 =  x124 &  x353 & ~x23 & ~x79 & ~x80 & ~x113 & ~x143 & ~x191 & ~x213 & ~x222 & ~x240 & ~x281 & ~x307 & ~x364 & ~x389 & ~x473 & ~x498 & ~x499 & ~x501 & ~x524 & ~x527 & ~x534 & ~x535 & ~x551 & ~x560 & ~x616 & ~x703 & ~x732 & ~x757;
assign c2188 =  x100 &  x127 &  x379 & ~x0 & ~x8 & ~x110 & ~x137 & ~x139 & ~x166 & ~x167 & ~x191 & ~x193 & ~x194 & ~x214 & ~x221 & ~x244 & ~x256 & ~x262 & ~x281 & ~x282 & ~x337 & ~x363 & ~x392 & ~x669 & ~x699 & ~x700 & ~x725 & ~x753 & ~x754;
assign c2190 =  x243 & ~x179 & ~x376 & ~x428 & ~x509 & ~x511;
assign c2192 =  x379 &  x406 & ~x3 & ~x27 & ~x57 & ~x60 & ~x80 & ~x81 & ~x83 & ~x84 & ~x85 & ~x87 & ~x110 & ~x113 & ~x116 & ~x136 & ~x137 & ~x138 & ~x139 & ~x141 & ~x143 & ~x144 & ~x157 & ~x172 & ~x184 & ~x196 & ~x198 & ~x199 & ~x224 & ~x251 & ~x254 & ~x281 & ~x282 & ~x305 & ~x336 & ~x360 & ~x362 & ~x390 & ~x415 & ~x419 & ~x447 & ~x471 & ~x491 & ~x492 & ~x500 & ~x519 & ~x529 & ~x531 & ~x699 & ~x700 & ~x728 & ~x729 & ~x755 & ~x756 & ~x757 & ~x758;
assign c2194 =  x618 & ~x537;
assign c2196 =  x478 & ~x463;
assign c2198 =  x156 &  x204 & ~x112 & ~x273 & ~x301 & ~x318 & ~x450 & ~x451 & ~x528 & ~x561 & ~x582 & ~x610 & ~x674 & ~x677 & ~x729;
assign c2200 =  x298 &  x551 & ~x5 & ~x391 & ~x419 & ~x428 & ~x482 & ~x700 & ~x712 & ~x739 & ~x741 & ~x754;
assign c2202 = ~x8 & ~x45 & ~x50 & ~x58 & ~x74 & ~x77 & ~x82 & ~x102 & ~x103 & ~x131 & ~x143 & ~x174 & ~x192 & ~x202 & ~x213 & ~x218 & ~x225 & ~x230 & ~x241 & ~x255 & ~x268 & ~x269 & ~x296 & ~x306 & ~x309 & ~x334 & ~x338 & ~x361 & ~x363 & ~x420 & ~x447 & ~x474 & ~x499 & ~x528 & ~x578 & ~x579 & ~x580 & ~x581 & ~x584 & ~x636 & ~x642 & ~x643 & ~x651 & ~x652 & ~x653 & ~x664 & ~x667 & ~x692 & ~x693 & ~x696 & ~x707 & ~x724 & ~x727 & ~x756 & ~x760;
assign c2204 = ~x1 & ~x56 & ~x85 & ~x136 & ~x194 & ~x225 & ~x243 & ~x269 & ~x276 & ~x296 & ~x310 & ~x323 & ~x357 & ~x363 & ~x385 & ~x386 & ~x387 & ~x452 & ~x564 & ~x579 & ~x604 & ~x608 & ~x662 & ~x667 & ~x719 & ~x747 & ~x754 & ~x755;
assign c2206 =  x231 &  x432 & ~x60 & ~x61 & ~x82 & ~x85 & ~x107 & ~x116 & ~x222 & ~x249 & ~x250 & ~x303 & ~x312 & ~x333 & ~x357 & ~x358 & ~x384 & ~x385 & ~x413 & ~x414 & ~x451 & ~x501 & ~x558 & ~x563 & ~x620 & ~x642 & ~x648 & ~x676 & ~x732;
assign c2208 =  x155 & ~x0 & ~x1 & ~x5 & ~x24 & ~x25 & ~x26 & ~x27 & ~x36 & ~x49 & ~x54 & ~x57 & ~x80 & ~x81 & ~x109 & ~x110 & ~x113 & ~x165 & ~x167 & ~x168 & ~x171 & ~x194 & ~x196 & ~x197 & ~x216 & ~x221 & ~x222 & ~x223 & ~x227 & ~x236 & ~x242 & ~x243 & ~x244 & ~x245 & ~x248 & ~x250 & ~x251 & ~x252 & ~x273 & ~x275 & ~x276 & ~x277 & ~x279 & ~x280 & ~x284 & ~x303 & ~x304 & ~x310 & ~x311 & ~x337 & ~x362 & ~x365 & ~x366 & ~x367 & ~x389 & ~x391 & ~x392 & ~x393 & ~x394 & ~x395 & ~x420 & ~x449 & ~x450 & ~x471 & ~x472 & ~x473 & ~x474 & ~x475 & ~x476 & ~x478 & ~x479 & ~x499 & ~x503 & ~x505 & ~x526 & ~x529 & ~x530 & ~x534 & ~x535 & ~x552 & ~x554 & ~x560 & ~x579 & ~x580 & ~x583 & ~x584 & ~x588 & ~x589 & ~x606 & ~x607 & ~x608 & ~x613 & ~x614 & ~x615 & ~x617 & ~x634 & ~x635 & ~x638 & ~x639 & ~x642 & ~x643 & ~x646 & ~x662 & ~x671 & ~x672 & ~x697 & ~x698 & ~x699 & ~x701 & ~x703 & ~x705 & ~x707 & ~x724 & ~x725 & ~x726 & ~x727 & ~x729 & ~x730 & ~x733 & ~x734 & ~x752 & ~x753 & ~x754 & ~x755 & ~x760 & ~x761 & ~x781;
assign c2210 = ~x5 & ~x24 & ~x25 & ~x54 & ~x153 & ~x349 & ~x374 & ~x387 & ~x388 & ~x389 & ~x401 & ~x416 & ~x426 & ~x427 & ~x428 & ~x446 & ~x455 & ~x480 & ~x481 & ~x483 & ~x500 & ~x505 & ~x507 & ~x510 & ~x528 & ~x530 & ~x537 & ~x556 & ~x559 & ~x561 & ~x564 & ~x565 & ~x590 & ~x594 & ~x616 & ~x622 & ~x623 & ~x640 & ~x641 & ~x646 & ~x654 & ~x668 & ~x674 & ~x675 & ~x704 & ~x758 & ~x761;
assign c2212 =  x99 &  x239 & ~x207 & ~x224 & ~x233 & ~x419 & ~x529 & ~x588 & ~x682 & ~x692 & ~x734 & ~x782;
assign c2214 = ~x10 & ~x26 & ~x29 & ~x52 & ~x54 & ~x110 & ~x166 & ~x249 & ~x280 & ~x356 & ~x412 & ~x421 & ~x447 & ~x454 & ~x466 & ~x467 & ~x482 & ~x497 & ~x522 & ~x523 & ~x526 & ~x531 & ~x534 & ~x538 & ~x550 & ~x554 & ~x567 & ~x578 & ~x582 & ~x590 & ~x593 & ~x613 & ~x623 & ~x645 & ~x652 & ~x690 & ~x697 & ~x699 & ~x703 & ~x716 & ~x732 & ~x734 & ~x746 & ~x754 & ~x756 & ~x757 & ~x780;
assign c2216 =  x468 & ~x0 & ~x1 & ~x4 & ~x28 & ~x55 & ~x58 & ~x60 & ~x168 & ~x261 & ~x263 & ~x474 & ~x559 & ~x645 & ~x672 & ~x698 & ~x704 & ~x727 & ~x729 & ~x737 & ~x754 & ~x760 & ~x763;
assign c2218 =  x133 & ~x5 & ~x277 & ~x346 & ~x428 & ~x700 & ~x702 & ~x728;
assign c2220 =  x353 &  x379 & ~x81 & ~x82 & ~x84 & ~x115 & ~x159 & ~x169 & ~x170 & ~x187 & ~x194 & ~x196 & ~x214 & ~x221 & ~x227 & ~x239 & ~x240 & ~x267 & ~x278 & ~x305 & ~x309 & ~x333 & ~x335 & ~x390 & ~x391 & ~x442 & ~x445 & ~x468 & ~x471 & ~x497 & ~x498 & ~x500 & ~x533 & ~x555 & ~x556 & ~x557 & ~x560 & ~x581 & ~x585 & ~x587 & ~x588 & ~x643 & ~x669 & ~x672 & ~x674 & ~x755 & ~x757 & ~x781;
assign c2222 =  x370 &  x398 & ~x1 & ~x2 & ~x3 & ~x22 & ~x23 & ~x26 & ~x31 & ~x49 & ~x51 & ~x52 & ~x53 & ~x58 & ~x79 & ~x81 & ~x85 & ~x87 & ~x110 & ~x113 & ~x114 & ~x115 & ~x136 & ~x137 & ~x138 & ~x143 & ~x169 & ~x193 & ~x198 & ~x199 & ~x223 & ~x225 & ~x248 & ~x249 & ~x252 & ~x253 & ~x280 & ~x282 & ~x283 & ~x306 & ~x307 & ~x309 & ~x338 & ~x364 & ~x389 & ~x392 & ~x394 & ~x448 & ~x449 & ~x473 & ~x498 & ~x503 & ~x504 & ~x505 & ~x528 & ~x529 & ~x530 & ~x560 & ~x561 & ~x575 & ~x586 & ~x589 & ~x602 & ~x603 & ~x614 & ~x644 & ~x670 & ~x673 & ~x700 & ~x726 & ~x728 & ~x729 & ~x730 & ~x759;
assign c2224 = ~x24 & ~x27 & ~x82 & ~x85 & ~x112 & ~x250 & ~x274 & ~x303 & ~x305 & ~x331 & ~x332 & ~x333 & ~x336 & ~x344 & ~x387 & ~x399 & ~x401 & ~x427 & ~x447 & ~x455 & ~x472 & ~x473 & ~x484 & ~x501 & ~x511 & ~x558 & ~x561 & ~x585 & ~x586 & ~x600 & ~x601 & ~x641 & ~x642 & ~x644 & ~x645 & ~x656 & ~x672 & ~x684 & ~x699 & ~x701 & ~x711 & ~x730 & ~x754 & ~x755 & ~x756;
assign c2226 =  x618 & ~x317 & ~x399 & ~x454 & ~x602;
assign c2228 =  x631 & ~x28 & ~x54 & ~x110 & ~x117 & ~x181 & ~x195 & ~x197 & ~x206 & ~x496 & ~x512 & ~x638 & ~x655 & ~x681 & ~x694;
assign c2230 =  x412 & ~x0 & ~x55 & ~x58 & ~x87 & ~x111 & ~x250 & ~x305 & ~x306 & ~x333 & ~x445 & ~x446 & ~x491 & ~x547 & ~x548 & ~x577 & ~x601 & ~x602 & ~x749 & ~x750;
assign c2232 =  x297 & ~x32 & ~x128 & ~x130 & ~x211 & ~x359 & ~x415 & ~x490 & ~x756;
assign c2234 =  x533;
assign c2236 =  x128 &  x155 &  x183 &  x323 & ~x8 & ~x53 & ~x59 & ~x63 & ~x109 & ~x167 & ~x298 & ~x326 & ~x360 & ~x450 & ~x530 & ~x561 & ~x583 & ~x585 & ~x614 & ~x664 & ~x671 & ~x692 & ~x694 & ~x698 & ~x706 & ~x726 & ~x731 & ~x734 & ~x783;
assign c2238 =  x477;
assign c2240 =  x292 &  x316 & ~x54 & ~x82 & ~x107 & ~x135 & ~x137 & ~x138 & ~x140 & ~x143 & ~x170 & ~x386 & ~x391 & ~x416 & ~x420 & ~x447 & ~x472 & ~x480 & ~x504 & ~x530 & ~x582 & ~x583 & ~x592 & ~x639 & ~x644 & ~x647 & ~x672 & ~x694 & ~x702 & ~x703 & ~x724 & ~x725 & ~x726 & ~x736 & ~x738 & ~x781;
assign c2242 =  x368 & ~x173 & ~x200 & ~x529 & ~x556 & ~x558 & ~x583 & ~x618 & ~x704;
assign c2244 =  x216 & ~x0 & ~x3 & ~x27 & ~x29 & ~x125 & ~x153 & ~x390 & ~x417 & ~x428 & ~x455 & ~x482 & ~x538 & ~x566 & ~x593;
assign c2246 = ~x23 & ~x24 & ~x28 & ~x29 & ~x70 & ~x97 & ~x98 & ~x223 & ~x251 & ~x279 & ~x280 & ~x351 & ~x352 & ~x360 & ~x362 & ~x372 & ~x379 & ~x380 & ~x390 & ~x407 & ~x419 & ~x434 & ~x725 & ~x727 & ~x782;
assign c2248 =  x434 &  x461 & ~x0 & ~x1 & ~x3 & ~x24 & ~x28 & ~x32 & ~x53 & ~x54 & ~x57 & ~x59 & ~x80 & ~x81 & ~x84 & ~x88 & ~x89 & ~x114 & ~x116 & ~x138 & ~x143 & ~x164 & ~x165 & ~x166 & ~x167 & ~x169 & ~x170 & ~x191 & ~x194 & ~x196 & ~x198 & ~x218 & ~x219 & ~x220 & ~x222 & ~x224 & ~x225 & ~x243 & ~x248 & ~x254 & ~x269 & ~x275 & ~x278 & ~x280 & ~x305 & ~x307 & ~x309 & ~x334 & ~x335 & ~x338 & ~x366 & ~x392 & ~x393 & ~x418 & ~x422 & ~x449 & ~x473 & ~x474 & ~x493 & ~x500 & ~x502 & ~x505 & ~x520 & ~x525 & ~x529 & ~x533 & ~x547 & ~x550 & ~x552 & ~x553 & ~x556 & ~x557 & ~x558 & ~x561 & ~x577 & ~x578 & ~x586 & ~x606 & ~x614 & ~x615 & ~x616 & ~x639 & ~x640 & ~x641 & ~x642 & ~x643 & ~x644 & ~x647 & ~x651 & ~x670 & ~x671 & ~x672 & ~x674 & ~x679 & ~x700 & ~x726 & ~x728 & ~x729 & ~x730 & ~x731 & ~x735 & ~x753 & ~x754 & ~x756 & ~x757 & ~x758 & ~x759 & ~x760 & ~x761 & ~x781;
assign c2250 = ~x0 & ~x1 & ~x26 & ~x29 & ~x112 & ~x204 & ~x206 & ~x208 & ~x256 & ~x390 & ~x418 & ~x474 & ~x500 & ~x501 & ~x505 & ~x507 & ~x534 & ~x563 & ~x583 & ~x627 & ~x640 & ~x653 & ~x654 & ~x675 & ~x680 & ~x682 & ~x684 & ~x693 & ~x696 & ~x708 & ~x710 & ~x711 & ~x722 & ~x724 & ~x733 & ~x734 & ~x766;
assign c2252 =  x232 & ~x9 & ~x33 & ~x35 & ~x113 & ~x139 & ~x146 & ~x167 & ~x318 & ~x346 & ~x418 & ~x420 & ~x475 & ~x506 & ~x534 & ~x584 & ~x586 & ~x589 & ~x611 & ~x674 & ~x701 & ~x781;
assign c2254 = ~x7 & ~x24 & ~x109 & ~x141 & ~x166 & ~x170 & ~x195 & ~x225 & ~x299 & ~x329 & ~x333 & ~x339 & ~x365 & ~x366 & ~x370 & ~x384 & ~x390 & ~x396 & ~x400 & ~x411 & ~x412 & ~x439 & ~x445 & ~x449 & ~x451 & ~x453 & ~x455 & ~x457 & ~x467 & ~x477 & ~x496 & ~x522 & ~x527 & ~x529 & ~x533 & ~x550 & ~x553 & ~x555 & ~x556 & ~x564 & ~x570 & ~x578 & ~x580 & ~x583 & ~x590 & ~x613 & ~x619 & ~x621 & ~x626 & ~x637 & ~x642 & ~x647 & ~x650 & ~x663 & ~x666 & ~x678 & ~x690 & ~x700 & ~x723 & ~x727 & ~x729 & ~x730 & ~x752;
assign c2256 =  x99 &  x408 & ~x3 & ~x24 & ~x52 & ~x111 & ~x168 & ~x418 & ~x526 & ~x531 & ~x551 & ~x553 & ~x554 & ~x556 & ~x562 & ~x585 & ~x595 & ~x597 & ~x611 & ~x617 & ~x623 & ~x640 & ~x646 & ~x650 & ~x652 & ~x668 & ~x698 & ~x700 & ~x704 & ~x705 & ~x712 & ~x725 & ~x738;
assign c2258 =  x181 & ~x54 & ~x114 & ~x137 & ~x141 & ~x143 & ~x242 & ~x298 & ~x363 & ~x392 & ~x419 & ~x497 & ~x523 & ~x563 & ~x578 & ~x632 & ~x641 & ~x662 & ~x692 & ~x719 & ~x755;
assign c2260 =  x455 & ~x6 & ~x55 & ~x79 & ~x81 & ~x106 & ~x108 & ~x132 & ~x134 & ~x160 & ~x170 & ~x198 & ~x216 & ~x228 & ~x245 & ~x253 & ~x255 & ~x269 & ~x270 & ~x277 & ~x278 & ~x447 & ~x506 & ~x562 & ~x589 & ~x590 & ~x607 & ~x610 & ~x635 & ~x636 & ~x640 & ~x665 & ~x666 & ~x696 & ~x697 & ~x699 & ~x725 & ~x728;
assign c2262 =  x713 &  x741 & ~x0 & ~x30 & ~x59 & ~x113 & ~x132 & ~x159 & ~x160 & ~x171 & ~x193 & ~x199 & ~x220 & ~x246 & ~x248 & ~x268 & ~x338 & ~x552 & ~x556 & ~x558 & ~x584 & ~x588 & ~x611 & ~x630 & ~x636 & ~x672 & ~x707 & ~x728 & ~x734 & ~x761 & ~x762 & ~x765;
assign c2264 = ~x1 & ~x8 & ~x26 & ~x30 & ~x31 & ~x35 & ~x53 & ~x59 & ~x61 & ~x81 & ~x87 & ~x109 & ~x114 & ~x117 & ~x138 & ~x140 & ~x142 & ~x169 & ~x173 & ~x174 & ~x186 & ~x193 & ~x198 & ~x199 & ~x201 & ~x202 & ~x225 & ~x251 & ~x252 & ~x254 & ~x255 & ~x277 & ~x281 & ~x283 & ~x308 & ~x309 & ~x311 & ~x332 & ~x333 & ~x360 & ~x364 & ~x389 & ~x390 & ~x391 & ~x418 & ~x455 & ~x474 & ~x500 & ~x501 & ~x502 & ~x527 & ~x530 & ~x587 & ~x655 & ~x656 & ~x684 & ~x711 & ~x737 & ~x739 & ~x765 & ~x782;
assign c2266 = ~x9 & ~x24 & ~x27 & ~x29 & ~x30 & ~x55 & ~x57 & ~x83 & ~x84 & ~x85 & ~x113 & ~x139 & ~x140 & ~x169 & ~x195 & ~x224 & ~x270 & ~x280 & ~x291 & ~x292 & ~x300 & ~x303 & ~x317 & ~x329 & ~x332 & ~x336 & ~x357 & ~x361 & ~x362 & ~x364 & ~x366 & ~x367 & ~x368 & ~x369 & ~x384 & ~x389 & ~x390 & ~x391 & ~x394 & ~x396 & ~x414 & ~x415 & ~x416 & ~x418 & ~x419 & ~x420 & ~x421 & ~x424 & ~x443 & ~x444 & ~x449 & ~x450 & ~x451 & ~x452 & ~x453 & ~x473 & ~x474 & ~x478 & ~x479 & ~x481 & ~x498 & ~x499 & ~x507 & ~x508 & ~x509 & ~x525 & ~x526 & ~x527 & ~x530 & ~x531 & ~x533 & ~x534 & ~x535 & ~x536 & ~x539 & ~x552 & ~x554 & ~x556 & ~x558 & ~x561 & ~x563 & ~x567 & ~x583 & ~x588 & ~x591 & ~x610 & ~x612 & ~x613 & ~x615 & ~x616 & ~x619 & ~x620 & ~x621 & ~x622 & ~x623 & ~x624 & ~x636 & ~x640 & ~x641 & ~x642 & ~x643 & ~x644 & ~x645 & ~x647 & ~x648 & ~x651 & ~x652 & ~x667 & ~x668 & ~x669 & ~x670 & ~x671 & ~x673 & ~x674 & ~x678 & ~x695 & ~x697 & ~x700 & ~x701 & ~x702 & ~x723 & ~x733 & ~x734 & ~x752 & ~x753 & ~x756 & ~x757 & ~x758 & ~x759 & ~x760 & ~x781;
assign c2268 = ~x0 & ~x2 & ~x6 & ~x27 & ~x28 & ~x29 & ~x31 & ~x33 & ~x45 & ~x51 & ~x53 & ~x54 & ~x56 & ~x58 & ~x72 & ~x78 & ~x81 & ~x85 & ~x88 & ~x89 & ~x107 & ~x110 & ~x114 & ~x116 & ~x133 & ~x138 & ~x164 & ~x165 & ~x167 & ~x169 & ~x188 & ~x190 & ~x191 & ~x193 & ~x228 & ~x246 & ~x248 & ~x250 & ~x253 & ~x278 & ~x279 & ~x282 & ~x303 & ~x304 & ~x306 & ~x309 & ~x311 & ~x330 & ~x331 & ~x333 & ~x334 & ~x335 & ~x339 & ~x357 & ~x359 & ~x362 & ~x366 & ~x388 & ~x390 & ~x393 & ~x396 & ~x415 & ~x417 & ~x419 & ~x423 & ~x442 & ~x443 & ~x444 & ~x445 & ~x448 & ~x449 & ~x471 & ~x475 & ~x477 & ~x529 & ~x530 & ~x532 & ~x533 & ~x534 & ~x558 & ~x562 & ~x587 & ~x589 & ~x590 & ~x617 & ~x630 & ~x643 & ~x644 & ~x658 & ~x668 & ~x670 & ~x673 & ~x674 & ~x698 & ~x702 & ~x723 & ~x728 & ~x752 & ~x754 & ~x760 & ~x768;
assign c2270 =  x551 & ~x25 & ~x57 & ~x125 & ~x361 & ~x373 & ~x399 & ~x400 & ~x417 & ~x419 & ~x427 & ~x482 & ~x768;
assign c2272 = ~x20 & ~x21 & ~x55 & ~x59 & ~x86 & ~x87 & ~x112 & ~x121 & ~x122 & ~x149 & ~x174 & ~x176 & ~x202 & ~x203 & ~x389 & ~x390 & ~x404 & ~x418 & ~x452 & ~x514 & ~x541 & ~x672 & ~x681 & ~x708 & ~x709 & ~x733 & ~x735 & ~x758 & ~x778 & ~x782;
assign c2274 =  x421;
assign c2276 =  x413 &  x563 & ~x577;
assign c2278 =  x182 & ~x27 & ~x28 & ~x60 & ~x88 & ~x104 & ~x140 & ~x142 & ~x144 & ~x189 & ~x214 & ~x218 & ~x221 & ~x254 & ~x422 & ~x500 & ~x537 & ~x558 & ~x608 & ~x622 & ~x648 & ~x654 & ~x655 & ~x667 & ~x668 & ~x669 & ~x700 & ~x748 & ~x754 & ~x780;
assign c2280 =  x327 & ~x109 & ~x204 & ~x205 & ~x231 & ~x445 & ~x740 & ~x741;
assign c2282 =  x293 &  x317 & ~x0 & ~x28 & ~x29 & ~x30 & ~x50 & ~x53 & ~x59 & ~x79 & ~x82 & ~x88 & ~x89 & ~x90 & ~x114 & ~x115 & ~x117 & ~x119 & ~x135 & ~x138 & ~x141 & ~x146 & ~x162 & ~x165 & ~x174 & ~x200 & ~x252 & ~x253 & ~x363 & ~x390 & ~x393 & ~x444 & ~x445 & ~x446 & ~x448 & ~x449 & ~x472 & ~x497 & ~x500 & ~x502 & ~x505 & ~x508 & ~x525 & ~x526 & ~x533 & ~x534 & ~x553 & ~x562 & ~x584 & ~x585 & ~x588 & ~x590 & ~x591 & ~x593 & ~x611 & ~x612 & ~x616 & ~x618 & ~x621 & ~x641 & ~x647 & ~x650 & ~x651 & ~x670 & ~x674 & ~x677 & ~x678 & ~x693 & ~x701 & ~x721 & ~x722 & ~x724 & ~x756 & ~x757 & ~x759 & ~x762 & ~x779 & ~x782;
assign c2284 =  x125 &  x153 &  x181 &  x209 &  x237 &  x265 &  x293 & ~x22 & ~x23 & ~x24 & ~x25 & ~x27 & ~x51 & ~x53 & ~x55 & ~x56 & ~x74 & ~x75 & ~x76 & ~x80 & ~x81 & ~x85 & ~x104 & ~x108 & ~x109 & ~x113 & ~x115 & ~x116 & ~x140 & ~x142 & ~x162 & ~x163 & ~x164 & ~x165 & ~x166 & ~x167 & ~x168 & ~x170 & ~x171 & ~x191 & ~x198 & ~x222 & ~x224 & ~x269 & ~x363 & ~x392 & ~x448 & ~x475 & ~x476 & ~x503 & ~x504 & ~x527 & ~x529 & ~x531 & ~x552 & ~x553 & ~x554 & ~x555 & ~x556 & ~x579 & ~x580 & ~x582 & ~x584 & ~x586 & ~x588 & ~x606 & ~x609 & ~x611 & ~x613 & ~x616 & ~x633 & ~x638 & ~x643 & ~x667 & ~x671 & ~x696 & ~x697 & ~x700 & ~x701 & ~x702 & ~x703 & ~x705 & ~x728 & ~x731 & ~x732 & ~x735 & ~x751 & ~x752 & ~x755 & ~x756 & ~x758 & ~x762 & ~x780 & ~x781 & ~x783;
assign c2286 =  x438 &  x464 &  x491 &  x517 &  x544 & ~x30 & ~x114 & ~x134 & ~x137 & ~x141 & ~x270 & ~x391 & ~x579 & ~x607 & ~x608 & ~x612 & ~x639 & ~x668 & ~x731 & ~x734;
assign c2288 = ~x139 & ~x274 & ~x279 & ~x292 & ~x293 & ~x306 & ~x330 & ~x336 & ~x337 & ~x369 & ~x370 & ~x373 & ~x386 & ~x388 & ~x417 & ~x423 & ~x426 & ~x427 & ~x446 & ~x449 & ~x452 & ~x455 & ~x479 & ~x481 & ~x483 & ~x499 & ~x504 & ~x511 & ~x527 & ~x538 & ~x558 & ~x562 & ~x563 & ~x567 & ~x586 & ~x587 & ~x591 & ~x620 & ~x622 & ~x623 & ~x624 & ~x626 & ~x638 & ~x640 & ~x643 & ~x645 & ~x652 & ~x653 & ~x678 & ~x694 & ~x701 & ~x707 & ~x725 & ~x726 & ~x751 & ~x756 & ~x757 & ~x782;
assign c2290 =  x515 & ~x24 & ~x49 & ~x82 & ~x104 & ~x128 & ~x136 & ~x141 & ~x155 & ~x166 & ~x173 & ~x195 & ~x251 & ~x266 & ~x280 & ~x305 & ~x306 & ~x414 & ~x417 & ~x533 & ~x554 & ~x584 & ~x588 & ~x620 & ~x666 & ~x672 & ~x756;
assign c2292 =  x182 & ~x3 & ~x4 & ~x24 & ~x27 & ~x28 & ~x33 & ~x45 & ~x48 & ~x51 & ~x57 & ~x59 & ~x60 & ~x76 & ~x77 & ~x83 & ~x85 & ~x86 & ~x87 & ~x106 & ~x107 & ~x110 & ~x112 & ~x114 & ~x116 & ~x138 & ~x140 & ~x143 & ~x165 & ~x167 & ~x170 & ~x171 & ~x191 & ~x192 & ~x194 & ~x195 & ~x197 & ~x219 & ~x221 & ~x223 & ~x224 & ~x225 & ~x226 & ~x227 & ~x249 & ~x250 & ~x270 & ~x276 & ~x278 & ~x279 & ~x282 & ~x283 & ~x299 & ~x302 & ~x305 & ~x310 & ~x327 & ~x332 & ~x334 & ~x335 & ~x337 & ~x338 & ~x352 & ~x353 & ~x361 & ~x364 & ~x366 & ~x390 & ~x421 & ~x422 & ~x446 & ~x447 & ~x476 & ~x477 & ~x531 & ~x532 & ~x555 & ~x556 & ~x557 & ~x558 & ~x560 & ~x580 & ~x581 & ~x583 & ~x588 & ~x613 & ~x616 & ~x633 & ~x634 & ~x645 & ~x661 & ~x664 & ~x670 & ~x671 & ~x692 & ~x695 & ~x697 & ~x698 & ~x700 & ~x723 & ~x727 & ~x753 & ~x757 & ~x781;
assign c2294 = ~x25 & ~x31 & ~x54 & ~x58 & ~x62 & ~x73 & ~x75 & ~x79 & ~x86 & ~x111 & ~x128 & ~x132 & ~x156 & ~x157 & ~x189 & ~x199 & ~x239 & ~x253 & ~x277 & ~x311 & ~x383 & ~x385 & ~x387 & ~x390 & ~x447 & ~x474 & ~x501 & ~x505 & ~x549 & ~x552 & ~x610 & ~x621 & ~x665 & ~x668 & ~x693 & ~x701 & ~x703 & ~x704 & ~x707 & ~x726 & ~x756 & ~x779;
assign c2296 = ~x30 & ~x33 & ~x35 & ~x55 & ~x57 & ~x93 & ~x223 & ~x359 & ~x387 & ~x390 & ~x416 & ~x428 & ~x429 & ~x447 & ~x455 & ~x457 & ~x472 & ~x483 & ~x511 & ~x514 & ~x534 & ~x537 & ~x538 & ~x542 & ~x543 & ~x558 & ~x592 & ~x614 & ~x615 & ~x627 & ~x628 & ~x654 & ~x670 & ~x699 & ~x711 & ~x733 & ~x757 & ~x759 & ~x765;
assign c2298 =  x374 & ~x2 & ~x28 & ~x53 & ~x60 & ~x84 & ~x85 & ~x106 & ~x107 & ~x111 & ~x113 & ~x116 & ~x141 & ~x165 & ~x168 & ~x171 & ~x192 & ~x195 & ~x198 & ~x227 & ~x228 & ~x250 & ~x278 & ~x279 & ~x306 & ~x332 & ~x356 & ~x362 & ~x363 & ~x382 & ~x383 & ~x384 & ~x385 & ~x387 & ~x417 & ~x441 & ~x470 & ~x471 & ~x476 & ~x498 & ~x503 & ~x527 & ~x529 & ~x535 & ~x554 & ~x555 & ~x556 & ~x558 & ~x562 & ~x582 & ~x586 & ~x590 & ~x592 & ~x606 & ~x608 & ~x610 & ~x612 & ~x620 & ~x633 & ~x642 & ~x645 & ~x646 & ~x649 & ~x663 & ~x670 & ~x673 & ~x674 & ~x676 & ~x698 & ~x700 & ~x718 & ~x721 & ~x724 & ~x725 & ~x727 & ~x728 & ~x756 & ~x758;
assign c2300 =  x125 &  x237 &  x265 &  x293 &  x321 & ~x0 & ~x1 & ~x3 & ~x25 & ~x29 & ~x50 & ~x53 & ~x54 & ~x55 & ~x78 & ~x79 & ~x81 & ~x82 & ~x84 & ~x86 & ~x107 & ~x108 & ~x110 & ~x116 & ~x133 & ~x136 & ~x137 & ~x139 & ~x140 & ~x141 & ~x142 & ~x143 & ~x145 & ~x162 & ~x164 & ~x166 & ~x167 & ~x169 & ~x172 & ~x193 & ~x194 & ~x195 & ~x196 & ~x198 & ~x221 & ~x223 & ~x227 & ~x228 & ~x243 & ~x246 & ~x247 & ~x248 & ~x250 & ~x251 & ~x255 & ~x268 & ~x277 & ~x279 & ~x282 & ~x283 & ~x296 & ~x297 & ~x306 & ~x312 & ~x337 & ~x338 & ~x393 & ~x419 & ~x420 & ~x421 & ~x502 & ~x503 & ~x505 & ~x531 & ~x533 & ~x556 & ~x579 & ~x580 & ~x581 & ~x584 & ~x586 & ~x587 & ~x608 & ~x610 & ~x611 & ~x612 & ~x613 & ~x614 & ~x638 & ~x640 & ~x642 & ~x667 & ~x668 & ~x669 & ~x670 & ~x696 & ~x698 & ~x699 & ~x701 & ~x724 & ~x728 & ~x729 & ~x756 & ~x758 & ~x781;
assign c2302 =  x401 & ~x137 & ~x159 & ~x217 & ~x220 & ~x578 & ~x587 & ~x603 & ~x608 & ~x611 & ~x633 & ~x634 & ~x646 & ~x736 & ~x753;
assign c2304 = ~x112 & ~x279 & ~x390 & ~x419 & ~x429 & ~x445 & ~x451 & ~x453 & ~x458 & ~x484 & ~x564 & ~x566 & ~x567 & ~x572 & ~x587 & ~x589 & ~x600 & ~x617 & ~x624 & ~x628 & ~x675 & ~x679 & ~x683 & ~x722 & ~x735 & ~x751;
assign c2306 =  x453 & ~x0 & ~x4 & ~x5 & ~x17 & ~x20 & ~x27 & ~x29 & ~x46 & ~x49 & ~x54 & ~x61 & ~x79 & ~x85 & ~x87 & ~x88 & ~x107 & ~x109 & ~x112 & ~x116 & ~x134 & ~x138 & ~x140 & ~x141 & ~x144 & ~x163 & ~x164 & ~x165 & ~x168 & ~x169 & ~x170 & ~x191 & ~x192 & ~x193 & ~x194 & ~x195 & ~x196 & ~x198 & ~x199 & ~x221 & ~x223 & ~x224 & ~x226 & ~x248 & ~x249 & ~x250 & ~x252 & ~x254 & ~x280 & ~x281 & ~x309 & ~x334 & ~x336 & ~x419 & ~x476 & ~x502 & ~x505 & ~x525 & ~x526 & ~x529 & ~x530 & ~x532 & ~x533 & ~x555 & ~x557 & ~x584 & ~x585 & ~x586 & ~x588 & ~x614 & ~x615 & ~x616 & ~x641 & ~x643 & ~x699 & ~x702 & ~x726 & ~x727 & ~x728 & ~x730 & ~x754 & ~x755 & ~x782;
assign c2308 =  x259 & ~x8 & ~x61 & ~x87 & ~x170 & ~x171 & ~x305 & ~x329 & ~x373 & ~x441 & ~x442 & ~x527 & ~x589 & ~x640 & ~x672 & ~x731;
assign c2310 =  x212 & ~x58 & ~x299 & ~x319 & ~x327 & ~x342 & ~x346 & ~x355 & ~x359 & ~x371 & ~x383 & ~x384 & ~x388 & ~x391 & ~x394 & ~x395 & ~x399 & ~x415 & ~x416 & ~x418 & ~x420 & ~x421 & ~x423 & ~x424 & ~x443 & ~x444 & ~x447 & ~x453 & ~x454 & ~x476 & ~x477 & ~x500 & ~x504 & ~x506 & ~x509 & ~x510 & ~x529 & ~x530 & ~x532 & ~x534 & ~x536 & ~x556 & ~x561 & ~x565 & ~x583 & ~x588 & ~x590 & ~x591 & ~x611 & ~x616 & ~x617 & ~x620 & ~x622 & ~x643 & ~x645 & ~x648 & ~x669 & ~x675 & ~x705 & ~x728 & ~x732 & ~x758 & ~x759;
assign c2312 =  x514 & ~x0 & ~x57 & ~x60 & ~x80 & ~x116 & ~x135 & ~x143 & ~x144 & ~x162 & ~x163 & ~x168 & ~x186 & ~x188 & ~x199 & ~x213 & ~x216 & ~x223 & ~x226 & ~x240 & ~x246 & ~x249 & ~x252 & ~x307 & ~x308 & ~x338 & ~x392 & ~x446 & ~x447 & ~x524 & ~x525 & ~x528 & ~x532 & ~x550 & ~x552 & ~x554 & ~x583 & ~x588 & ~x616 & ~x623 & ~x639 & ~x676 & ~x678 & ~x698 & ~x699 & ~x705 & ~x707 & ~x725 & ~x726;
assign c2314 =  x212 & ~x28 & ~x82 & ~x152 & ~x328 & ~x330 & ~x331 & ~x346 & ~x357 & ~x359 & ~x362 & ~x363 & ~x372 & ~x398 & ~x414 & ~x440 & ~x451 & ~x468 & ~x473 & ~x476 & ~x478 & ~x504 & ~x561 & ~x642 & ~x670 & ~x693 & ~x720 & ~x756 & ~x758 & ~x759;
assign c2316 =  x152 &  x655 & ~x1 & ~x3 & ~x24 & ~x25 & ~x27 & ~x28 & ~x29 & ~x31 & ~x53 & ~x56 & ~x57 & ~x59 & ~x78 & ~x81 & ~x83 & ~x86 & ~x108 & ~x113 & ~x114 & ~x136 & ~x138 & ~x140 & ~x141 & ~x161 & ~x162 & ~x163 & ~x164 & ~x166 & ~x167 & ~x169 & ~x170 & ~x190 & ~x191 & ~x193 & ~x195 & ~x197 & ~x198 & ~x199 & ~x217 & ~x220 & ~x222 & ~x224 & ~x225 & ~x227 & ~x242 & ~x244 & ~x245 & ~x246 & ~x253 & ~x254 & ~x269 & ~x270 & ~x275 & ~x279 & ~x307 & ~x308 & ~x334 & ~x337 & ~x390 & ~x391 & ~x392 & ~x393 & ~x446 & ~x448 & ~x472 & ~x473 & ~x475 & ~x476 & ~x502 & ~x504 & ~x526 & ~x532 & ~x552 & ~x555 & ~x556 & ~x557 & ~x558 & ~x581 & ~x583 & ~x584 & ~x585 & ~x587 & ~x605 & ~x609 & ~x610 & ~x613 & ~x615 & ~x616 & ~x637 & ~x639 & ~x669 & ~x671 & ~x672 & ~x697 & ~x699 & ~x700 & ~x725 & ~x728 & ~x729 & ~x730 & ~x753 & ~x754 & ~x756 & ~x757 & ~x760;
assign c2318 =  x183 &  x294 &  x349 & ~x3 & ~x19 & ~x21 & ~x31 & ~x32 & ~x47 & ~x53 & ~x60 & ~x81 & ~x115 & ~x168 & ~x170 & ~x196 & ~x201 & ~x244 & ~x269 & ~x270 & ~x272 & ~x280 & ~x282 & ~x283 & ~x297 & ~x301 & ~x334 & ~x337 & ~x420 & ~x422 & ~x502 & ~x530 & ~x534 & ~x561 & ~x585 & ~x612 & ~x616 & ~x636 & ~x670 & ~x705 & ~x731 & ~x732 & ~x734 & ~x753 & ~x756 & ~x781 & ~x782;
assign c2320 =  x297 & ~x56 & ~x81 & ~x208 & ~x448 & ~x456 & ~x473 & ~x498 & ~x509 & ~x540 & ~x541 & ~x558 & ~x565 & ~x566 & ~x598 & ~x652 & ~x667 & ~x680 & ~x706 & ~x728 & ~x753;
assign c2322 = ~x180 & ~x376 & ~x400 & ~x401 & ~x428 & ~x451 & ~x452 & ~x456 & ~x484 & ~x506 & ~x508 & ~x512 & ~x534 & ~x564 & ~x567 & ~x591 & ~x614 & ~x624 & ~x672 & ~x674;
assign c2324 =  x130 & ~x3 & ~x4 & ~x31 & ~x52 & ~x55 & ~x70 & ~x96 & ~x97 & ~x273 & ~x302 & ~x336 & ~x357 & ~x358 & ~x360 & ~x385 & ~x386 & ~x387 & ~x475 & ~x503 & ~x532 & ~x560 & ~x561 & ~x644 & ~x672 & ~x698 & ~x727 & ~x750 & ~x755;
assign c2326 = ~x0 & ~x1 & ~x26 & ~x28 & ~x31 & ~x110 & ~x303 & ~x305 & ~x332 & ~x333 & ~x334 & ~x359 & ~x400 & ~x444 & ~x446 & ~x455 & ~x516 & ~x544 & ~x599 & ~x601 & ~x627 & ~x629 & ~x655 & ~x682 & ~x713 & ~x728 & ~x759 & ~x766;
assign c2328 =  x208 & ~x0 & ~x1 & ~x20 & ~x24 & ~x25 & ~x28 & ~x29 & ~x30 & ~x31 & ~x46 & ~x52 & ~x53 & ~x59 & ~x73 & ~x74 & ~x76 & ~x77 & ~x79 & ~x80 & ~x101 & ~x102 & ~x105 & ~x106 & ~x107 & ~x109 & ~x110 & ~x112 & ~x114 & ~x115 & ~x129 & ~x130 & ~x135 & ~x136 & ~x140 & ~x141 & ~x142 & ~x159 & ~x160 & ~x164 & ~x166 & ~x170 & ~x186 & ~x193 & ~x199 & ~x218 & ~x220 & ~x223 & ~x224 & ~x227 & ~x239 & ~x249 & ~x254 & ~x255 & ~x267 & ~x276 & ~x278 & ~x280 & ~x282 & ~x283 & ~x307 & ~x308 & ~x310 & ~x334 & ~x335 & ~x336 & ~x363 & ~x365 & ~x389 & ~x391 & ~x417 & ~x420 & ~x421 & ~x422 & ~x443 & ~x445 & ~x447 & ~x449 & ~x471 & ~x472 & ~x478 & ~x506 & ~x526 & ~x528 & ~x530 & ~x531 & ~x535 & ~x551 & ~x552 & ~x557 & ~x560 & ~x561 & ~x562 & ~x579 & ~x582 & ~x583 & ~x586 & ~x587 & ~x589 & ~x590 & ~x610 & ~x615 & ~x618 & ~x619 & ~x620 & ~x637 & ~x638 & ~x640 & ~x643 & ~x664 & ~x667 & ~x670 & ~x672 & ~x673 & ~x676 & ~x693 & ~x694 & ~x695 & ~x700 & ~x701 & ~x705 & ~x726 & ~x729 & ~x730 & ~x731 & ~x732 & ~x733 & ~x734 & ~x755 & ~x756 & ~x757 & ~x759 & ~x762 & ~x781 & ~x782 & ~x783;
assign c2330 =  x542 &  x597 & ~x24 & ~x26 & ~x28 & ~x30 & ~x31 & ~x50 & ~x53 & ~x54 & ~x57 & ~x79 & ~x83 & ~x84 & ~x110 & ~x112 & ~x115 & ~x136 & ~x137 & ~x142 & ~x165 & ~x166 & ~x167 & ~x171 & ~x172 & ~x197 & ~x199 & ~x200 & ~x221 & ~x222 & ~x226 & ~x250 & ~x306 & ~x334 & ~x338 & ~x391 & ~x418 & ~x447 & ~x477 & ~x501 & ~x503 & ~x504 & ~x519 & ~x530 & ~x531 & ~x558 & ~x561 & ~x573 & ~x574 & ~x575 & ~x587 & ~x588 & ~x589 & ~x603 & ~x614 & ~x673 & ~x729 & ~x754 & ~x757;
assign c2332 = ~x0 & ~x1 & ~x2 & ~x4 & ~x5 & ~x16 & ~x17 & ~x23 & ~x24 & ~x25 & ~x27 & ~x28 & ~x29 & ~x30 & ~x31 & ~x32 & ~x33 & ~x50 & ~x51 & ~x52 & ~x54 & ~x55 & ~x56 & ~x57 & ~x58 & ~x60 & ~x61 & ~x80 & ~x81 & ~x83 & ~x84 & ~x85 & ~x107 & ~x108 & ~x110 & ~x113 & ~x114 & ~x115 & ~x116 & ~x134 & ~x135 & ~x136 & ~x137 & ~x138 & ~x140 & ~x141 & ~x143 & ~x144 & ~x162 & ~x163 & ~x164 & ~x166 & ~x168 & ~x169 & ~x171 & ~x172 & ~x191 & ~x192 & ~x193 & ~x194 & ~x196 & ~x197 & ~x198 & ~x218 & ~x219 & ~x220 & ~x221 & ~x222 & ~x223 & ~x224 & ~x226 & ~x228 & ~x246 & ~x247 & ~x249 & ~x251 & ~x254 & ~x255 & ~x274 & ~x275 & ~x276 & ~x277 & ~x278 & ~x279 & ~x281 & ~x282 & ~x306 & ~x307 & ~x308 & ~x309 & ~x334 & ~x335 & ~x336 & ~x337 & ~x363 & ~x365 & ~x391 & ~x392 & ~x393 & ~x419 & ~x420 & ~x421 & ~x422 & ~x444 & ~x446 & ~x447 & ~x473 & ~x476 & ~x501 & ~x502 & ~x503 & ~x504 & ~x505 & ~x530 & ~x532 & ~x533 & ~x557 & ~x558 & ~x560 & ~x561 & ~x585 & ~x586 & ~x587 & ~x588 & ~x589 & ~x614 & ~x615 & ~x616 & ~x617 & ~x640 & ~x641 & ~x642 & ~x644 & ~x645 & ~x670 & ~x671 & ~x672 & ~x673 & ~x674 & ~x697 & ~x698 & ~x699 & ~x701 & ~x702 & ~x726 & ~x728 & ~x755 & ~x756 & ~x782;
assign c2334 = ~x5 & ~x6 & ~x7 & ~x21 & ~x25 & ~x34 & ~x37 & ~x47 & ~x53 & ~x55 & ~x56 & ~x61 & ~x76 & ~x82 & ~x83 & ~x103 & ~x114 & ~x117 & ~x118 & ~x121 & ~x168 & ~x169 & ~x174 & ~x175 & ~x180 & ~x196 & ~x391 & ~x417 & ~x418 & ~x422 & ~x446 & ~x454 & ~x472 & ~x474 & ~x478 & ~x481 & ~x483 & ~x505 & ~x506 & ~x511 & ~x528 & ~x529 & ~x539 & ~x557 & ~x560 & ~x561 & ~x564 & ~x565 & ~x567 & ~x584 & ~x591 & ~x595 & ~x596 & ~x597 & ~x611 & ~x615 & ~x617 & ~x620 & ~x626 & ~x639 & ~x643 & ~x644 & ~x648 & ~x649 & ~x653 & ~x668 & ~x672 & ~x675 & ~x680 & ~x682 & ~x694 & ~x697 & ~x702 & ~x706 & ~x722 & ~x723 & ~x724 & ~x725 & ~x726 & ~x727 & ~x728 & ~x731 & ~x735 & ~x750 & ~x751 & ~x756 & ~x757 & ~x759 & ~x778 & ~x779 & ~x782;
assign c2336 =  x510 &  x598 & ~x49 & ~x112 & ~x114 & ~x170 & ~x196 & ~x419 & ~x580 & ~x612 & ~x667 & ~x754 & ~x756;
assign c2338 =  x67 & ~x22 & ~x100 & ~x102 & ~x138 & ~x165 & ~x183 & ~x239 & ~x337 & ~x365 & ~x386 & ~x387 & ~x440 & ~x465 & ~x468 & ~x564 & ~x672 & ~x676 & ~x727;
assign c2340 =  x239 & ~x4 & ~x24 & ~x29 & ~x176 & ~x178 & ~x180 & ~x208 & ~x363 & ~x446 & ~x469 & ~x473 & ~x504 & ~x525 & ~x530 & ~x552 & ~x612 & ~x613 & ~x615 & ~x623 & ~x639 & ~x667 & ~x680 & ~x733 & ~x735;
assign c2342 = ~x5 & ~x24 & ~x26 & ~x48 & ~x79 & ~x83 & ~x102 & ~x104 & ~x113 & ~x130 & ~x132 & ~x158 & ~x170 & ~x189 & ~x219 & ~x222 & ~x241 & ~x243 & ~x247 & ~x251 & ~x254 & ~x256 & ~x259 & ~x268 & ~x283 & ~x303 & ~x323 & ~x363 & ~x366 & ~x395 & ~x414 & ~x444 & ~x448 & ~x473 & ~x500 & ~x504 & ~x534 & ~x551 & ~x553 & ~x561 & ~x589 & ~x608 & ~x634 & ~x639 & ~x641 & ~x663 & ~x666 & ~x671 & ~x707 & ~x732 & ~x777 & ~x780 & ~x782 & ~x783;
assign c2344 =  x343 & ~x3 & ~x6 & ~x24 & ~x28 & ~x30 & ~x32 & ~x61 & ~x78 & ~x79 & ~x82 & ~x83 & ~x87 & ~x105 & ~x107 & ~x133 & ~x137 & ~x140 & ~x141 & ~x165 & ~x166 & ~x168 & ~x169 & ~x171 & ~x189 & ~x191 & ~x195 & ~x196 & ~x197 & ~x198 & ~x199 & ~x222 & ~x225 & ~x227 & ~x251 & ~x281 & ~x307 & ~x336 & ~x365 & ~x386 & ~x388 & ~x389 & ~x390 & ~x391 & ~x414 & ~x419 & ~x420 & ~x421 & ~x442 & ~x448 & ~x450 & ~x470 & ~x471 & ~x473 & ~x474 & ~x475 & ~x499 & ~x503 & ~x504 & ~x505 & ~x525 & ~x527 & ~x530 & ~x553 & ~x554 & ~x558 & ~x559 & ~x561 & ~x581 & ~x582 & ~x586 & ~x589 & ~x608 & ~x610 & ~x612 & ~x615 & ~x638 & ~x643 & ~x649 & ~x670 & ~x671 & ~x673 & ~x675 & ~x695 & ~x696 & ~x727 & ~x761 & ~x780 & ~x781;
assign c2346 =  x317 & ~x54 & ~x63 & ~x76 & ~x117 & ~x131 & ~x195 & ~x384 & ~x386 & ~x399 & ~x500 & ~x509 & ~x522 & ~x524 & ~x533 & ~x580 & ~x596 & ~x637 & ~x641 & ~x723 & ~x781;
assign c2348 =  x285 & ~x26 & ~x27 & ~x54 & ~x82 & ~x83 & ~x110 & ~x111 & ~x114 & ~x140 & ~x331 & ~x359 & ~x360 & ~x362 & ~x373 & ~x387 & ~x390 & ~x391 & ~x415 & ~x419 & ~x444 & ~x445 & ~x446 & ~x447 & ~x453 & ~x473 & ~x482 & ~x503 & ~x509 & ~x755;
assign c2350 =  x132 &  x412 & ~x390 & ~x685 & ~x739;
assign c2352 = ~x57 & ~x69 & ~x82 & ~x111 & ~x140 & ~x277 & ~x279 & ~x305 & ~x343 & ~x363 & ~x388 & ~x391 & ~x398 & ~x399 & ~x426 & ~x454 & ~x473 & ~x482 & ~x503 & ~x509 & ~x544 & ~x572 & ~x599 & ~x600 & ~x655 & ~x681 & ~x717 & ~x745;
assign c2354 =  x45 &  x127 & ~x53 & ~x55 & ~x166 & ~x421 & ~x474 & ~x475 & ~x498 & ~x499 & ~x636 & ~x644 & ~x669 & ~x672 & ~x679 & ~x696 & ~x726 & ~x777;
assign c2356 =  x153 &  x410 &  x436 & ~x30 & ~x54 & ~x165 & ~x220 & ~x268 & ~x418 & ~x526 & ~x554 & ~x556 & ~x579 & ~x706;
assign c2358 =  x508 & ~x0 & ~x2 & ~x16 & ~x22 & ~x23 & ~x24 & ~x26 & ~x27 & ~x29 & ~x30 & ~x52 & ~x53 & ~x54 & ~x55 & ~x57 & ~x80 & ~x81 & ~x82 & ~x83 & ~x85 & ~x86 & ~x108 & ~x109 & ~x110 & ~x111 & ~x112 & ~x115 & ~x135 & ~x136 & ~x138 & ~x139 & ~x141 & ~x142 & ~x163 & ~x164 & ~x165 & ~x166 & ~x168 & ~x169 & ~x191 & ~x193 & ~x198 & ~x199 & ~x219 & ~x220 & ~x221 & ~x248 & ~x249 & ~x250 & ~x275 & ~x277 & ~x278 & ~x280 & ~x307 & ~x308 & ~x333 & ~x335 & ~x362 & ~x364 & ~x365 & ~x391 & ~x418 & ~x420 & ~x448 & ~x475 & ~x501 & ~x503 & ~x504 & ~x532 & ~x533 & ~x561 & ~x588 & ~x589 & ~x614 & ~x616 & ~x617 & ~x644 & ~x670 & ~x671 & ~x672 & ~x698 & ~x727 & ~x728 & ~x754 & ~x755 & ~x756;
assign c2360 =  x103 & ~x332 & ~x346 & ~x415 & ~x428 & ~x455 & ~x484 & ~x511 & ~x532 & ~x533 & ~x567 & ~x729;
assign c2362 =  x545 & ~x6 & ~x7 & ~x33 & ~x107 & ~x150 & ~x179 & ~x376 & ~x443 & ~x500 & ~x505 & ~x556 & ~x562 & ~x566 & ~x584 & ~x623 & ~x668;
assign c2364 =  x349 & ~x25 & ~x59 & ~x83 & ~x90 & ~x110 & ~x112 & ~x113 & ~x114 & ~x117 & ~x130 & ~x136 & ~x141 & ~x158 & ~x165 & ~x171 & ~x197 & ~x219 & ~x224 & ~x226 & ~x250 & ~x254 & ~x255 & ~x256 & ~x305 & ~x335 & ~x336 & ~x365 & ~x382 & ~x408 & ~x447 & ~x475 & ~x502 & ~x505 & ~x530 & ~x534 & ~x552 & ~x580 & ~x586 & ~x588 & ~x614 & ~x616 & ~x635 & ~x638 & ~x640 & ~x645 & ~x672 & ~x693 & ~x695 & ~x703 & ~x708 & ~x730 & ~x731 & ~x733 & ~x753 & ~x756 & ~x779 & ~x780;
assign c2366 =  x367 & ~x55 & ~x193 & ~x250 & ~x426 & ~x446 & ~x490;
assign c2368 =  x520 & ~x28 & ~x29 & ~x64 & ~x81 & ~x86 & ~x141 & ~x166 & ~x169 & ~x171 & ~x172 & ~x199 & ~x243 & ~x272 & ~x291 & ~x303 & ~x326 & ~x330 & ~x331 & ~x332 & ~x333 & ~x334 & ~x335 & ~x363 & ~x478 & ~x504 & ~x506 & ~x579 & ~x582 & ~x609 & ~x613 & ~x667 & ~x699 & ~x701 & ~x726 & ~x755 & ~x764 & ~x781;
assign c2370 =  x38 &  x376 & ~x491 & ~x518 & ~x575;
assign c2372 =  x123 & ~x2 & ~x21 & ~x28 & ~x29 & ~x51 & ~x54 & ~x55 & ~x58 & ~x80 & ~x82 & ~x84 & ~x87 & ~x106 & ~x110 & ~x113 & ~x114 & ~x132 & ~x139 & ~x140 & ~x143 & ~x158 & ~x167 & ~x170 & ~x186 & ~x188 & ~x190 & ~x192 & ~x193 & ~x194 & ~x196 & ~x198 & ~x199 & ~x218 & ~x222 & ~x247 & ~x252 & ~x253 & ~x276 & ~x277 & ~x310 & ~x335 & ~x336 & ~x389 & ~x392 & ~x447 & ~x470 & ~x471 & ~x472 & ~x473 & ~x474 & ~x476 & ~x497 & ~x498 & ~x499 & ~x500 & ~x501 & ~x502 & ~x503 & ~x504 & ~x523 & ~x526 & ~x527 & ~x529 & ~x550 & ~x551 & ~x555 & ~x557 & ~x577 & ~x580 & ~x582 & ~x583 & ~x584 & ~x585 & ~x586 & ~x604 & ~x610 & ~x611 & ~x613 & ~x615 & ~x617 & ~x619 & ~x634 & ~x637 & ~x641 & ~x643 & ~x646 & ~x648 & ~x649 & ~x666 & ~x670 & ~x671 & ~x675 & ~x676 & ~x677 & ~x695 & ~x702 & ~x705 & ~x709 & ~x729 & ~x730 & ~x734 & ~x735 & ~x754 & ~x759 & ~x761 & ~x781 & ~x782 & ~x783;
assign c2374 =  x104 & ~x69 & ~x82 & ~x112 & ~x217 & ~x218 & ~x220 & ~x223 & ~x247 & ~x274 & ~x275 & ~x277 & ~x278 & ~x305 & ~x308 & ~x316 & ~x331 & ~x334 & ~x359 & ~x414 & ~x415 & ~x446 & ~x473;
assign c2376 = ~x1 & ~x21 & ~x29 & ~x32 & ~x33 & ~x34 & ~x51 & ~x52 & ~x53 & ~x79 & ~x85 & ~x86 & ~x88 & ~x107 & ~x109 & ~x110 & ~x111 & ~x141 & ~x142 & ~x167 & ~x168 & ~x169 & ~x170 & ~x171 & ~x193 & ~x194 & ~x195 & ~x196 & ~x197 & ~x199 & ~x219 & ~x224 & ~x226 & ~x228 & ~x241 & ~x243 & ~x249 & ~x268 & ~x269 & ~x276 & ~x277 & ~x278 & ~x282 & ~x295 & ~x305 & ~x306 & ~x323 & ~x336 & ~x337 & ~x338 & ~x392 & ~x421 & ~x448 & ~x450 & ~x502 & ~x503 & ~x504 & ~x526 & ~x527 & ~x528 & ~x529 & ~x530 & ~x531 & ~x553 & ~x554 & ~x557 & ~x559 & ~x561 & ~x576 & ~x581 & ~x583 & ~x586 & ~x587 & ~x588 & ~x589 & ~x602 & ~x603 & ~x609 & ~x614 & ~x615 & ~x639 & ~x640 & ~x642 & ~x645 & ~x667 & ~x671 & ~x672 & ~x673 & ~x698 & ~x702 & ~x729 & ~x730 & ~x731 & ~x754 & ~x758;
assign c2378 =  x131 & ~x0 & ~x28 & ~x96 & ~x359 & ~x387 & ~x389 & ~x391 & ~x415 & ~x444 & ~x445 & ~x446 & ~x451 & ~x471 & ~x472 & ~x474 & ~x475 & ~x506 & ~x509 & ~x511 & ~x532 & ~x533 & ~x537 & ~x559 & ~x563 & ~x564 & ~x588 & ~x591 & ~x595 & ~x620 & ~x647 & ~x648 & ~x669 & ~x674 & ~x675 & ~x679 & ~x700 & ~x702 & ~x729 & ~x730 & ~x781;
assign c2380 = ~x0 & ~x2 & ~x17 & ~x18 & ~x19 & ~x22 & ~x23 & ~x25 & ~x26 & ~x28 & ~x29 & ~x30 & ~x47 & ~x52 & ~x57 & ~x76 & ~x79 & ~x87 & ~x89 & ~x103 & ~x107 & ~x112 & ~x113 & ~x114 & ~x115 & ~x130 & ~x133 & ~x136 & ~x143 & ~x144 & ~x163 & ~x164 & ~x165 & ~x168 & ~x172 & ~x189 & ~x194 & ~x197 & ~x199 & ~x200 & ~x201 & ~x216 & ~x230 & ~x243 & ~x244 & ~x245 & ~x246 & ~x249 & ~x250 & ~x253 & ~x269 & ~x280 & ~x281 & ~x299 & ~x306 & ~x308 & ~x309 & ~x325 & ~x326 & ~x327 & ~x330 & ~x333 & ~x337 & ~x352 & ~x360 & ~x363 & ~x366 & ~x388 & ~x389 & ~x393 & ~x419 & ~x421 & ~x446 & ~x447 & ~x474 & ~x475 & ~x476 & ~x477 & ~x502 & ~x503 & ~x506 & ~x528 & ~x531 & ~x533 & ~x561 & ~x579 & ~x580 & ~x581 & ~x605 & ~x607 & ~x609 & ~x610 & ~x614 & ~x619 & ~x634 & ~x637 & ~x638 & ~x642 & ~x664 & ~x668 & ~x672 & ~x696 & ~x701 & ~x705 & ~x724 & ~x726 & ~x727 & ~x728 & ~x729 & ~x732 & ~x734 & ~x753 & ~x755 & ~x756 & ~x759 & ~x761 & ~x762 & ~x763 & ~x782 & ~x783;
assign c2382 =  x484 & ~x1 & ~x26 & ~x51 & ~x53 & ~x78 & ~x81 & ~x108 & ~x109 & ~x111 & ~x112 & ~x113 & ~x114 & ~x134 & ~x138 & ~x139 & ~x140 & ~x142 & ~x189 & ~x191 & ~x193 & ~x196 & ~x197 & ~x199 & ~x213 & ~x214 & ~x216 & ~x226 & ~x243 & ~x250 & ~x253 & ~x334 & ~x337 & ~x417 & ~x418 & ~x419 & ~x444 & ~x445 & ~x446 & ~x496 & ~x497 & ~x500 & ~x524 & ~x527 & ~x529 & ~x530 & ~x552 & ~x559 & ~x581 & ~x584 & ~x617 & ~x621 & ~x644 & ~x646 & ~x648 & ~x649 & ~x699 & ~x700 & ~x701 & ~x704 & ~x728 & ~x729 & ~x730 & ~x757 & ~x759;
assign c2384 =  x353 &  x380 &  x407 & ~x27 & ~x54 & ~x115 & ~x169 & ~x194 & ~x240 & ~x248 & ~x295 & ~x305 & ~x413 & ~x419 & ~x420 & ~x526 & ~x672 & ~x759;
assign c2386 =  x326 &  x339 & ~x418;
assign c2388 =  x98 &  x239 & ~x11 & ~x60 & ~x146 & ~x387 & ~x416 & ~x418 & ~x452 & ~x453 & ~x455 & ~x484 & ~x505 & ~x506 & ~x508 & ~x530 & ~x536 & ~x555 & ~x563 & ~x593 & ~x595 & ~x611 & ~x613 & ~x619 & ~x620 & ~x624 & ~x626 & ~x646 & ~x652 & ~x654 & ~x671 & ~x674 & ~x677 & ~x695 & ~x707 & ~x708 & ~x725 & ~x762 & ~x778;
assign c2390 =  x133 & ~x29 & ~x248 & ~x249 & ~x275 & ~x276 & ~x277 & ~x291 & ~x303 & ~x304 & ~x318 & ~x335 & ~x360 & ~x361 & ~x372 & ~x399 & ~x418 & ~x447 & ~x475 & ~x482 & ~x756;
assign c2392 = ~x1 & ~x6 & ~x8 & ~x10 & ~x22 & ~x25 & ~x27 & ~x31 & ~x32 & ~x51 & ~x58 & ~x59 & ~x79 & ~x84 & ~x86 & ~x90 & ~x107 & ~x108 & ~x109 & ~x111 & ~x132 & ~x135 & ~x136 & ~x140 & ~x158 & ~x159 & ~x163 & ~x165 & ~x167 & ~x170 & ~x172 & ~x174 & ~x190 & ~x191 & ~x192 & ~x194 & ~x197 & ~x198 & ~x200 & ~x217 & ~x221 & ~x224 & ~x225 & ~x230 & ~x251 & ~x278 & ~x279 & ~x282 & ~x286 & ~x305 & ~x312 & ~x337 & ~x360 & ~x361 & ~x362 & ~x392 & ~x394 & ~x417 & ~x421 & ~x445 & ~x447 & ~x448 & ~x449 & ~x474 & ~x478 & ~x498 & ~x499 & ~x501 & ~x502 & ~x504 & ~x505 & ~x525 & ~x527 & ~x528 & ~x530 & ~x531 & ~x533 & ~x551 & ~x553 & ~x555 & ~x558 & ~x561 & ~x577 & ~x579 & ~x583 & ~x584 & ~x587 & ~x590 & ~x606 & ~x608 & ~x610 & ~x612 & ~x617 & ~x619 & ~x620 & ~x635 & ~x641 & ~x642 & ~x645 & ~x646 & ~x647 & ~x649 & ~x654 & ~x679 & ~x694 & ~x695 & ~x696 & ~x703 & ~x704 & ~x705 & ~x709 & ~x723 & ~x725 & ~x726 & ~x728 & ~x730 & ~x731 & ~x734 & ~x753 & ~x756 & ~x761 & ~x762 & ~x776 & ~x777;
assign c2394 = ~x43 & ~x165 & ~x192 & ~x246 & ~x361 & ~x416 & ~x417 & ~x419 & ~x434 & ~x435 & ~x463 & ~x473 & ~x544 & ~x627 & ~x682 & ~x720 & ~x746 & ~x747;
assign c2396 =  x678 &  x705 & ~x137 & ~x165 & ~x220 & ~x250 & ~x718 & ~x719 & ~x748;
assign c2398 =  x439 & ~x5 & ~x81 & ~x139 & ~x190 & ~x192 & ~x198 & ~x216 & ~x245 & ~x254 & ~x270 & ~x271 & ~x279 & ~x297 & ~x298 & ~x299 & ~x325 & ~x335 & ~x337 & ~x353 & ~x364 & ~x504 & ~x580 & ~x582 & ~x583 & ~x608 & ~x609 & ~x647 & ~x667 & ~x700 & ~x729 & ~x733 & ~x735;
assign c2400 =  x438 & ~x164 & ~x197 & ~x200 & ~x229 & ~x241 & ~x243 & ~x245 & ~x246 & ~x261 & ~x269 & ~x271 & ~x296 & ~x352 & ~x532 & ~x551 & ~x578 & ~x605 & ~x609 & ~x612 & ~x641;
assign c2402 =  x618 & ~x454;
assign c2404 =  x158 &  x410 &  x438 & ~x0 & ~x414 & ~x415 & ~x622 & ~x625 & ~x650 & ~x677 & ~x678 & ~x701 & ~x728 & ~x732 & ~x757 & ~x783;
assign c2406 = ~x0 & ~x1 & ~x3 & ~x5 & ~x23 & ~x25 & ~x27 & ~x29 & ~x30 & ~x53 & ~x55 & ~x57 & ~x58 & ~x84 & ~x85 & ~x86 & ~x96 & ~x124 & ~x140 & ~x150 & ~x168 & ~x332 & ~x333 & ~x334 & ~x335 & ~x346 & ~x359 & ~x360 & ~x361 & ~x362 & ~x363 & ~x372 & ~x373 & ~x387 & ~x389 & ~x399 & ~x400 & ~x416 & ~x417 & ~x418 & ~x419 & ~x426 & ~x443 & ~x445 & ~x447 & ~x472 & ~x474 & ~x475 & ~x481 & ~x482 & ~x503 & ~x510 & ~x511 & ~x531 & ~x538 & ~x588 & ~x696 & ~x698 & ~x727 & ~x728 & ~x754 & ~x755 & ~x756 & ~x757 & ~x759 & ~x760;
assign c2408 = ~x0 & ~x4 & ~x5 & ~x6 & ~x21 & ~x24 & ~x27 & ~x30 & ~x32 & ~x46 & ~x47 & ~x49 & ~x53 & ~x56 & ~x57 & ~x59 & ~x61 & ~x76 & ~x77 & ~x78 & ~x79 & ~x107 & ~x112 & ~x113 & ~x114 & ~x115 & ~x116 & ~x132 & ~x135 & ~x137 & ~x166 & ~x167 & ~x168 & ~x172 & ~x188 & ~x217 & ~x219 & ~x221 & ~x222 & ~x223 & ~x246 & ~x248 & ~x252 & ~x275 & ~x277 & ~x280 & ~x302 & ~x309 & ~x310 & ~x311 & ~x312 & ~x336 & ~x337 & ~x338 & ~x362 & ~x363 & ~x366 & ~x380 & ~x391 & ~x394 & ~x419 & ~x420 & ~x421 & ~x422 & ~x444 & ~x473 & ~x474 & ~x476 & ~x502 & ~x503 & ~x504 & ~x528 & ~x531 & ~x534 & ~x555 & ~x557 & ~x560 & ~x562 & ~x577 & ~x581 & ~x584 & ~x586 & ~x603 & ~x604 & ~x606 & ~x609 & ~x610 & ~x611 & ~x614 & ~x615 & ~x617 & ~x633 & ~x635 & ~x636 & ~x637 & ~x638 & ~x639 & ~x644 & ~x646 & ~x665 & ~x667 & ~x671 & ~x672 & ~x674 & ~x675 & ~x693 & ~x694 & ~x697 & ~x698 & ~x703 & ~x705 & ~x707 & ~x723 & ~x726 & ~x729 & ~x731 & ~x734 & ~x751 & ~x752 & ~x756 & ~x757 & ~x760 & ~x779 & ~x781 & ~x782 & ~x783;
assign c2410 = ~x18 & ~x22 & ~x25 & ~x26 & ~x47 & ~x48 & ~x51 & ~x52 & ~x54 & ~x55 & ~x59 & ~x62 & ~x77 & ~x82 & ~x84 & ~x85 & ~x105 & ~x106 & ~x107 & ~x108 & ~x109 & ~x115 & ~x134 & ~x135 & ~x143 & ~x144 & ~x147 & ~x163 & ~x165 & ~x168 & ~x172 & ~x186 & ~x190 & ~x191 & ~x193 & ~x194 & ~x199 & ~x213 & ~x215 & ~x217 & ~x218 & ~x220 & ~x225 & ~x226 & ~x228 & ~x241 & ~x243 & ~x246 & ~x248 & ~x249 & ~x251 & ~x254 & ~x273 & ~x275 & ~x276 & ~x277 & ~x283 & ~x302 & ~x305 & ~x306 & ~x307 & ~x308 & ~x334 & ~x335 & ~x359 & ~x361 & ~x362 & ~x363 & ~x366 & ~x367 & ~x368 & ~x386 & ~x387 & ~x388 & ~x389 & ~x390 & ~x391 & ~x392 & ~x394 & ~x416 & ~x418 & ~x419 & ~x420 & ~x423 & ~x443 & ~x449 & ~x451 & ~x472 & ~x477 & ~x480 & ~x498 & ~x499 & ~x503 & ~x505 & ~x506 & ~x526 & ~x529 & ~x530 & ~x531 & ~x532 & ~x533 & ~x550 & ~x552 & ~x554 & ~x557 & ~x558 & ~x559 & ~x563 & ~x580 & ~x582 & ~x583 & ~x588 & ~x592 & ~x606 & ~x609 & ~x610 & ~x611 & ~x615 & ~x616 & ~x638 & ~x641 & ~x648 & ~x649 & ~x653 & ~x664 & ~x665 & ~x667 & ~x670 & ~x672 & ~x675 & ~x681 & ~x695 & ~x698 & ~x699 & ~x701 & ~x703 & ~x705 & ~x706 & ~x709 & ~x722 & ~x723 & ~x726 & ~x727 & ~x729 & ~x731 & ~x733 & ~x737 & ~x750 & ~x751 & ~x754 & ~x755 & ~x757 & ~x759 & ~x760 & ~x761 & ~x763 & ~x776 & ~x778 & ~x779 & ~x781 & ~x783;
assign c2412 = ~x35 & ~x55 & ~x62 & ~x126 & ~x361 & ~x399 & ~x400 & ~x447 & ~x454 & ~x482 & ~x483 & ~x510 & ~x511 & ~x758;
assign c2414 =  x184 & ~x27 & ~x30 & ~x31 & ~x54 & ~x56 & ~x57 & ~x59 & ~x84 & ~x85 & ~x110 & ~x111 & ~x112 & ~x140 & ~x169 & ~x225 & ~x243 & ~x251 & ~x254 & ~x264 & ~x272 & ~x275 & ~x278 & ~x280 & ~x300 & ~x302 & ~x328 & ~x329 & ~x332 & ~x357 & ~x358 & ~x362 & ~x366 & ~x386 & ~x389 & ~x393 & ~x423 & ~x446 & ~x447 & ~x475 & ~x530 & ~x558 & ~x588 & ~x638 & ~x640 & ~x667 & ~x673 & ~x692 & ~x697 & ~x700 & ~x726 & ~x728 & ~x731 & ~x754 & ~x755 & ~x781;
assign c2416 =  x100 & ~x24 & ~x30 & ~x82 & ~x83 & ~x84 & ~x111 & ~x196 & ~x252 & ~x253 & ~x298 & ~x300 & ~x301 & ~x330 & ~x336 & ~x365 & ~x391 & ~x394 & ~x397 & ~x416 & ~x419 & ~x444 & ~x449 & ~x450 & ~x470 & ~x472 & ~x479 & ~x498 & ~x505 & ~x524 & ~x527 & ~x531 & ~x533 & ~x535 & ~x537 & ~x550 & ~x552 & ~x554 & ~x561 & ~x579 & ~x582 & ~x584 & ~x592 & ~x606 & ~x609 & ~x619 & ~x622 & ~x623 & ~x642 & ~x647 & ~x669 & ~x677 & ~x689 & ~x694 & ~x703 & ~x707 & ~x724 & ~x725 & ~x727 & ~x733 & ~x734 & ~x735 & ~x751 & ~x752 & ~x753 & ~x757 & ~x758 & ~x779 & ~x782;
assign c2418 =  x394 & ~x58 & ~x180 & ~x287 & ~x490;
assign c2420 = ~x320 & ~x332 & ~x392 & ~x399 & ~x400 & ~x401 & ~x428 & ~x442 & ~x444 & ~x452 & ~x456 & ~x474 & ~x483 & ~x485 & ~x503 & ~x511 & ~x512 & ~x514 & ~x529 & ~x530 & ~x532 & ~x534 & ~x535 & ~x542 & ~x543 & ~x569 & ~x590 & ~x592 & ~x596 & ~x599 & ~x626 & ~x639 & ~x649 & ~x654 & ~x670 & ~x680;
assign c2422 =  x316 & ~x33 & ~x61 & ~x81 & ~x82 & ~x85 & ~x105 & ~x106 & ~x108 & ~x114 & ~x117 & ~x131 & ~x146 & ~x159 & ~x164 & ~x196 & ~x198 & ~x391 & ~x393 & ~x413 & ~x414 & ~x416 & ~x443 & ~x471 & ~x479 & ~x506 & ~x531 & ~x538 & ~x557 & ~x585 & ~x592 & ~x593 & ~x615 & ~x621 & ~x622 & ~x650 & ~x651 & ~x692 & ~x723 & ~x752 & ~x778 & ~x780;
assign c2424 =  x76 & ~x24 & ~x390 & ~x399 & ~x427 & ~x446 & ~x455 & ~x566;
assign c2426 =  x478 &  x646;
assign c2428 = ~x25 & ~x27 & ~x28 & ~x33 & ~x55 & ~x58 & ~x60 & ~x61 & ~x99 & ~x110 & ~x127 & ~x138 & ~x142 & ~x143 & ~x169 & ~x196 & ~x248 & ~x250 & ~x275 & ~x276 & ~x305 & ~x332 & ~x334 & ~x335 & ~x391 & ~x417 & ~x436 & ~x437 & ~x444 & ~x490 & ~x501 & ~x510 & ~x737 & ~x780;
assign c2430 =  x382 & ~x0 & ~x22 & ~x24 & ~x32 & ~x50 & ~x55 & ~x56 & ~x77 & ~x81 & ~x106 & ~x107 & ~x108 & ~x110 & ~x111 & ~x134 & ~x137 & ~x140 & ~x144 & ~x161 & ~x164 & ~x167 & ~x168 & ~x172 & ~x190 & ~x193 & ~x196 & ~x213 & ~x219 & ~x220 & ~x222 & ~x223 & ~x243 & ~x253 & ~x269 & ~x270 & ~x279 & ~x280 & ~x297 & ~x309 & ~x335 & ~x390 & ~x420 & ~x445 & ~x473 & ~x496 & ~x498 & ~x502 & ~x504 & ~x524 & ~x547 & ~x552 & ~x553 & ~x555 & ~x581 & ~x583 & ~x584 & ~x586 & ~x588 & ~x589 & ~x611 & ~x614 & ~x639 & ~x671 & ~x672 & ~x677 & ~x699 & ~x703 & ~x706 & ~x725 & ~x727 & ~x732 & ~x733 & ~x734 & ~x753 & ~x754 & ~x758;
assign c2432 = ~x111 & ~x112 & ~x197 & ~x225 & ~x245 & ~x251 & ~x266 & ~x291 & ~x300 & ~x319 & ~x331 & ~x386 & ~x390 & ~x414 & ~x416 & ~x417 & ~x471 & ~x535 & ~x560 & ~x580 & ~x619 & ~x642 & ~x673 & ~x748 & ~x751 & ~x776;
assign c2434 =  x155 &  x182 & ~x31 & ~x55 & ~x114 & ~x224 & ~x242 & ~x270 & ~x271 & ~x277 & ~x302 & ~x354 & ~x362 & ~x367 & ~x370 & ~x389 & ~x416 & ~x422 & ~x443 & ~x473 & ~x476 & ~x479 & ~x552 & ~x606 & ~x609 & ~x617 & ~x673 & ~x698 & ~x705 & ~x719 & ~x723 & ~x728 & ~x730 & ~x751 & ~x758 & ~x779 & ~x780;
assign c2436 = ~x28 & ~x29 & ~x84 & ~x251 & ~x352 & ~x359 & ~x389 & ~x399 & ~x408 & ~x425 & ~x427 & ~x435 & ~x453 & ~x461 & ~x530 & ~x558 & ~x682;
assign c2438 = ~x86 & ~x157 & ~x199 & ~x238 & ~x278 & ~x307 & ~x389 & ~x466 & ~x467 & ~x474 & ~x491 & ~x518 & ~x757;
assign c2440 = ~x3 & ~x43 & ~x54 & ~x59 & ~x98 & ~x207 & ~x221 & ~x222 & ~x248 & ~x262 & ~x274 & ~x277 & ~x289 & ~x317 & ~x334 & ~x344 & ~x363 & ~x462 & ~x473 & ~x490 & ~x491 & ~x517 & ~x545 & ~x628 & ~x728 & ~x748 & ~x775;
assign c2442 =  x590 & ~x454;
assign c2444 =  x324 &  x377 & ~x133 & ~x157 & ~x185 & ~x437 & ~x467;
assign c2446 =  x69 &  x354 &  x380 &  x381 &  x407 & ~x53 & ~x54 & ~x56 & ~x78 & ~x103 & ~x108 & ~x165 & ~x169 & ~x194 & ~x195 & ~x196 & ~x240 & ~x253 & ~x418 & ~x475 & ~x530 & ~x531 & ~x552 & ~x556;
assign c2448 =  x339 & ~x389 & ~x407 & ~x736;
assign c2450 =  x72 &  x491 & ~x53 & ~x54 & ~x85 & ~x86 & ~x137 & ~x167 & ~x224 & ~x270 & ~x279 & ~x363 & ~x390 & ~x392 & ~x475 & ~x477 & ~x502 & ~x504 & ~x527 & ~x584 & ~x585 & ~x609 & ~x613 & ~x614 & ~x634 & ~x646 & ~x647 & ~x672 & ~x674 & ~x676 & ~x680 & ~x681 & ~x703 & ~x705 & ~x706 & ~x761 & ~x783;
assign c2452 =  x98 &  x154 &  x266 & ~x18 & ~x91 & ~x138 & ~x141 & ~x194 & ~x196 & ~x201 & ~x216 & ~x217 & ~x225 & ~x242 & ~x244 & ~x245 & ~x269 & ~x334 & ~x364 & ~x416 & ~x417 & ~x446 & ~x473 & ~x507 & ~x529 & ~x535 & ~x579 & ~x608 & ~x641 & ~x653 & ~x664 & ~x692 & ~x702 & ~x708;
assign c2454 = ~x8 & ~x24 & ~x84 & ~x124 & ~x251 & ~x279 & ~x321 & ~x345 & ~x359 & ~x362 & ~x363 & ~x373 & ~x392 & ~x396 & ~x398 & ~x416 & ~x424 & ~x425 & ~x426 & ~x448 & ~x452 & ~x454 & ~x455 & ~x475 & ~x477 & ~x482 & ~x502 & ~x529 & ~x530 & ~x536 & ~x538 & ~x561 & ~x564 & ~x565 & ~x568 & ~x593 & ~x595 & ~x615 & ~x616 & ~x620 & ~x644 & ~x650 & ~x668 & ~x670 & ~x672 & ~x677 & ~x697 & ~x703 & ~x731 & ~x756 & ~x757 & ~x760 & ~x761 & ~x781;
assign c2456 =  x449 & ~x424;
assign c2458 =  x184 & ~x0 & ~x2 & ~x29 & ~x30 & ~x32 & ~x54 & ~x140 & ~x271 & ~x277 & ~x292 & ~x300 & ~x318 & ~x327 & ~x330 & ~x363 & ~x365 & ~x388 & ~x392 & ~x396 & ~x413 & ~x414 & ~x415 & ~x422 & ~x423 & ~x446 & ~x447 & ~x449 & ~x451 & ~x452 & ~x471 & ~x472 & ~x505 & ~x526 & ~x528 & ~x532 & ~x552 & ~x556 & ~x559 & ~x582 & ~x587 & ~x610 & ~x615 & ~x641 & ~x645 & ~x647 & ~x648 & ~x649 & ~x670 & ~x675 & ~x697 & ~x704 & ~x726 & ~x727 & ~x729 & ~x754 & ~x756;
assign c2460 =  x216 & ~x148 & ~x388 & ~x416 & ~x533 & ~x534 & ~x555 & ~x558 & ~x564 & ~x583 & ~x591 & ~x594 & ~x595 & ~x644 & ~x651 & ~x653 & ~x672 & ~x673 & ~x705 & ~x735 & ~x782;
assign c2462 = ~x26 & ~x125 & ~x350 & ~x375 & ~x388 & ~x403 & ~x426 & ~x448 & ~x453 & ~x472 & ~x485 & ~x532 & ~x563 & ~x590 & ~x616 & ~x780;
assign c2464 =  x759;
assign c2466 = ~x2 & ~x30 & ~x32 & ~x34 & ~x50 & ~x51 & ~x54 & ~x56 & ~x57 & ~x61 & ~x82 & ~x83 & ~x90 & ~x112 & ~x113 & ~x139 & ~x173 & ~x193 & ~x196 & ~x197 & ~x200 & ~x221 & ~x225 & ~x275 & ~x303 & ~x305 & ~x331 & ~x334 & ~x360 & ~x361 & ~x372 & ~x388 & ~x391 & ~x392 & ~x415 & ~x420 & ~x428 & ~x444 & ~x456 & ~x477 & ~x484 & ~x503 & ~x505 & ~x506 & ~x511 & ~x532 & ~x533 & ~x538 & ~x539 & ~x561 & ~x627 & ~x645 & ~x670 & ~x671 & ~x673 & ~x698 & ~x744 & ~x745 & ~x746 & ~x755 & ~x770 & ~x774 & ~x775 & ~x781 & ~x782 & ~x783;
assign c2468 =  x185 &  x213 & ~x84 & ~x300 & ~x319 & ~x333 & ~x346 & ~x356 & ~x387 & ~x418 & ~x451 & ~x455 & ~x473 & ~x479 & ~x500 & ~x504 & ~x509 & ~x564 & ~x567 & ~x588 & ~x589 & ~x593 & ~x621 & ~x622 & ~x651 & ~x675 & ~x676 & ~x679 & ~x705;
assign c2470 = ~x51 & ~x89 & ~x92 & ~x130 & ~x135 & ~x189 & ~x211 & ~x228 & ~x280 & ~x393 & ~x438 & ~x464 & ~x478 & ~x499 & ~x594 & ~x610;
assign c2472 =  x287 & ~x52 & ~x76 & ~x84 & ~x104 & ~x105 & ~x111 & ~x135 & ~x137 & ~x140 & ~x165 & ~x197 & ~x278 & ~x330 & ~x358 & ~x364 & ~x385 & ~x387 & ~x396 & ~x424 & ~x445 & ~x451 & ~x475 & ~x476 & ~x501 & ~x528 & ~x534 & ~x553 & ~x556 & ~x559 & ~x584 & ~x591 & ~x616 & ~x671 & ~x696 & ~x700 & ~x702 & ~x725 & ~x736 & ~x763 & ~x781;
assign c2474 =  x648 & ~x125 & ~x261 & ~x407 & ~x491 & ~x546 & ~x656;
assign c2476 =  x405 & ~x110 & ~x139 & ~x140 & ~x157 & ~x171 & ~x198 & ~x249 & ~x281 & ~x304 & ~x332 & ~x360 & ~x415 & ~x445 & ~x465 & ~x471 & ~x520 & ~x530 & ~x729;
assign c2478 =  x454 &  x482 &  x515 & ~x59 & ~x85 & ~x164 & ~x167 & ~x171 & ~x194 & ~x221 & ~x248 & ~x249 & ~x446 & ~x554 & ~x582 & ~x644 & ~x697 & ~x703 & ~x759;
assign c2480 =  x186 & ~x3 & ~x54 & ~x55 & ~x152 & ~x391 & ~x418 & ~x420 & ~x428 & ~x450 & ~x452 & ~x455 & ~x473 & ~x479 & ~x482 & ~x483 & ~x506 & ~x508 & ~x511 & ~x534 & ~x535 & ~x536 & ~x588 & ~x592 & ~x593 & ~x614 & ~x615 & ~x641 & ~x648 & ~x649 & ~x652 & ~x673 & ~x680 & ~x696 & ~x700 & ~x701 & ~x731 & ~x732 & ~x733 & ~x753 & ~x759;
assign c2482 =  x231 & ~x3 & ~x23 & ~x24 & ~x26 & ~x56 & ~x82 & ~x85 & ~x86 & ~x111 & ~x137 & ~x168 & ~x300 & ~x328 & ~x331 & ~x334 & ~x356 & ~x364 & ~x366 & ~x388 & ~x389 & ~x390 & ~x392 & ~x413 & ~x415 & ~x417 & ~x419 & ~x420 & ~x442 & ~x443 & ~x470 & ~x471 & ~x475 & ~x478 & ~x483 & ~x500 & ~x503 & ~x504 & ~x505 & ~x527 & ~x555 & ~x584 & ~x586 & ~x610 & ~x613 & ~x673 & ~x674 & ~x675 & ~x699 & ~x752 & ~x754;
assign c2484 =  x561 & ~x425;
assign c2486 = ~x0 & ~x7 & ~x26 & ~x28 & ~x54 & ~x147 & ~x208 & ~x446 & ~x456 & ~x472 & ~x484 & ~x485 & ~x503 & ~x504 & ~x509 & ~x530 & ~x533 & ~x535 & ~x539 & ~x561 & ~x562 & ~x564 & ~x565 & ~x566 & ~x567 & ~x588 & ~x589 & ~x597 & ~x621 & ~x624 & ~x644 & ~x645 & ~x672 & ~x677 & ~x699 & ~x705 & ~x706 & ~x711 & ~x712 & ~x724 & ~x726 & ~x731 & ~x732 & ~x737 & ~x738 & ~x758 & ~x759 & ~x761;
assign c2488 = ~x26 & ~x51 & ~x53 & ~x57 & ~x113 & ~x136 & ~x169 & ~x222 & ~x305 & ~x307 & ~x310 & ~x311 & ~x327 & ~x328 & ~x335 & ~x338 & ~x354 & ~x380 & ~x389 & ~x390 & ~x418 & ~x476 & ~x525 & ~x527 & ~x528 & ~x531 & ~x560 & ~x577 & ~x579 & ~x585 & ~x606 & ~x631 & ~x646 & ~x648 & ~x660 & ~x662 & ~x667 & ~x668 & ~x693 & ~x708 & ~x721 & ~x752 & ~x777;
assign c2490 = ~x2 & ~x3 & ~x27 & ~x29 & ~x33 & ~x177 & ~x178 & ~x378 & ~x390 & ~x404 & ~x405 & ~x431 & ~x479 & ~x652 & ~x709 & ~x723 & ~x737 & ~x756 & ~x757 & ~x764 & ~x767 & ~x769;
assign c2492 =  x547 & ~x57 & ~x84 & ~x242 & ~x243 & ~x271 & ~x275 & ~x281 & ~x302 & ~x306 & ~x316 & ~x341 & ~x344 & ~x388 & ~x411 & ~x446 & ~x588 & ~x609 & ~x634 & ~x661 & ~x668 & ~x680 & ~x700 & ~x701;
assign c2494 =  x384 & ~x0 & ~x1 & ~x21 & ~x27 & ~x30 & ~x33 & ~x51 & ~x52 & ~x53 & ~x55 & ~x58 & ~x78 & ~x80 & ~x81 & ~x82 & ~x84 & ~x88 & ~x108 & ~x111 & ~x114 & ~x135 & ~x136 & ~x163 & ~x166 & ~x167 & ~x169 & ~x191 & ~x192 & ~x193 & ~x196 & ~x219 & ~x220 & ~x245 & ~x246 & ~x249 & ~x272 & ~x273 & ~x274 & ~x276 & ~x278 & ~x279 & ~x305 & ~x307 & ~x391 & ~x418 & ~x447 & ~x472 & ~x473 & ~x500 & ~x501 & ~x528 & ~x531 & ~x548 & ~x549 & ~x575 & ~x577 & ~x604;
assign c2496 =  x676 & ~x454;
assign c2498 =  x5 & ~x54 & ~x87 & ~x111 & ~x118 & ~x145 & ~x170 & ~x194 & ~x302 & ~x305 & ~x332 & ~x334 & ~x451 & ~x478 & ~x538 & ~x551 & ~x583 & ~x585 & ~x638 & ~x639 & ~x761;
assign c21 =  x296 &  x408 & ~x2 & ~x27 & ~x47 & ~x52 & ~x57 & ~x59 & ~x84 & ~x133 & ~x134 & ~x138 & ~x162 & ~x167 & ~x227 & ~x247 & ~x275 & ~x278 & ~x285 & ~x302 & ~x303 & ~x307 & ~x313 & ~x332 & ~x339 & ~x358 & ~x368 & ~x369 & ~x390 & ~x396 & ~x423 & ~x447 & ~x448 & ~x450 & ~x454 & ~x474 & ~x476 & ~x498 & ~x501 & ~x510 & ~x528 & ~x534 & ~x562 & ~x619 & ~x639 & ~x672 & ~x695 & ~x701 & ~x733 & ~x760 & ~x779 & ~x781;
assign c23 = ~x2 & ~x20 & ~x24 & ~x45 & ~x83 & ~x108 & ~x111 & ~x113 & ~x137 & ~x143 & ~x165 & ~x194 & ~x198 & ~x225 & ~x254 & ~x391 & ~x416 & ~x449 & ~x460 & ~x461 & ~x487 & ~x488 & ~x544 & ~x700 & ~x705 & ~x731 & ~x755 & ~x778 & ~x779 & ~x783;
assign c25 =  x251;
assign c27 = ~x0 & ~x25 & ~x50 & ~x54 & ~x83 & ~x105 & ~x116 & ~x120 & ~x133 & ~x134 & ~x140 & ~x143 & ~x148 & ~x163 & ~x165 & ~x189 & ~x201 & ~x202 & ~x221 & ~x228 & ~x231 & ~x232 & ~x252 & ~x254 & ~x262 & ~x277 & ~x312 & ~x333 & ~x339 & ~x343 & ~x365 & ~x368 & ~x371 & ~x389 & ~x395 & ~x397 & ~x399 & ~x400 & ~x401 & ~x419 & ~x420 & ~x427 & ~x453 & ~x476 & ~x481 & ~x495 & ~x504 & ~x505 & ~x526 & ~x536 & ~x588 & ~x612 & ~x618 & ~x671 & ~x672 & ~x698 & ~x699 & ~x704 & ~x706 & ~x733 & ~x762;
assign c29 =  x115;
assign c211 = ~x716;
assign c213 = ~x1 & ~x28 & ~x79 & ~x171 & ~x196 & ~x214 & ~x323 & ~x435 & ~x464 & ~x466 & ~x728 & ~x729;
assign c215 =  x479 & ~x12 & ~x373 & ~x514;
assign c217 =  x700;
assign c219 = ~x1 & ~x23 & ~x28 & ~x53 & ~x55 & ~x58 & ~x77 & ~x78 & ~x80 & ~x81 & ~x105 & ~x107 & ~x109 & ~x112 & ~x118 & ~x140 & ~x142 & ~x162 & ~x167 & ~x168 & ~x170 & ~x174 & ~x197 & ~x198 & ~x199 & ~x202 & ~x222 & ~x225 & ~x230 & ~x245 & ~x247 & ~x250 & ~x252 & ~x255 & ~x257 & ~x259 & ~x280 & ~x283 & ~x284 & ~x285 & ~x286 & ~x302 & ~x304 & ~x305 & ~x306 & ~x311 & ~x330 & ~x333 & ~x336 & ~x339 & ~x340 & ~x341 & ~x358 & ~x362 & ~x363 & ~x368 & ~x389 & ~x400 & ~x401 & ~x416 & ~x417 & ~x419 & ~x420 & ~x421 & ~x428 & ~x429 & ~x431 & ~x448 & ~x452 & ~x453 & ~x454 & ~x455 & ~x457 & ~x469 & ~x471 & ~x473 & ~x480 & ~x481 & ~x484 & ~x498 & ~x501 & ~x511 & ~x526 & ~x537 & ~x583 & ~x584 & ~x585 & ~x590 & ~x593 & ~x614 & ~x644 & ~x646 & ~x669 & ~x675 & ~x679 & ~x697 & ~x701 & ~x706 & ~x735 & ~x751 & ~x755 & ~x757 & ~x760 & ~x764 & ~x774 & ~x780;
assign c221 =  x757;
assign c223 =  x150 &  x178 &  x233 & ~x241 & ~x479 & ~x481 & ~x482;
assign c225 =  x719 & ~x381 & ~x410 & ~x412 & ~x468;
assign c227 =  x324 &  x553 & ~x613;
assign c229 =  x681 & ~x137 & ~x162 & ~x169 & ~x282 & ~x284 & ~x371 & ~x399 & ~x421 & ~x424 & ~x425 & ~x507 & ~x759;
assign c231 =  x418;
assign c233 =  x554 &  x594;
assign c235 = ~x22 & ~x33 & ~x59 & ~x64 & ~x80 & ~x88 & ~x107 & ~x134 & ~x140 & ~x146 & ~x165 & ~x203 & ~x230 & ~x252 & ~x253 & ~x259 & ~x303 & ~x306 & ~x313 & ~x335 & ~x339 & ~x368 & ~x430 & ~x431 & ~x445 & ~x455 & ~x456 & ~x457 & ~x459 & ~x469 & ~x472 & ~x477 & ~x479 & ~x482 & ~x484 & ~x527 & ~x528 & ~x531 & ~x539 & ~x554 & ~x563 & ~x594 & ~x621 & ~x641 & ~x645 & ~x647 & ~x649 & ~x702 & ~x726 & ~x750 & ~x761;
assign c237 =  x418;
assign c239 =  x738 & ~x452 & ~x658 & ~x683;
assign c241 =  x408 & ~x75 & ~x104 & ~x158 & ~x161 & ~x188 & ~x216 & ~x244 & ~x361 & ~x429 & ~x456 & ~x482 & ~x508 & ~x563 & ~x672;
assign c243 =  x375 &  x429 & ~x310 & ~x421 & ~x528 & ~x598 & ~x683;
assign c245 =  x55;
assign c247 =  x295 &  x353 & ~x25 & ~x103 & ~x159 & ~x188 & ~x272 & ~x335 & ~x358 & ~x362 & ~x416 & ~x452 & ~x476 & ~x478 & ~x534 & ~x561;
assign c251 = ~x22 & ~x67 & ~x82 & ~x108 & ~x112 & ~x123 & ~x152 & ~x159 & ~x190 & ~x220 & ~x370 & ~x372 & ~x425 & ~x448 & ~x500 & ~x503 & ~x558 & ~x613 & ~x614 & ~x694 & ~x697 & ~x725 & ~x732 & ~x760 & ~x763 & ~x780 & ~x783;
assign c253 = ~x1 & ~x22 & ~x23 & ~x28 & ~x30 & ~x32 & ~x33 & ~x37 & ~x49 & ~x78 & ~x79 & ~x80 & ~x82 & ~x89 & ~x104 & ~x105 & ~x106 & ~x112 & ~x115 & ~x135 & ~x140 & ~x163 & ~x164 & ~x168 & ~x173 & ~x190 & ~x195 & ~x200 & ~x201 & ~x222 & ~x224 & ~x231 & ~x249 & ~x250 & ~x257 & ~x259 & ~x260 & ~x273 & ~x275 & ~x276 & ~x279 & ~x281 & ~x283 & ~x286 & ~x288 & ~x289 & ~x305 & ~x309 & ~x313 & ~x314 & ~x315 & ~x325 & ~x332 & ~x335 & ~x336 & ~x339 & ~x340 & ~x354 & ~x355 & ~x362 & ~x367 & ~x383 & ~x387 & ~x389 & ~x391 & ~x394 & ~x397 & ~x398 & ~x412 & ~x418 & ~x421 & ~x424 & ~x425 & ~x439 & ~x442 & ~x449 & ~x450 & ~x454 & ~x466 & ~x468 & ~x476 & ~x478 & ~x479 & ~x481 & ~x500 & ~x502 & ~x503 & ~x508 & ~x522 & ~x525 & ~x530 & ~x531 & ~x551 & ~x555 & ~x556 & ~x562 & ~x563 & ~x584 & ~x587 & ~x588 & ~x589 & ~x591 & ~x609 & ~x612 & ~x620 & ~x644 & ~x645 & ~x647 & ~x671 & ~x672 & ~x674 & ~x698 & ~x729 & ~x730 & ~x752 & ~x753 & ~x755 & ~x759 & ~x765;
assign c255 = ~x37 & ~x54 & ~x69 & ~x81 & ~x112 & ~x126 & ~x154 & ~x282 & ~x283 & ~x394 & ~x420 & ~x503 & ~x523 & ~x733 & ~x739 & ~x740;
assign c257 = ~x158 & ~x184 & ~x237 & ~x429 & ~x563 & ~x664 & ~x705 & ~x726;
assign c259 = ~x1 & ~x23 & ~x28 & ~x79 & ~x84 & ~x89 & ~x115 & ~x117 & ~x139 & ~x149 & ~x161 & ~x170 & ~x175 & ~x190 & ~x201 & ~x220 & ~x225 & ~x226 & ~x227 & ~x230 & ~x246 & ~x257 & ~x279 & ~x290 & ~x310 & ~x317 & ~x339 & ~x344 & ~x358 & ~x362 & ~x371 & ~x372 & ~x394 & ~x425 & ~x426 & ~x440 & ~x499 & ~x500 & ~x506 & ~x510 & ~x554 & ~x565 & ~x590 & ~x593 & ~x596 & ~x621 & ~x623 & ~x650 & ~x668 & ~x676 & ~x677 & ~x698 & ~x728 & ~x736 & ~x759 & ~x765;
assign c261 =  x203 & ~x184 & ~x272 & ~x320;
assign c263 =  x502;
assign c265 = ~x105 & ~x155 & ~x773;
assign c267 =  x205 &  x289 &  x317 & ~x365 & ~x404;
assign c269 =  x270 & ~x5 & ~x29 & ~x30 & ~x47 & ~x160 & ~x248 & ~x274 & ~x278 & ~x280 & ~x287 & ~x288 & ~x332 & ~x388 & ~x421 & ~x614 & ~x699 & ~x762 & ~x779;
assign c271 = ~x6 & ~x23 & ~x26 & ~x48 & ~x50 & ~x56 & ~x60 & ~x61 & ~x62 & ~x64 & ~x83 & ~x88 & ~x106 & ~x120 & ~x143 & ~x161 & ~x164 & ~x166 & ~x167 & ~x202 & ~x245 & ~x248 & ~x251 & ~x258 & ~x260 & ~x261 & ~x275 & ~x280 & ~x285 & ~x331 & ~x333 & ~x334 & ~x341 & ~x357 & ~x364 & ~x366 & ~x391 & ~x418 & ~x447 & ~x449 & ~x454 & ~x458 & ~x469 & ~x482 & ~x485 & ~x497 & ~x502 & ~x503 & ~x510 & ~x512 & ~x513 & ~x527 & ~x530 & ~x531 & ~x536 & ~x537 & ~x556 & ~x558 & ~x562 & ~x565 & ~x568 & ~x582 & ~x585 & ~x595 & ~x611 & ~x612 & ~x613 & ~x668 & ~x669 & ~x671 & ~x695 & ~x699 & ~x723 & ~x725;
assign c273 =  x196;
assign c275 =  x602 & ~x101 & ~x129 & ~x293;
assign c277 =  x56;
assign c279 =  x323 & ~x33 & ~x76 & ~x104 & ~x144 & ~x161 & ~x165 & ~x167 & ~x204 & ~x223 & ~x246 & ~x247 & ~x255 & ~x276 & ~x281 & ~x303 & ~x330 & ~x342 & ~x358 & ~x372 & ~x424 & ~x425 & ~x454 & ~x476 & ~x556 & ~x557 & ~x560 & ~x582 & ~x645 & ~x700 & ~x781;
assign c281 =  x168;
assign c283 =  x417 &  x502;
assign c285 =  x579 & ~x20 & ~x77 & ~x107 & ~x136 & ~x199 & ~x278 & ~x334 & ~x369 & ~x416 & ~x417 & ~x734;
assign c287 = ~x0 & ~x2 & ~x3 & ~x32 & ~x49 & ~x50 & ~x51 & ~x52 & ~x55 & ~x56 & ~x59 & ~x77 & ~x79 & ~x84 & ~x86 & ~x88 & ~x106 & ~x111 & ~x113 & ~x114 & ~x133 & ~x135 & ~x138 & ~x141 & ~x143 & ~x164 & ~x169 & ~x172 & ~x173 & ~x191 & ~x192 & ~x193 & ~x194 & ~x196 & ~x198 & ~x199 & ~x220 & ~x223 & ~x225 & ~x228 & ~x247 & ~x253 & ~x254 & ~x255 & ~x258 & ~x274 & ~x275 & ~x282 & ~x285 & ~x288 & ~x289 & ~x302 & ~x303 & ~x305 & ~x310 & ~x312 & ~x314 & ~x315 & ~x331 & ~x332 & ~x333 & ~x334 & ~x336 & ~x339 & ~x340 & ~x342 & ~x343 & ~x384 & ~x388 & ~x390 & ~x394 & ~x395 & ~x396 & ~x415 & ~x416 & ~x418 & ~x421 & ~x423 & ~x424 & ~x439 & ~x440 & ~x441 & ~x442 & ~x443 & ~x445 & ~x449 & ~x450 & ~x469 & ~x470 & ~x471 & ~x472 & ~x474 & ~x475 & ~x496 & ~x499 & ~x502 & ~x504 & ~x505 & ~x525 & ~x529 & ~x531 & ~x532 & ~x533 & ~x535 & ~x559 & ~x584 & ~x586 & ~x639 & ~x640 & ~x641 & ~x698 & ~x699 & ~x700 & ~x702 & ~x727 & ~x729 & ~x730 & ~x733 & ~x756 & ~x760 & ~x761;
assign c289 =  x138;
assign c291 =  x473;
assign c293 = ~x11 & ~x12 & ~x13 & ~x18 & ~x28 & ~x40 & ~x41 & ~x44 & ~x50 & ~x54 & ~x58 & ~x68 & ~x71 & ~x82 & ~x83 & ~x151 & ~x392 & ~x670 & ~x679 & ~x699 & ~x708 & ~x726 & ~x778 & ~x782 & ~x783;
assign c295 =  x390;
assign c297 =  x177 & ~x74 & ~x108 & ~x250 & ~x402 & ~x429 & ~x618 & ~x724 & ~x760;
assign c299 =  x328 & ~x30 & ~x49 & ~x53 & ~x54 & ~x57 & ~x83 & ~x115 & ~x135 & ~x136 & ~x139 & ~x165 & ~x195 & ~x221 & ~x226 & ~x304 & ~x305 & ~x307 & ~x333 & ~x334 & ~x336 & ~x340 & ~x361 & ~x389 & ~x395 & ~x396 & ~x397 & ~x421 & ~x445 & ~x446 & ~x449 & ~x450 & ~x478 & ~x503 & ~x559 & ~x759;
assign c2101 =  x397 & ~x597 & ~x625 & ~x629 & ~x658 & ~x689 & ~x717;
assign c2103 =  x0;
assign c2105 =  x230 &  x332;
assign c2107 =  x419;
assign c2109 =  x272 & ~x48 & ~x52 & ~x53 & ~x55 & ~x87 & ~x106 & ~x108 & ~x109 & ~x110 & ~x164 & ~x219 & ~x220 & ~x224 & ~x247 & ~x251 & ~x252 & ~x276 & ~x280 & ~x303 & ~x305 & ~x333 & ~x334 & ~x335 & ~x360 & ~x421 & ~x445 & ~x446 & ~x474 & ~x724 & ~x726 & ~x751 & ~x765 & ~x778 & ~x779 & ~x781;
assign c2111 =  x447 & ~x100;
assign c2115 = ~x4 & ~x11 & ~x68 & ~x75 & ~x98 & ~x106 & ~x111 & ~x132 & ~x134 & ~x365 & ~x711 & ~x736 & ~x754 & ~x763 & ~x773;
assign c2117 =  x350 &  x683 & ~x336 & ~x428 & ~x563 & ~x764 & ~x765;
assign c2119 =  x375 &  x429 & ~x46 & ~x368 & ~x394 & ~x395;
assign c2121 = ~x138 & ~x154 & ~x376 & ~x515 & ~x566 & ~x645 & ~x746;
assign c2123 =  x756;
assign c2125 =  x712 & ~x162 & ~x302 & ~x313 & ~x512 & ~x514 & ~x515 & ~x537 & ~x538 & ~x620;
assign c2127 = ~x4 & ~x31 & ~x54 & ~x56 & ~x112 & ~x169 & ~x191 & ~x201 & ~x218 & ~x227 & ~x256 & ~x274 & ~x310 & ~x334 & ~x338 & ~x341 & ~x342 & ~x343 & ~x370 & ~x398 & ~x416 & ~x424 & ~x454 & ~x456 & ~x459 & ~x460 & ~x470 & ~x473 & ~x483 & ~x485 & ~x499 & ~x507 & ~x510 & ~x537 & ~x563 & ~x564 & ~x565 & ~x566 & ~x587 & ~x592 & ~x593 & ~x616 & ~x618 & ~x621 & ~x677 & ~x678 & ~x679 & ~x728 & ~x731 & ~x736 & ~x759 & ~x762 & ~x764 & ~x766;
assign c2129 =  x672;
assign c2131 = ~x20 & ~x30 & ~x32 & ~x48 & ~x49 & ~x50 & ~x57 & ~x63 & ~x75 & ~x78 & ~x80 & ~x81 & ~x85 & ~x89 & ~x104 & ~x111 & ~x112 & ~x115 & ~x134 & ~x138 & ~x141 & ~x143 & ~x146 & ~x160 & ~x161 & ~x170 & ~x193 & ~x200 & ~x201 & ~x217 & ~x218 & ~x219 & ~x220 & ~x221 & ~x223 & ~x226 & ~x227 & ~x229 & ~x247 & ~x277 & ~x282 & ~x283 & ~x312 & ~x341 & ~x343 & ~x344 & ~x345 & ~x357 & ~x359 & ~x361 & ~x362 & ~x363 & ~x364 & ~x368 & ~x369 & ~x371 & ~x374 & ~x392 & ~x393 & ~x396 & ~x397 & ~x398 & ~x400 & ~x416 & ~x418 & ~x419 & ~x420 & ~x442 & ~x446 & ~x450 & ~x455 & ~x478 & ~x500 & ~x504 & ~x507 & ~x528 & ~x530 & ~x534 & ~x535 & ~x536 & ~x537 & ~x557 & ~x558 & ~x559 & ~x585 & ~x586 & ~x590 & ~x592 & ~x609 & ~x613 & ~x615 & ~x617 & ~x637 & ~x639 & ~x647 & ~x649 & ~x676 & ~x677 & ~x693 & ~x696 & ~x723 & ~x757 & ~x761 & ~x764 & ~x780 & ~x783;
assign c2133 =  x127 &  x207 &  x262 &  x317;
assign c2135 =  x710 &  x739 & ~x1 & ~x50 & ~x87 & ~x110 & ~x132 & ~x161 & ~x168 & ~x169 & ~x171 & ~x191 & ~x222 & ~x248 & ~x391 & ~x417 & ~x427 & ~x428 & ~x452 & ~x455 & ~x508 & ~x534 & ~x560 & ~x616 & ~x618 & ~x670 & ~x782;
assign c2137 = ~x60 & ~x77 & ~x80 & ~x86 & ~x87 & ~x114 & ~x226 & ~x254 & ~x295 & ~x297 & ~x299 & ~x324 & ~x352 & ~x353 & ~x409 & ~x466 & ~x532 & ~x589 & ~x643 & ~x699 & ~x765 & ~x766 & ~x783;
assign c2139 =  x599 & ~x5 & ~x28 & ~x57 & ~x164 & ~x226 & ~x228 & ~x283 & ~x310 & ~x369 & ~x391 & ~x422 & ~x424 & ~x430 & ~x453 & ~x457 & ~x474 & ~x477 & ~x484 & ~x504 & ~x510 & ~x529 & ~x531 & ~x532 & ~x534 & ~x537 & ~x559 & ~x611 & ~x620 & ~x726 & ~x751 & ~x753 & ~x754 & ~x755 & ~x761 & ~x781;
assign c2141 =  x672;
assign c2143 =  x359;
assign c2145 = ~x20 & ~x22 & ~x24 & ~x29 & ~x30 & ~x32 & ~x48 & ~x53 & ~x60 & ~x61 & ~x62 & ~x63 & ~x84 & ~x85 & ~x106 & ~x140 & ~x145 & ~x164 & ~x166 & ~x172 & ~x173 & ~x190 & ~x191 & ~x192 & ~x197 & ~x200 & ~x202 & ~x222 & ~x223 & ~x225 & ~x227 & ~x229 & ~x232 & ~x249 & ~x279 & ~x304 & ~x308 & ~x309 & ~x313 & ~x314 & ~x331 & ~x334 & ~x335 & ~x338 & ~x340 & ~x357 & ~x360 & ~x364 & ~x403 & ~x416 & ~x419 & ~x426 & ~x428 & ~x429 & ~x430 & ~x442 & ~x446 & ~x447 & ~x448 & ~x454 & ~x472 & ~x481 & ~x501 & ~x534 & ~x535 & ~x560 & ~x561 & ~x562 & ~x564 & ~x583 & ~x591 & ~x594 & ~x610 & ~x618 & ~x620 & ~x640 & ~x675 & ~x679 & ~x701 & ~x704 & ~x721 & ~x729 & ~x732 & ~x748 & ~x749 & ~x754 & ~x757 & ~x758 & ~x760 & ~x761 & ~x779;
assign c2147 =  x454 & ~x42 & ~x71 & ~x432 & ~x459 & ~x460;
assign c2149 =  x389;
assign c2151 =  x244 & ~x162 & ~x165 & ~x254 & ~x258 & ~x310 & ~x313 & ~x340 & ~x504;
assign c2153 =  x201 & ~x236 & ~x265 & ~x293;
assign c2155 =  x718 & ~x32 & ~x54 & ~x84 & ~x88 & ~x105 & ~x164 & ~x228 & ~x250 & ~x251 & ~x339 & ~x369 & ~x383 & ~x445 & ~x467 & ~x499 & ~x578 & ~x588 & ~x698;
assign c2157 =  x418;
assign c2159 =  x136;
assign c2161 =  x725;
assign c2163 =  x360;
assign c2165 =  x496 & ~x584 & ~x635 & ~x718;
assign c2167 =  x439 & ~x130 & ~x167 & ~x222 & ~x481 & ~x536 & ~x726 & ~x746;
assign c2169 =  x700;
assign c2171 = ~x29 & ~x31 & ~x32 & ~x52 & ~x61 & ~x80 & ~x88 & ~x92 & ~x106 & ~x134 & ~x135 & ~x146 & ~x148 & ~x164 & ~x165 & ~x166 & ~x176 & ~x177 & ~x191 & ~x192 & ~x231 & ~x248 & ~x253 & ~x260 & ~x277 & ~x278 & ~x280 & ~x287 & ~x288 & ~x289 & ~x300 & ~x307 & ~x308 & ~x318 & ~x330 & ~x343 & ~x357 & ~x371 & ~x397 & ~x422 & ~x423 & ~x447 & ~x451 & ~x474 & ~x477 & ~x481 & ~x482 & ~x497 & ~x502 & ~x509 & ~x524 & ~x527 & ~x557 & ~x560 & ~x562 & ~x614 & ~x617 & ~x621 & ~x646 & ~x667 & ~x700 & ~x731 & ~x734 & ~x761 & ~x780;
assign c2173 = ~x54 & ~x321 & ~x353 & ~x463 & ~x466 & ~x493 & ~x732;
assign c2175 =  x473;
assign c2177 = ~x72 & ~x73 & ~x156 & ~x270 & ~x308 & ~x456 & ~x478 & ~x511 & ~x632 & ~x633 & ~x660;
assign c2179 =  x737 & ~x482 & ~x483 & ~x509 & ~x510;
assign c2181 =  x264 & ~x23 & ~x28 & ~x29 & ~x57 & ~x61 & ~x77 & ~x80 & ~x86 & ~x88 & ~x89 & ~x114 & ~x115 & ~x164 & ~x170 & ~x190 & ~x192 & ~x204 & ~x223 & ~x229 & ~x247 & ~x259 & ~x260 & ~x278 & ~x281 & ~x283 & ~x285 & ~x289 & ~x313 & ~x315 & ~x316 & ~x330 & ~x337 & ~x340 & ~x343 & ~x386 & ~x390 & ~x393 & ~x399 & ~x416 & ~x422 & ~x424 & ~x443 & ~x445 & ~x470 & ~x471 & ~x498 & ~x500 & ~x535 & ~x559 & ~x584 & ~x617 & ~x640 & ~x646 & ~x700;
assign c2183 = ~x6 & ~x20 & ~x51 & ~x83 & ~x84 & ~x107 & ~x115 & ~x135 & ~x145 & ~x172 & ~x195 & ~x198 & ~x219 & ~x222 & ~x224 & ~x228 & ~x251 & ~x252 & ~x258 & ~x283 & ~x284 & ~x285 & ~x309 & ~x312 & ~x313 & ~x315 & ~x336 & ~x342 & ~x364 & ~x367 & ~x385 & ~x396 & ~x416 & ~x422 & ~x426 & ~x427 & ~x430 & ~x431 & ~x432 & ~x441 & ~x443 & ~x444 & ~x446 & ~x448 & ~x451 & ~x454 & ~x455 & ~x456 & ~x457 & ~x458 & ~x469 & ~x476 & ~x481 & ~x502 & ~x510 & ~x537 & ~x555 & ~x588 & ~x592 & ~x615 & ~x621 & ~x639 & ~x643 & ~x664 & ~x671 & ~x680 & ~x693 & ~x694 & ~x699 & ~x702 & ~x721 & ~x725 & ~x727 & ~x728 & ~x753 & ~x756 & ~x758 & ~x759 & ~x765 & ~x778;
assign c2185 =  x482 & ~x181 & ~x405 & ~x422;
assign c2187 =  x268 & ~x18 & ~x76 & ~x104 & ~x132 & ~x160 & ~x217 & ~x278 & ~x311 & ~x330 & ~x336 & ~x343 & ~x345 & ~x449 & ~x470 & ~x509;
assign c2189 = ~x24 & ~x55 & ~x56 & ~x57 & ~x79 & ~x86 & ~x88 & ~x89 & ~x110 & ~x115 & ~x138 & ~x162 & ~x174 & ~x190 & ~x217 & ~x226 & ~x227 & ~x281 & ~x283 & ~x311 & ~x313 & ~x330 & ~x338 & ~x363 & ~x364 & ~x388 & ~x402 & ~x404 & ~x430 & ~x431 & ~x432 & ~x447 & ~x473 & ~x483 & ~x484 & ~x504 & ~x509 & ~x510 & ~x533 & ~x582 & ~x585 & ~x613 & ~x619 & ~x641 & ~x678 & ~x723 & ~x755 & ~x761;
assign c2191 =  x140;
assign c2193 =  x194;
assign c2195 = ~x54 & ~x57 & ~x77 & ~x135 & ~x137 & ~x143 & ~x165 & ~x194 & ~x198 & ~x223 & ~x249 & ~x255 & ~x278 & ~x332 & ~x334 & ~x335 & ~x363 & ~x382 & ~x393 & ~x401 & ~x402 & ~x403 & ~x404 & ~x429 & ~x431 & ~x432 & ~x456 & ~x474 & ~x507 & ~x512 & ~x530 & ~x559 & ~x567 & ~x584 & ~x594 & ~x595 & ~x618 & ~x646 & ~x668 & ~x706 & ~x724 & ~x726 & ~x729 & ~x736 & ~x765;
assign c2197 =  x231 & ~x100 & ~x270;
assign c2199 =  x85;
assign c2201 =  x397 & ~x11 & ~x40 & ~x41 & ~x349;
assign c2203 =  x334;
assign c2205 =  x184 &  x325 & ~x2 & ~x28 & ~x120 & ~x161 & ~x171 & ~x256 & ~x282 & ~x283 & ~x307 & ~x310 & ~x314 & ~x389 & ~x455 & ~x750 & ~x761 & ~x778;
assign c2207 =  x376 &  x403 & ~x20 & ~x26 & ~x61 & ~x77 & ~x78 & ~x79 & ~x107 & ~x143 & ~x173 & ~x201 & ~x221 & ~x223 & ~x230 & ~x252 & ~x261 & ~x288 & ~x303 & ~x312 & ~x339 & ~x342 & ~x343 & ~x359 & ~x362 & ~x367 & ~x370 & ~x371 & ~x399 & ~x422 & ~x451 & ~x469 & ~x471 & ~x478 & ~x480 & ~x505 & ~x558 & ~x614 & ~x641 & ~x645 & ~x671 & ~x701 & ~x702 & ~x728 & ~x783;
assign c2209 =  x154 &  x180 &  x235 & ~x75 & ~x76 & ~x170 & ~x198 & ~x254 & ~x256 & ~x417 & ~x594 & ~x648;
assign c2211 =  x151 &  x206 & ~x17 & ~x18 & ~x432 & ~x731 & ~x752;
assign c2213 = ~x0 & ~x54 & ~x77 & ~x79 & ~x108 & ~x115 & ~x116 & ~x137 & ~x191 & ~x196 & ~x200 & ~x219 & ~x222 & ~x247 & ~x311 & ~x346 & ~x375 & ~x376 & ~x402 & ~x417 & ~x512 & ~x587 & ~x669 & ~x697 & ~x705 & ~x729 & ~x751 & ~x756 & ~x765 & ~x773 & ~x778 & ~x779;
assign c2215 =  x147 & ~x11 & ~x152 & ~x180 & ~x441 & ~x448 & ~x671;
assign c2217 =  x88;
assign c2219 =  x424 & ~x13 & ~x430 & ~x541 & ~x542;
assign c2221 = ~x20 & ~x27 & ~x36 & ~x58 & ~x78 & ~x84 & ~x108 & ~x113 & ~x170 & ~x192 & ~x221 & ~x276 & ~x306 & ~x310 & ~x332 & ~x335 & ~x362 & ~x366 & ~x392 & ~x393 & ~x394 & ~x395 & ~x419 & ~x421 & ~x422 & ~x448 & ~x462 & ~x475 & ~x477 & ~x515 & ~x543 & ~x559 & ~x571 & ~x599 & ~x732 & ~x754 & ~x755 & ~x758 & ~x761 & ~x762 & ~x766 & ~x778 & ~x780;
assign c2223 =  x575 &  x626 & ~x306 & ~x595;
assign c2225 =  x152 &  x179 &  x234 & ~x6 & ~x256 & ~x284 & ~x446 & ~x475 & ~x482 & ~x506 & ~x509 & ~x535 & ~x671;
assign c2227 =  x178 &  x206 &  x233 &  x575;
assign c2229 =  x417;
assign c2231 = ~x134 & ~x167 & ~x275 & ~x360 & ~x368 & ~x371 & ~x373 & ~x384 & ~x398 & ~x449 & ~x509 & ~x547 & ~x555 & ~x557 & ~x573;
assign c2233 =  x391;
assign c2235 =  x406 &  x434 &  x491 & ~x28 & ~x33 & ~x53 & ~x56 & ~x82 & ~x89 & ~x105 & ~x115 & ~x131 & ~x188 & ~x245 & ~x256 & ~x331 & ~x336 & ~x368 & ~x391 & ~x392 & ~x393 & ~x419 & ~x421 & ~x445 & ~x477 & ~x479 & ~x484 & ~x505 & ~x509 & ~x536 & ~x538 & ~x669 & ~x695 & ~x751;
assign c2237 = ~x19 & ~x55 & ~x104 & ~x205 & ~x206 & ~x253 & ~x392 & ~x570 & ~x595 & ~x596 & ~x599 & ~x623 & ~x630 & ~x657;
assign c2239 =  x444;
assign c2241 =  x728;
assign c2243 = ~x0 & ~x50 & ~x84 & ~x89 & ~x136 & ~x139 & ~x167 & ~x234 & ~x311 & ~x329 & ~x357 & ~x370 & ~x407 & ~x464 & ~x468 & ~x469 & ~x615 & ~x698 & ~x702;
assign c2245 =  x335;
assign c2247 =  x680 & ~x459 & ~x460 & ~x752;
assign c2249 =  x475;
assign c2251 =  x135 & ~x244;
assign c2253 = ~x1 & ~x20 & ~x24 & ~x46 & ~x69 & ~x74 & ~x75 & ~x80 & ~x96 & ~x97 & ~x98 & ~x102 & ~x103 & ~x104 & ~x108 & ~x188 & ~x421 & ~x445 & ~x642 & ~x667 & ~x668 & ~x707 & ~x753 & ~x755 & ~x757 & ~x763 & ~x764 & ~x778 & ~x782;
assign c2255 = ~x2 & ~x7 & ~x27 & ~x79 & ~x90 & ~x140 & ~x248 & ~x253 & ~x322 & ~x323 & ~x337 & ~x379 & ~x408 & ~x492 & ~x521 & ~x674 & ~x701 & ~x703 & ~x727 & ~x732 & ~x754;
assign c2257 =  x203 &  x317 & ~x15 & ~x725 & ~x740;
assign c2259 =  x251;
assign c2261 = ~x1 & ~x18 & ~x24 & ~x48 & ~x49 & ~x50 & ~x59 & ~x78 & ~x80 & ~x105 & ~x140 & ~x223 & ~x309 & ~x365 & ~x374 & ~x390 & ~x393 & ~x429 & ~x456 & ~x484 & ~x539 & ~x603 & ~x674 & ~x679 & ~x698 & ~x707 & ~x722 & ~x724 & ~x731 & ~x733 & ~x734 & ~x736 & ~x759 & ~x761 & ~x764 & ~x782;
assign c2263 =  x122 & ~x101 & ~x129 & ~x401 & ~x428 & ~x480 & ~x481 & ~x536 & ~x590;
assign c2265 =  x179 &  x234 &  x262 &  x289 &  x317 & ~x2 & ~x26 & ~x30 & ~x32 & ~x140 & ~x311 & ~x340 & ~x422 & ~x447 & ~x530 & ~x783;
assign c2267 =  x447;
assign c2269 =  x757;
assign c2271 =  x174 &  x230 & ~x542;
assign c2273 = ~x69 & ~x99 & ~x126 & ~x158 & ~x337 & ~x476 & ~x529 & ~x714 & ~x741 & ~x746 & ~x756;
assign c2275 =  x27;
assign c2277 =  x692 & ~x368 & ~x370;
assign c2279 =  x530;
assign c2281 =  x328 & ~x51 & ~x77 & ~x78 & ~x79 & ~x108 & ~x109 & ~x168 & ~x278 & ~x332 & ~x361 & ~x366 & ~x393 & ~x421 & ~x433 & ~x728 & ~x759;
assign c2283 = ~x22 & ~x23 & ~x27 & ~x33 & ~x79 & ~x82 & ~x84 & ~x104 & ~x107 & ~x111 & ~x114 & ~x138 & ~x165 & ~x224 & ~x281 & ~x304 & ~x310 & ~x377 & ~x406 & ~x463 & ~x465 & ~x521 & ~x643;
assign c2285 =  x582 & ~x337 & ~x676;
assign c2287 =  x554 & ~x159 & ~x761;
assign c2289 =  x539 & ~x5 & ~x58 & ~x59 & ~x86 & ~x99 & ~x224 & ~x280 & ~x309 & ~x363 & ~x392 & ~x504 & ~x505 & ~x570 & ~x598 & ~x626 & ~x682 & ~x710;
assign c2291 =  x718 &  x720 & ~x53 & ~x326 & ~x384 & ~x467;
assign c2293 =  x191;
assign c2295 =  x264 &  x319 & ~x1 & ~x5 & ~x6 & ~x50 & ~x54 & ~x77 & ~x78 & ~x79 & ~x85 & ~x105 & ~x106 & ~x114 & ~x116 & ~x117 & ~x138 & ~x143 & ~x145 & ~x164 & ~x166 & ~x174 & ~x227 & ~x248 & ~x252 & ~x256 & ~x280 & ~x283 & ~x303 & ~x305 & ~x307 & ~x309 & ~x313 & ~x315 & ~x331 & ~x341 & ~x342 & ~x344 & ~x368 & ~x371 & ~x395 & ~x425 & ~x453 & ~x479 & ~x480 & ~x501 & ~x505 & ~x529 & ~x534 & ~x555 & ~x563 & ~x585 & ~x588 & ~x589 & ~x614 & ~x616 & ~x669 & ~x674 & ~x675 & ~x676 & ~x694 & ~x700 & ~x704 & ~x705 & ~x723 & ~x724 & ~x727 & ~x734 & ~x735 & ~x760 & ~x762 & ~x763 & ~x764;
assign c2297 =  x739 &  x740 &  x743 & ~x104 & ~x229 & ~x256 & ~x399 & ~x426 & ~x453 & ~x507 & ~x533 & ~x673;
assign c2299 =  x43 &  x240 & ~x113 & ~x137 & ~x160 & ~x189 & ~x245 & ~x313 & ~x333 & ~x369 & ~x388 & ~x476 & ~x506 & ~x508 & ~x533 & ~x646 & ~x758 & ~x759;
assign c2301 =  x193;
assign c2303 =  x305;
assign c2305 =  x57;
assign c2307 =  x32;
assign c2309 = ~x0 & ~x1 & ~x28 & ~x47 & ~x49 & ~x50 & ~x51 & ~x54 & ~x56 & ~x60 & ~x62 & ~x63 & ~x83 & ~x88 & ~x90 & ~x105 & ~x108 & ~x113 & ~x118 & ~x134 & ~x135 & ~x138 & ~x140 & ~x145 & ~x168 & ~x170 & ~x171 & ~x177 & ~x191 & ~x193 & ~x200 & ~x203 & ~x204 & ~x218 & ~x219 & ~x222 & ~x225 & ~x226 & ~x246 & ~x249 & ~x256 & ~x271 & ~x274 & ~x277 & ~x280 & ~x282 & ~x283 & ~x309 & ~x312 & ~x317 & ~x318 & ~x330 & ~x331 & ~x335 & ~x340 & ~x344 & ~x345 & ~x358 & ~x362 & ~x365 & ~x368 & ~x385 & ~x390 & ~x396 & ~x397 & ~x398 & ~x414 & ~x415 & ~x419 & ~x441 & ~x448 & ~x452 & ~x453 & ~x474 & ~x478 & ~x505 & ~x509 & ~x555 & ~x582 & ~x583 & ~x584 & ~x593 & ~x611 & ~x612 & ~x616 & ~x617 & ~x638 & ~x667 & ~x672 & ~x673 & ~x694 & ~x697 & ~x700 & ~x701 & ~x703 & ~x704 & ~x723 & ~x729 & ~x734 & ~x749 & ~x752 & ~x760 & ~x779;
assign c2311 =  x452 & ~x11 & ~x13 & ~x402 & ~x430;
assign c2313 =  x738 & ~x683 & ~x685;
assign c2315 = ~x9 & ~x27 & ~x110 & ~x196 & ~x351 & ~x380 & ~x393 & ~x408 & ~x437 & ~x520 & ~x553 & ~x615 & ~x641 & ~x674 & ~x709 & ~x752 & ~x757 & ~x765;
assign c2317 =  x454 & ~x28 & ~x30 & ~x59 & ~x85 & ~x360 & ~x392 & ~x393 & ~x422 & ~x449 & ~x487 & ~x542 & ~x543 & ~x598 & ~x682;
assign c2319 =  x501;
assign c2321 =  x235 &  x262 &  x290 & ~x8 & ~x27 & ~x37 & ~x39 & ~x57 & ~x81 & ~x226 & ~x253 & ~x256 & ~x285 & ~x307 & ~x338 & ~x361 & ~x418 & ~x445 & ~x532 & ~x642 & ~x700 & ~x757;
assign c2323 =  x682 & ~x485 & ~x486 & ~x567 & ~x764;
assign c2325 = ~x2 & ~x3 & ~x27 & ~x29 & ~x50 & ~x54 & ~x55 & ~x57 & ~x59 & ~x60 & ~x73 & ~x78 & ~x82 & ~x108 & ~x165 & ~x167 & ~x194 & ~x225 & ~x226 & ~x248 & ~x255 & ~x285 & ~x308 & ~x333 & ~x334 & ~x337 & ~x364 & ~x419 & ~x445 & ~x448 & ~x458 & ~x459 & ~x475 & ~x484 & ~x485 & ~x528 & ~x539 & ~x560 & ~x566 & ~x567 & ~x593 & ~x594 & ~x595 & ~x613 & ~x616 & ~x618 & ~x645 & ~x646 & ~x670 & ~x694 & ~x700 & ~x703 & ~x704 & ~x721 & ~x726 & ~x728 & ~x732 & ~x733 & ~x760 & ~x764;
assign c2327 =  x528;
assign c2329 =  x178 &  x233 &  x261 &  x288 & ~x352;
assign c2331 =  x502;
assign c2333 =  x303 & ~x321;
assign c2335 = ~x4 & ~x20 & ~x26 & ~x35 & ~x63 & ~x88 & ~x92 & ~x105 & ~x107 & ~x115 & ~x146 & ~x147 & ~x148 & ~x162 & ~x173 & ~x189 & ~x190 & ~x193 & ~x202 & ~x245 & ~x253 & ~x257 & ~x274 & ~x275 & ~x316 & ~x317 & ~x318 & ~x332 & ~x344 & ~x345 & ~x361 & ~x372 & ~x387 & ~x390 & ~x399 & ~x445 & ~x456 & ~x469 & ~x470 & ~x479 & ~x499 & ~x506 & ~x509 & ~x526 & ~x529 & ~x533 & ~x536 & ~x539 & ~x554 & ~x555 & ~x582 & ~x584 & ~x589 & ~x591 & ~x610 & ~x613 & ~x641 & ~x643 & ~x644 & ~x662 & ~x675 & ~x676 & ~x695 & ~x701 & ~x703 & ~x723 & ~x732 & ~x749 & ~x780;
assign c2337 = ~x1 & ~x5 & ~x19 & ~x30 & ~x57 & ~x59 & ~x108 & ~x137 & ~x138 & ~x139 & ~x158 & ~x304 & ~x323 & ~x334 & ~x337 & ~x391 & ~x392 & ~x417 & ~x421 & ~x448 & ~x487 & ~x515 & ~x531 & ~x543 & ~x568 & ~x570 & ~x571 & ~x699 & ~x708 & ~x765 & ~x783;
assign c2339 =  x429 &  x483 &  x510 & ~x450 & ~x478;
assign c2341 =  x325 &  x438 & ~x158 & ~x244 & ~x254 & ~x273 & ~x280;
assign c2343 =  x551 & ~x105 & ~x137 & ~x195 & ~x219 & ~x254 & ~x284 & ~x312 & ~x368 & ~x762;
assign c2345 = ~x14 & ~x21 & ~x40 & ~x70 & ~x126 & ~x184 & ~x496 & ~x497;
assign c2347 =  x359 & ~x40;
assign c2349 =  x297 & ~x26 & ~x30 & ~x77 & ~x116 & ~x118 & ~x123 & ~x124 & ~x161 & ~x171 & ~x190 & ~x192 & ~x196 & ~x197 & ~x229 & ~x255 & ~x283 & ~x308 & ~x314 & ~x331 & ~x422 & ~x477 & ~x501 & ~x618 & ~x647 & ~x671 & ~x705 & ~x752 & ~x781;
assign c2351 = ~x29 & ~x79 & ~x81 & ~x115 & ~x143 & ~x163 & ~x168 & ~x197 & ~x228 & ~x278 & ~x339 & ~x350 & ~x351 & ~x379 & ~x392 & ~x407 & ~x421 & ~x422 & ~x425 & ~x504 & ~x558 & ~x585 & ~x611 & ~x612 & ~x613 & ~x649 & ~x677 & ~x705 & ~x706 & ~x726 & ~x734 & ~x735 & ~x759 & ~x763;
assign c2353 =  x581;
assign c2355 = ~x40 & ~x42 & ~x55 & ~x98 & ~x102 & ~x183 & ~x184 & ~x393 & ~x418 & ~x421 & ~x692 & ~x698 & ~x699 & ~x721;
assign c2357 =  x359 & ~x41;
assign c2359 =  x485 &  x512 &  x539 & ~x449 & ~x453 & ~x507 & ~x533 & ~x586;
assign c2361 = ~x4 & ~x25 & ~x32 & ~x33 & ~x54 & ~x55 & ~x59 & ~x61 & ~x78 & ~x82 & ~x109 & ~x115 & ~x136 & ~x143 & ~x170 & ~x172 & ~x175 & ~x177 & ~x190 & ~x195 & ~x200 & ~x201 & ~x202 & ~x228 & ~x229 & ~x232 & ~x245 & ~x246 & ~x256 & ~x278 & ~x287 & ~x303 & ~x306 & ~x312 & ~x313 & ~x341 & ~x344 & ~x366 & ~x373 & ~x374 & ~x391 & ~x416 & ~x422 & ~x426 & ~x429 & ~x443 & ~x445 & ~x447 & ~x451 & ~x453 & ~x473 & ~x474 & ~x481 & ~x482 & ~x483 & ~x501 & ~x507 & ~x534 & ~x535 & ~x555 & ~x558 & ~x563 & ~x564 & ~x643 & ~x728 & ~x729 & ~x730 & ~x731 & ~x762 & ~x782;
assign c2363 =  x621 & ~x14 & ~x236 & ~x393 & ~x597;
assign c2365 =  x232 &  x287 & ~x14 & ~x15 & ~x45 & ~x110 & ~x322;
assign c2367 =  x628 & ~x12 & ~x142 & ~x165 & ~x195 & ~x310 & ~x331 & ~x333 & ~x394 & ~x402 & ~x455 & ~x456 & ~x482 & ~x483 & ~x560 & ~x615;
assign c2369 =  x204 & ~x18 & ~x44 & ~x371 & ~x393 & ~x425 & ~x451 & ~x508 & ~x645;
assign c2371 = ~x14 & ~x15 & ~x30 & ~x42 & ~x43 & ~x44 & ~x51 & ~x52 & ~x79 & ~x100 & ~x101 & ~x166 & ~x252 & ~x254 & ~x282 & ~x309 & ~x310 & ~x363 & ~x364 & ~x377 & ~x461 & ~x721 & ~x724 & ~x781;
assign c2373 =  x598 & ~x334 & ~x425 & ~x458 & ~x467 & ~x511;
assign c2375 =  x361;
assign c2377 =  x540 & ~x3 & ~x30 & ~x53 & ~x86 & ~x157 & ~x163 & ~x199 & ~x225 & ~x247 & ~x252 & ~x276 & ~x278 & ~x335 & ~x394 & ~x396 & ~x399 & ~x421 & ~x426 & ~x450 & ~x480 & ~x531 & ~x557 & ~x755;
assign c2379 =  x527;
assign c2381 =  x502;
assign c2383 =  x195;
assign c2385 =  x498 & ~x131;
assign c2387 =  x250;
assign c2389 =  x535 & ~x514 & ~x597;
assign c2391 = ~x0 & ~x49 & ~x70 & ~x73 & ~x84 & ~x101 & ~x102 & ~x187 & ~x252 & ~x334 & ~x365 & ~x372 & ~x389 & ~x397 & ~x422 & ~x424 & ~x445 & ~x452 & ~x453 & ~x454 & ~x476 & ~x506 & ~x559 & ~x699;
assign c2393 =  x332;
assign c2395 =  x554 & ~x104 & ~x561;
assign c2397 =  x174 & ~x181 & ~x459;
assign c2399 =  x745 & ~x29 & ~x111 & ~x170 & ~x198 & ~x200 & ~x220 & ~x282 & ~x339 & ~x340 & ~x355 & ~x381 & ~x412 & ~x422 & ~x440 & ~x506 & ~x521 & ~x522 & ~x532 & ~x550 & ~x758;
assign c2401 =  x202 & ~x11 & ~x152 & ~x180 & ~x181 & ~x188;
assign c2403 =  x274 & ~x279 & ~x306 & ~x307 & ~x367 & ~x421 & ~x423 & ~x478;
assign c2405 =  x208 & ~x58 & ~x79 & ~x168 & ~x199 & ~x225 & ~x254 & ~x256 & ~x304 & ~x426 & ~x453 & ~x458 & ~x459 & ~x485 & ~x510 & ~x511 & ~x512 & ~x563 & ~x642 & ~x757;
assign c2407 =  x333;
assign c2409 =  x379 & ~x24 & ~x75 & ~x104 & ~x113 & ~x138 & ~x158 & ~x166 & ~x338 & ~x372 & ~x373 & ~x394 & ~x399 & ~x480 & ~x501 & ~x764;
assign c2411 =  x595 & ~x201 & ~x305 & ~x339 & ~x363 & ~x422 & ~x427 & ~x454 & ~x481 & ~x533 & ~x534 & ~x726;
assign c2413 =  x379 &  x407 &  x491 & ~x75 & ~x104 & ~x162 & ~x196 & ~x280 & ~x425 & ~x481 & ~x483 & ~x485 & ~x509 & ~x511 & ~x539 & ~x562 & ~x591 & ~x646 & ~x736 & ~x765;
assign c2415 =  x418;
assign c2417 =  x179 &  x290 & ~x9 & ~x29 & ~x312;
assign c2419 =  x320 &  x745 & ~x48 & ~x53 & ~x57 & ~x78 & ~x81 & ~x108 & ~x113 & ~x168 & ~x199 & ~x282 & ~x283 & ~x338 & ~x345 & ~x372 & ~x398 & ~x415 & ~x421 & ~x425 & ~x427 & ~x472 & ~x474 & ~x585 & ~x587 & ~x643 & ~x757;
assign c2421 =  x390;
assign c2423 =  x224;
assign c2425 = ~x7 & ~x11 & ~x20 & ~x40 & ~x77 & ~x125 & ~x206 & ~x336 & ~x337 & ~x392 & ~x416 & ~x449 & ~x615 & ~x744 & ~x763 & ~x773 & ~x783;
assign c2427 =  x582 & ~x337 & ~x386 & ~x761 & ~x762;
assign c2429 =  x234 & ~x20 & ~x22 & ~x34 & ~x140 & ~x200 & ~x201 & ~x224 & ~x226 & ~x227 & ~x428 & ~x450 & ~x454 & ~x458 & ~x477 & ~x481 & ~x503 & ~x507 & ~x561 & ~x584 & ~x643 & ~x674 & ~x675 & ~x696 & ~x699 & ~x732 & ~x764 & ~x766;
assign c2431 =  x59;
assign c2433 =  x30;
assign c2435 =  x206 &  x290 & ~x1 & ~x66 & ~x83 & ~x195 & ~x284 & ~x287 & ~x480 & ~x759;
assign c2437 =  x307;
assign c2439 =  x709 & ~x456 & ~x508 & ~x510 & ~x535;
assign c2441 =  x26;
assign c2443 = ~x33 & ~x54 & ~x270 & ~x379 & ~x408 & ~x435 & ~x464 & ~x493 & ~x648 & ~x671 & ~x701 & ~x702 & ~x731 & ~x755 & ~x759 & ~x764 & ~x767;
assign c2445 = ~x2 & ~x5 & ~x6 & ~x22 & ~x25 & ~x29 & ~x33 & ~x34 & ~x49 & ~x58 & ~x61 & ~x62 & ~x77 & ~x80 & ~x85 & ~x89 & ~x113 & ~x114 & ~x116 & ~x133 & ~x143 & ~x145 & ~x162 & ~x165 & ~x174 & ~x190 & ~x199 & ~x200 & ~x222 & ~x225 & ~x227 & ~x228 & ~x231 & ~x246 & ~x250 & ~x255 & ~x258 & ~x275 & ~x276 & ~x280 & ~x283 & ~x302 & ~x304 & ~x310 & ~x312 & ~x314 & ~x331 & ~x334 & ~x337 & ~x339 & ~x358 & ~x367 & ~x390 & ~x395 & ~x422 & ~x423 & ~x424 & ~x427 & ~x428 & ~x444 & ~x448 & ~x453 & ~x455 & ~x458 & ~x459 & ~x460 & ~x472 & ~x475 & ~x476 & ~x477 & ~x481 & ~x483 & ~x484 & ~x485 & ~x486 & ~x500 & ~x508 & ~x510 & ~x528 & ~x529 & ~x530 & ~x534 & ~x536 & ~x537 & ~x556 & ~x559 & ~x562 & ~x582 & ~x588 & ~x593 & ~x609 & ~x610 & ~x612 & ~x645 & ~x649 & ~x667 & ~x668 & ~x671 & ~x672 & ~x697 & ~x700 & ~x702 & ~x721 & ~x724 & ~x730 & ~x750 & ~x762 & ~x763 & ~x764 & ~x779 & ~x781 & ~x783;
assign c2449 =  x638 &  x731;
assign c2451 = ~x18 & ~x47 & ~x52 & ~x68 & ~x72 & ~x95 & ~x105 & ~x212 & ~x365 & ~x393 & ~x419 & ~x450 & ~x749 & ~x750 & ~x753 & ~x761;
assign c2453 =  x553;
assign c2455 = ~x49 & ~x59 & ~x76 & ~x88 & ~x109 & ~x115 & ~x144 & ~x193 & ~x220 & ~x226 & ~x228 & ~x277 & ~x308 & ~x313 & ~x340 & ~x342 & ~x368 & ~x372 & ~x399 & ~x401 & ~x402 & ~x403 & ~x454 & ~x456 & ~x504 & ~x507 & ~x556 & ~x592 & ~x616 & ~x641 & ~x672 & ~x737;
assign c2457 =  x0;
assign c2459 =  x150 &  x233 & ~x352;
assign c2461 =  x624 & ~x456 & ~x479 & ~x510;
assign c2463 =  x112;
assign c2465 = ~x49 & ~x164 & ~x171 & ~x232 & ~x261 & ~x284 & ~x339 & ~x352 & ~x353 & ~x437 & ~x465 & ~x522 & ~x698 & ~x765;
assign c2467 =  x482 & ~x450 & ~x477 & ~x542 & ~x596 & ~x597 & ~x624;
assign c2469 = ~x21 & ~x65 & ~x79 & ~x81 & ~x111 & ~x227 & ~x247 & ~x489 & ~x515 & ~x538 & ~x569 & ~x570 & ~x595 & ~x734 & ~x758 & ~x779;
assign c2471 =  x503;
assign c2473 =  x619 & ~x365 & ~x421 & ~x449 & ~x569 & ~x625 & ~x681;
assign c2475 =  x700;
assign c2477 = ~x4 & ~x25 & ~x82 & ~x85 & ~x102 & ~x138 & ~x158 & ~x222 & ~x246 & ~x255 & ~x277 & ~x308 & ~x332 & ~x345 & ~x346 & ~x372 & ~x417 & ~x426 & ~x484 & ~x533 & ~x588 & ~x614 & ~x621 & ~x637 & ~x673 & ~x732 & ~x765;
assign c2479 = ~x4 & ~x20 & ~x25 & ~x53 & ~x64 & ~x87 & ~x89 & ~x105 & ~x108 & ~x109 & ~x111 & ~x137 & ~x143 & ~x145 & ~x148 & ~x149 & ~x160 & ~x163 & ~x164 & ~x166 & ~x172 & ~x220 & ~x231 & ~x278 & ~x279 & ~x287 & ~x290 & ~x305 & ~x307 & ~x313 & ~x316 & ~x317 & ~x331 & ~x332 & ~x336 & ~x342 & ~x362 & ~x371 & ~x393 & ~x418 & ~x427 & ~x442 & ~x444 & ~x445 & ~x451 & ~x467 & ~x469 & ~x471 & ~x474 & ~x479 & ~x480 & ~x498 & ~x531 & ~x553 & ~x559 & ~x585 & ~x610 & ~x614 & ~x619 & ~x640 & ~x672 & ~x727 & ~x728 & ~x734 & ~x754 & ~x761;
assign c2481 =  x351 & ~x101 & ~x129 & ~x185 & ~x219 & ~x245 & ~x272 & ~x363;
assign c2483 =  x295 &  x408 & ~x47 & ~x78 & ~x102 & ~x103 & ~x133 & ~x137 & ~x168 & ~x217 & ~x222 & ~x227 & ~x229 & ~x306 & ~x341 & ~x363 & ~x397 & ~x425 & ~x537 & ~x586 & ~x592 & ~x702 & ~x783;
assign c2485 = ~x75 & ~x106 & ~x132 & ~x189 & ~x246 & ~x318 & ~x400 & ~x401 & ~x482 & ~x588 & ~x638 & ~x714 & ~x763;
assign c2487 =  x0 &  x783;
assign c2489 =  x718 & ~x286 & ~x325 & ~x354 & ~x440 & ~x442 & ~x466 & ~x495;
assign c2491 = ~x2 & ~x29 & ~x32 & ~x53 & ~x58 & ~x77 & ~x85 & ~x86 & ~x90 & ~x116 & ~x132 & ~x139 & ~x143 & ~x160 & ~x162 & ~x164 & ~x197 & ~x199 & ~x202 & ~x218 & ~x229 & ~x230 & ~x248 & ~x256 & ~x257 & ~x273 & ~x285 & ~x304 & ~x305 & ~x306 & ~x312 & ~x313 & ~x336 & ~x344 & ~x365 & ~x369 & ~x371 & ~x372 & ~x387 & ~x401 & ~x402 & ~x403 & ~x420 & ~x425 & ~x442 & ~x444 & ~x445 & ~x450 & ~x452 & ~x475 & ~x479 & ~x481 & ~x483 & ~x484 & ~x500 & ~x505 & ~x506 & ~x527 & ~x560 & ~x583 & ~x593 & ~x613 & ~x615 & ~x619 & ~x636 & ~x645 & ~x677 & ~x698 & ~x720 & ~x735 & ~x750 & ~x759 & ~x781;
assign c2493 = ~x1 & ~x26 & ~x29 & ~x30 & ~x31 & ~x52 & ~x53 & ~x55 & ~x57 & ~x58 & ~x59 & ~x76 & ~x77 & ~x79 & ~x81 & ~x92 & ~x105 & ~x114 & ~x116 & ~x117 & ~x118 & ~x120 & ~x139 & ~x144 & ~x148 & ~x163 & ~x164 & ~x165 & ~x168 & ~x191 & ~x193 & ~x196 & ~x198 & ~x201 & ~x219 & ~x221 & ~x222 & ~x224 & ~x225 & ~x227 & ~x229 & ~x230 & ~x247 & ~x249 & ~x250 & ~x253 & ~x255 & ~x256 & ~x257 & ~x274 & ~x275 & ~x276 & ~x277 & ~x278 & ~x280 & ~x281 & ~x288 & ~x303 & ~x313 & ~x314 & ~x330 & ~x336 & ~x340 & ~x341 & ~x343 & ~x358 & ~x361 & ~x365 & ~x366 & ~x371 & ~x387 & ~x394 & ~x398 & ~x399 & ~x421 & ~x423 & ~x428 & ~x446 & ~x447 & ~x448 & ~x453 & ~x454 & ~x473 & ~x480 & ~x502 & ~x504 & ~x528 & ~x529 & ~x533 & ~x534 & ~x536 & ~x558 & ~x559 & ~x560 & ~x563 & ~x585 & ~x587 & ~x588 & ~x590 & ~x591 & ~x611 & ~x612 & ~x613 & ~x614 & ~x616 & ~x617 & ~x639 & ~x640 & ~x646 & ~x668 & ~x670 & ~x697 & ~x700 & ~x724 & ~x726 & ~x727 & ~x729 & ~x733 & ~x754 & ~x756 & ~x760 & ~x761 & ~x765 & ~x779;
assign c2495 =  x333;
assign c2497 =  x314 & ~x14 & ~x264 & ~x514;
assign c2499 =  x390;
assign c30 =  x211 &  x498 & ~x300 & ~x406 & ~x433 & ~x461 & ~x488 & ~x589 & ~x616;
assign c32 = ~x98 & ~x109 & ~x389 & ~x493 & ~x520 & ~x534 & ~x572 & ~x573 & ~x596 & ~x704 & ~x705 & ~x733;
assign c34 = ~x1 & ~x12 & ~x19 & ~x23 & ~x26 & ~x28 & ~x30 & ~x49 & ~x55 & ~x67 & ~x68 & ~x88 & ~x109 & ~x111 & ~x115 & ~x134 & ~x194 & ~x198 & ~x220 & ~x225 & ~x281 & ~x335 & ~x391 & ~x392 & ~x395 & ~x415 & ~x416 & ~x417 & ~x418 & ~x419 & ~x443 & ~x448 & ~x471 & ~x472 & ~x532 & ~x533 & ~x559 & ~x560 & ~x572 & ~x612 & ~x613 & ~x640 & ~x646 & ~x668 & ~x669 & ~x697 & ~x698 & ~x703 & ~x711 & ~x724 & ~x726 & ~x731 & ~x751;
assign c36 =  x157 &  x158 &  x186 & ~x27 & ~x38 & ~x39 & ~x56 & ~x83 & ~x85 & ~x123 & ~x140 & ~x141 & ~x167 & ~x170 & ~x221 & ~x250 & ~x251 & ~x253 & ~x279 & ~x306 & ~x308 & ~x392 & ~x474 & ~x476 & ~x502 & ~x557 & ~x642 & ~x701 & ~x757;
assign c38 = ~x0 & ~x12 & ~x85 & ~x196 & ~x197 & ~x224 & ~x291 & ~x292 & ~x375 & ~x392 & ~x398 & ~x445 & ~x446 & ~x457 & ~x481 & ~x513 & ~x568 & ~x569 & ~x596 & ~x616 & ~x643 & ~x717;
assign c310 = ~x110 & ~x318 & ~x369 & ~x377 & ~x378 & ~x407 & ~x434 & ~x461 & ~x489 & ~x504 & ~x533 & ~x661 & ~x688;
assign c312 =  x692 & ~x53 & ~x86 & ~x110 & ~x139 & ~x224 & ~x225 & ~x249 & ~x251 & ~x277 & ~x282 & ~x306 & ~x307 & ~x308 & ~x309 & ~x391 & ~x532 & ~x587 & ~x603 & ~x630 & ~x659 & ~x660 & ~x670 & ~x696 & ~x700 & ~x703 & ~x727 & ~x753;
assign c314 =  x662 & ~x21 & ~x23 & ~x27 & ~x112 & ~x139 & ~x166 & ~x195 & ~x249 & ~x278 & ~x334 & ~x486 & ~x514 & ~x544 & ~x600 & ~x630 & ~x669 & ~x726 & ~x777 & ~x779;
assign c316 = ~x274 & ~x358 & ~x380 & ~x381 & ~x384 & ~x399 & ~x405 & ~x410 & ~x411 & ~x439 & ~x453;
assign c318 = ~x82 & ~x85 & ~x86 & ~x114 & ~x138 & ~x141 & ~x142 & ~x167 & ~x195 & ~x250 & ~x251 & ~x254 & ~x262 & ~x281 & ~x418 & ~x446 & ~x447 & ~x474 & ~x491 & ~x506 & ~x531 & ~x540 & ~x561 & ~x562 & ~x588 & ~x596 & ~x615 & ~x616 & ~x617 & ~x645 & ~x647 & ~x670 & ~x700 & ~x730 & ~x747 & ~x754 & ~x783;
assign c320 = ~x30 & ~x322 & ~x323 & ~x325 & ~x348 & ~x379 & ~x381 & ~x432 & ~x460 & ~x478 & ~x488 & ~x507 & ~x532 & ~x535 & ~x565 & ~x587 & ~x666 & ~x692 & ~x697 & ~x723 & ~x777;
assign c322 =  x323 & ~x24 & ~x85 & ~x86 & ~x308 & ~x410 & ~x438 & ~x463 & ~x466 & ~x493 & ~x494 & ~x517 & ~x519 & ~x520 & ~x547 & ~x572 & ~x575 & ~x629 & ~x656 & ~x700;
assign c324 = ~x7 & ~x25 & ~x38 & ~x42 & ~x114 & ~x141 & ~x151 & ~x168 & ~x206 & ~x226 & ~x233 & ~x282 & ~x337 & ~x343 & ~x371 & ~x390 & ~x419 & ~x447 & ~x462 & ~x503 & ~x531 & ~x546 & ~x559 & ~x603 & ~x614 & ~x727;
assign c326 = ~x92 & ~x147 & ~x162 & ~x250 & ~x279 & ~x450 & ~x464 & ~x471 & ~x615 & ~x618 & ~x640 & ~x707 & ~x709 & ~x730;
assign c328 = ~x6 & ~x56 & ~x60 & ~x83 & ~x112 & ~x172 & ~x199 & ~x223 & ~x226 & ~x253 & ~x358 & ~x437 & ~x442 & ~x463 & ~x493 & ~x681 & ~x683 & ~x685 & ~x707 & ~x708 & ~x761 & ~x762;
assign c330 = ~x2 & ~x15 & ~x81 & ~x141 & ~x251 & ~x407 & ~x408 & ~x459 & ~x462 & ~x465 & ~x491 & ~x514 & ~x542 & ~x562 & ~x587 & ~x618 & ~x646 & ~x649 & ~x652 & ~x754 & ~x757 & ~x758;
assign c332 =  x240 &  x267 & ~x1 & ~x82 & ~x139 & ~x289 & ~x344 & ~x404 & ~x428 & ~x455 & ~x484;
assign c334 = ~x53 & ~x385 & ~x411 & ~x413 & ~x441 & ~x467 & ~x468 & ~x510 & ~x561 & ~x598 & ~x599;
assign c336 =  x257 & ~x6 & ~x12 & ~x26 & ~x37 & ~x39 & ~x50 & ~x67 & ~x68 & ~x81 & ~x94 & ~x111 & ~x112 & ~x114 & ~x122 & ~x139 & ~x140 & ~x142 & ~x143 & ~x166 & ~x167 & ~x170 & ~x171 & ~x198 & ~x199 & ~x392 & ~x448 & ~x476 & ~x504 & ~x515 & ~x531 & ~x532 & ~x543 & ~x559 & ~x560 & ~x588 & ~x616 & ~x627 & ~x642 & ~x671 & ~x700 & ~x729 & ~x755 & ~x756 & ~x757 & ~x759;
assign c338 = ~x0 & ~x5 & ~x7 & ~x25 & ~x37 & ~x134 & ~x135 & ~x139 & ~x220 & ~x221 & ~x246 & ~x247 & ~x250 & ~x278 & ~x306 & ~x308 & ~x448 & ~x520 & ~x548 & ~x574 & ~x604 & ~x615 & ~x643 & ~x670 & ~x683 & ~x685 & ~x709 & ~x724 & ~x737 & ~x753 & ~x757 & ~x781 & ~x783;
assign c340 =  x71 &  x72 & ~x167 & ~x207 & ~x236 & ~x262 & ~x263 & ~x430;
assign c342 = ~x60 & ~x85 & ~x115 & ~x381 & ~x405 & ~x435 & ~x462 & ~x503 & ~x537 & ~x565 & ~x594 & ~x595 & ~x644 & ~x679 & ~x718 & ~x747 & ~x754 & ~x772 & ~x774 & ~x783;
assign c344 = ~x53 & ~x243 & ~x402 & ~x409 & ~x423 & ~x436 & ~x490 & ~x532 & ~x589 & ~x674;
assign c346 =  x749 & ~x196 & ~x271 & ~x299 & ~x336 & ~x420 & ~x550;
assign c348 =  x306 &  x334 & ~x330 & ~x354 & ~x359 & ~x387 & ~x414 & ~x439 & ~x440 & ~x441 & ~x458 & ~x469 & ~x485 & ~x568;
assign c350 =  x270 & ~x55 & ~x80 & ~x81 & ~x114 & ~x140 & ~x195 & ~x223 & ~x224 & ~x226 & ~x252 & ~x335 & ~x361 & ~x363 & ~x402 & ~x486 & ~x501 & ~x542 & ~x548 & ~x587 & ~x598 & ~x616 & ~x642 & ~x672 & ~x724 & ~x729 & ~x782;
assign c352 = ~x6 & ~x7 & ~x8 & ~x35 & ~x54 & ~x139 & ~x381 & ~x408 & ~x431 & ~x464 & ~x570 & ~x595 & ~x624 & ~x625 & ~x626 & ~x652 & ~x672 & ~x727 & ~x728;
assign c354 =  x192 &  x221 &  x305 & ~x349 & ~x376 & ~x403 & ~x645;
assign c356 = ~x27 & ~x30 & ~x58 & ~x416 & ~x461 & ~x464 & ~x526 & ~x553 & ~x554 & ~x566 & ~x648 & ~x728 & ~x749;
assign c358 =  x497 & ~x438 & ~x462 & ~x486 & ~x542 & ~x588 & ~x595 & ~x724 & ~x778;
assign c360 = ~x60 & ~x61 & ~x114 & ~x141 & ~x197 & ~x358 & ~x385 & ~x386 & ~x409 & ~x414 & ~x440 & ~x467 & ~x469 & ~x486 & ~x494 & ~x512 & ~x595 & ~x616 & ~x620 & ~x644 & ~x723 & ~x727 & ~x729 & ~x739 & ~x740 & ~x749 & ~x760 & ~x772;
assign c362 =  x276 & ~x27 & ~x56 & ~x354 & ~x392 & ~x407 & ~x432 & ~x436 & ~x448 & ~x458 & ~x459 & ~x461 & ~x560 & ~x616 & ~x645 & ~x646 & ~x701 & ~x729 & ~x756;
assign c364 =  x453 &  x481 & ~x21 & ~x28 & ~x51 & ~x54 & ~x56 & ~x58 & ~x86 & ~x108 & ~x109 & ~x110 & ~x114 & ~x139 & ~x164 & ~x167 & ~x168 & ~x169 & ~x193 & ~x194 & ~x221 & ~x224 & ~x250 & ~x276 & ~x278 & ~x282 & ~x308 & ~x309 & ~x310 & ~x334 & ~x365 & ~x417 & ~x419 & ~x449 & ~x475 & ~x502 & ~x516 & ~x530 & ~x531 & ~x533 & ~x558 & ~x561 & ~x572 & ~x585 & ~x586 & ~x589 & ~x590 & ~x617 & ~x642 & ~x644 & ~x668 & ~x669 & ~x673 & ~x674 & ~x699 & ~x726 & ~x729 & ~x732 & ~x754 & ~x756 & ~x760 & ~x783;
assign c366 =  x611 & ~x0 & ~x4 & ~x54 & ~x61 & ~x112 & ~x195 & ~x307 & ~x495 & ~x496 & ~x521 & ~x548 & ~x599 & ~x600 & ~x643 & ~x654 & ~x736;
assign c368 = ~x3 & ~x60 & ~x114 & ~x172 & ~x275 & ~x360 & ~x436 & ~x462 & ~x463 & ~x479 & ~x519 & ~x545 & ~x547 & ~x601 & ~x673 & ~x680 & ~x703;
assign c370 =  x265 & ~x27 & ~x57 & ~x61 & ~x62 & ~x72 & ~x85 & ~x89 & ~x98 & ~x113 & ~x114 & ~x139 & ~x308 & ~x354 & ~x436 & ~x437 & ~x462 & ~x465 & ~x646 & ~x755 & ~x758 & ~x783;
assign c372 =  x314 &  x342 & ~x2 & ~x9 & ~x29 & ~x31 & ~x53 & ~x59 & ~x86 & ~x107 & ~x111 & ~x139 & ~x165 & ~x166 & ~x167 & ~x194 & ~x197 & ~x199 & ~x223 & ~x224 & ~x228 & ~x251 & ~x255 & ~x278 & ~x284 & ~x308 & ~x310 & ~x312 & ~x336 & ~x363 & ~x365 & ~x366 & ~x393 & ~x419 & ~x474 & ~x478 & ~x533 & ~x557 & ~x559 & ~x641 & ~x642 & ~x644 & ~x645 & ~x670 & ~x671 & ~x672 & ~x674 & ~x698 & ~x701 & ~x730 & ~x739 & ~x759 & ~x782 & ~x783;
assign c374 =  x740 & ~x6 & ~x319 & ~x375 & ~x403 & ~x487;
assign c376 = ~x22 & ~x23 & ~x352 & ~x353 & ~x379 & ~x381 & ~x395 & ~x407 & ~x435 & ~x451 & ~x452 & ~x509 & ~x532 & ~x563 & ~x566 & ~x706 & ~x780;
assign c378 =  x611 & ~x111 & ~x238 & ~x485 & ~x532 & ~x550 & ~x626;
assign c380 = ~x54 & ~x119 & ~x174 & ~x204 & ~x286 & ~x313 & ~x341 & ~x542 & ~x575 & ~x677 & ~x681 & ~x707 & ~x729 & ~x735 & ~x760;
assign c382 =  x302 & ~x29 & ~x109 & ~x140 & ~x165 & ~x221 & ~x222 & ~x223 & ~x224 & ~x251 & ~x253 & ~x317 & ~x334 & ~x363 & ~x446 & ~x448 & ~x463 & ~x473 & ~x475 & ~x490 & ~x501 & ~x586 & ~x613 & ~x674 & ~x726 & ~x729 & ~x730;
assign c384 =  x380 &  x534 &  x562 & ~x56 & ~x168 & ~x195 & ~x281 & ~x307 & ~x516 & ~x570 & ~x654;
assign c386 =  x268 &  x269 &  x295 & ~x47 & ~x140 & ~x169 & ~x252 & ~x385 & ~x440 & ~x460 & ~x468 & ~x488 & ~x517 & ~x544 & ~x545 & ~x700 & ~x701 & ~x729;
assign c388 =  x501 & ~x3 & ~x30 & ~x33 & ~x34 & ~x56 & ~x58 & ~x114 & ~x115 & ~x117 & ~x141 & ~x142 & ~x143 & ~x145 & ~x170 & ~x171 & ~x173 & ~x196 & ~x200 & ~x227 & ~x228 & ~x252 & ~x255 & ~x280 & ~x282 & ~x309 & ~x469 & ~x494 & ~x495 & ~x496 & ~x523 & ~x547 & ~x575 & ~x599;
assign c390 = ~x6 & ~x22 & ~x39 & ~x55 & ~x63 & ~x64 & ~x82 & ~x108 & ~x110 & ~x113 & ~x138 & ~x149 & ~x152 & ~x166 & ~x178 & ~x193 & ~x206 & ~x233 & ~x234 & ~x251 & ~x289 & ~x319 & ~x334 & ~x335 & ~x389 & ~x417 & ~x447 & ~x475 & ~x504 & ~x751 & ~x755 & ~x756 & ~x779 & ~x781 & ~x783;
assign c392 =  x327 &  x353 &  x355 &  x480 & ~x22 & ~x109 & ~x170 & ~x193 & ~x199 & ~x253 & ~x279 & ~x282 & ~x308 & ~x391 & ~x393;
assign c394 = ~x4 & ~x7 & ~x8 & ~x9 & ~x63 & ~x64 & ~x89 & ~x115 & ~x300 & ~x353 & ~x379 & ~x483 & ~x562 & ~x613 & ~x689 & ~x699 & ~x716;
assign c396 =  x267 &  x566 & ~x196 & ~x252 & ~x403 & ~x420 & ~x542 & ~x543 & ~x681 & ~x701 & ~x729;
assign c398 =  x473 & ~x27 & ~x59 & ~x85 & ~x116 & ~x245 & ~x246 & ~x273 & ~x274 & ~x301 & ~x521 & ~x522 & ~x547 & ~x653 & ~x738;
assign c3100 = ~x37 & ~x52 & ~x79 & ~x82 & ~x133 & ~x141 & ~x167 & ~x181 & ~x197 & ~x225 & ~x277 & ~x308 & ~x375 & ~x387 & ~x389 & ~x418 & ~x502 & ~x504 & ~x533 & ~x626 & ~x641 & ~x645 & ~x655 & ~x695 & ~x697 & ~x709 & ~x721 & ~x750 & ~x753 & ~x783;
assign c3102 = ~x278 & ~x299 & ~x306 & ~x455 & ~x464 & ~x465 & ~x468 & ~x491 & ~x549 & ~x588 & ~x757;
assign c3104 =  x663 & ~x5 & ~x6 & ~x60 & ~x85 & ~x107 & ~x114 & ~x135 & ~x166 & ~x168 & ~x191 & ~x224 & ~x307 & ~x476 & ~x574 & ~x588 & ~x627 & ~x683 & ~x725 & ~x729 & ~x782;
assign c3106 = ~x0 & ~x1 & ~x3 & ~x57 & ~x58 & ~x78 & ~x85 & ~x86 & ~x97 & ~x197 & ~x250 & ~x281 & ~x364 & ~x404 & ~x419 & ~x433 & ~x445 & ~x476 & ~x501 & ~x502 & ~x518 & ~x528 & ~x532 & ~x547 & ~x572 & ~x573 & ~x584 & ~x585 & ~x588 & ~x600 & ~x612 & ~x682 & ~x698 & ~x700 & ~x726 & ~x757 & ~x780;
assign c3108 =  x250 & ~x378 & ~x405 & ~x425;
assign c3110 = ~x7 & ~x31 & ~x52 & ~x54 & ~x98 & ~x190 & ~x254 & ~x303 & ~x339 & ~x362 & ~x396 & ~x445 & ~x473 & ~x474 & ~x501 & ~x529 & ~x555 & ~x562 & ~x591 & ~x641 & ~x649 & ~x734 & ~x751 & ~x759;
assign c3112 =  x102 &  x185 &  x622 &  x678 & ~x27 & ~x139 & ~x277 & ~x281 & ~x364 & ~x501 & ~x528 & ~x586 & ~x700 & ~x712 & ~x755;
assign c3114 =  x246 &  x422 & ~x0 & ~x1 & ~x23 & ~x26 & ~x27 & ~x52 & ~x53 & ~x54 & ~x57 & ~x84 & ~x110 & ~x111 & ~x168 & ~x195 & ~x224 & ~x252 & ~x432 & ~x458 & ~x461 & ~x462 & ~x463 & ~x486 & ~x489 & ~x490 & ~x491 & ~x514 & ~x517 & ~x531 & ~x559 & ~x615 & ~x616 & ~x700 & ~x727 & ~x729 & ~x757 & ~x783;
assign c3116 =  x258 & ~x40 & ~x144 & ~x195 & ~x248 & ~x505 & ~x560 & ~x589 & ~x673 & ~x702 & ~x722 & ~x724 & ~x755;
assign c3118 =  x380 &  x407 &  x691 & ~x112 & ~x114 & ~x166 & ~x307 & ~x333 & ~x628 & ~x655 & ~x684 & ~x739;
assign c3120 = ~x2 & ~x3 & ~x4 & ~x30 & ~x31 & ~x32 & ~x39 & ~x83 & ~x84 & ~x264 & ~x265 & ~x291 & ~x292 & ~x320 & ~x345 & ~x347 & ~x348 & ~x404 & ~x422 & ~x429 & ~x431 & ~x475 & ~x476 & ~x503 & ~x531 & ~x532 & ~x558 & ~x559 & ~x560 & ~x561 & ~x588 & ~x670 & ~x672 & ~x724 & ~x727 & ~x753 & ~x754 & ~x755 & ~x774;
assign c3122 =  x260 & ~x2 & ~x6 & ~x35 & ~x54 & ~x227 & ~x228 & ~x406 & ~x489 & ~x504 & ~x557 & ~x589 & ~x590 & ~x591 & ~x640 & ~x643 & ~x672 & ~x722 & ~x752 & ~x757;
assign c3124 =  x334 & ~x52 & ~x59 & ~x354 & ~x356 & ~x382 & ~x385 & ~x412 & ~x434 & ~x438 & ~x485 & ~x513 & ~x566 & ~x746 & ~x764 & ~x778;
assign c3126 =  x287 &  x370 & ~x226 & ~x305 & ~x368 & ~x395 & ~x423 & ~x648 & ~x705;
assign c3128 =  x397 &  x508 &  x536 & ~x33 & ~x55 & ~x194 & ~x198 & ~x281 & ~x393 & ~x394 & ~x412 & ~x474 & ~x477 & ~x491 & ~x533 & ~x586 & ~x588 & ~x673;
assign c3130 =  x324 & ~x78 & ~x111 & ~x194 & ~x223 & ~x318 & ~x346 & ~x373 & ~x516 & ~x549 & ~x559 & ~x572 & ~x588 & ~x700 & ~x757;
assign c3132 = ~x1 & ~x57 & ~x141 & ~x357 & ~x385 & ~x411 & ~x435 & ~x439 & ~x441 & ~x490 & ~x493 & ~x495 & ~x522 & ~x548 & ~x575 & ~x628 & ~x654 & ~x708 & ~x709 & ~x710 & ~x775;
assign c3134 =  x331 &  x695 & ~x504 & ~x587;
assign c3136 = ~x1 & ~x3 & ~x5 & ~x57 & ~x84 & ~x85 & ~x145 & ~x169 & ~x170 & ~x171 & ~x226 & ~x227 & ~x228 & ~x255 & ~x283 & ~x308 & ~x336 & ~x440 & ~x468 & ~x492 & ~x494 & ~x495 & ~x521 & ~x522 & ~x548 & ~x575 & ~x597 & ~x600 & ~x601 & ~x602 & ~x625 & ~x627 & ~x628 & ~x630 & ~x651 & ~x654 & ~x655 & ~x656 & ~x658 & ~x679 & ~x680 & ~x681 & ~x682 & ~x683 & ~x707 & ~x708 & ~x734 & ~x762;
assign c3138 = ~x53 & ~x56 & ~x83 & ~x166 & ~x271 & ~x299 & ~x350 & ~x355 & ~x377 & ~x466 & ~x477 & ~x495 & ~x503 & ~x505 & ~x518 & ~x586 & ~x589 & ~x617 & ~x698 & ~x780 & ~x783;
assign c3140 =  x417 & ~x217 & ~x245 & ~x246 & ~x299 & ~x302 & ~x449 & ~x486 & ~x514 & ~x542 & ~x595 & ~x596 & ~x699 & ~x727;
assign c3142 = ~x7 & ~x35 & ~x78 & ~x197 & ~x306 & ~x464 & ~x504 & ~x516 & ~x521 & ~x533 & ~x575 & ~x656 & ~x701 & ~x707 & ~x708 & ~x709 & ~x736;
assign c3144 =  x331 & ~x0 & ~x177 & ~x195 & ~x293 & ~x321 & ~x348 & ~x473 & ~x474 & ~x503 & ~x716;
assign c3146 =  x187 & ~x11 & ~x39 & ~x65 & ~x95 & ~x125 & ~x142 & ~x151 & ~x197 & ~x233 & ~x250 & ~x261 & ~x293 & ~x306 & ~x316 & ~x446 & ~x503 & ~x572 & ~x783;
assign c3148 = ~x6 & ~x27 & ~x52 & ~x60 & ~x63 & ~x79 & ~x82 & ~x86 & ~x87 & ~x89 & ~x91 & ~x110 & ~x142 & ~x144 & ~x145 & ~x146 & ~x162 & ~x163 & ~x171 & ~x172 & ~x188 & ~x190 & ~x193 & ~x212 & ~x221 & ~x228 & ~x251 & ~x308 & ~x521 & ~x545 & ~x575 & ~x601 & ~x626 & ~x629 & ~x651 & ~x653 & ~x657 & ~x678 & ~x707 & ~x709 & ~x733 & ~x760;
assign c3150 =  x44 &  x100 & ~x38 & ~x52 & ~x196 & ~x292 & ~x519 & ~x631 & ~x710 & ~x711;
assign c3152 = ~x34 & ~x56 & ~x111 & ~x138 & ~x142 & ~x151 & ~x164 & ~x167 & ~x180 & ~x182 & ~x194 & ~x195 & ~x196 & ~x309 & ~x317 & ~x362 & ~x363 & ~x373 & ~x415 & ~x473 & ~x475 & ~x499 & ~x543 & ~x560 & ~x729 & ~x783;
assign c3154 = ~x96 & ~x143 & ~x409 & ~x434 & ~x460 & ~x511 & ~x530 & ~x533 & ~x539 & ~x590 & ~x662 & ~x689;
assign c3156 = ~x23 & ~x270 & ~x407 & ~x421 & ~x452 & ~x477 & ~x478 & ~x531 & ~x561 & ~x562 & ~x640 & ~x678 & ~x679 & ~x727 & ~x730 & ~x731 & ~x762;
assign c3158 =  x185 & ~x1 & ~x2 & ~x4 & ~x9 & ~x23 & ~x24 & ~x27 & ~x31 & ~x56 & ~x67 & ~x78 & ~x83 & ~x84 & ~x109 & ~x111 & ~x137 & ~x166 & ~x167 & ~x196 & ~x197 & ~x223 & ~x224 & ~x249 & ~x251 & ~x266 & ~x280 & ~x307 & ~x308 & ~x337 & ~x419 & ~x420 & ~x447 & ~x473 & ~x475 & ~x476 & ~x502 & ~x504 & ~x516 & ~x544 & ~x558 & ~x559 & ~x587 & ~x588 & ~x628 & ~x671 & ~x699 & ~x700 & ~x757 & ~x782;
assign c3160 =  x157 &  x268 & ~x20 & ~x41 & ~x109 & ~x151 & ~x222 & ~x224 & ~x445 & ~x502 & ~x530 & ~x586 & ~x588 & ~x616 & ~x642 & ~x669 & ~x670 & ~x758;
assign c3162 =  x360 &  x388 &  x416 &  x444 & ~x1 & ~x57 & ~x465 & ~x491 & ~x492 & ~x493 & ~x494 & ~x504 & ~x516 & ~x520 & ~x521 & ~x531 & ~x532 & ~x547 & ~x548 & ~x701 & ~x728 & ~x756;
assign c3164 = ~x42 & ~x377 & ~x409 & ~x432 & ~x433 & ~x464 & ~x475 & ~x491 & ~x506 & ~x518 & ~x536 & ~x537 & ~x562 & ~x585 & ~x586 & ~x594 & ~x644 & ~x666 & ~x727;
assign c3166 =  x474 & ~x0 & ~x16 & ~x28 & ~x56 & ~x57 & ~x58 & ~x63 & ~x89 & ~x112 & ~x117 & ~x470 & ~x485 & ~x495 & ~x539 & ~x566 & ~x567 & ~x594 & ~x595 & ~x597 & ~x623 & ~x767 & ~x773;
assign c3168 =  x219 & ~x206 & ~x234 & ~x261 & ~x288 & ~x306 & ~x343 & ~x427;
assign c3170 =  x501 & ~x27 & ~x58 & ~x84 & ~x86 & ~x169 & ~x274 & ~x301 & ~x302 & ~x551 & ~x569 & ~x570 & ~x596 & ~x597 & ~x625 & ~x679 & ~x680 & ~x682 & ~x736;
assign c3172 =  x479 &  x720 & ~x67 & ~x122 & ~x287;
assign c3174 =  x324 & ~x13 & ~x111 & ~x135 & ~x137 & ~x140 & ~x195 & ~x198 & ~x223 & ~x253 & ~x335 & ~x486 & ~x514 & ~x546 & ~x574 & ~x616 & ~x631 & ~x657 & ~x658 & ~x685 & ~x710 & ~x728 & ~x729 & ~x765 & ~x766;
assign c3176 =  x323 &  x636 & ~x38 & ~x79 & ~x109 & ~x420 & ~x545 & ~x573 & ~x587 & ~x600 & ~x601 & ~x628 & ~x701;
assign c3178 =  x713 & ~x381 & ~x408 & ~x434 & ~x436 & ~x462 & ~x490 & ~x491 & ~x518 & ~x542 & ~x626;
assign c3180 =  x585 & ~x440 & ~x442 & ~x497 & ~x552 & ~x554 & ~x570 & ~x579 & ~x581 & ~x608 & ~x625 & ~x681;
assign c3182 =  x332 &  x360 & ~x83 & ~x273 & ~x301 & ~x436 & ~x437 & ~x459 & ~x462 & ~x477 & ~x490 & ~x646;
assign c3184 = ~x2 & ~x9 & ~x11 & ~x37 & ~x39 & ~x67 & ~x152 & ~x180 & ~x233 & ~x237 & ~x277 & ~x279 & ~x419 & ~x432 & ~x460 & ~x476 & ~x501 & ~x531 & ~x557 & ~x673 & ~x757 & ~x782;
assign c3186 = ~x28 & ~x37 & ~x83 & ~x108 & ~x110 & ~x138 & ~x249 & ~x252 & ~x253 & ~x310 & ~x311 & ~x335 & ~x390 & ~x405 & ~x473 & ~x533 & ~x539 & ~x567 & ~x580 & ~x608;
assign c3188 = ~x16 & ~x17 & ~x18 & ~x19 & ~x44 & ~x48 & ~x56 & ~x115 & ~x140 & ~x170 & ~x197 & ~x224 & ~x330 & ~x385 & ~x386 & ~x440 & ~x442 & ~x467 & ~x469 & ~x496 & ~x515 & ~x542 & ~x598 & ~x599 & ~x652 & ~x654 & ~x763;
assign c3190 =  x509 &  x537 & ~x117 & ~x173 & ~x199 & ~x438 & ~x466 & ~x549 & ~x615 & ~x702;
assign c3192 =  x352 &  x635 & ~x22 & ~x98 & ~x107 & ~x278 & ~x306 & ~x446 & ~x599;
assign c3194 =  x324 & ~x12 & ~x52 & ~x83 & ~x135 & ~x138 & ~x224 & ~x308 & ~x335 & ~x475 & ~x487 & ~x500 & ~x532 & ~x543 & ~x573 & ~x588 & ~x602 & ~x643 & ~x654 & ~x657 & ~x659 & ~x684 & ~x710 & ~x755 & ~x782;
assign c3196 = ~x3 & ~x25 & ~x51 & ~x82 & ~x325 & ~x351 & ~x353 & ~x380 & ~x405 & ~x432 & ~x502 & ~x529 & ~x531 & ~x532 & ~x533 & ~x559 & ~x584 & ~x586 & ~x588 & ~x589 & ~x616 & ~x641 & ~x674 & ~x701 & ~x705 & ~x716 & ~x753 & ~x754 & ~x755 & ~x783;
assign c3198 =  x474 & ~x23 & ~x31 & ~x58 & ~x199 & ~x227 & ~x442 & ~x443 & ~x469 & ~x495 & ~x541 & ~x542 & ~x623 & ~x729;
assign c3200 = ~x7 & ~x21 & ~x28 & ~x30 & ~x35 & ~x36 & ~x79 & ~x111 & ~x115 & ~x119 & ~x162 & ~x168 & ~x174 & ~x195 & ~x200 & ~x201 & ~x224 & ~x284 & ~x307 & ~x308 & ~x337 & ~x491 & ~x520 & ~x548 & ~x642 & ~x679 & ~x706 & ~x778 & ~x782;
assign c3202 =  x474 & ~x58 & ~x443 & ~x498 & ~x576 & ~x580;
assign c3204 =  x269 &  x296 &  x479 & ~x114 & ~x138 & ~x139 & ~x140 & ~x170 & ~x197 & ~x224 & ~x226 & ~x281 & ~x491 & ~x518 & ~x545 & ~x588 & ~x699;
assign c3206 = ~x0 & ~x4 & ~x24 & ~x26 & ~x50 & ~x58 & ~x78 & ~x191 & ~x192 & ~x224 & ~x363 & ~x433 & ~x461 & ~x462 & ~x474 & ~x490 & ~x492 & ~x502 & ~x530 & ~x533 & ~x545 & ~x560 & ~x561 & ~x584 & ~x612 & ~x615 & ~x617 & ~x626 & ~x627 & ~x674 & ~x695 & ~x697 & ~x709 & ~x729 & ~x781;
assign c3208 =  x221 &  x361 &  x501 & ~x83 & ~x302 & ~x384;
assign c3210 = ~x83 & ~x86 & ~x171 & ~x188 & ~x190 & ~x212 & ~x214 & ~x219 & ~x240 & ~x248 & ~x267 & ~x280 & ~x522 & ~x547 & ~x570 & ~x571 & ~x596 & ~x597 & ~x603 & ~x625 & ~x653 & ~x654 & ~x707 & ~x709;
assign c3212 =  x342 &  x453 & ~x0 & ~x21 & ~x28 & ~x32 & ~x54 & ~x55 & ~x59 & ~x82 & ~x83 & ~x113 & ~x114 & ~x140 & ~x143 & ~x165 & ~x170 & ~x193 & ~x195 & ~x196 & ~x199 & ~x200 & ~x224 & ~x225 & ~x249 & ~x253 & ~x277 & ~x282 & ~x283 & ~x309 & ~x311 & ~x363 & ~x364 & ~x389 & ~x392 & ~x418 & ~x421 & ~x445 & ~x472 & ~x475 & ~x479 & ~x507 & ~x528 & ~x534 & ~x560 & ~x589 & ~x591 & ~x615 & ~x616 & ~x617 & ~x672 & ~x702 & ~x725 & ~x729 & ~x755 & ~x756 & ~x779 & ~x781;
assign c3214 = ~x82 & ~x84 & ~x108 & ~x112 & ~x136 & ~x148 & ~x168 & ~x176 & ~x203 & ~x235 & ~x236 & ~x259 & ~x264 & ~x265 & ~x287 & ~x292 & ~x319 & ~x348 & ~x375 & ~x403 & ~x418 & ~x419 & ~x430 & ~x471 & ~x475 & ~x542 & ~x570 & ~x598;
assign c3216 =  x610 & ~x55 & ~x83 & ~x138 & ~x477 & ~x491 & ~x505 & ~x519 & ~x545 & ~x548 & ~x549 & ~x571 & ~x572 & ~x574 & ~x589 & ~x601 & ~x626 & ~x642 & ~x654 & ~x697 & ~x699 & ~x700 & ~x701 & ~x729 & ~x754;
assign c3218 =  x269 &  x295 & ~x1 & ~x19 & ~x28 & ~x29 & ~x57 & ~x111 & ~x135 & ~x142 & ~x159 & ~x226 & ~x254 & ~x280 & ~x459 & ~x460 & ~x515 & ~x560 & ~x574 & ~x614 & ~x643 & ~x729 & ~x730 & ~x757;
assign c3220 =  x160 & ~x72 & ~x86 & ~x197 & ~x234 & ~x336 & ~x504 & ~x577 & ~x587 & ~x628;
assign c3222 = ~x109 & ~x223 & ~x306 & ~x381 & ~x489 & ~x493 & ~x546 & ~x548 & ~x562 & ~x564 & ~x676 & ~x700 & ~x781;
assign c3224 =  x528 & ~x4 & ~x54 & ~x141 & ~x384 & ~x413 & ~x437 & ~x442 & ~x496 & ~x497 & ~x515;
assign c3226 =  x418 & ~x142 & ~x412 & ~x440 & ~x488 & ~x517 & ~x521 & ~x542 & ~x546 & ~x547;
assign c3228 =  x184 & ~x2 & ~x23 & ~x24 & ~x31 & ~x81 & ~x98 & ~x109 & ~x137 & ~x167 & ~x223 & ~x252 & ~x406 & ~x489 & ~x517 & ~x518 & ~x533 & ~x545 & ~x587 & ~x589 & ~x616 & ~x647 & ~x671 & ~x674 & ~x701 & ~x731 & ~x732;
assign c3230 =  x267 & ~x29 & ~x166 & ~x168 & ~x327 & ~x383 & ~x410 & ~x411 & ~x435 & ~x437 & ~x438 & ~x439 & ~x462 & ~x464 & ~x465 & ~x493 & ~x494 & ~x645 & ~x672 & ~x730 & ~x781 & ~x782;
assign c3232 = ~x5 & ~x8 & ~x66 & ~x77 & ~x78 & ~x80 & ~x82 & ~x87 & ~x106 & ~x113 & ~x170 & ~x179 & ~x181 & ~x182 & ~x196 & ~x208 & ~x224 & ~x250 & ~x251 & ~x303 & ~x308 & ~x362 & ~x390 & ~x420 & ~x500 & ~x531 & ~x587 & ~x644 & ~x724 & ~x727 & ~x782;
assign c3234 = ~x323 & ~x377 & ~x378 & ~x380 & ~x408 & ~x429 & ~x477 & ~x613 & ~x637 & ~x640 & ~x643 & ~x672 & ~x691 & ~x745;
assign c3236 =  x469 &  x497 & ~x462 & ~x491 & ~x535 & ~x567 & ~x589 & ~x591;
assign c3238 = ~x351 & ~x406 & ~x431 & ~x432 & ~x450 & ~x458 & ~x514 & ~x530 & ~x531 & ~x533 & ~x534 & ~x557 & ~x560 & ~x566 & ~x619 & ~x669 & ~x689 & ~x690 & ~x718 & ~x744 & ~x745 & ~x772 & ~x773 & ~x775 & ~x780;
assign c3240 =  x562 &  x647 &  x677 & ~x38 & ~x66 & ~x113 & ~x599 & ~x672;
assign c3242 =  x350 & ~x47 & ~x56 & ~x140 & ~x156 & ~x516 & ~x520 & ~x596 & ~x625 & ~x650 & ~x703;
assign c3244 = ~x4 & ~x5 & ~x20 & ~x27 & ~x58 & ~x84 & ~x85 & ~x106 & ~x111 & ~x112 & ~x168 & ~x251 & ~x307 & ~x357 & ~x385 & ~x413 & ~x433 & ~x434 & ~x435 & ~x460 & ~x492 & ~x518 & ~x520 & ~x548 & ~x595 & ~x624 & ~x651 & ~x700 & ~x727 & ~x728 & ~x755 & ~x756;
assign c3246 = ~x8 & ~x37 & ~x109 & ~x147 & ~x162 & ~x172 & ~x203 & ~x275 & ~x422 & ~x603 & ~x627 & ~x651 & ~x679 & ~x705 & ~x734;
assign c3248 = ~x1 & ~x59 & ~x139 & ~x326 & ~x350 & ~x380 & ~x410 & ~x431 & ~x432 & ~x437 & ~x505 & ~x507 & ~x564 & ~x592 & ~x596 & ~x616 & ~x643 & ~x693 & ~x720 & ~x721 & ~x748 & ~x752 & ~x778;
assign c3250 =  x528 & ~x18 & ~x168 & ~x357 & ~x414 & ~x459 & ~x469 & ~x524 & ~x615;
assign c3252 = ~x355 & ~x381 & ~x434 & ~x436 & ~x456 & ~x461 & ~x483 & ~x529 & ~x748 & ~x783;
assign c3254 =  x474 & ~x97 & ~x331 & ~x382;
assign c3256 =  x453 &  x481 &  x509 & ~x1 & ~x26 & ~x29 & ~x31 & ~x52 & ~x56 & ~x58 & ~x60 & ~x83 & ~x87 & ~x89 & ~x115 & ~x138 & ~x167 & ~x168 & ~x171 & ~x193 & ~x226 & ~x248 & ~x276 & ~x279 & ~x281 & ~x332 & ~x335 & ~x394 & ~x421 & ~x444 & ~x445 & ~x446 & ~x501 & ~x505 & ~x507 & ~x556 & ~x591 & ~x612 & ~x614 & ~x616 & ~x617 & ~x619 & ~x640 & ~x648 & ~x672 & ~x674 & ~x675 & ~x758 & ~x759;
assign c3258 =  x278 &  x362 & ~x301 & ~x358 & ~x382 & ~x385 & ~x412 & ~x438 & ~x459 & ~x463 & ~x466;
assign c3260 =  x318 &  x474 & ~x141 & ~x199 & ~x496 & ~x570 & ~x625 & ~x628 & ~x651;
assign c3262 =  x562 &  x590 & ~x6 & ~x84 & ~x113 & ~x280 & ~x287 & ~x342 & ~x370 & ~x425 & ~x453 & ~x458 & ~x515 & ~x542 & ~x544 & ~x570 & ~x700;
assign c3264 = ~x5 & ~x33 & ~x167 & ~x327 & ~x363 & ~x365 & ~x410 & ~x420 & ~x435 & ~x489 & ~x504 & ~x529 & ~x557 & ~x560 & ~x635 & ~x725 & ~x753;
assign c3266 =  x306 &  x334 & ~x56 & ~x115 & ~x359 & ~x380 & ~x385 & ~x386 & ~x411 & ~x413 & ~x440 & ~x467;
assign c3268 = ~x2 & ~x22 & ~x84 & ~x139 & ~x243 & ~x297 & ~x327 & ~x420 & ~x423 & ~x437 & ~x451 & ~x452 & ~x506 & ~x560 & ~x563 & ~x619 & ~x704 & ~x728;
assign c3270 = ~x50 & ~x52 & ~x141 & ~x145 & ~x171 & ~x253 & ~x433 & ~x471 & ~x604 & ~x619 & ~x639 & ~x684 & ~x705 & ~x710 & ~x739 & ~x756;
assign c3272 =  x379 & ~x1 & ~x30 & ~x77 & ~x78 & ~x79 & ~x110 & ~x111 & ~x114 & ~x138 & ~x141 & ~x142 & ~x164 & ~x165 & ~x167 & ~x198 & ~x220 & ~x248 & ~x253 & ~x276 & ~x277 & ~x281 & ~x282 & ~x306 & ~x334 & ~x362 & ~x447 & ~x572 & ~x599 & ~x628 & ~x642 & ~x656 & ~x670 & ~x684 & ~x685 & ~x698 & ~x699 & ~x711 & ~x713 & ~x714 & ~x728 & ~x738 & ~x739 & ~x754 & ~x756 & ~x781;
assign c3274 =  x160 &  x328 & ~x7 & ~x22 & ~x24 & ~x52 & ~x57 & ~x79 & ~x108 & ~x114 & ~x139 & ~x197 & ~x222 & ~x224 & ~x249 & ~x252 & ~x253 & ~x279 & ~x305 & ~x311 & ~x363 & ~x365 & ~x418 & ~x421 & ~x473 & ~x499 & ~x505 & ~x530 & ~x531 & ~x555 & ~x558 & ~x585 & ~x616 & ~x645 & ~x670 & ~x673 & ~x699 & ~x727 & ~x729;
assign c3276 =  x245 & ~x0 & ~x22 & ~x39 & ~x52 & ~x79 & ~x85 & ~x112 & ~x113 & ~x181 & ~x195 & ~x224 & ~x281 & ~x304 & ~x388 & ~x405 & ~x444 & ~x503 & ~x531 & ~x613 & ~x641 & ~x700 & ~x727;
assign c3278 =  x425 &  x453 & ~x0 & ~x1 & ~x3 & ~x25 & ~x30 & ~x55 & ~x57 & ~x58 & ~x60 & ~x81 & ~x112 & ~x113 & ~x116 & ~x143 & ~x165 & ~x166 & ~x168 & ~x172 & ~x194 & ~x197 & ~x222 & ~x249 & ~x252 & ~x253 & ~x254 & ~x277 & ~x280 & ~x307 & ~x310 & ~x334 & ~x335 & ~x336 & ~x361 & ~x363 & ~x393 & ~x417 & ~x445 & ~x446 & ~x447 & ~x448 & ~x449 & ~x450 & ~x473 & ~x474 & ~x476 & ~x501 & ~x504 & ~x505 & ~x529 & ~x530 & ~x557 & ~x558 & ~x561 & ~x562 & ~x574 & ~x585 & ~x586 & ~x587 & ~x589 & ~x590 & ~x613 & ~x614 & ~x616 & ~x617 & ~x631 & ~x642 & ~x644 & ~x669 & ~x670 & ~x685 & ~x712 & ~x725 & ~x726 & ~x727 & ~x728 & ~x730 & ~x731 & ~x752 & ~x753;
assign c3280 =  x388 &  x416 &  x556 & ~x58 & ~x59 & ~x111 & ~x114 & ~x170 & ~x196 & ~x504 & ~x522 & ~x548 & ~x727;
assign c3282 =  x418 & ~x46 & ~x329 & ~x411 & ~x560 & ~x566 & ~x721;
assign c3284 =  x721 & ~x521 & ~x522 & ~x544 & ~x574 & ~x602 & ~x683 & ~x767;
assign c3286 =  x552 &  x553 &  x580 & ~x3 & ~x4 & ~x26 & ~x27 & ~x53 & ~x54 & ~x57 & ~x112 & ~x113 & ~x195 & ~x487 & ~x514 & ~x542 & ~x543 & ~x558 & ~x571 & ~x597 & ~x723 & ~x724 & ~x725 & ~x727 & ~x728 & ~x751 & ~x754 & ~x773 & ~x774;
assign c3288 =  x296 & ~x327 & ~x411 & ~x435 & ~x461 & ~x492 & ~x494;
assign c3290 = ~x140 & ~x290 & ~x381 & ~x382 & ~x401 & ~x425 & ~x448 & ~x539 & ~x564;
assign c3292 = ~x98 & ~x140 & ~x413 & ~x414 & ~x443 & ~x469 & ~x489 & ~x490 & ~x519 & ~x520 & ~x521 & ~x547 & ~x553 & ~x572 & ~x573 & ~x576 & ~x604 & ~x627 & ~x682 & ~x758;
assign c3294 =  x323 & ~x30 & ~x84 & ~x160 & ~x194 & ~x436 & ~x546 & ~x574 & ~x628 & ~x656 & ~x707 & ~x709 & ~x711;
assign c3296 =  x425 &  x537 & ~x0 & ~x26 & ~x109 & ~x110 & ~x112 & ~x139 & ~x141 & ~x144 & ~x194 & ~x199 & ~x200 & ~x221 & ~x222 & ~x223 & ~x227 & ~x277 & ~x281 & ~x304 & ~x305 & ~x333 & ~x334 & ~x335 & ~x339 & ~x360 & ~x366 & ~x392 & ~x394 & ~x416 & ~x417 & ~x418 & ~x421 & ~x444 & ~x445 & ~x449 & ~x450 & ~x473 & ~x474 & ~x476 & ~x477 & ~x478 & ~x500 & ~x505 & ~x506 & ~x529 & ~x530 & ~x531 & ~x534 & ~x556 & ~x557 & ~x558 & ~x560 & ~x561 & ~x562 & ~x586 & ~x588 & ~x589 & ~x617 & ~x618 & ~x641 & ~x642 & ~x643 & ~x644 & ~x647 & ~x669 & ~x671 & ~x672 & ~x675 & ~x697 & ~x702 & ~x703 & ~x725 & ~x726 & ~x731 & ~x752;
assign c3298 =  x319 &  x390 & ~x170 & ~x494;
assign c3300 = ~x272 & ~x297 & ~x319 & ~x323 & ~x352 & ~x374 & ~x378 & ~x379 & ~x449 & ~x507 & ~x508 & ~x539 & ~x614 & ~x724;
assign c3302 =  x412 & ~x22 & ~x36 & ~x37 & ~x64 & ~x65 & ~x84 & ~x93 & ~x94 & ~x110 & ~x111 & ~x122 & ~x138 & ~x167 & ~x195 & ~x224 & ~x249 & ~x251 & ~x276 & ~x304 & ~x306 & ~x308 & ~x391 & ~x476 & ~x543 & ~x571 & ~x627 & ~x628 & ~x656 & ~x670 & ~x671 & ~x685 & ~x711;
assign c3304 = ~x28 & ~x52 & ~x85 & ~x383 & ~x438 & ~x439 & ~x458 & ~x512 & ~x561 & ~x562 & ~x565 & ~x588 & ~x589 & ~x592 & ~x595 & ~x614 & ~x615 & ~x667 & ~x672 & ~x693 & ~x718 & ~x719 & ~x727 & ~x729 & ~x748 & ~x769 & ~x777 & ~x781;
assign c3306 =  x128 & ~x23 & ~x28 & ~x57 & ~x58 & ~x109 & ~x110 & ~x112 & ~x138 & ~x168 & ~x264 & ~x291 & ~x374 & ~x402 & ~x430 & ~x447 & ~x458 & ~x475 & ~x504 & ~x529 & ~x542 & ~x560 & ~x616 & ~x701 & ~x757;
assign c3308 =  x352 &  x356 & ~x81 & ~x86 & ~x164 & ~x165 & ~x194 & ~x195 & ~x265 & ~x278 & ~x545 & ~x573 & ~x643 & ~x657;
assign c3310 =  x159 & ~x3 & ~x12 & ~x21 & ~x22 & ~x84 & ~x293 & ~x308 & ~x309 & ~x321 & ~x349 & ~x371 & ~x391 & ~x399 & ~x432 & ~x475 & ~x476 & ~x515 & ~x543 & ~x559 & ~x571 & ~x642 & ~x643;
assign c3312 =  x370 &  x552 & ~x24 & ~x53 & ~x82 & ~x107 & ~x530 & ~x585 & ~x586 & ~x611 & ~x614 & ~x642 & ~x674 & ~x695 & ~x753 & ~x758 & ~x779;
assign c3314 =  x239 & ~x14 & ~x24 & ~x353 & ~x381 & ~x559 & ~x678 & ~x689 & ~x698;
assign c3316 = ~x5 & ~x7 & ~x30 & ~x38 & ~x50 & ~x65 & ~x66 & ~x94 & ~x135 & ~x138 & ~x141 & ~x149 & ~x161 & ~x222 & ~x223 & ~x282 & ~x283 & ~x338 & ~x416 & ~x626 & ~x642 & ~x681 & ~x698 & ~x736 & ~x737;
assign c3318 =  x185 &  x186 & ~x0 & ~x2 & ~x30 & ~x39 & ~x52 & ~x55 & ~x56 & ~x57 & ~x68 & ~x69 & ~x83 & ~x166 & ~x167 & ~x198 & ~x224 & ~x251 & ~x376 & ~x503 & ~x531 & ~x558 & ~x559 & ~x585 & ~x586 & ~x587 & ~x588 & ~x613 & ~x615 & ~x641 & ~x671 & ~x672 & ~x673 & ~x728 & ~x730 & ~x738 & ~x739 & ~x754 & ~x757 & ~x782;
assign c3320 = ~x0 & ~x2 & ~x23 & ~x24 & ~x25 & ~x30 & ~x31 & ~x106 & ~x111 & ~x141 & ~x143 & ~x144 & ~x164 & ~x167 & ~x192 & ~x193 & ~x195 & ~x196 & ~x207 & ~x219 & ~x223 & ~x225 & ~x226 & ~x254 & ~x276 & ~x304 & ~x308 & ~x334 & ~x361 & ~x362 & ~x388 & ~x392 & ~x394 & ~x414 & ~x420 & ~x432 & ~x442 & ~x444 & ~x448 & ~x472 & ~x473 & ~x477 & ~x479 & ~x500 & ~x501 & ~x531 & ~x532 & ~x557 & ~x559 & ~x562 & ~x572 & ~x591 & ~x601 & ~x613 & ~x617 & ~x618 & ~x619 & ~x642 & ~x644 & ~x646 & ~x672 & ~x700 & ~x701 & ~x722 & ~x725 & ~x726 & ~x731 & ~x732 & ~x750 & ~x754 & ~x758 & ~x779;
assign c3322 = ~x0 & ~x4 & ~x9 & ~x65 & ~x86 & ~x94 & ~x107 & ~x109 & ~x165 & ~x198 & ~x304 & ~x307 & ~x486 & ~x500 & ~x533 & ~x548 & ~x571 & ~x615 & ~x724 & ~x752 & ~x756;
assign c3324 =  x387 &  x443 & ~x54 & ~x82 & ~x300 & ~x460 & ~x465 & ~x476 & ~x502 & ~x531 & ~x533 & ~x560 & ~x588 & ~x701;
assign c3326 =  x278 & ~x274 & ~x319 & ~x458 & ~x481 & ~x515;
assign c3328 =  x352 &  x383 & ~x37 & ~x49 & ~x54 & ~x66 & ~x93 & ~x167 & ~x198 & ~x221 & ~x277;
assign c3330 =  x554 &  x582 & ~x0 & ~x29 & ~x85 & ~x87 & ~x111 & ~x140 & ~x171 & ~x197 & ~x225 & ~x251 & ~x252 & ~x467 & ~x491 & ~x493 & ~x505 & ~x522 & ~x549 & ~x558 & ~x559 & ~x562 & ~x586 & ~x614 & ~x641 & ~x670 & ~x698 & ~x725 & ~x726;
assign c3332 =  x479 &  x507 & ~x169 & ~x224 & ~x468 & ~x497 & ~x552 & ~x580;
assign c3334 =  x696 & ~x33 & ~x142 & ~x169 & ~x280 & ~x496 & ~x525 & ~x552 & ~x581;
assign c3336 =  x413 & ~x24 & ~x56 & ~x80 & ~x110 & ~x115 & ~x227 & ~x248 & ~x279 & ~x281 & ~x362 & ~x390 & ~x391 & ~x421 & ~x477 & ~x516 & ~x555 & ~x557 & ~x642 & ~x725;
assign c3338 =  x74 & ~x25 & ~x28 & ~x29 & ~x53 & ~x55 & ~x58 & ~x59 & ~x82 & ~x289 & ~x296 & ~x297 & ~x365 & ~x377 & ~x394 & ~x420 & ~x422 & ~x447 & ~x448 & ~x504 & ~x505 & ~x533 & ~x561 & ~x589 & ~x672 & ~x702;
assign c3340 = ~x33 & ~x110 & ~x116 & ~x200 & ~x223 & ~x255 & ~x278 & ~x450 & ~x461 & ~x473 & ~x505 & ~x528 & ~x557 & ~x589 & ~x601 & ~x617 & ~x644 & ~x646 & ~x670 & ~x683 & ~x705 & ~x709 & ~x755;
assign c3342 = ~x34 & ~x86 & ~x167 & ~x325 & ~x379 & ~x506 & ~x509 & ~x535 & ~x542 & ~x567 & ~x690;
assign c3344 = ~x22 & ~x30 & ~x107 & ~x114 & ~x135 & ~x164 & ~x173 & ~x201 & ~x213 & ~x221 & ~x226 & ~x251 & ~x309 & ~x311 & ~x491 & ~x519 & ~x595 & ~x648 & ~x649 & ~x650 & ~x654 & ~x681 & ~x706 & ~x709;
assign c3346 =  x340 &  x396 &  x479 &  x507 & ~x0 & ~x1 & ~x2 & ~x3 & ~x29 & ~x56 & ~x57 & ~x83 & ~x87 & ~x111 & ~x138 & ~x139 & ~x168 & ~x170 & ~x195 & ~x199 & ~x224 & ~x226 & ~x279 & ~x281 & ~x309 & ~x310 & ~x336 & ~x337 & ~x363 & ~x365 & ~x392 & ~x446 & ~x447 & ~x448 & ~x474 & ~x477 & ~x502 & ~x505 & ~x530 & ~x533 & ~x561 & ~x588 & ~x616 & ~x642 & ~x644 & ~x645 & ~x670 & ~x671 & ~x672 & ~x673 & ~x698 & ~x701 & ~x727 & ~x728 & ~x755 & ~x757 & ~x782 & ~x783;
assign c3348 =  x398 &  x426 & ~x29 & ~x80 & ~x277 & ~x312 & ~x332 & ~x396 & ~x506 & ~x545 & ~x615 & ~x642 & ~x704 & ~x780;
assign c3350 =  x47 & ~x2 & ~x293 & ~x321 & ~x323 & ~x419;
assign c3352 =  x125 &  x126 & ~x319 & ~x346 & ~x430 & ~x432 & ~x435 & ~x457 & ~x491 & ~x728;
assign c3354 =  x156 & ~x50 & ~x57 & ~x82 & ~x83 & ~x85 & ~x86 & ~x112 & ~x124 & ~x246 & ~x293 & ~x532 & ~x585 & ~x639 & ~x640 & ~x641 & ~x644 & ~x698 & ~x711 & ~x728 & ~x756 & ~x766 & ~x783;
assign c3356 =  x524 & ~x8 & ~x12 & ~x50 & ~x67 & ~x97 & ~x98 & ~x432 & ~x478 & ~x533 & ~x643 & ~x673 & ~x724 & ~x759;
assign c3358 =  x292 & ~x34 & ~x72 & ~x117 & ~x410 & ~x488 & ~x573 & ~x616 & ~x642 & ~x647 & ~x703 & ~x704 & ~x760;
assign c3360 =  x162 &  x358 & ~x25 & ~x138 & ~x393 & ~x449 & ~x477 & ~x529 & ~x585 & ~x586 & ~x588 & ~x614 & ~x615 & ~x700 & ~x758;
assign c3362 = ~x1 & ~x3 & ~x26 & ~x60 & ~x82 & ~x87 & ~x114 & ~x117 & ~x173 & ~x201 & ~x226 & ~x227 & ~x229 & ~x253 & ~x254 & ~x256 & ~x283 & ~x384 & ~x410 & ~x440 & ~x462 & ~x464 & ~x465 & ~x467 & ~x491 & ~x493 & ~x518 & ~x520 & ~x701 & ~x705 & ~x712 & ~x731 & ~x773;
assign c3364 =  x241 &  x451 & ~x26 & ~x140 & ~x357 & ~x410;
assign c3366 =  x380 & ~x36 & ~x40 & ~x122 & ~x320 & ~x363 & ~x445 & ~x543 & ~x556 & ~x655 & ~x698 & ~x757;
assign c3368 = ~x6 & ~x83 & ~x326 & ~x354 & ~x409 & ~x435 & ~x457 & ~x464 & ~x484 & ~x490 & ~x512 & ~x531 & ~x560 & ~x562 & ~x566 & ~x568 & ~x592 & ~x616 & ~x622 & ~x643 & ~x652 & ~x671 & ~x677 & ~x694 & ~x725;
assign c3370 =  x562 &  x697 & ~x554;
assign c3372 = ~x291 & ~x292 & ~x325 & ~x347 & ~x375 & ~x376 & ~x380 & ~x398 & ~x408 & ~x426 & ~x436 & ~x448 & ~x503 & ~x504 & ~x510 & ~x667 & ~x672 & ~x693 & ~x783;
assign c3374 = ~x111 & ~x144 & ~x172 & ~x273 & ~x351 & ~x379 & ~x409 & ~x411 & ~x468 & ~x562 & ~x589 & ~x616;
assign c3376 =  x378 & ~x84 & ~x138 & ~x164 & ~x487 & ~x491 & ~x547 & ~x575 & ~x627 & ~x682 & ~x737;
assign c3378 = ~x35 & ~x98 & ~x200 & ~x227 & ~x465 & ~x474 & ~x547 & ~x561 & ~x644 & ~x648 & ~x651 & ~x672 & ~x732;
assign c3380 = ~x2 & ~x8 & ~x9 & ~x22 & ~x23 & ~x25 & ~x28 & ~x55 & ~x78 & ~x81 & ~x83 & ~x84 & ~x140 & ~x141 & ~x167 & ~x169 & ~x192 & ~x251 & ~x252 & ~x307 & ~x337 & ~x364 & ~x463 & ~x474 & ~x504 & ~x516 & ~x517 & ~x518 & ~x531 & ~x546 & ~x559 & ~x626 & ~x627 & ~x629 & ~x644 & ~x680 & ~x698 & ~x709 & ~x728 & ~x753 & ~x756 & ~x758 & ~x781;
assign c3382 = ~x6 & ~x51 & ~x55 & ~x56 & ~x82 & ~x87 & ~x88 & ~x110 & ~x113 & ~x115 & ~x117 & ~x141 & ~x164 & ~x168 & ~x171 & ~x172 & ~x194 & ~x200 & ~x224 & ~x278 & ~x280 & ~x307 & ~x308 & ~x312 & ~x333 & ~x335 & ~x338 & ~x339 & ~x361 & ~x364 & ~x365 & ~x395 & ~x417 & ~x422 & ~x450 & ~x472 & ~x476 & ~x477 & ~x489 & ~x501 & ~x503 & ~x506 & ~x532 & ~x533 & ~x545 & ~x557 & ~x573 & ~x586 & ~x590 & ~x642 & ~x671 & ~x696 & ~x701 & ~x739 & ~x751 & ~x755 & ~x779 & ~x782;
assign c3384 =  x211 & ~x7 & ~x201 & ~x302 & ~x468 & ~x489 & ~x547 & ~x654 & ~x739;
assign c3386 =  x508 & ~x0 & ~x32 & ~x58 & ~x59 & ~x86 & ~x91 & ~x172 & ~x198 & ~x199 & ~x200 & ~x201 & ~x225 & ~x227 & ~x252 & ~x254 & ~x255 & ~x256 & ~x282 & ~x283 & ~x311 & ~x364 & ~x542 & ~x570 & ~x623 & ~x652 & ~x655 & ~x679 & ~x682 & ~x709 & ~x736 & ~x755;
assign c3388 =  x268 & ~x27 & ~x31 & ~x61 & ~x87 & ~x170 & ~x198 & ~x225 & ~x327 & ~x355 & ~x381 & ~x382 & ~x406 & ~x411 & ~x461 & ~x729;
assign c3390 = ~x1 & ~x43 & ~x70 & ~x86 & ~x112 & ~x115 & ~x152 & ~x381 & ~x435 & ~x442 & ~x463 & ~x465 & ~x470 & ~x490 & ~x520 & ~x523 & ~x525 & ~x547 & ~x550;
assign c3392 =  x205 & ~x29 & ~x34 & ~x58 & ~x108 & ~x114 & ~x167 & ~x491 & ~x519 & ~x575 & ~x576 & ~x600 & ~x678;
assign c3394 =  x359 &  x638 & ~x293 & ~x307 & ~x572 & ~x575 & ~x599 & ~x604 & ~x628 & ~x632 & ~x783;
assign c3396 =  x220 & ~x44 & ~x168 & ~x371 & ~x404 & ~x405 & ~x475 & ~x476 & ~x588 & ~x701;
assign c3398 =  x425 & ~x9 & ~x39 & ~x94 & ~x142 & ~x311 & ~x388 & ~x389 & ~x392 & ~x432 & ~x445 & ~x460 & ~x543 & ~x558 & ~x560 & ~x616 & ~x672 & ~x701;
assign c3400 = ~x0 & ~x2 & ~x24 & ~x25 & ~x26 & ~x27 & ~x28 & ~x29 & ~x30 & ~x42 & ~x50 & ~x51 & ~x52 & ~x53 & ~x54 & ~x57 & ~x58 & ~x59 & ~x60 & ~x78 & ~x81 & ~x82 & ~x84 & ~x87 & ~x113 & ~x115 & ~x139 & ~x140 & ~x141 & ~x142 & ~x143 & ~x144 & ~x165 & ~x166 & ~x170 & ~x171 & ~x193 & ~x194 & ~x196 & ~x198 & ~x199 & ~x221 & ~x222 & ~x224 & ~x225 & ~x247 & ~x248 & ~x249 & ~x251 & ~x253 & ~x254 & ~x281 & ~x282 & ~x303 & ~x304 & ~x305 & ~x306 & ~x307 & ~x310 & ~x311 & ~x332 & ~x333 & ~x335 & ~x338 & ~x339 & ~x361 & ~x365 & ~x366 & ~x390 & ~x391 & ~x393 & ~x394 & ~x416 & ~x417 & ~x419 & ~x446 & ~x447 & ~x448 & ~x449 & ~x474 & ~x475 & ~x476 & ~x478 & ~x502 & ~x503 & ~x505 & ~x527 & ~x528 & ~x529 & ~x530 & ~x532 & ~x555 & ~x556 & ~x557 & ~x559 & ~x560 & ~x583 & ~x584 & ~x585 & ~x586 & ~x587 & ~x588 & ~x601 & ~x612 & ~x616 & ~x617 & ~x629 & ~x641 & ~x642 & ~x644 & ~x645 & ~x668 & ~x669 & ~x670 & ~x671 & ~x696 & ~x697 & ~x702 & ~x703 & ~x704 & ~x723 & ~x724 & ~x725 & ~x729 & ~x731 & ~x751 & ~x754 & ~x758 & ~x760 & ~x761 & ~x779 & ~x780 & ~x782;
assign c3402 =  x355 & ~x12 & ~x168 & ~x224 & ~x236 & ~x291 & ~x343 & ~x389 & ~x416 & ~x418 & ~x446 & ~x559 & ~x644 & ~x727 & ~x756 & ~x783;
assign c3404 =  x669 & ~x301 & ~x553 & ~x554 & ~x682;
assign c3406 =  x578 & ~x6 & ~x433 & ~x434 & ~x490 & ~x491 & ~x548 & ~x567 & ~x569 & ~x587 & ~x641 & ~x748;
assign c3408 =  x472 & ~x324 & ~x380 & ~x383 & ~x429 & ~x561 & ~x565 & ~x566;
assign c3410 =  x555 & ~x45 & ~x329 & ~x357 & ~x412 & ~x467 & ~x538;
assign c3412 =  x585 & ~x29 & ~x58 & ~x84 & ~x141 & ~x440 & ~x467 & ~x469 & ~x470 & ~x498 & ~x520 & ~x525 & ~x526 & ~x548 & ~x552 & ~x573 & ~x580 & ~x629 & ~x654;
assign c3414 =  x229 &  x312 & ~x1 & ~x84 & ~x112 & ~x113 & ~x142 & ~x169 & ~x195 & ~x223 & ~x225 & ~x251 & ~x307 & ~x370 & ~x398 & ~x420 & ~x426 & ~x431 & ~x487 & ~x531 & ~x546 & ~x559 & ~x560 & ~x574 & ~x615 & ~x626 & ~x672 & ~x783;
assign c3416 =  x526 & ~x28 & ~x29 & ~x33 & ~x109 & ~x112 & ~x355 & ~x406 & ~x411 & ~x437 & ~x495 & ~x506 & ~x562 & ~x589 & ~x674 & ~x697;
assign c3418 = ~x24 & ~x32 & ~x55 & ~x56 & ~x83 & ~x110 & ~x378 & ~x391 & ~x394 & ~x407 & ~x434 & ~x450 & ~x503 & ~x507 & ~x516 & ~x518 & ~x536 & ~x617 & ~x639 & ~x705 & ~x716 & ~x717 & ~x728 & ~x729 & ~x743 & ~x754;
assign c3420 =  x526 & ~x26 & ~x115 & ~x116 & ~x356 & ~x435 & ~x437 & ~x440 & ~x613 & ~x645 & ~x646 & ~x669 & ~x670 & ~x699;
assign c3422 = ~x14 & ~x112 & ~x273 & ~x399 & ~x425 & ~x426 & ~x439 & ~x466 & ~x491 & ~x672 & ~x700 & ~x711 & ~x729 & ~x759;
assign c3424 =  x424 & ~x113 & ~x144 & ~x197 & ~x223 & ~x227 & ~x254 & ~x256 & ~x283 & ~x310 & ~x311 & ~x412 & ~x439 & ~x465 & ~x468 & ~x489 & ~x494 & ~x496 & ~x524 & ~x548;
assign c3426 =  x648 &  x676 & ~x9 & ~x22 & ~x25 & ~x55 & ~x81 & ~x94 & ~x113 & ~x167 & ~x196 & ~x224 & ~x252 & ~x292 & ~x348 & ~x375 & ~x447 & ~x514 & ~x515 & ~x542 & ~x543 & ~x571 & ~x572 & ~x615 & ~x626 & ~x644 & ~x671 & ~x700 & ~x728 & ~x729;
assign c3428 =  x422 & ~x0 & ~x6 & ~x141 & ~x142 & ~x168 & ~x169 & ~x170 & ~x198 & ~x226 & ~x253 & ~x414 & ~x442 & ~x486 & ~x541 & ~x545 & ~x672;
assign c3430 =  x43 & ~x111 & ~x138 & ~x260 & ~x292 & ~x472 & ~x516;
assign c3432 =  x74 &  x274 & ~x292 & ~x320 & ~x321 & ~x348 & ~x363 & ~x431 & ~x444 & ~x500 & ~x501 & ~x529 & ~x530 & ~x616 & ~x672;
assign c3434 = ~x0 & ~x26 & ~x57 & ~x61 & ~x83 & ~x85 & ~x86 & ~x112 & ~x115 & ~x244 & ~x246 & ~x270 & ~x271 & ~x273 & ~x275 & ~x279 & ~x301 & ~x303 & ~x523 & ~x524 & ~x601 & ~x628 & ~x651 & ~x652 & ~x679 & ~x680 & ~x699 & ~x705 & ~x708 & ~x709 & ~x761 & ~x762 & ~x765 & ~x783;
assign c3436 =  x320 &  x423 & ~x100 & ~x116 & ~x438 & ~x439 & ~x467 & ~x516 & ~x616;
assign c3438 =  x324 &  x637 & ~x1 & ~x21 & ~x28 & ~x29 & ~x55 & ~x94 & ~x113 & ~x138 & ~x166 & ~x194 & ~x222 & ~x223 & ~x573 & ~x616 & ~x700 & ~x712 & ~x728 & ~x755;
assign c3440 =  x326 &  x506 &  x534 & ~x85 & ~x252 & ~x516 & ~x570 & ~x598 & ~x672;
assign c3442 =  x178 & ~x3 & ~x28 & ~x31 & ~x34 & ~x402 & ~x484 & ~x485 & ~x486 & ~x542 & ~x719 & ~x720;
assign c3444 = ~x5 & ~x62 & ~x107 & ~x135 & ~x464 & ~x465 & ~x504 & ~x509 & ~x519 & ~x535 & ~x537 & ~x545 & ~x546 & ~x547 & ~x562 & ~x572 & ~x601 & ~x621 & ~x622 & ~x645 & ~x655 & ~x678 & ~x751;
assign c3446 =  x356 &  x411 & ~x27 & ~x80 & ~x81 & ~x84 & ~x85 & ~x110 & ~x166 & ~x167 & ~x252 & ~x292 & ~x370 & ~x445 & ~x446 & ~x475 & ~x499 & ~x502 & ~x527 & ~x529 & ~x530 & ~x643 & ~x755 & ~x783;
assign c3448 =  x352 &  x383 &  x663 & ~x66 & ~x306 & ~x307 & ~x308 & ~x392 & ~x504 & ~x644 & ~x671 & ~x672 & ~x683;
assign c3450 =  x293 &  x553 & ~x0 & ~x559 & ~x652 & ~x671 & ~x701;
assign c3452 = ~x89 & ~x377 & ~x408 & ~x409 & ~x420 & ~x434 & ~x478 & ~x492 & ~x510 & ~x537 & ~x621 & ~x623 & ~x729 & ~x745;
assign c3454 =  x534 &  x562 &  x613 & ~x141 & ~x168 & ~x169 & ~x197 & ~x253 & ~x441 & ~x470 & ~x626;
assign c3456 = ~x5 & ~x117 & ~x129 & ~x142 & ~x144 & ~x196 & ~x199 & ~x200 & ~x201 & ~x226 & ~x245 & ~x467 & ~x493 & ~x519 & ~x521 & ~x654 & ~x655 & ~x681 & ~x699 & ~x708 & ~x709 & ~x728;
assign c3458 = ~x97 & ~x424 & ~x453 & ~x480 & ~x491 & ~x510 & ~x520 & ~x674 & ~x675 & ~x768;
assign c3460 = ~x1 & ~x29 & ~x36 & ~x57 & ~x64 & ~x92 & ~x100 & ~x156 & ~x162 & ~x174 & ~x183 & ~x196 & ~x228 & ~x283 & ~x284 & ~x578 & ~x598 & ~x650 & ~x652 & ~x653 & ~x654 & ~x678 & ~x679 & ~x680 & ~x705 & ~x708;
assign c3462 =  x306 & ~x350 & ~x378 & ~x407 & ~x465;
assign c3464 =  x186 &  x650 & ~x2 & ~x8 & ~x95 & ~x320 & ~x348 & ~x376 & ~x615 & ~x684 & ~x701 & ~x728 & ~x757 & ~x758;
assign c3466 =  x241 &  x594 & ~x22 & ~x31 & ~x34 & ~x39 & ~x49 & ~x58 & ~x67 & ~x81 & ~x82 & ~x85 & ~x110 & ~x115 & ~x138 & ~x170 & ~x198 & ~x224 & ~x253 & ~x280 & ~x281 & ~x336 & ~x447 & ~x474 & ~x475 & ~x531 & ~x560 & ~x587 & ~x644 & ~x655 & ~x672 & ~x701 & ~x730 & ~x738 & ~x755 & ~x783;
assign c3468 =  x102 &  x622 & ~x37 & ~x38 & ~x168 & ~x471 & ~x502 & ~x557 & ~x615 & ~x728 & ~x759;
assign c3470 = ~x0 & ~x2 & ~x9 & ~x25 & ~x26 & ~x27 & ~x29 & ~x30 & ~x36 & ~x38 & ~x39 & ~x55 & ~x57 & ~x81 & ~x82 & ~x84 & ~x85 & ~x87 & ~x94 & ~x109 & ~x114 & ~x137 & ~x138 & ~x139 & ~x140 & ~x142 & ~x143 & ~x150 & ~x166 & ~x168 & ~x194 & ~x196 & ~x197 & ~x223 & ~x224 & ~x249 & ~x250 & ~x252 & ~x253 & ~x279 & ~x280 & ~x282 & ~x305 & ~x306 & ~x307 & ~x309 & ~x334 & ~x362 & ~x363 & ~x390 & ~x391 & ~x417 & ~x418 & ~x419 & ~x420 & ~x474 & ~x475 & ~x477 & ~x501 & ~x505 & ~x529 & ~x532 & ~x533 & ~x558 & ~x561 & ~x571 & ~x587 & ~x588 & ~x614 & ~x615 & ~x616 & ~x617 & ~x627 & ~x643 & ~x655 & ~x670 & ~x672 & ~x673 & ~x699 & ~x726 & ~x727 & ~x728 & ~x729 & ~x782 & ~x783;
assign c3472 =  x611 & ~x88 & ~x493 & ~x496 & ~x544 & ~x561 & ~x644 & ~x645 & ~x674;
assign c3474 =  x410 &  x411 &  x438 &  x465 & ~x23 & ~x24 & ~x108 & ~x109 & ~x110 & ~x137 & ~x140 & ~x168 & ~x169 & ~x197 & ~x222 & ~x251 & ~x280 & ~x281 & ~x306 & ~x333 & ~x348 & ~x530 & ~x543 & ~x557 & ~x727;
assign c3476 =  x387 &  x722 & ~x56 & ~x81 & ~x142 & ~x168 & ~x279 & ~x364 & ~x476;
assign c3478 = ~x8 & ~x27 & ~x232 & ~x252 & ~x286 & ~x291 & ~x320 & ~x342 & ~x348 & ~x369 & ~x370 & ~x374 & ~x402 & ~x419 & ~x426 & ~x430 & ~x447 & ~x458 & ~x514 & ~x597;
assign c3480 =  x233 &  x288 & ~x57 & ~x119 & ~x488 & ~x596 & ~x773;
assign c3482 = ~x0 & ~x2 & ~x26 & ~x31 & ~x139 & ~x432 & ~x506 & ~x507 & ~x517 & ~x518 & ~x540 & ~x564 & ~x568 & ~x585 & ~x593 & ~x598 & ~x612 & ~x623 & ~x624 & ~x650 & ~x669 & ~x696 & ~x697 & ~x745 & ~x776;
assign c3484 = ~x25 & ~x118 & ~x134 & ~x145 & ~x146 & ~x168 & ~x169 & ~x174 & ~x202 & ~x229 & ~x281 & ~x284 & ~x295 & ~x310 & ~x335 & ~x339 & ~x653 & ~x678 & ~x680 & ~x706 & ~x709 & ~x736;
assign c3486 = ~x6 & ~x29 & ~x36 & ~x52 & ~x114 & ~x141 & ~x197 & ~x278 & ~x416 & ~x419 & ~x489 & ~x516 & ~x561 & ~x613 & ~x631 & ~x682 & ~x734 & ~x752 & ~x780;
assign c3488 =  x610 & ~x86 & ~x114 & ~x142 & ~x468 & ~x522 & ~x544 & ~x550 & ~x551 & ~x645 & ~x656 & ~x674 & ~x700 & ~x732;
assign c3490 =  x203 & ~x117 & ~x172 & ~x344 & ~x521 & ~x523;
assign c3492 =  x371 & ~x27 & ~x35 & ~x88 & ~x142 & ~x144 & ~x173 & ~x229 & ~x284 & ~x490 & ~x596 & ~x622 & ~x625 & ~x627 & ~x648 & ~x676 & ~x677 & ~x678 & ~x705 & ~x728 & ~x733 & ~x773 & ~x780;
assign c3494 =  x637 & ~x112 & ~x139 & ~x165 & ~x194 & ~x250 & ~x434 & ~x518 & ~x562 & ~x574 & ~x576 & ~x590 & ~x603 & ~x632 & ~x644 & ~x647 & ~x729 & ~x732 & ~x753 & ~x780;
assign c3496 =  x355 & ~x6 & ~x22 & ~x34 & ~x38 & ~x52 & ~x55 & ~x56 & ~x108 & ~x111 & ~x112 & ~x139 & ~x164 & ~x168 & ~x170 & ~x236 & ~x263 & ~x265 & ~x291 & ~x319 & ~x320 & ~x348 & ~x517 & ~x572;
assign c3498 =  x442 &  x722 & ~x280 & ~x327 & ~x362 & ~x754;
assign c31 = ~x19 & ~x23 & ~x28 & ~x39 & ~x42 & ~x44 & ~x111 & ~x138 & ~x207 & ~x234 & ~x293 & ~x392 & ~x487 & ~x572 & ~x718 & ~x726 & ~x736 & ~x750 & ~x752 & ~x757 & ~x760 & ~x774 & ~x782;
assign c33 = ~x23 & ~x30 & ~x82 & ~x112 & ~x219 & ~x245 & ~x246 & ~x247 & ~x272 & ~x273 & ~x277 & ~x305 & ~x307 & ~x328 & ~x329 & ~x330 & ~x332 & ~x333 & ~x335 & ~x360 & ~x443 & ~x461 & ~x470 & ~x672 & ~x690 & ~x757;
assign c35 =  x145 &  x342 & ~x97 & ~x123 & ~x124;
assign c37 =  x285;
assign c39 = ~x12 & ~x15 & ~x24 & ~x30 & ~x52 & ~x79 & ~x88 & ~x101 & ~x125 & ~x127 & ~x129 & ~x220 & ~x225 & ~x227 & ~x279 & ~x405 & ~x448 & ~x732 & ~x756 & ~x769;
assign c311 =  x323 &  x518 & ~x678;
assign c313 =  x507 & ~x22 & ~x294 & ~x295 & ~x322 & ~x379 & ~x518 & ~x545 & ~x771;
assign c315 = ~x8 & ~x12 & ~x45 & ~x78 & ~x79 & ~x80 & ~x105 & ~x130 & ~x137 & ~x225 & ~x252 & ~x483 & ~x529 & ~x531 & ~x558 & ~x591 & ~x616 & ~x730;
assign c317 = ~x24 & ~x40 & ~x41 & ~x97 & ~x124 & ~x211 & ~x266 & ~x268 & ~x323 & ~x353 & ~x403 & ~x571 & ~x599 & ~x669 & ~x670 & ~x779;
assign c319 =  x321 &  x430 & ~x451;
assign c321 = ~x428 & ~x451 & ~x456 & ~x469 & ~x470 & ~x471 & ~x478 & ~x500 & ~x506 & ~x510 & ~x529 & ~x537 & ~x558 & ~x559 & ~x597 & ~x733 & ~x766;
assign c323 =  x571 & ~x26 & ~x47 & ~x49 & ~x391 & ~x559;
assign c325 =  x538 & ~x17 & ~x52 & ~x112 & ~x212 & ~x239 & ~x379 & ~x777;
assign c327 = ~x18 & ~x71 & ~x80 & ~x96 & ~x109 & ~x138 & ~x139 & ~x207 & ~x208 & ~x234 & ~x263 & ~x336 & ~x380 & ~x462 & ~x600 & ~x627 & ~x656 & ~x747 & ~x778;
assign c329 =  x547 & ~x5 & ~x335 & ~x485 & ~x683;
assign c331 = ~x13 & ~x14 & ~x17 & ~x43 & ~x55 & ~x100 & ~x248 & ~x250 & ~x251 & ~x279 & ~x303 & ~x309 & ~x331 & ~x334 & ~x359 & ~x365 & ~x379 & ~x416 & ~x431;
assign c333 =  x553 &  x639 & ~x45;
assign c335 =  x486 & ~x130 & ~x157 & ~x589 & ~x613 & ~x641 & ~x697 & ~x747 & ~x750 & ~x752;
assign c337 = ~x14 & ~x19 & ~x39 & ~x49 & ~x51 & ~x57 & ~x68 & ~x73 & ~x179 & ~x235 & ~x320 & ~x707;
assign c339 = ~x9 & ~x51 & ~x65 & ~x69 & ~x96 & ~x139 & ~x294 & ~x336 & ~x349 & ~x374 & ~x448 & ~x626 & ~x650 & ~x651 & ~x652 & ~x669 & ~x680 & ~x721 & ~x736 & ~x740;
assign c341 =  x179 &  x716 & ~x368;
assign c343 =  x518 & ~x278 & ~x281 & ~x307 & ~x364 & ~x511 & ~x641 & ~x651 & ~x706 & ~x733 & ~x738 & ~x755 & ~x777;
assign c345 =  x92 & ~x11 & ~x136 & ~x162;
assign c347 =  x351 &  x573;
assign c349 = ~x1 & ~x43 & ~x55 & ~x76 & ~x126 & ~x145 & ~x195 & ~x280 & ~x420 & ~x576 & ~x579 & ~x611 & ~x640 & ~x690 & ~x691 & ~x698 & ~x721 & ~x732 & ~x749 & ~x754;
assign c351 =  x569 & ~x721;
assign c353 =  x372 &  x456 & ~x268 & ~x408 & ~x519;
assign c355 =  x545 & ~x76 & ~x77 & ~x494 & ~x586;
assign c357 =  x417 &  x444 & ~x1 & ~x20 & ~x50 & ~x79 & ~x164 & ~x193 & ~x235 & ~x262 & ~x667 & ~x722 & ~x723 & ~x762;
assign c359 =  x592 &  x620 & ~x17 & ~x44 & ~x125 & ~x360 & ~x443;
assign c361 = ~x16 & ~x24 & ~x54 & ~x111 & ~x360 & ~x387 & ~x390 & ~x391 & ~x417 & ~x418 & ~x420 & ~x444 & ~x445 & ~x448 & ~x474 & ~x475 & ~x516 & ~x652 & ~x708 & ~x719 & ~x720 & ~x736 & ~x737 & ~x738 & ~x746 & ~x749 & ~x777 & ~x780;
assign c363 =  x397 &  x399 &  x454 & ~x206 & ~x448 & ~x458 & ~x682;
assign c365 =  x480 & ~x21 & ~x76 & ~x124 & ~x126 & ~x392 & ~x600 & ~x683 & ~x751;
assign c367 =  x434 &  x515;
assign c369 = ~x53 & ~x125 & ~x211 & ~x240 & ~x241 & ~x325 & ~x349 & ~x382 & ~x520;
assign c371 =  x374 &  x401 &  x538 &  x566;
assign c373 = ~x24 & ~x125 & ~x182 & ~x242 & ~x266 & ~x296 & ~x309 & ~x364 & ~x379 & ~x380 & ~x407 & ~x409 & ~x490 & ~x546 & ~x573;
assign c375 =  x541 & ~x61 & ~x112 & ~x163 & ~x192 & ~x281 & ~x454 & ~x750 & ~x769 & ~x778;
assign c377 =  x203 &  x371 &  x372 & ~x14 & ~x15 & ~x28 & ~x40 & ~x41 & ~x55 & ~x59 & ~x280 & ~x364 & ~x366 & ~x392 & ~x672 & ~x700 & ~x710;
assign c379 =  x94 &  x622 & ~x240 & ~x389;
assign c381 =  x570 & ~x45 & ~x46 & ~x107 & ~x643;
assign c383 =  x599 & ~x48 & ~x103 & ~x108 & ~x132 & ~x419;
assign c385 =  x238 &  x435 & ~x633;
assign c387 = ~x3 & ~x6 & ~x30 & ~x91 & ~x228 & ~x229 & ~x247 & ~x276 & ~x279 & ~x283 & ~x286 & ~x315 & ~x316 & ~x344 & ~x367 & ~x422 & ~x423 & ~x444 & ~x476 & ~x500 & ~x502 & ~x507 & ~x614 & ~x616 & ~x643 & ~x671 & ~x727 & ~x759;
assign c389 =  x455 & ~x101 & ~x263 & ~x450 & ~x477 & ~x741;
assign c391 =  x516 & ~x147 & ~x587;
assign c393 = ~x3 & ~x23 & ~x42 & ~x44 & ~x110 & ~x222 & ~x251 & ~x302 & ~x331 & ~x335 & ~x391 & ~x415 & ~x443 & ~x444 & ~x445 & ~x446 & ~x448 & ~x474 & ~x498 & ~x501 & ~x530 & ~x727 & ~x747 & ~x764;
assign c395 =  x375 &  x512 & ~x352;
assign c397 =  x541 &  x627;
assign c399 = ~x24 & ~x40 & ~x53 & ~x336 & ~x445 & ~x456 & ~x474 & ~x480 & ~x481 & ~x482 & ~x483 & ~x507 & ~x508 & ~x517 & ~x560 & ~x589 & ~x619 & ~x703 & ~x725 & ~x764;
assign c3101 =  x203 &  x455 & ~x479;
assign c3103 =  x568 & ~x109 & ~x137 & ~x157 & ~x215 & ~x243 & ~x308 & ~x408 & ~x749;
assign c3105 = ~x17 & ~x51 & ~x97 & ~x108 & ~x154 & ~x177 & ~x208 & ~x235 & ~x420 & ~x431 & ~x514 & ~x628 & ~x656 & ~x711 & ~x746 & ~x766 & ~x771;
assign c3107 =  x408 & ~x134 & ~x530 & ~x539 & ~x566 & ~x584 & ~x624;
assign c3109 = ~x11 & ~x39 & ~x47 & ~x137 & ~x265 & ~x291 & ~x350 & ~x379 & ~x655 & ~x695 & ~x720 & ~x744 & ~x747 & ~x763;
assign c3111 =  x398 & ~x103 & ~x366 & ~x590 & ~x637 & ~x736;
assign c3113 =  x368 & ~x206 & ~x209 & ~x268 & ~x290 & ~x297 & ~x326 & ~x681 & ~x707;
assign c3115 = ~x3 & ~x47 & ~x54 & ~x137 & ~x410 & ~x521 & ~x532 & ~x552 & ~x553 & ~x555 & ~x580 & ~x612 & ~x638 & ~x667 & ~x670 & ~x676 & ~x702 & ~x781;
assign c3117 =  x432 & ~x501 & ~x617 & ~x635 & ~x638;
assign c3119 =  x439 & ~x16 & ~x18 & ~x19 & ~x379 & ~x386 & ~x747;
assign c3121 =  x484 &  x485 & ~x451 & ~x669 & ~x686 & ~x696;
assign c3123 = ~x0 & ~x54 & ~x198 & ~x280 & ~x281 & ~x329 & ~x471 & ~x472 & ~x474 & ~x475 & ~x498 & ~x502 & ~x717 & ~x718 & ~x744 & ~x746 & ~x749 & ~x757 & ~x761 & ~x764 & ~x772 & ~x774 & ~x775;
assign c3125 =  x314 & ~x22 & ~x102 & ~x130 & ~x159 & ~x219 & ~x530 & ~x735 & ~x770;
assign c3127 = ~x165 & ~x173 & ~x190 & ~x197 & ~x393 & ~x420 & ~x611 & ~x613 & ~x638 & ~x659 & ~x662 & ~x664 & ~x718;
assign c3129 =  x128 &  x319 & ~x473 & ~x607;
assign c3131 = ~x26 & ~x35 & ~x108 & ~x139 & ~x420 & ~x421 & ~x438 & ~x523 & ~x552 & ~x553 & ~x580 & ~x588 & ~x607 & ~x610 & ~x667 & ~x753 & ~x755;
assign c3133 = ~x19 & ~x66 & ~x128 & ~x149 & ~x180 & ~x263 & ~x348 & ~x353 & ~x431 & ~x434 & ~x602 & ~x698;
assign c3135 =  x536 &  x646 & ~x720 & ~x751;
assign c3137 =  x90 & ~x274 & ~x302 & ~x388 & ~x416 & ~x445 & ~x690;
assign c3139 =  x69 & ~x47 & ~x75 & ~x76 & ~x397 & ~x477 & ~x783;
assign c3141 =  x348 & ~x80 & ~x393 & ~x444 & ~x530 & ~x719 & ~x720;
assign c3143 =  x628 &  x689 & ~x162;
assign c3145 = ~x45 & ~x80 & ~x85 & ~x252 & ~x281 & ~x382 & ~x419 & ~x434 & ~x548 & ~x579 & ~x606 & ~x632 & ~x723 & ~x769;
assign c3147 =  x459 & ~x672 & ~x692 & ~x716 & ~x747;
assign c3149 =  x515 &  x541 & ~x481;
assign c3151 =  x343 &  x372 & ~x11 & ~x393 & ~x408;
assign c3153 =  x215 &  x376 & ~x473;
assign c3155 =  x710 & ~x230;
assign c3157 =  x317 &  x318 & ~x530 & ~x551 & ~x580 & ~x581 & ~x583 & ~x588;
assign c3159 =  x179 & ~x164 & ~x246 & ~x483 & ~x510;
assign c3161 =  x149 & ~x294 & ~x421 & ~x473 & ~x559 & ~x684 & ~x736 & ~x740;
assign c3163 = ~x19 & ~x36 & ~x63 & ~x135 & ~x142 & ~x173 & ~x202 & ~x474 & ~x484 & ~x498 & ~x501 & ~x510 & ~x592 & ~x670 & ~x759 & ~x764;
assign c3165 = ~x17 & ~x18 & ~x19 & ~x23 & ~x48 & ~x72 & ~x110 & ~x223 & ~x323 & ~x364 & ~x392 & ~x464 & ~x492 & ~x574 & ~x578 & ~x685 & ~x687 & ~x692 & ~x693 & ~x723 & ~x746 & ~x751 & ~x756 & ~x757 & ~x778 & ~x783;
assign c3167 =  x295 &  x518 & ~x678;
assign c3169 = ~x27 & ~x29 & ~x55 & ~x111 & ~x113 & ~x116 & ~x143 & ~x171 & ~x172 & ~x175 & ~x279 & ~x361 & ~x363 & ~x364 & ~x366 & ~x388 & ~x389 & ~x393 & ~x397 & ~x398 & ~x399 & ~x400 & ~x415 & ~x416 & ~x417 & ~x418 & ~x422 & ~x423 & ~x424 & ~x444 & ~x445 & ~x450 & ~x451 & ~x452 & ~x453 & ~x473 & ~x478 & ~x479 & ~x503 & ~x505 & ~x507 & ~x533 & ~x535 & ~x560 & ~x589 & ~x590 & ~x642 & ~x646 & ~x671 & ~x672 & ~x697 & ~x757 & ~x760 & ~x761;
assign c3171 = ~x35 & ~x252 & ~x383 & ~x412 & ~x416 & ~x417 & ~x440 & ~x441 & ~x459 & ~x499 & ~x502 & ~x503 & ~x525 & ~x527 & ~x528;
assign c3173 = ~x88 & ~x115 & ~x122 & ~x129 & ~x160 & ~x163 & ~x165 & ~x216 & ~x279 & ~x585 & ~x688;
assign c3175 = ~x25 & ~x55 & ~x56 & ~x140 & ~x168 & ~x244 & ~x245 & ~x246 & ~x247 & ~x273 & ~x274 & ~x302 & ~x303 & ~x388 & ~x516 & ~x586 & ~x587 & ~x615 & ~x634 & ~x643 & ~x663 & ~x760;
assign c3177 =  x344 &  x484 & ~x55 & ~x380 & ~x436;
assign c3179 =  x399 & ~x12 & ~x14 & ~x16 & ~x21 & ~x24 & ~x33 & ~x73 & ~x74 & ~x83 & ~x336 & ~x394 & ~x604 & ~x615;
assign c3181 =  x481 & ~x5 & ~x14 & ~x21 & ~x97 & ~x306 & ~x459 & ~x460 & ~x655 & ~x682 & ~x710 & ~x714 & ~x768 & ~x775;
assign c3183 =  x94 & ~x55 & ~x73 & ~x74 & ~x113 & ~x348 & ~x362 & ~x364 & ~x391;
assign c3185 =  x486 & ~x480 & ~x663;
assign c3187 = ~x29 & ~x446 & ~x451 & ~x473 & ~x497 & ~x499 & ~x503 & ~x512 & ~x531 & ~x532 & ~x570 & ~x595 & ~x726 & ~x746 & ~x762 & ~x763 & ~x765 & ~x767;
assign c3189 =  x463 &  x489 &  x515;
assign c3191 = ~x20 & ~x31 & ~x53 & ~x79 & ~x87 & ~x180 & ~x294 & ~x404 & ~x405 & ~x489 & ~x543 & ~x573 & ~x630 & ~x740 & ~x745 & ~x746 & ~x747 & ~x750 & ~x764 & ~x771;
assign c3193 = ~x26 & ~x106 & ~x175 & ~x177 & ~x552 & ~x589 & ~x607 & ~x620 & ~x666 & ~x678 & ~x698;
assign c3195 =  x599 & ~x19 & ~x189;
assign c3197 =  x325 &  x710 & ~x367;
assign c3199 =  x712 & ~x189 & ~x220;
assign c3201 =  x270 & ~x0 & ~x4 & ~x5 & ~x223 & ~x224 & ~x364 & ~x426 & ~x448 & ~x450 & ~x451 & ~x453 & ~x502 & ~x508 & ~x534 & ~x557 & ~x559 & ~x614 & ~x645 & ~x671 & ~x730;
assign c3203 =  x482 &  x591;
assign c3205 =  x569 & ~x375;
assign c3207 = ~x1 & ~x17 & ~x44 & ~x46 & ~x47 & ~x53 & ~x56 & ~x57 & ~x73 & ~x99 & ~x111 & ~x140 & ~x153 & ~x387 & ~x388 & ~x390 & ~x414 & ~x416 & ~x419 & ~x442 & ~x472 & ~x474 & ~x502 & ~x559 & ~x764 & ~x766;
assign c3209 =  x400 & ~x411 & ~x479 & ~x499;
assign c3211 =  x575 &  x576 & ~x79 & ~x111 & ~x164 & ~x167 & ~x559 & ~x615 & ~x700 & ~x708 & ~x767 & ~x768;
assign c3213 =  x299 &  x356 & ~x87 & ~x352 & ~x394 & ~x629;
assign c3217 =  x426 & ~x24 & ~x138 & ~x266 & ~x296 & ~x336 & ~x365 & ~x380 & ~x671 & ~x749;
assign c3219 = ~x12 & ~x72 & ~x128 & ~x129 & ~x131 & ~x132 & ~x158 & ~x248 & ~x250 & ~x278 & ~x322 & ~x364 & ~x378 & ~x752;
assign c3221 =  x373 & ~x47 & ~x103 & ~x465 & ~x501 & ~x617 & ~x643 & ~x669;
assign c3223 =  x65 &  x92 & ~x248;
assign c3225 = ~x17 & ~x21 & ~x271 & ~x356 & ~x474 & ~x498 & ~x499 & ~x500 & ~x530 & ~x557 & ~x558 & ~x559 & ~x586 & ~x624 & ~x651 & ~x652 & ~x735 & ~x764 & ~x769 & ~x770;
assign c3227 = ~x2 & ~x50 & ~x54 & ~x55 & ~x70 & ~x86 & ~x169 & ~x224 & ~x364 & ~x504 & ~x575 & ~x588 & ~x597 & ~x604 & ~x632 & ~x633 & ~x662 & ~x702 & ~x725 & ~x741 & ~x742 & ~x746 & ~x747 & ~x760 & ~x774 & ~x778 & ~x782;
assign c3229 =  x238 &  x296 & ~x35 & ~x148 & ~x734;
assign c3231 =  x489 & ~x162 & ~x585 & ~x719;
assign c3233 = ~x2 & ~x7 & ~x8 & ~x87 & ~x140 & ~x223 & ~x225 & ~x253 & ~x254 & ~x279 & ~x280 & ~x385 & ~x386 & ~x401 & ~x402 & ~x428 & ~x446 & ~x485 & ~x502 & ~x504 & ~x558 & ~x614 & ~x619 & ~x683 & ~x699 & ~x752 & ~x783;
assign c3235 =  x303 &  x474 & ~x553;
assign c3237 =  x458 & ~x508 & ~x719;
assign c3239 = ~x169 & ~x194 & ~x202 & ~x255 & ~x274 & ~x306 & ~x334 & ~x335 & ~x360 & ~x371 & ~x372 & ~x387 & ~x399 & ~x415 & ~x418 & ~x419 & ~x472 & ~x500 & ~x503 & ~x529 & ~x531 & ~x658 & ~x758;
assign c3241 =  x123 &  x124 & ~x23 & ~x75 & ~x102 & ~x145 & ~x425 & ~x559;
assign c3243 = ~x301 & ~x649 & ~x690;
assign c3245 = ~x0 & ~x12 & ~x18 & ~x23 & ~x24 & ~x49 & ~x79 & ~x81 & ~x85 & ~x94 & ~x98 & ~x110 & ~x136 & ~x263 & ~x281 & ~x292 & ~x323 & ~x351 & ~x364 & ~x598 & ~x685 & ~x693 & ~x719 & ~x722 & ~x749 & ~x752 & ~x756;
assign c3247 =  x485 &  x486 & ~x16 & ~x17 & ~x237;
assign c3249 =  x509 &  x563 & ~x294 & ~x351;
assign c3251 = ~x8 & ~x86 & ~x227 & ~x228 & ~x230 & ~x248 & ~x253 & ~x286 & ~x287 & ~x310 & ~x313 & ~x315 & ~x316 & ~x334 & ~x337 & ~x386 & ~x394 & ~x501 & ~x584 & ~x585 & ~x614 & ~x615 & ~x731 & ~x762;
assign c3253 =  x380 &  x516 &  x543;
assign c3255 =  x320 & ~x387 & ~x400 & ~x406 & ~x427 & ~x444 & ~x446;
assign c3257 =  x276 &  x461;
assign c3259 =  x211 &  x374 & ~x61 & ~x88;
assign c3261 =  x66 & ~x46 & ~x47 & ~x55 & ~x112 & ~x420 & ~x421 & ~x587 & ~x670 & ~x727 & ~x728;
assign c3263 = ~x3 & ~x6 & ~x16 & ~x17 & ~x24 & ~x25 & ~x47 & ~x53 & ~x56 & ~x110 & ~x167 & ~x267 & ~x297 & ~x322 & ~x325 & ~x350 & ~x378 & ~x382 & ~x407 & ~x433 & ~x698 & ~x699 & ~x711 & ~x754 & ~x767 & ~x782 & ~x783;
assign c3265 =  x125 & ~x20 & ~x21 & ~x23 & ~x29 & ~x32 & ~x34 & ~x60 & ~x141 & ~x168 & ~x363 & ~x391 & ~x418 & ~x447 & ~x475 & ~x501 & ~x558 & ~x586 & ~x673 & ~x674 & ~x704 & ~x729 & ~x733 & ~x760 & ~x761 & ~x763 & ~x764;
assign c3267 = ~x33 & ~x110 & ~x117 & ~x165 & ~x192 & ~x194 & ~x342 & ~x372 & ~x373 & ~x394 & ~x397 & ~x402 & ~x420 & ~x421 & ~x422 & ~x483 & ~x511 & ~x557 & ~x671 & ~x763;
assign c3269 =  x324 & ~x169 & ~x217 & ~x244 & ~x245 & ~x272 & ~x274 & ~x301 & ~x303 & ~x386 & ~x387 & ~x414 & ~x417;
assign c3271 =  x425 &  x427 & ~x24 & ~x306 & ~x335 & ~x349 & ~x781;
assign c3273 = ~x139 & ~x245 & ~x304 & ~x305 & ~x308 & ~x309 & ~x318 & ~x335 & ~x360 & ~x386 & ~x427 & ~x453 & ~x455 & ~x472 & ~x474;
assign c3275 = ~x0 & ~x4 & ~x16 & ~x98 & ~x125 & ~x245 & ~x275 & ~x305 & ~x364 & ~x475 & ~x606 & ~x720;
assign c3277 = ~x125 & ~x150 & ~x264 & ~x296 & ~x325 & ~x434 & ~x492 & ~x600 & ~x721 & ~x725;
assign c3279 = ~x279 & ~x306 & ~x358 & ~x385 & ~x413 & ~x414 & ~x415 & ~x430 & ~x443 & ~x444 & ~x446 & ~x447 & ~x502 & ~x513 & ~x540 & ~x557 & ~x558 & ~x585 & ~x650 & ~x763 & ~x767 & ~x768;
assign c3281 =  x431 & ~x635 & ~x665 & ~x694 & ~x723 & ~x750;
assign c3283 =  x382 &  x605 & ~x322 & ~x378 & ~x385 & ~x735;
assign c3285 = ~x9 & ~x19 & ~x20 & ~x96 & ~x149 & ~x293 & ~x337 & ~x460 & ~x651 & ~x683 & ~x710 & ~x734 & ~x747 & ~x753 & ~x754 & ~x778;
assign c3287 =  x460 & ~x16 & ~x18 & ~x613;
assign c3289 = ~x61 & ~x199 & ~x247 & ~x273 & ~x286 & ~x287 & ~x311 & ~x316 & ~x332 & ~x344 & ~x360 & ~x372;
assign c3291 = ~x26 & ~x29 & ~x138 & ~x216 & ~x278 & ~x334 & ~x366 & ~x413 & ~x640 & ~x728 & ~x746 & ~x767 & ~x774;
assign c3293 = ~x23 & ~x45 & ~x60 & ~x199 & ~x224 & ~x226 & ~x303 & ~x474 & ~x516 & ~x544 & ~x575 & ~x634 & ~x718 & ~x720 & ~x747 & ~x782;
assign c3295 =  x403 & ~x691 & ~x692 & ~x693 & ~x694 & ~x721 & ~x722 & ~x751 & ~x776 & ~x777 & ~x779 & ~x780;
assign c3297 =  x659 & ~x426 & ~x447 & ~x506 & ~x739;
assign c3299 = ~x22 & ~x25 & ~x27 & ~x115 & ~x335 & ~x389 & ~x545 & ~x559 & ~x635 & ~x637 & ~x663 & ~x690 & ~x693 & ~x736 & ~x747 & ~x749 & ~x760 & ~x777;
assign c3301 =  x426 & ~x23 & ~x108 & ~x266 & ~x337 & ~x636 & ~x722;
assign c3303 = ~x202 & ~x203 & ~x288 & ~x330 & ~x334 & ~x358 & ~x360 & ~x453 & ~x485 & ~x488;
assign c3305 =  x631 & ~x137 & ~x250 & ~x422 & ~x567 & ~x587 & ~x735 & ~x767;
assign c3307 =  x369 &  x398 & ~x14 & ~x336 & ~x365 & ~x392 & ~x406 & ~x658 & ~x682 & ~x690 & ~x736 & ~x739 & ~x764 & ~x774;
assign c3309 =  x370 &  x455 & ~x17 & ~x394 & ~x422 & ~x756;
assign c3311 = ~x17 & ~x19 & ~x45 & ~x84 & ~x165 & ~x185 & ~x193 & ~x194 & ~x222 & ~x268 & ~x297 & ~x325 & ~x353 & ~x392 & ~x409 & ~x521;
assign c3313 = ~x2 & ~x12 & ~x21 & ~x25 & ~x34 & ~x113 & ~x115 & ~x139 & ~x171 & ~x434 & ~x547 & ~x634 & ~x662 & ~x719 & ~x741 & ~x750 & ~x776 & ~x777;
assign c3315 = ~x15 & ~x20 & ~x24 & ~x99 & ~x237 & ~x280 & ~x296 & ~x309 & ~x319 & ~x392 & ~x407 & ~x654 & ~x710 & ~x712 & ~x741 & ~x753 & ~x767 & ~x780;
assign c3317 = ~x15 & ~x23 & ~x38 & ~x65 & ~x96 & ~x123 & ~x265 & ~x319 & ~x353 & ~x354 & ~x488 & ~x603 & ~x655 & ~x726;
assign c3319 =  x516;
assign c3321 = ~x5 & ~x60 & ~x85 & ~x307 & ~x362 & ~x363 & ~x391 & ~x467 & ~x609 & ~x633 & ~x640 & ~x666 & ~x764 & ~x765 & ~x766 & ~x782;
assign c3323 =  x346 & ~x328 & ~x359 & ~x529;
assign c3325 =  x319 &  x321 & ~x2 & ~x506 & ~x552 & ~x565 & ~x585 & ~x586;
assign c3327 = ~x10 & ~x25 & ~x40 & ~x108 & ~x180 & ~x239 & ~x264 & ~x268 & ~x296 & ~x380 & ~x734 & ~x766 & ~x768;
assign c3329 =  x595 & ~x44 & ~x235 & ~x297 & ~x353 & ~x360 & ~x770;
assign c3331 =  x155 & ~x107 & ~x678 & ~x705;
assign c3333 = ~x2 & ~x16 & ~x17 & ~x19 & ~x44 & ~x194 & ~x277 & ~x282 & ~x301 & ~x302 & ~x309 & ~x333 & ~x337 & ~x361 & ~x362 & ~x388 & ~x418 & ~x419 & ~x473 & ~x691 & ~x783;
assign c3335 =  x520 &  x547 &  x638;
assign c3337 = ~x6 & ~x29 & ~x222 & ~x273 & ~x280 & ~x308 & ~x329 & ~x331 & ~x390 & ~x420 & ~x442 & ~x446 & ~x447 & ~x473 & ~x476 & ~x500 & ~x516 & ~x630 & ~x746 & ~x775;
assign c3339 = ~x104 & ~x133 & ~x454;
assign c3341 = ~x8 & ~x28 & ~x29 & ~x141 & ~x363 & ~x416 & ~x417 & ~x418 & ~x419 & ~x444 & ~x474 & ~x483 & ~x503 & ~x537 & ~x538 & ~x562 & ~x589 & ~x644 & ~x651 & ~x703 & ~x708 & ~x734 & ~x736 & ~x738 & ~x759 & ~x767;
assign c3343 =  x151 &  x714 & ~x103 & ~x563 & ~x591;
assign c3345 = ~x29 & ~x39 & ~x40 & ~x95 & ~x123 & ~x264 & ~x291 & ~x321 & ~x349 & ~x351 & ~x352 & ~x377 & ~x378 & ~x408 & ~x460 & ~x572 & ~x573 & ~x721 & ~x722 & ~x770;
assign c3347 = ~x163 & ~x165 & ~x220 & ~x250 & ~x538 & ~x539 & ~x565 & ~x770;
assign c3349 = ~x17 & ~x384 & ~x495 & ~x498 & ~x534 & ~x563 & ~x581 & ~x585;
assign c3351 =  x469 & ~x17 & ~x360 & ~x603 & ~x692;
assign c3353 = ~x35 & ~x63 & ~x201 & ~x316 & ~x341 & ~x343 & ~x361 & ~x363 & ~x372 & ~x399 & ~x400 & ~x425 & ~x446 & ~x455 & ~x505 & ~x534 & ~x646 & ~x675 & ~x730 & ~x760;
assign c3355 =  x177 &  x456 & ~x40 & ~x778;
assign c3357 =  x120 &  x483 &  x484;
assign c3359 =  x152 & ~x47 & ~x75 & ~x170 & ~x419 & ~x449 & ~x479 & ~x480 & ~x506 & ~x532 & ~x533;
assign c3361 =  x206 &  x207 & ~x23 & ~x26 & ~x80 & ~x86 & ~x112 & ~x137 & ~x168 & ~x225 & ~x363 & ~x452 & ~x453 & ~x454 & ~x563 & ~x643 & ~x673 & ~x759 & ~x760 & ~x762;
assign c3363 =  x215 &  x262 & ~x582 & ~x610;
assign c3365 = ~x14 & ~x95 & ~x109 & ~x211 & ~x238 & ~x294 & ~x349 & ~x375 & ~x543 & ~x544 & ~x693 & ~x750;
assign c3367 =  x288 &  x484 &  x485 & ~x559;
assign c3369 =  x484 & ~x263 & ~x632 & ~x633 & ~x691 & ~x718 & ~x749 & ~x765;
assign c3371 = ~x97 & ~x512 & ~x540 & ~x541 & ~x567 & ~x622 & ~x677 & ~x680 & ~x732 & ~x736 & ~x760;
assign c3373 = ~x11 & ~x47 & ~x48 & ~x73 & ~x351 & ~x391 & ~x406 & ~x467 & ~x504 & ~x606 & ~x638 & ~x695 & ~x763;
assign c3375 =  x459 &  x460 & ~x721;
assign c3377 =  x258 & ~x335 & ~x379 & ~x710 & ~x737;
assign c3379 =  x404 & ~x390 & ~x454 & ~x473 & ~x481 & ~x500 & ~x504 & ~x505 & ~x506 & ~x530;
assign c3381 =  x729;
assign c3383 =  x297 & ~x0 & ~x335 & ~x399 & ~x420 & ~x422 & ~x423 & ~x425 & ~x427 & ~x445 & ~x451 & ~x452 & ~x534 & ~x562 & ~x617 & ~x643;
assign c3385 = ~x24 & ~x27 & ~x63 & ~x73 & ~x74 & ~x223 & ~x338 & ~x440 & ~x474 & ~x529 & ~x554 & ~x582 & ~x584 & ~x756;
assign c3387 = ~x0 & ~x22 & ~x59 & ~x88 & ~x111 & ~x453 & ~x454 & ~x472 & ~x474 & ~x479 & ~x481 & ~x500 & ~x501 & ~x530 & ~x532 & ~x534 & ~x559 & ~x561 & ~x562 & ~x563 & ~x564 & ~x573;
assign c3389 =  x389 & ~x720;
assign c3391 = ~x32 & ~x35 & ~x54 & ~x81 & ~x115 & ~x139 & ~x440 & ~x467 & ~x496 & ~x498 & ~x499 & ~x500 & ~x502 & ~x527 & ~x553 & ~x582 & ~x610 & ~x611 & ~x650 & ~x733;
assign c3393 =  x543 & ~x19 & ~x50 & ~x108 & ~x135 & ~x165 & ~x615 & ~x642;
assign c3395 =  x149 &  x428 &  x456 & ~x15;
assign c3397 =  x343 &  x455 &  x565 & ~x460 & ~x487 & ~x754;
assign c3399 = ~x21 & ~x27 & ~x79 & ~x81 & ~x252 & ~x448 & ~x495 & ~x496 & ~x497 & ~x502 & ~x524 & ~x528 & ~x530 & ~x552 & ~x557 & ~x558 & ~x560 & ~x580 & ~x581 & ~x582 & ~x585 & ~x592 & ~x610 & ~x611 & ~x613 & ~x614 & ~x618 & ~x642 & ~x646 & ~x670 & ~x673 & ~x755;
assign c3401 =  x709 & ~x313 & ~x370 & ~x397;
assign c3403 =  x69 & ~x104 & ~x508;
assign c3405 =  x517 & ~x136 & ~x189 & ~x279 & ~x614 & ~x749;
assign c3407 =  x535 & ~x295 & ~x323 & ~x336 & ~x380 & ~x433 & ~x436 & ~x604 & ~x752 & ~x778;
assign c3409 = ~x0 & ~x1 & ~x2 & ~x15 & ~x18 & ~x20 & ~x23 & ~x24 & ~x55 & ~x81 & ~x108 & ~x112 & ~x277 & ~x278 & ~x279 & ~x306 & ~x438 & ~x587 & ~x617 & ~x642 & ~x645 & ~x671 & ~x693 & ~x700 & ~x707 & ~x723 & ~x736 & ~x749 & ~x750 & ~x751 & ~x753 & ~x762 & ~x764 & ~x775 & ~x781 & ~x782;
assign c3411 =  x438 & ~x15 & ~x61 & ~x129 & ~x162 & ~x733;
assign c3413 = ~x361 & ~x386 & ~x390 & ~x413 & ~x415 & ~x451 & ~x473 & ~x477 & ~x501 & ~x504 & ~x553 & ~x581 & ~x597 & ~x680 & ~x707 & ~x737 & ~x763 & ~x768;
assign c3415 =  x228 &  x425 & ~x18 & ~x337 & ~x764 & ~x768;
assign c3417 =  x578 & ~x33 & ~x112 & ~x277 & ~x304 & ~x332 & ~x359 & ~x379 & ~x436 & ~x473 & ~x656 & ~x765;
assign c3419 =  x170 &  x481 &  x483;
assign c3421 = ~x27 & ~x34 & ~x90 & ~x222 & ~x248 & ~x250 & ~x255 & ~x285 & ~x314 & ~x315 & ~x316 & ~x455 & ~x477 & ~x482 & ~x613 & ~x732;
assign c3423 =  x230 &  x257 & ~x23 & ~x39 & ~x123 & ~x211 & ~x239 & ~x336 & ~x680;
assign c3425 =  x370 & ~x17 & ~x54 & ~x81 & ~x150 & ~x308 & ~x336 & ~x350 & ~x604 & ~x680;
assign c3427 = ~x112 & ~x168 & ~x196 & ~x225 & ~x276 & ~x304 & ~x334 & ~x335 & ~x336 & ~x388 & ~x502 & ~x587 & ~x606 & ~x629 & ~x631 & ~x632 & ~x634 & ~x635 & ~x662 & ~x663 & ~x691 & ~x692 & ~x721;
assign c3429 =  x109 & ~x332 & ~x390;
assign c3431 =  x455 & ~x53 & ~x125 & ~x239 & ~x324 & ~x351 & ~x380;
assign c3433 = ~x230 & ~x335 & ~x361 & ~x373 & ~x392 & ~x399 & ~x426 & ~x483 & ~x507 & ~x619 & ~x764 & ~x765;
assign c3435 = ~x52 & ~x169 & ~x224 & ~x253 & ~x323 & ~x364 & ~x373 & ~x380 & ~x519 & ~x520 & ~x574 & ~x576 & ~x720 & ~x765 & ~x781;
assign c3437 =  x265 &  x430 & ~x21 & ~x30 & ~x196 & ~x475 & ~x588;
assign c3439 =  x379 &  x712;
assign c3441 = ~x17 & ~x28 & ~x47 & ~x54 & ~x72 & ~x116 & ~x149 & ~x234 & ~x265 & ~x662 & ~x720 & ~x742 & ~x756;
assign c3443 =  x343 &  x426 &  x508 & ~x153 & ~x324 & ~x449;
assign c3445 = ~x16 & ~x47 & ~x83 & ~x123 & ~x165 & ~x205 & ~x264 & ~x406 & ~x407 & ~x548 & ~x601 & ~x771 & ~x777;
assign c3447 =  x464 & ~x144 & ~x222 & ~x453 & ~x481 & ~x706 & ~x764;
assign c3449 = ~x50 & ~x128 & ~x268 & ~x317 & ~x336 & ~x467 & ~x525 & ~x756;
assign c3451 =  x374 & ~x419 & ~x446 & ~x470 & ~x501 & ~x516 & ~x588;
assign c3453 = ~x14 & ~x19 & ~x20 & ~x26 & ~x45 & ~x47 & ~x123 & ~x223 & ~x308 & ~x322 & ~x347 & ~x351 & ~x364 & ~x374 & ~x487 & ~x489 & ~x514 & ~x571 & ~x684 & ~x686 & ~x699 & ~x700 & ~x740 & ~x751 & ~x752 & ~x753 & ~x771 & ~x772 & ~x779;
assign c3455 =  x177 &  x456 & ~x424 & ~x479 & ~x770;
assign c3457 = ~x43 & ~x45 & ~x125 & ~x126 & ~x277 & ~x309 & ~x331 & ~x682 & ~x683 & ~x689 & ~x699 & ~x716 & ~x718 & ~x772;
assign c3459 =  x155 & ~x47 & ~x84 & ~x104 & ~x131 & ~x132 & ~x133 & ~x134 & ~x135 & ~x504 & ~x586 & ~x706 & ~x731 & ~x761;
assign c3461 = ~x17 & ~x18 & ~x290 & ~x322 & ~x348 & ~x364 & ~x517 & ~x652 & ~x680 & ~x682 & ~x737 & ~x741 & ~x742 & ~x750 & ~x769 & ~x770 & ~x776 & ~x778;
assign c3463 =  x378 &  x573 & ~x411 & ~x762;
assign c3465 = ~x394 & ~x586;
assign c3467 = ~x17 & ~x18 & ~x44 & ~x53 & ~x57 & ~x125 & ~x126 & ~x140 & ~x168 & ~x180 & ~x225 & ~x337 & ~x557 & ~x558 & ~x600 & ~x718 & ~x737 & ~x739 & ~x740 & ~x741 & ~x742 & ~x743 & ~x744 & ~x764 & ~x771 & ~x772 & ~x773;
assign c3469 =  x661 & ~x116 & ~x136 & ~x454 & ~x580 & ~x589 & ~x732;
assign c3471 = ~x8 & ~x12 & ~x24 & ~x140 & ~x167 & ~x470 & ~x474 & ~x497 & ~x498 & ~x499 & ~x500 & ~x511 & ~x512 & ~x529 & ~x555 & ~x556 & ~x558 & ~x559 & ~x611 & ~x612 & ~x617 & ~x645 & ~x646 & ~x647 & ~x649 & ~x668 & ~x673 & ~x676 & ~x705 & ~x735 & ~x761 & ~x764;
assign c3473 =  x479 & ~x70 & ~x180 & ~x379 & ~x749 & ~x776;
assign c3475 = ~x19 & ~x56 & ~x59 & ~x138 & ~x166 & ~x300 & ~x441 & ~x502 & ~x532 & ~x533 & ~x553 & ~x555 & ~x581 & ~x582 & ~x583 & ~x585 & ~x587 & ~x610 & ~x640 & ~x641 & ~x667 & ~x671 & ~x707 & ~x723 & ~x759 & ~x764 & ~x783;
assign c3477 =  x509 & ~x88 & ~x350 & ~x691 & ~x692 & ~x693 & ~x695 & ~x722 & ~x733 & ~x746 & ~x751 & ~x753 & ~x767 & ~x768 & ~x769 & ~x776;
assign c3479 = ~x26 & ~x415 & ~x419 & ~x443 & ~x473 & ~x477 & ~x479 & ~x499 & ~x500 & ~x541 & ~x557 & ~x568 & ~x623 & ~x644 & ~x650 & ~x654 & ~x711 & ~x737 & ~x756 & ~x762 & ~x763 & ~x765 & ~x766 & ~x769;
assign c3481 = ~x8 & ~x29 & ~x72 & ~x264 & ~x323 & ~x376 & ~x432 & ~x521 & ~x725 & ~x743 & ~x762 & ~x767;
assign c3483 =  x296 &  x324 &  x464 & ~x44 & ~x707 & ~x708;
assign c3485 = ~x26 & ~x359 & ~x361 & ~x399 & ~x401 & ~x402 & ~x403 & ~x417 & ~x430 & ~x474 & ~x475 & ~x512 & ~x536 & ~x557 & ~x586 & ~x645 & ~x646 & ~x648 & ~x649 & ~x677 & ~x680 & ~x703 & ~x704 & ~x711 & ~x730 & ~x735 & ~x760 & ~x765 & ~x778;
assign c3487 =  x376 &  x596 & ~x46 & ~x746;
assign c3489 =  x455 &  x537 & ~x193 & ~x476 & ~x489 & ~x514;
assign c3491 =  x267 & ~x173 & ~x196 & ~x225 & ~x248 & ~x607 & ~x759;
assign c3493 = ~x25 & ~x28 & ~x53 & ~x84 & ~x88 & ~x113 & ~x115 & ~x144 & ~x168 & ~x420 & ~x455 & ~x482 & ~x484 & ~x503 & ~x506 & ~x509 & ~x527 & ~x528 & ~x529 & ~x532 & ~x557 & ~x559 & ~x569 & ~x596 & ~x597 & ~x616 & ~x623 & ~x624 & ~x644 & ~x650 & ~x654 & ~x668 & ~x670 & ~x671 & ~x679 & ~x680 & ~x705 & ~x706 & ~x707 & ~x708 & ~x736 & ~x738 & ~x759 & ~x760 & ~x762 & ~x763 & ~x764 & ~x767;
assign c3495 = ~x9 & ~x15 & ~x23 & ~x30 & ~x181 & ~x209 & ~x322 & ~x379 & ~x544 & ~x548 & ~x631 & ~x722 & ~x723 & ~x743 & ~x745 & ~x747 & ~x758 & ~x771 & ~x776;
assign c3497 = ~x18 & ~x46 & ~x48 & ~x222 & ~x265 & ~x307 & ~x323 & ~x347 & ~x352 & ~x495 & ~x640 & ~x778;
assign c3499 =  x388 & ~x42 & ~x120 & ~x127 & ~x149 & ~x552 & ~x597 & ~x693;
assign c40 =  x204 & ~x29 & ~x44 & ~x45 & ~x72 & ~x74 & ~x100 & ~x170 & ~x344 & ~x398 & ~x451 & ~x615 & ~x699 & ~x743;
assign c42 =  x311 &  x365 & ~x11 & ~x39 & ~x97 & ~x101 & ~x559 & ~x608 & ~x613 & ~x615 & ~x668 & ~x669 & ~x755;
assign c44 =  x491 & ~x4 & ~x15 & ~x31 & ~x82 & ~x109 & ~x143 & ~x166 & ~x169 & ~x192 & ~x200 & ~x275 & ~x307 & ~x322 & ~x453 & ~x454 & ~x504 & ~x532 & ~x643 & ~x726 & ~x756;
assign c46 =  x442 & ~x103 & ~x140 & ~x401 & ~x426 & ~x478 & ~x506 & ~x532 & ~x589 & ~x643 & ~x645 & ~x751 & ~x778 & ~x780;
assign c48 =  x152 &  x382 &  x411 & ~x18 & ~x22 & ~x46 & ~x49 & ~x75 & ~x278 & ~x279 & ~x643 & ~x699;
assign c410 = ~x24 & ~x25 & ~x53 & ~x55 & ~x60 & ~x86 & ~x112 & ~x113 & ~x117 & ~x185 & ~x224 & ~x252 & ~x279 & ~x304 & ~x311 & ~x337 & ~x338 & ~x423 & ~x474 & ~x488 & ~x500 & ~x504 & ~x528 & ~x560 & ~x563 & ~x587 & ~x590 & ~x613 & ~x624 & ~x641 & ~x643 & ~x650 & ~x670 & ~x694 & ~x699 & ~x702 & ~x703 & ~x727 & ~x735 & ~x761 & ~x765 & ~x769 & ~x778;
assign c412 =  x582 & ~x47 & ~x163 & ~x447 & ~x503 & ~x532 & ~x563 & ~x619 & ~x757;
assign c414 =  x653 &  x681 & ~x25 & ~x27 & ~x29 & ~x83 & ~x86 & ~x98 & ~x197 & ~x224 & ~x411 & ~x439 & ~x692 & ~x726 & ~x757 & ~x763 & ~x774 & ~x780 & ~x781;
assign c416 =  x603 &  x631 &  x685 & ~x75 & ~x482 & ~x504 & ~x507 & ~x600;
assign c418 =  x150 & ~x4 & ~x12 & ~x72 & ~x332 & ~x389 & ~x392 & ~x417 & ~x447 & ~x539 & ~x557 & ~x585 & ~x680 & ~x741;
assign c420 =  x146 & ~x19 & ~x53 & ~x111 & ~x137 & ~x156 & ~x157 & ~x400 & ~x455 & ~x664 & ~x700 & ~x719 & ~x748 & ~x756 & ~x758 & ~x759;
assign c422 =  x181 &  x208 &  x235 &  x688 & ~x461;
assign c424 = ~x2 & ~x8 & ~x9 & ~x19 & ~x21 & ~x22 & ~x23 & ~x27 & ~x29 & ~x30 & ~x32 & ~x45 & ~x49 & ~x51 & ~x52 & ~x54 & ~x56 & ~x81 & ~x85 & ~x86 & ~x87 & ~x108 & ~x109 & ~x114 & ~x115 & ~x137 & ~x138 & ~x139 & ~x140 & ~x168 & ~x195 & ~x197 & ~x222 & ~x223 & ~x225 & ~x246 & ~x273 & ~x274 & ~x299 & ~x302 & ~x308 & ~x329 & ~x330 & ~x331 & ~x332 & ~x337 & ~x387 & ~x388 & ~x417 & ~x474 & ~x475 & ~x502 & ~x503 & ~x504 & ~x531 & ~x586 & ~x587 & ~x588 & ~x616 & ~x644 & ~x675 & ~x676 & ~x719 & ~x729 & ~x732 & ~x746 & ~x747 & ~x749 & ~x755 & ~x757 & ~x771 & ~x773 & ~x775 & ~x777 & ~x783;
assign c426 = ~x305 & ~x364 & ~x366 & ~x440 & ~x467 & ~x476 & ~x477 & ~x494 & ~x502 & ~x522 & ~x531 & ~x558 & ~x605 & ~x625 & ~x652 & ~x661 & ~x755 & ~x760 & ~x765 & ~x777;
assign c428 =  x597 &  x625 &  x651 & ~x36 & ~x52 & ~x136 & ~x198 & ~x225 & ~x634 & ~x754;
assign c430 =  x123 &  x177 & ~x16 & ~x84 & ~x114 & ~x142 & ~x168 & ~x252 & ~x398 & ~x448 & ~x533 & ~x615 & ~x616 & ~x618 & ~x619 & ~x707 & ~x708 & ~x725 & ~x731 & ~x733 & ~x751 & ~x754 & ~x755 & ~x756 & ~x760;
assign c432 =  x630 &  x685 &  x709 &  x737 & ~x142 & ~x670 & ~x729 & ~x756;
assign c434 =  x283 & ~x11 & ~x13 & ~x28 & ~x56 & ~x132 & ~x139 & ~x239 & ~x252 & ~x491 & ~x671;
assign c436 =  x652 & ~x14 & ~x42 & ~x87 & ~x459 & ~x633;
assign c438 =  x680 &  x783;
assign c440 =  x459 & ~x29 & ~x57 & ~x81 & ~x112 & ~x198 & ~x280 & ~x401 & ~x481 & ~x489 & ~x534 & ~x535 & ~x617;
assign c442 =  x27;
assign c444 =  x756;
assign c446 =  x97 &  x151 &  x152 &  x206 & ~x219 & ~x293 & ~x294;
assign c448 = ~x45 & ~x47 & ~x59 & ~x108 & ~x142 & ~x166 & ~x246 & ~x305 & ~x418 & ~x532 & ~x587 & ~x619 & ~x642 & ~x648 & ~x672 & ~x678 & ~x685 & ~x689 & ~x711 & ~x713 & ~x735 & ~x737 & ~x738 & ~x740 & ~x765 & ~x781;
assign c450 =  x547 & ~x23 & ~x54 & ~x99 & ~x130 & ~x195 & ~x373 & ~x399 & ~x400 & ~x588 & ~x673 & ~x694 & ~x699 & ~x700 & ~x769;
assign c452 =  x323 & ~x0 & ~x81 & ~x140 & ~x168 & ~x238 & ~x555 & ~x608 & ~x615 & ~x635 & ~x662 & ~x663 & ~x691 & ~x757 & ~x771 & ~x776 & ~x783;
assign c454 =  x263 &  x318 & ~x376 & ~x587 & ~x600 & ~x707 & ~x753 & ~x767 & ~x776;
assign c456 =  x637 & ~x103 & ~x350 & ~x534 & ~x564;
assign c458 =  x337 &  x599;
assign c460 =  x234 &  x566 & ~x224 & ~x308 & ~x447 & ~x667 & ~x669 & ~x670 & ~x699 & ~x749 & ~x754 & ~x762 & ~x778 & ~x779;
assign c462 = ~x91 & ~x185 & ~x277 & ~x308 & ~x414 & ~x421 & ~x499 & ~x596 & ~x607 & ~x690 & ~x745 & ~x746 & ~x767 & ~x777;
assign c464 =  x125 & ~x4 & ~x86 & ~x278 & ~x349 & ~x392 & ~x432 & ~x543 & ~x560 & ~x588 & ~x709 & ~x731 & ~x734 & ~x737 & ~x761;
assign c466 =  x493 &  x660 & ~x45 & ~x46 & ~x462 & ~x540 & ~x725;
assign c468 =  x711 & ~x2 & ~x76 & ~x77 & ~x104 & ~x105 & ~x111 & ~x112 & ~x139 & ~x161 & ~x213 & ~x217 & ~x276 & ~x277 & ~x306 & ~x504 & ~x716 & ~x769;
assign c470 =  x655 &  x709 & ~x27 & ~x55 & ~x71 & ~x111 & ~x170 & ~x224 & ~x714 & ~x742;
assign c472 =  x283 &  x338 & ~x97 & ~x604;
assign c474 =  x66 &  x358 & ~x397;
assign c476 =  x148 &  x175 & ~x18 & ~x23 & ~x30 & ~x46 & ~x70 & ~x72 & ~x102 & ~x115 & ~x129 & ~x447 & ~x476 & ~x505 & ~x562 & ~x645 & ~x664 & ~x672 & ~x696 & ~x729;
assign c478 = ~x180 & ~x236 & ~x298 & ~x456 & ~x466 & ~x522 & ~x587 & ~x605 & ~x615 & ~x700 & ~x715 & ~x743 & ~x771;
assign c480 =  x234 &  x553 & ~x115 & ~x281 & ~x295 & ~x446;
assign c482 =  x231 &  x257 & ~x13 & ~x27 & ~x28 & ~x29 & ~x46 & ~x55 & ~x71 & ~x72 & ~x73 & ~x103 & ~x113 & ~x167 & ~x195 & ~x197 & ~x420 & ~x426 & ~x453 & ~x670 & ~x671 & ~x725 & ~x726 & ~x728 & ~x755;
assign c484 =  x179 &  x263 & ~x4 & ~x14 & ~x224 & ~x418 & ~x452 & ~x618 & ~x643 & ~x646 & ~x750 & ~x758 & ~x763;
assign c486 =  x177 &  x575 &  x659 & ~x238 & ~x588 & ~x781;
assign c488 = ~x11 & ~x12 & ~x30 & ~x40 & ~x43 & ~x70 & ~x98 & ~x100 & ~x101 & ~x127 & ~x194 & ~x197 & ~x199 & ~x221 & ~x222 & ~x225 & ~x278 & ~x362 & ~x447 & ~x559 & ~x592 & ~x614 & ~x616 & ~x622 & ~x672 & ~x731;
assign c490 = ~x0 & ~x183 & ~x237 & ~x320 & ~x329 & ~x430 & ~x442 & ~x471 & ~x475 & ~x486 & ~x501 & ~x503 & ~x556 & ~x700 & ~x728 & ~x758 & ~x759;
assign c492 = ~x9 & ~x11 & ~x30 & ~x56 & ~x57 & ~x81 & ~x97 & ~x111 & ~x138 & ~x167 & ~x270 & ~x271 & ~x274 & ~x298 & ~x300 & ~x301 & ~x302 & ~x327 & ~x356 & ~x390 & ~x549 & ~x729 & ~x756 & ~x758 & ~x773;
assign c494 =  x655 & ~x55 & ~x57 & ~x71 & ~x82 & ~x98 & ~x139 & ~x167 & ~x195 & ~x468 & ~x559 & ~x578 & ~x606 & ~x615 & ~x634 & ~x644 & ~x661 & ~x672 & ~x727;
assign c496 =  x470 &  x625 &  x653 & ~x22 & ~x50 & ~x169 & ~x517 & ~x670 & ~x699 & ~x727 & ~x755 & ~x781 & ~x783;
assign c498 = ~x52 & ~x59 & ~x67 & ~x95 & ~x169 & ~x243 & ~x280 & ~x327 & ~x335 & ~x431 & ~x545 & ~x572 & ~x605 & ~x752 & ~x757;
assign c4100 =  x654 &  x681 & ~x71 & ~x316 & ~x743 & ~x770;
assign c4102 = ~x12 & ~x56 & ~x72 & ~x167 & ~x182 & ~x209 & ~x383 & ~x410 & ~x411 & ~x430 & ~x438 & ~x441 & ~x457 & ~x466 & ~x469 & ~x501 & ~x557 & ~x558 & ~x615 & ~x700;
assign c4104 =  x66 &  x95 & ~x4 & ~x22 & ~x75 & ~x76 & ~x87 & ~x143 & ~x318 & ~x399;
assign c4106 = ~x6 & ~x35 & ~x48 & ~x59 & ~x83 & ~x92 & ~x141 & ~x169 & ~x251 & ~x362 & ~x388 & ~x489 & ~x504 & ~x533 & ~x544 & ~x626 & ~x652 & ~x679 & ~x726 & ~x750 & ~x756 & ~x762;
assign c4108 =  x179 & ~x0 & ~x2 & ~x16 & ~x24 & ~x28 & ~x30 & ~x32 & ~x52 & ~x59 & ~x85 & ~x88 & ~x110 & ~x168 & ~x197 & ~x223 & ~x278 & ~x282 & ~x304 & ~x306 & ~x310 & ~x332 & ~x339 & ~x359 & ~x389 & ~x391 & ~x392 & ~x394 & ~x395 & ~x416 & ~x418 & ~x423 & ~x444 & ~x445 & ~x447 & ~x448 & ~x472 & ~x474 & ~x503 & ~x529 & ~x530 & ~x532 & ~x586 & ~x653 & ~x654 & ~x666 & ~x680 & ~x693 & ~x694 & ~x699 & ~x707 & ~x710 & ~x724 & ~x727 & ~x728 & ~x736 & ~x737 & ~x738 & ~x749 & ~x750 & ~x755 & ~x763 & ~x765 & ~x782;
assign c4110 =  x400 & ~x196 & ~x363 & ~x385 & ~x415 & ~x416 & ~x417 & ~x431 & ~x470 & ~x486 & ~x499 & ~x514 & ~x529 & ~x583 & ~x764;
assign c4112 =  x0;
assign c4114 =  x631 & ~x101 & ~x239 & ~x334 & ~x405 & ~x416 & ~x420 & ~x755;
assign c4116 =  x659 & ~x247 & ~x277 & ~x278 & ~x280 & ~x433 & ~x489 & ~x569 & ~x617 & ~x652 & ~x673 & ~x680 & ~x697 & ~x698 & ~x726 & ~x763;
assign c4118 =  x687 & ~x23 & ~x91 & ~x214 & ~x280 & ~x421 & ~x442 & ~x461 & ~x541;
assign c4120 = ~x28 & ~x53 & ~x60 & ~x112 & ~x115 & ~x168 & ~x281 & ~x283 & ~x307 & ~x309 & ~x311 & ~x335 & ~x336 & ~x360 & ~x361 & ~x365 & ~x387 & ~x389 & ~x390 & ~x414 & ~x418 & ~x441 & ~x448 & ~x460 & ~x471 & ~x500 & ~x515 & ~x526 & ~x531 & ~x532 & ~x534 & ~x570 & ~x581 & ~x583 & ~x585 & ~x588 & ~x590 & ~x597 & ~x608 & ~x615 & ~x668 & ~x672 & ~x673 & ~x693 & ~x721 & ~x725 & ~x754 & ~x755 & ~x757 & ~x761 & ~x765 & ~x779 & ~x780 & ~x782;
assign c4122 =  x180 &  x233 &  x438 & ~x391 & ~x406 & ~x614 & ~x752;
assign c4124 =  x577 &  x660 &  x687 & ~x72 & ~x85 & ~x172 & ~x505 & ~x563 & ~x588 & ~x595;
assign c4126 =  x376 & ~x43 & ~x169 & ~x197 & ~x379 & ~x409 & ~x718 & ~x719 & ~x727;
assign c4128 =  x93 &  x599 &  x626 & ~x197 & ~x224 & ~x409 & ~x465 & ~x503 & ~x693 & ~x776;
assign c4130 =  x180 &  x692;
assign c4132 =  x209 &  x292 & ~x25 & ~x52 & ~x79 & ~x138 & ~x188 & ~x217 & ~x275 & ~x405 & ~x458 & ~x486;
assign c4134 =  x147 & ~x16 & ~x43 & ~x101 & ~x141 & ~x168 & ~x196 & ~x197 & ~x252 & ~x280 & ~x447 & ~x534 & ~x561 & ~x588 & ~x589 & ~x614 & ~x646 & ~x727 & ~x732 & ~x758 & ~x763 & ~x770;
assign c4136 =  x97 & ~x256 & ~x349 & ~x530 & ~x618 & ~x677 & ~x700;
assign c4138 =  x94 &  x203 & ~x19 & ~x73 & ~x142 & ~x170 & ~x197 & ~x343 & ~x344 & ~x503 & ~x642 & ~x698;
assign c4140 =  x497 & ~x51 & ~x190 & ~x228 & ~x245 & ~x253 & ~x254 & ~x445 & ~x447 & ~x522 & ~x550 & ~x645 & ~x670;
assign c4142 =  x230 &  x312 & ~x12 & ~x26 & ~x48 & ~x69 & ~x75 & ~x77 & ~x81 & ~x280 & ~x452 & ~x615;
assign c4144 = ~x4 & ~x9 & ~x109 & ~x186 & ~x187 & ~x217 & ~x246 & ~x278 & ~x281 & ~x301 & ~x402 & ~x454 & ~x482 & ~x483 & ~x680 & ~x745 & ~x773;
assign c4146 =  x683 &  x709 & ~x31 & ~x57 & ~x113 & ~x114 & ~x137 & ~x141 & ~x167 & ~x169 & ~x191 & ~x484 & ~x717;
assign c4148 =  x494 &  x661 & ~x26 & ~x46 & ~x434 & ~x461 & ~x532 & ~x559 & ~x588 & ~x642 & ~x698 & ~x754;
assign c4150 = ~x27 & ~x52 & ~x60 & ~x82 & ~x167 & ~x180 & ~x183 & ~x184 & ~x210 & ~x211 & ~x237 & ~x239 & ~x325 & ~x383 & ~x440 & ~x441 & ~x469 & ~x633 & ~x661 & ~x756 & ~x760;
assign c4152 = ~x27 & ~x129 & ~x138 & ~x141 & ~x166 & ~x193 & ~x222 & ~x225 & ~x375 & ~x399 & ~x401 & ~x402 & ~x426 & ~x428 & ~x454 & ~x504 & ~x508 & ~x533 & ~x560 & ~x561 & ~x615 & ~x618 & ~x670 & ~x672 & ~x673 & ~x696 & ~x700 & ~x703 & ~x724 & ~x740 & ~x753 & ~x756 & ~x764 & ~x767 & ~x779;
assign c4154 =  x237 &  x292 & ~x75 & ~x133 & ~x187 & ~x190 & ~x225 & ~x247 & ~x278 & ~x279 & ~x333 & ~x391 & ~x405 & ~x447 & ~x561 & ~x590 & ~x730 & ~x758;
assign c4156 = ~x0 & ~x15 & ~x26 & ~x27 & ~x100 & ~x110 & ~x114 & ~x198 & ~x221 & ~x224 & ~x276 & ~x278 & ~x279 & ~x307 & ~x310 & ~x468 & ~x475 & ~x503 & ~x505 & ~x531 & ~x551 & ~x559 & ~x560 & ~x563 & ~x591 & ~x611 & ~x613 & ~x614 & ~x644 & ~x645 & ~x646 & ~x652 & ~x676 & ~x679 & ~x703 & ~x704 & ~x725 & ~x730 & ~x733 & ~x736 & ~x749 & ~x757 & ~x760 & ~x762 & ~x766 & ~x771 & ~x776 & ~x777 & ~x781;
assign c4158 =  x402 & ~x0 & ~x2 & ~x3 & ~x13 & ~x26 & ~x113 & ~x141 & ~x197 & ~x225 & ~x406 & ~x475 & ~x489 & ~x615 & ~x641 & ~x667 & ~x669 & ~x696 & ~x724 & ~x726 & ~x727 & ~x728 & ~x732 & ~x750 & ~x760;
assign c4160 = ~x0 & ~x1 & ~x4 & ~x53 & ~x54 & ~x86 & ~x112 & ~x194 & ~x327 & ~x391 & ~x459 & ~x504 & ~x554 & ~x561 & ~x606 & ~x610 & ~x615 & ~x616 & ~x618 & ~x643 & ~x669 & ~x722 & ~x747 & ~x759 & ~x762 & ~x775 & ~x782;
assign c4162 =  x347 &  x597 & ~x111 & ~x407 & ~x420 & ~x434 & ~x724 & ~x734 & ~x770 & ~x783;
assign c4164 =  x628 & ~x156 & ~x330 & ~x335 & ~x348 & ~x355 & ~x447 & ~x562 & ~x673 & ~x701;
assign c4166 = ~x32 & ~x57 & ~x138 & ~x213 & ~x240 & ~x273 & ~x274 & ~x301 & ~x302 & ~x329 & ~x363 & ~x446 & ~x475 & ~x511 & ~x512 & ~x645 & ~x701 & ~x729 & ~x770;
assign c4168 = ~x30 & ~x53 & ~x82 & ~x157 & ~x196 & ~x340 & ~x376 & ~x388 & ~x467 & ~x486 & ~x513 & ~x558 & ~x560 & ~x720 & ~x725 & ~x727 & ~x747 & ~x753;
assign c4170 =  x554 & ~x135 & ~x578 & ~x647;
assign c4172 =  x179 &  x329 & ~x47 & ~x317 & ~x370 & ~x425 & ~x699;
assign c4174 =  x0;
assign c4176 = ~x5 & ~x13 & ~x29 & ~x32 & ~x44 & ~x58 & ~x112 & ~x167 & ~x168 & ~x169 & ~x209 & ~x252 & ~x305 & ~x307 & ~x332 & ~x333 & ~x337 & ~x447 & ~x532 & ~x533 & ~x557 & ~x559 & ~x562 & ~x616 & ~x617 & ~x646 & ~x666 & ~x672 & ~x691 & ~x693 & ~x700 & ~x720 & ~x722 & ~x731 & ~x733 & ~x747 & ~x752 & ~x754 & ~x760 & ~x761 & ~x778 & ~x779;
assign c4178 =  x632 &  x715 & ~x21 & ~x184 & ~x563 & ~x579 & ~x722;
assign c4180 = ~x25 & ~x28 & ~x35 & ~x88 & ~x108 & ~x138 & ~x139 & ~x157 & ~x169 & ~x192 & ~x194 & ~x223 & ~x227 & ~x309 & ~x338 & ~x425 & ~x501 & ~x509 & ~x536 & ~x565 & ~x584 & ~x592 & ~x618 & ~x623 & ~x648 & ~x673 & ~x677 & ~x708 & ~x713 & ~x721 & ~x723 & ~x735 & ~x738 & ~x765 & ~x781;
assign c4182 =  x178 &  x605 & ~x25 & ~x52 & ~x73 & ~x74 & ~x101 & ~x102 & ~x140 & ~x251 & ~x505 & ~x586 & ~x588 & ~x696 & ~x783;
assign c4184 =  x471 &  x498 &  x679 &  x709;
assign c4186 =  x574 & ~x5 & ~x29 & ~x59 & ~x101 & ~x128 & ~x168 & ~x428 & ~x467 & ~x577 & ~x605 & ~x724;
assign c4188 = ~x50 & ~x83 & ~x110 & ~x168 & ~x185 & ~x195 & ~x308 & ~x339 & ~x348 & ~x391 & ~x404 & ~x459 & ~x502 & ~x531 & ~x643 & ~x677 & ~x735 & ~x764;
assign c4190 = ~x2 & ~x3 & ~x8 & ~x21 & ~x28 & ~x31 & ~x56 & ~x60 & ~x81 & ~x85 & ~x89 & ~x112 & ~x166 & ~x170 & ~x197 & ~x224 & ~x306 & ~x308 & ~x309 & ~x333 & ~x335 & ~x336 & ~x359 & ~x360 & ~x366 & ~x388 & ~x395 & ~x414 & ~x419 & ~x420 & ~x421 & ~x422 & ~x448 & ~x473 & ~x474 & ~x475 & ~x499 & ~x505 & ~x529 & ~x531 & ~x543 & ~x557 & ~x586 & ~x625 & ~x648 & ~x650 & ~x652 & ~x653 & ~x673 & ~x680 & ~x701 & ~x702 & ~x706 & ~x723 & ~x731 & ~x732 & ~x733 & ~x748 & ~x761 & ~x765 & ~x775 & ~x778 & ~x781;
assign c4192 =  x140;
assign c4196 =  x257 & ~x13 & ~x44 & ~x70 & ~x71 & ~x83 & ~x126 & ~x224 & ~x425 & ~x605 & ~x688 & ~x698 & ~x730 & ~x741 & ~x754 & ~x761;
assign c4198 = ~x4 & ~x6 & ~x27 & ~x30 & ~x52 & ~x53 & ~x54 & ~x83 & ~x84 & ~x86 & ~x87 & ~x111 & ~x139 & ~x140 & ~x169 & ~x223 & ~x250 & ~x253 & ~x279 & ~x283 & ~x306 & ~x336 & ~x339 & ~x358 & ~x359 & ~x360 & ~x364 & ~x365 & ~x367 & ~x391 & ~x393 & ~x414 & ~x416 & ~x420 & ~x423 & ~x433 & ~x443 & ~x444 & ~x446 & ~x447 & ~x448 & ~x469 & ~x472 & ~x474 & ~x479 & ~x504 & ~x505 & ~x506 & ~x529 & ~x533 & ~x556 & ~x557 & ~x558 & ~x559 & ~x562 & ~x584 & ~x588 & ~x597 & ~x615 & ~x618 & ~x624 & ~x640 & ~x641 & ~x642 & ~x643 & ~x651 & ~x652 & ~x669 & ~x670 & ~x673 & ~x675 & ~x677 & ~x695 & ~x698 & ~x699 & ~x703 & ~x707 & ~x722 & ~x723 & ~x725 & ~x731 & ~x749 & ~x750 & ~x751 & ~x753 & ~x754 & ~x757 & ~x760 & ~x761 & ~x763 & ~x765 & ~x777 & ~x780;
assign c4200 =  x125 & ~x30 & ~x48 & ~x75 & ~x251 & ~x252 & ~x391 & ~x393 & ~x406 & ~x420 & ~x422 & ~x433 & ~x445 & ~x446 & ~x487 & ~x541 & ~x728 & ~x757 & ~x763;
assign c4202 =  x521 &  x604 & ~x45 & ~x75 & ~x378 & ~x442 & ~x502 & ~x559;
assign c4204 =  x95 &  x152 &  x179 & ~x74 & ~x372 & ~x399 & ~x425 & ~x454 & ~x478 & ~x563;
assign c4206 =  x264 &  x526 & ~x108 & ~x189 & ~x190 & ~x274;
assign c4208 =  x365;
assign c4210 =  x124 &  x629 & ~x278 & ~x335 & ~x544 & ~x748;
assign c4212 =  x311 & ~x70 & ~x209 & ~x580 & ~x698 & ~x725;
assign c4214 = ~x1 & ~x18 & ~x25 & ~x28 & ~x30 & ~x52 & ~x53 & ~x54 & ~x56 & ~x57 & ~x81 & ~x82 & ~x85 & ~x111 & ~x112 & ~x137 & ~x138 & ~x140 & ~x164 & ~x165 & ~x166 & ~x167 & ~x168 & ~x169 & ~x187 & ~x188 & ~x189 & ~x191 & ~x194 & ~x198 & ~x214 & ~x215 & ~x216 & ~x217 & ~x220 & ~x223 & ~x225 & ~x243 & ~x244 & ~x245 & ~x250 & ~x252 & ~x273 & ~x274 & ~x275 & ~x276 & ~x277 & ~x279 & ~x301 & ~x302 & ~x303 & ~x308 & ~x330 & ~x332 & ~x359 & ~x361 & ~x362 & ~x364 & ~x418 & ~x446 & ~x474 & ~x475 & ~x503 & ~x532 & ~x577 & ~x587 & ~x700 & ~x755 & ~x756 & ~x760 & ~x773 & ~x783;
assign c4216 =  x259 &  x459 & ~x253 & ~x373 & ~x592 & ~x615;
assign c4218 =  x144 &  x680;
assign c4220 = ~x0 & ~x1 & ~x2 & ~x5 & ~x15 & ~x27 & ~x44 & ~x54 & ~x55 & ~x114 & ~x165 & ~x167 & ~x192 & ~x197 & ~x216 & ~x217 & ~x219 & ~x220 & ~x221 & ~x246 & ~x252 & ~x277 & ~x304 & ~x307 & ~x309 & ~x310 & ~x331 & ~x337 & ~x392 & ~x502 & ~x508 & ~x534 & ~x557 & ~x586 & ~x588 & ~x590 & ~x591 & ~x614 & ~x657 & ~x670 & ~x672 & ~x673 & ~x684 & ~x703 & ~x708 & ~x732 & ~x735 & ~x738 & ~x750 & ~x755 & ~x756 & ~x763 & ~x775 & ~x777 & ~x780 & ~x783;
assign c4222 =  x679 & ~x20 & ~x33 & ~x52 & ~x280 & ~x329 & ~x351 & ~x510 & ~x777;
assign c4224 =  x128 &  x182 &  x263 &  x291 &  x318 & ~x5 & ~x90 & ~x112 & ~x253 & ~x331 & ~x699 & ~x725 & ~x757;
assign c4226 =  x95 &  x96 &  x520 & ~x17 & ~x46 & ~x47 & ~x84 & ~x140 & ~x280 & ~x405 & ~x504 & ~x588 & ~x671 & ~x782;
assign c4228 =  x408 &  x547 & ~x4 & ~x52 & ~x54 & ~x161 & ~x220 & ~x221 & ~x245 & ~x268 & ~x304 & ~x503 & ~x642 & ~x697 & ~x726 & ~x755 & ~x760;
assign c4230 = ~x16 & ~x18 & ~x24 & ~x25 & ~x26 & ~x55 & ~x73 & ~x80 & ~x85 & ~x105 & ~x133 & ~x139 & ~x169 & ~x191 & ~x192 & ~x196 & ~x214 & ~x221 & ~x224 & ~x242 & ~x243 & ~x247 & ~x248 & ~x272 & ~x277 & ~x392 & ~x430 & ~x481 & ~x483 & ~x745 & ~x769;
assign c4232 =  x29;
assign c4234 = ~x1 & ~x3 & ~x30 & ~x54 & ~x55 & ~x83 & ~x84 & ~x86 & ~x110 & ~x139 & ~x152 & ~x223 & ~x237 & ~x280 & ~x298 & ~x330 & ~x353 & ~x355 & ~x357 & ~x384 & ~x385 & ~x413 & ~x440 & ~x701 & ~x702 & ~x722 & ~x728 & ~x730 & ~x751 & ~x756 & ~x757 & ~x760 & ~x761 & ~x780 & ~x782;
assign c4236 = ~x29 & ~x223 & ~x321 & ~x359 & ~x361 & ~x376 & ~x387 & ~x416 & ~x438 & ~x441 & ~x486 & ~x497 & ~x501 & ~x514 & ~x533 & ~x705 & ~x732;
assign c4238 = ~x24 & ~x25 & ~x27 & ~x29 & ~x54 & ~x57 & ~x111 & ~x139 & ~x155 & ~x167 & ~x250 & ~x304 & ~x329 & ~x331 & ~x348 & ~x357 & ~x359 & ~x361 & ~x388 & ~x390 & ~x417 & ~x551 & ~x607 & ~x662 & ~x698 & ~x718;
assign c4240 =  x401 & ~x7 & ~x56 & ~x308 & ~x322 & ~x336 & ~x349 & ~x378 & ~x517 & ~x572 & ~x600 & ~x601 & ~x628 & ~x684 & ~x697 & ~x712 & ~x734 & ~x761 & ~x762;
assign c4242 =  x200 &  x625 & ~x587 & ~x605 & ~x633 & ~x660 & ~x714 & ~x725 & ~x728 & ~x729 & ~x730 & ~x733 & ~x758 & ~x768 & ~x779;
assign c4244 =  x55;
assign c4246 =  x553 & ~x82 & ~x133 & ~x134 & ~x227 & ~x273 & ~x331 & ~x389 & ~x393 & ~x620;
assign c4248 = ~x20 & ~x21 & ~x24 & ~x28 & ~x87 & ~x113 & ~x134 & ~x195 & ~x225 & ~x266 & ~x428 & ~x506 & ~x533 & ~x615 & ~x698 & ~x700 & ~x714 & ~x729 & ~x734 & ~x742 & ~x747 & ~x757 & ~x761 & ~x762;
assign c4250 =  x560;
assign c4252 = ~x1 & ~x9 & ~x32 & ~x34 & ~x53 & ~x58 & ~x86 & ~x113 & ~x167 & ~x169 & ~x196 & ~x226 & ~x252 & ~x254 & ~x266 & ~x275 & ~x279 & ~x304 & ~x305 & ~x309 & ~x312 & ~x331 & ~x333 & ~x334 & ~x337 & ~x359 & ~x360 & ~x364 & ~x388 & ~x417 & ~x418 & ~x420 & ~x445 & ~x449 & ~x450 & ~x475 & ~x476 & ~x477 & ~x479 & ~x504 & ~x531 & ~x560 & ~x561 & ~x562 & ~x619 & ~x640 & ~x669 & ~x680 & ~x700 & ~x725 & ~x726 & ~x728 & ~x738 & ~x746 & ~x753 & ~x754 & ~x757 & ~x761 & ~x776 & ~x777 & ~x779 & ~x781;
assign c4254 = ~x6 & ~x15 & ~x16 & ~x85 & ~x138 & ~x155 & ~x167 & ~x196 & ~x237 & ~x246 & ~x250 & ~x279 & ~x305 & ~x306 & ~x336 & ~x392 & ~x532 & ~x534 & ~x562 & ~x589 & ~x647 & ~x676 & ~x731 & ~x733 & ~x748 & ~x749 & ~x754 & ~x777;
assign c4256 =  x496 & ~x0 & ~x18 & ~x19 & ~x50 & ~x75 & ~x79 & ~x80 & ~x103 & ~x104 & ~x107 & ~x133 & ~x135 & ~x166 & ~x169 & ~x195 & ~x319 & ~x345 & ~x346 & ~x372 & ~x426 & ~x427 & ~x453 & ~x477 & ~x534 & ~x561 & ~x563 & ~x588 & ~x591 & ~x617 & ~x645 & ~x647 & ~x671 & ~x674 & ~x675 & ~x755 & ~x760 & ~x781 & ~x783;
assign c4258 =  x435 &  x463 & ~x56 & ~x183 & ~x357 & ~x375 & ~x389 & ~x430 & ~x760;
assign c4260 =  x173 &  x653 & ~x12 & ~x426;
assign c4262 =  x434 & ~x26 & ~x57 & ~x70 & ~x71 & ~x99 & ~x225 & ~x252 & ~x382 & ~x410 & ~x419 & ~x531 & ~x561 & ~x562 & ~x643 & ~x702 & ~x720 & ~x731 & ~x747 & ~x758 & ~x759 & ~x761;
assign c4264 =  x376 & ~x13 & ~x14 & ~x23 & ~x57 & ~x84 & ~x87 & ~x112 & ~x224 & ~x345 & ~x397 & ~x450 & ~x451 & ~x560 & ~x561 & ~x615 & ~x645 & ~x668 & ~x670 & ~x671 & ~x702 & ~x724 & ~x733 & ~x755 & ~x762 & ~x763;
assign c4266 =  x195;
assign c4268 =  x148 &  x176 &  x597 & ~x17 & ~x53 & ~x111 & ~x169 & ~x197 & ~x308 & ~x349 & ~x670 & ~x698 & ~x725 & ~x726 & ~x750 & ~x755;
assign c4270 =  x468 & ~x5 & ~x30 & ~x76 & ~x106 & ~x363 & ~x451 & ~x505 & ~x534 & ~x535 & ~x592 & ~x614 & ~x621 & ~x707 & ~x726 & ~x729 & ~x736;
assign c4272 = ~x22 & ~x39 & ~x44 & ~x47 & ~x56 & ~x58 & ~x102 & ~x166 & ~x373 & ~x526 & ~x528 & ~x585 & ~x587 & ~x615 & ~x636 & ~x668 & ~x691 & ~x699 & ~x756 & ~x759 & ~x767 & ~x772 & ~x778;
assign c4274 = ~x0 & ~x1 & ~x2 & ~x3 & ~x17 & ~x22 & ~x23 & ~x25 & ~x47 & ~x48 & ~x50 & ~x75 & ~x78 & ~x105 & ~x106 & ~x108 & ~x109 & ~x113 & ~x114 & ~x135 & ~x138 & ~x158 & ~x162 & ~x163 & ~x167 & ~x168 & ~x169 & ~x188 & ~x191 & ~x193 & ~x197 & ~x214 & ~x216 & ~x217 & ~x224 & ~x225 & ~x226 & ~x246 & ~x247 & ~x251 & ~x274 & ~x280 & ~x308 & ~x392 & ~x504 & ~x531 & ~x532 & ~x587 & ~x615 & ~x689 & ~x702 & ~x716 & ~x728 & ~x744 & ~x757 & ~x758 & ~x759 & ~x760 & ~x768;
assign c4276 =  x319 & ~x212 & ~x245 & ~x303 & ~x330 & ~x331 & ~x358 & ~x769 & ~x770;
assign c4278 = ~x5 & ~x17 & ~x43 & ~x47 & ~x48 & ~x58 & ~x75 & ~x141 & ~x276 & ~x306 & ~x332 & ~x337 & ~x361 & ~x416 & ~x502 & ~x509 & ~x534 & ~x537 & ~x562 & ~x572 & ~x599 & ~x692 & ~x764;
assign c4280 =  x178 &  x330 & ~x142 & ~x371 & ~x372 & ~x397 & ~x452;
assign c4282 =  x602 &  x657 & ~x186 & ~x503 & ~x561 & ~x572 & ~x587 & ~x589 & ~x590 & ~x614 & ~x669 & ~x750 & ~x751;
assign c4284 =  x778;
assign c4286 =  x94 &  x683 & ~x634 & ~x715 & ~x772;
assign c4288 =  x151 &  x205 &  x632 &  x660 &  x688 & ~x420 & ~x462;
assign c4290 = ~x0 & ~x20 & ~x21 & ~x23 & ~x27 & ~x28 & ~x48 & ~x49 & ~x50 & ~x51 & ~x52 & ~x56 & ~x58 & ~x59 & ~x77 & ~x78 & ~x81 & ~x84 & ~x85 & ~x86 & ~x87 & ~x103 & ~x104 & ~x105 & ~x111 & ~x113 & ~x114 & ~x132 & ~x135 & ~x136 & ~x137 & ~x140 & ~x162 & ~x165 & ~x167 & ~x169 & ~x170 & ~x194 & ~x195 & ~x196 & ~x197 & ~x223 & ~x225 & ~x253 & ~x280 & ~x346 & ~x398 & ~x399 & ~x425 & ~x448 & ~x478 & ~x479 & ~x481 & ~x504 & ~x506 & ~x533 & ~x534 & ~x560 & ~x561 & ~x563 & ~x564 & ~x588 & ~x590 & ~x591 & ~x592 & ~x617 & ~x619 & ~x620 & ~x641 & ~x643 & ~x648 & ~x653 & ~x678 & ~x699 & ~x700 & ~x702 & ~x704 & ~x709 & ~x724 & ~x727 & ~x730 & ~x731 & ~x732 & ~x733 & ~x735 & ~x736 & ~x754 & ~x755 & ~x760 & ~x765 & ~x779;
assign c4292 =  x631 &  x658 &  x685 & ~x0 & ~x1 & ~x27 & ~x56 & ~x85 & ~x86 & ~x112 & ~x137 & ~x139 & ~x166 & ~x197 & ~x219 & ~x247 & ~x250 & ~x255 & ~x277 & ~x282 & ~x305 & ~x306 & ~x308 & ~x391 & ~x476 & ~x587 & ~x591 & ~x661 & ~x670 & ~x672 & ~x702 & ~x752 & ~x759 & ~x760 & ~x781;
assign c4294 =  x38 &  x271 & ~x74 & ~x335 & ~x336 & ~x561 & ~x590 & ~x733;
assign c4296 =  x468 &  x579 & ~x56 & ~x132 & ~x533 & ~x590 & ~x622 & ~x646 & ~x649 & ~x674;
assign c4298 =  x678 &  x737 & ~x3 & ~x50 & ~x112 & ~x138 & ~x169 & ~x218 & ~x219 & ~x770;
assign c4300 =  x289 &  x343 &  x370 & ~x3 & ~x19 & ~x21 & ~x23 & ~x30 & ~x45 & ~x46 & ~x109 & ~x111 & ~x135 & ~x136 & ~x138 & ~x161 & ~x162 & ~x164 & ~x169 & ~x171 & ~x189 & ~x193 & ~x225 & ~x281 & ~x335 & ~x364 & ~x418 & ~x419 & ~x560 & ~x616 & ~x672;
assign c4302 =  x427 & ~x247 & ~x251 & ~x274 & ~x363 & ~x388 & ~x417 & ~x475 & ~x485 & ~x503 & ~x561 & ~x589 & ~x616 & ~x673 & ~x728 & ~x729;
assign c4304 = ~x154 & ~x181 & ~x237 & ~x291 & ~x293 & ~x301 & ~x412 & ~x468 & ~x534 & ~x562 & ~x762;
assign c4306 =  x575 & ~x5 & ~x26 & ~x31 & ~x54 & ~x224 & ~x251 & ~x253 & ~x334 & ~x505 & ~x522 & ~x572 & ~x587 & ~x615 & ~x640 & ~x668 & ~x700 & ~x722 & ~x724 & ~x750 & ~x774;
assign c4308 =  x94 &  x549 & ~x16 & ~x45 & ~x211 & ~x417 & ~x527 & ~x555 & ~x582 & ~x583 & ~x610 & ~x616 & ~x638 & ~x643 & ~x694 & ~x722 & ~x735 & ~x738 & ~x748;
assign c4310 =  x494 &  x632 & ~x3 & ~x18 & ~x54 & ~x56 & ~x225 & ~x280 & ~x471 & ~x503 & ~x504 & ~x526 & ~x527 & ~x529 & ~x559 & ~x562 & ~x586 & ~x614 & ~x617 & ~x672 & ~x673 & ~x696 & ~x697 & ~x729 & ~x756 & ~x757 & ~x758 & ~x762 & ~x782 & ~x783;
assign c4312 =  x550 &  x605 &  x633 &  x660 & ~x5 & ~x19 & ~x23 & ~x167 & ~x280 & ~x563 & ~x567 & ~x592 & ~x618 & ~x647 & ~x649 & ~x673 & ~x674 & ~x700 & ~x703 & ~x731 & ~x732 & ~x758;
assign c4314 = ~x1 & ~x18 & ~x22 & ~x23 & ~x33 & ~x52 & ~x58 & ~x106 & ~x117 & ~x134 & ~x142 & ~x189 & ~x191 & ~x196 & ~x219 & ~x225 & ~x266 & ~x278 & ~x281 & ~x309 & ~x362 & ~x446 & ~x502 & ~x504 & ~x543 & ~x635 & ~x663 & ~x692 & ~x695 & ~x719 & ~x721 & ~x728 & ~x731 & ~x746 & ~x752 & ~x775 & ~x778;
assign c4316 =  x179 &  x232 & ~x57 & ~x76 & ~x131 & ~x141 & ~x279 & ~x307 & ~x344 & ~x398 & ~x425 & ~x452 & ~x478 & ~x532;
assign c4318 =  x527 & ~x51 & ~x55 & ~x113 & ~x227 & ~x302 & ~x309 & ~x418 & ~x446 & ~x672 & ~x697 & ~x698 & ~x699 & ~x700;
assign c4320 = ~x184 & ~x209 & ~x237 & ~x385 & ~x440 & ~x456 & ~x467 & ~x495 & ~x579 & ~x582 & ~x634 & ~x640 & ~x670 & ~x746 & ~x754 & ~x776;
assign c4322 =  x94 &  x574 &  x601 & ~x44 & ~x53 & ~x54 & ~x113 & ~x168 & ~x197 & ~x504 & ~x558 & ~x586 & ~x643 & ~x644 & ~x669 & ~x673 & ~x700 & ~x701 & ~x724 & ~x725 & ~x729 & ~x730 & ~x748 & ~x752 & ~x753 & ~x754 & ~x755 & ~x756 & ~x773 & ~x782;
assign c4324 =  x182 &  x292 & ~x255 & ~x281 & ~x333 & ~x433 & ~x447 & ~x621 & ~x782;
assign c4326 =  x122 &  x575 & ~x73 & ~x100 & ~x291 & ~x319 & ~x644 & ~x723 & ~x726 & ~x760;
assign c4328 =  x133 & ~x302 & ~x415 & ~x418 & ~x526 & ~x586 & ~x749;
assign c4330 =  x121 &  x176 &  x603 & ~x263 & ~x264 & ~x419 & ~x588 & ~x668 & ~x751 & ~x752;
assign c4332 =  x522 &  x577 &  x632 & ~x18 & ~x55 & ~x57 & ~x73 & ~x104 & ~x137 & ~x483 & ~x509 & ~x562 & ~x566 & ~x587 & ~x590 & ~x591 & ~x619 & ~x642 & ~x647 & ~x701 & ~x726 & ~x727 & ~x753 & ~x754;
assign c4334 = ~x2 & ~x3 & ~x15 & ~x29 & ~x30 & ~x40 & ~x56 & ~x72 & ~x110 & ~x138 & ~x280 & ~x298 & ~x301 & ~x326 & ~x327 & ~x355 & ~x357 & ~x410 & ~x411 & ~x606 & ~x633 & ~x634 & ~x662 & ~x701 & ~x702 & ~x717 & ~x718 & ~x745 & ~x748 & ~x758 & ~x761;
assign c4336 =  x652 & ~x301 & ~x356 & ~x410 & ~x521 & ~x662;
assign c4338 =  x399 &  x598 &  x653 & ~x224 & ~x484 & ~x540;
assign c4340 =  x526 & ~x162 & ~x223 & ~x274 & ~x308 & ~x448 & ~x509 & ~x729 & ~x762;
assign c4342 =  x365 & ~x156 & ~x580;
assign c4344 =  x161 & ~x183 & ~x237 & ~x388 & ~x415 & ~x444 & ~x583 & ~x585 & ~x722 & ~x760;
assign c4346 =  x634 &  x690 & ~x364 & ~x378 & ~x405 & ~x488 & ~x515 & ~x615;
assign c4348 =  x499 & ~x19 & ~x134 & ~x138 & ~x165 & ~x197 & ~x252 & ~x479 & ~x484 & ~x757;
assign c4350 =  x64 &  x67 & ~x18 & ~x44 & ~x45 & ~x56 & ~x83 & ~x84 & ~x85 & ~x100 & ~x115 & ~x673;
assign c4352 =  x493 &  x632 & ~x1 & ~x351 & ~x461 & ~x563 & ~x727;
assign c4354 = ~x25 & ~x195 & ~x196 & ~x224 & ~x266 & ~x321 & ~x338 & ~x349 & ~x364 & ~x365 & ~x366 & ~x450 & ~x460 & ~x587 & ~x589 & ~x651 & ~x668 & ~x695 & ~x700 & ~x705 & ~x706 & ~x708 & ~x728 & ~x731 & ~x736 & ~x750 & ~x777 & ~x778;
assign c4356 =  x56;
assign c4358 = ~x18 & ~x90 & ~x93 & ~x115 & ~x137 & ~x159 & ~x282 & ~x304 & ~x311 & ~x336 & ~x455 & ~x554 & ~x559 & ~x586 & ~x646 & ~x696 & ~x748 & ~x769 & ~x776;
assign c4360 =  x463 & ~x209 & ~x264 & ~x335 & ~x529 & ~x613 & ~x705;
assign c4362 =  x575 &  x658 & ~x14 & ~x29 & ~x43 & ~x55 & ~x139 & ~x475 & ~x529 & ~x560 & ~x579 & ~x588 & ~x617 & ~x637 & ~x691 & ~x701 & ~x721 & ~x776;
assign c4364 =  x150 & ~x31 & ~x55 & ~x278 & ~x294 & ~x305 & ~x307 & ~x333 & ~x349 & ~x362 & ~x390 & ~x446 & ~x449 & ~x450 & ~x477 & ~x503 & ~x504 & ~x529 & ~x595 & ~x640 & ~x650 & ~x668 & ~x669 & ~x680 & ~x706 & ~x723 & ~x727 & ~x732 & ~x733 & ~x735 & ~x754 & ~x760 & ~x763 & ~x779;
assign c4366 =  x102 &  x681;
assign c4368 =  x520 &  x548 &  x603 & ~x20 & ~x25 & ~x43 & ~x44 & ~x45 & ~x82 & ~x85 & ~x102 & ~x196 & ~x224 & ~x479 & ~x504 & ~x505 & ~x532 & ~x563 & ~x702 & ~x721 & ~x723 & ~x724 & ~x748 & ~x759;
assign c4370 =  x346 & ~x0 & ~x3 & ~x6 & ~x29 & ~x32 & ~x55 & ~x56 & ~x81 & ~x84 & ~x86 & ~x140 & ~x166 & ~x169 & ~x198 & ~x280 & ~x281 & ~x308 & ~x309 & ~x433 & ~x461 & ~x516 & ~x544 & ~x670 & ~x671 & ~x706 & ~x752 & ~x753 & ~x763 & ~x764 & ~x779;
assign c4372 =  x315 &  x343 & ~x101 & ~x183 & ~x308 & ~x430 & ~x431 & ~x486 & ~x533 & ~x755 & ~x757;
assign c4374 =  x371 & ~x6 & ~x19 & ~x28 & ~x29 & ~x32 & ~x55 & ~x56 & ~x110 & ~x167 & ~x223 & ~x251 & ~x253 & ~x279 & ~x281 & ~x302 & ~x304 & ~x305 & ~x334 & ~x484 & ~x511 & ~x532 & ~x537 & ~x560 & ~x565 & ~x751;
assign c4376 =  x175 & ~x2 & ~x21 & ~x25 & ~x28 & ~x42 & ~x43 & ~x44 & ~x54 & ~x57 & ~x58 & ~x70 & ~x71 & ~x73 & ~x85 & ~x99 & ~x136 & ~x137 & ~x164 & ~x195 & ~x223 & ~x224 & ~x252 & ~x336 & ~x447 & ~x502 & ~x503 & ~x532 & ~x671 & ~x700 & ~x731 & ~x733 & ~x734 & ~x735 & ~x758 & ~x760 & ~x769 & ~x782;
assign c4378 =  x571 &  x598 & ~x2 & ~x30 & ~x59 & ~x83 & ~x85 & ~x142 & ~x196 & ~x222 & ~x225 & ~x249 & ~x506 & ~x614 & ~x699 & ~x715 & ~x726 & ~x742;
assign c4380 =  x495 &  x606 &  x661 & ~x130 & ~x158 & ~x563;
assign c4382 =  x226 &  x650;
assign c4384 = ~x0 & ~x4 & ~x18 & ~x22 & ~x81 & ~x131 & ~x139 & ~x162 & ~x165 & ~x278 & ~x279 & ~x283 & ~x309 & ~x336 & ~x361 & ~x389 & ~x416 & ~x444 & ~x472 & ~x474 & ~x531 & ~x585 & ~x587 & ~x621 & ~x628 & ~x644 & ~x655 & ~x681 & ~x703 & ~x708 & ~x718 & ~x729 & ~x730 & ~x740 & ~x780;
assign c4386 =  x386 & ~x77 & ~x170 & ~x196 & ~x317 & ~x343 & ~x370 & ~x371 & ~x397 & ~x452 & ~x476 & ~x504 & ~x561 & ~x590 & ~x618 & ~x673 & ~x674;
assign c4388 =  x373 & ~x0 & ~x1 & ~x7 & ~x57 & ~x86 & ~x112 & ~x360 & ~x361 & ~x362 & ~x363 & ~x391 & ~x404 & ~x415 & ~x416 & ~x443 & ~x444 & ~x459 & ~x469 & ~x473 & ~x528 & ~x533 & ~x697 & ~x721 & ~x727 & ~x728 & ~x751 & ~x760 & ~x762 & ~x763 & ~x779;
assign c4390 =  x394 & ~x13;
assign c4392 =  x180 &  x236 & ~x51 & ~x81 & ~x165 & ~x279 & ~x350 & ~x377 & ~x432 & ~x476 & ~x729 & ~x757;
assign c4394 =  x175 & ~x11 & ~x83 & ~x84 & ~x182 & ~x209 & ~x419 & ~x469 & ~x553 & ~x555 & ~x561 & ~x581 & ~x615 & ~x616 & ~x666;
assign c4396 = ~x27 & ~x64 & ~x110 & ~x119 & ~x143 & ~x144 & ~x164 & ~x198 & ~x227 & ~x309 & ~x328 & ~x331 & ~x337 & ~x446 & ~x448 & ~x499 & ~x614 & ~x635 & ~x643 & ~x653 & ~x732 & ~x750 & ~x767 & ~x778;
assign c4398 =  x662 & ~x351 & ~x434 & ~x447 & ~x461 & ~x476 & ~x488 & ~x558 & ~x615 & ~x707 & ~x735 & ~x781;
assign c4400 =  x548 &  x632 & ~x18 & ~x462 & ~x489 & ~x587 & ~x615 & ~x673;
assign c4402 =  x651 &  x658 &  x737;
assign c4404 =  x174 &  x651 & ~x486 & ~x662;
assign c4406 = ~x0 & ~x4 & ~x20 & ~x21 & ~x25 & ~x27 & ~x28 & ~x45 & ~x47 & ~x48 & ~x52 & ~x55 & ~x75 & ~x82 & ~x85 & ~x105 & ~x106 & ~x107 & ~x109 & ~x113 & ~x133 & ~x134 & ~x141 & ~x160 & ~x162 & ~x165 & ~x167 & ~x187 & ~x188 & ~x190 & ~x192 & ~x195 & ~x197 & ~x219 & ~x221 & ~x244 & ~x248 & ~x272 & ~x274 & ~x277 & ~x299 & ~x300 & ~x302 & ~x308 & ~x309 & ~x330 & ~x336 & ~x362 & ~x388 & ~x504 & ~x587 & ~x588 & ~x615 & ~x643 & ~x672 & ~x691 & ~x700 & ~x701 & ~x719 & ~x729 & ~x742 & ~x746 & ~x756 & ~x759 & ~x769;
assign c4408 =  x180 &  x182 & ~x5 & ~x6 & ~x19 & ~x20 & ~x31 & ~x84 & ~x109 & ~x113 & ~x133 & ~x139 & ~x142 & ~x162 & ~x167 & ~x168 & ~x170 & ~x197 & ~x200 & ~x225 & ~x228 & ~x281 & ~x282 & ~x306 & ~x307 & ~x322 & ~x333 & ~x391 & ~x419 & ~x421 & ~x446 & ~x447 & ~x502 & ~x503 & ~x617 & ~x618 & ~x726 & ~x730 & ~x780;
assign c4410 = ~x22 & ~x46 & ~x81 & ~x162 & ~x163 & ~x168 & ~x169 & ~x251 & ~x252 & ~x278 & ~x307 & ~x402 & ~x429 & ~x457 & ~x484 & ~x579 & ~x607 & ~x615 & ~x636 & ~x670 & ~x689 & ~x691 & ~x716 & ~x744 & ~x745 & ~x758;
assign c4412 =  x365 & ~x97 & ~x184 & ~x252 & ~x615 & ~x670 & ~x781;
assign c4414 =  x383 &  x633 & ~x609;
assign c4416 =  x492 &  x548 &  x631 & ~x27 & ~x84 & ~x168 & ~x185 & ~x448 & ~x591 & ~x733 & ~x775;
assign c4418 = ~x56 & ~x115 & ~x279 & ~x294 & ~x337 & ~x385 & ~x432 & ~x471 & ~x487 & ~x504 & ~x542 & ~x612 & ~x615 & ~x638 & ~x639 & ~x667 & ~x701 & ~x724 & ~x753 & ~x755 & ~x762 & ~x778;
assign c4420 =  x201 &  x228 & ~x82 & ~x169 & ~x183 & ~x196 & ~x441 & ~x525 & ~x641 & ~x670;
assign c4422 =  x92 &  x119 &  x709 & ~x183 & ~x197;
assign c4424 =  x546 &  x573 & ~x14 & ~x19 & ~x22 & ~x29 & ~x30 & ~x43 & ~x45 & ~x46 & ~x52 & ~x53 & ~x57 & ~x141 & ~x168 & ~x195 & ~x196 & ~x197 & ~x225 & ~x448 & ~x478 & ~x501 & ~x506 & ~x507 & ~x530 & ~x560 & ~x585 & ~x586 & ~x589 & ~x590 & ~x612 & ~x613 & ~x641 & ~x644 & ~x646 & ~x665 & ~x668 & ~x675 & ~x692 & ~x697 & ~x700 & ~x721 & ~x727 & ~x728 & ~x732 & ~x733 & ~x746 & ~x747 & ~x748 & ~x749 & ~x751 & ~x775;
assign c4426 =  x371 & ~x56 & ~x280 & ~x357 & ~x360 & ~x362 & ~x384 & ~x386 & ~x388 & ~x412 & ~x458 & ~x474 & ~x485 & ~x501 & ~x530 & ~x587 & ~x589 & ~x645 & ~x702 & ~x704 & ~x730 & ~x777;
assign c4428 =  x93 &  x603 & ~x72 & ~x210 & ~x236 & ~x319 & ~x347 & ~x616 & ~x645 & ~x698 & ~x727 & ~x750 & ~x753 & ~x760;
assign c4430 = ~x1 & ~x20 & ~x26 & ~x28 & ~x29 & ~x56 & ~x57 & ~x60 & ~x84 & ~x104 & ~x110 & ~x114 & ~x139 & ~x141 & ~x142 & ~x158 & ~x162 & ~x164 & ~x167 & ~x191 & ~x220 & ~x251 & ~x279 & ~x281 & ~x373 & ~x400 & ~x424 & ~x427 & ~x455 & ~x477 & ~x480 & ~x534 & ~x536 & ~x563 & ~x564 & ~x588 & ~x619 & ~x645 & ~x667 & ~x670 & ~x675 & ~x679 & ~x683 & ~x709 & ~x712 & ~x723 & ~x725 & ~x728 & ~x730 & ~x734 & ~x737 & ~x739 & ~x753 & ~x775;
assign c4432 =  x547 &  x575 & ~x2 & ~x21 & ~x193 & ~x273 & ~x304 & ~x361 & ~x419 & ~x422 & ~x449 & ~x537 & ~x561 & ~x578 & ~x633 & ~x773 & ~x775;
assign c4434 =  x229 &  x257 &  x283 & ~x57 & ~x368 & ~x369 & ~x448 & ~x669;
assign c4436 = ~x37 & ~x110 & ~x160 & ~x167 & ~x170 & ~x195 & ~x391 & ~x422 & ~x423 & ~x530 & ~x562 & ~x602 & ~x629 & ~x667 & ~x684 & ~x697 & ~x739 & ~x750 & ~x754 & ~x764;
assign c4438 =  x629 & ~x23 & ~x57 & ~x195 & ~x328 & ~x356 & ~x385 & ~x441 & ~x459 & ~x471 & ~x487 & ~x543 & ~x569 & ~x750;
assign c4440 =  x206 &  x234 &  x262 & ~x15 & ~x21 & ~x25 & ~x27 & ~x84 & ~x86 & ~x169 & ~x278 & ~x279 & ~x301 & ~x306 & ~x307 & ~x308 & ~x332 & ~x333 & ~x361 & ~x389 & ~x417 & ~x419 & ~x446 & ~x588 & ~x645 & ~x674 & ~x680 & ~x730 & ~x736 & ~x748 & ~x749 & ~x757 & ~x762 & ~x763;
assign c4442 =  x152 &  x382 & ~x55 & ~x371 & ~x425 & ~x531 & ~x621;
assign c4444 = ~x1 & ~x4 & ~x52 & ~x59 & ~x83 & ~x195 & ~x223 & ~x311 & ~x321 & ~x339 & ~x359 & ~x392 & ~x419 & ~x423 & ~x446 & ~x474 & ~x495 & ~x531 & ~x533 & ~x577 & ~x605 & ~x614 & ~x642 & ~x645 & ~x670 & ~x671 & ~x672 & ~x733 & ~x746 & ~x747 & ~x749 & ~x752 & ~x764 & ~x781;
assign c4446 =  x491 &  x603 &  x684 & ~x24 & ~x335 & ~x562 & ~x722 & ~x777;
assign c4448 =  x120 &  x653 &  x681 & ~x43 & ~x70 & ~x169 & ~x196 & ~x197 & ~x198 & ~x224 & ~x225 & ~x691 & ~x756 & ~x773;
assign c4450 =  x519 &  x546 & ~x56 & ~x58 & ~x84 & ~x114 & ~x165 & ~x242 & ~x247 & ~x302 & ~x307 & ~x362 & ~x392 & ~x418 & ~x421 & ~x450 & ~x474 & ~x529 & ~x587 & ~x588 & ~x616 & ~x672 & ~x674 & ~x721 & ~x745 & ~x746 & ~x773 & ~x781;
assign c4452 =  x67 &  x96 &  x549 & ~x462;
assign c4454 =  x65 &  x521 & ~x533 & ~x646;
assign c4456 = ~x2 & ~x23 & ~x28 & ~x42 & ~x58 & ~x99 & ~x111 & ~x112 & ~x139 & ~x154 & ~x208 & ~x211 & ~x252 & ~x301 & ~x327 & ~x329 & ~x355 & ~x357 & ~x383 & ~x385 & ~x411 & ~x498 & ~x555 & ~x587 & ~x763 & ~x779 & ~x780;
assign c4458 =  x29;
assign c4460 =  x679;
assign c4462 =  x94 &  x441 & ~x12 & ~x200 & ~x464 & ~x645;
assign c4464 =  x610 & ~x0 & ~x29 & ~x108 & ~x135 & ~x165 & ~x222 & ~x393 & ~x394 & ~x477 & ~x537 & ~x562;
assign c4466 =  x610 &  x626 & ~x194 & ~x198 & ~x280 & ~x323 & ~x531 & ~x723;
assign c4468 =  x497 &  x552 &  x579 &  x634 & ~x48 & ~x114 & ~x426 & ~x533 & ~x535 & ~x644 & ~x675;
assign c4470 = ~x24 & ~x25 & ~x40 & ~x69 & ~x71 & ~x80 & ~x82 & ~x109 & ~x252 & ~x412 & ~x548 & ~x559 & ~x604 & ~x632 & ~x633 & ~x688 & ~x715 & ~x751 & ~x756 & ~x758 & ~x769 & ~x778;
assign c4472 =  x439 &  x608 &  x663 & ~x132 & ~x477 & ~x674;
assign c4474 =  x688 & ~x4 & ~x112 & ~x225 & ~x350 & ~x420 & ~x422 & ~x515 & ~x650 & ~x671 & ~x673 & ~x757 & ~x763;
assign c4476 =  x628 & ~x154 & ~x466 & ~x522 & ~x548;
assign c4478 = ~x0 & ~x17 & ~x19 & ~x58 & ~x73 & ~x87 & ~x114 & ~x136 & ~x192 & ~x193 & ~x195 & ~x252 & ~x276 & ~x279 & ~x280 & ~x306 & ~x310 & ~x394 & ~x418 & ~x421 & ~x449 & ~x505 & ~x557 & ~x613 & ~x615 & ~x633 & ~x643 & ~x660 & ~x671 & ~x704 & ~x715 & ~x726 & ~x733 & ~x742;
assign c4480 =  x91 & ~x71 & ~x101 & ~x113 & ~x127 & ~x142 & ~x221 & ~x400 & ~x506 & ~x754 & ~x767;
assign c4482 =  x182 &  x208 &  x497 & ~x145;
assign c4484 =  x123 & ~x16 & ~x18 & ~x86 & ~x306 & ~x312 & ~x335 & ~x535 & ~x541 & ~x564 & ~x746 & ~x766;
assign c4486 =  x400 & ~x279 & ~x363 & ~x403 & ~x413 & ~x431 & ~x475 & ~x479 & ~x497 & ~x500 & ~x530 & ~x555 & ~x557 & ~x558 & ~x587 & ~x727 & ~x763 & ~x764 & ~x765;
assign c4488 =  x602 &  x629 &  x656 &  x683 & ~x0 & ~x44 & ~x74 & ~x102 & ~x308 & ~x418 & ~x446 & ~x503 & ~x504 & ~x533 & ~x618 & ~x756 & ~x783;
assign c4490 =  x263 &  x315 &  x316 &  x317 & ~x26 & ~x169 & ~x196 & ~x228 & ~x275 & ~x307 & ~x309 & ~x336 & ~x503 & ~x534 & ~x562 & ~x589 & ~x645 & ~x646;
assign c4492 =  x484 & ~x84 & ~x167 & ~x252 & ~x359 & ~x390 & ~x391 & ~x418 & ~x441 & ~x444 & ~x460 & ~x475 & ~x488 & ~x502 & ~x503 & ~x528 & ~x703 & ~x731 & ~x750 & ~x760 & ~x777;
assign c4494 =  x630 & ~x2 & ~x25 & ~x27 & ~x83 & ~x168 & ~x184 & ~x377 & ~x391 & ~x416 & ~x459 & ~x561 & ~x589 & ~x673 & ~x730 & ~x731 & ~x751 & ~x761 & ~x762;
assign c4496 =  x523 &  x551 &  x606 &  x661 & ~x23 & ~x24 & ~x47 & ~x168 & ~x224 & ~x452 & ~x533 & ~x679 & ~x699 & ~x727 & ~x757 & ~x783;
assign c4498 =  x92 &  x93 & ~x12 & ~x13 & ~x14 & ~x15 & ~x16 & ~x18 & ~x42 & ~x44 & ~x55 & ~x141 & ~x168 & ~x461 & ~x474 & ~x475 & ~x479 & ~x504 & ~x505 & ~x557 & ~x558 & ~x559 & ~x560 & ~x614 & ~x616 & ~x617 & ~x642 & ~x645 & ~x670 & ~x671;
assign c41 = ~x51 & ~x105 & ~x145 & ~x179 & ~x292 & ~x365 & ~x448 & ~x473;
assign c43 =  x397 &  x426 &  x453 & ~x66 & ~x106 & ~x697 & ~x727 & ~x755;
assign c45 = ~x292 & ~x294 & ~x319 & ~x347 & ~x350 & ~x351 & ~x375 & ~x376 & ~x379 & ~x420 & ~x448 & ~x449 & ~x749 & ~x755 & ~x756 & ~x772;
assign c47 = ~x0 & ~x1 & ~x33 & ~x41 & ~x94 & ~x149 & ~x150 & ~x651 & ~x678 & ~x707 & ~x770 & ~x771;
assign c49 =  x663 & ~x1 & ~x49 & ~x50 & ~x53 & ~x78 & ~x79 & ~x80 & ~x106 & ~x133 & ~x393 & ~x417 & ~x447 & ~x448 & ~x472 & ~x475 & ~x476 & ~x497 & ~x499 & ~x524 & ~x526 & ~x528 & ~x553 & ~x782;
assign c411 =  x211 &  x267 & ~x0 & ~x4 & ~x26 & ~x27 & ~x53 & ~x79 & ~x80 & ~x82 & ~x112 & ~x139 & ~x140 & ~x141 & ~x168 & ~x427 & ~x428 & ~x457 & ~x559 & ~x587 & ~x643 & ~x669 & ~x670 & ~x671 & ~x700 & ~x756;
assign c413 =  x326 &  x353 &  x378 & ~x0 & ~x359 & ~x471 & ~x499;
assign c415 =  x194 & ~x680;
assign c417 = ~x55 & ~x222 & ~x223 & ~x226 & ~x249 & ~x305 & ~x314 & ~x390 & ~x415 & ~x490 & ~x658 & ~x688;
assign c419 =  x731 & ~x681 & ~x709;
assign c421 =  x388 & ~x356 & ~x357 & ~x557 & ~x559 & ~x586 & ~x639 & ~x641 & ~x671 & ~x703 & ~x757 & ~x783;
assign c423 =  x350 & ~x24 & ~x110 & ~x314 & ~x390 & ~x392 & ~x411 & ~x427 & ~x475 & ~x498 & ~x508 & ~x525 & ~x618 & ~x704;
assign c425 =  x324 &  x352 & ~x53 & ~x77 & ~x369 & ~x390 & ~x392 & ~x398 & ~x414 & ~x415 & ~x417 & ~x441 & ~x455 & ~x468 & ~x470 & ~x528 & ~x533 & ~x555 & ~x583 & ~x591 & ~x675 & ~x755;
assign c427 = ~x2 & ~x26 & ~x32 & ~x52 & ~x59 & ~x372 & ~x402 & ~x458 & ~x459 & ~x488 & ~x489 & ~x569 & ~x617 & ~x646;
assign c429 =  x249 & ~x467 & ~x539 & ~x566 & ~x624;
assign c431 =  x745 & ~x528 & ~x662 & ~x663;
assign c433 =  x160 & ~x26 & ~x56 & ~x84 & ~x109 & ~x167 & ~x560 & ~x599;
assign c435 =  x269 &  x324 &  x352 & ~x23 & ~x50 & ~x198 & ~x257 & ~x284 & ~x340 & ~x507 & ~x754 & ~x755;
assign c437 = ~x9 & ~x10 & ~x19 & ~x22 & ~x27 & ~x598 & ~x599 & ~x626 & ~x649 & ~x652 & ~x653 & ~x654 & ~x668 & ~x707 & ~x708 & ~x724 & ~x726 & ~x734 & ~x744 & ~x745 & ~x746 & ~x747 & ~x752 & ~x770 & ~x774 & ~x775 & ~x776;
assign c439 =  x103 & ~x0 & ~x25 & ~x625 & ~x680;
assign c441 =  x265 &  x516 & ~x1 & ~x23 & ~x27 & ~x134 & ~x199 & ~x249 & ~x308 & ~x734 & ~x779;
assign c443 = ~x0 & ~x2 & ~x17 & ~x21 & ~x30 & ~x31 & ~x46 & ~x53 & ~x56 & ~x77 & ~x78 & ~x79 & ~x81 & ~x83 & ~x104 & ~x106 & ~x108 & ~x137 & ~x159 & ~x160 & ~x161 & ~x191 & ~x214 & ~x215 & ~x216 & ~x242 & ~x252 & ~x269 & ~x270 & ~x271 & ~x297 & ~x335 & ~x338 & ~x339 & ~x366 & ~x394 & ~x420 & ~x421 & ~x445 & ~x448 & ~x452 & ~x453 & ~x472 & ~x477 & ~x478 & ~x479 & ~x497 & ~x500 & ~x502 & ~x505 & ~x528 & ~x532 & ~x533 & ~x552 & ~x554 & ~x557 & ~x563 & ~x583 & ~x586 & ~x588 & ~x589 & ~x591 & ~x616 & ~x640 & ~x641 & ~x646 & ~x648 & ~x671 & ~x696 & ~x699 & ~x700 & ~x727 & ~x728 & ~x731 & ~x752 & ~x755 & ~x760 & ~x782 & ~x783;
assign c445 =  x241 & ~x0 & ~x23 & ~x38 & ~x65 & ~x82 & ~x84 & ~x93 & ~x140 & ~x175 & ~x756 & ~x759 & ~x775;
assign c447 =  x714 &  x715 & ~x160 & ~x611 & ~x632 & ~x634 & ~x636;
assign c449 = ~x54 & ~x87 & ~x88 & ~x244 & ~x273 & ~x298 & ~x300 & ~x380 & ~x584 & ~x585 & ~x589 & ~x591 & ~x611 & ~x637 & ~x651 & ~x676 & ~x679 & ~x708 & ~x727 & ~x728 & ~x730 & ~x733 & ~x781;
assign c451 = ~x26 & ~x106 & ~x107 & ~x213 & ~x240 & ~x308 & ~x336 & ~x444 & ~x447 & ~x449 & ~x474 & ~x497 & ~x498 & ~x501 & ~x522 & ~x524 & ~x526 & ~x531 & ~x536 & ~x551 & ~x552 & ~x554 & ~x558 & ~x560 & ~x563 & ~x593 & ~x640 & ~x642 & ~x646 & ~x648 & ~x697 & ~x698 & ~x699 & ~x700 & ~x702 & ~x727 & ~x728 & ~x729 & ~x732 & ~x753 & ~x759 & ~x763 & ~x781;
assign c453 =  x267 & ~x337 & ~x627 & ~x658 & ~x780;
assign c455 = ~x5 & ~x23 & ~x27 & ~x55 & ~x139 & ~x300 & ~x325 & ~x328 & ~x329 & ~x566 & ~x594 & ~x597 & ~x622 & ~x623 & ~x624 & ~x653 & ~x665 & ~x667 & ~x668 & ~x682 & ~x698 & ~x723 & ~x782;
assign c457 =  x459 & ~x541 & ~x550 & ~x552 & ~x597 & ~x648;
assign c459 = ~x25 & ~x50 & ~x53 & ~x77 & ~x79 & ~x106 & ~x112 & ~x130 & ~x184 & ~x186 & ~x187 & ~x240 & ~x241 & ~x268 & ~x365 & ~x394 & ~x395 & ~x421 & ~x448 & ~x471 & ~x472 & ~x476 & ~x496 & ~x497 & ~x498 & ~x499 & ~x501 & ~x505 & ~x506 & ~x507 & ~x525 & ~x528 & ~x531 & ~x555 & ~x556 & ~x557 & ~x558 & ~x559 & ~x585 & ~x586 & ~x588 & ~x617 & ~x698 & ~x699 & ~x731;
assign c461 =  x324 & ~x22 & ~x57 & ~x195 & ~x287 & ~x303 & ~x336 & ~x370 & ~x414 & ~x429;
assign c463 = ~x24 & ~x35 & ~x458 & ~x476 & ~x482 & ~x516 & ~x561 & ~x590 & ~x591 & ~x595 & ~x596 & ~x617 & ~x618 & ~x670 & ~x752 & ~x773 & ~x776 & ~x783;
assign c465 = ~x2 & ~x21 & ~x22 & ~x25 & ~x42 & ~x51 & ~x52 & ~x69 & ~x122 & ~x337 & ~x365 & ~x366 & ~x420 & ~x560 & ~x613 & ~x615 & ~x641 & ~x671 & ~x753 & ~x760 & ~x765;
assign c467 =  x740 & ~x132 & ~x658 & ~x760;
assign c469 =  x446 & ~x668 & ~x681 & ~x706 & ~x722 & ~x776;
assign c471 =  x457 &  x487 & ~x78 & ~x161 & ~x553;
assign c473 =  x717 & ~x524 & ~x527 & ~x549 & ~x551 & ~x580;
assign c475 = ~x20 & ~x21 & ~x29 & ~x39 & ~x42 & ~x79 & ~x88 & ~x106 & ~x615 & ~x625 & ~x643 & ~x678 & ~x697 & ~x704 & ~x719 & ~x750 & ~x752 & ~x755 & ~x768 & ~x770 & ~x771 & ~x782;
assign c477 =  x405 &  x428 &  x459;
assign c479 =  x342 &  x427 & ~x262 & ~x392 & ~x449;
assign c481 = ~x0 & ~x3 & ~x29 & ~x30 & ~x55 & ~x59 & ~x60 & ~x82 & ~x112 & ~x134 & ~x147 & ~x168 & ~x174 & ~x196 & ~x202 & ~x208 & ~x672 & ~x700 & ~x755 & ~x756 & ~x773 & ~x777;
assign c483 = ~x37 & ~x55 & ~x79 & ~x126 & ~x154 & ~x337 & ~x363 & ~x364 & ~x393 & ~x445 & ~x447 & ~x449 & ~x456 & ~x472 & ~x501 & ~x528 & ~x560 & ~x618 & ~x671 & ~x697 & ~x698 & ~x728 & ~x754 & ~x782;
assign c485 = ~x0 & ~x52 & ~x54 & ~x350 & ~x433 & ~x434 & ~x436 & ~x464 & ~x477 & ~x504 & ~x560 & ~x644 & ~x715 & ~x717 & ~x729;
assign c487 =  x140;
assign c489 =  x130 &  x131 & ~x2 & ~x24 & ~x25 & ~x28 & ~x85 & ~x196 & ~x625;
assign c491 = ~x1 & ~x25 & ~x27 & ~x28 & ~x83 & ~x113 & ~x114 & ~x141 & ~x166 & ~x281 & ~x477 & ~x493 & ~x571 & ~x598 & ~x599 & ~x600 & ~x627 & ~x654 & ~x714 & ~x756 & ~x782 & ~x783;
assign c493 = ~x125 & ~x127 & ~x347 & ~x380 & ~x406 & ~x421 & ~x743 & ~x744 & ~x759 & ~x774 & ~x778;
assign c495 = ~x461 & ~x489 & ~x490 & ~x518 & ~x519 & ~x520 & ~x588 & ~x590 & ~x643 & ~x645 & ~x698 & ~x703 & ~x724 & ~x746 & ~x757 & ~x776 & ~x780;
assign c497 =  x723 & ~x62 & ~x419;
assign c499 = ~x205 & ~x206 & ~x232 & ~x316 & ~x322 & ~x362 & ~x371 & ~x389 & ~x390 & ~x417 & ~x475;
assign c4101 =  x743 &  x745 & ~x633 & ~x634;
assign c4103 =  x343 &  x456 & ~x55 & ~x421 & ~x583 & ~x584 & ~x640 & ~x699 & ~x717 & ~x772;
assign c4105 =  x425 & ~x7 & ~x9 & ~x26 & ~x27 & ~x57 & ~x114 & ~x115 & ~x168 & ~x617 & ~x645 & ~x646 & ~x673 & ~x681 & ~x701 & ~x754 & ~x764 & ~x783;
assign c4107 =  x210 & ~x30 & ~x551 & ~x567 & ~x584 & ~x586 & ~x609 & ~x728 & ~x755;
assign c4109 =  x315 &  x428 & ~x10 & ~x21 & ~x74 & ~x77 & ~x111 & ~x128 & ~x449;
assign c4111 =  x745 & ~x364 & ~x549 & ~x551 & ~x552 & ~x578 & ~x579 & ~x580 & ~x609 & ~x672;
assign c4113 = ~x124 & ~x180 & ~x319 & ~x348 & ~x393 & ~x421 & ~x738 & ~x744 & ~x757 & ~x777;
assign c4115 =  x488 & ~x5 & ~x50 & ~x196 & ~x414 & ~x437 & ~x440 & ~x442 & ~x450 & ~x505 & ~x643 & ~x679 & ~x763;
assign c4117 =  x239 &  x295 &  x380 & ~x28 & ~x62 & ~x86 & ~x281;
assign c4119 =  x717 & ~x524 & ~x549 & ~x555;
assign c4121 =  x371 &  x418 & ~x21 & ~x48 & ~x51 & ~x75 & ~x77 & ~x103 & ~x705;
assign c4123 =  x430 &  x459 &  x488 & ~x79 & ~x106 & ~x109 & ~x448 & ~x643 & ~x703 & ~x705;
assign c4125 =  x457 &  x486 &  x487 &  x516 & ~x0 & ~x28 & ~x84 & ~x110 & ~x111 & ~x764;
assign c4127 =  x287 &  x370 & ~x12 & ~x39 & ~x50 & ~x54 & ~x122;
assign c4129 = ~x30 & ~x322 & ~x375 & ~x377 & ~x406 & ~x449 & ~x476 & ~x576 & ~x605 & ~x696 & ~x737 & ~x752;
assign c4131 = ~x0 & ~x26 & ~x54 & ~x84 & ~x136 & ~x139 & ~x220 & ~x254 & ~x255 & ~x257 & ~x281 & ~x284 & ~x304 & ~x305 & ~x309 & ~x311 & ~x336 & ~x338 & ~x339 & ~x343 & ~x361 & ~x362 & ~x365 & ~x368 & ~x369 & ~x370 & ~x389 & ~x394 & ~x395 & ~x400 & ~x412 & ~x413 & ~x416 & ~x417 & ~x419 & ~x424 & ~x425 & ~x427 & ~x428 & ~x442 & ~x458 & ~x480 & ~x500 & ~x501 & ~x503 & ~x508 & ~x531 & ~x556 & ~x560 & ~x582 & ~x584 & ~x588 & ~x591 & ~x613 & ~x617 & ~x643 & ~x673 & ~x696 & ~x697 & ~x702 & ~x725 & ~x727 & ~x729 & ~x730 & ~x732 & ~x752 & ~x755 & ~x760;
assign c4133 = ~x418 & ~x449 & ~x478 & ~x530 & ~x532 & ~x573 & ~x574 & ~x575 & ~x603 & ~x606 & ~x617 & ~x632 & ~x644 & ~x645 & ~x727 & ~x728;
assign c4135 =  x183 &  x239 &  x379 & ~x106 & ~x754 & ~x777 & ~x782;
assign c4137 =  x744 & ~x27 & ~x162 & ~x227 & ~x310 & ~x476 & ~x586 & ~x588 & ~x634 & ~x635 & ~x637;
assign c4139 =  x301 & ~x94 & ~x334 & ~x360 & ~x389 & ~x773;
assign c4141 =  x296 & ~x30 & ~x51 & ~x66 & ~x224 & ~x334 & ~x556 & ~x560 & ~x586 & ~x617 & ~x698 & ~x747;
assign c4143 = ~x26 & ~x252 & ~x305 & ~x371 & ~x463 & ~x615 & ~x672;
assign c4145 =  x480 &  x508 & ~x10 & ~x19 & ~x38 & ~x74 & ~x365 & ~x641 & ~x775 & ~x777 & ~x780;
assign c4147 =  x12 & ~x35 & ~x166 & ~x299 & ~x300 & ~x353 & ~x473 & ~x672 & ~x758;
assign c4149 = ~x538 & ~x548 & ~x549 & ~x550 & ~x567 & ~x595 & ~x623 & ~x652 & ~x679 & ~x680 & ~x772;
assign c4151 =  x249 & ~x271 & ~x567;
assign c4153 = ~x347 & ~x350 & ~x374 & ~x393 & ~x407 & ~x434 & ~x435 & ~x449 & ~x463 & ~x476 & ~x715 & ~x754;
assign c4155 = ~x27 & ~x28 & ~x55 & ~x112 & ~x409 & ~x411 & ~x412 & ~x436 & ~x438 & ~x439 & ~x463 & ~x464 & ~x465 & ~x490 & ~x491 & ~x492 & ~x560 & ~x589 & ~x617 & ~x671 & ~x673 & ~x702 & ~x728 & ~x729 & ~x756;
assign c4157 = ~x15 & ~x80 & ~x86 & ~x164 & ~x168 & ~x281 & ~x291 & ~x292 & ~x310 & ~x338 & ~x387 & ~x394 & ~x447 & ~x472 & ~x503 & ~x615 & ~x671 & ~x752 & ~x783;
assign c4159 =  x620 & ~x177 & ~x232 & ~x260 & ~x307;
assign c4161 =  x156 &  x324 & ~x23 & ~x138 & ~x309 & ~x483;
assign c4163 =  x553 & ~x234 & ~x443 & ~x655;
assign c4165 = ~x49 & ~x103 & ~x106 & ~x165 & ~x188 & ~x217 & ~x242 & ~x270 & ~x445 & ~x473 & ~x480 & ~x495 & ~x498 & ~x501 & ~x505 & ~x522 & ~x524 & ~x527 & ~x536 & ~x552 & ~x561 & ~x564 & ~x588 & ~x589 & ~x590 & ~x592 & ~x617 & ~x642 & ~x676;
assign c4167 =  x742 & ~x167 & ~x392 & ~x476 & ~x587 & ~x612 & ~x633 & ~x659 & ~x661 & ~x662 & ~x673 & ~x699 & ~x701;
assign c4169 = ~x5 & ~x6 & ~x23 & ~x53 & ~x60 & ~x61 & ~x63 & ~x86 & ~x88 & ~x116 & ~x118 & ~x127 & ~x144 & ~x145 & ~x146 & ~x172 & ~x200 & ~x305 & ~x313 & ~x365 & ~x421 & ~x422 & ~x472 & ~x491 & ~x731 & ~x760 & ~x780 & ~x783;
assign c4171 =  x315 & ~x10 & ~x35 & ~x39 & ~x65 & ~x93 & ~x94 & ~x144 & ~x172 & ~x586 & ~x675 & ~x701 & ~x757 & ~x775;
assign c4173 =  x371 &  x483 &  x512 & ~x101 & ~x392 & ~x422 & ~x423;
assign c4175 = ~x17 & ~x43 & ~x60 & ~x68 & ~x83 & ~x153 & ~x154 & ~x210 & ~x364 & ~x422 & ~x476 & ~x713 & ~x738 & ~x745 & ~x755 & ~x768 & ~x774;
assign c4177 = ~x290 & ~x317 & ~x464 & ~x600 & ~x603 & ~x604;
assign c4179 = ~x206 & ~x287 & ~x302 & ~x544 & ~x572 & ~x573 & ~x624;
assign c4181 =  x378 & ~x4 & ~x27 & ~x79 & ~x81 & ~x83 & ~x107 & ~x130 & ~x131 & ~x133 & ~x159 & ~x280 & ~x339 & ~x389 & ~x390 & ~x414 & ~x421 & ~x425 & ~x440 & ~x441 & ~x448 & ~x451 & ~x469 & ~x526 & ~x529 & ~x558 & ~x582 & ~x641 & ~x642 & ~x644 & ~x700 & ~x702 & ~x726 & ~x761 & ~x781;
assign c4183 = ~x1 & ~x3 & ~x25 & ~x86 & ~x143 & ~x171 & ~x199 & ~x223 & ~x224 & ~x226 & ~x229 & ~x282 & ~x284 & ~x307 & ~x337 & ~x340 & ~x391 & ~x419 & ~x488 & ~x491 & ~x517 & ~x519 & ~x520 & ~x728 & ~x731 & ~x758 & ~x780;
assign c4185 = ~x3 & ~x123 & ~x314 & ~x342 & ~x370 & ~x447 & ~x456 & ~x709;
assign c4187 =  x75 & ~x558 & ~x598;
assign c4189 = ~x207 & ~x316 & ~x517 & ~x545 & ~x573;
assign c4191 =  x334 & ~x586 & ~x590 & ~x592;
assign c4193 = ~x356 & ~x624 & ~x625 & ~x677 & ~x749;
assign c4195 = ~x3 & ~x24 & ~x29 & ~x31 & ~x59 & ~x141 & ~x169 & ~x195 & ~x251 & ~x278 & ~x281 & ~x307 & ~x337 & ~x396 & ~x398 & ~x422 & ~x425 & ~x427 & ~x445 & ~x451 & ~x452 & ~x455 & ~x458 & ~x470 & ~x472 & ~x473 & ~x485 & ~x486 & ~x487 & ~x499 & ~x500 & ~x509 & ~x511 & ~x512 & ~x515 & ~x527 & ~x528 & ~x534 & ~x536 & ~x538 & ~x560 & ~x590 & ~x673 & ~x675 & ~x726 & ~x730;
assign c4197 =  x509 &  x510 & ~x40 & ~x69 & ~x393 & ~x615 & ~x666 & ~x717 & ~x720 & ~x723 & ~x743 & ~x775 & ~x777 & ~x778;
assign c4199 =  x500 & ~x437 & ~x772;
assign c4201 = ~x27 & ~x289 & ~x318 & ~x401 & ~x544 & ~x573 & ~x699 & ~x772 & ~x773 & ~x776;
assign c4203 =  x288 &  x289 &  x316 & ~x5 & ~x10 & ~x39 & ~x48 & ~x137 & ~x378 & ~x421 & ~x765 & ~x774 & ~x777;
assign c4205 = ~x122 & ~x150 & ~x205 & ~x288 & ~x516 & ~x761;
assign c4207 =  x710 & ~x56 & ~x80 & ~x221 & ~x255 & ~x280 & ~x310 & ~x312 & ~x399 & ~x446 & ~x455;
assign c4209 =  x239 &  x323 & ~x0 & ~x122;
assign c4211 =  x129 &  x157 & ~x483 & ~x566 & ~x586;
assign c4213 =  x250 & ~x624;
assign c4215 =  x274 & ~x65 & ~x335 & ~x745 & ~x775;
assign c4217 =  x405 & ~x2 & ~x3 & ~x131 & ~x452 & ~x481 & ~x496 & ~x498 & ~x507 & ~x522 & ~x524 & ~x527 & ~x529 & ~x532 & ~x553 & ~x565 & ~x591 & ~x592 & ~x593 & ~x619 & ~x621 & ~x645 & ~x673 & ~x676 & ~x703 & ~x726 & ~x729 & ~x732 & ~x756 & ~x759 & ~x760;
assign c4219 =  x380 &  x405 & ~x0 & ~x51 & ~x442 & ~x445 & ~x470 & ~x497 & ~x498 & ~x528 & ~x700;
assign c4221 =  x539 & ~x91 & ~x92 & ~x148 & ~x176 & ~x287;
assign c4223 =  x617;
assign c4225 = ~x25 & ~x27 & ~x55 & ~x206 & ~x281 & ~x309 & ~x317 & ~x334 & ~x335 & ~x337 & ~x363 & ~x392 & ~x393 & ~x448 & ~x475 & ~x476 & ~x503 & ~x559 & ~x587 & ~x644 & ~x781 & ~x782 & ~x783;
assign c4227 =  x428 &  x484 &  x513 &  x569 & ~x85 & ~x111 & ~x250 & ~x421 & ~x422 & ~x423 & ~x783;
assign c4229 =  x540 & ~x0 & ~x57 & ~x60 & ~x108 & ~x119 & ~x137 & ~x138 & ~x147 & ~x173 & ~x174 & ~x199 & ~x201 & ~x202 & ~x228 & ~x229 & ~x230 & ~x250 & ~x251 & ~x257 & ~x279 & ~x284 & ~x285 & ~x310 & ~x336 & ~x393 & ~x530 & ~x532 & ~x728 & ~x756 & ~x760;
assign c4231 = ~x6 & ~x23 & ~x25 & ~x27 & ~x95 & ~x107 & ~x108 & ~x133 & ~x237 & ~x266 & ~x336 & ~x339 & ~x394 & ~x420 & ~x588 & ~x670 & ~x728;
assign c4233 =  x533 & ~x145 & ~x249 & ~x280;
assign c4235 =  x240 &  x295 &  x324 & ~x27 & ~x64;
assign c4237 =  x691 & ~x0 & ~x1 & ~x474 & ~x498 & ~x501 & ~x523 & ~x527 & ~x556 & ~x560;
assign c4239 = ~x56 & ~x224 & ~x229 & ~x286 & ~x314 & ~x341 & ~x342 & ~x363 & ~x368 & ~x424 & ~x474 & ~x475 & ~x502 & ~x602 & ~x603 & ~x631 & ~x632 & ~x727 & ~x755;
assign c4241 =  x487 &  x488 &  x489 & ~x131 & ~x477 & ~x497 & ~x498 & ~x523 & ~x555;
assign c4243 =  x509 & ~x16 & ~x31 & ~x45 & ~x46 & ~x111 & ~x133 & ~x155 & ~x336 & ~x365 & ~x366 & ~x392 & ~x393 & ~x420 & ~x421 & ~x671 & ~x699 & ~x754 & ~x759 & ~x778;
assign c4245 =  x305 & ~x593 & ~x594 & ~x623 & ~x624 & ~x650 & ~x775;
assign c4247 =  x16 &  x150;
assign c4249 =  x455 & ~x124 & ~x144 & ~x292 & ~x365;
assign c4251 =  x468 & ~x94 & ~x95 & ~x121 & ~x308 & ~x586 & ~x727;
assign c4253 = ~x79 & ~x107 & ~x240 & ~x246 & ~x271 & ~x298 & ~x299 & ~x351 & ~x498 & ~x499 & ~x504 & ~x523 & ~x525 & ~x552 & ~x588 & ~x609 & ~x729;
assign c4255 =  x212 &  x240 & ~x56 & ~x113 & ~x168 & ~x223 & ~x624 & ~x652 & ~x653 & ~x773 & ~x776;
assign c4257 = ~x26 & ~x83 & ~x122 & ~x123 & ~x125 & ~x365 & ~x367 & ~x419 & ~x473 & ~x501 & ~x710;
assign c4259 =  x185 & ~x24 & ~x66 & ~x83 & ~x320 & ~x338 & ~x371 & ~x614 & ~x615 & ~x782;
assign c4261 =  x43 & ~x59 & ~x113 & ~x114 & ~x142 & ~x171 & ~x524 & ~x588 & ~x758;
assign c4263 = ~x35 & ~x289 & ~x346 & ~x374 & ~x399 & ~x403 & ~x425 & ~x538;
assign c4265 =  x370 &  x398 &  x482 & ~x74 & ~x83 & ~x449 & ~x737 & ~x771;
assign c4267 =  x189 & ~x94 & ~x149 & ~x588;
assign c4269 = ~x261 & ~x280 & ~x289 & ~x336 & ~x344 & ~x461 & ~x462 & ~x491;
assign c4271 =  x343 & ~x0 & ~x1 & ~x19 & ~x23 & ~x28 & ~x38 & ~x41 & ~x42 & ~x44 & ~x49 & ~x53 & ~x54 & ~x69 & ~x73 & ~x74 & ~x392 & ~x420 & ~x642 & ~x670 & ~x671 & ~x697 & ~x701 & ~x719 & ~x727 & ~x728 & ~x746 & ~x748 & ~x766 & ~x767 & ~x768 & ~x772 & ~x777 & ~x778 & ~x780;
assign c4273 =  x156 & ~x25 & ~x83 & ~x84 & ~x196 & ~x402 & ~x515 & ~x537 & ~x645 & ~x667 & ~x673 & ~x702 & ~x755;
assign c4275 =  x13 & ~x1 & ~x26 & ~x35 & ~x53 & ~x62 & ~x83 & ~x126 & ~x616;
assign c4277 =  x293 &  x715 & ~x89 & ~x355;
assign c4279 =  x395 & ~x597 & ~x651 & ~x654 & ~x679 & ~x706;
assign c4281 =  x216 & ~x176;
assign c4283 =  x744 & ~x83 & ~x130 & ~x140 & ~x164 & ~x250 & ~x447 & ~x633 & ~x662 & ~x663;
assign c4285 =  x428 & ~x75 & ~x105 & ~x107 & ~x109 & ~x156 & ~x348 & ~x393 & ~x421 & ~x422 & ~x766;
assign c4287 =  x157 & ~x35 & ~x37 & ~x54 & ~x224 & ~x593 & ~x594 & ~x620 & ~x672 & ~x696 & ~x727;
assign c4289 = ~x18 & ~x19 & ~x104 & ~x157 & ~x187 & ~x213 & ~x215 & ~x240 & ~x362 & ~x447 & ~x448 & ~x474 & ~x501 & ~x526 & ~x530 & ~x552 & ~x554 & ~x561 & ~x577 & ~x578 & ~x579 & ~x580 & ~x583 & ~x591 & ~x606 & ~x607 & ~x668 & ~x671 & ~x700 & ~x753 & ~x755 & ~x758 & ~x781 & ~x783;
assign c4291 = ~x0 & ~x85 & ~x96 & ~x97 & ~x117 & ~x143 & ~x145 & ~x172 & ~x375 & ~x468 & ~x699 & ~x703 & ~x722 & ~x724 & ~x756 & ~x771;
assign c4293 = ~x20 & ~x27 & ~x152 & ~x153 & ~x179 & ~x360 & ~x418 & ~x419 & ~x420;
assign c4295 = ~x51 & ~x83 & ~x150 & ~x153 & ~x154 & ~x178 & ~x252 & ~x254 & ~x283 & ~x284 & ~x422 & ~x449 & ~x504 & ~x505 & ~x781;
assign c4297 = ~x8 & ~x91 & ~x126 & ~x459 & ~x541 & ~x596 & ~x597 & ~x626 & ~x773 & ~x776;
assign c4299 =  x405 &  x408 & ~x367 & ~x395 & ~x442 & ~x446 & ~x450 & ~x468 & ~x477 & ~x500 & ~x530 & ~x556 & ~x759;
assign c4301 =  x675 & ~x233 & ~x709;
assign c4303 =  x183 &  x239 &  x295 &  x379 & ~x26 & ~x250 & ~x755 & ~x777;
assign c4305 = ~x1 & ~x3 & ~x57 & ~x84 & ~x111 & ~x168 & ~x180 & ~x290 & ~x336 & ~x449 & ~x573 & ~x684;
assign c4307 = ~x192 & ~x202 & ~x231 & ~x249 & ~x370 & ~x462 & ~x659;
assign c4309 =  x210 &  x322 &  x350 & ~x0 & ~x5 & ~x26 & ~x36 & ~x82 & ~x84 & ~x88 & ~x140 & ~x170 & ~x252 & ~x253 & ~x308 & ~x336 & ~x776;
assign c4311 =  x156 &  x297 & ~x303 & ~x313 & ~x341;
assign c4313 = ~x3 & ~x24 & ~x55 & ~x56 & ~x57 & ~x59 & ~x140 & ~x167 & ~x198 & ~x226 & ~x281 & ~x283 & ~x309 & ~x312 & ~x334 & ~x337 & ~x360 & ~x363 & ~x391 & ~x420 & ~x421 & ~x447 & ~x448 & ~x473 & ~x475 & ~x476 & ~x503 & ~x600 & ~x602 & ~x603 & ~x630 & ~x632 & ~x727;
assign c4315 =  x742 & ~x55 & ~x134 & ~x161 & ~x190 & ~x222 & ~x271 & ~x326 & ~x363 & ~x394 & ~x446 & ~x448 & ~x450 & ~x527 & ~x556 & ~x581 & ~x610 & ~x669 & ~x672;
assign c4317 =  x239 &  x267 & ~x59 & ~x87 & ~x103 & ~x116 & ~x171 & ~x198 & ~x278 & ~x283 & ~x309 & ~x726 & ~x781;
assign c4319 = ~x2 & ~x3 & ~x19 & ~x27 & ~x31 & ~x57 & ~x78 & ~x106 & ~x111 & ~x112 & ~x136 & ~x167 & ~x195 & ~x270 & ~x271 & ~x475 & ~x499 & ~x501 & ~x524 & ~x525 & ~x528 & ~x537 & ~x554 & ~x558 & ~x577 & ~x578 & ~x580 & ~x582 & ~x583 & ~x584 & ~x586 & ~x588 & ~x589 & ~x590 & ~x592 & ~x593 & ~x611 & ~x616 & ~x617 & ~x621 & ~x638 & ~x645 & ~x646 & ~x647 & ~x649 & ~x671 & ~x676 & ~x678 & ~x702 & ~x704 & ~x728 & ~x756 & ~x760 & ~x763 & ~x782;
assign c4321 =  x743 & ~x106 & ~x162 & ~x187 & ~x215 & ~x271 & ~x555 & ~x583 & ~x609 & ~x611 & ~x639;
assign c4323 =  x417 &  x445 & ~x39 & ~x49 & ~x357 & ~x641 & ~x670;
assign c4325 =  x594 & ~x25 & ~x53 & ~x81 & ~x140 & ~x142 & ~x165 & ~x171 & ~x192 & ~x193 & ~x225 & ~x227 & ~x229 & ~x250 & ~x251 & ~x276 & ~x277 & ~x304 & ~x309 & ~x311 & ~x335 & ~x336 & ~x337 & ~x363 & ~x369 & ~x394 & ~x419 & ~x423 & ~x424 & ~x478 & ~x615 & ~x641 & ~x753 & ~x754;
assign c4327 =  x667 & ~x26 & ~x56 & ~x84 & ~x224 & ~x390 & ~x420 & ~x529 & ~x558 & ~x727 & ~x775 & ~x776 & ~x783;
assign c4329 =  x299 & ~x27 & ~x28 & ~x56 & ~x69 & ~x95 & ~x123 & ~x333 & ~x334 & ~x335 & ~x363 & ~x755;
assign c4331 = ~x158 & ~x268 & ~x393 & ~x504 & ~x575 & ~x577 & ~x579 & ~x607 & ~x619 & ~x642 & ~x643 & ~x698 & ~x727;
assign c4333 =  x290 &  x459 &  x460 &  x489 & ~x526 & ~x560;
assign c4335 =  x236 & ~x27 & ~x49 & ~x50 & ~x192 & ~x298 & ~x364 & ~x467 & ~x470 & ~x493 & ~x497 & ~x639 & ~x640 & ~x695 & ~x729;
assign c4337 = ~x1 & ~x5 & ~x20 & ~x24 & ~x25 & ~x26 & ~x48 & ~x49 & ~x50 & ~x53 & ~x77 & ~x79 & ~x80 & ~x103 & ~x104 & ~x105 & ~x133 & ~x364 & ~x393 & ~x420 & ~x421 & ~x449 & ~x465 & ~x466 & ~x468 & ~x469 & ~x471 & ~x504 & ~x615 & ~x642 & ~x676 & ~x703 & ~x727 & ~x729 & ~x754 & ~x757 & ~x782 & ~x783;
assign c4339 = ~x32 & ~x112 & ~x194 & ~x423 & ~x428 & ~x448 & ~x449 & ~x487 & ~x489 & ~x563 & ~x564 & ~x585 & ~x612 & ~x646 & ~x783;
assign c4341 = ~x490 & ~x491 & ~x493 & ~x519 & ~x520 & ~x522 & ~x532 & ~x597 & ~x625 & ~x644 & ~x775 & ~x778;
assign c4343 = ~x52 & ~x69 & ~x82 & ~x98 & ~x139 & ~x140 & ~x309 & ~x348 & ~x365 & ~x420 & ~x474 & ~x476 & ~x502 & ~x559 & ~x682 & ~x685;
assign c4345 = ~x131 & ~x248 & ~x393 & ~x631 & ~x632 & ~x633 & ~x635 & ~x636 & ~x637 & ~x646 & ~x667 & ~x753;
assign c4347 =  x508 &  x536 &  x564 & ~x65 & ~x421 & ~x774;
assign c4349 = ~x43 & ~x69 & ~x71 & ~x96 & ~x206 & ~x625 & ~x653 & ~x682 & ~x708 & ~x709;
assign c4351 = ~x3 & ~x32 & ~x81 & ~x84 & ~x85 & ~x111 & ~x112 & ~x139 & ~x140 & ~x168 & ~x193 & ~x196 & ~x222 & ~x249 & ~x253 & ~x277 & ~x279 & ~x280 & ~x309 & ~x333 & ~x338 & ~x339 & ~x363 & ~x366 & ~x394 & ~x395 & ~x419 & ~x450 & ~x559 & ~x599 & ~x601 & ~x614 & ~x616 & ~x630 & ~x631 & ~x643 & ~x644 & ~x672 & ~x728 & ~x752 & ~x755 & ~x758 & ~x781 & ~x782 & ~x783;
assign c4353 =  x611 &  x648 & ~x654 & ~x710;
assign c4355 = ~x56 & ~x97 & ~x168 & ~x170 & ~x261 & ~x316 & ~x654 & ~x710;
assign c4357 = ~x25 & ~x26 & ~x28 & ~x35 & ~x53 & ~x58 & ~x91 & ~x110 & ~x116 & ~x119 & ~x120 & ~x145 & ~x146 & ~x147 & ~x172 & ~x175 & ~x181 & ~x182 & ~x199 & ~x230 & ~x252 & ~x254 & ~x281 & ~x282 & ~x310 & ~x728 & ~x754 & ~x755 & ~x782;
assign c4359 =  x301 & ~x27 & ~x83 & ~x154 & ~x365 & ~x415;
assign c4361 =  x239 &  x351 & ~x138 & ~x428 & ~x432 & ~x455;
assign c4363 =  x185 &  x213 & ~x3 & ~x29 & ~x55 & ~x56 & ~x60 & ~x111 & ~x138 & ~x455 & ~x456 & ~x484 & ~x587 & ~x642 & ~x725 & ~x726;
assign c4365 =  x323 &  x349 &  x351 & ~x19 & ~x21 & ~x28 & ~x29 & ~x32 & ~x33 & ~x34 & ~x35 & ~x54 & ~x57 & ~x61 & ~x83 & ~x85 & ~x113 & ~x199 & ~x252 & ~x305 & ~x308 & ~x560 & ~x587 & ~x617 & ~x644 & ~x757;
assign c4367 =  x743 &  x745 & ~x8 & ~x163 & ~x168 & ~x638;
assign c4369 = ~x1 & ~x2 & ~x6 & ~x30 & ~x49 & ~x51 & ~x54 & ~x77 & ~x82 & ~x83 & ~x107 & ~x131 & ~x138 & ~x156 & ~x157 & ~x159 & ~x161 & ~x167 & ~x186 & ~x188 & ~x189 & ~x212 & ~x214 & ~x215 & ~x223 & ~x240 & ~x242 & ~x243 & ~x244 & ~x269 & ~x270 & ~x297 & ~x324 & ~x337 & ~x394 & ~x472 & ~x476 & ~x498 & ~x504 & ~x526 & ~x529 & ~x554 & ~x556 & ~x557 & ~x559 & ~x582 & ~x583 & ~x584 & ~x610 & ~x613 & ~x618 & ~x644 & ~x646 & ~x674 & ~x696 & ~x702 & ~x755 & ~x758 & ~x761 & ~x783;
assign c4371 = ~x262 & ~x514 & ~x597 & ~x628 & ~x658;
assign c4373 =  x269 &  x321 & ~x413 & ~x705 & ~x734 & ~x779;
assign c4375 = ~x1 & ~x2 & ~x21 & ~x25 & ~x26 & ~x28 & ~x47 & ~x50 & ~x53 & ~x54 & ~x58 & ~x80 & ~x81 & ~x83 & ~x111 & ~x437 & ~x438 & ~x440 & ~x441 & ~x442 & ~x455 & ~x466 & ~x467 & ~x470 & ~x481 & ~x482 & ~x496 & ~x506 & ~x524 & ~x531 & ~x535 & ~x537 & ~x563 & ~x587 & ~x591 & ~x594 & ~x614 & ~x617 & ~x619 & ~x621 & ~x644 & ~x645 & ~x648 & ~x649 & ~x650 & ~x651 & ~x700 & ~x701 & ~x702 & ~x706 & ~x726 & ~x729 & ~x730 & ~x734 & ~x752 & ~x783;
assign c4377 = ~x0 & ~x1 & ~x23 & ~x26 & ~x69 & ~x112 & ~x290 & ~x303 & ~x309 & ~x318 & ~x319 & ~x364 & ~x655 & ~x684;
assign c4379 =  x268 &  x294 &  x296 & ~x118 & ~x251 & ~x356 & ~x645 & ~x701;
assign c4381 =  x316 &  x361 & ~x8 & ~x27 & ~x48 & ~x694 & ~x704 & ~x705 & ~x758;
assign c4383 = ~x1 & ~x26 & ~x56 & ~x58 & ~x59 & ~x79 & ~x88 & ~x407 & ~x434 & ~x435 & ~x536 & ~x576 & ~x589 & ~x592 & ~x646 & ~x648 & ~x673 & ~x721 & ~x749;
assign c4385 =  x267 &  x324 &  x352 &  x380 & ~x30 & ~x53 & ~x112 & ~x141 & ~x145 & ~x171 & ~x252 & ~x277 & ~x308 & ~x761 & ~x781;
assign c4387 = ~x96 & ~x123 & ~x151 & ~x178 & ~x363 & ~x390 & ~x418 & ~x421 & ~x475 & ~x476 & ~x681;
assign c4389 =  x741 &  x742 & ~x84 & ~x106 & ~x161 & ~x248 & ~x249 & ~x307 & ~x309 & ~x529 & ~x661;
assign c4391 = ~x77 & ~x97 & ~x112 & ~x125 & ~x126 & ~x151 & ~x153 & ~x395 & ~x472 & ~x504 & ~x528 & ~x616 & ~x671 & ~x700 & ~x709;
assign c4393 =  x566 & ~x7 & ~x76 & ~x86 & ~x192 & ~x201 & ~x220 & ~x249 & ~x278 & ~x334 & ~x335 & ~x338 & ~x340 & ~x364 & ~x393 & ~x394 & ~x421 & ~x443 & ~x643 & ~x755;
assign c4395 = ~x114 & ~x252 & ~x312 & ~x363 & ~x532 & ~x600 & ~x603 & ~x613 & ~x632 & ~x633 & ~x697 & ~x781;
assign c4397 =  x399 &  x446 & ~x48;
assign c4399 =  x268 & ~x151 & ~x316;
assign c4401 = ~x230 & ~x256 & ~x259 & ~x286 & ~x345 & ~x363 & ~x365 & ~x373 & ~x375 & ~x392 & ~x450 & ~x502 & ~x557 & ~x558 & ~x559 & ~x615 & ~x616 & ~x698 & ~x699;
assign c4403 =  x344 & ~x9 & ~x11 & ~x37 & ~x38 & ~x48 & ~x79 & ~x116 & ~x133 & ~x167 & ~x172 & ~x678 & ~x699 & ~x712 & ~x756 & ~x766 & ~x779;
assign c4405 =  x315 &  x343 &  x388 & ~x30 & ~x705;
assign c4407 =  x480 &  x515 &  x544;
assign c4409 = ~x2 & ~x5 & ~x21 & ~x27 & ~x32 & ~x59 & ~x400 & ~x427 & ~x455 & ~x457 & ~x458 & ~x484 & ~x486 & ~x513 & ~x515 & ~x516 & ~x536 & ~x541 & ~x564 & ~x568 & ~x616 & ~x621 & ~x644 & ~x648 & ~x667 & ~x668 & ~x669 & ~x672 & ~x694 & ~x697 & ~x700 & ~x702 & ~x726 & ~x727 & ~x728 & ~x782;
assign c4411 = ~x0 & ~x27 & ~x29 & ~x54 & ~x168 & ~x280 & ~x309 & ~x335 & ~x363 & ~x391 & ~x394 & ~x446 & ~x448 & ~x449 & ~x460 & ~x626 & ~x657 & ~x686 & ~x687 & ~x688;
assign c4413 = ~x78 & ~x105 & ~x187 & ~x422 & ~x448 & ~x452 & ~x498 & ~x500 & ~x507 & ~x508 & ~x527 & ~x529 & ~x548 & ~x549 & ~x550 & ~x551 & ~x562 & ~x580 & ~x581 & ~x582 & ~x589 & ~x591 & ~x617 & ~x675 & ~x705 & ~x728 & ~x732 & ~x734 & ~x757 & ~x783;
assign c4415 =  x278 & ~x624;
assign c4417 =  x286 & ~x503 & ~x599 & ~x600 & ~x627;
assign c4419 = ~x23 & ~x27 & ~x223 & ~x224 & ~x280 & ~x335 & ~x343 & ~x371 & ~x400 & ~x424 & ~x429 & ~x452 & ~x458 & ~x459 & ~x461 & ~x473 & ~x476 & ~x483 & ~x499 & ~x502 & ~x556 & ~x588 & ~x590 & ~x611 & ~x613 & ~x616 & ~x619 & ~x642 & ~x643 & ~x646 & ~x647 & ~x672 & ~x673 & ~x702 & ~x704 & ~x727 & ~x728 & ~x758;
assign c4421 =  x674 & ~x346 & ~x678;
assign c4423 =  x263 &  x461 & ~x31 & ~x336 & ~x496 & ~x497 & ~x524 & ~x532 & ~x587 & ~x671;
assign c4425 = ~x4 & ~x8 & ~x25 & ~x28 & ~x33 & ~x47 & ~x48 & ~x73 & ~x75 & ~x76 & ~x103 & ~x482 & ~x501 & ~x508 & ~x522 & ~x523 & ~x524 & ~x525 & ~x531 & ~x552 & ~x563 & ~x564 & ~x581 & ~x589 & ~x591 & ~x593 & ~x645 & ~x652 & ~x668 & ~x669 & ~x680 & ~x696 & ~x699 & ~x700 & ~x705 & ~x706 & ~x726 & ~x731 & ~x737 & ~x751 & ~x753;
assign c4427 = ~x17 & ~x27 & ~x44 & ~x54 & ~x55 & ~x77 & ~x78 & ~x79 & ~x80 & ~x104 & ~x106 & ~x140 & ~x167 & ~x507 & ~x528 & ~x529 & ~x536 & ~x548 & ~x549 & ~x551 & ~x553 & ~x557 & ~x563 & ~x583 & ~x590 & ~x612 & ~x615 & ~x620 & ~x642 & ~x668 & ~x723 & ~x754 & ~x761 & ~x783;
assign c4429 = ~x3 & ~x26 & ~x28 & ~x31 & ~x37 & ~x63 & ~x91 & ~x117 & ~x546 & ~x547 & ~x548 & ~x591 & ~x617 & ~x672 & ~x756 & ~x757;
assign c4431 =  x647 & ~x233 & ~x335;
assign c4433 =  x128 & ~x25 & ~x27 & ~x513 & ~x536 & ~x542 & ~x597 & ~x623;
assign c4435 =  x716 & ~x0 & ~x27 & ~x50 & ~x54 & ~x105 & ~x308 & ~x336 & ~x364 & ~x392 & ~x501 & ~x504 & ~x529 & ~x585 & ~x605 & ~x611 & ~x612 & ~x634 & ~x642 & ~x728 & ~x729 & ~x755 & ~x759 & ~x783;
assign c4437 =  x259 &  x483 &  x508 &  x509 & ~x448 & ~x476;
assign c4439 =  x194 & ~x744;
assign c4441 = ~x1 & ~x13 & ~x22 & ~x26 & ~x28 & ~x29 & ~x37 & ~x39 & ~x41 & ~x55 & ~x60 & ~x65 & ~x69 & ~x80 & ~x86 & ~x106 & ~x137 & ~x138 & ~x142 & ~x145 & ~x196 & ~x559 & ~x561 & ~x563 & ~x616 & ~x645 & ~x646 & ~x647 & ~x673 & ~x704 & ~x728 & ~x756 & ~x774 & ~x783;
assign c4443 = ~x24 & ~x25 & ~x55 & ~x56 & ~x223 & ~x224 & ~x226 & ~x445 & ~x447 & ~x474 & ~x475 & ~x502 & ~x504 & ~x531 & ~x533 & ~x544 & ~x560 & ~x584 & ~x588 & ~x600 & ~x616 & ~x617 & ~x627 & ~x628 & ~x630 & ~x643 & ~x644 & ~x657 & ~x698 & ~x782 & ~x783;
assign c4445 =  x515 & ~x25 & ~x50 & ~x60 & ~x62 & ~x105 & ~x134 & ~x193 & ~x223 & ~x408 & ~x552 & ~x678 & ~x705 & ~x728 & ~x733 & ~x734 & ~x756;
assign c4447 = ~x77 & ~x159 & ~x217 & ~x244 & ~x532 & ~x564 & ~x586 & ~x620 & ~x631 & ~x632 & ~x638 & ~x643 & ~x661 & ~x664;
assign c4449 = ~x9 & ~x24 & ~x27 & ~x34 & ~x56 & ~x61 & ~x89 & ~x485 & ~x514 & ~x541 & ~x570 & ~x572 & ~x596 & ~x597 & ~x601 & ~x624 & ~x643 & ~x670 & ~x671 & ~x727 & ~x782;
assign c4451 = ~x1 & ~x8 & ~x26 & ~x29 & ~x49 & ~x61 & ~x112 & ~x356 & ~x379 & ~x565 & ~x617 & ~x621 & ~x622 & ~x643 & ~x644 & ~x651 & ~x673 & ~x699 & ~x703 & ~x704 & ~x722 & ~x724 & ~x753 & ~x772 & ~x773 & ~x777 & ~x779 & ~x781;
assign c4453 = ~x112 & ~x139 & ~x196 & ~x229 & ~x314 & ~x385 & ~x420 & ~x434 & ~x435 & ~x442 & ~x455 & ~x533 & ~x584 & ~x586 & ~x699;
assign c4455 =  x322 &  x323 & ~x132 & ~x168 & ~x310 & ~x410 & ~x732 & ~x754 & ~x762;
assign c4457 = ~x344 & ~x372 & ~x545 & ~x548 & ~x573 & ~x576;
assign c4459 =  x373 &  x389 & ~x680 & ~x681;
assign c4461 = ~x0 & ~x2 & ~x21 & ~x83 & ~x112 & ~x195 & ~x341 & ~x361 & ~x369 & ~x393 & ~x397 & ~x400 & ~x414 & ~x441 & ~x444 & ~x446 & ~x447 & ~x448 & ~x451 & ~x452 & ~x455 & ~x456 & ~x458 & ~x460 & ~x477 & ~x501 & ~x560 & ~x561 & ~x587 & ~x639 & ~x671 & ~x695 & ~x728 & ~x729 & ~x760;
assign c4463 =  x452 &  x508 &  x535 & ~x75 & ~x103 & ~x133 & ~x309 & ~x393 & ~x777;
assign c4465 =  x713 & ~x159 & ~x631 & ~x634 & ~x647;
assign c4467 =  x219 & ~x243 & ~x529;
assign c4469 = ~x1 & ~x24 & ~x47 & ~x74 & ~x81 & ~x83 & ~x105 & ~x107 & ~x132 & ~x133 & ~x135 & ~x138 & ~x139 & ~x160 & ~x162 & ~x191 & ~x242 & ~x244 & ~x297 & ~x422 & ~x472 & ~x474 & ~x499 & ~x501 & ~x502 & ~x503 & ~x524 & ~x529 & ~x530 & ~x531 & ~x550 & ~x553 & ~x555 & ~x644 & ~x646 & ~x703 & ~x728 & ~x731 & ~x781;
assign c4471 =  x333 & ~x63 & ~x593 & ~x649 & ~x731 & ~x771;
assign c4473 = ~x2 & ~x4 & ~x5 & ~x18 & ~x20 & ~x21 & ~x22 & ~x24 & ~x25 & ~x29 & ~x32 & ~x39 & ~x42 & ~x47 & ~x52 & ~x54 & ~x57 & ~x75 & ~x156 & ~x392 & ~x393 & ~x720 & ~x722 & ~x733 & ~x739 & ~x741 & ~x744 & ~x745 & ~x746 & ~x756 & ~x763 & ~x770 & ~x771 & ~x772 & ~x776 & ~x779 & ~x780 & ~x781 & ~x782;
assign c4475 =  x434 &  x604 & ~x653;
assign c4477 = ~x2 & ~x3 & ~x5 & ~x7 & ~x8 & ~x21 & ~x23 & ~x32 & ~x33 & ~x36 & ~x53 & ~x55 & ~x62 & ~x80 & ~x86 & ~x87 & ~x106 & ~x107 & ~x138 & ~x166 & ~x197 & ~x198 & ~x224 & ~x256 & ~x308 & ~x309 & ~x311 & ~x333 & ~x364 & ~x421 & ~x446 & ~x447 & ~x450 & ~x452 & ~x471 & ~x473 & ~x474 & ~x475 & ~x479 & ~x501 & ~x503 & ~x508 & ~x523 & ~x526 & ~x534 & ~x552 & ~x553 & ~x557 & ~x558 & ~x560 & ~x563 & ~x611 & ~x613 & ~x615 & ~x616 & ~x619 & ~x621 & ~x639 & ~x642 & ~x645 & ~x646 & ~x647 & ~x674 & ~x677 & ~x699 & ~x701 & ~x702 & ~x706 & ~x733 & ~x753 & ~x755 & ~x782 & ~x783;
assign c4479 = ~x8 & ~x21 & ~x35 & ~x69 & ~x598 & ~x627 & ~x667 & ~x679 & ~x734 & ~x744;
assign c4481 =  x713 &  x742 & ~x222 & ~x365 & ~x444 & ~x585 & ~x661;
assign c4483 =  x596 & ~x3 & ~x22 & ~x23 & ~x25 & ~x26 & ~x28 & ~x31 & ~x52 & ~x53 & ~x59 & ~x79 & ~x80 & ~x81 & ~x106 & ~x108 & ~x110 & ~x111 & ~x113 & ~x138 & ~x142 & ~x195 & ~x223 & ~x224 & ~x226 & ~x228 & ~x251 & ~x252 & ~x255 & ~x256 & ~x257 & ~x281 & ~x284 & ~x305 & ~x306 & ~x309 & ~x310 & ~x312 & ~x335 & ~x338 & ~x340 & ~x341 & ~x342 & ~x362 & ~x365 & ~x366 & ~x370 & ~x389 & ~x392 & ~x395 & ~x397 & ~x415 & ~x424 & ~x425 & ~x443 & ~x445 & ~x448 & ~x449 & ~x451 & ~x471 & ~x472 & ~x473 & ~x479 & ~x480 & ~x504 & ~x558 & ~x561 & ~x588 & ~x640 & ~x643 & ~x697 & ~x726 & ~x727 & ~x728 & ~x780 & ~x782;
assign c4485 = ~x13 & ~x25 & ~x27 & ~x49 & ~x80 & ~x134 & ~x160 & ~x203 & ~x255 & ~x271 & ~x279 & ~x311 & ~x339 & ~x471 & ~x496 & ~x498 & ~x501 & ~x502 & ~x524 & ~x529 & ~x563 & ~x564 & ~x582 & ~x585 & ~x592 & ~x638 & ~x676 & ~x696 & ~x702 & ~x704 & ~x781;
assign c4487 =  x239 &  x267 &  x351 & ~x4 & ~x24 & ~x28 & ~x51 & ~x54 & ~x55 & ~x79 & ~x106 & ~x108 & ~x109 & ~x112 & ~x136 & ~x164 & ~x166 & ~x169 & ~x194 & ~x226 & ~x251 & ~x283 & ~x309 & ~x310 & ~x505 & ~x560 & ~x672 & ~x697 & ~x700 & ~x727 & ~x755 & ~x779 & ~x780 & ~x781;
assign c4489 = ~x189 & ~x242 & ~x386 & ~x519 & ~x524 & ~x619;
assign c4491 =  x376 &  x433 & ~x338 & ~x368 & ~x473 & ~x498 & ~x532 & ~x590 & ~x593 & ~x620 & ~x705;
assign c4493 =  x484 &  x486 &  x488 &  x513 & ~x25 & ~x46 & ~x48 & ~x49 & ~x74 & ~x280 & ~x763 & ~x778 & ~x783;
assign c4495 =  x457 & ~x11 & ~x104 & ~x134 & ~x156 & ~x379 & ~x422 & ~x727 & ~x773 & ~x776;
assign c4497 =  x433 &  x435 &  x436 & ~x336 & ~x421 & ~x448 & ~x470 & ~x472 & ~x505 & ~x554 & ~x757 & ~x783;
assign c4499 =  x741 &  x743 & ~x506 & ~x660 & ~x730;
assign c50 =  x27;
assign c52 = ~x0 & ~x26 & ~x55 & ~x77 & ~x81 & ~x82 & ~x87 & ~x106 & ~x138 & ~x146 & ~x163 & ~x193 & ~x224 & ~x247 & ~x248 & ~x252 & ~x308 & ~x326 & ~x334 & ~x336 & ~x352 & ~x355 & ~x379 & ~x381 & ~x407 & ~x408 & ~x409 & ~x414 & ~x435 & ~x439 & ~x464 & ~x465 & ~x469 & ~x471 & ~x494 & ~x495 & ~x496 & ~x498 & ~x499 & ~x502 & ~x527 & ~x588 & ~x672 & ~x727;
assign c54 =  x308;
assign c56 = ~x21 & ~x23 & ~x29 & ~x52 & ~x54 & ~x55 & ~x57 & ~x78 & ~x79 & ~x81 & ~x82 & ~x87 & ~x106 & ~x107 & ~x109 & ~x110 & ~x111 & ~x113 & ~x134 & ~x137 & ~x140 & ~x142 & ~x163 & ~x164 & ~x165 & ~x166 & ~x169 & ~x170 & ~x192 & ~x195 & ~x196 & ~x197 & ~x198 & ~x200 & ~x219 & ~x220 & ~x221 & ~x222 & ~x223 & ~x224 & ~x248 & ~x249 & ~x277 & ~x279 & ~x282 & ~x302 & ~x306 & ~x309 & ~x312 & ~x330 & ~x331 & ~x335 & ~x337 & ~x357 & ~x358 & ~x359 & ~x362 & ~x364 & ~x378 & ~x379 & ~x380 & ~x381 & ~x387 & ~x388 & ~x409 & ~x415 & ~x422 & ~x436 & ~x443 & ~x444 & ~x465 & ~x470 & ~x473 & ~x498 & ~x499 & ~x502 & ~x527 & ~x528 & ~x530 & ~x555 & ~x558 & ~x561 & ~x585 & ~x586 & ~x587 & ~x612 & ~x640 & ~x645 & ~x670 & ~x673 & ~x699 & ~x727 & ~x729 & ~x754 & ~x757 & ~x783;
assign c58 = ~x0 & ~x20 & ~x21 & ~x23 & ~x24 & ~x25 & ~x26 & ~x27 & ~x32 & ~x33 & ~x34 & ~x56 & ~x62 & ~x81 & ~x82 & ~x86 & ~x88 & ~x90 & ~x106 & ~x110 & ~x111 & ~x112 & ~x114 & ~x116 & ~x134 & ~x138 & ~x142 & ~x163 & ~x190 & ~x192 & ~x193 & ~x199 & ~x218 & ~x244 & ~x246 & ~x247 & ~x252 & ~x272 & ~x276 & ~x277 & ~x279 & ~x335 & ~x338 & ~x361 & ~x388 & ~x390 & ~x392 & ~x393 & ~x418 & ~x422 & ~x423 & ~x474 & ~x504 & ~x508 & ~x532 & ~x543 & ~x544 & ~x558 & ~x560 & ~x571 & ~x583 & ~x589 & ~x591 & ~x592 & ~x594 & ~x599 & ~x614 & ~x615 & ~x616 & ~x618 & ~x619 & ~x624 & ~x626 & ~x640 & ~x643 & ~x653 & ~x655 & ~x678 & ~x699 & ~x702 & ~x703 & ~x708 & ~x728 & ~x731 & ~x733 & ~x754 & ~x755 & ~x758 & ~x783;
assign c510 =  x425 & ~x1 & ~x41 & ~x42 & ~x54 & ~x69 & ~x113 & ~x122 & ~x142 & ~x254 & ~x281 & ~x309 & ~x310 & ~x319 & ~x320 & ~x321 & ~x322 & ~x323 & ~x349 & ~x350 & ~x365 & ~x375 & ~x376 & ~x377 & ~x402 & ~x403 & ~x404 & ~x405 & ~x407 & ~x430 & ~x476 & ~x589 & ~x615 & ~x616 & ~x642 & ~x643 & ~x739 & ~x756;
assign c512 =  x684 & ~x245 & ~x247 & ~x296 & ~x329 & ~x330 & ~x351 & ~x360 & ~x361 & ~x387 & ~x518 & ~x558 & ~x650;
assign c514 = ~x142 & ~x200 & ~x312 & ~x360 & ~x361 & ~x378 & ~x380 & ~x381 & ~x382 & ~x383 & ~x396 & ~x416 & ~x519 & ~x529 & ~x546 & ~x762;
assign c516 = ~x109 & ~x166 & ~x222 & ~x295 & ~x298 & ~x350 & ~x380 & ~x409 & ~x411 & ~x421 & ~x519 & ~x623 & ~x640 & ~x735;
assign c518 =  x228 &  x302 &  x416;
assign c520 =  x691 &  x718 & ~x37 & ~x81 & ~x166 & ~x192 & ~x220 & ~x250 & ~x275 & ~x276 & ~x334 & ~x360 & ~x381 & ~x409 & ~x443 & ~x465 & ~x466 & ~x472 & ~x473 & ~x502 & ~x527 & ~x528;
assign c522 = ~x52 & ~x354 & ~x406 & ~x448 & ~x462 & ~x497 & ~x526 & ~x555 & ~x579 & ~x580 & ~x611 & ~x687 & ~x689 & ~x690 & ~x718;
assign c524 = ~x28 & ~x65 & ~x79 & ~x87 & ~x122 & ~x150 & ~x292 & ~x293 & ~x308 & ~x337 & ~x350 & ~x458 & ~x485 & ~x486 & ~x540 & ~x595 & ~x596 & ~x655 & ~x656 & ~x685 & ~x711 & ~x740 & ~x769;
assign c526 =  x275 & ~x92 & ~x205 & ~x267 & ~x292 & ~x298 & ~x486;
assign c528 =  x209 &  x292 &  x319 &  x347 & ~x19 & ~x54 & ~x78 & ~x90 & ~x92 & ~x134 & ~x165 & ~x197 & ~x219 & ~x249 & ~x253 & ~x270 & ~x271 & ~x272 & ~x282 & ~x308 & ~x329 & ~x336 & ~x343 & ~x367 & ~x370 & ~x396 & ~x449 & ~x475 & ~x478 & ~x528 & ~x529 & ~x556 & ~x559 & ~x561 & ~x597 & ~x649 & ~x652 & ~x697 & ~x706 & ~x724 & ~x734 & ~x756;
assign c530 =  x371 & ~x20 & ~x32 & ~x47 & ~x53 & ~x80 & ~x113 & ~x152 & ~x180 & ~x336 & ~x351 & ~x366 & ~x377 & ~x393 & ~x407 & ~x422 & ~x434 & ~x435 & ~x488 & ~x504 & ~x624 & ~x679 & ~x680 & ~x709 & ~x725 & ~x737 & ~x738 & ~x740 & ~x750 & ~x752 & ~x769 & ~x772 & ~x782;
assign c532 =  x415 & ~x20 & ~x32 & ~x34 & ~x103 & ~x437 & ~x549 & ~x576 & ~x656 & ~x658 & ~x666 & ~x712 & ~x743 & ~x744 & ~x751 & ~x754;
assign c534 = ~x4 & ~x6 & ~x45 & ~x46 & ~x52 & ~x57 & ~x59 & ~x77 & ~x79 & ~x85 & ~x109 & ~x165 & ~x166 & ~x280 & ~x467 & ~x496 & ~x523 & ~x549 & ~x553 & ~x578 & ~x605 & ~x628 & ~x636 & ~x638 & ~x639 & ~x665 & ~x666 & ~x680 & ~x685 & ~x737 & ~x757 & ~x769;
assign c536 =  x330 &  x359 &  x444 & ~x235 & ~x407;
assign c538 =  x372 & ~x1 & ~x19 & ~x22 & ~x25 & ~x78 & ~x79 & ~x409 & ~x421 & ~x439 & ~x504 & ~x602 & ~x667 & ~x706 & ~x707 & ~x758 & ~x759;
assign c540 = ~x30 & ~x45 & ~x54 & ~x59 & ~x82 & ~x111 & ~x121 & ~x150 & ~x177 & ~x180 & ~x205 & ~x209 & ~x233 & ~x235 & ~x261 & ~x262 & ~x263 & ~x346 & ~x347 & ~x401 & ~x403 & ~x458 & ~x540 & ~x706 & ~x709 & ~x711 & ~x739;
assign c542 =  x484 & ~x50 & ~x517 & ~x545 & ~x574 & ~x607 & ~x722 & ~x741 & ~x763 & ~x768 & ~x776;
assign c544 =  x760;
assign c546 = ~x6 & ~x49 & ~x81 & ~x82 & ~x83 & ~x106 & ~x135 & ~x136 & ~x140 & ~x307 & ~x435 & ~x517 & ~x522 & ~x523 & ~x546 & ~x547 & ~x552 & ~x579 & ~x609 & ~x632 & ~x658 & ~x661 & ~x663 & ~x688 & ~x711 & ~x720 & ~x721 & ~x769;
assign c548 =  x717 & ~x4 & ~x21 & ~x28 & ~x29 & ~x50 & ~x55 & ~x58 & ~x81 & ~x82 & ~x107 & ~x108 & ~x109 & ~x110 & ~x111 & ~x113 & ~x163 & ~x165 & ~x167 & ~x170 & ~x191 & ~x193 & ~x196 & ~x199 & ~x223 & ~x225 & ~x226 & ~x249 & ~x250 & ~x253 & ~x278 & ~x281 & ~x302 & ~x304 & ~x305 & ~x306 & ~x307 & ~x311 & ~x333 & ~x334 & ~x337 & ~x359 & ~x360 & ~x363 & ~x365 & ~x381 & ~x390 & ~x392 & ~x393 & ~x409 & ~x414 & ~x415 & ~x419 & ~x421 & ~x437 & ~x443 & ~x444 & ~x448 & ~x449 & ~x470 & ~x471 & ~x472 & ~x474 & ~x475 & ~x476 & ~x499 & ~x500 & ~x501 & ~x504 & ~x505 & ~x530 & ~x556 & ~x558 & ~x561 & ~x562 & ~x586 & ~x588 & ~x614 & ~x617 & ~x641 & ~x643 & ~x671 & ~x673 & ~x682 & ~x699 & ~x710 & ~x726 & ~x764;
assign c550 =  x279;
assign c552 = ~x2 & ~x10 & ~x23 & ~x63 & ~x86 & ~x87 & ~x91 & ~x114 & ~x119 & ~x121 & ~x145 & ~x150 & ~x157 & ~x183 & ~x184 & ~x203 & ~x267 & ~x299 & ~x458 & ~x671 & ~x682 & ~x721 & ~x726 & ~x756 & ~x764 & ~x778;
assign c554 = ~x8 & ~x18 & ~x20 & ~x26 & ~x31 & ~x47 & ~x51 & ~x75 & ~x84 & ~x364 & ~x392 & ~x448 & ~x467 & ~x494 & ~x522 & ~x553 & ~x580 & ~x598 & ~x626 & ~x636 & ~x638 & ~x654 & ~x661 & ~x671 & ~x688 & ~x695 & ~x698 & ~x707 & ~x712 & ~x713 & ~x726 & ~x751 & ~x767 & ~x770;
assign c556 =  x484 &  x485 &  x512 & ~x48 & ~x60 & ~x77 & ~x112 & ~x132 & ~x196 & ~x493 & ~x519 & ~x560 & ~x606 & ~x735;
assign c558 =  x692 &  x718 & ~x192 & ~x249 & ~x304 & ~x306 & ~x408 & ~x415 & ~x417 & ~x436 & ~x464 & ~x465 & ~x499 & ~x500 & ~x561 & ~x588;
assign c560 =  x348 &  x431 & ~x24 & ~x36 & ~x88 & ~x283 & ~x300 & ~x315 & ~x344 & ~x370 & ~x394 & ~x556 & ~x653 & ~x708;
assign c562 =  x301 &  x473 & ~x718;
assign c564 =  x568 &  x742 &  x744 & ~x359 & ~x410 & ~x735;
assign c566 = ~x3 & ~x32 & ~x47 & ~x79 & ~x80 & ~x83 & ~x114 & ~x142 & ~x144 & ~x191 & ~x201 & ~x223 & ~x249 & ~x251 & ~x256 & ~x283 & ~x296 & ~x298 & ~x335 & ~x336 & ~x339 & ~x341 & ~x353 & ~x358 & ~x364 & ~x379 & ~x381 & ~x394 & ~x407 & ~x409 & ~x411 & ~x415 & ~x438 & ~x442 & ~x469 & ~x470 & ~x555 & ~x584 & ~x673 & ~x675 & ~x705 & ~x732 & ~x781;
assign c568 = ~x3 & ~x20 & ~x21 & ~x23 & ~x47 & ~x48 & ~x49 & ~x51 & ~x52 & ~x54 & ~x55 & ~x60 & ~x75 & ~x76 & ~x78 & ~x81 & ~x84 & ~x88 & ~x107 & ~x109 & ~x111 & ~x116 & ~x134 & ~x137 & ~x140 & ~x164 & ~x166 & ~x171 & ~x195 & ~x219 & ~x220 & ~x222 & ~x247 & ~x248 & ~x284 & ~x285 & ~x305 & ~x339 & ~x342 & ~x354 & ~x357 & ~x360 & ~x364 & ~x366 & ~x380 & ~x381 & ~x384 & ~x387 & ~x394 & ~x396 & ~x411 & ~x416 & ~x421 & ~x423 & ~x440 & ~x442 & ~x443 & ~x444 & ~x451 & ~x452 & ~x471 & ~x474 & ~x479 & ~x500 & ~x503 & ~x505 & ~x507 & ~x528 & ~x531 & ~x533 & ~x535 & ~x562 & ~x586 & ~x589 & ~x592 & ~x617 & ~x619 & ~x647 & ~x670 & ~x675 & ~x681 & ~x682 & ~x683 & ~x696 & ~x732 & ~x736 & ~x753 & ~x758 & ~x759 & ~x761 & ~x764 & ~x765;
assign c570 =  x760 & ~x322 & ~x430 & ~x457;
assign c572 =  x0 &  x30;
assign c574 = ~x15 & ~x22 & ~x28 & ~x42 & ~x46 & ~x52 & ~x80 & ~x181 & ~x182 & ~x263 & ~x265 & ~x292 & ~x347 & ~x353 & ~x376 & ~x382 & ~x403 & ~x458 & ~x459 & ~x542 & ~x671 & ~x676 & ~x700 & ~x726 & ~x727 & ~x738 & ~x753;
assign c576 =  x460 &  x515 &  x745 & ~x174 & ~x231 & ~x329 & ~x381 & ~x385 & ~x409 & ~x435 & ~x440;
assign c578 =  x717 & ~x191 & ~x248 & ~x382 & ~x409 & ~x435 & ~x463 & ~x491 & ~x501 & ~x521 & ~x528;
assign c580 =  x307;
assign c582 =  x601 &  x745 & ~x55 & ~x138 & ~x165 & ~x194 & ~x248 & ~x249 & ~x437 & ~x465 & ~x492 & ~x527;
assign c584 =  x112;
assign c586 =  x699;
assign c588 =  x0 &  x759;
assign c590 =  x16 &  x757;
assign c592 =  x264 &  x319 & ~x186 & ~x222 & ~x242 & ~x299 & ~x328 & ~x384 & ~x451 & ~x600 & ~x622 & ~x625 & ~x666;
assign c594 =  x606 & ~x140 & ~x147 & ~x167 & ~x205 & ~x221 & ~x223 & ~x232 & ~x247 & ~x297 & ~x337 & ~x366 & ~x682;
assign c596 =  x515 &  x600 & ~x192 & ~x200 & ~x227 & ~x303 & ~x365 & ~x366 & ~x410 & ~x443 & ~x463 & ~x465 & ~x466 & ~x519;
assign c598 =  x154 &  x689 & ~x436 & ~x438;
assign c5100 =  x744 & ~x5 & ~x33 & ~x46 & ~x49 & ~x50 & ~x60 & ~x142 & ~x143 & ~x165 & ~x229 & ~x255 & ~x303 & ~x304 & ~x306 & ~x310 & ~x333 & ~x340 & ~x354 & ~x357 & ~x359 & ~x365 & ~x385 & ~x416 & ~x422 & ~x469 & ~x471 & ~x491 & ~x533 & ~x605 & ~x616 & ~x709 & ~x735 & ~x754;
assign c5102 =  x415 & ~x84 & ~x236 & ~x280 & ~x463 & ~x466 & ~x467 & ~x597 & ~x779;
assign c5104 = ~x5 & ~x20 & ~x22 & ~x31 & ~x59 & ~x75 & ~x80 & ~x84 & ~x107 & ~x113 & ~x130 & ~x138 & ~x158 & ~x225 & ~x254 & ~x336 & ~x365 & ~x394 & ~x409 & ~x420 & ~x476 & ~x514 & ~x542 & ~x543 & ~x570 & ~x572 & ~x600 & ~x628 & ~x641 & ~x642 & ~x655 & ~x670 & ~x696 & ~x700 & ~x757 & ~x759 & ~x760 & ~x762 & ~x775;
assign c5106 =  x127 &  x239 &  x773 & ~x439;
assign c5108 =  x657 &  x747 & ~x492 & ~x493;
assign c5110 = ~x119 & ~x150 & ~x280 & ~x292 & ~x465 & ~x595 & ~x634 & ~x661 & ~x712;
assign c5112 =  x372 & ~x78 & ~x337 & ~x350 & ~x381 & ~x405 & ~x433 & ~x450 & ~x464 & ~x465 & ~x467 & ~x489 & ~x494 & ~x518 & ~x758;
assign c5114 =  x245 &  x331 &  x475;
assign c5116 =  x228 &  x285 &  x302 &  x331 &  x342 & ~x489;
assign c5118 =  x431 &  x459 &  x513 & ~x34 & ~x65 & ~x80 & ~x90 & ~x92 & ~x139 & ~x521 & ~x533 & ~x616 & ~x709;
assign c5120 = ~x4 & ~x12 & ~x15 & ~x16 & ~x26 & ~x28 & ~x29 & ~x41 & ~x56 & ~x69 & ~x84 & ~x85 & ~x111 & ~x112 & ~x123 & ~x141 & ~x151 & ~x197 & ~x224 & ~x235 & ~x263 & ~x264 & ~x292 & ~x294 & ~x295 & ~x308 & ~x319 & ~x320 & ~x336 & ~x347 & ~x378 & ~x403 & ~x406 & ~x430 & ~x432 & ~x433 & ~x458 & ~x459 & ~x514 & ~x615 & ~x650 & ~x706 & ~x726 & ~x751 & ~x754 & ~x756 & ~x757 & ~x758 & ~x779;
assign c5122 =  x196;
assign c5124 = ~x1 & ~x27 & ~x29 & ~x30 & ~x51 & ~x61 & ~x85 & ~x89 & ~x136 & ~x158 & ~x197 & ~x215 & ~x217 & ~x244 & ~x297 & ~x302 & ~x327 & ~x380 & ~x383 & ~x393 & ~x397 & ~x446 & ~x449 & ~x535 & ~x588 & ~x600 & ~x627 & ~x654 & ~x667 & ~x680 & ~x699 & ~x705 & ~x753;
assign c5126 =  x531;
assign c5128 = ~x76 & ~x108 & ~x110 & ~x138 & ~x198 & ~x220 & ~x223 & ~x246 & ~x252 & ~x277 & ~x284 & ~x296 & ~x300 & ~x303 & ~x325 & ~x327 & ~x328 & ~x334 & ~x354 & ~x355 & ~x358 & ~x362 & ~x379 & ~x380 & ~x387 & ~x417 & ~x422 & ~x464 & ~x476 & ~x491 & ~x558 & ~x707 & ~x735;
assign c5130 = ~x57 & ~x186 & ~x241 & ~x251 & ~x273 & ~x309 & ~x352 & ~x353 & ~x381 & ~x393 & ~x409 & ~x410 & ~x415 & ~x436 & ~x528 & ~x650 & ~x655 & ~x678 & ~x707;
assign c5132 =  x348 &  x403 &  x457 & ~x20 & ~x34 & ~x54 & ~x55 & ~x92 & ~x106 & ~x287 & ~x425 & ~x507 & ~x534 & ~x652 & ~x697 & ~x708 & ~x759 & ~x762;
assign c5134 =  x84;
assign c5136 = ~x10 & ~x13 & ~x36 & ~x37 & ~x41 & ~x92 & ~x140 & ~x141 & ~x206 & ~x234 & ~x252 & ~x262 & ~x320 & ~x322 & ~x347 & ~x349 & ~x376 & ~x403 & ~x456 & ~x457 & ~x485 & ~x510 & ~x512 & ~x513 & ~x514 & ~x540 & ~x566 & ~x586 & ~x594 & ~x623 & ~x699 & ~x726 & ~x755;
assign c5138 =  x419 & ~x93 & ~x241 & ~x270 & ~x437;
assign c5140 =  x756;
assign c5142 = ~x151 & ~x234 & ~x324 & ~x325 & ~x721;
assign c5144 =  x472 &  x529 & ~x548 & ~x551 & ~x633 & ~x684;
assign c5146 = ~x1 & ~x10 & ~x23 & ~x30 & ~x52 & ~x54 & ~x55 & ~x77 & ~x79 & ~x81 & ~x83 & ~x105 & ~x108 & ~x116 & ~x117 & ~x139 & ~x162 & ~x167 & ~x194 & ~x196 & ~x255 & ~x309 & ~x310 & ~x325 & ~x339 & ~x352 & ~x354 & ~x364 & ~x365 & ~x368 & ~x381 & ~x395 & ~x422 & ~x449 & ~x465 & ~x466 & ~x467 & ~x497 & ~x525 & ~x589 & ~x654 & ~x681 & ~x708 & ~x754 & ~x759 & ~x760 & ~x761;
assign c5148 =  x426 &  x481 &  x536 & ~x50 & ~x436 & ~x438 & ~x487 & ~x488 & ~x493 & ~x518 & ~x547 & ~x572 & ~x678 & ~x680 & ~x707;
assign c5150 = ~x26 & ~x48 & ~x351 & ~x382 & ~x410 & ~x440 & ~x449 & ~x463 & ~x491 & ~x517 & ~x525 & ~x526 & ~x554 & ~x555 & ~x610 & ~x612 & ~x636 & ~x681 & ~x725 & ~x754 & ~x764;
assign c5152 =  x27 &  x420;
assign c5154 =  x386 &  x415 & ~x627 & ~x684;
assign c5156 =  x431 &  x459 &  x513 & ~x34 & ~x93 & ~x145 & ~x505 & ~x519 & ~x582 & ~x589 & ~x609 & ~x634 & ~x707;
assign c5158 =  x397 &  x417 & ~x65 & ~x380 & ~x541;
assign c5160 = ~x18 & ~x21 & ~x48 & ~x85 & ~x86 & ~x87 & ~x110 & ~x115 & ~x143 & ~x158 & ~x190 & ~x192 & ~x202 & ~x228 & ~x229 & ~x247 & ~x254 & ~x256 & ~x279 & ~x284 & ~x301 & ~x303 & ~x307 & ~x309 & ~x339 & ~x355 & ~x356 & ~x361 & ~x367 & ~x384 & ~x385 & ~x388 & ~x394 & ~x413 & ~x414 & ~x419 & ~x424 & ~x425 & ~x443 & ~x446 & ~x450 & ~x474 & ~x476 & ~x478 & ~x479 & ~x481 & ~x501 & ~x502 & ~x528 & ~x529 & ~x561 & ~x573 & ~x583 & ~x626 & ~x627 & ~x643 & ~x653 & ~x675 & ~x680 & ~x706 & ~x707 & ~x709 & ~x753 & ~x754 & ~x755;
assign c5162 =  x728;
assign c5164 = ~x10 & ~x28 & ~x84 & ~x139 & ~x168 & ~x177 & ~x179 & ~x209 & ~x213 & ~x234 & ~x353 & ~x407 & ~x485 & ~x595 & ~x621 & ~x648 & ~x671 & ~x679 & ~x680 & ~x691 & ~x697 & ~x705 & ~x732 & ~x754 & ~x778;
assign c5166 =  x26;
assign c5168 =  x756;
assign c5170 =  x303 &  x360 & ~x578;
assign c5172 =  x348 &  x375 &  x430 & ~x3 & ~x5 & ~x6 & ~x8 & ~x30 & ~x50 & ~x53 & ~x58 & ~x76 & ~x77 & ~x79 & ~x81 & ~x82 & ~x86 & ~x87 & ~x105 & ~x107 & ~x113 & ~x114 & ~x118 & ~x134 & ~x136 & ~x139 & ~x140 & ~x141 & ~x143 & ~x144 & ~x168 & ~x171 & ~x193 & ~x201 & ~x255 & ~x277 & ~x280 & ~x282 & ~x306 & ~x308 & ~x309 & ~x310 & ~x312 & ~x330 & ~x332 & ~x337 & ~x340 & ~x341 & ~x342 & ~x359 & ~x365 & ~x368 & ~x369 & ~x388 & ~x389 & ~x392 & ~x393 & ~x394 & ~x395 & ~x396 & ~x421 & ~x424 & ~x449 & ~x452 & ~x475 & ~x476 & ~x504 & ~x505 & ~x527 & ~x529 & ~x531 & ~x533 & ~x535 & ~x559 & ~x562 & ~x587 & ~x589 & ~x611 & ~x612 & ~x625 & ~x641 & ~x642 & ~x652 & ~x653 & ~x679 & ~x680 & ~x681 & ~x697 & ~x708 & ~x725 & ~x729 & ~x732 & ~x734 & ~x736 & ~x755 & ~x756 & ~x758 & ~x760 & ~x761 & ~x762 & ~x763 & ~x780 & ~x783;
assign c5174 =  x524 & ~x10 & ~x18 & ~x27 & ~x82 & ~x85 & ~x87 & ~x109 & ~x110 & ~x111 & ~x115 & ~x121 & ~x138 & ~x166 & ~x177 & ~x204 & ~x226 & ~x246 & ~x249 & ~x250 & ~x279 & ~x281 & ~x282 & ~x302 & ~x304 & ~x307 & ~x330 & ~x331 & ~x360 & ~x362 & ~x392 & ~x416 & ~x417 & ~x445 & ~x446 & ~x447 & ~x476 & ~x533 & ~x560 & ~x561 & ~x586 & ~x613 & ~x614 & ~x643 & ~x644 & ~x698 & ~x727;
assign c5176 =  x274 &  x302 &  x331 &  x388 & ~x69 & ~x325 & ~x381 & ~x487 & ~x489 & ~x680 & ~x720 & ~x748;
assign c5178 =  x0;
assign c5180 =  x375 & ~x19 & ~x87 & ~x107 & ~x136 & ~x197 & ~x224 & ~x242 & ~x259 & ~x272 & ~x299 & ~x362 & ~x384 & ~x393 & ~x413 & ~x416 & ~x449 & ~x452 & ~x564 & ~x567 & ~x585 & ~x598 & ~x622 & ~x625 & ~x648 & ~x654 & ~x666 & ~x733;
assign c5182 =  x773 & ~x81 & ~x107 & ~x173 & ~x360 & ~x380 & ~x385 & ~x411 & ~x412 & ~x418 & ~x419 & ~x443 & ~x548 & ~x761 & ~x782;
assign c5184 =  x374 & ~x3 & ~x24 & ~x31 & ~x84 & ~x309 & ~x324 & ~x325 & ~x367 & ~x381 & ~x392 & ~x395 & ~x421 & ~x437 & ~x450 & ~x467 & ~x493 & ~x615 & ~x624 & ~x643 & ~x764;
assign c5186 =  x496 &  x552 &  x580 & ~x18 & ~x57 & ~x68 & ~x137 & ~x141 & ~x165 & ~x166 & ~x197 & ~x222 & ~x225 & ~x253 & ~x278 & ~x309 & ~x346 & ~x347 & ~x348 & ~x358 & ~x374 & ~x389 & ~x390 & ~x402 & ~x431 & ~x445 & ~x458 & ~x472 & ~x476 & ~x502 & ~x727 & ~x739;
assign c5188 =  x27;
assign c5190 = ~x6 & ~x30 & ~x54 & ~x55 & ~x61 & ~x86 & ~x88 & ~x108 & ~x116 & ~x220 & ~x224 & ~x228 & ~x245 & ~x269 & ~x273 & ~x279 & ~x280 & ~x296 & ~x307 & ~x313 & ~x314 & ~x324 & ~x325 & ~x326 & ~x352 & ~x359 & ~x360 & ~x380 & ~x388 & ~x396 & ~x408 & ~x410 & ~x412 & ~x416 & ~x419 & ~x421 & ~x436 & ~x446 & ~x449 & ~x465 & ~x466 & ~x467 & ~x468 & ~x472 & ~x476 & ~x498 & ~x528 & ~x531 & ~x532 & ~x554 & ~x557 & ~x586 & ~x640 & ~x642 & ~x676 & ~x678 & ~x681 & ~x696 & ~x728 & ~x756;
assign c5192 =  x287 &  x315 &  x398 &  x453 & ~x41 & ~x96 & ~x321 & ~x351 & ~x403 & ~x458 & ~x567;
assign c5194 =  x472 &  x499 & ~x79 & ~x80 & ~x130 & ~x161 & ~x656 & ~x657 & ~x714 & ~x717;
assign c5196 =  x392;
assign c5198 = ~x18 & ~x23 & ~x33 & ~x60 & ~x81 & ~x106 & ~x183 & ~x225 & ~x364 & ~x486 & ~x514 & ~x592 & ~x624 & ~x643 & ~x678 & ~x683 & ~x684 & ~x715 & ~x733 & ~x743 & ~x753 & ~x755 & ~x759;
assign c5200 =  x263 &  x318 & ~x191 & ~x211 & ~x215 & ~x239 & ~x240 & ~x269 & ~x272 & ~x299 & ~x307 & ~x312 & ~x390 & ~x596 & ~x597 & ~x623 & ~x624 & ~x679 & ~x704 & ~x705;
assign c5202 =  x25 &  x447;
assign c5204 =  x319 & ~x144 & ~x225 & ~x270 & ~x295 & ~x323 & ~x353 & ~x354 & ~x366 & ~x367 & ~x383 & ~x506 & ~x557 & ~x653 & ~x681 & ~x700 & ~x706 & ~x733 & ~x736;
assign c5206 = ~x7 & ~x10 & ~x11 & ~x27 & ~x41 & ~x53 & ~x57 & ~x58 & ~x65 & ~x83 & ~x112 & ~x280 & ~x298 & ~x324 & ~x325 & ~x336 & ~x352 & ~x353 & ~x364 & ~x381 & ~x527 & ~x543 & ~x556 & ~x570 & ~x572 & ~x584 & ~x585 & ~x598 & ~x615 & ~x626 & ~x627 & ~x639 & ~x652 & ~x672 & ~x750 & ~x780 & ~x783;
assign c5208 =  x783;
assign c5210 = ~x30 & ~x91 & ~x109 & ~x161 & ~x165 & ~x171 & ~x186 & ~x190 & ~x192 & ~x213 & ~x214 & ~x216 & ~x220 & ~x229 & ~x244 & ~x272 & ~x360 & ~x363 & ~x398 & ~x505 & ~x532 & ~x573 & ~x598 & ~x616 & ~x624 & ~x626 & ~x627 & ~x644 & ~x651 & ~x678 & ~x681 & ~x704 & ~x705 & ~x731 & ~x762 & ~x781;
assign c5212 =  x26;
assign c5214 = ~x2 & ~x19 & ~x39 & ~x42 & ~x43 & ~x53 & ~x67 & ~x83 & ~x91 & ~x96 & ~x100 & ~x108 & ~x113 & ~x126 & ~x129 & ~x135 & ~x140 & ~x164 & ~x166 & ~x364 & ~x406 & ~x421 & ~x432 & ~x459 & ~x490 & ~x518 & ~x543 & ~x627 & ~x656 & ~x666 & ~x671 & ~x694 & ~x698 & ~x712 & ~x730 & ~x739 & ~x747;
assign c5216 = ~x0 & ~x27 & ~x48 & ~x50 & ~x56 & ~x83 & ~x393 & ~x404 & ~x405 & ~x432 & ~x459 & ~x460 & ~x516 & ~x518 & ~x583 & ~x585 & ~x612 & ~x638 & ~x655 & ~x667 & ~x669 & ~x686 & ~x696 & ~x704 & ~x723 & ~x728 & ~x730 & ~x732 & ~x758 & ~x770;
assign c5218 =  x386 &  x471 & ~x604 & ~x633;
assign c5220 =  x487 & ~x36 & ~x85 & ~x143 & ~x198 & ~x200 & ~x248 & ~x304 & ~x312 & ~x329 & ~x352 & ~x380 & ~x384 & ~x385 & ~x407 & ~x409 & ~x412 & ~x435 & ~x437 & ~x438 & ~x439 & ~x470 & ~x471 & ~x475 & ~x505 & ~x530 & ~x558 & ~x562;
assign c5222 =  x385 &  x443 &  x471 & ~x212 & ~x602 & ~x627;
assign c5224 =  x292 &  x405 & ~x65 & ~x93 & ~x120 & ~x134 & ~x143 & ~x162 & ~x172 & ~x175 & ~x227 & ~x277 & ~x287 & ~x315 & ~x330 & ~x331 & ~x333 & ~x337 & ~x371 & ~x397 & ~x423 & ~x449 & ~x589 & ~x654 & ~x655 & ~x708;
assign c5226 =  x0;
assign c5228 =  x388 &  x426 &  x481 & ~x461 & ~x653 & ~x712;
assign c5230 = ~x18 & ~x21 & ~x22 & ~x30 & ~x50 & ~x56 & ~x57 & ~x69 & ~x79 & ~x83 & ~x87 & ~x109 & ~x113 & ~x126 & ~x139 & ~x142 & ~x143 & ~x169 & ~x170 & ~x192 & ~x194 & ~x195 & ~x198 & ~x199 & ~x221 & ~x224 & ~x225 & ~x248 & ~x251 & ~x252 & ~x253 & ~x303 & ~x304 & ~x309 & ~x310 & ~x321 & ~x323 & ~x331 & ~x333 & ~x334 & ~x338 & ~x348 & ~x349 & ~x351 & ~x358 & ~x360 & ~x362 & ~x365 & ~x366 & ~x376 & ~x378 & ~x379 & ~x386 & ~x387 & ~x388 & ~x391 & ~x393 & ~x394 & ~x405 & ~x407 & ~x414 & ~x415 & ~x416 & ~x417 & ~x421 & ~x432 & ~x433 & ~x443 & ~x446 & ~x471 & ~x472 & ~x474 & ~x475 & ~x477 & ~x478 & ~x500 & ~x501 & ~x505 & ~x506 & ~x530 & ~x533 & ~x534 & ~x558 & ~x559 & ~x560 & ~x561 & ~x562 & ~x588 & ~x590 & ~x613 & ~x614 & ~x644 & ~x645 & ~x646 & ~x672 & ~x673 & ~x701 & ~x726 & ~x729 & ~x754 & ~x756 & ~x768;
assign c5232 =  x341 &  x369 &  x397 & ~x2 & ~x3 & ~x13 & ~x18 & ~x19 & ~x21 & ~x23 & ~x40 & ~x41 & ~x42 & ~x50 & ~x66 & ~x68 & ~x69 & ~x70 & ~x80 & ~x84 & ~x96 & ~x98 & ~x110 & ~x113 & ~x121 & ~x122 & ~x149 & ~x150 & ~x168 & ~x196 & ~x252 & ~x280 & ~x281 & ~x308 & ~x321 & ~x322 & ~x336 & ~x337 & ~x349 & ~x350 & ~x364 & ~x375 & ~x376 & ~x392 & ~x404 & ~x405 & ~x430 & ~x431 & ~x432 & ~x433 & ~x458 & ~x459 & ~x487 & ~x558 & ~x586 & ~x587 & ~x614 & ~x642 & ~x670 & ~x672 & ~x699 & ~x700 & ~x701 & ~x729 & ~x738 & ~x739 & ~x754 & ~x757 & ~x766 & ~x781 & ~x782;
assign c5234 = ~x50 & ~x114 & ~x140 & ~x196 & ~x197 & ~x219 & ~x223 & ~x277 & ~x278 & ~x282 & ~x326 & ~x334 & ~x352 & ~x360 & ~x362 & ~x364 & ~x407 & ~x412 & ~x413 & ~x438 & ~x440 & ~x443 & ~x467 & ~x469 & ~x471 & ~x476 & ~x492 & ~x506 & ~x616 & ~x644 & ~x728 & ~x734;
assign c5236 = ~x8 & ~x19 & ~x27 & ~x84 & ~x85 & ~x104 & ~x144 & ~x158 & ~x186 & ~x188 & ~x191 & ~x196 & ~x229 & ~x244 & ~x300 & ~x362 & ~x386 & ~x389 & ~x544 & ~x598 & ~x647 & ~x648 & ~x650 & ~x655 & ~x670 & ~x675 & ~x680 & ~x683 & ~x696 & ~x700 & ~x726 & ~x754;
assign c5238 = ~x54 & ~x421 & ~x438 & ~x600 & ~x603 & ~x610 & ~x630 & ~x661 & ~x665 & ~x684;
assign c5240 =  x425 &  x453 &  x480 & ~x293 & ~x377 & ~x431 & ~x486 & ~x514 & ~x541 & ~x596 & ~x597 & ~x650;
assign c5242 =  x531;
assign c5244 = ~x23 & ~x28 & ~x52 & ~x86 & ~x144 & ~x165 & ~x201 & ~x218 & ~x228 & ~x253 & ~x271 & ~x274 & ~x277 & ~x285 & ~x305 & ~x311 & ~x324 & ~x332 & ~x354 & ~x359 & ~x360 & ~x381 & ~x389 & ~x391 & ~x412 & ~x419 & ~x437 & ~x438 & ~x465 & ~x529 & ~x555 & ~x557 & ~x558 & ~x583 & ~x590 & ~x645 & ~x682 & ~x698 & ~x699 & ~x706 & ~x709 & ~x734 & ~x735 & ~x758 & ~x763;
assign c5248 =  x500 & ~x107 & ~x110 & ~x521 & ~x547 & ~x606 & ~x631 & ~x688 & ~x689 & ~x747 & ~x767 & ~x769;
assign c5250 = ~x52 & ~x134 & ~x173 & ~x190 & ~x200 & ~x239 & ~x304 & ~x332 & ~x361 & ~x363 & ~x364 & ~x380 & ~x418 & ~x561 & ~x564 & ~x570 & ~x597 & ~x616 & ~x619 & ~x620 & ~x624 & ~x653 & ~x655 & ~x680 & ~x683 & ~x708;
assign c5252 = ~x17 & ~x23 & ~x83 & ~x91 & ~x93 & ~x236 & ~x263 & ~x291 & ~x346 & ~x347 & ~x354 & ~x376 & ~x402 & ~x538 & ~x650 & ~x736;
assign c5254 =  x425 & ~x152 & ~x364 & ~x375 & ~x376 & ~x458 & ~x514;
assign c5256 =  x256 &  x285 &  x315 &  x342 & ~x522 & ~x631;
assign c5258 =  x783;
assign c5260 =  x27;
assign c5262 = ~x11 & ~x65 & ~x68 & ~x154 & ~x184 & ~x225 & ~x235 & ~x263 & ~x319 & ~x376 & ~x403 & ~x431 & ~x432 & ~x458 & ~x459 & ~x513 & ~x515 & ~x540 & ~x541 & ~x566 & ~x649 & ~x650 & ~x725 & ~x726 & ~x744 & ~x773;
assign c5264 =  x1;
assign c5266 =  x168;
assign c5268 =  x347 &  x430 &  x485 & ~x33 & ~x296 & ~x299 & ~x325 & ~x330 & ~x423 & ~x610 & ~x704 & ~x705;
assign c5270 =  x531;
assign c5272 = ~x65 & ~x66 & ~x100 & ~x124 & ~x292 & ~x318 & ~x320 & ~x373 & ~x402 & ~x430 & ~x566 & ~x620 & ~x623 & ~x693 & ~x721 & ~x769;
assign c5274 =  x284 &  x340 & ~x9 & ~x37 & ~x38 & ~x93 & ~x212 & ~x292 & ~x294 & ~x297 & ~x319 & ~x375 & ~x429 & ~x430 & ~x431 & ~x488 & ~x514 & ~x543;
assign c5276 =  x286 &  x371 & ~x177 & ~x410 & ~x433 & ~x517 & ~x734;
assign c5278 =  x414 &  x472 &  x500 & ~x658 & ~x687 & ~x714 & ~x718;
assign c5280 = ~x33 & ~x135 & ~x142 & ~x270 & ~x271 & ~x296 & ~x310 & ~x322 & ~x323 & ~x351 & ~x352 & ~x357 & ~x383 & ~x394 & ~x438 & ~x449 & ~x498 & ~x527 & ~x650 & ~x733 & ~x751;
assign c5282 =  x746 &  x747 &  x775 & ~x49 & ~x59 & ~x61 & ~x139 & ~x221 & ~x249 & ~x275 & ~x277 & ~x342 & ~x357 & ~x367 & ~x558 & ~x738;
assign c5284 = ~x2 & ~x86 & ~x94 & ~x95 & ~x207 & ~x236 & ~x264 & ~x267 & ~x320 & ~x322 & ~x325 & ~x405 & ~x459 & ~x460 & ~x544 & ~x598 & ~x599 & ~x600 & ~x615 & ~x624 & ~x626 & ~x650 & ~x651 & ~x697 & ~x723;
assign c5286 =  x26;
assign c5288 =  x384 &  x471 & ~x656 & ~x686 & ~x744;
assign c5290 =  x745 & ~x47 & ~x79 & ~x163 & ~x164 & ~x189 & ~x194 & ~x227 & ~x249 & ~x274 & ~x275 & ~x302 & ~x326 & ~x328 & ~x333 & ~x334 & ~x358 & ~x360 & ~x367 & ~x368 & ~x475 & ~x491 & ~x529 & ~x557 & ~x560 & ~x734;
assign c5292 =  x414 &  x442 &  x499 & ~x107 & ~x657 & ~x661 & ~x662 & ~x719;
assign c5294 = ~x19 & ~x22 & ~x77 & ~x79 & ~x83 & ~x106 & ~x466 & ~x550 & ~x588 & ~x602 & ~x632 & ~x637 & ~x654 & ~x656 & ~x690 & ~x715 & ~x748 & ~x750 & ~x776;
assign c5296 = ~x133 & ~x135 & ~x239 & ~x268 & ~x279 & ~x324 & ~x326 & ~x363 & ~x382 & ~x384 & ~x440 & ~x447 & ~x584 & ~x627 & ~x679 & ~x703;
assign c5298 =  x223 &  x392;
assign c5300 = ~x6 & ~x35 & ~x62 & ~x64 & ~x93 & ~x128 & ~x149 & ~x156 & ~x159 & ~x197 & ~x239 & ~x364 & ~x543 & ~x570 & ~x571 & ~x597 & ~x642 & ~x646 & ~x647 & ~x648 & ~x664 & ~x666 & ~x678 & ~x730 & ~x749 & ~x752 & ~x783;
assign c5302 =  x188 &  x275 &  x447;
assign c5304 =  x212 &  x237 &  x266 & ~x361 & ~x398 & ~x439 & ~x500 & ~x521;
assign c5306 =  x265 &  x292 &  x540 & ~x370 & ~x372;
assign c5308 = ~x10 & ~x12 & ~x23 & ~x42 & ~x55 & ~x111 & ~x112 & ~x140 & ~x168 & ~x169 & ~x179 & ~x180 & ~x197 & ~x207 & ~x208 & ~x209 & ~x237 & ~x265 & ~x292 & ~x293 & ~x319 & ~x323 & ~x374 & ~x375 & ~x402 & ~x403 & ~x458 & ~x459 & ~x487 & ~x593 & ~x650 & ~x679 & ~x699 & ~x706 & ~x733 & ~x755 & ~x772;
assign c5310 =  x212 &  x515 & ~x408 & ~x439 & ~x470 & ~x497 & ~x520;
assign c5314 = ~x105 & ~x106 & ~x110 & ~x141 & ~x161 & ~x163 & ~x200 & ~x216 & ~x219 & ~x221 & ~x223 & ~x225 & ~x247 & ~x252 & ~x274 & ~x277 & ~x302 & ~x305 & ~x306 & ~x328 & ~x332 & ~x334 & ~x352 & ~x353 & ~x366 & ~x382 & ~x411 & ~x414 & ~x436 & ~x439 & ~x440 & ~x466 & ~x469 & ~x476 & ~x556 & ~x613 & ~x696 & ~x702 & ~x708 & ~x760 & ~x761 & ~x781;
assign c5316 =  x633 & ~x115 & ~x160 & ~x213 & ~x241 & ~x242 & ~x254 & ~x297 & ~x326 & ~x382 & ~x417 & ~x703;
assign c5318 =  x266 &  x292 &  x404 &  x460 &  x567;
assign c5320 = ~x25 & ~x29 & ~x30 & ~x55 & ~x83 & ~x84 & ~x85 & ~x86 & ~x113 & ~x212 & ~x223 & ~x267 & ~x280 & ~x296 & ~x322 & ~x323 & ~x325 & ~x352 & ~x354 & ~x381 & ~x382 & ~x422 & ~x499 & ~x504 & ~x531 & ~x557 & ~x596 & ~x597 & ~x614 & ~x615 & ~x625 & ~x643 & ~x680 & ~x694 & ~x722 & ~x727 & ~x751 & ~x753 & ~x754 & ~x757 & ~x761 & ~x780;
assign c5322 =  x376 & ~x4 & ~x47 & ~x58 & ~x86 & ~x106 & ~x115 & ~x137 & ~x200 & ~x222 & ~x226 & ~x230 & ~x256 & ~x288 & ~x301 & ~x303 & ~x328 & ~x357 & ~x363 & ~x387 & ~x392 & ~x398 & ~x419 & ~x469 & ~x474 & ~x509 & ~x536 & ~x598 & ~x617 & ~x645 & ~x653 & ~x654 & ~x675 & ~x736 & ~x755 & ~x778;
assign c5324 =  x479 & ~x16 & ~x42 & ~x111 & ~x147 & ~x149 & ~x175 & ~x204 & ~x205 & ~x263 & ~x349 & ~x351 & ~x352 & ~x353 & ~x374 & ~x376 & ~x429;
assign c5326 = ~x50 & ~x57 & ~x83 & ~x107 & ~x114 & ~x161 & ~x190 & ~x198 & ~x225 & ~x227 & ~x250 & ~x266 & ~x268 & ~x270 & ~x272 & ~x283 & ~x298 & ~x308 & ~x313 & ~x327 & ~x340 & ~x354 & ~x357 & ~x414 & ~x555 & ~x556 & ~x652 & ~x675 & ~x679 & ~x729 & ~x734 & ~x735 & ~x782 & ~x783;
assign c5328 =  x1 &  x3;
assign c5330 =  x563 & ~x9 & ~x11 & ~x36 & ~x52 & ~x65 & ~x97 & ~x176 & ~x178 & ~x353 & ~x377 & ~x379 & ~x404 & ~x405 & ~x406 & ~x433 & ~x434 & ~x487 & ~x671 & ~x680;
assign c5332 = ~x2 & ~x3 & ~x17 & ~x18 & ~x28 & ~x35 & ~x38 & ~x45 & ~x49 & ~x50 & ~x119 & ~x148 & ~x177 & ~x206 & ~x280 & ~x365 & ~x436 & ~x437 & ~x466 & ~x494 & ~x569 & ~x598 & ~x600 & ~x627 & ~x644 & ~x666 & ~x694 & ~x712 & ~x762 & ~x777 & ~x782;
assign c5334 =  x746 &  x747 & ~x18 & ~x135 & ~x192 & ~x219 & ~x333 & ~x389 & ~x408 & ~x437 & ~x492 & ~x493;
assign c5336 = ~x0 & ~x22 & ~x30 & ~x68 & ~x80 & ~x85 & ~x143 & ~x169 & ~x171 & ~x199 & ~x255 & ~x282 & ~x292 & ~x295 & ~x320 & ~x321 & ~x338 & ~x346 & ~x348 & ~x375 & ~x402 & ~x403 & ~x404 & ~x430 & ~x431 & ~x432 & ~x458 & ~x505 & ~x506 & ~x507 & ~x532 & ~x533 & ~x561 & ~x642 & ~x670 & ~x672 & ~x701 & ~x712 & ~x739 & ~x741 & ~x754;
assign c5338 =  x341 & ~x3 & ~x22 & ~x47 & ~x50 & ~x53 & ~x72 & ~x233 & ~x392 & ~x406 & ~x434 & ~x438 & ~x488 & ~x542 & ~x599 & ~x629 & ~x714 & ~x729 & ~x741 & ~x762 & ~x768 & ~x769;
assign c5340 =  x246 &  x419;
assign c5342 = ~x2 & ~x6 & ~x23 & ~x46 & ~x58 & ~x80 & ~x169 & ~x229 & ~x239 & ~x265 & ~x269 & ~x286 & ~x295 & ~x322 & ~x326 & ~x379 & ~x380 & ~x437 & ~x670;
assign c5344 =  x237 &  x293 &  x431 & ~x230 & ~x283 & ~x373 & ~x653 & ~x680;
assign c5346 =  x357 &  x472 & ~x630 & ~x686 & ~x688 & ~x714;
assign c5348 =  x302 &  x331 & ~x497 & ~x636 & ~x690 & ~x693;
assign c5350 =  x460 &  x659 &  x687 &  x746 & ~x249 & ~x328;
assign c5352 =  x662 & ~x2 & ~x84 & ~x110 & ~x111 & ~x139 & ~x165 & ~x194 & ~x197 & ~x280 & ~x296 & ~x304 & ~x305 & ~x307 & ~x308 & ~x324 & ~x325 & ~x326 & ~x331 & ~x333 & ~x334 & ~x352 & ~x361 & ~x382 & ~x392 & ~x409 & ~x416 & ~x417 & ~x418 & ~x446 & ~x448 & ~x500 & ~x557 & ~x558 & ~x754;
assign c5354 =  x224;
assign c5356 =  x347 &  x429 &  x430 &  x456 & ~x3 & ~x5 & ~x109 & ~x138 & ~x139 & ~x421 & ~x422 & ~x477 & ~x479 & ~x533 & ~x560 & ~x561 & ~x608 & ~x609 & ~x664 & ~x692 & ~x756 & ~x777 & ~x782;
assign c5358 =  x348 &  x405 & ~x7 & ~x35 & ~x187 & ~x194 & ~x200 & ~x216 & ~x218 & ~x285 & ~x334 & ~x342 & ~x395 & ~x422 & ~x426 & ~x507 & ~x584 & ~x599 & ~x680 & ~x736;
assign c5360 =  x432 &  x686 &  x743 &  x772 & ~x120 & ~x201 & ~x372;
assign c5362 =  x27;
assign c5364 =  x451 & ~x23 & ~x120 & ~x121 & ~x209 & ~x320 & ~x376 & ~x404 & ~x431 & ~x457 & ~x512 & ~x538 & ~x541 & ~x568 & ~x569;
assign c5366 =  x188 & ~x2 & ~x22 & ~x26 & ~x43 & ~x80 & ~x112 & ~x113 & ~x165 & ~x167 & ~x224 & ~x280 & ~x293 & ~x294 & ~x319 & ~x320 & ~x323 & ~x324 & ~x337 & ~x349 & ~x350 & ~x365 & ~x378 & ~x401 & ~x402 & ~x430 & ~x458 & ~x529 & ~x531 & ~x614 & ~x711 & ~x741;
assign c5368 =  x550 & ~x42 & ~x56 & ~x69 & ~x70 & ~x112 & ~x252 & ~x253 & ~x280 & ~x281 & ~x292 & ~x293 & ~x320 & ~x321 & ~x322 & ~x323 & ~x324 & ~x347 & ~x348 & ~x349 & ~x350 & ~x351 & ~x375 & ~x376 & ~x377 & ~x378 & ~x379 & ~x380 & ~x402 & ~x403 & ~x405 & ~x406 & ~x407 & ~x431 & ~x432 & ~x457 & ~x458 & ~x459 & ~x485 & ~x513 & ~x530 & ~x558 & ~x559 & ~x587 & ~x778;
assign c5370 = ~x1 & ~x20 & ~x27 & ~x48 & ~x49 & ~x80 & ~x81 & ~x84 & ~x86 & ~x88 & ~x106 & ~x110 & ~x137 & ~x167 & ~x170 & ~x194 & ~x195 & ~x197 & ~x199 & ~x220 & ~x226 & ~x249 & ~x282 & ~x283 & ~x296 & ~x297 & ~x303 & ~x305 & ~x308 & ~x313 & ~x324 & ~x330 & ~x331 & ~x332 & ~x334 & ~x335 & ~x340 & ~x353 & ~x357 & ~x360 & ~x364 & ~x385 & ~x391 & ~x393 & ~x395 & ~x409 & ~x420 & ~x421 & ~x437 & ~x446 & ~x450 & ~x470 & ~x500 & ~x503 & ~x506 & ~x507 & ~x528 & ~x532 & ~x534 & ~x535 & ~x556 & ~x562 & ~x586 & ~x588 & ~x590 & ~x614 & ~x615 & ~x655 & ~x672 & ~x682 & ~x683 & ~x710 & ~x728 & ~x735 & ~x754 & ~x757;
assign c5372 =  x302 & ~x497 & ~x524 & ~x581 & ~x667 & ~x721 & ~x723;
assign c5374 = ~x11 & ~x16 & ~x18 & ~x22 & ~x43 & ~x44 & ~x46 & ~x47 & ~x53 & ~x54 & ~x68 & ~x79 & ~x81 & ~x83 & ~x109 & ~x110 & ~x121 & ~x167 & ~x318 & ~x337 & ~x348 & ~x349 & ~x364 & ~x374 & ~x402 & ~x404 & ~x405 & ~x430 & ~x432 & ~x458 & ~x512 & ~x540 & ~x622 & ~x651 & ~x670 & ~x679 & ~x720 & ~x729 & ~x783;
assign c5376 = ~x11 & ~x13 & ~x23 & ~x24 & ~x29 & ~x40 & ~x68 & ~x86 & ~x110 & ~x111 & ~x139 & ~x225 & ~x235 & ~x262 & ~x291 & ~x292 & ~x294 & ~x296 & ~x317 & ~x318 & ~x320 & ~x323 & ~x324 & ~x345 & ~x346 & ~x352 & ~x400 & ~x401 & ~x402 & ~x404 & ~x428 & ~x429 & ~x431 & ~x456 & ~x458 & ~x484 & ~x503 & ~x531 & ~x540 & ~x560 & ~x588 & ~x671 & ~x698 & ~x711 & ~x727 & ~x768;
assign c5378 =  x756;
assign c5380 =  x285 & ~x11 & ~x210 & ~x211 & ~x347 & ~x375 & ~x377 & ~x403 & ~x459 & ~x486 & ~x564 & ~x587;
assign c5382 =  x112;
assign c5384 =  x1;
assign c5386 =  x370 & ~x0 & ~x17 & ~x21 & ~x27 & ~x41 & ~x42 & ~x43 & ~x44 & ~x49 & ~x69 & ~x124 & ~x125 & ~x309 & ~x336 & ~x337 & ~x350 & ~x375 & ~x376 & ~x379 & ~x403 & ~x407 & ~x430 & ~x458 & ~x459 & ~x476 & ~x485 & ~x540 & ~x567 & ~x643 & ~x729 & ~x782;
assign c5388 = ~x9 & ~x11 & ~x24 & ~x69 & ~x208 & ~x225 & ~x237 & ~x238 & ~x267 & ~x281 & ~x292 & ~x297 & ~x318 & ~x336 & ~x375 & ~x430 & ~x514 & ~x539 & ~x541 & ~x566 & ~x621 & ~x695 & ~x734 & ~x752;
assign c5390 =  x487 &  x541 &  x713 & ~x372 & ~x708 & ~x763;
assign c5392 =  x593 &  x662 & ~x51 & ~x110 & ~x137 & ~x198 & ~x199 & ~x220 & ~x249 & ~x250 & ~x255 & ~x283 & ~x304 & ~x311 & ~x332 & ~x359 & ~x379 & ~x386 & ~x387 & ~x390 & ~x394 & ~x407 & ~x419 & ~x421 & ~x443 & ~x445 & ~x471 & ~x472 & ~x500 & ~x505 & ~x701;
assign c5394 =  x755;
assign c5396 =  x217 & ~x495 & ~x498 & ~x527 & ~x528 & ~x549 & ~x555;
assign c5398 = ~x1 & ~x23 & ~x29 & ~x41 & ~x42 & ~x65 & ~x84 & ~x93 & ~x122 & ~x196 & ~x253 & ~x263 & ~x293 & ~x348 & ~x349 & ~x374 & ~x376 & ~x401 & ~x402 & ~x403 & ~x457 & ~x458 & ~x539 & ~x540 & ~x569 & ~x623 & ~x644 & ~x650 & ~x699 & ~x728 & ~x735 & ~x741 & ~x753 & ~x769 & ~x773 & ~x782;
assign c5400 =  x629 &  x720 & ~x493;
assign c5402 =  x443 &  x472 & ~x129 & ~x160 & ~x661 & ~x686 & ~x687 & ~x738 & ~x740 & ~x741 & ~x743;
assign c5404 = ~x11 & ~x29 & ~x54 & ~x85 & ~x111 & ~x168 & ~x181 & ~x209 & ~x236 & ~x237 & ~x238 & ~x263 & ~x264 & ~x266 & ~x291 & ~x319 & ~x375 & ~x376 & ~x377 & ~x378 & ~x403 & ~x405 & ~x430 & ~x432 & ~x434 & ~x459 & ~x486 & ~x487 & ~x514 & ~x538 & ~x592 & ~x594 & ~x595 & ~x620 & ~x623 & ~x649 & ~x731 & ~x735 & ~x753 & ~x754 & ~x762 & ~x783;
assign c5406 =  x387 &  x416 &  x445 & ~x518 & ~x694 & ~x740;
assign c5408 =  x196 &  x279;
assign c5410 =  x127 & ~x3 & ~x112 & ~x138 & ~x194 & ~x297 & ~x309 & ~x325 & ~x327 & ~x352 & ~x356 & ~x360 & ~x382 & ~x384 & ~x409 & ~x411 & ~x415 & ~x418 & ~x437 & ~x445 & ~x465 & ~x471 & ~x496 & ~x558 & ~x587 & ~x615 & ~x616 & ~x644 & ~x648 & ~x698 & ~x706 & ~x782;
assign c5412 = ~x8 & ~x21 & ~x24 & ~x33 & ~x83 & ~x103 & ~x135 & ~x143 & ~x159 & ~x162 & ~x167 & ~x169 & ~x171 & ~x174 & ~x199 & ~x232 & ~x249 & ~x277 & ~x299 & ~x308 & ~x309 & ~x384 & ~x391 & ~x419 & ~x448 & ~x452 & ~x479 & ~x559 & ~x561 & ~x571 & ~x587 & ~x617 & ~x624 & ~x627 & ~x649 & ~x654 & ~x668 & ~x672 & ~x677 & ~x679 & ~x683 & ~x695 & ~x696 & ~x708 & ~x722 & ~x730 & ~x754;
assign c5414 =  x361 &  x390 & ~x149 & ~x240 & ~x324 & ~x348 & ~x376 & ~x486;
assign c5416 =  x55;
assign c5418 =  x264 &  x348 & ~x49 & ~x63 & ~x115 & ~x133 & ~x143 & ~x164 & ~x243 & ~x255 & ~x257 & ~x258 & ~x287 & ~x364 & ~x398 & ~x448 & ~x481 & ~x529 & ~x591 & ~x626 & ~x680 & ~x735 & ~x759;
assign c5420 =  x140;
assign c5422 =  x643;
assign c5424 =  x291 &  x319 & ~x18 & ~x19 & ~x54 & ~x55 & ~x60 & ~x105 & ~x107 & ~x130 & ~x135 & ~x160 & ~x162 & ~x168 & ~x173 & ~x189 & ~x214 & ~x215 & ~x227 & ~x252 & ~x255 & ~x258 & ~x273 & ~x279 & ~x280 & ~x282 & ~x306 & ~x309 & ~x310 & ~x311 & ~x338 & ~x341 & ~x342 & ~x358 & ~x359 & ~x364 & ~x391 & ~x392 & ~x394 & ~x420 & ~x422 & ~x445 & ~x474 & ~x504 & ~x535 & ~x562 & ~x571 & ~x583 & ~x585 & ~x597 & ~x598 & ~x617 & ~x638 & ~x639 & ~x671 & ~x679 & ~x680 & ~x697 & ~x723 & ~x724 & ~x733 & ~x758 & ~x760 & ~x763 & ~x780;
assign c5426 =  x0;
assign c5428 = ~x1 & ~x2 & ~x25 & ~x28 & ~x30 & ~x31 & ~x38 & ~x54 & ~x57 & ~x66 & ~x81 & ~x82 & ~x84 & ~x94 & ~x95 & ~x108 & ~x109 & ~x112 & ~x113 & ~x123 & ~x139 & ~x140 & ~x142 & ~x144 & ~x150 & ~x165 & ~x170 & ~x171 & ~x192 & ~x195 & ~x196 & ~x199 & ~x219 & ~x224 & ~x226 & ~x249 & ~x250 & ~x251 & ~x252 & ~x254 & ~x255 & ~x275 & ~x276 & ~x279 & ~x280 & ~x301 & ~x302 & ~x305 & ~x308 & ~x309 & ~x310 & ~x330 & ~x332 & ~x338 & ~x345 & ~x358 & ~x360 & ~x361 & ~x362 & ~x363 & ~x374 & ~x386 & ~x389 & ~x390 & ~x392 & ~x400 & ~x414 & ~x416 & ~x417 & ~x444 & ~x445 & ~x449 & ~x472 & ~x475 & ~x477 & ~x478 & ~x500 & ~x502 & ~x503 & ~x505 & ~x506 & ~x529 & ~x530 & ~x531 & ~x533 & ~x534 & ~x557 & ~x558 & ~x561 & ~x585 & ~x586 & ~x590 & ~x614 & ~x615 & ~x616 & ~x645 & ~x670 & ~x681 & ~x728 & ~x735 & ~x737 & ~x756 & ~x763 & ~x764 & ~x765 & ~x783;
assign c5430 = ~x11 & ~x41 & ~x81 & ~x83 & ~x96 & ~x99 & ~x141 & ~x225 & ~x235 & ~x266 & ~x323 & ~x376 & ~x431 & ~x435 & ~x458 & ~x485 & ~x513 & ~x593 & ~x723 & ~x755 & ~x781 & ~x782;
assign c5432 =  x240 &  x265 & ~x361 & ~x409 & ~x412 & ~x521;
assign c5434 = ~x4 & ~x52 & ~x88 & ~x109 & ~x322 & ~x337 & ~x348 & ~x349 & ~x350 & ~x376 & ~x377 & ~x394 & ~x403 & ~x404 & ~x407 & ~x477 & ~x507 & ~x534 & ~x562 & ~x613 & ~x616 & ~x617 & ~x642 & ~x645 & ~x646 & ~x669 & ~x673 & ~x710 & ~x711 & ~x712 & ~x740 & ~x746 & ~x754 & ~x766 & ~x767 & ~x768 & ~x769 & ~x771 & ~x772 & ~x775;
assign c5436 =  x348 &  x376 &  x403 & ~x38 & ~x48 & ~x49 & ~x53 & ~x57 & ~x61 & ~x85 & ~x90 & ~x114 & ~x117 & ~x167 & ~x218 & ~x242 & ~x249 & ~x252 & ~x280 & ~x313 & ~x339 & ~x342 & ~x366 & ~x389 & ~x391 & ~x449 & ~x474 & ~x478 & ~x626 & ~x652 & ~x666 & ~x668 & ~x676 & ~x678 & ~x681 & ~x696 & ~x708 & ~x781;
assign c5438 =  x719 & ~x0 & ~x6 & ~x17 & ~x46 & ~x53 & ~x58 & ~x108 & ~x110 & ~x113 & ~x141 & ~x193 & ~x277 & ~x305 & ~x332 & ~x333 & ~x336 & ~x359 & ~x364 & ~x393 & ~x408 & ~x436 & ~x437 & ~x446 & ~x465 & ~x471 & ~x474 & ~x492 & ~x493 & ~x527;
assign c5440 = ~x16 & ~x17 & ~x23 & ~x25 & ~x28 & ~x53 & ~x56 & ~x58 & ~x67 & ~x84 & ~x95 & ~x96 & ~x112 & ~x122 & ~x177 & ~x224 & ~x225 & ~x281 & ~x317 & ~x345 & ~x401 & ~x429 & ~x458 & ~x485 & ~x513 & ~x531 & ~x540 & ~x643 & ~x671 & ~x680 & ~x682 & ~x693 & ~x707 & ~x708 & ~x710 & ~x723 & ~x739 & ~x753 & ~x757 & ~x764 & ~x767 & ~x768 & ~x782;
assign c5442 =  x140;
assign c5444 =  x266 &  x514 & ~x95 & ~x122 & ~x506;
assign c5446 = ~x20 & ~x31 & ~x46 & ~x58 & ~x63 & ~x110 & ~x129 & ~x139 & ~x178 & ~x179 & ~x183 & ~x210 & ~x211 & ~x234 & ~x543 & ~x572 & ~x627 & ~x654 & ~x657 & ~x678 & ~x684 & ~x722 & ~x767 & ~x777;
assign c5448 = ~x56 & ~x66 & ~x93 & ~x97 & ~x122 & ~x123 & ~x125 & ~x149 & ~x151 & ~x263 & ~x293 & ~x323 & ~x348 & ~x379 & ~x381 & ~x403 & ~x405 & ~x458 & ~x460 & ~x515 & ~x668 & ~x722 & ~x757;
assign c5450 =  x744 & ~x18 & ~x25 & ~x47 & ~x48 & ~x50 & ~x59 & ~x90 & ~x95 & ~x110 & ~x112 & ~x123 & ~x141 & ~x162 & ~x225 & ~x254 & ~x277 & ~x300 & ~x309 & ~x334 & ~x338 & ~x361 & ~x363 & ~x370 & ~x371 & ~x384 & ~x385 & ~x399 & ~x412 & ~x422 & ~x445 & ~x477 & ~x482 & ~x502 & ~x532 & ~x700 & ~x728 & ~x730 & ~x733 & ~x735;
assign c5452 =  x460 &  x486 & ~x17 & ~x142 & ~x174 & ~x202 & ~x219 & ~x329 & ~x343 & ~x372 & ~x398 & ~x399 & ~x584 & ~x585 & ~x588 & ~x681 & ~x738;
assign c5454 =  x388 & ~x50 & ~x233 & ~x380 & ~x436 & ~x466 & ~x520 & ~x570 & ~x686 & ~x742 & ~x747;
assign c5456 =  x749 & ~x409 & ~x438;
assign c5458 =  x455 & ~x8 & ~x19 & ~x21 & ~x24 & ~x26 & ~x48 & ~x79 & ~x110 & ~x392 & ~x492 & ~x518 & ~x521 & ~x533 & ~x680 & ~x681 & ~x708 & ~x709 & ~x763 & ~x768 & ~x769 & ~x779;
assign c5460 =  x274 & ~x29 & ~x392 & ~x497 & ~x552 & ~x579 & ~x582 & ~x583 & ~x608 & ~x611 & ~x632 & ~x633 & ~x636 & ~x637 & ~x694 & ~x722 & ~x746 & ~x748 & ~x751 & ~x752 & ~x773;
assign c5462 = ~x0 & ~x4 & ~x12 & ~x14 & ~x15 & ~x24 & ~x27 & ~x28 & ~x29 & ~x38 & ~x41 & ~x43 & ~x44 & ~x51 & ~x52 & ~x54 & ~x56 & ~x66 & ~x68 & ~x79 & ~x80 & ~x82 & ~x85 & ~x97 & ~x98 & ~x109 & ~x122 & ~x123 & ~x124 & ~x125 & ~x139 & ~x140 & ~x141 & ~x150 & ~x168 & ~x195 & ~x196 & ~x224 & ~x252 & ~x253 & ~x281 & ~x295 & ~x309 & ~x320 & ~x321 & ~x322 & ~x324 & ~x337 & ~x349 & ~x364 & ~x376 & ~x380 & ~x392 & ~x404 & ~x406 & ~x420 & ~x431 & ~x432 & ~x434 & ~x531 & ~x558 & ~x559 & ~x586 & ~x615 & ~x616 & ~x642 & ~x643 & ~x644 & ~x683 & ~x699 & ~x726 & ~x728 & ~x729 & ~x756 & ~x767 & ~x782 & ~x783;
assign c5464 =  x460 &  x688 & ~x105 & ~x195 & ~x231 & ~x245 & ~x258 & ~x297 & ~x304 & ~x331 & ~x353 & ~x361 & ~x370 & ~x533;
assign c5466 =  x223;
assign c5468 = ~x84 & ~x135 & ~x251 & ~x296 & ~x301 & ~x313 & ~x322 & ~x325 & ~x351 & ~x387 & ~x408 & ~x414 & ~x437 & ~x465 & ~x470 & ~x474 & ~x502 & ~x528 & ~x554 & ~x555;
assign c5470 =  x376 & ~x23 & ~x51 & ~x60 & ~x61 & ~x76 & ~x84 & ~x137 & ~x141 & ~x163 & ~x196 & ~x222 & ~x256 & ~x283 & ~x355 & ~x356 & ~x359 & ~x368 & ~x370 & ~x371 & ~x413 & ~x444 & ~x448 & ~x450 & ~x476 & ~x477 & ~x505 & ~x506 & ~x508 & ~x528 & ~x556 & ~x583 & ~x619 & ~x627 & ~x640 & ~x654 & ~x672 & ~x682 & ~x683 & ~x699 & ~x702 & ~x705 & ~x707 & ~x708 & ~x710 & ~x735;
assign c5472 =  x375 &  x402 &  x429 & ~x270 & ~x313 & ~x324 & ~x327 & ~x624 & ~x735 & ~x782;
assign c5474 = ~x7 & ~x22 & ~x25 & ~x59 & ~x67 & ~x77 & ~x88 & ~x105 & ~x170 & ~x189 & ~x224 & ~x229 & ~x246 & ~x272 & ~x275 & ~x300 & ~x301 & ~x329 & ~x335 & ~x337 & ~x342 & ~x354 & ~x355 & ~x372 & ~x387 & ~x472 & ~x530 & ~x586 & ~x627 & ~x681 & ~x683 & ~x693 & ~x694 & ~x707 & ~x737 & ~x778;
assign c5476 =  x347 &  x374 &  x375 & ~x0 & ~x6 & ~x20 & ~x33 & ~x60 & ~x80 & ~x88 & ~x113 & ~x116 & ~x117 & ~x133 & ~x140 & ~x165 & ~x190 & ~x199 & ~x216 & ~x225 & ~x228 & ~x230 & ~x285 & ~x299 & ~x311 & ~x338 & ~x358 & ~x362 & ~x366 & ~x387 & ~x394 & ~x419 & ~x421 & ~x425 & ~x443 & ~x501 & ~x502 & ~x530 & ~x532 & ~x585 & ~x586 & ~x590 & ~x615 & ~x623 & ~x624 & ~x625 & ~x640 & ~x650 & ~x666 & ~x669 & ~x672 & ~x702 & ~x727 & ~x733 & ~x760 & ~x761;
assign c5478 =  x387 &  x445 & ~x633 & ~x660 & ~x686 & ~x689 & ~x690 & ~x694 & ~x715;
assign c5480 = ~x48 & ~x242 & ~x248 & ~x273 & ~x278 & ~x296 & ~x298 & ~x313 & ~x323 & ~x326 & ~x328 & ~x351 & ~x353 & ~x363 & ~x445 & ~x491 & ~x492 & ~x585 & ~x640 & ~x707 & ~x734 & ~x783;
assign c5482 =  x387 &  x530;
assign c5484 =  x187 &  x425 &  x453 &  x481 & ~x68 & ~x96 & ~x321 & ~x324 & ~x350 & ~x351 & ~x379 & ~x432 & ~x433 & ~x556 & ~x585 & ~x586 & ~x614 & ~x670 & ~x767 & ~x783;
assign c5486 =  x425 & ~x13 & ~x40 & ~x51 & ~x80 & ~x83 & ~x111 & ~x112 & ~x114 & ~x115 & ~x122 & ~x252 & ~x280 & ~x281 & ~x321 & ~x322 & ~x349 & ~x350 & ~x351 & ~x375 & ~x376 & ~x377 & ~x392 & ~x403 & ~x404 & ~x431 & ~x432 & ~x458 & ~x459 & ~x486 & ~x487 & ~x558 & ~x559 & ~x586 & ~x587 & ~x614 & ~x699 & ~x710 & ~x711 & ~x728 & ~x755 & ~x756 & ~x769;
assign c5488 = ~x84 & ~x93 & ~x120 & ~x139 & ~x308 & ~x355 & ~x410 & ~x412 & ~x441 & ~x467 & ~x541 & ~x569 & ~x584 & ~x628 & ~x658 & ~x696;
assign c5490 = ~x8 & ~x21 & ~x22 & ~x32 & ~x91 & ~x100 & ~x365 & ~x380 & ~x392 & ~x468 & ~x597 & ~x598 & ~x599 & ~x643 & ~x655 & ~x656 & ~x657 & ~x660 & ~x666 & ~x709 & ~x728 & ~x729 & ~x731 & ~x740 & ~x753;
assign c5492 = ~x27 & ~x31 & ~x55 & ~x64 & ~x85 & ~x91 & ~x92 & ~x115 & ~x118 & ~x119 & ~x137 & ~x176 & ~x177 & ~x267 & ~x336 & ~x381 & ~x382 & ~x411 & ~x412 & ~x572 & ~x584 & ~x612 & ~x626 & ~x638 & ~x782;
assign c5494 =  x756;
assign c5496 =  x213 &  x243 & ~x51 & ~x88 & ~x438 & ~x476 & ~x494 & ~x495 & ~x576;
assign c5498 =  x373 &  x510 & ~x50 & ~x465 & ~x466 & ~x519 & ~x520 & ~x546 & ~x551 & ~x735;
assign c51 =  x158 & ~x275 & ~x634 & ~x636 & ~x692 & ~x717;
assign c53 = ~x97 & ~x195 & ~x308 & ~x353 & ~x388 & ~x389 & ~x462 & ~x489 & ~x517 & ~x518 & ~x575 & ~x605 & ~x630 & ~x756;
assign c55 =  x438 & ~x2 & ~x4 & ~x10 & ~x37 & ~x459 & ~x671 & ~x703 & ~x732 & ~x734 & ~x736 & ~x758 & ~x759 & ~x761 & ~x765 & ~x766 & ~x779;
assign c57 = ~x302 & ~x426 & ~x521 & ~x684 & ~x718 & ~x744;
assign c59 =  x93 & ~x24 & ~x27 & ~x55 & ~x56 & ~x139 & ~x454 & ~x483 & ~x700 & ~x702 & ~x758;
assign c511 =  x439 &  x542 & ~x669;
assign c513 =  x681 & ~x369 & ~x615 & ~x751 & ~x753 & ~x755 & ~x758 & ~x778;
assign c515 =  x285 &  x430 & ~x0 & ~x56 & ~x530 & ~x531 & ~x557 & ~x616 & ~x756;
assign c517 =  x285 & ~x443 & ~x446 & ~x448 & ~x656;
assign c519 =  x401 &  x461 & ~x10 & ~x29 & ~x56 & ~x109 & ~x139 & ~x142 & ~x167 & ~x674 & ~x724 & ~x725 & ~x727 & ~x728 & ~x759 & ~x780;
assign c521 =  x205 & ~x113 & ~x119 & ~x589 & ~x672 & ~x673 & ~x684 & ~x705;
assign c523 =  x294 & ~x27 & ~x58 & ~x109 & ~x166 & ~x201 & ~x251 & ~x253 & ~x627 & ~x632 & ~x633 & ~x660 & ~x661 & ~x775;
assign c525 =  x269 &  x494 & ~x27 & ~x196 & ~x280 & ~x734 & ~x761 & ~x762;
assign c527 = ~x72 & ~x183 & ~x389 & ~x399 & ~x438 & ~x522;
assign c529 =  x599 & ~x7 & ~x13 & ~x18 & ~x25 & ~x49 & ~x50 & ~x157 & ~x722 & ~x775;
assign c531 =  x266 & ~x0 & ~x2 & ~x29 & ~x30 & ~x45 & ~x298 & ~x531 & ~x563 & ~x706 & ~x743 & ~x745;
assign c533 = ~x350 & ~x367 & ~x372 & ~x398 & ~x426 & ~x452 & ~x453 & ~x534;
assign c535 = ~x25 & ~x52 & ~x72 & ~x138 & ~x146 & ~x438 & ~x441 & ~x480 & ~x481 & ~x483 & ~x505 & ~x509 & ~x535 & ~x536 & ~x564 & ~x567 & ~x588 & ~x595 & ~x596 & ~x619 & ~x621 & ~x623 & ~x624 & ~x777;
assign c537 =  x369 &  x406;
assign c539 =  x380 & ~x50 & ~x469 & ~x680 & ~x687;
assign c541 = ~x2 & ~x8 & ~x9 & ~x25 & ~x31 & ~x33 & ~x36 & ~x62 & ~x83 & ~x116 & ~x385 & ~x405 & ~x455 & ~x482 & ~x483 & ~x484 & ~x506 & ~x532 & ~x533 & ~x537 & ~x539 & ~x540 & ~x560 & ~x561 & ~x563 & ~x569 & ~x587 & ~x588 & ~x674 & ~x731 & ~x762 & ~x768;
assign c543 = ~x130 & ~x156 & ~x157 & ~x195 & ~x269 & ~x271 & ~x276 & ~x296 & ~x299 & ~x324 & ~x352 & ~x495 & ~x549 & ~x634;
assign c545 =  x550 & ~x634 & ~x635 & ~x636 & ~x662 & ~x663 & ~x781;
assign c547 =  x186 & ~x8 & ~x27 & ~x34 & ~x223 & ~x244 & ~x616 & ~x653 & ~x700 & ~x702 & ~x732;
assign c549 =  x534 & ~x0 & ~x1 & ~x28 & ~x29 & ~x32 & ~x56 & ~x57 & ~x83 & ~x86 & ~x111 & ~x139 & ~x143 & ~x170 & ~x195 & ~x198 & ~x199 & ~x223 & ~x224 & ~x253 & ~x279 & ~x308 & ~x335 & ~x363 & ~x364 & ~x420 & ~x448 & ~x521 & ~x548 & ~x574 & ~x604 & ~x605;
assign c551 =  x206 &  x211 & ~x110 & ~x140 & ~x483 & ~x615 & ~x671;
assign c553 =  x102 & ~x4 & ~x31 & ~x99 & ~x188;
assign c555 =  x297 &  x553 & ~x252;
assign c557 =  x108 & ~x274 & ~x448;
assign c559 =  x94 & ~x490 & ~x645 & ~x646 & ~x684;
assign c561 = ~x0 & ~x23 & ~x26 & ~x71 & ~x186 & ~x212 & ~x240 & ~x249 & ~x250 & ~x299 & ~x364 & ~x383 & ~x411 & ~x466 & ~x697 & ~x776;
assign c563 =  x186 & ~x427 & ~x503 & ~x659;
assign c565 =  x573 & ~x3 & ~x27 & ~x31 & ~x158 & ~x214 & ~x394 & ~x421 & ~x699 & ~x727 & ~x758 & ~x762 & ~x780;
assign c567 =  x259 &  x460 & ~x725 & ~x756 & ~x761 & ~x782 & ~x783;
assign c569 =  x434 & ~x3 & ~x10 & ~x37 & ~x350 & ~x782;
assign c571 =  x264 & ~x23 & ~x52 & ~x141 & ~x253 & ~x433 & ~x458 & ~x672 & ~x737 & ~x750 & ~x761 & ~x763 & ~x766 & ~x776 & ~x779;
assign c573 =  x376 & ~x15 & ~x23 & ~x69 & ~x70 & ~x71 & ~x97 & ~x98 & ~x124 & ~x280 & ~x308 & ~x559 & ~x587 & ~x616;
assign c575 =  x426 & ~x56 & ~x188 & ~x733 & ~x761;
assign c577 =  x432 & ~x11 & ~x19 & ~x38 & ~x128 & ~x743 & ~x756 & ~x764;
assign c579 =  x294 & ~x25 & ~x26 & ~x326 & ~x405 & ~x560 & ~x561 & ~x608 & ~x673;
assign c581 =  x379 & ~x26 & ~x27 & ~x53 & ~x54 & ~x55 & ~x77 & ~x83 & ~x86 & ~x475 & ~x501 & ~x504 & ~x671 & ~x687 & ~x699 & ~x727;
assign c583 =  x262 &  x263 & ~x10 & ~x11 & ~x12 & ~x13 & ~x35 & ~x39 & ~x143 & ~x198 & ~x704 & ~x748 & ~x749 & ~x750 & ~x751 & ~x761;
assign c585 =  x628 & ~x3 & ~x47 & ~x52 & ~x59 & ~x158 & ~x496 & ~x667 & ~x699 & ~x706 & ~x730 & ~x748 & ~x749 & ~x750 & ~x758 & ~x763 & ~x776 & ~x780;
assign c587 =  x185 &  x291 & ~x567 & ~x656 & ~x680 & ~x684 & ~x709 & ~x733;
assign c589 = ~x29 & ~x53 & ~x56 & ~x88 & ~x104 & ~x167 & ~x195 & ~x281 & ~x333 & ~x337 & ~x361 & ~x409 & ~x416 & ~x436 & ~x444 & ~x448 & ~x606 & ~x660 & ~x662 & ~x777 & ~x778 & ~x779 & ~x780 & ~x783;
assign c591 =  x380 & ~x20 & ~x472 & ~x528 & ~x554 & ~x601;
assign c593 =  x69 & ~x377 & ~x429 & ~x457 & ~x704;
assign c595 =  x260 & ~x5 & ~x7 & ~x12 & ~x23 & ~x24 & ~x26 & ~x27 & ~x39 & ~x51 & ~x55 & ~x56 & ~x84 & ~x130 & ~x140 & ~x614 & ~x640 & ~x641 & ~x668 & ~x669 & ~x672 & ~x675 & ~x695 & ~x697 & ~x699 & ~x700 & ~x703 & ~x722 & ~x724 & ~x727 & ~x730 & ~x734 & ~x750 & ~x753 & ~x755 & ~x756 & ~x757 & ~x758 & ~x759 & ~x760 & ~x761 & ~x764 & ~x776 & ~x783;
assign c597 =  x201 & ~x0 & ~x5 & ~x18 & ~x161 & ~x585 & ~x757 & ~x783;
assign c599 = ~x226 & ~x228 & ~x254 & ~x256 & ~x438 & ~x485 & ~x515 & ~x548 & ~x616 & ~x647 & ~x723 & ~x750 & ~x776;
assign c5101 =  x80;
assign c5103 =  x174 &  x461 & ~x19 & ~x25 & ~x46;
assign c5105 =  x429 &  x506 & ~x59 & ~x83 & ~x167 & ~x364 & ~x727 & ~x758 & ~x759;
assign c5107 =  x305 & ~x24 & ~x25 & ~x26 & ~x30 & ~x50 & ~x78 & ~x82 & ~x109 & ~x167 & ~x483 & ~x504 & ~x510 & ~x532 & ~x560 & ~x561 & ~x562 & ~x572 & ~x588 & ~x589 & ~x618 & ~x621 & ~x645 & ~x651 & ~x673 & ~x676 & ~x677 & ~x701 & ~x730 & ~x733 & ~x759 & ~x760 & ~x765 & ~x781;
assign c5109 =  x260 & ~x21 & ~x77 & ~x113 & ~x114 & ~x143 & ~x411 & ~x645 & ~x674 & ~x693 & ~x700 & ~x721 & ~x732 & ~x734;
assign c5111 = ~x55 & ~x203 & ~x231 & ~x313 & ~x369 & ~x526 & ~x599 & ~x601 & ~x603 & ~x615 & ~x628;
assign c5113 =  x241 & ~x28 & ~x92 & ~x138 & ~x139 & ~x142 & ~x167 & ~x454 & ~x508 & ~x615 & ~x755 & ~x777 & ~x780;
assign c5115 =  x379 & ~x28 & ~x45 & ~x53 & ~x111 & ~x167 & ~x412 & ~x504 & ~x650 & ~x700 & ~x727 & ~x760 & ~x774 & ~x776;
assign c5117 =  x191 & ~x16 & ~x19 & ~x341 & ~x616 & ~x673;
assign c5119 =  x517 &  x518 &  x546 & ~x8 & ~x609 & ~x635 & ~x695 & ~x761 & ~x762 & ~x777;
assign c5121 =  x242 & ~x272 & ~x273 & ~x488;
assign c5123 = ~x27 & ~x55 & ~x196 & ~x224 & ~x252 & ~x281 & ~x399 & ~x427 & ~x435 & ~x490 & ~x518 & ~x519 & ~x545 & ~x547 & ~x657;
assign c5125 =  x293 &  x439 & ~x10 & ~x12;
assign c5127 =  x370 &  x544 & ~x3 & ~x760 & ~x761;
assign c5129 = ~x3 & ~x89 & ~x168 & ~x441 & ~x460 & ~x461 & ~x482 & ~x485 & ~x490 & ~x507 & ~x513 & ~x619;
assign c5131 =  x581 & ~x471 & ~x605 & ~x663;
assign c5133 = ~x19 & ~x22 & ~x42 & ~x424 & ~x451 & ~x456 & ~x512 & ~x593 & ~x616 & ~x652 & ~x754 & ~x766;
assign c5135 =  x527 & ~x195 & ~x477 & ~x496 & ~x585 & ~x615;
assign c5137 =  x266 & ~x25 & ~x27 & ~x114 & ~x224 & ~x241 & ~x269 & ~x475 & ~x531 & ~x553 & ~x632 & ~x752;
assign c5139 =  x317 &  x583 & ~x172;
assign c5141 = ~x8 & ~x20 & ~x404 & ~x405 & ~x450 & ~x453 & ~x454 & ~x511 & ~x616 & ~x617 & ~x620 & ~x776;
assign c5143 =  x556 & ~x168 & ~x199 & ~x224 & ~x470;
assign c5145 =  x379 & ~x26 & ~x212 & ~x309 & ~x411 & ~x607 & ~x783;
assign c5147 =  x120 & ~x167 & ~x187 & ~x309 & ~x364 & ~x448 & ~x759;
assign c5149 =  x180 &  x208 & ~x7 & ~x33 & ~x141 & ~x169 & ~x428 & ~x466 & ~x484 & ~x644 & ~x727 & ~x732 & ~x733 & ~x753 & ~x755;
assign c5151 =  x155 &  x409 & ~x1 & ~x23 & ~x24 & ~x26 & ~x27 & ~x52 & ~x53 & ~x54 & ~x55 & ~x56 & ~x57 & ~x79 & ~x84 & ~x109 & ~x138 & ~x139 & ~x195 & ~x223 & ~x308 & ~x671 & ~x761;
assign c5153 = ~x43 & ~x281 & ~x288 & ~x445 & ~x446 & ~x521 & ~x601 & ~x656 & ~x661;
assign c5155 =  x324 & ~x279 & ~x475 & ~x526 & ~x545 & ~x573 & ~x777;
assign c5157 =  x418 & ~x4 & ~x28 & ~x83 & ~x112 & ~x358 & ~x560 & ~x589 & ~x617 & ~x619 & ~x644 & ~x645 & ~x649 & ~x700;
assign c5159 =  x50;
assign c5161 =  x710 & ~x52 & ~x252 & ~x511 & ~x783;
assign c5163 =  x178 & ~x3 & ~x55 & ~x403 & ~x511 & ~x702 & ~x727 & ~x760;
assign c5165 =  x208 &  x499 & ~x26;
assign c5167 =  x352 & ~x384 & ~x440 & ~x573 & ~x615;
assign c5169 = ~x54 & ~x409 & ~x428 & ~x493 & ~x506 & ~x531 & ~x534 & ~x640 & ~x663 & ~x719 & ~x730 & ~x747;
assign c5171 =  x324 &  x551 & ~x587;
assign c5173 =  x358 &  x519 & ~x26 & ~x192 & ~x587;
assign c5175 =  x484 & ~x21 & ~x23 & ~x25 & ~x139 & ~x167 & ~x391 & ~x418 & ~x444 & ~x471 & ~x473 & ~x744 & ~x746;
assign c5177 =  x599 & ~x13 & ~x19 & ~x101 & ~x184 & ~x466;
assign c5179 =  x416 &  x490;
assign c5181 =  x66 & ~x0 & ~x28 & ~x112 & ~x169 & ~x195 & ~x225 & ~x252 & ~x406 & ~x419 & ~x515 & ~x728;
assign c5183 =  x261 &  x288 & ~x19 & ~x27 & ~x29 & ~x32 & ~x56 & ~x57 & ~x60 & ~x168 & ~x170 & ~x197 & ~x203 & ~x511 & ~x748 & ~x760 & ~x761;
assign c5185 =  x108 & ~x302 & ~x783;
assign c5187 = ~x174 & ~x282 & ~x358 & ~x436 & ~x544 & ~x550 & ~x578 & ~x764 & ~x777;
assign c5189 =  x325 & ~x442 & ~x553 & ~x650 & ~x675 & ~x676 & ~x706 & ~x732 & ~x777;
assign c5191 =  x680 & ~x251 & ~x409;
assign c5193 = ~x65 & ~x313 & ~x339 & ~x433 & ~x509 & ~x534 & ~x559 & ~x562 & ~x710 & ~x755 & ~x765 & ~x777 & ~x782;
assign c5195 =  x267 & ~x168 & ~x327 & ~x328 & ~x599 & ~x605 & ~x625;
assign c5197 = ~x194 & ~x333 & ~x408 & ~x415 & ~x528 & ~x576 & ~x603 & ~x741;
assign c5199 =  x38 & ~x28 & ~x29 & ~x627 & ~x628 & ~x702;
assign c5201 =  x244 &  x350 & ~x134 & ~x691 & ~x780;
assign c5203 = ~x370 & ~x376 & ~x383 & ~x395 & ~x433 & ~x541;
assign c5205 =  x292 & ~x199 & ~x330 & ~x463 & ~x512 & ~x519 & ~x575 & ~x604;
assign c5207 = ~x21 & ~x24 & ~x46 & ~x47 & ~x104 & ~x128 & ~x298 & ~x299 & ~x324 & ~x326 & ~x352 & ~x353 & ~x391 & ~x497 & ~x523 & ~x549 & ~x551 & ~x671 & ~x698 & ~x721 & ~x727 & ~x777;
assign c5209 = ~x140 & ~x224 & ~x252 & ~x264 & ~x335 & ~x364 & ~x441 & ~x447 & ~x521 & ~x571 & ~x578 & ~x663;
assign c5211 =  x236 &  x287 & ~x27 & ~x53 & ~x81 & ~x108 & ~x110 & ~x139 & ~x140 & ~x143 & ~x509 & ~x536 & ~x537 & ~x561 & ~x615 & ~x728 & ~x755 & ~x757 & ~x758;
assign c5213 =  x710 & ~x26 & ~x111 & ~x364 & ~x392 & ~x587 & ~x615 & ~x626 & ~x699 & ~x755;
assign c5215 =  x191 & ~x62 & ~x304 & ~x332;
assign c5217 = ~x1 & ~x23 & ~x27 & ~x33 & ~x54 & ~x55 & ~x59 & ~x115 & ~x165 & ~x171 & ~x194 & ~x196 & ~x197 & ~x228 & ~x279 & ~x306 & ~x308 & ~x311 & ~x336 & ~x337 & ~x362 & ~x420 & ~x421 & ~x443 & ~x475 & ~x577 & ~x599 & ~x601 & ~x602 & ~x604 & ~x605 & ~x782 & ~x783;
assign c5219 = ~x26 & ~x35 & ~x84 & ~x111 & ~x112 & ~x168 & ~x276 & ~x526 & ~x601 & ~x603 & ~x618 & ~x626 & ~x628;
assign c5221 =  x430 & ~x41 & ~x42 & ~x318 & ~x615 & ~x699;
assign c5223 =  x261 &  x311 & ~x130;
assign c5225 =  x563 &  x651;
assign c5227 =  x512 &  x520 &  x539 & ~x0 & ~x20 & ~x26 & ~x27 & ~x54 & ~x55;
assign c5229 =  x143 & ~x388;
assign c5231 =  x77 & ~x357 & ~x448;
assign c5233 =  x654 & ~x140 & ~x410 & ~x643 & ~x748 & ~x766 & ~x777 & ~x781;
assign c5235 =  x435 & ~x190 & ~x496 & ~x575 & ~x580;
assign c5237 =  x344 &  x407 & ~x23 & ~x30 & ~x586 & ~x782;
assign c5239 =  x432 & ~x24 & ~x419 & ~x587 & ~x615 & ~x616 & ~x715 & ~x716 & ~x743 & ~x755 & ~x762 & ~x772;
assign c5241 =  x653 & ~x26 & ~x45 & ~x214 & ~x672 & ~x757;
assign c5243 = ~x61 & ~x63 & ~x348 & ~x392 & ~x395 & ~x503 & ~x506 & ~x539 & ~x561 & ~x594 & ~x609 & ~x610 & ~x612 & ~x623 & ~x652 & ~x668 & ~x681 & ~x736;
assign c5245 =  x354 &  x381 & ~x23 & ~x25 & ~x54 & ~x83 & ~x441 & ~x443 & ~x733 & ~x734 & ~x764 & ~x782;
assign c5247 =  x436 &  x572 & ~x23 & ~x25 & ~x106;
assign c5249 =  x258 &  x283 & ~x199 & ~x420;
assign c5251 =  x205 & ~x0 & ~x7 & ~x27 & ~x29 & ~x31 & ~x380 & ~x408 & ~x409 & ~x415 & ~x503 & ~x616 & ~x698 & ~x699 & ~x703 & ~x722 & ~x726 & ~x727 & ~x750 & ~x757 & ~x758 & ~x761 & ~x762;
assign c5253 =  x324 & ~x196 & ~x384 & ~x713 & ~x720;
assign c5255 = ~x1 & ~x3 & ~x5 & ~x7 & ~x11 & ~x12 & ~x22 & ~x27 & ~x31 & ~x55 & ~x56 & ~x62 & ~x65 & ~x80 & ~x112 & ~x224 & ~x231 & ~x232 & ~x252 & ~x253 & ~x254 & ~x258 & ~x281 & ~x285 & ~x309 & ~x615 & ~x642 & ~x643 & ~x706 & ~x727 & ~x732 & ~x734 & ~x735 & ~x741 & ~x742 & ~x749 & ~x750 & ~x751 & ~x755 & ~x756 & ~x761 & ~x775 & ~x776;
assign c5257 =  x657 & ~x139 & ~x185 & ~x392 & ~x466 & ~x694 & ~x695 & ~x696 & ~x722 & ~x749;
assign c5259 = ~x313 & ~x352 & ~x428 & ~x432 & ~x433 & ~x478 & ~x535 & ~x649 & ~x734 & ~x761;
assign c5261 =  x361 & ~x134 & ~x161 & ~x503 & ~x532 & ~x561 & ~x617 & ~x670 & ~x735 & ~x751 & ~x765 & ~x776;
assign c5263 =  x324 &  x351 & ~x252 & ~x309 & ~x384 & ~x409 & ~x410 & ~x615 & ~x777;
assign c5265 = ~x40 & ~x49 & ~x259 & ~x275 & ~x415 & ~x642 & ~x643 & ~x660 & ~x687 & ~x688 & ~x783;
assign c5267 =  x707 & ~x83 & ~x244 & ~x336;
assign c5269 =  x380 &  x430 & ~x495 & ~x698 & ~x733 & ~x760;
assign c5271 =  x508 &  x595 & ~x336 & ~x778;
assign c5273 =  x234 & ~x172 & ~x465 & ~x494 & ~x511 & ~x745;
assign c5275 =  x201 &  x202 & ~x83 & ~x309 & ~x342 & ~x447;
assign c5277 = ~x22 & ~x31 & ~x135 & ~x137 & ~x165 & ~x168 & ~x192 & ~x204 & ~x221 & ~x223 & ~x390 & ~x392 & ~x418 & ~x446 & ~x472 & ~x474 & ~x499 & ~x501 & ~x559 & ~x602 & ~x603 & ~x630 & ~x661 & ~x662;
assign c5279 = ~x142 & ~x430 & ~x532 & ~x551 & ~x559 & ~x561 & ~x562 & ~x587 & ~x590 & ~x594 & ~x649 & ~x652 & ~x738 & ~x776;
assign c5281 =  x625 & ~x22 & ~x72 & ~x643 & ~x718 & ~x757 & ~x760 & ~x761;
assign c5283 =  x299 & ~x1 & ~x55 & ~x224 & ~x251 & ~x387 & ~x689 & ~x717 & ~x718 & ~x763;
assign c5285 =  x358 & ~x0 & ~x1 & ~x25 & ~x58 & ~x84 & ~x112 & ~x164 & ~x169 & ~x171 & ~x201 & ~x226 & ~x251 & ~x308 & ~x560 & ~x616;
assign c5287 =  x230 & ~x2 & ~x5 & ~x25 & ~x27 & ~x57 & ~x69 & ~x316 & ~x338 & ~x392 & ~x736 & ~x737 & ~x764 & ~x765 & ~x783;
assign c5289 = ~x8 & ~x56 & ~x129 & ~x195 & ~x246 & ~x413 & ~x615 & ~x636 & ~x663 & ~x666 & ~x713 & ~x746 & ~x752 & ~x763 & ~x781;
assign c5291 =  x255 &  x256 & ~x74 & ~x301;
assign c5293 =  x269 &  x346 & ~x644;
assign c5295 =  x322 & ~x0 & ~x18 & ~x25 & ~x26 & ~x41 & ~x42 & ~x503 & ~x504 & ~x529 & ~x644 & ~x699 & ~x755;
assign c5297 = ~x40 & ~x201 & ~x202 & ~x483 & ~x533 & ~x534 & ~x540 & ~x544 & ~x560 & ~x561 & ~x574 & ~x589 & ~x645 & ~x646 & ~x761;
assign c5299 =  x406 & ~x10 & ~x19 & ~x24 & ~x25 & ~x49 & ~x50 & ~x83 & ~x476 & ~x530 & ~x557 & ~x672 & ~x729 & ~x748 & ~x752 & ~x758 & ~x772 & ~x773 & ~x774 & ~x776;
assign c5301 =  x462 & ~x73 & ~x138 & ~x212 & ~x522 & ~x550 & ~x551 & ~x733 & ~x751;
assign c5303 =  x259 & ~x26 & ~x58 & ~x127 & ~x128 & ~x154 & ~x193 & ~x221 & ~x222 & ~x251 & ~x279 & ~x327 & ~x644 & ~x645 & ~x700 & ~x757;
assign c5305 =  x562 &  x622 & ~x5 & ~x56 & ~x335;
assign c5307 = ~x77 & ~x345 & ~x396 & ~x449 & ~x457 & ~x482 & ~x511 & ~x513 & ~x590 & ~x766;
assign c5309 =  x408 & ~x234 & ~x280 & ~x575;
assign c5311 =  x402 &  x520 & ~x1 & ~x28 & ~x29 & ~x236 & ~x252 & ~x727 & ~x781 & ~x782;
assign c5313 =  x610 & ~x117 & ~x198 & ~x199 & ~x381 & ~x518 & ~x521 & ~x780;
assign c5315 = ~x22 & ~x178 & ~x304 & ~x331 & ~x429 & ~x486 & ~x551 & ~x732;
assign c5317 =  x175 &  x507 & ~x753;
assign c5319 = ~x9 & ~x55 & ~x235 & ~x244 & ~x336 & ~x392 & ~x671 & ~x761 & ~x783;
assign c5321 =  x260 &  x287 & ~x74 & ~x101 & ~x106 & ~x128 & ~x345 & ~x420 & ~x755;
assign c5323 =  x555 & ~x33 & ~x441 & ~x475;
assign c5325 =  x627 &  x628 & ~x157 & ~x587 & ~x748 & ~x749 & ~x750;
assign c5327 =  x491 & ~x46 & ~x106 & ~x269 & ~x270 & ~x297 & ~x325 & ~x421 & ~x476 & ~x579 & ~x581 & ~x608;
assign c5329 =  x261 &  x718 & ~x455 & ~x538 & ~x644 & ~x776;
assign c5331 =  x204 & ~x8 & ~x24 & ~x142 & ~x382 & ~x644 & ~x669 & ~x702 & ~x718 & ~x759;
assign c5333 = ~x8 & ~x19 & ~x318 & ~x368 & ~x396 & ~x398 & ~x450 & ~x485 & ~x562 & ~x588 & ~x616 & ~x623 & ~x641 & ~x648 & ~x699 & ~x724;
assign c5335 =  x109;
assign c5337 =  x437 & ~x0 & ~x26 & ~x189 & ~x233 & ~x497 & ~x644;
assign c5339 =  x708 & ~x0 & ~x244 & ~x615;
assign c5341 =  x288 &  x311 & ~x3 & ~x441;
assign c5343 =  x352 & ~x0 & ~x8 & ~x56 & ~x178 & ~x504 & ~x586 & ~x596 & ~x643 & ~x761;
assign c5345 =  x151 & ~x2 & ~x7 & ~x8 & ~x25 & ~x33 & ~x34 & ~x37 & ~x171 & ~x587 & ~x617 & ~x644 & ~x669 & ~x698 & ~x733 & ~x747 & ~x762 & ~x774;
assign c5347 =  x221 & ~x196 & ~x442 & ~x764;
assign c5349 =  x434 &  x572 & ~x1 & ~x4 & ~x27 & ~x49 & ~x51 & ~x55 & ~x56 & ~x83 & ~x113 & ~x135 & ~x138 & ~x224 & ~x308 & ~x448 & ~x476 & ~x727;
assign c5351 =  x404 & ~x84 & ~x85 & ~x280 & ~x291 & ~x319 & ~x476 & ~x531 & ~x559 & ~x587 & ~x642 & ~x643 & ~x670 & ~x727;
assign c5353 =  x740 & ~x3 & ~x112 & ~x744 & ~x756;
assign c5355 =  x381 & ~x0 & ~x179 & ~x180 & ~x733;
assign c5357 =  x529 & ~x31 & ~x57 & ~x84 & ~x443 & ~x471;
assign c5359 =  x175 &  x201 & ~x24 & ~x43 & ~x55 & ~x58 & ~x82 & ~x448 & ~x761;
assign c5361 =  x488 & ~x10 & ~x12 & ~x94 & ~x105 & ~x733 & ~x759 & ~x760 & ~x761 & ~x770 & ~x771 & ~x773 & ~x778;
assign c5363 = ~x84 & ~x138 & ~x165 & ~x222 & ~x280 & ~x281 & ~x307 & ~x333 & ~x361 & ~x418 & ~x472 & ~x574 & ~x575 & ~x576 & ~x600 & ~x601 & ~x603 & ~x606 & ~x627;
assign c5365 =  x299 & ~x103 & ~x415 & ~x447 & ~x705;
assign c5367 =  x516 & ~x21 & ~x39 & ~x40 & ~x52 & ~x53 & ~x614 & ~x636 & ~x643 & ~x776;
assign c5369 =  x709 & ~x83 & ~x453 & ~x699;
assign c5371 =  x230 & ~x1 & ~x16 & ~x29 & ~x81 & ~x108 & ~x131 & ~x267 & ~x557 & ~x699;
assign c5373 =  x150 &  x260 & ~x118 & ~x626;
assign c5375 = ~x168 & ~x261 & ~x280 & ~x388 & ~x389 & ~x569 & ~x587 & ~x599 & ~x604 & ~x632 & ~x745 & ~x746;
assign c5377 =  x491 &  x519 &  x520 & ~x2 & ~x3 & ~x134 & ~x139 & ~x219 & ~x580 & ~x699;
assign c5379 =  x260 &  x310 & ~x112 & ~x448;
assign c5381 =  x518 & ~x500 & ~x558 & ~x581 & ~x582 & ~x658 & ~x664 & ~x761;
assign c5383 =  x353 & ~x167 & ~x470 & ~x572 & ~x600 & ~x626;
assign c5385 = ~x5 & ~x22 & ~x25 & ~x26 & ~x27 & ~x114 & ~x140 & ~x196 & ~x224 & ~x276 & ~x304 & ~x472 & ~x547 & ~x576 & ~x605 & ~x630 & ~x632 & ~x633 & ~x634 & ~x741;
assign c5387 =  x264 & ~x197 & ~x376 & ~x377 & ~x534 & ~x718 & ~x762 & ~x777;
assign c5389 =  x190 & ~x468 & ~x562 & ~x563 & ~x591 & ~x677 & ~x705 & ~x728;
assign c5391 =  x137;
assign c5393 =  x128 & ~x6 & ~x20 & ~x26 & ~x27 & ~x37 & ~x132 & ~x159 & ~x160 & ~x196 & ~x708 & ~x734 & ~x753 & ~x761 & ~x762 & ~x763 & ~x776 & ~x781 & ~x782 & ~x783;
assign c5395 =  x463 &  x491 &  x519 &  x547 &  x575 & ~x25 & ~x26 & ~x27 & ~x55 & ~x80 & ~x82 & ~x392 & ~x504 & ~x560;
assign c5397 =  x178 & ~x28 & ~x409 & ~x437 & ~x464 & ~x564 & ~x747 & ~x762;
assign c5399 =  x562 &  x594 & ~x778;
assign c5401 =  x462 & ~x16 & ~x73 & ~x74 & ~x272 & ~x523 & ~x579 & ~x766;
assign c5403 =  x266 & ~x73 & ~x196 & ~x229 & ~x383 & ~x410 & ~x540 & ~x620 & ~x648 & ~x650;
assign c5405 =  x121 & ~x5 & ~x26 & ~x55 & ~x83 & ~x482 & ~x644 & ~x674;
assign c5407 =  x638 & ~x30 & ~x53 & ~x115 & ~x143 & ~x280 & ~x489 & ~x545 & ~x574;
assign c5409 =  x183 &  x410 & ~x28 & ~x59 & ~x732 & ~x757 & ~x759 & ~x779;
assign c5411 = ~x159 & ~x213 & ~x214 & ~x222 & ~x224 & ~x228 & ~x374 & ~x732;
assign c5413 =  x176 &  x204 &  x428 & ~x26 & ~x115 & ~x116 & ~x338 & ~x765;
assign c5415 =  x248 &  x249 & ~x32 & ~x137 & ~x563 & ~x591 & ~x649;
assign c5417 =  x624 & ~x21 & ~x32 & ~x59 & ~x114 & ~x142 & ~x171 & ~x198 & ~x199 & ~x226 & ~x756 & ~x757 & ~x760 & ~x772 & ~x783;
assign c5419 =  x154 &  x178 &  x180 & ~x5 & ~x7 & ~x139 & ~x171 & ~x726 & ~x732 & ~x755;
assign c5421 =  x343 & ~x130 & ~x733;
assign c5423 =  x203 & ~x16 & ~x29 & ~x30 & ~x316 & ~x336 & ~x337 & ~x366 & ~x392 & ~x655 & ~x682 & ~x699;
assign c5425 =  x177 &  x204 & ~x7 & ~x27 & ~x28 & ~x29 & ~x32 & ~x55 & ~x56 & ~x391 & ~x392 & ~x643 & ~x733 & ~x753 & ~x759 & ~x764;
assign c5427 =  x295 & ~x14 & ~x26 & ~x260 & ~x623 & ~x758;
assign c5429 = ~x83 & ~x87 & ~x138 & ~x139 & ~x169 & ~x248 & ~x309 & ~x444 & ~x602 & ~x626 & ~x634 & ~x639 & ~x657 & ~x700;
assign c5431 =  x296 & ~x14 & ~x22 & ~x50 & ~x308 & ~x356 & ~x624 & ~x652 & ~x723 & ~x724 & ~x752 & ~x756;
assign c5433 =  x319 &  x425 & ~x3 & ~x85 & ~x114 & ~x137 & ~x167 & ~x170 & ~x171 & ~x193 & ~x198 & ~x223 & ~x228 & ~x251 & ~x253 & ~x255 & ~x643 & ~x760;
assign c5435 =  x492 & ~x19 & ~x26 & ~x27 & ~x28 & ~x30 & ~x49 & ~x56 & ~x74 & ~x261 & ~x504 & ~x552 & ~x759;
assign c5437 =  x460 & ~x20 & ~x22 & ~x25 & ~x50 & ~x184 & ~x212 & ~x394 & ~x467 & ~x494 & ~x523 & ~x578 & ~x697 & ~x700 & ~x704 & ~x725 & ~x727 & ~x754;
assign c5439 =  x707 & ~x299;
assign c5441 =  x183 &  x468 & ~x7 & ~x27 & ~x143 & ~x167 & ~x223 & ~x757;
assign c5443 = ~x17 & ~x45 & ~x65 & ~x84 & ~x359 & ~x457 & ~x562 & ~x639 & ~x707 & ~x729 & ~x733 & ~x739 & ~x774 & ~x780;
assign c5445 =  x709 &  x710 &  x711 & ~x757;
assign c5447 = ~x1 & ~x29 & ~x78 & ~x195 & ~x196 & ~x276 & ~x279 & ~x305 & ~x308 & ~x362 & ~x363 & ~x392 & ~x444 & ~x471 & ~x473 & ~x499 & ~x501 & ~x604 & ~x631 & ~x632 & ~x658 & ~x659 & ~x661 & ~x683 & ~x727;
assign c5449 =  x312 & ~x104 & ~x196 & ~x307 & ~x443 & ~x471 & ~x653 & ~x763;
assign c5451 =  x66 & ~x57 & ~x85 & ~x454 & ~x517 & ~x701 & ~x783;
assign c5453 = ~x5 & ~x7 & ~x19 & ~x60 & ~x340 & ~x381 & ~x401 & ~x415 & ~x508 & ~x522 & ~x550 & ~x615 & ~x700 & ~x718 & ~x746 & ~x774;
assign c5455 = ~x68 & ~x82 & ~x83 & ~x185 & ~x238 & ~x239 & ~x373 & ~x385 & ~x394 & ~x438;
assign c5457 =  x291 & ~x68 & ~x70 & ~x97 & ~x140 & ~x223 & ~x225 & ~x233 & ~x260 & ~x679;
assign c5459 =  x416 & ~x195 & ~x223 & ~x251 & ~x357 & ~x475 & ~x502 & ~x589 & ~x701;
assign c5461 =  x333 & ~x26 & ~x51 & ~x53 & ~x54 & ~x82 & ~x168 & ~x346 & ~x396 & ~x397 & ~x422 & ~x503 & ~x532 & ~x560 & ~x672 & ~x728 & ~x729 & ~x732;
assign c5463 =  x534 &  x678;
assign c5465 =  x151 & ~x114 & ~x145 & ~x460 & ~x676;
assign c5467 =  x646 & ~x0 & ~x28 & ~x112 & ~x140 & ~x253 & ~x363 & ~x391 & ~x419 & ~x685;
assign c5469 =  x323 & ~x528 & ~x530 & ~x531 & ~x587 & ~x616 & ~x744 & ~x762 & ~x772;
assign c5471 =  x205 & ~x26 & ~x54 & ~x482 & ~x509 & ~x625 & ~x626 & ~x749 & ~x765 & ~x778;
assign c5473 =  x414 & ~x0 & ~x1 & ~x26 & ~x56 & ~x84 & ~x86 & ~x113 & ~x116 & ~x140 & ~x193 & ~x196 & ~x223 & ~x224 & ~x447 & ~x473 & ~x529 & ~x559 & ~x587 & ~x728 & ~x756;
assign c5475 = ~x8 & ~x73 & ~x79 & ~x100 & ~x129 & ~x185 & ~x215 & ~x325 & ~x477 & ~x495 & ~x496 & ~x523 & ~x531 & ~x612 & ~x728 & ~x748 & ~x750 & ~x757;
assign c5477 =  x261 & ~x493 & ~x511 & ~x522 & ~x693 & ~x695;
assign c5479 = ~x26 & ~x84 & ~x109 & ~x115 & ~x165 & ~x223 & ~x360 & ~x380 & ~x463 & ~x464 & ~x528 & ~x576 & ~x631 & ~x688 & ~x689 & ~x783;
assign c5481 =  x435 &  x571 & ~x4 & ~x19 & ~x587 & ~x642 & ~x756 & ~x783;
assign c5483 = ~x2 & ~x3 & ~x7 & ~x12 & ~x23 & ~x26 & ~x31 & ~x32 & ~x40 & ~x52 & ~x83 & ~x420 & ~x450 & ~x451 & ~x453 & ~x455 & ~x479 & ~x480 & ~x508 & ~x509 & ~x536 & ~x539 & ~x564 & ~x567 & ~x586 & ~x588 & ~x590 & ~x591 & ~x616 & ~x621 & ~x625 & ~x670 & ~x672 & ~x674 & ~x678 & ~x723 & ~x725 & ~x729 & ~x736 & ~x757 & ~x760 & ~x761;
assign c5485 =  x527 & ~x168 & ~x383 & ~x396 & ~x760;
assign c5487 = ~x95 & ~x363 & ~x391 & ~x434 & ~x445 & ~x471 & ~x576 & ~x632 & ~x716;
assign c5489 =  x264 & ~x83 & ~x350 & ~x375 & ~x403 & ~x508 & ~x733;
assign c5491 =  x491 &  x684 & ~x75 & ~x756 & ~x783;
assign c5493 =  x517 & ~x104 & ~x105 & ~x130 & ~x353 & ~x404;
assign c5495 =  x737 & ~x26 & ~x453;
assign c5497 = ~x28 & ~x85 & ~x275 & ~x297 & ~x414 & ~x493 & ~x636 & ~x673 & ~x733 & ~x746 & ~x771;
assign c5499 =  x231 &  x488 & ~x109 & ~x696 & ~x751 & ~x760;
assign c60 =  x516 &  x517 & ~x2 & ~x27 & ~x54 & ~x82 & ~x85 & ~x87 & ~x106 & ~x108 & ~x111 & ~x112 & ~x114 & ~x117 & ~x136 & ~x138 & ~x139 & ~x170 & ~x196 & ~x199 & ~x200 & ~x201 & ~x218 & ~x219 & ~x224 & ~x228 & ~x230 & ~x247 & ~x255 & ~x275 & ~x277 & ~x280 & ~x283 & ~x286 & ~x302 & ~x303 & ~x310 & ~x312 & ~x339 & ~x341 & ~x342 & ~x360 & ~x362 & ~x416 & ~x417 & ~x445 & ~x470 & ~x472 & ~x500 & ~x502 & ~x504 & ~x528 & ~x536 & ~x555 & ~x558 & ~x561 & ~x562 & ~x563 & ~x582 & ~x587 & ~x588 & ~x590 & ~x608 & ~x611 & ~x614 & ~x663 & ~x690 & ~x692 & ~x695 & ~x696 & ~x703 & ~x718 & ~x726 & ~x730 & ~x745 & ~x750 & ~x753 & ~x756 & ~x760 & ~x773;
assign c62 =  x638 & ~x25 & ~x55 & ~x84 & ~x111 & ~x113 & ~x138 & ~x139 & ~x140 & ~x142 & ~x167 & ~x168 & ~x170 & ~x197 & ~x224 & ~x225 & ~x671 & ~x749 & ~x776 & ~x783;
assign c64 =  x414 & ~x65 & ~x167 & ~x251 & ~x355 & ~x391 & ~x776;
assign c66 =  x464 & ~x3 & ~x4 & ~x5 & ~x19 & ~x22 & ~x25 & ~x26 & ~x27 & ~x28 & ~x29 & ~x30 & ~x34 & ~x53 & ~x68 & ~x69 & ~x80 & ~x81 & ~x82 & ~x84 & ~x85 & ~x86 & ~x87 & ~x110 & ~x112 & ~x114 & ~x137 & ~x141 & ~x165 & ~x168 & ~x195 & ~x197 & ~x225 & ~x252 & ~x336 & ~x377 & ~x403 & ~x404 & ~x643 & ~x699 & ~x700 & ~x727 & ~x753 & ~x754 & ~x756 & ~x780 & ~x781 & ~x783;
assign c68 =  x514 &  x550 & ~x0 & ~x2 & ~x25 & ~x27 & ~x28 & ~x30 & ~x53 & ~x58 & ~x84 & ~x86 & ~x89 & ~x90 & ~x111 & ~x139 & ~x141 & ~x143 & ~x197 & ~x252 & ~x354 & ~x588 & ~x701 & ~x748 & ~x755 & ~x775;
assign c610 = ~x1 & ~x23 & ~x50 & ~x58 & ~x83 & ~x108 & ~x115 & ~x140 & ~x142 & ~x170 & ~x172 & ~x190 & ~x218 & ~x219 & ~x220 & ~x221 & ~x224 & ~x227 & ~x229 & ~x238 & ~x247 & ~x248 & ~x251 & ~x252 & ~x255 & ~x256 & ~x278 & ~x283 & ~x312 & ~x313 & ~x359 & ~x364 & ~x367 & ~x378 & ~x388 & ~x390 & ~x391 & ~x417 & ~x422 & ~x425 & ~x450 & ~x451 & ~x508 & ~x610 & ~x639 & ~x642 & ~x669 & ~x700 & ~x701 & ~x745 & ~x753 & ~x771 & ~x782;
assign c612 =  x185 & ~x23 & ~x25 & ~x53 & ~x81 & ~x83 & ~x105 & ~x106 & ~x108 & ~x110 & ~x115 & ~x162 & ~x170 & ~x173 & ~x189 & ~x190 & ~x197 & ~x204 & ~x217 & ~x222 & ~x223 & ~x224 & ~x247 & ~x250 & ~x254 & ~x275 & ~x277 & ~x278 & ~x305 & ~x309 & ~x331 & ~x340 & ~x341 & ~x390 & ~x421 & ~x425 & ~x444 & ~x445 & ~x450 & ~x468 & ~x477 & ~x479 & ~x499 & ~x509 & ~x512 & ~x532 & ~x538 & ~x554 & ~x556 & ~x562 & ~x583 & ~x590 & ~x591 & ~x594 & ~x611 & ~x617 & ~x670 & ~x676 & ~x677 & ~x703 & ~x705 & ~x753 & ~x755 & ~x760 & ~x783;
assign c614 =  x185 & ~x1 & ~x2 & ~x3 & ~x15 & ~x22 & ~x25 & ~x26 & ~x27 & ~x28 & ~x32 & ~x49 & ~x50 & ~x51 & ~x52 & ~x54 & ~x56 & ~x58 & ~x59 & ~x60 & ~x78 & ~x79 & ~x80 & ~x83 & ~x85 & ~x88 & ~x106 & ~x107 & ~x108 & ~x110 & ~x112 & ~x113 & ~x115 & ~x137 & ~x139 & ~x141 & ~x165 & ~x168 & ~x171 & ~x189 & ~x190 & ~x194 & ~x195 & ~x199 & ~x200 & ~x220 & ~x221 & ~x222 & ~x225 & ~x226 & ~x228 & ~x248 & ~x249 & ~x251 & ~x253 & ~x254 & ~x255 & ~x277 & ~x280 & ~x282 & ~x306 & ~x308 & ~x333 & ~x334 & ~x335 & ~x337 & ~x340 & ~x362 & ~x364 & ~x366 & ~x395 & ~x417 & ~x418 & ~x420 & ~x445 & ~x448 & ~x449 & ~x450 & ~x474 & ~x475 & ~x500 & ~x501 & ~x502 & ~x504 & ~x529 & ~x530 & ~x541 & ~x556 & ~x558 & ~x559 & ~x560 & ~x564 & ~x586 & ~x587 & ~x588 & ~x591 & ~x612 & ~x613 & ~x618 & ~x638 & ~x639 & ~x641 & ~x643 & ~x644 & ~x667 & ~x669 & ~x671 & ~x672 & ~x673 & ~x675 & ~x697 & ~x700 & ~x726 & ~x729 & ~x753 & ~x754 & ~x756 & ~x758 & ~x759 & ~x762 & ~x780 & ~x781 & ~x783;
assign c616 =  x462 &  x605 & ~x6 & ~x21 & ~x25 & ~x27 & ~x29 & ~x35 & ~x51 & ~x53 & ~x54 & ~x57 & ~x62 & ~x78 & ~x79 & ~x80 & ~x81 & ~x83 & ~x84 & ~x106 & ~x107 & ~x108 & ~x109 & ~x110 & ~x112 & ~x133 & ~x134 & ~x135 & ~x136 & ~x137 & ~x138 & ~x139 & ~x140 & ~x141 & ~x163 & ~x164 & ~x165 & ~x166 & ~x167 & ~x168 & ~x192 & ~x193 & ~x194 & ~x195 & ~x220 & ~x221 & ~x224 & ~x225 & ~x226 & ~x251 & ~x253 & ~x277 & ~x278 & ~x281 & ~x309 & ~x335 & ~x364 & ~x365 & ~x391 & ~x392 & ~x419 & ~x447 & ~x476 & ~x503 & ~x531 & ~x532 & ~x615 & ~x642 & ~x644 & ~x671 & ~x672 & ~x728 & ~x729 & ~x748 & ~x776 & ~x777 & ~x783;
assign c618 =  x397 &  x489 & ~x28 & ~x55 & ~x82 & ~x83 & ~x92 & ~x93 & ~x112 & ~x121 & ~x148 & ~x167 & ~x195 & ~x196 & ~x251 & ~x254 & ~x392 & ~x756 & ~x757;
assign c620 =  x154 &  x574 & ~x24 & ~x103 & ~x112 & ~x274 & ~x283 & ~x393 & ~x423 & ~x449 & ~x474 & ~x504 & ~x530 & ~x533 & ~x644 & ~x650 & ~x663 & ~x694 & ~x697 & ~x756 & ~x760 & ~x781;
assign c622 =  x323 &  x519 &  x637 & ~x27 & ~x85 & ~x110 & ~x138 & ~x141 & ~x166 & ~x169 & ~x194 & ~x280 & ~x763;
assign c624 =  x124 &  x188 & ~x3 & ~x33 & ~x55 & ~x61 & ~x84 & ~x85 & ~x86 & ~x138 & ~x164 & ~x168 & ~x196 & ~x222 & ~x224 & ~x253 & ~x280 & ~x334 & ~x391 & ~x419 & ~x446 & ~x504 & ~x616 & ~x673 & ~x700 & ~x729 & ~x754 & ~x757 & ~x759;
assign c626 =  x388 &  x675;
assign c628 = ~x28 & ~x29 & ~x30 & ~x52 & ~x55 & ~x56 & ~x79 & ~x83 & ~x106 & ~x107 & ~x108 & ~x133 & ~x136 & ~x140 & ~x141 & ~x152 & ~x162 & ~x167 & ~x188 & ~x189 & ~x190 & ~x191 & ~x194 & ~x195 & ~x222 & ~x224 & ~x225 & ~x226 & ~x281 & ~x305 & ~x333 & ~x335 & ~x338 & ~x363 & ~x365 & ~x366 & ~x390 & ~x394 & ~x395 & ~x396 & ~x420 & ~x422 & ~x443 & ~x445 & ~x446 & ~x449 & ~x471 & ~x500 & ~x504 & ~x505 & ~x512 & ~x517 & ~x534 & ~x541 & ~x542 & ~x544 & ~x557 & ~x568 & ~x589 & ~x595 & ~x597 & ~x619 & ~x624 & ~x642 & ~x647 & ~x649 & ~x651 & ~x669 & ~x673 & ~x677 & ~x695 & ~x699 & ~x703 & ~x704 & ~x705 & ~x726 & ~x782;
assign c630 =  x664 &  x691 & ~x27 & ~x34 & ~x66 & ~x67 & ~x81 & ~x83 & ~x93 & ~x111 & ~x140 & ~x167 & ~x176 & ~x587 & ~x615 & ~x643 & ~x727;
assign c632 = ~x203 & ~x218 & ~x231 & ~x302 & ~x373 & ~x542 & ~x548 & ~x576 & ~x605 & ~x634 & ~x661;
assign c634 = ~x23 & ~x46 & ~x68 & ~x88 & ~x119 & ~x132 & ~x165 & ~x193 & ~x199 & ~x202 & ~x218 & ~x259 & ~x287 & ~x331 & ~x360 & ~x387 & ~x413 & ~x416 & ~x419 & ~x429 & ~x568 & ~x569 & ~x620 & ~x624 & ~x648 & ~x680 & ~x710;
assign c636 = ~x1 & ~x2 & ~x3 & ~x20 & ~x21 & ~x22 & ~x23 & ~x25 & ~x26 & ~x27 & ~x29 & ~x30 & ~x31 & ~x32 & ~x33 & ~x49 & ~x50 & ~x53 & ~x55 & ~x56 & ~x57 & ~x58 & ~x59 & ~x77 & ~x78 & ~x80 & ~x82 & ~x83 & ~x86 & ~x87 & ~x89 & ~x106 & ~x107 & ~x110 & ~x111 & ~x112 & ~x113 & ~x115 & ~x132 & ~x133 & ~x135 & ~x136 & ~x137 & ~x140 & ~x143 & ~x144 & ~x151 & ~x152 & ~x160 & ~x161 & ~x163 & ~x164 & ~x165 & ~x166 & ~x167 & ~x168 & ~x171 & ~x172 & ~x188 & ~x189 & ~x193 & ~x194 & ~x195 & ~x196 & ~x197 & ~x198 & ~x199 & ~x200 & ~x216 & ~x217 & ~x218 & ~x220 & ~x222 & ~x224 & ~x225 & ~x226 & ~x227 & ~x228 & ~x244 & ~x245 & ~x246 & ~x247 & ~x249 & ~x251 & ~x252 & ~x253 & ~x254 & ~x255 & ~x273 & ~x274 & ~x275 & ~x276 & ~x277 & ~x278 & ~x279 & ~x280 & ~x281 & ~x283 & ~x303 & ~x304 & ~x305 & ~x306 & ~x308 & ~x309 & ~x310 & ~x311 & ~x313 & ~x332 & ~x333 & ~x334 & ~x335 & ~x337 & ~x338 & ~x339 & ~x340 & ~x361 & ~x362 & ~x363 & ~x364 & ~x366 & ~x367 & ~x368 & ~x389 & ~x390 & ~x391 & ~x392 & ~x393 & ~x394 & ~x395 & ~x397 & ~x416 & ~x417 & ~x418 & ~x421 & ~x422 & ~x424 & ~x446 & ~x447 & ~x448 & ~x450 & ~x471 & ~x472 & ~x475 & ~x476 & ~x501 & ~x503 & ~x504 & ~x505 & ~x525 & ~x528 & ~x530 & ~x531 & ~x532 & ~x535 & ~x538 & ~x540 & ~x554 & ~x555 & ~x557 & ~x558 & ~x559 & ~x560 & ~x562 & ~x567 & ~x569 & ~x583 & ~x584 & ~x585 & ~x586 & ~x587 & ~x589 & ~x596 & ~x597 & ~x609 & ~x610 & ~x611 & ~x612 & ~x614 & ~x615 & ~x616 & ~x617 & ~x618 & ~x619 & ~x620 & ~x625 & ~x638 & ~x639 & ~x640 & ~x641 & ~x642 & ~x643 & ~x644 & ~x646 & ~x647 & ~x650 & ~x652 & ~x653 & ~x665 & ~x667 & ~x668 & ~x670 & ~x671 & ~x672 & ~x673 & ~x674 & ~x675 & ~x676 & ~x677 & ~x679 & ~x680 & ~x693 & ~x694 & ~x695 & ~x696 & ~x697 & ~x698 & ~x699 & ~x700 & ~x701 & ~x702 & ~x704 & ~x705 & ~x708 & ~x722 & ~x724 & ~x725 & ~x726 & ~x727 & ~x728 & ~x729 & ~x730 & ~x731 & ~x733 & ~x734 & ~x736 & ~x751 & ~x755 & ~x756 & ~x757 & ~x758 & ~x759 & ~x763 & ~x778 & ~x779 & ~x780 & ~x781 & ~x782 & ~x783;
assign c638 = ~x125 & ~x133 & ~x188 & ~x246 & ~x312 & ~x313 & ~x333 & ~x462 & ~x480 & ~x569 & ~x625 & ~x653;
assign c640 =  x600 &  x601 &  x627 &  x628 &  x629 &  x679 & ~x24 & ~x29 & ~x53 & ~x55 & ~x56 & ~x59 & ~x83 & ~x85 & ~x86 & ~x113 & ~x139 & ~x168 & ~x197 & ~x225 & ~x252 & ~x254 & ~x281 & ~x391 & ~x644 & ~x699 & ~x727 & ~x730 & ~x755 & ~x783;
assign c642 =  x338 &  x366 &  x394;
assign c644 =  x395 &  x515 & ~x25 & ~x167;
assign c646 =  x14 &  x42 &  x576 &  x604 & ~x1 & ~x2 & ~x26 & ~x28 & ~x29 & ~x30 & ~x37 & ~x54 & ~x56 & ~x57 & ~x64 & ~x80 & ~x81 & ~x82 & ~x83 & ~x86 & ~x110 & ~x111 & ~x138 & ~x140 & ~x166 & ~x167 & ~x168 & ~x169 & ~x170 & ~x171 & ~x195 & ~x196 & ~x225 & ~x252 & ~x253 & ~x279 & ~x282 & ~x308 & ~x309 & ~x335 & ~x363 & ~x364 & ~x366 & ~x421 & ~x445 & ~x446 & ~x448 & ~x473 & ~x475 & ~x501 & ~x504 & ~x529 & ~x531 & ~x532 & ~x557 & ~x558 & ~x560 & ~x586 & ~x587 & ~x589 & ~x617 & ~x669 & ~x672 & ~x673 & ~x698 & ~x699 & ~x700 & ~x702 & ~x725 & ~x726 & ~x729 & ~x755 & ~x781 & ~x782 & ~x783;
assign c648 =  x356 &  x601 & ~x1 & ~x27 & ~x57 & ~x67 & ~x85 & ~x94 & ~x95 & ~x110 & ~x111 & ~x113 & ~x142 & ~x222 & ~x278 & ~x282 & ~x308 & ~x389 & ~x422 & ~x447 & ~x473 & ~x475 & ~x557 & ~x559 & ~x560 & ~x614 & ~x618 & ~x640 & ~x673 & ~x699 & ~x702 & ~x728 & ~x756 & ~x781 & ~x782;
assign c650 =  x367 &  x395 &  x489 & ~x24 & ~x112 & ~x195 & ~x735 & ~x756 & ~x764;
assign c652 =  x464 &  x556 & ~x63 & ~x90;
assign c654 =  x179 &  x551 & ~x2 & ~x25 & ~x26 & ~x66 & ~x67 & ~x94 & ~x111 & ~x112 & ~x113 & ~x121 & ~x141 & ~x167 & ~x252 & ~x308 & ~x336 & ~x364 & ~x392 & ~x532 & ~x756 & ~x762 & ~x782;
assign c656 =  x505 &  x590;
assign c658 =  x663 & ~x0 & ~x5 & ~x23 & ~x25 & ~x26 & ~x30 & ~x32 & ~x57 & ~x85 & ~x108 & ~x110 & ~x140 & ~x165 & ~x168 & ~x193 & ~x221 & ~x226 & ~x250 & ~x308 & ~x335 & ~x337 & ~x363 & ~x393 & ~x432 & ~x440 & ~x441 & ~x559 & ~x560 & ~x586 & ~x614 & ~x616 & ~x644 & ~x756 & ~x757;
assign c660 =  x368 &  x489 & ~x55 & ~x63 & ~x91 & ~x109 & ~x118 & ~x196 & ~x224 & ~x308 & ~x756 & ~x757 & ~x783;
assign c662 = ~x112 & ~x134 & ~x144 & ~x151 & ~x161 & ~x162 & ~x188 & ~x194 & ~x208 & ~x209 & ~x216 & ~x228 & ~x311 & ~x394 & ~x396 & ~x418 & ~x444 & ~x511 & ~x561 & ~x597 & ~x642 & ~x652 & ~x653 & ~x679 & ~x698 & ~x749;
assign c664 =  x294 &  x434 &  x462 &  x544 & ~x6 & ~x26 & ~x28 & ~x33 & ~x54 & ~x58 & ~x80 & ~x82 & ~x87 & ~x114 & ~x139 & ~x168 & ~x195 & ~x226 & ~x253 & ~x254 & ~x465 & ~x503 & ~x556 & ~x558 & ~x560 & ~x587 & ~x616 & ~x618 & ~x645 & ~x671 & ~x755 & ~x758;
assign c666 =  x602 &  x684 &  x711 & ~x26 & ~x58 & ~x139 & ~x140 & ~x141 & ~x142 & ~x253 & ~x305 & ~x339 & ~x390 & ~x499 & ~x505 & ~x554 & ~x557 & ~x582 & ~x584 & ~x644 & ~x757 & ~x758 & ~x783;
assign c668 =  x408 &  x609 & ~x110 & ~x112 & ~x252;
assign c670 =  x333 &  x527 &  x554;
assign c672 = ~x31 & ~x51 & ~x53 & ~x54 & ~x57 & ~x59 & ~x79 & ~x80 & ~x111 & ~x113 & ~x114 & ~x115 & ~x139 & ~x144 & ~x168 & ~x169 & ~x191 & ~x195 & ~x197 & ~x200 & ~x226 & ~x248 & ~x250 & ~x255 & ~x276 & ~x278 & ~x281 & ~x284 & ~x306 & ~x310 & ~x312 & ~x313 & ~x330 & ~x331 & ~x337 & ~x367 & ~x389 & ~x391 & ~x393 & ~x397 & ~x398 & ~x408 & ~x416 & ~x419 & ~x421 & ~x427 & ~x430 & ~x440 & ~x452 & ~x453 & ~x469 & ~x471 & ~x476 & ~x478 & ~x481 & ~x482 & ~x499 & ~x526 & ~x531 & ~x534 & ~x535 & ~x553 & ~x561 & ~x565 & ~x581 & ~x587 & ~x588 & ~x590 & ~x611 & ~x668 & ~x670 & ~x699 & ~x702 & ~x705 & ~x717 & ~x754 & ~x756 & ~x760 & ~x762;
assign c674 =  x479 &  x507 &  x563 &  x647;
assign c676 = ~x11 & ~x38 & ~x39 & ~x53 & ~x83 & ~x138 & ~x167 & ~x198 & ~x220 & ~x221 & ~x222 & ~x223 & ~x307 & ~x362 & ~x364 & ~x366 & ~x420 & ~x425 & ~x452 & ~x458 & ~x461 & ~x470 & ~x477 & ~x481 & ~x489 & ~x495 & ~x551 & ~x563 & ~x586 & ~x590 & ~x610 & ~x611 & ~x644 & ~x647 & ~x770;
assign c678 =  x129 & ~x61 & ~x106 & ~x108 & ~x111 & ~x134 & ~x140 & ~x141 & ~x163 & ~x165 & ~x210 & ~x221 & ~x222 & ~x252 & ~x253 & ~x279 & ~x280 & ~x306 & ~x307 & ~x309 & ~x475 & ~x560 & ~x587 & ~x616 & ~x716 & ~x729 & ~x744 & ~x770 & ~x782;
assign c680 =  x271 & ~x33 & ~x52 & ~x57 & ~x115 & ~x139 & ~x143 & ~x165 & ~x194 & ~x197 & ~x225 & ~x227 & ~x228 & ~x279 & ~x282 & ~x284 & ~x311 & ~x313 & ~x314 & ~x335 & ~x336 & ~x339 & ~x366 & ~x367 & ~x394 & ~x395 & ~x397 & ~x399 & ~x412 & ~x418 & ~x419 & ~x420 & ~x422 & ~x425 & ~x426 & ~x443 & ~x446 & ~x451 & ~x472 & ~x474 & ~x481 & ~x502 & ~x525 & ~x528 & ~x532 & ~x555 & ~x559 & ~x589 & ~x591 & ~x610 & ~x615 & ~x640 & ~x643 & ~x668 & ~x670 & ~x672 & ~x698 & ~x699 & ~x700 & ~x702 & ~x726 & ~x779;
assign c682 =  x130 &  x605 & ~x27 & ~x28 & ~x54 & ~x61 & ~x80 & ~x83 & ~x84 & ~x108 & ~x109 & ~x137 & ~x138 & ~x140 & ~x249 & ~x252 & ~x254 & ~x278 & ~x307 & ~x391 & ~x418 & ~x419 & ~x474 & ~x501 & ~x589 & ~x644 & ~x671 & ~x702 & ~x728 & ~x730 & ~x758 & ~x759 & ~x769 & ~x783;
assign c684 =  x435 &  x452 &  x480 & ~x106 & ~x251 & ~x253 & ~x281 & ~x559 & ~x756;
assign c686 =  x572 &  x637 &  x664 & ~x23 & ~x25 & ~x27 & ~x80 & ~x81 & ~x82 & ~x83 & ~x112 & ~x139 & ~x168 & ~x195 & ~x196 & ~x224 & ~x225 & ~x252 & ~x587 & ~x671 & ~x672 & ~x700 & ~x766;
assign c688 = ~x21 & ~x33 & ~x54 & ~x133 & ~x161 & ~x252 & ~x284 & ~x304 & ~x305 & ~x341 & ~x347 & ~x481 & ~x536 & ~x713 & ~x728 & ~x767 & ~x768 & ~x769 & ~x779;
assign c690 =  x516 &  x577 & ~x27 & ~x28 & ~x29 & ~x80 & ~x83 & ~x86 & ~x107 & ~x117 & ~x169 & ~x197 & ~x277 & ~x278 & ~x334 & ~x364 & ~x365 & ~x389 & ~x391 & ~x474 & ~x502 & ~x557 & ~x559 & ~x613 & ~x699 & ~x729 & ~x773;
assign c692 =  x352 & ~x26 & ~x53 & ~x57 & ~x77 & ~x86 & ~x106 & ~x124 & ~x138 & ~x162 & ~x190 & ~x197 & ~x226 & ~x250 & ~x252 & ~x277 & ~x337 & ~x360 & ~x422 & ~x506 & ~x554 & ~x568 & ~x569 & ~x700 & ~x701 & ~x751 & ~x758 & ~x779;
assign c694 =  x354 & ~x2 & ~x3 & ~x30 & ~x56 & ~x58 & ~x61 & ~x78 & ~x83 & ~x86 & ~x88 & ~x107 & ~x109 & ~x113 & ~x115 & ~x135 & ~x137 & ~x162 & ~x166 & ~x167 & ~x170 & ~x171 & ~x190 & ~x191 & ~x194 & ~x218 & ~x224 & ~x226 & ~x246 & ~x253 & ~x254 & ~x276 & ~x283 & ~x285 & ~x311 & ~x313 & ~x332 & ~x338 & ~x390 & ~x392 & ~x422 & ~x444 & ~x446 & ~x454 & ~x473 & ~x476 & ~x477 & ~x483 & ~x498 & ~x499 & ~x501 & ~x531 & ~x532 & ~x536 & ~x557 & ~x560 & ~x567 & ~x588 & ~x594 & ~x595 & ~x611 & ~x620 & ~x621 & ~x624 & ~x640 & ~x642 & ~x645 & ~x648 & ~x667 & ~x672 & ~x699 & ~x705 & ~x706 & ~x727 & ~x728 & ~x730 & ~x759 & ~x783;
assign c696 = ~x8 & ~x87 & ~x102 & ~x110 & ~x118 & ~x130 & ~x133 & ~x141 & ~x160 & ~x165 & ~x167 & ~x190 & ~x194 & ~x199 & ~x220 & ~x225 & ~x281 & ~x332 & ~x367 & ~x390 & ~x415 & ~x418 & ~x425 & ~x444 & ~x453 & ~x458 & ~x484 & ~x486 & ~x488 & ~x494 & ~x500 & ~x504 & ~x506 & ~x522 & ~x523 & ~x536 & ~x538 & ~x556 & ~x564 & ~x668 & ~x674 & ~x722 & ~x727 & ~x752 & ~x756;
assign c698 =  x367 &  x417 & ~x386;
assign c6100 = ~x21 & ~x48 & ~x49 & ~x56 & ~x84 & ~x131 & ~x135 & ~x140 & ~x169 & ~x170 & ~x196 & ~x197 & ~x213 & ~x219 & ~x223 & ~x224 & ~x225 & ~x229 & ~x248 & ~x280 & ~x284 & ~x305 & ~x310 & ~x313 & ~x339 & ~x340 & ~x359 & ~x387 & ~x389 & ~x394 & ~x418 & ~x427 & ~x455 & ~x457 & ~x477 & ~x483 & ~x501 & ~x506 & ~x531 & ~x577 & ~x587 & ~x605 & ~x611 & ~x621 & ~x622 & ~x633 & ~x664 & ~x674 & ~x695 & ~x697 & ~x705 & ~x728 & ~x729 & ~x773;
assign c6102 =  x501 &  x556 &  x637;
assign c6104 =  x720 & ~x35 & ~x61 & ~x80 & ~x81 & ~x82 & ~x109 & ~x123 & ~x138 & ~x195 & ~x504 & ~x643 & ~x728 & ~x762;
assign c6106 =  x70 &  x154 &  x182 &  x266 &  x351 &  x407 &  x463 &  x491 & ~x169 & ~x253 & ~x308 & ~x474 & ~x475 & ~x588 & ~x616 & ~x648 & ~x676 & ~x783;
assign c6108 =  x425 &  x453 & ~x0 & ~x26 & ~x29 & ~x53 & ~x54 & ~x56 & ~x80 & ~x82 & ~x83 & ~x85 & ~x112 & ~x135 & ~x136 & ~x137 & ~x139 & ~x142 & ~x162 & ~x165 & ~x166 & ~x192 & ~x197 & ~x198 & ~x223 & ~x225 & ~x226 & ~x251 & ~x278 & ~x281 & ~x308 & ~x335 & ~x363 & ~x419 & ~x475 & ~x477 & ~x504 & ~x532 & ~x533 & ~x560 & ~x561 & ~x589 & ~x644 & ~x645 & ~x700 & ~x749 & ~x777;
assign c6110 =  x298 &  x575 & ~x2 & ~x5 & ~x33 & ~x54 & ~x85 & ~x86 & ~x97 & ~x107 & ~x108 & ~x110 & ~x137 & ~x138 & ~x144 & ~x163 & ~x172 & ~x191 & ~x221 & ~x248 & ~x254 & ~x284 & ~x304 & ~x305 & ~x310 & ~x311 & ~x312 & ~x359 & ~x368 & ~x394 & ~x417 & ~x420 & ~x447 & ~x450 & ~x452 & ~x476 & ~x505 & ~x528 & ~x530 & ~x555 & ~x558 & ~x559 & ~x584 & ~x590 & ~x614 & ~x673 & ~x700 & ~x732 & ~x759;
assign c6112 =  x211 &  x239 &  x295 &  x379 &  x491 &  x631 &  x687 & ~x86 & ~x110 & ~x138 & ~x278 & ~x280 & ~x307 & ~x310 & ~x335 & ~x367 & ~x394 & ~x525 & ~x530 & ~x532 & ~x534 & ~x536 & ~x551 & ~x555 & ~x580 & ~x585 & ~x592 & ~x595 & ~x783;
assign c6114 =  x235 &  x326 & ~x53 & ~x59 & ~x87 & ~x109 & ~x111 & ~x136 & ~x141 & ~x165 & ~x168 & ~x193 & ~x223 & ~x228 & ~x254 & ~x279 & ~x280 & ~x282 & ~x310 & ~x313 & ~x314 & ~x335 & ~x363 & ~x395 & ~x425 & ~x448 & ~x471 & ~x472 & ~x473 & ~x475 & ~x479 & ~x511 & ~x525 & ~x535 & ~x537 & ~x538 & ~x539 & ~x554 & ~x562 & ~x564 & ~x583 & ~x611 & ~x613 & ~x616 & ~x648 & ~x670 & ~x698 & ~x755 & ~x782;
assign c6116 = ~x10 & ~x11 & ~x53 & ~x54 & ~x55 & ~x56 & ~x76 & ~x80 & ~x84 & ~x89 & ~x91 & ~x108 & ~x118 & ~x135 & ~x146 & ~x173 & ~x196 & ~x203 & ~x221 & ~x223 & ~x229 & ~x250 & ~x252 & ~x259 & ~x275 & ~x288 & ~x309 & ~x329 & ~x331 & ~x334 & ~x339 & ~x341 & ~x343 & ~x361 & ~x364 & ~x384 & ~x387 & ~x392 & ~x416 & ~x417 & ~x419 & ~x420 & ~x426 & ~x446 & ~x447 & ~x451 & ~x454 & ~x479 & ~x480 & ~x525 & ~x532 & ~x535 & ~x559 & ~x580 & ~x586 & ~x588 & ~x605 & ~x609 & ~x611 & ~x615 & ~x616 & ~x638 & ~x671 & ~x695 & ~x700 & ~x701 & ~x717 & ~x735 & ~x752 & ~x757 & ~x758 & ~x762 & ~x763 & ~x772 & ~x778 & ~x780;
assign c6118 =  x324 &  x661 & ~x58 & ~x87 & ~x111 & ~x139 & ~x141 & ~x143 & ~x195 & ~x196 & ~x197 & ~x223 & ~x309 & ~x311 & ~x341 & ~x364 & ~x389 & ~x391 & ~x396 & ~x424 & ~x452 & ~x497 & ~x532 & ~x537 & ~x540 & ~x564 & ~x566 & ~x568 & ~x612 & ~x613 & ~x618 & ~x639 & ~x668 & ~x708 & ~x725 & ~x730 & ~x754 & ~x761 & ~x779;
assign c6120 = ~x1 & ~x23 & ~x53 & ~x55 & ~x82 & ~x83 & ~x114 & ~x142 & ~x143 & ~x192 & ~x197 & ~x199 & ~x223 & ~x228 & ~x252 & ~x253 & ~x256 & ~x257 & ~x258 & ~x307 & ~x308 & ~x313 & ~x342 & ~x389 & ~x393 & ~x447 & ~x450 & ~x451 & ~x508 & ~x560 & ~x561 & ~x565 & ~x581 & ~x589 & ~x620 & ~x630 & ~x658 & ~x675 & ~x684 & ~x699 & ~x702 & ~x712 & ~x726 & ~x747 & ~x749 & ~x757 & ~x758 & ~x780;
assign c6122 = ~x4 & ~x9 & ~x19 & ~x23 & ~x24 & ~x31 & ~x33 & ~x62 & ~x78 & ~x83 & ~x90 & ~x102 & ~x105 & ~x111 & ~x114 & ~x131 & ~x132 & ~x137 & ~x139 & ~x141 & ~x145 & ~x161 & ~x166 & ~x171 & ~x188 & ~x189 & ~x190 & ~x193 & ~x201 & ~x221 & ~x222 & ~x246 & ~x256 & ~x271 & ~x273 & ~x275 & ~x303 & ~x313 & ~x358 & ~x367 & ~x368 & ~x383 & ~x387 & ~x388 & ~x395 & ~x419 & ~x424 & ~x442 & ~x473 & ~x499 & ~x506 & ~x507 & ~x535 & ~x537 & ~x540 & ~x556 & ~x560 & ~x584 & ~x586 & ~x593 & ~x598 & ~x609 & ~x617 & ~x624 & ~x626 & ~x634 & ~x642 & ~x645 & ~x653 & ~x662 & ~x665 & ~x666 & ~x670 & ~x678 & ~x698 & ~x722 & ~x731 & ~x735 & ~x762 & ~x763 & ~x780 & ~x783;
assign c6124 = ~x22 & ~x76 & ~x105 & ~x135 & ~x148 & ~x161 & ~x188 & ~x217 & ~x260 & ~x261 & ~x262 & ~x313 & ~x340 & ~x559 & ~x605 & ~x653 & ~x690 & ~x744;
assign c6126 =  x291 &  x602 &  x629 &  x630 & ~x27 & ~x28 & ~x32 & ~x56 & ~x59 & ~x60 & ~x78 & ~x108 & ~x110 & ~x113 & ~x140 & ~x142 & ~x163 & ~x191 & ~x218 & ~x221 & ~x227 & ~x248 & ~x276 & ~x277 & ~x282 & ~x283 & ~x310 & ~x333 & ~x340 & ~x363 & ~x393 & ~x396 & ~x424 & ~x470 & ~x500 & ~x501 & ~x526 & ~x527 & ~x564 & ~x581 & ~x582 & ~x583 & ~x590 & ~x593 & ~x610 & ~x615 & ~x618 & ~x642 & ~x645 & ~x647 & ~x725 & ~x727 & ~x732 & ~x758 & ~x761 & ~x762 & ~x775;
assign c6128 =  x244 & ~x25 & ~x38 & ~x108 & ~x137 & ~x139 & ~x167 & ~x194 & ~x223 & ~x224 & ~x253 & ~x257 & ~x276 & ~x278 & ~x279 & ~x280 & ~x281 & ~x282 & ~x283 & ~x284 & ~x336 & ~x338 & ~x340 & ~x363 & ~x419 & ~x440 & ~x445 & ~x451 & ~x508 & ~x534 & ~x586 & ~x591 & ~x643 & ~x648 & ~x676 & ~x705 & ~x729 & ~x754 & ~x755 & ~x757 & ~x759;
assign c6130 =  x602 &  x658 &  x683 & ~x3 & ~x25 & ~x30 & ~x32 & ~x51 & ~x56 & ~x57 & ~x59 & ~x110 & ~x112 & ~x114 & ~x136 & ~x138 & ~x139 & ~x165 & ~x191 & ~x225 & ~x250 & ~x332 & ~x333 & ~x335 & ~x392 & ~x421 & ~x422 & ~x423 & ~x447 & ~x474 & ~x476 & ~x478 & ~x480 & ~x499 & ~x500 & ~x508 & ~x528 & ~x532 & ~x533 & ~x558 & ~x588 & ~x639 & ~x645 & ~x673 & ~x699;
assign c6132 =  x599 &  x627 &  x636 & ~x26 & ~x27 & ~x28 & ~x29 & ~x34 & ~x53 & ~x63 & ~x82 & ~x83 & ~x89 & ~x90 & ~x112 & ~x168 & ~x196 & ~x224 & ~x252 & ~x280 & ~x765;
assign c6134 =  x606 &  x663 & ~x22 & ~x24 & ~x25 & ~x26 & ~x30 & ~x59 & ~x109 & ~x140 & ~x168 & ~x196 & ~x197 & ~x252 & ~x253 & ~x475 & ~x531 & ~x532 & ~x587 & ~x588 & ~x615 & ~x672 & ~x698 & ~x699 & ~x729 & ~x756 & ~x757 & ~x783;
assign c6136 =  x571 &  x636 & ~x3 & ~x37 & ~x62 & ~x111 & ~x120 & ~x139 & ~x140 & ~x147 & ~x224 & ~x776 & ~x783;
assign c6138 =  x505 & ~x482 & ~x778;
assign c6140 =  x433 &  x461 & ~x27 & ~x33 & ~x61 & ~x62 & ~x80 & ~x82 & ~x86 & ~x110 & ~x118 & ~x135 & ~x140 & ~x169 & ~x171 & ~x202 & ~x223 & ~x225 & ~x256 & ~x257 & ~x258 & ~x278 & ~x282 & ~x285 & ~x304 & ~x305 & ~x310 & ~x314 & ~x336 & ~x339 & ~x342 & ~x362 & ~x393 & ~x419 & ~x442 & ~x444 & ~x471 & ~x472 & ~x479 & ~x505 & ~x506 & ~x525 & ~x529 & ~x557 & ~x562 & ~x579 & ~x611 & ~x633 & ~x637 & ~x641 & ~x645 & ~x661 & ~x670 & ~x671 & ~x689 & ~x702 & ~x716 & ~x745 & ~x755 & ~x776 & ~x779 & ~x781;
assign c6142 =  x394 &  x534 &  x590;
assign c6144 =  x238 &  x547 &  x603 &  x687 & ~x3 & ~x26 & ~x57 & ~x82 & ~x86 & ~x113 & ~x144 & ~x166 & ~x191 & ~x219 & ~x254 & ~x255 & ~x282 & ~x307 & ~x338 & ~x340 & ~x341 & ~x451 & ~x470 & ~x476 & ~x504 & ~x527 & ~x538 & ~x563 & ~x581 & ~x584 & ~x593 & ~x608 & ~x609 & ~x611 & ~x640 & ~x697 & ~x727;
assign c6146 =  x562 & ~x399 & ~x454;
assign c6148 = ~x1 & ~x27 & ~x28 & ~x51 & ~x53 & ~x56 & ~x78 & ~x96 & ~x124 & ~x162 & ~x190 & ~x192 & ~x225 & ~x227 & ~x247 & ~x252 & ~x285 & ~x311 & ~x313 & ~x417 & ~x421 & ~x444 & ~x476 & ~x479 & ~x486 & ~x488 & ~x498 & ~x514 & ~x557 & ~x566 & ~x569 & ~x586 & ~x587 & ~x589 & ~x592 & ~x595 & ~x725 & ~x728 & ~x731 & ~x759;
assign c6150 =  x552 & ~x0 & ~x24 & ~x40 & ~x53 & ~x56 & ~x81 & ~x83 & ~x110 & ~x138 & ~x141 & ~x254 & ~x281 & ~x335 & ~x336 & ~x363 & ~x391 & ~x392 & ~x446 & ~x473 & ~x475 & ~x529 & ~x530 & ~x531 & ~x559 & ~x588 & ~x615 & ~x652 & ~x681 & ~x700 & ~x701 & ~x708 & ~x709 & ~x728 & ~x736 & ~x754 & ~x755 & ~x779;
assign c6152 =  x464 &  x528 & ~x83 & ~x357 & ~x385;
assign c6154 =  x544 & ~x1 & ~x32 & ~x54 & ~x69 & ~x108 & ~x112 & ~x165 & ~x195 & ~x260 & ~x376 & ~x401 & ~x728 & ~x775 & ~x777;
assign c6156 =  x434 &  x581 & ~x0 & ~x4 & ~x5 & ~x25 & ~x34 & ~x51 & ~x53 & ~x55 & ~x62 & ~x81 & ~x82 & ~x109 & ~x110 & ~x112 & ~x139 & ~x140 & ~x195 & ~x196 & ~x252 & ~x503 & ~x700 & ~x734 & ~x756 & ~x757 & ~x763 & ~x764 & ~x783;
assign c6158 =  x461 &  x489 & ~x2 & ~x5 & ~x6 & ~x11 & ~x20 & ~x21 & ~x22 & ~x23 & ~x24 & ~x25 & ~x26 & ~x50 & ~x51 & ~x54 & ~x55 & ~x58 & ~x60 & ~x77 & ~x80 & ~x82 & ~x83 & ~x85 & ~x87 & ~x105 & ~x106 & ~x107 & ~x112 & ~x113 & ~x115 & ~x133 & ~x134 & ~x135 & ~x136 & ~x138 & ~x140 & ~x141 & ~x142 & ~x163 & ~x165 & ~x167 & ~x198 & ~x218 & ~x219 & ~x223 & ~x227 & ~x229 & ~x254 & ~x255 & ~x258 & ~x310 & ~x333 & ~x335 & ~x339 & ~x360 & ~x365 & ~x366 & ~x389 & ~x394 & ~x416 & ~x418 & ~x419 & ~x420 & ~x421 & ~x422 & ~x447 & ~x448 & ~x476 & ~x477 & ~x479 & ~x502 & ~x526 & ~x527 & ~x529 & ~x531 & ~x532 & ~x534 & ~x554 & ~x555 & ~x556 & ~x559 & ~x561 & ~x562 & ~x563 & ~x581 & ~x585 & ~x586 & ~x613 & ~x619 & ~x633 & ~x639 & ~x644 & ~x673 & ~x693 & ~x695 & ~x696 & ~x699 & ~x702 & ~x724 & ~x746 & ~x747 & ~x757 & ~x763 & ~x774 & ~x782;
assign c6160 =  x458 &  x522 & ~x21 & ~x24 & ~x25 & ~x29 & ~x35 & ~x53 & ~x56 & ~x58 & ~x62 & ~x81 & ~x111 & ~x112 & ~x118 & ~x137 & ~x139 & ~x140 & ~x141 & ~x194 & ~x195 & ~x197 & ~x224 & ~x280 & ~x363 & ~x474 & ~x502 & ~x616 & ~x707 & ~x728 & ~x729 & ~x735 & ~x757 & ~x783;
assign c6162 =  x674;
assign c6164 = ~x8 & ~x24 & ~x53 & ~x54 & ~x60 & ~x80 & ~x81 & ~x83 & ~x89 & ~x108 & ~x110 & ~x111 & ~x112 & ~x139 & ~x162 & ~x168 & ~x195 & ~x198 & ~x221 & ~x231 & ~x256 & ~x257 & ~x280 & ~x301 & ~x303 & ~x304 & ~x331 & ~x334 & ~x338 & ~x339 & ~x341 & ~x386 & ~x390 & ~x392 & ~x394 & ~x396 & ~x407 & ~x408 & ~x414 & ~x419 & ~x426 & ~x442 & ~x446 & ~x473 & ~x479 & ~x500 & ~x584 & ~x594 & ~x611 & ~x613 & ~x616 & ~x621 & ~x633 & ~x641 & ~x662 & ~x732 & ~x733 & ~x762;
assign c6166 =  x70 &  x433 &  x461 & ~x1 & ~x3 & ~x5 & ~x26 & ~x30 & ~x33 & ~x52 & ~x56 & ~x61 & ~x81 & ~x108 & ~x144 & ~x164 & ~x167 & ~x169 & ~x198 & ~x223 & ~x225 & ~x251 & ~x280 & ~x308 & ~x362 & ~x391 & ~x419 & ~x475 & ~x501 & ~x559 & ~x644 & ~x663 & ~x717 & ~x724 & ~x725 & ~x744 & ~x745 & ~x757 & ~x760;
assign c6168 =  x517 & ~x195 & ~x255 & ~x402 & ~x429 & ~x431 & ~x439 & ~x502 & ~x685 & ~x739;
assign c6170 =  x185 & ~x1 & ~x2 & ~x6 & ~x20 & ~x21 & ~x26 & ~x49 & ~x53 & ~x54 & ~x57 & ~x77 & ~x84 & ~x106 & ~x109 & ~x110 & ~x113 & ~x134 & ~x136 & ~x137 & ~x139 & ~x161 & ~x164 & ~x165 & ~x189 & ~x190 & ~x197 & ~x198 & ~x217 & ~x218 & ~x220 & ~x222 & ~x226 & ~x248 & ~x251 & ~x254 & ~x279 & ~x280 & ~x287 & ~x306 & ~x333 & ~x337 & ~x364 & ~x370 & ~x391 & ~x448 & ~x475 & ~x476 & ~x483 & ~x501 & ~x532 & ~x538 & ~x554 & ~x558 & ~x560 & ~x567 & ~x584 & ~x594 & ~x595 & ~x612 & ~x622 & ~x624 & ~x639 & ~x641 & ~x643 & ~x648 & ~x672 & ~x679 & ~x681 & ~x696 & ~x698 & ~x703 & ~x706 & ~x723 & ~x724 & ~x725 & ~x727 & ~x728 & ~x729 & ~x734 & ~x752 & ~x753 & ~x754 & ~x762 & ~x781;
assign c6172 =  x152 &  x266 & ~x27 & ~x110 & ~x137 & ~x196 & ~x197 & ~x250 & ~x335 & ~x336 & ~x343 & ~x344 & ~x361 & ~x363 & ~x370 & ~x375 & ~x392 & ~x399 & ~x401 & ~x418 & ~x470 & ~x474 & ~x479 & ~x500 & ~x501 & ~x508 & ~x526 & ~x528 & ~x533 & ~x555 & ~x560 & ~x563 & ~x586 & ~x640 & ~x695 & ~x697 & ~x758 & ~x782;
assign c6174 =  x547 &  x637 &  x666 & ~x1 & ~x2 & ~x26 & ~x27 & ~x28 & ~x30 & ~x52 & ~x56 & ~x58 & ~x63 & ~x80 & ~x82 & ~x84 & ~x86 & ~x90 & ~x114 & ~x139 & ~x140 & ~x168 & ~x196 & ~x281 & ~x308 & ~x336 & ~x532 & ~x671 & ~x672 & ~x700 & ~x756;
assign c6176 =  x572 &  x573 &  x637 & ~x3 & ~x4 & ~x26 & ~x27 & ~x28 & ~x32 & ~x63 & ~x64 & ~x82 & ~x110 & ~x111 & ~x137 & ~x138 & ~x140 & ~x195 & ~x559 & ~x756 & ~x765;
assign c6178 =  x350 &  x494 &  x582 & ~x144 & ~x224;
assign c6180 =  x263 &  x434 & ~x25 & ~x33 & ~x58 & ~x87 & ~x94 & ~x95 & ~x108 & ~x122 & ~x131 & ~x132 & ~x141 & ~x250 & ~x304 & ~x334 & ~x339 & ~x390 & ~x419 & ~x502 & ~x552 & ~x580 & ~x608 & ~x617 & ~x726 & ~x759;
assign c6182 =  x434 &  x542 &  x578 & ~x25 & ~x27 & ~x54 & ~x67 & ~x79 & ~x80 & ~x82 & ~x84 & ~x111 & ~x138 & ~x140 & ~x196 & ~x756 & ~x761;
assign c6184 =  x562 &  x618 &  x646 & ~x106 & ~x166 & ~x195 & ~x735 & ~x751 & ~x762;
assign c6186 =  x178 &  x604 & ~x17 & ~x19 & ~x25 & ~x27 & ~x28 & ~x51 & ~x108 & ~x111 & ~x136 & ~x163 & ~x165 & ~x166 & ~x195 & ~x200 & ~x249 & ~x252 & ~x257 & ~x280 & ~x308 & ~x361 & ~x390 & ~x438 & ~x446 & ~x671 & ~x728 & ~x730 & ~x754 & ~x758;
assign c6188 =  x589 & ~x454;
assign c6190 = ~x1 & ~x79 & ~x82 & ~x85 & ~x108 & ~x154 & ~x169 & ~x172 & ~x247 & ~x255 & ~x283 & ~x323 & ~x334 & ~x360 & ~x393 & ~x449 & ~x478 & ~x482 & ~x499 & ~x556 & ~x588 & ~x593 & ~x616 & ~x725;
assign c6192 =  x685 &  x738 &  x739 & ~x1 & ~x26 & ~x29 & ~x30 & ~x81 & ~x85 & ~x108 & ~x113 & ~x136 & ~x139 & ~x141 & ~x164 & ~x167 & ~x194 & ~x195 & ~x252 & ~x253 & ~x254 & ~x278 & ~x281 & ~x363 & ~x366 & ~x391 & ~x392 & ~x416 & ~x417 & ~x419 & ~x472 & ~x474 & ~x499 & ~x500 & ~x501 & ~x502 & ~x503 & ~x506 & ~x525 & ~x529 & ~x531 & ~x536 & ~x560 & ~x565 & ~x585 & ~x590 & ~x616 & ~x618 & ~x619 & ~x641 & ~x644 & ~x645 & ~x671 & ~x672 & ~x673 & ~x700 & ~x730 & ~x755 & ~x756 & ~x759;
assign c6194 = ~x176 & ~x204 & ~x218 & ~x228 & ~x261 & ~x280 & ~x344 & ~x374 & ~x391 & ~x569 & ~x596 & ~x599 & ~x652 & ~x653 & ~x696 & ~x706 & ~x708 & ~x746 & ~x752;
assign c6196 =  x573 & ~x0 & ~x11 & ~x22 & ~x24 & ~x26 & ~x28 & ~x39 & ~x50 & ~x53 & ~x56 & ~x60 & ~x67 & ~x108 & ~x110 & ~x112 & ~x113 & ~x136 & ~x169 & ~x193 & ~x196 & ~x199 & ~x200 & ~x219 & ~x221 & ~x224 & ~x247 & ~x249 & ~x310 & ~x332 & ~x334 & ~x363 & ~x366 & ~x390 & ~x391 & ~x420 & ~x422 & ~x431 & ~x450 & ~x459 & ~x474 & ~x501 & ~x557 & ~x616 & ~x697 & ~x757;
assign c6198 =  x219 &  x322 &  x350 & ~x167 & ~x223 & ~x642;
assign c6200 = ~x19 & ~x22 & ~x29 & ~x31 & ~x48 & ~x51 & ~x62 & ~x104 & ~x112 & ~x115 & ~x136 & ~x159 & ~x164 & ~x166 & ~x169 & ~x188 & ~x192 & ~x218 & ~x223 & ~x226 & ~x247 & ~x254 & ~x274 & ~x276 & ~x277 & ~x278 & ~x284 & ~x312 & ~x313 & ~x341 & ~x359 & ~x366 & ~x368 & ~x387 & ~x389 & ~x396 & ~x418 & ~x478 & ~x498 & ~x525 & ~x536 & ~x561 & ~x572 & ~x583 & ~x586 & ~x592 & ~x594 & ~x596 & ~x599 & ~x600 & ~x607 & ~x608 & ~x610 & ~x613 & ~x619 & ~x623 & ~x624 & ~x635 & ~x637 & ~x644 & ~x646 & ~x653 & ~x663 & ~x670 & ~x672 & ~x673 & ~x699 & ~x706 & ~x726 & ~x751 & ~x755 & ~x758 & ~x760 & ~x764;
assign c6202 =  x658 & ~x1 & ~x26 & ~x29 & ~x30 & ~x56 & ~x57 & ~x81 & ~x85 & ~x86 & ~x109 & ~x114 & ~x115 & ~x133 & ~x139 & ~x140 & ~x161 & ~x166 & ~x189 & ~x195 & ~x199 & ~x221 & ~x226 & ~x227 & ~x247 & ~x248 & ~x274 & ~x278 & ~x335 & ~x337 & ~x338 & ~x340 & ~x362 & ~x363 & ~x366 & ~x367 & ~x388 & ~x390 & ~x393 & ~x417 & ~x420 & ~x450 & ~x479 & ~x480 & ~x496 & ~x500 & ~x501 & ~x502 & ~x511 & ~x512 & ~x513 & ~x514 & ~x515 & ~x516 & ~x523 & ~x524 & ~x525 & ~x527 & ~x531 & ~x538 & ~x541 & ~x550 & ~x552 & ~x559 & ~x562 & ~x563 & ~x566 & ~x567 & ~x583 & ~x585 & ~x592 & ~x620 & ~x621 & ~x637 & ~x642 & ~x643 & ~x669 & ~x696 & ~x697 & ~x698 & ~x701 & ~x703 & ~x705 & ~x729 & ~x762;
assign c6204 =  x323 &  x489 &  x578 &  x579 &  x606 & ~x224;
assign c6206 =  x488 & ~x4 & ~x23 & ~x24 & ~x57 & ~x60 & ~x85 & ~x107 & ~x141 & ~x164 & ~x168 & ~x173 & ~x200 & ~x201 & ~x276 & ~x281 & ~x308 & ~x363 & ~x381 & ~x390 & ~x557 & ~x560 & ~x615 & ~x662 & ~x690 & ~x717 & ~x719 & ~x745 & ~x746 & ~x750 & ~x774;
assign c6208 = ~x39 & ~x53 & ~x54 & ~x58 & ~x80 & ~x82 & ~x106 & ~x115 & ~x164 & ~x166 & ~x170 & ~x191 & ~x225 & ~x227 & ~x257 & ~x276 & ~x281 & ~x284 & ~x313 & ~x314 & ~x334 & ~x396 & ~x398 & ~x416 & ~x417 & ~x432 & ~x433 & ~x442 & ~x444 & ~x453 & ~x461 & ~x468 & ~x476 & ~x477 & ~x494 & ~x511 & ~x513 & ~x514 & ~x525 & ~x564 & ~x640 & ~x672 & ~x703 & ~x705 & ~x729 & ~x730 & ~x753 & ~x759;
assign c6210 =  x489 &  x552 & ~x1 & ~x23 & ~x28 & ~x38 & ~x54 & ~x57 & ~x81 & ~x85 & ~x138 & ~x165 & ~x167 & ~x748 & ~x782;
assign c6212 =  x240 &  x633 & ~x5 & ~x21 & ~x61 & ~x110 & ~x141 & ~x168 & ~x252 & ~x283 & ~x306 & ~x312 & ~x334 & ~x340 & ~x365 & ~x445 & ~x512 & ~x528 & ~x531 & ~x539 & ~x596 & ~x610 & ~x651 & ~x673 & ~x762;
assign c6214 =  x152 & ~x1 & ~x6 & ~x24 & ~x25 & ~x27 & ~x29 & ~x30 & ~x31 & ~x34 & ~x37 & ~x52 & ~x54 & ~x55 & ~x58 & ~x60 & ~x66 & ~x79 & ~x83 & ~x84 & ~x85 & ~x86 & ~x87 & ~x89 & ~x90 & ~x93 & ~x112 & ~x113 & ~x116 & ~x117 & ~x138 & ~x139 & ~x143 & ~x168 & ~x170 & ~x173 & ~x194 & ~x195 & ~x196 & ~x197 & ~x223 & ~x224 & ~x225 & ~x226 & ~x251 & ~x279 & ~x280 & ~x282 & ~x307 & ~x308 & ~x335 & ~x363 & ~x364 & ~x381 & ~x382 & ~x391 & ~x392 & ~x419 & ~x476 & ~x499 & ~x501 & ~x503 & ~x504 & ~x531 & ~x532 & ~x588 & ~x589 & ~x617 & ~x645 & ~x646 & ~x671 & ~x673 & ~x674 & ~x675 & ~x702 & ~x704 & ~x730 & ~x731 & ~x732 & ~x756 & ~x757 & ~x759 & ~x760 & ~x761 & ~x776 & ~x777;
assign c6216 = ~x90 & ~x104 & ~x113 & ~x147 & ~x159 & ~x171 & ~x192 & ~x195 & ~x231 & ~x246 & ~x315 & ~x317 & ~x395 & ~x397 & ~x473 & ~x484 & ~x529 & ~x558 & ~x568 & ~x570 & ~x592 & ~x605 & ~x614 & ~x615 & ~x622 & ~x624 & ~x625 & ~x695 & ~x727 & ~x760;
assign c6218 =  x664 & ~x0 & ~x27 & ~x35 & ~x53 & ~x54 & ~x55 & ~x56 & ~x57 & ~x78 & ~x80 & ~x84 & ~x85 & ~x107 & ~x110 & ~x114 & ~x139 & ~x165 & ~x166 & ~x167 & ~x170 & ~x194 & ~x197 & ~x251 & ~x252 & ~x282 & ~x308 & ~x336 & ~x363 & ~x431 & ~x440 & ~x476 & ~x671 & ~x699 & ~x700 & ~x728 & ~x729;
assign c6220 =  x647 & ~x223 & ~x400 & ~x594 & ~x696 & ~x707 & ~x735;
assign c6222 =  x459 &  x497 &  x525 &  x552 &  x553 & ~x64 & ~x91 & ~x92 & ~x168;
assign c6224 = ~x55 & ~x77 & ~x79 & ~x82 & ~x114 & ~x115 & ~x134 & ~x141 & ~x164 & ~x224 & ~x229 & ~x250 & ~x257 & ~x337 & ~x370 & ~x387 & ~x389 & ~x391 & ~x396 & ~x418 & ~x422 & ~x441 & ~x464 & ~x528 & ~x530 & ~x534 & ~x586 & ~x587 & ~x615 & ~x622 & ~x638 & ~x660 & ~x673 & ~x675 & ~x688 & ~x695 & ~x707 & ~x715 & ~x743;
assign c6226 =  x551 & ~x330 & ~x357 & ~x734;
assign c6228 = ~x1 & ~x20 & ~x59 & ~x84 & ~x87 & ~x107 & ~x141 & ~x162 & ~x165 & ~x200 & ~x219 & ~x225 & ~x275 & ~x276 & ~x318 & ~x335 & ~x347 & ~x352 & ~x423 & ~x443 & ~x448 & ~x470 & ~x472 & ~x473 & ~x502 & ~x554 & ~x585 & ~x611 & ~x725 & ~x730 & ~x745 & ~x747 & ~x754 & ~x755 & ~x776 & ~x782;
assign c6230 =  x239 &  x267 &  x324 & ~x0 & ~x104 & ~x139 & ~x193 & ~x197 & ~x250 & ~x254 & ~x279 & ~x285 & ~x339 & ~x366 & ~x395 & ~x420 & ~x421 & ~x424 & ~x466 & ~x494 & ~x495 & ~x507 & ~x512 & ~x594;
assign c6232 =  x102 &  x103 &  x632 &  x661 & ~x281 & ~x448 & ~x758;
assign c6234 =  x351 & ~x3 & ~x5 & ~x28 & ~x130 & ~x169 & ~x192 & ~x217 & ~x246 & ~x255 & ~x340 & ~x499 & ~x503 & ~x508 & ~x514 & ~x523 & ~x540 & ~x542 & ~x543 & ~x544 & ~x550 & ~x551 & ~x552 & ~x564 & ~x615 & ~x676;
assign c6236 = ~x3 & ~x7 & ~x20 & ~x21 & ~x23 & ~x26 & ~x31 & ~x35 & ~x48 & ~x57 & ~x60 & ~x62 & ~x77 & ~x89 & ~x91 & ~x92 & ~x106 & ~x107 & ~x108 & ~x120 & ~x132 & ~x135 & ~x137 & ~x144 & ~x146 & ~x161 & ~x162 & ~x189 & ~x199 & ~x200 & ~x202 & ~x224 & ~x249 & ~x251 & ~x273 & ~x275 & ~x276 & ~x303 & ~x306 & ~x307 & ~x312 & ~x313 & ~x340 & ~x368 & ~x386 & ~x387 & ~x397 & ~x421 & ~x423 & ~x426 & ~x447 & ~x448 & ~x451 & ~x455 & ~x474 & ~x483 & ~x497 & ~x498 & ~x499 & ~x500 & ~x508 & ~x510 & ~x531 & ~x534 & ~x535 & ~x538 & ~x555 & ~x558 & ~x562 & ~x564 & ~x565 & ~x569 & ~x590 & ~x595 & ~x600 & ~x611 & ~x619 & ~x635 & ~x639 & ~x643 & ~x652 & ~x665 & ~x676 & ~x680 & ~x701 & ~x707 & ~x708 & ~x730 & ~x731 & ~x760 & ~x761;
assign c6238 =  x523 & ~x21 & ~x51 & ~x58 & ~x81 & ~x83 & ~x109 & ~x138 & ~x383 & ~x652 & ~x681 & ~x724 & ~x728 & ~x765 & ~x782;
assign c6240 =  x296 &  x632 & ~x108 & ~x113 & ~x312 & ~x313 & ~x364 & ~x415 & ~x488 & ~x489 & ~x495 & ~x499 & ~x512 & ~x513 & ~x528 & ~x729;
assign c6242 =  x688 & ~x25 & ~x30 & ~x74 & ~x83 & ~x88 & ~x106 & ~x136 & ~x143 & ~x196 & ~x221 & ~x249 & ~x254 & ~x276 & ~x279 & ~x310 & ~x360 & ~x362 & ~x390 & ~x424 & ~x482 & ~x483 & ~x503 & ~x513 & ~x516 & ~x524 & ~x529 & ~x559 & ~x565 & ~x581 & ~x582 & ~x609 & ~x668 & ~x724 & ~x752 & ~x760;
assign c6244 =  x156 &  x606 & ~x54 & ~x112 & ~x168 & ~x252 & ~x263 & ~x307 & ~x308 & ~x335 & ~x363 & ~x440;
assign c6246 =  x206 &  x350 &  x574 &  x603 & ~x23 & ~x24 & ~x26 & ~x52 & ~x55 & ~x56 & ~x80 & ~x85 & ~x110 & ~x142 & ~x197 & ~x222 & ~x225 & ~x251 & ~x252 & ~x281 & ~x282 & ~x307 & ~x335 & ~x362 & ~x363 & ~x364 & ~x366 & ~x389 & ~x390 & ~x417 & ~x418 & ~x419 & ~x446 & ~x450 & ~x475 & ~x562 & ~x586 & ~x587 & ~x588 & ~x589 & ~x611 & ~x614 & ~x615 & ~x669 & ~x672 & ~x701 & ~x729 & ~x781;
assign c6248 = ~x0 & ~x22 & ~x28 & ~x85 & ~x106 & ~x108 & ~x112 & ~x115 & ~x134 & ~x168 & ~x171 & ~x173 & ~x190 & ~x198 & ~x223 & ~x246 & ~x278 & ~x309 & ~x311 & ~x334 & ~x337 & ~x363 & ~x368 & ~x388 & ~x393 & ~x449 & ~x473 & ~x477 & ~x478 & ~x501 & ~x503 & ~x537 & ~x566 & ~x588 & ~x590 & ~x591 & ~x603 & ~x639 & ~x640 & ~x668 & ~x670 & ~x672 & ~x673 & ~x688 & ~x725 & ~x750 & ~x752 & ~x753 & ~x771;
assign c6250 = ~x22 & ~x26 & ~x27 & ~x29 & ~x31 & ~x33 & ~x34 & ~x52 & ~x61 & ~x82 & ~x86 & ~x87 & ~x88 & ~x107 & ~x112 & ~x141 & ~x143 & ~x169 & ~x197 & ~x219 & ~x221 & ~x224 & ~x258 & ~x260 & ~x276 & ~x277 & ~x278 & ~x286 & ~x308 & ~x311 & ~x316 & ~x333 & ~x337 & ~x340 & ~x342 & ~x361 & ~x368 & ~x369 & ~x386 & ~x388 & ~x389 & ~x390 & ~x394 & ~x397 & ~x416 & ~x418 & ~x442 & ~x447 & ~x452 & ~x454 & ~x470 & ~x472 & ~x475 & ~x535 & ~x555 & ~x563 & ~x582 & ~x585 & ~x609 & ~x611 & ~x619 & ~x639 & ~x645 & ~x667 & ~x670 & ~x672 & ~x675 & ~x686 & ~x698 & ~x701 & ~x714 & ~x741 & ~x752 & ~x761 & ~x767 & ~x781;
assign c6252 =  x211 &  x547 &  x631 & ~x5 & ~x16 & ~x52 & ~x53 & ~x80 & ~x277 & ~x285 & ~x342 & ~x391 & ~x419 & ~x421 & ~x482 & ~x537 & ~x552 & ~x564 & ~x618 & ~x645 & ~x733 & ~x734 & ~x752 & ~x777;
assign c6254 =  x544 & ~x2 & ~x6 & ~x7 & ~x20 & ~x25 & ~x30 & ~x32 & ~x33 & ~x35 & ~x43 & ~x51 & ~x54 & ~x55 & ~x56 & ~x57 & ~x59 & ~x62 & ~x71 & ~x79 & ~x80 & ~x81 & ~x106 & ~x109 & ~x111 & ~x113 & ~x115 & ~x137 & ~x165 & ~x166 & ~x167 & ~x168 & ~x223 & ~x252 & ~x336 & ~x429 & ~x504 & ~x588 & ~x615 & ~x670 & ~x671 & ~x699 & ~x728 & ~x729 & ~x763 & ~x774 & ~x783;
assign c6256 =  x186 &  x214 & ~x0 & ~x23 & ~x32 & ~x54 & ~x58 & ~x61 & ~x86 & ~x87 & ~x88 & ~x114 & ~x115 & ~x134 & ~x139 & ~x164 & ~x170 & ~x173 & ~x195 & ~x198 & ~x199 & ~x200 & ~x219 & ~x223 & ~x224 & ~x248 & ~x250 & ~x255 & ~x256 & ~x257 & ~x274 & ~x276 & ~x278 & ~x285 & ~x308 & ~x310 & ~x331 & ~x338 & ~x339 & ~x361 & ~x366 & ~x367 & ~x393 & ~x413 & ~x419 & ~x481 & ~x506 & ~x528 & ~x529 & ~x537 & ~x557 & ~x559 & ~x562 & ~x588 & ~x589 & ~x591 & ~x617 & ~x618 & ~x641 & ~x645 & ~x648 & ~x650 & ~x667 & ~x672 & ~x675 & ~x679 & ~x699 & ~x700 & ~x701 & ~x729 & ~x732 & ~x733 & ~x759 & ~x760 & ~x762;
assign c6258 =  x233 &  x237 & ~x50 & ~x57 & ~x79 & ~x110 & ~x141 & ~x172 & ~x224 & ~x256 & ~x285 & ~x364 & ~x471 & ~x473 & ~x508 & ~x531 & ~x533 & ~x555 & ~x557 & ~x560 & ~x565 & ~x620 & ~x703 & ~x780;
assign c6260 = ~x19 & ~x52 & ~x72 & ~x86 & ~x111 & ~x117 & ~x165 & ~x171 & ~x201 & ~x254 & ~x281 & ~x313 & ~x387 & ~x389 & ~x401 & ~x430 & ~x437 & ~x438 & ~x445 & ~x458 & ~x473 & ~x475 & ~x477 & ~x478 & ~x501 & ~x536 & ~x560 & ~x582 & ~x586 & ~x611 & ~x618 & ~x698 & ~x729 & ~x757;
assign c6262 =  x240 &  x268 &  x660 & ~x188 & ~x282 & ~x419 & ~x506 & ~x526 & ~x533 & ~x567 & ~x751;
assign c6264 =  x183 &  x211 &  x239 &  x323 &  x351 & ~x76 & ~x80 & ~x101 & ~x103 & ~x108 & ~x140 & ~x280 & ~x335 & ~x339 & ~x445 & ~x474 & ~x503 & ~x523 & ~x526 & ~x556 & ~x566 & ~x595 & ~x618 & ~x667 & ~x701;
assign c6266 =  x658 & ~x4 & ~x194 & ~x304 & ~x390 & ~x480 & ~x512 & ~x516 & ~x517 & ~x572 & ~x586 & ~x598 & ~x642 & ~x652 & ~x727 & ~x736 & ~x783;
assign c6268 =  x490 &  x609 & ~x0 & ~x24 & ~x27 & ~x34 & ~x52 & ~x53 & ~x56 & ~x57 & ~x64 & ~x79 & ~x81 & ~x87 & ~x91 & ~x108 & ~x109 & ~x167 & ~x195 & ~x224 & ~x252 & ~x756 & ~x764;
assign c6270 =  x293 &  x656 & ~x142 & ~x482 & ~x521 & ~x641 & ~x780;
assign c6272 =  x155 &  x211 & ~x26 & ~x32 & ~x61 & ~x79 & ~x103 & ~x159 & ~x193 & ~x259 & ~x308 & ~x314 & ~x336 & ~x363 & ~x397 & ~x499 & ~x505 & ~x510 & ~x513 & ~x524 & ~x746;
assign c6274 =  x69 &  x350 &  x406 &  x490 & ~x60 & ~x163 & ~x168 & ~x219 & ~x220 & ~x252 & ~x255 & ~x282 & ~x306 & ~x363 & ~x391 & ~x422 & ~x473 & ~x537 & ~x612 & ~x643 & ~x701 & ~x703 & ~x719 & ~x758;
assign c6276 =  x445 &  x473 &  x638;
assign c6278 =  x240 &  x605 & ~x26 & ~x52 & ~x53 & ~x54 & ~x55 & ~x56 & ~x79 & ~x81 & ~x82 & ~x85 & ~x107 & ~x110 & ~x112 & ~x137 & ~x141 & ~x163 & ~x165 & ~x166 & ~x168 & ~x169 & ~x192 & ~x195 & ~x220 & ~x222 & ~x225 & ~x250 & ~x251 & ~x252 & ~x253 & ~x255 & ~x278 & ~x279 & ~x280 & ~x281 & ~x283 & ~x285 & ~x306 & ~x309 & ~x312 & ~x338 & ~x364 & ~x367 & ~x391 & ~x392 & ~x417 & ~x419 & ~x420 & ~x421 & ~x422 & ~x448 & ~x449 & ~x450 & ~x470 & ~x472 & ~x473 & ~x475 & ~x483 & ~x498 & ~x502 & ~x505 & ~x506 & ~x509 & ~x526 & ~x527 & ~x528 & ~x537 & ~x538 & ~x553 & ~x555 & ~x556 & ~x557 & ~x558 & ~x559 & ~x589 & ~x592 & ~x614 & ~x618 & ~x639 & ~x641 & ~x642 & ~x647 & ~x668 & ~x674 & ~x676 & ~x698 & ~x725 & ~x731 & ~x733 & ~x753 & ~x758 & ~x760 & ~x762 & ~x780 & ~x783;
assign c6280 = ~x8 & ~x15 & ~x24 & ~x43 & ~x71 & ~x89 & ~x163 & ~x281 & ~x364 & ~x367 & ~x393 & ~x394 & ~x422 & ~x424 & ~x425 & ~x449 & ~x472 & ~x502 & ~x510 & ~x563 & ~x581 & ~x593 & ~x621 & ~x623 & ~x668 & ~x698 & ~x730;
assign c6282 =  x184 & ~x2 & ~x3 & ~x25 & ~x28 & ~x30 & ~x49 & ~x51 & ~x53 & ~x82 & ~x112 & ~x113 & ~x138 & ~x142 & ~x189 & ~x190 & ~x200 & ~x201 & ~x217 & ~x219 & ~x225 & ~x252 & ~x253 & ~x279 & ~x280 & ~x308 & ~x312 & ~x331 & ~x334 & ~x337 & ~x363 & ~x396 & ~x418 & ~x453 & ~x470 & ~x478 & ~x527 & ~x529 & ~x531 & ~x536 & ~x541 & ~x565 & ~x566 & ~x567 & ~x568 & ~x573 & ~x587 & ~x610 & ~x613 & ~x620 & ~x637 & ~x644 & ~x670 & ~x674 & ~x702 & ~x727 & ~x755;
assign c6284 = ~x2 & ~x30 & ~x33 & ~x89 & ~x132 & ~x171 & ~x218 & ~x256 & ~x258 & ~x310 & ~x312 & ~x444 & ~x474 & ~x479 & ~x581 & ~x585 & ~x605 & ~x612 & ~x715 & ~x725 & ~x756 & ~x758;
assign c6286 =  x301 & ~x21 & ~x22 & ~x27 & ~x30 & ~x51 & ~x54 & ~x56 & ~x58 & ~x65 & ~x66 & ~x81 & ~x82 & ~x84 & ~x86 & ~x108 & ~x109 & ~x111 & ~x113 & ~x121 & ~x137 & ~x141 & ~x167 & ~x168 & ~x169 & ~x225 & ~x252 & ~x253 & ~x254 & ~x279 & ~x280 & ~x305 & ~x306 & ~x307 & ~x308 & ~x309 & ~x333 & ~x334 & ~x335 & ~x336 & ~x337 & ~x361 & ~x365 & ~x390 & ~x392 & ~x418 & ~x421 & ~x475 & ~x502 & ~x504 & ~x532 & ~x559 & ~x560 & ~x590 & ~x615 & ~x617 & ~x673 & ~x698 & ~x730 & ~x756 & ~x758;
assign c6288 =  x394 &  x562;
assign c6290 =  x239 &  x265 &  x350 &  x406 & ~x32 & ~x225 & ~x252 & ~x391 & ~x502 & ~x531 & ~x700 & ~x747 & ~x749 & ~x774 & ~x775 & ~x776 & ~x777;
assign c6292 =  x75 &  x551 & ~x0 & ~x1 & ~x23 & ~x25 & ~x28 & ~x113 & ~x114 & ~x142 & ~x166 & ~x197 & ~x253 & ~x254 & ~x280 & ~x335 & ~x392 & ~x418 & ~x528 & ~x531 & ~x583 & ~x584 & ~x612 & ~x617 & ~x645 & ~x696 & ~x756 & ~x758 & ~x759 & ~x783;
assign c6294 =  x577 &  x633 & ~x0 & ~x25 & ~x29 & ~x40 & ~x53 & ~x56 & ~x66 & ~x106 & ~x112 & ~x114 & ~x138 & ~x139 & ~x140 & ~x169 & ~x191 & ~x221 & ~x306 & ~x334 & ~x362 & ~x418 & ~x449 & ~x474 & ~x615 & ~x698 & ~x729 & ~x732;
assign c6296 =  x204 &  x321 & ~x0 & ~x1 & ~x5 & ~x7 & ~x24 & ~x25 & ~x26 & ~x28 & ~x29 & ~x35 & ~x55 & ~x56 & ~x58 & ~x60 & ~x61 & ~x84 & ~x85 & ~x112 & ~x114 & ~x117 & ~x139 & ~x140 & ~x142 & ~x169 & ~x196 & ~x197 & ~x224 & ~x280 & ~x307 & ~x335 & ~x337 & ~x363 & ~x588 & ~x704 & ~x728 & ~x730 & ~x733 & ~x759 & ~x782 & ~x783;
assign c6298 = ~x52 & ~x79 & ~x162 & ~x189 & ~x190 & ~x277 & ~x285 & ~x303 & ~x311 & ~x316 & ~x369 & ~x397 & ~x450 & ~x455 & ~x483 & ~x499 & ~x505 & ~x509 & ~x512 & ~x515 & ~x548 & ~x554 & ~x568 & ~x596 & ~x645 & ~x647 & ~x676 & ~x725 & ~x730 & ~x773;
assign c6300 =  x546 &  x573 & ~x4 & ~x25 & ~x54 & ~x79 & ~x82 & ~x84 & ~x87 & ~x110 & ~x111 & ~x112 & ~x113 & ~x140 & ~x167 & ~x168 & ~x196 & ~x197 & ~x278 & ~x308 & ~x316 & ~x402 & ~x404 & ~x431 & ~x440 & ~x476 & ~x560 & ~x697 & ~x700 & ~x725 & ~x726 & ~x755 & ~x781;
assign c6302 =  x571 &  x572 &  x599 & ~x2 & ~x6 & ~x59 & ~x109 & ~x112 & ~x116 & ~x140 & ~x142 & ~x167 & ~x169 & ~x170 & ~x196 & ~x197 & ~x222 & ~x224 & ~x226 & ~x227 & ~x248 & ~x254 & ~x276 & ~x283 & ~x362 & ~x390 & ~x392 & ~x411 & ~x419 & ~x420 & ~x438 & ~x449 & ~x456 & ~x457 & ~x466 & ~x467 & ~x474 & ~x477 & ~x483 & ~x533 & ~x558 & ~x561 & ~x585 & ~x586 & ~x589 & ~x616 & ~x643 & ~x756 & ~x757 & ~x759;
assign c6304 = ~x0 & ~x92 & ~x137 & ~x148 & ~x165 & ~x166 & ~x168 & ~x197 & ~x224 & ~x237 & ~x250 & ~x262 & ~x289 & ~x290 & ~x344 & ~x345 & ~x348 & ~x623 & ~x667 & ~x679 & ~x697 & ~x698 & ~x725 & ~x726 & ~x753 & ~x761 & ~x779 & ~x781 & ~x782;
assign c6306 =  x493 &  x637 & ~x66 & ~x92 & ~x119 & ~x782;
assign c6308 = ~x1 & ~x3 & ~x8 & ~x32 & ~x50 & ~x58 & ~x81 & ~x103 & ~x109 & ~x135 & ~x139 & ~x141 & ~x160 & ~x166 & ~x172 & ~x187 & ~x189 & ~x195 & ~x199 & ~x217 & ~x226 & ~x228 & ~x246 & ~x253 & ~x260 & ~x281 & ~x283 & ~x303 & ~x305 & ~x313 & ~x314 & ~x315 & ~x336 & ~x363 & ~x372 & ~x400 & ~x418 & ~x454 & ~x457 & ~x471 & ~x475 & ~x484 & ~x508 & ~x512 & ~x525 & ~x528 & ~x536 & ~x551 & ~x561 & ~x568 & ~x570 & ~x580 & ~x582 & ~x583 & ~x585 & ~x597 & ~x598 & ~x609 & ~x634 & ~x640 & ~x663 & ~x666 & ~x669 & ~x693 & ~x709 & ~x724 & ~x751 & ~x764;
assign c6310 =  x489 &  x609 & ~x40 & ~x94 & ~x121 & ~x149 & ~x176;
assign c6312 =  x294 &  x574 &  x602 &  x657 &  x658 & ~x169 & ~x197 & ~x285 & ~x366 & ~x367 & ~x395 & ~x396 & ~x423 & ~x498 & ~x507 & ~x528 & ~x537 & ~x559 & ~x584 & ~x593;
assign c6314 =  x601 &  x629 &  x655 &  x657 & ~x26 & ~x111 & ~x172 & ~x192 & ~x223 & ~x226 & ~x228 & ~x249 & ~x255 & ~x279 & ~x307 & ~x338 & ~x339 & ~x340 & ~x396 & ~x416 & ~x446 & ~x472 & ~x473 & ~x478 & ~x482 & ~x500 & ~x565 & ~x580 & ~x583 & ~x671 & ~x732 & ~x757 & ~x779 & ~x780;
assign c6316 = ~x6 & ~x19 & ~x59 & ~x106 & ~x189 & ~x203 & ~x230 & ~x248 & ~x250 & ~x260 & ~x305 & ~x308 & ~x314 & ~x317 & ~x335 & ~x424 & ~x426 & ~x541 & ~x570 & ~x591 & ~x597 & ~x604 & ~x681;
assign c6318 = ~x24 & ~x25 & ~x79 & ~x110 & ~x137 & ~x145 & ~x228 & ~x252 & ~x277 & ~x305 & ~x331 & ~x335 & ~x342 & ~x368 & ~x387 & ~x416 & ~x444 & ~x449 & ~x477 & ~x481 & ~x530 & ~x534 & ~x556 & ~x562 & ~x568 & ~x585 & ~x612 & ~x614 & ~x618 & ~x621 & ~x630 & ~x658 & ~x669 & ~x670 & ~x697 & ~x729 & ~x742 & ~x757 & ~x762 & ~x770;
assign c6320 =  x405 &  x600 &  x627 & ~x1 & ~x26 & ~x31 & ~x58 & ~x108 & ~x137 & ~x195 & ~x224 & ~x251 & ~x334 & ~x336 & ~x363 & ~x391 & ~x393 & ~x505 & ~x514 & ~x529 & ~x559 & ~x589 & ~x590 & ~x614 & ~x617 & ~x645 & ~x670 & ~x701;
assign c6322 = ~x26 & ~x29 & ~x144 & ~x145 & ~x164 & ~x190 & ~x194 & ~x201 & ~x307 & ~x342 & ~x388 & ~x415 & ~x419 & ~x482 & ~x492 & ~x513 & ~x523 & ~x561 & ~x576 & ~x620 & ~x622 & ~x632 & ~x650 & ~x669 & ~x779;
assign c6324 =  x233 &  x349 & ~x1 & ~x24 & ~x30 & ~x52 & ~x81 & ~x83 & ~x113 & ~x114 & ~x136 & ~x140 & ~x141 & ~x165 & ~x168 & ~x169 & ~x194 & ~x197 & ~x252 & ~x254 & ~x281 & ~x311 & ~x337 & ~x339 & ~x361 & ~x389 & ~x391 & ~x416 & ~x421 & ~x444 & ~x449 & ~x453 & ~x472 & ~x473 & ~x474 & ~x478 & ~x499 & ~x504 & ~x528 & ~x529 & ~x557 & ~x562 & ~x584 & ~x585 & ~x616 & ~x617 & ~x701 & ~x703 & ~x704 & ~x719 & ~x729 & ~x730 & ~x754 & ~x755 & ~x758 & ~x760 & ~x783;
assign c6326 =  x546 &  x608 & ~x52 & ~x54 & ~x82 & ~x108 & ~x137 & ~x195 & ~x196 & ~x384 & ~x735 & ~x736 & ~x764 & ~x767;
assign c6328 = ~x15 & ~x25 & ~x52 & ~x57 & ~x60 & ~x85 & ~x140 & ~x194 & ~x198 & ~x219 & ~x259 & ~x286 & ~x303 & ~x313 & ~x330 & ~x342 & ~x359 & ~x360 & ~x364 & ~x367 & ~x391 & ~x395 & ~x408 & ~x416 & ~x422 & ~x427 & ~x445 & ~x451 & ~x452 & ~x454 & ~x480 & ~x503 & ~x536 & ~x537 & ~x548 & ~x565 & ~x567 & ~x620 & ~x649 & ~x723 & ~x751 & ~x777;
assign c6330 = ~x22 & ~x25 & ~x30 & ~x53 & ~x59 & ~x79 & ~x81 & ~x106 & ~x109 & ~x110 & ~x114 & ~x137 & ~x138 & ~x140 & ~x142 & ~x145 & ~x191 & ~x192 & ~x193 & ~x201 & ~x220 & ~x222 & ~x230 & ~x246 & ~x250 & ~x255 & ~x258 & ~x275 & ~x276 & ~x281 & ~x285 & ~x307 & ~x309 & ~x311 & ~x337 & ~x338 & ~x340 & ~x371 & ~x380 & ~x389 & ~x390 & ~x397 & ~x403 & ~x413 & ~x417 & ~x418 & ~x423 & ~x427 & ~x442 & ~x443 & ~x472 & ~x478 & ~x482 & ~x501 & ~x502 & ~x526 & ~x537 & ~x554 & ~x562 & ~x563 & ~x564 & ~x565 & ~x584 & ~x588 & ~x595 & ~x610 & ~x617 & ~x619 & ~x620 & ~x638 & ~x639 & ~x646 & ~x668 & ~x671 & ~x675 & ~x697 & ~x703 & ~x722 & ~x728 & ~x730 & ~x732 & ~x733 & ~x754 & ~x779 & ~x783;
assign c6332 =  x182 &  x208 &  x434 &  x574 & ~x0 & ~x2 & ~x30 & ~x76 & ~x102 & ~x113 & ~x642 & ~x756;
assign c6334 =  x212 &  x240 &  x577 & ~x0 & ~x23 & ~x27 & ~x29 & ~x50 & ~x56 & ~x81 & ~x83 & ~x105 & ~x107 & ~x110 & ~x114 & ~x139 & ~x141 & ~x162 & ~x164 & ~x165 & ~x166 & ~x189 & ~x190 & ~x191 & ~x198 & ~x199 & ~x249 & ~x253 & ~x282 & ~x308 & ~x311 & ~x337 & ~x338 & ~x390 & ~x394 & ~x395 & ~x417 & ~x418 & ~x419 & ~x420 & ~x421 & ~x474 & ~x477 & ~x479 & ~x497 & ~x525 & ~x533 & ~x557 & ~x558 & ~x562 & ~x579 & ~x581 & ~x584 & ~x589 & ~x612 & ~x614 & ~x619 & ~x623 & ~x641 & ~x642 & ~x651 & ~x652 & ~x678 & ~x706 & ~x729;
assign c6336 =  x183 &  x323 & ~x21 & ~x139 & ~x142 & ~x143 & ~x163 & ~x169 & ~x221 & ~x254 & ~x311 & ~x337 & ~x362 & ~x418 & ~x430 & ~x431 & ~x437 & ~x446 & ~x448 & ~x467 & ~x504 & ~x559 & ~x585 & ~x673 & ~x700;
assign c6338 =  x405 & ~x9 & ~x22 & ~x23 & ~x29 & ~x37 & ~x38 & ~x52 & ~x53 & ~x56 & ~x59 & ~x85 & ~x87 & ~x91 & ~x92 & ~x109 & ~x138 & ~x171 & ~x172 & ~x195 & ~x200 & ~x251 & ~x335 & ~x353 & ~x362 & ~x363 & ~x381 & ~x503 & ~x700 & ~x720 & ~x721 & ~x746 & ~x748 & ~x758 & ~x783;
assign c6340 =  x296 &  x605 & ~x1 & ~x24 & ~x27 & ~x51 & ~x55 & ~x79 & ~x81 & ~x106 & ~x108 & ~x109 & ~x136 & ~x141 & ~x166 & ~x167 & ~x170 & ~x250 & ~x251 & ~x253 & ~x277 & ~x278 & ~x282 & ~x284 & ~x308 & ~x309 & ~x310 & ~x312 & ~x363 & ~x364 & ~x367 & ~x390 & ~x417 & ~x419 & ~x424 & ~x449 & ~x451 & ~x467 & ~x476 & ~x495 & ~x499 & ~x534 & ~x555 & ~x559 & ~x590 & ~x612 & ~x643 & ~x671 & ~x672 & ~x674 & ~x754 & ~x756 & ~x759 & ~x761;
assign c6342 =  x534 &  x674;
assign c6344 =  x211 &  x239 &  x267 &  x657 &  x684 & ~x0 & ~x28 & ~x52 & ~x56 & ~x57 & ~x82 & ~x107 & ~x137 & ~x223 & ~x279 & ~x307 & ~x336 & ~x365 & ~x419 & ~x471 & ~x472 & ~x473 & ~x502 & ~x530 & ~x584 & ~x586 & ~x588 & ~x589 & ~x616 & ~x645 & ~x701 & ~x727 & ~x754 & ~x757;
assign c6346 =  x322 &  x547 &  x658 & ~x58 & ~x130 & ~x197 & ~x366 & ~x424 & ~x448 & ~x451 & ~x469 & ~x502 & ~x536 & ~x560 & ~x645 & ~x672 & ~x725 & ~x757 & ~x760;
assign c6348 =  x462 &  x515 & ~x3 & ~x5 & ~x22 & ~x27 & ~x30 & ~x53 & ~x56 & ~x60 & ~x81 & ~x83 & ~x84 & ~x136 & ~x137 & ~x139 & ~x166 & ~x167 & ~x168 & ~x196 & ~x252 & ~x503 & ~x531 & ~x680 & ~x700 & ~x729 & ~x747 & ~x764 & ~x781 & ~x782;
assign c6350 = ~x5 & ~x111 & ~x227 & ~x258 & ~x304 & ~x309 & ~x417 & ~x426 & ~x474 & ~x604 & ~x624 & ~x695 & ~x742;
assign c6352 =  x663 & ~x0 & ~x25 & ~x27 & ~x28 & ~x96 & ~x123 & ~x137 & ~x165 & ~x166 & ~x192 & ~x193 & ~x194 & ~x196 & ~x220 & ~x221 & ~x278 & ~x305 & ~x307 & ~x363 & ~x476 & ~x560 & ~x588 & ~x616 & ~x668 & ~x698 & ~x700 & ~x726 & ~x755;
assign c6354 =  x325 &  x604 &  x689 & ~x0 & ~x3 & ~x24 & ~x82 & ~x108 & ~x167 & ~x254 & ~x277 & ~x334 & ~x336 & ~x340 & ~x418 & ~x420 & ~x445 & ~x449 & ~x504 & ~x508 & ~x511 & ~x512 & ~x536 & ~x590 & ~x639 & ~x782;
assign c6356 =  x437 &  x529;
assign c6358 = ~x2 & ~x5 & ~x8 & ~x9 & ~x37 & ~x51 & ~x52 & ~x53 & ~x78 & ~x79 & ~x105 & ~x137 & ~x145 & ~x159 & ~x169 & ~x188 & ~x217 & ~x218 & ~x223 & ~x224 & ~x225 & ~x226 & ~x228 & ~x248 & ~x249 & ~x274 & ~x285 & ~x302 & ~x306 & ~x307 & ~x310 & ~x332 & ~x333 & ~x338 & ~x339 & ~x362 & ~x364 & ~x366 & ~x473 & ~x476 & ~x477 & ~x501 & ~x504 & ~x505 & ~x523 & ~x533 & ~x554 & ~x555 & ~x556 & ~x559 & ~x560 & ~x564 & ~x566 & ~x578 & ~x582 & ~x589 & ~x593 & ~x594 & ~x610 & ~x611 & ~x612 & ~x621 & ~x642 & ~x643 & ~x647 & ~x672 & ~x677 & ~x694 & ~x695 & ~x697 & ~x715 & ~x721 & ~x723 & ~x724 & ~x727 & ~x730 & ~x732 & ~x759 & ~x770;
assign c6360 =  x442 &  x550 & ~x307 & ~x327 & ~x473;
assign c6362 = ~x4 & ~x25 & ~x28 & ~x50 & ~x53 & ~x55 & ~x110 & ~x112 & ~x132 & ~x133 & ~x141 & ~x146 & ~x150 & ~x161 & ~x163 & ~x165 & ~x169 & ~x173 & ~x195 & ~x197 & ~x219 & ~x228 & ~x229 & ~x248 & ~x257 & ~x279 & ~x285 & ~x286 & ~x329 & ~x335 & ~x336 & ~x339 & ~x342 & ~x358 & ~x363 & ~x364 & ~x418 & ~x443 & ~x444 & ~x450 & ~x481 & ~x507 & ~x511 & ~x528 & ~x535 & ~x539 & ~x564 & ~x584 & ~x586 & ~x594 & ~x606 & ~x611 & ~x615 & ~x621 & ~x623 & ~x633 & ~x637 & ~x661 & ~x671 & ~x678 & ~x690 & ~x700 & ~x704 & ~x730 & ~x732 & ~x743 & ~x748 & ~x749 & ~x762 & ~x777 & ~x779 & ~x781;
assign c6364 =  x488 &  x578 & ~x0 & ~x3 & ~x23 & ~x27 & ~x37 & ~x51 & ~x57 & ~x62 & ~x63 & ~x80 & ~x84 & ~x85 & ~x86 & ~x90 & ~x91 & ~x92 & ~x106 & ~x107 & ~x111 & ~x112 & ~x138 & ~x165 & ~x169 & ~x225 & ~x226 & ~x250 & ~x251 & ~x279 & ~x281 & ~x306 & ~x308 & ~x309 & ~x334 & ~x335 & ~x391 & ~x419 & ~x475 & ~x532 & ~x762;
assign c6366 =  x297 & ~x78 & ~x83 & ~x85 & ~x97 & ~x98 & ~x137 & ~x161 & ~x165 & ~x190 & ~x196 & ~x219 & ~x220 & ~x222 & ~x227 & ~x254 & ~x284 & ~x285 & ~x286 & ~x305 & ~x313 & ~x335 & ~x417 & ~x451 & ~x497 & ~x498 & ~x508 & ~x527 & ~x538 & ~x540 & ~x555 & ~x556 & ~x563 & ~x565 & ~x668 & ~x704 & ~x759;
assign c6368 =  x352 &  x660 & ~x24 & ~x112 & ~x123 & ~x143 & ~x168 & ~x169 & ~x196 & ~x197 & ~x281 & ~x306 & ~x333 & ~x339 & ~x364 & ~x395 & ~x416 & ~x446 & ~x447 & ~x478 & ~x529 & ~x568 & ~x587 & ~x590 & ~x616 & ~x624 & ~x645 & ~x696 & ~x697 & ~x698 & ~x726 & ~x757;
assign c6370 =  x470 &  x579 & ~x57 & ~x81 & ~x112 & ~x120 & ~x196 & ~x225 & ~x391 & ~x419 & ~x447 & ~x474 & ~x531 & ~x532 & ~x736 & ~x737 & ~x765;
assign c6372 =  x573 &  x636 &  x637 & ~x0 & ~x1 & ~x3 & ~x26 & ~x27 & ~x53 & ~x54 & ~x55 & ~x56 & ~x57 & ~x58 & ~x77 & ~x80 & ~x83 & ~x84 & ~x86 & ~x87 & ~x108 & ~x109 & ~x110 & ~x111 & ~x113 & ~x140 & ~x141 & ~x167 & ~x168 & ~x169 & ~x170 & ~x195 & ~x196 & ~x198 & ~x224 & ~x252 & ~x253 & ~x587 & ~x616 & ~x756 & ~x757 & ~x777;
assign c6374 =  x212 &  x240 &  x548 & ~x18 & ~x24 & ~x50 & ~x57 & ~x76 & ~x105 & ~x109 & ~x111 & ~x132 & ~x161 & ~x162 & ~x165 & ~x166 & ~x169 & ~x189 & ~x192 & ~x219 & ~x220 & ~x245 & ~x247 & ~x253 & ~x255 & ~x274 & ~x277 & ~x280 & ~x281 & ~x305 & ~x312 & ~x331 & ~x336 & ~x363 & ~x368 & ~x390 & ~x393 & ~x394 & ~x418 & ~x423 & ~x424 & ~x443 & ~x474 & ~x478 & ~x496 & ~x499 & ~x508 & ~x511 & ~x527 & ~x529 & ~x539 & ~x559 & ~x562 & ~x566 & ~x567 & ~x584 & ~x593 & ~x615 & ~x617 & ~x623 & ~x638 & ~x639 & ~x640 & ~x650 & ~x666 & ~x668 & ~x673 & ~x694 & ~x695 & ~x701 & ~x703 & ~x705 & ~x726 & ~x752 & ~x755 & ~x756 & ~x780 & ~x782;
assign c6376 =  x488 &  x527 & ~x24 & ~x26 & ~x357 & ~x681;
assign c6378 = ~x6 & ~x10 & ~x29 & ~x34 & ~x49 & ~x54 & ~x59 & ~x78 & ~x79 & ~x81 & ~x135 & ~x139 & ~x141 & ~x143 & ~x168 & ~x251 & ~x253 & ~x255 & ~x256 & ~x282 & ~x285 & ~x313 & ~x335 & ~x385 & ~x387 & ~x388 & ~x389 & ~x390 & ~x399 & ~x400 & ~x403 & ~x417 & ~x427 & ~x428 & ~x429 & ~x432 & ~x438 & ~x440 & ~x445 & ~x449 & ~x458 & ~x473 & ~x477 & ~x478 & ~x497 & ~x503 & ~x505 & ~x506 & ~x507 & ~x530 & ~x589 & ~x591 & ~x593 & ~x613 & ~x644 & ~x673 & ~x726 & ~x753 & ~x756 & ~x758 & ~x778;
assign c6380 =  x628 &  x656 &  x683 & ~x57 & ~x81 & ~x105 & ~x113 & ~x137 & ~x163 & ~x222 & ~x283 & ~x310 & ~x333 & ~x336 & ~x366 & ~x370 & ~x390 & ~x395 & ~x416 & ~x419 & ~x442 & ~x529 & ~x530 & ~x533 & ~x534 & ~x536 & ~x538 & ~x552 & ~x553 & ~x555 & ~x563 & ~x589 & ~x607 & ~x666 & ~x675 & ~x695 & ~x701 & ~x725 & ~x731 & ~x757 & ~x761 & ~x762;
assign c6382 = ~x2 & ~x23 & ~x24 & ~x62 & ~x93 & ~x101 & ~x192 & ~x221 & ~x222 & ~x223 & ~x224 & ~x225 & ~x227 & ~x248 & ~x250 & ~x335 & ~x347 & ~x364 & ~x375 & ~x381 & ~x391 & ~x445 & ~x448 & ~x702 & ~x748 & ~x754;
assign c6384 = ~x1 & ~x2 & ~x4 & ~x5 & ~x19 & ~x21 & ~x22 & ~x27 & ~x30 & ~x32 & ~x47 & ~x54 & ~x55 & ~x59 & ~x68 & ~x77 & ~x83 & ~x106 & ~x107 & ~x110 & ~x114 & ~x134 & ~x136 & ~x140 & ~x161 & ~x162 & ~x163 & ~x164 & ~x165 & ~x166 & ~x169 & ~x170 & ~x189 & ~x192 & ~x194 & ~x220 & ~x221 & ~x222 & ~x225 & ~x226 & ~x250 & ~x251 & ~x252 & ~x254 & ~x255 & ~x277 & ~x278 & ~x282 & ~x283 & ~x306 & ~x307 & ~x308 & ~x334 & ~x336 & ~x338 & ~x339 & ~x364 & ~x366 & ~x367 & ~x393 & ~x394 & ~x395 & ~x405 & ~x411 & ~x418 & ~x420 & ~x431 & ~x450 & ~x456 & ~x472 & ~x476 & ~x501 & ~x529 & ~x530 & ~x531 & ~x558 & ~x559 & ~x562 & ~x585 & ~x588 & ~x612 & ~x613 & ~x615 & ~x616 & ~x640 & ~x645 & ~x670 & ~x672 & ~x674 & ~x698 & ~x699 & ~x700 & ~x701 & ~x702 & ~x724 & ~x725 & ~x728 & ~x729 & ~x755 & ~x758 & ~x780 & ~x782 & ~x783;
assign c6386 =  x660 &  x688 & ~x25 & ~x27 & ~x28 & ~x51 & ~x54 & ~x81 & ~x87 & ~x111 & ~x138 & ~x142 & ~x194 & ~x221 & ~x222 & ~x248 & ~x254 & ~x255 & ~x279 & ~x280 & ~x281 & ~x310 & ~x312 & ~x337 & ~x338 & ~x339 & ~x361 & ~x364 & ~x416 & ~x454 & ~x455 & ~x456 & ~x470 & ~x489 & ~x496 & ~x504 & ~x512 & ~x513 & ~x514 & ~x527 & ~x529 & ~x530 & ~x532 & ~x537 & ~x552 & ~x553 & ~x587 & ~x588 & ~x589 & ~x590 & ~x591 & ~x613 & ~x615 & ~x616 & ~x641 & ~x647 & ~x673 & ~x725 & ~x729 & ~x757;
assign c6388 =  x572 & ~x3 & ~x30 & ~x33 & ~x83 & ~x87 & ~x88 & ~x111 & ~x116 & ~x138 & ~x139 & ~x162 & ~x166 & ~x167 & ~x189 & ~x196 & ~x209 & ~x216 & ~x217 & ~x244 & ~x245 & ~x254 & ~x278 & ~x283 & ~x309 & ~x350 & ~x529 & ~x698 & ~x715;
assign c6390 =  x451 &  x601 & ~x1 & ~x3 & ~x24 & ~x25 & ~x26 & ~x27 & ~x35 & ~x53 & ~x54 & ~x63 & ~x90 & ~x111 & ~x728 & ~x756;
assign c6392 =  x328 & ~x0 & ~x23 & ~x24 & ~x28 & ~x29 & ~x30 & ~x31 & ~x54 & ~x57 & ~x58 & ~x81 & ~x85 & ~x86 & ~x87 & ~x111 & ~x112 & ~x113 & ~x114 & ~x140 & ~x141 & ~x142 & ~x164 & ~x166 & ~x167 & ~x170 & ~x192 & ~x193 & ~x194 & ~x196 & ~x197 & ~x221 & ~x222 & ~x224 & ~x227 & ~x249 & ~x250 & ~x254 & ~x277 & ~x278 & ~x280 & ~x283 & ~x304 & ~x305 & ~x307 & ~x309 & ~x310 & ~x311 & ~x338 & ~x360 & ~x361 & ~x364 & ~x365 & ~x368 & ~x395 & ~x416 & ~x420 & ~x422 & ~x423 & ~x424 & ~x444 & ~x445 & ~x446 & ~x448 & ~x449 & ~x451 & ~x452 & ~x474 & ~x475 & ~x476 & ~x501 & ~x502 & ~x503 & ~x505 & ~x506 & ~x508 & ~x529 & ~x533 & ~x534 & ~x536 & ~x552 & ~x556 & ~x559 & ~x561 & ~x585 & ~x590 & ~x591 & ~x613 & ~x614 & ~x615 & ~x616 & ~x617 & ~x641 & ~x642 & ~x643 & ~x645 & ~x668 & ~x669 & ~x671 & ~x672 & ~x674 & ~x698 & ~x701 & ~x726 & ~x727 & ~x754 & ~x758 & ~x776 & ~x782;
assign c6394 =  x269 & ~x0 & ~x1 & ~x19 & ~x22 & ~x54 & ~x78 & ~x80 & ~x95 & ~x134 & ~x139 & ~x162 & ~x163 & ~x165 & ~x168 & ~x193 & ~x194 & ~x219 & ~x220 & ~x224 & ~x246 & ~x248 & ~x280 & ~x333 & ~x337 & ~x338 & ~x390 & ~x446 & ~x477 & ~x532 & ~x557 & ~x596 & ~x597 & ~x615 & ~x619 & ~x641 & ~x668 & ~x671 & ~x700;
assign c6396 =  x154 &  x294 &  x350 &  x550 & ~x53 & ~x85 & ~x89 & ~x391 & ~x700 & ~x783;
assign c6398 =  x434 &  x462 &  x516 &  x551 & ~x0 & ~x1 & ~x5 & ~x21 & ~x22 & ~x23 & ~x24 & ~x25 & ~x28 & ~x29 & ~x50 & ~x51 & ~x52 & ~x54 & ~x55 & ~x56 & ~x58 & ~x79 & ~x80 & ~x81 & ~x82 & ~x83 & ~x85 & ~x109 & ~x111 & ~x113 & ~x138 & ~x141 & ~x169 & ~x194 & ~x195 & ~x223 & ~x224 & ~x251 & ~x252 & ~x253 & ~x280 & ~x335 & ~x391 & ~x475 & ~x503 & ~x560 & ~x586 & ~x588 & ~x700 & ~x757 & ~x774 & ~x783;
assign c6400 =  x238 &  x601 &  x655 & ~x54 & ~x86 & ~x446 & ~x448 & ~x476 & ~x493 & ~x502 & ~x561 & ~x645 & ~x647 & ~x669 & ~x697 & ~x781;
assign c6402 =  x329 & ~x29 & ~x50 & ~x94 & ~x110 & ~x111 & ~x197 & ~x311 & ~x367 & ~x391 & ~x417 & ~x449 & ~x586 & ~x589 & ~x613;
assign c6404 =  x542 &  x579 &  x607 &  x635 & ~x2 & ~x24 & ~x25 & ~x26 & ~x27 & ~x28 & ~x30 & ~x33 & ~x51 & ~x56 & ~x81 & ~x82 & ~x83 & ~x86 & ~x110 & ~x112 & ~x138 & ~x139 & ~x141 & ~x169 & ~x196 & ~x197 & ~x224 & ~x251 & ~x252 & ~x280 & ~x281 & ~x475 & ~x503 & ~x559 & ~x586 & ~x587 & ~x614 & ~x616 & ~x670 & ~x671 & ~x672 & ~x699 & ~x728 & ~x756 & ~x763 & ~x764;
assign c6406 =  x463 &  x507 &  x535 &  x563 & ~x26 & ~x140 & ~x252 & ~x559 & ~x587;
assign c6408 =  x434 &  x495 & ~x2 & ~x29 & ~x31 & ~x55 & ~x83 & ~x138 & ~x169 & ~x197 & ~x253 & ~x447 & ~x475 & ~x531 & ~x652 & ~x680 & ~x709 & ~x719 & ~x736 & ~x746 & ~x783;
assign c6410 =  x579 & ~x27 & ~x30 & ~x81 & ~x85 & ~x107 & ~x112 & ~x169 & ~x250 & ~x308 & ~x502 & ~x559 & ~x586 & ~x595 & ~x625 & ~x653 & ~x711 & ~x780;
assign c6412 =  x449 &  x477 & ~x77 & ~x80 & ~x761;
assign c6414 =  x417 &  x528 & ~x358 & ~x385;
assign c6416 = ~x1 & ~x26 & ~x27 & ~x29 & ~x30 & ~x51 & ~x52 & ~x57 & ~x79 & ~x121 & ~x134 & ~x138 & ~x140 & ~x149 & ~x169 & ~x171 & ~x188 & ~x189 & ~x194 & ~x223 & ~x226 & ~x252 & ~x277 & ~x278 & ~x279 & ~x293 & ~x307 & ~x332 & ~x365 & ~x394 & ~x395 & ~x419 & ~x420 & ~x422 & ~x474 & ~x503 & ~x530 & ~x557 & ~x558 & ~x559 & ~x590 & ~x624 & ~x641 & ~x653 & ~x674 & ~x681 & ~x697 & ~x699 & ~x701 & ~x712 & ~x728 & ~x730 & ~x750 & ~x759 & ~x779 & ~x782;
assign c6418 =  x442 & ~x110 & ~x137 & ~x141 & ~x142 & ~x167 & ~x168 & ~x170 & ~x198 & ~x224 & ~x253 & ~x278 & ~x307 & ~x335 & ~x391 & ~x446 & ~x473 & ~x474 & ~x501 & ~x503 & ~x530 & ~x531 & ~x588 & ~x728 & ~x748 & ~x749 & ~x755 & ~x756 & ~x757 & ~x777 & ~x780;
assign c6420 =  x500 & ~x63 & ~x83 & ~x168 & ~x196 & ~x385 & ~x455;
assign c6422 =  x294 &  x518 &  x546 & ~x25 & ~x31 & ~x72 & ~x83 & ~x103 & ~x111 & ~x166 & ~x250 & ~x253 & ~x304 & ~x334 & ~x336 & ~x338 & ~x339 & ~x390 & ~x392 & ~x447 & ~x474 & ~x477 & ~x494 & ~x532 & ~x535 & ~x561 & ~x587 & ~x590 & ~x640 & ~x671 & ~x698 & ~x782;
assign c6424 = ~x9 & ~x171 & ~x227 & ~x232 & ~x280 & ~x420 & ~x429 & ~x499 & ~x535 & ~x595 & ~x598 & ~x632 & ~x652 & ~x723 & ~x736 & ~x755 & ~x773 & ~x775;
assign c6426 =  x242 &  x293 &  x602 & ~x24 & ~x51 & ~x55 & ~x142 & ~x221 & ~x222 & ~x252 & ~x253 & ~x280 & ~x335 & ~x390 & ~x391 & ~x419 & ~x559;
assign c6428 = ~x1 & ~x5 & ~x25 & ~x36 & ~x77 & ~x84 & ~x85 & ~x107 & ~x132 & ~x138 & ~x159 & ~x172 & ~x173 & ~x194 & ~x225 & ~x229 & ~x243 & ~x286 & ~x300 & ~x306 & ~x307 & ~x310 & ~x338 & ~x340 & ~x420 & ~x425 & ~x512 & ~x514 & ~x515 & ~x516 & ~x521 & ~x522 & ~x529 & ~x551 & ~x555 & ~x558 & ~x578 & ~x612 & ~x614 & ~x667 & ~x694 & ~x704 & ~x724 & ~x749 & ~x782;
assign c6430 =  x631 &  x659 &  x712 & ~x1 & ~x28 & ~x29 & ~x30 & ~x56 & ~x57 & ~x77 & ~x85 & ~x109 & ~x137 & ~x163 & ~x167 & ~x169 & ~x253 & ~x278 & ~x306 & ~x307 & ~x309 & ~x313 & ~x334 & ~x338 & ~x364 & ~x394 & ~x421 & ~x447 & ~x450 & ~x471 & ~x472 & ~x476 & ~x481 & ~x497 & ~x498 & ~x502 & ~x503 & ~x505 & ~x506 & ~x507 & ~x524 & ~x526 & ~x534 & ~x538 & ~x552 & ~x589 & ~x592 & ~x612 & ~x668 & ~x697 & ~x699 & ~x704 & ~x757 & ~x763;
assign c6432 =  x603 &  x658 &  x686 & ~x0 & ~x1 & ~x22 & ~x23 & ~x25 & ~x27 & ~x55 & ~x57 & ~x79 & ~x84 & ~x87 & ~x107 & ~x108 & ~x109 & ~x110 & ~x113 & ~x133 & ~x134 & ~x139 & ~x141 & ~x142 & ~x144 & ~x161 & ~x164 & ~x167 & ~x191 & ~x195 & ~x197 & ~x199 & ~x219 & ~x223 & ~x224 & ~x249 & ~x250 & ~x254 & ~x257 & ~x278 & ~x279 & ~x281 & ~x282 & ~x309 & ~x312 & ~x332 & ~x338 & ~x340 & ~x360 & ~x365 & ~x367 & ~x368 & ~x388 & ~x389 & ~x390 & ~x391 & ~x393 & ~x420 & ~x423 & ~x450 & ~x454 & ~x470 & ~x471 & ~x477 & ~x481 & ~x500 & ~x501 & ~x505 & ~x507 & ~x508 & ~x509 & ~x524 & ~x528 & ~x531 & ~x536 & ~x537 & ~x553 & ~x554 & ~x556 & ~x558 & ~x559 & ~x560 & ~x561 & ~x579 & ~x583 & ~x587 & ~x588 & ~x595 & ~x608 & ~x610 & ~x613 & ~x618 & ~x640 & ~x643 & ~x649 & ~x670 & ~x675 & ~x697 & ~x698 & ~x705 & ~x724 & ~x725 & ~x730 & ~x731 & ~x733 & ~x753 & ~x756 & ~x757 & ~x758 & ~x759 & ~x760 & ~x781;
assign c6434 = ~x55 & ~x80 & ~x106 & ~x114 & ~x169 & ~x192 & ~x224 & ~x228 & ~x230 & ~x246 & ~x251 & ~x255 & ~x257 & ~x258 & ~x275 & ~x284 & ~x285 & ~x307 & ~x311 & ~x333 & ~x337 & ~x341 & ~x358 & ~x359 & ~x364 & ~x389 & ~x390 & ~x391 & ~x394 & ~x398 & ~x418 & ~x419 & ~x420 & ~x424 & ~x425 & ~x426 & ~x427 & ~x434 & ~x447 & ~x452 & ~x455 & ~x458 & ~x469 & ~x485 & ~x486 & ~x494 & ~x496 & ~x498 & ~x504 & ~x510 & ~x511 & ~x528 & ~x554 & ~x561 & ~x615 & ~x616 & ~x639 & ~x640 & ~x646 & ~x648 & ~x671 & ~x723 & ~x728 & ~x779;
assign c6436 =  x368 &  x540 & ~x63 & ~x64 & ~x82 & ~x91 & ~x118 & ~x145 & ~x146 & ~x167 & ~x756 & ~x776 & ~x783;
assign c6438 = ~x23 & ~x24 & ~x27 & ~x84 & ~x86 & ~x109 & ~x135 & ~x136 & ~x140 & ~x168 & ~x193 & ~x197 & ~x199 & ~x225 & ~x248 & ~x255 & ~x305 & ~x306 & ~x311 & ~x314 & ~x333 & ~x335 & ~x340 & ~x416 & ~x421 & ~x429 & ~x430 & ~x437 & ~x445 & ~x448 & ~x468 & ~x480 & ~x493 & ~x496 & ~x508 & ~x510 & ~x528 & ~x529 & ~x533 & ~x561 & ~x584 & ~x613 & ~x645 & ~x727 & ~x731 & ~x732 & ~x759;
assign c6440 =  x518 &  x579 & ~x3 & ~x4 & ~x5 & ~x7 & ~x27 & ~x35 & ~x51 & ~x81 & ~x111 & ~x137 & ~x139 & ~x165 & ~x194 & ~x252 & ~x278 & ~x279 & ~x280 & ~x307 & ~x335 & ~x383 & ~x737 & ~x756 & ~x764;
assign c6442 =  x213 &  x292 &  x632 & ~x23 & ~x25 & ~x54 & ~x108 & ~x109 & ~x113 & ~x136 & ~x140 & ~x166 & ~x198 & ~x219 & ~x225 & ~x247 & ~x249 & ~x253 & ~x283 & ~x305 & ~x312 & ~x334 & ~x339 & ~x367 & ~x391 & ~x470 & ~x475 & ~x476 & ~x498 & ~x503 & ~x526 & ~x538 & ~x588 & ~x643 & ~x644 & ~x646 & ~x647 & ~x728 & ~x754 & ~x756 & ~x781;
assign c6444 =  x443 &  x592 & ~x419 & ~x474 & ~x475;
assign c6446 =  x434 & ~x0 & ~x1 & ~x25 & ~x26 & ~x81 & ~x82 & ~x109 & ~x162 & ~x163 & ~x166 & ~x168 & ~x220 & ~x224 & ~x225 & ~x226 & ~x390 & ~x419 & ~x545 & ~x554 & ~x558 & ~x572 & ~x596 & ~x597 & ~x598 & ~x614 & ~x624 & ~x641 & ~x680 & ~x753 & ~x776;
assign c6448 =  x304 &  x436 & ~x251 & ~x279 & ~x307 & ~x335;
assign c6450 = ~x1 & ~x5 & ~x30 & ~x33 & ~x36 & ~x53 & ~x62 & ~x79 & ~x86 & ~x87 & ~x91 & ~x103 & ~x111 & ~x114 & ~x115 & ~x117 & ~x131 & ~x133 & ~x136 & ~x160 & ~x165 & ~x171 & ~x192 & ~x196 & ~x222 & ~x228 & ~x251 & ~x255 & ~x257 & ~x275 & ~x287 & ~x308 & ~x311 & ~x315 & ~x317 & ~x362 & ~x363 & ~x368 & ~x391 & ~x392 & ~x394 & ~x414 & ~x418 & ~x419 & ~x453 & ~x470 & ~x494 & ~x495 & ~x503 & ~x506 & ~x526 & ~x541 & ~x549 & ~x553 & ~x564 & ~x577 & ~x584 & ~x588 & ~x589 & ~x592 & ~x594 & ~x595 & ~x606 & ~x615 & ~x623 & ~x646 & ~x664 & ~x700 & ~x721 & ~x729 & ~x753 & ~x754 & ~x755 & ~x756 & ~x780;
assign c6452 =  x600 &  x626 & ~x5 & ~x27 & ~x31 & ~x56 & ~x138 & ~x194 & ~x195 & ~x251 & ~x280 & ~x281 & ~x311 & ~x442 & ~x446 & ~x466 & ~x467 & ~x468 & ~x472 & ~x476 & ~x523 & ~x699 & ~x760;
assign c6454 =  x269 &  x297 &  x606 & ~x1 & ~x2 & ~x30 & ~x53 & ~x55 & ~x56 & ~x81 & ~x82 & ~x107 & ~x108 & ~x113 & ~x136 & ~x140 & ~x166 & ~x168 & ~x169 & ~x196 & ~x224 & ~x249 & ~x278 & ~x282 & ~x283 & ~x305 & ~x306 & ~x311 & ~x312 & ~x335 & ~x337 & ~x363 & ~x392 & ~x393 & ~x420 & ~x421 & ~x449 & ~x474 & ~x475 & ~x498 & ~x501 & ~x503 & ~x504 & ~x505 & ~x508 & ~x509 & ~x525 & ~x560 & ~x588 & ~x591 & ~x612 & ~x613 & ~x618 & ~x643 & ~x644 & ~x670 & ~x671 & ~x673 & ~x675 & ~x699 & ~x702 & ~x704 & ~x726 & ~x727 & ~x730 & ~x754 & ~x755 & ~x760 & ~x783;
assign c6456 = ~x3 & ~x4 & ~x19 & ~x24 & ~x51 & ~x58 & ~x116 & ~x143 & ~x162 & ~x191 & ~x203 & ~x247 & ~x251 & ~x257 & ~x274 & ~x277 & ~x279 & ~x333 & ~x336 & ~x337 & ~x338 & ~x392 & ~x395 & ~x396 & ~x444 & ~x445 & ~x451 & ~x474 & ~x503 & ~x505 & ~x512 & ~x537 & ~x558 & ~x612 & ~x616 & ~x623 & ~x650 & ~x659 & ~x687 & ~x700 & ~x718 & ~x728 & ~x743 & ~x752 & ~x757 & ~x761 & ~x770 & ~x772 & ~x776 & ~x781;
assign c6458 =  x328 & ~x1 & ~x2 & ~x4 & ~x26 & ~x31 & ~x53 & ~x55 & ~x56 & ~x57 & ~x65 & ~x82 & ~x86 & ~x108 & ~x114 & ~x116 & ~x137 & ~x141 & ~x143 & ~x168 & ~x170 & ~x193 & ~x221 & ~x222 & ~x223 & ~x249 & ~x277 & ~x279 & ~x281 & ~x304 & ~x305 & ~x307 & ~x334 & ~x360 & ~x361 & ~x363 & ~x366 & ~x391 & ~x416 & ~x443 & ~x444 & ~x446 & ~x447 & ~x478 & ~x480 & ~x501 & ~x504 & ~x505 & ~x527 & ~x528 & ~x534 & ~x535 & ~x555 & ~x561 & ~x562 & ~x615 & ~x645 & ~x648 & ~x673 & ~x674 & ~x699 & ~x703 & ~x704 & ~x753 & ~x754;
assign c6460 =  x442 &  x551 & ~x170 & ~x196 & ~x253 & ~x299 & ~x391 & ~x729;
assign c6462 =  x604 & ~x2 & ~x49 & ~x78 & ~x87 & ~x105 & ~x106 & ~x107 & ~x165 & ~x171 & ~x193 & ~x195 & ~x196 & ~x223 & ~x308 & ~x474 & ~x475 & ~x476 & ~x504 & ~x505 & ~x533 & ~x557 & ~x782;
assign c6464 =  x394 &  x488 &  x555;
assign c6466 =  x434 &  x450 & ~x49 & ~x50 & ~x52 & ~x55 & ~x80 & ~x83 & ~x112 & ~x762;
assign c6468 =  x551 &  x664 & ~x1 & ~x4 & ~x7 & ~x23 & ~x24 & ~x28 & ~x35 & ~x52 & ~x61 & ~x81 & ~x82 & ~x83 & ~x116 & ~x117 & ~x169 & ~x196 & ~x254 & ~x281 & ~x706 & ~x707 & ~x756 & ~x764 & ~x766;
assign c6470 =  x182 &  x237 &  x322 &  x406 & ~x44 & ~x45 & ~x397 & ~x589 & ~x593;
assign c6472 =  x238 &  x657 &  x684 & ~x31 & ~x57 & ~x139 & ~x224 & ~x338 & ~x367 & ~x422 & ~x445 & ~x472 & ~x514 & ~x524 & ~x561 & ~x563 & ~x568 & ~x587 & ~x619 & ~x670 & ~x781;
assign c6474 = ~x3 & ~x25 & ~x26 & ~x27 & ~x32 & ~x83 & ~x109 & ~x113 & ~x114 & ~x136 & ~x138 & ~x141 & ~x193 & ~x195 & ~x196 & ~x198 & ~x221 & ~x225 & ~x252 & ~x256 & ~x258 & ~x277 & ~x278 & ~x303 & ~x306 & ~x309 & ~x312 & ~x334 & ~x337 & ~x339 & ~x341 & ~x357 & ~x358 & ~x362 & ~x370 & ~x388 & ~x390 & ~x393 & ~x394 & ~x399 & ~x409 & ~x416 & ~x418 & ~x420 & ~x427 & ~x431 & ~x432 & ~x437 & ~x443 & ~x445 & ~x450 & ~x454 & ~x482 & ~x483 & ~x484 & ~x497 & ~x500 & ~x504 & ~x506 & ~x527 & ~x534 & ~x535 & ~x559 & ~x560 & ~x583 & ~x586 & ~x591 & ~x594 & ~x610 & ~x615 & ~x643 & ~x646 & ~x699 & ~x726 & ~x730 & ~x731 & ~x732 & ~x751 & ~x753 & ~x755 & ~x756 & ~x759 & ~x778 & ~x780;
assign c6476 =  x461 &  x542 &  x578 & ~x0 & ~x7 & ~x23 & ~x24 & ~x27 & ~x52 & ~x82 & ~x90 & ~x118 & ~x138 & ~x195 & ~x252 & ~x749 & ~x756;
assign c6478 =  x352 & ~x0 & ~x55 & ~x78 & ~x88 & ~x103 & ~x105 & ~x110 & ~x116 & ~x159 & ~x162 & ~x187 & ~x197 & ~x220 & ~x222 & ~x224 & ~x226 & ~x244 & ~x247 & ~x254 & ~x279 & ~x313 & ~x332 & ~x336 & ~x389 & ~x391 & ~x396 & ~x443 & ~x475 & ~x482 & ~x503 & ~x512 & ~x513 & ~x523 & ~x524 & ~x542 & ~x560 & ~x563 & ~x567 & ~x579 & ~x591 & ~x597 & ~x608 & ~x610 & ~x619 & ~x621 & ~x624 & ~x644 & ~x668 & ~x674 & ~x677 & ~x729 & ~x735 & ~x750 & ~x781;
assign c6480 =  x572 &  x574 &  x604 &  x633 & ~x27 & ~x249 & ~x279 & ~x334 & ~x523 & ~x641 & ~x643 & ~x669;
assign c6482 =  x44 & ~x0 & ~x22 & ~x24 & ~x27 & ~x29 & ~x38 & ~x39 & ~x40 & ~x66 & ~x68 & ~x79 & ~x82 & ~x84 & ~x106 & ~x108 & ~x109 & ~x110 & ~x112 & ~x113 & ~x114 & ~x132 & ~x133 & ~x134 & ~x136 & ~x137 & ~x138 & ~x139 & ~x141 & ~x142 & ~x143 & ~x161 & ~x166 & ~x190 & ~x191 & ~x193 & ~x195 & ~x196 & ~x197 & ~x198 & ~x199 & ~x221 & ~x222 & ~x223 & ~x224 & ~x248 & ~x249 & ~x250 & ~x251 & ~x255 & ~x277 & ~x278 & ~x281 & ~x282 & ~x305 & ~x306 & ~x307 & ~x308 & ~x309 & ~x333 & ~x334 & ~x335 & ~x336 & ~x337 & ~x363 & ~x365 & ~x390 & ~x391 & ~x417 & ~x418 & ~x419 & ~x447 & ~x475 & ~x477 & ~x501 & ~x502 & ~x504 & ~x505 & ~x527 & ~x530 & ~x531 & ~x532 & ~x533 & ~x559 & ~x586 & ~x587 & ~x589 & ~x590 & ~x614 & ~x616 & ~x617 & ~x642 & ~x643 & ~x644 & ~x645 & ~x646 & ~x672 & ~x675 & ~x676 & ~x698 & ~x699 & ~x700 & ~x701 & ~x702 & ~x703 & ~x704 & ~x727 & ~x729 & ~x746 & ~x753 & ~x756 & ~x757 & ~x781;
assign c6484 =  x156 &  x379 &  x606 & ~x25 & ~x26 & ~x28 & ~x54 & ~x55 & ~x111 & ~x112 & ~x139 & ~x141 & ~x252 & ~x559 & ~x643 & ~x670 & ~x672 & ~x698 & ~x700 & ~x726;
assign c6486 = ~x114 & ~x163 & ~x192 & ~x256 & ~x313 & ~x336 & ~x395 & ~x407 & ~x426 & ~x447 & ~x463 & ~x471 & ~x481 & ~x528 & ~x539 & ~x557 & ~x582 & ~x588 & ~x730 & ~x771 & ~x773;
assign c6488 =  x233 &  x604 & ~x4 & ~x8 & ~x23 & ~x27 & ~x28 & ~x37 & ~x52 & ~x53 & ~x57 & ~x78 & ~x81 & ~x82 & ~x84 & ~x86 & ~x111 & ~x112 & ~x167 & ~x171 & ~x224 & ~x226 & ~x281 & ~x338 & ~x391 & ~x420 & ~x444 & ~x446 & ~x448 & ~x473 & ~x475 & ~x477 & ~x531 & ~x533 & ~x554 & ~x616 & ~x640 & ~x701 & ~x727 & ~x782 & ~x783;
assign c6490 =  x243 & ~x1 & ~x2 & ~x5 & ~x25 & ~x66 & ~x112 & ~x136 & ~x140 & ~x142 & ~x167 & ~x168 & ~x199 & ~x224 & ~x225 & ~x228 & ~x248 & ~x278 & ~x280 & ~x284 & ~x285 & ~x337 & ~x339 & ~x340 & ~x368 & ~x394 & ~x448 & ~x449 & ~x452 & ~x476 & ~x505 & ~x553 & ~x561 & ~x589 & ~x611 & ~x613 & ~x615 & ~x620 & ~x639 & ~x701 & ~x751 & ~x756 & ~x782;
assign c6492 =  x212 &  x463 &  x491 &  x636 & ~x0 & ~x1 & ~x25 & ~x26 & ~x29 & ~x51 & ~x52 & ~x80 & ~x84 & ~x138 & ~x166 & ~x167 & ~x168 & ~x194 & ~x224 & ~x252 & ~x699 & ~x782 & ~x783;
assign c6494 =  x181 & ~x45 & ~x72 & ~x87 & ~x88 & ~x116 & ~x117 & ~x145 & ~x319 & ~x334 & ~x340 & ~x453 & ~x471 & ~x501 & ~x551 & ~x584 & ~x698 & ~x732 & ~x754;
assign c6496 = ~x4 & ~x22 & ~x23 & ~x53 & ~x54 & ~x55 & ~x56 & ~x78 & ~x85 & ~x87 & ~x107 & ~x112 & ~x115 & ~x141 & ~x165 & ~x168 & ~x169 & ~x193 & ~x198 & ~x223 & ~x226 & ~x227 & ~x228 & ~x251 & ~x254 & ~x255 & ~x306 & ~x312 & ~x333 & ~x335 & ~x336 & ~x363 & ~x368 & ~x386 & ~x412 & ~x417 & ~x422 & ~x430 & ~x436 & ~x445 & ~x456 & ~x479 & ~x480 & ~x495 & ~x497 & ~x502 & ~x503 & ~x510 & ~x533 & ~x534 & ~x553 & ~x559 & ~x561 & ~x564 & ~x567 & ~x584 & ~x594 & ~x617 & ~x618 & ~x619 & ~x620 & ~x622 & ~x640 & ~x670 & ~x674 & ~x701 & ~x720 & ~x725 & ~x728 & ~x730 & ~x749 & ~x753 & ~x777;
assign c6498 =  x158 &  x578 & ~x25 & ~x30 & ~x55 & ~x56 & ~x78 & ~x81 & ~x86 & ~x90 & ~x91 & ~x108 & ~x109 & ~x112 & ~x138 & ~x139 & ~x140 & ~x142 & ~x166 & ~x168 & ~x170 & ~x197 & ~x223 & ~x335 & ~x419 & ~x559 & ~x728 & ~x734 & ~x735 & ~x756 & ~x757 & ~x761 & ~x783;
assign c61 =  x195;
assign c63 =  x467 & ~x158 & ~x202 & ~x460;
assign c65 =  x292 & ~x105 & ~x134 & ~x214 & ~x245 & ~x268 & ~x269 & ~x450 & ~x678 & ~x737 & ~x764 & ~x780;
assign c67 =  x485 & ~x393 & ~x461 & ~x479;
assign c69 =  x41 &  x98 &  x743 & ~x7 & ~x22 & ~x34 & ~x86 & ~x103 & ~x104 & ~x108 & ~x137 & ~x145 & ~x160 & ~x162 & ~x172 & ~x189 & ~x192 & ~x202 & ~x252 & ~x281 & ~x303 & ~x366 & ~x423 & ~x477 & ~x478 & ~x480 & ~x506 & ~x530 & ~x532 & ~x533 & ~x587 & ~x642 & ~x725 & ~x754 & ~x759;
assign c611 =  x211 & ~x197 & ~x218 & ~x247 & ~x302 & ~x305 & ~x308 & ~x332 & ~x334 & ~x359 & ~x361 & ~x389 & ~x604 & ~x605 & ~x606 & ~x627 & ~x632;
assign c613 =  x783;
assign c615 =  x756;
assign c617 =  x354 &  x381 & ~x25 & ~x275 & ~x306 & ~x333 & ~x334 & ~x335 & ~x359 & ~x601 & ~x602;
assign c619 =  x117;
assign c621 =  x318 &  x373 &  x374 & ~x78 & ~x597 & ~x655;
assign c623 =  x360 & ~x567 & ~x569 & ~x592 & ~x625 & ~x674;
assign c625 =  x463 & ~x1 & ~x22 & ~x26 & ~x27 & ~x30 & ~x50 & ~x52 & ~x77 & ~x81 & ~x140 & ~x166 & ~x168 & ~x197 & ~x295 & ~x429 & ~x447 & ~x457 & ~x481 & ~x504 & ~x510 & ~x511 & ~x512 & ~x532 & ~x535 & ~x540 & ~x561 & ~x587 & ~x589 & ~x590 & ~x614 & ~x641 & ~x647 & ~x668 & ~x672 & ~x675 & ~x696 & ~x723 & ~x725 & ~x727 & ~x728 & ~x731 & ~x748 & ~x751 & ~x754 & ~x758 & ~x779;
assign c627 =  x742 & ~x26 & ~x277 & ~x363 & ~x389 & ~x423 & ~x533 & ~x637 & ~x639 & ~x642 & ~x659 & ~x660 & ~x662 & ~x666 & ~x671;
assign c629 =  x326 & ~x333 & ~x573 & ~x602;
assign c631 =  x252;
assign c633 =  x119 & ~x99 & ~x156 & ~x237;
assign c635 = ~x0 & ~x12 & ~x15 & ~x16 & ~x77 & ~x80 & ~x81 & ~x131 & ~x141 & ~x163 & ~x165 & ~x184 & ~x185 & ~x189 & ~x336 & ~x448 & ~x565 & ~x585 & ~x620 & ~x645 & ~x673 & ~x700 & ~x729 & ~x730 & ~x732 & ~x733;
assign c637 =  x742 &  x743 & ~x22 & ~x608 & ~x633 & ~x660;
assign c639 =  x126 & ~x3 & ~x10 & ~x25 & ~x31 & ~x52 & ~x53 & ~x83 & ~x114 & ~x170 & ~x214 & ~x245 & ~x247 & ~x252 & ~x271 & ~x280 & ~x302 & ~x330 & ~x358 & ~x359 & ~x386 & ~x388 & ~x393 & ~x422 & ~x449 & ~x457 & ~x585 & ~x627 & ~x641 & ~x642 & ~x644 & ~x656 & ~x703 & ~x723 & ~x725 & ~x727 & ~x728 & ~x758;
assign c641 =  x625 & ~x88 & ~x276 & ~x503 & ~x600;
assign c643 =  x111;
assign c645 =  x234 & ~x55 & ~x103 & ~x614 & ~x621 & ~x643 & ~x649 & ~x668 & ~x701 & ~x703 & ~x722 & ~x723 & ~x742 & ~x749 & ~x773 & ~x774;
assign c647 = ~x70 & ~x113 & ~x164 & ~x674 & ~x686 & ~x690 & ~x703 & ~x709 & ~x747 & ~x760;
assign c649 =  x97 &  x659 & ~x118 & ~x159 & ~x170 & ~x172 & ~x176 & ~x189 & ~x221 & ~x428 & ~x481 & ~x613;
assign c651 =  x316 &  x343 & ~x6 & ~x7 & ~x540 & ~x566 & ~x567 & ~x594 & ~x648 & ~x651 & ~x677 & ~x679 & ~x702 & ~x726 & ~x730;
assign c653 =  x372 &  x418 & ~x690;
assign c655 = ~x29 & ~x48 & ~x80 & ~x86 & ~x88 & ~x89 & ~x110 & ~x138 & ~x142 & ~x224 & ~x225 & ~x447 & ~x468 & ~x469 & ~x496 & ~x525 & ~x543 & ~x564 & ~x570 & ~x572 & ~x588 & ~x589 & ~x592 & ~x598 & ~x619 & ~x627 & ~x628 & ~x645 & ~x657 & ~x671 & ~x672 & ~x697 & ~x712 & ~x729 & ~x730 & ~x757 & ~x778 & ~x779;
assign c657 =  x296 & ~x24 & ~x26 & ~x169 & ~x225 & ~x633 & ~x659 & ~x661 & ~x663 & ~x664 & ~x721 & ~x774;
assign c659 =  x404 &  x745 & ~x176 & ~x298 & ~x333 & ~x386;
assign c661 =  x274 &  x427;
assign c663 =  x415 &  x474;
assign c665 =  x93 &  x151 & ~x321;
assign c667 =  x154 &  x182 & ~x23 & ~x50 & ~x65 & ~x77 & ~x87 & ~x113 & ~x141 & ~x146 & ~x164 & ~x192 & ~x215 & ~x221 & ~x223 & ~x229 & ~x242 & ~x244 & ~x259 & ~x269 & ~x284 & ~x297 & ~x299 & ~x309 & ~x311 & ~x312 & ~x328 & ~x355 & ~x368 & ~x385 & ~x391 & ~x394 & ~x532 & ~x533 & ~x557 & ~x586 & ~x590 & ~x614 & ~x732 & ~x755;
assign c669 =  x69 & ~x31 & ~x55 & ~x56 & ~x58 & ~x81 & ~x139 & ~x168 & ~x252 & ~x432 & ~x433 & ~x435;
assign c671 =  x154 &  x345 &  x400 & ~x654;
assign c673 =  x360 & ~x551;
assign c675 = ~x180 & ~x181 & ~x353 & ~x409 & ~x655 & ~x739;
assign c677 =  x632 & ~x56 & ~x216 & ~x227 & ~x240 & ~x270 & ~x329 & ~x333 & ~x384;
assign c679 =  x124 &  x318 & ~x22 & ~x25 & ~x31 & ~x47 & ~x48 & ~x55 & ~x60 & ~x81 & ~x86 & ~x106 & ~x108 & ~x136 & ~x166 & ~x191 & ~x197 & ~x214 & ~x216 & ~x246 & ~x249 & ~x255 & ~x256 & ~x280 & ~x283 & ~x307 & ~x560 & ~x672 & ~x703 & ~x752 & ~x779;
assign c681 =  x566 & ~x550;
assign c683 =  x603 & ~x19 & ~x22 & ~x24 & ~x28 & ~x47 & ~x55 & ~x58 & ~x65 & ~x66 & ~x81 & ~x109 & ~x145 & ~x170 & ~x224 & ~x279 & ~x308 & ~x356 & ~x510 & ~x537 & ~x559 & ~x566 & ~x569 & ~x570 & ~x580 & ~x581 & ~x585 & ~x587 & ~x594 & ~x615 & ~x617 & ~x620 & ~x626 & ~x637 & ~x645 & ~x648 & ~x651 & ~x652 & ~x654 & ~x666 & ~x668 & ~x673 & ~x683 & ~x697 & ~x698 & ~x699 & ~x703 & ~x721 & ~x730 & ~x733 & ~x734 & ~x736 & ~x756 & ~x764;
assign c685 =  x66 &  x95 &  x123 & ~x0 & ~x17 & ~x18 & ~x22 & ~x23 & ~x25 & ~x50 & ~x75 & ~x102 & ~x105 & ~x137 & ~x143 & ~x252 & ~x253 & ~x615 & ~x730;
assign c687 = ~x414 & ~x442 & ~x488 & ~x571 & ~x573 & ~x654 & ~x656 & ~x713;
assign c689 =  x276 & ~x379 & ~x406;
assign c691 = ~x29 & ~x34 & ~x47 & ~x57 & ~x76 & ~x78 & ~x115 & ~x140 & ~x162 & ~x170 & ~x188 & ~x189 & ~x198 & ~x201 & ~x214 & ~x240 & ~x269 & ~x295 & ~x391 & ~x392 & ~x422 & ~x448 & ~x699 & ~x703 & ~x733 & ~x761 & ~x781;
assign c695 = ~x44 & ~x128 & ~x156 & ~x265 & ~x721 & ~x768;
assign c697 = ~x17 & ~x46 & ~x56 & ~x74 & ~x157 & ~x211 & ~x393 & ~x643 & ~x680 & ~x740 & ~x761;
assign c699 =  x110;
assign c6101 =  x441 & ~x323;
assign c6103 = ~x55 & ~x99 & ~x121 & ~x572 & ~x628 & ~x686;
assign c6105 =  x347 & ~x13 & ~x16 & ~x43 & ~x653;
assign c6107 =  x66 &  x150 &  x179 & ~x101;
assign c6109 =  x210 & ~x324 & ~x378 & ~x446 & ~x698;
assign c6111 =  x112 & ~x488;
assign c6113 = ~x17 & ~x47 & ~x102 & ~x158 & ~x211 & ~x420 & ~x455 & ~x647 & ~x671 & ~x697;
assign c6115 =  x94 & ~x102 & ~x129 & ~x184 & ~x448 & ~x724 & ~x760;
assign c6117 =  x137;
assign c6119 =  x64 &  x121 & ~x100;
assign c6121 =  x64;
assign c6123 =  x469 & ~x102 & ~x407;
assign c6125 =  x374 &  x431 & ~x408 & ~x523;
assign c6127 =  x94 &  x151 & ~x108 & ~x129;
assign c6129 =  x111;
assign c6131 =  x14 & ~x602 & ~x603 & ~x632;
assign c6133 =  x1;
assign c6135 =  x120 &  x121 &  x232 & ~x71 & ~x346;
assign c6137 =  x351 & ~x334 & ~x360 & ~x392 & ~x416 & ~x478 & ~x530 & ~x627 & ~x632 & ~x633 & ~x634 & ~x656;
assign c6139 = ~x4 & ~x26 & ~x40 & ~x59 & ~x84 & ~x94 & ~x253 & ~x386 & ~x414 & ~x415 & ~x459 & ~x486 & ~x487 & ~x515 & ~x570 & ~x571 & ~x598 & ~x616 & ~x629 & ~x671 & ~x730 & ~x755 & ~x759;
assign c6141 =  x98 & ~x7 & ~x21 & ~x77 & ~x87 & ~x103 & ~x131 & ~x159 & ~x198 & ~x199 & ~x276 & ~x280 & ~x307 & ~x332 & ~x404 & ~x430 & ~x455 & ~x458 & ~x617;
assign c6143 =  x783;
assign c6145 =  x383 & ~x517 & ~x631;
assign c6147 =  x347 & ~x469 & ~x521 & ~x522 & ~x550 & ~x597 & ~x680;
assign c6149 =  x357 &  x359;
assign c6151 =  x232 & ~x13 & ~x14 & ~x31 & ~x41 & ~x42 & ~x139 & ~x587 & ~x588 & ~x621 & ~x642 & ~x643 & ~x649 & ~x668 & ~x696 & ~x697 & ~x703 & ~x704 & ~x725 & ~x757 & ~x759 & ~x766 & ~x776;
assign c6153 =  x430 &  x573 & ~x9 & ~x440 & ~x682;
assign c6155 = ~x45 & ~x74 & ~x101 & ~x159 & ~x240 & ~x267 & ~x484 & ~x561 & ~x672 & ~x723;
assign c6157 =  x118 & ~x354 & ~x493 & ~x494;
assign c6159 =  x90 &  x559;
assign c6161 = ~x35 & ~x408 & ~x435 & ~x437 & ~x464 & ~x542 & ~x654 & ~x709;
assign c6163 =  x116 &  x134;
assign c6165 =  x140;
assign c6167 =  x296 & ~x81 & ~x85 & ~x169 & ~x573 & ~x575 & ~x604;
assign c6169 =  x621 & ~x549 & ~x634;
assign c6171 =  x702 & ~x634;
assign c6173 =  x427 & ~x580 & ~x583;
assign c6175 =  x456 & ~x432 & ~x461 & ~x469;
assign c6177 = ~x72 & ~x95 & ~x96 & ~x693 & ~x714 & ~x719 & ~x731 & ~x744;
assign c6179 =  x494 & ~x32 & ~x47 & ~x53 & ~x57 & ~x85 & ~x102 & ~x105 & ~x111 & ~x112 & ~x134 & ~x145 & ~x172 & ~x175 & ~x192 & ~x196 & ~x215 & ~x219 & ~x251 & ~x253 & ~x276 & ~x281 & ~x332 & ~x337 & ~x361 & ~x392 & ~x482 & ~x616 & ~x643 & ~x754 & ~x778 & ~x783;
assign c6181 =  x743 &  x771 & ~x31 & ~x104 & ~x105 & ~x110 & ~x131 & ~x146 & ~x160 & ~x172 & ~x202 & ~x206 & ~x256 & ~x283 & ~x287 & ~x307 & ~x342 & ~x392 & ~x427 & ~x452 & ~x734 & ~x763;
assign c6183 =  x37 &  x94 &  x95;
assign c6185 =  x715 & ~x24 & ~x114 & ~x140 & ~x255 & ~x451 & ~x528 & ~x550 & ~x551 & ~x576 & ~x643 & ~x704 & ~x709 & ~x725 & ~x738;
assign c6187 =  x265 & ~x134 & ~x406 & ~x435;
assign c6189 =  x162 & ~x263;
assign c6191 =  x741 & ~x58 & ~x300 & ~x304 & ~x472 & ~x657 & ~x666;
assign c6193 =  x262 & ~x521 & ~x599;
assign c6195 =  x266 & ~x130 & ~x406 & ~x433 & ~x718 & ~x720;
assign c6197 =  x594 & ~x388 & ~x632 & ~x633;
assign c6199 =  x352 & ~x25 & ~x29 & ~x305 & ~x516 & ~x629 & ~x658;
assign c6201 =  x98 &  x153 & ~x294 & ~x295 & ~x533 & ~x614;
assign c6203 =  x600 & ~x24 & ~x62 & ~x252 & ~x534 & ~x535 & ~x624 & ~x625 & ~x633 & ~x634 & ~x636 & ~x643 & ~x654 & ~x710 & ~x726 & ~x739 & ~x758;
assign c6205 =  x487 &  x514 & ~x31 & ~x392 & ~x448 & ~x576 & ~x578 & ~x579 & ~x580 & ~x582 & ~x643 & ~x755;
assign c6207 =  x379 & ~x73 & ~x101 & ~x102 & ~x157 & ~x185 & ~x239 & ~x455;
assign c6209 =  x437 & ~x157 & ~x216 & ~x406;
assign c6211 = ~x99 & ~x154 & ~x184 & ~x242 & ~x694 & ~x721 & ~x768;
assign c6213 =  x542 & ~x46 & ~x132 & ~x134 & ~x256 & ~x549 & ~x551 & ~x552 & ~x554 & ~x576 & ~x578 & ~x643 & ~x756;
assign c6215 =  x140;
assign c6217 =  x154 &  x347 & ~x466;
assign c6219 =  x491 & ~x56 & ~x459 & ~x542 & ~x571 & ~x572 & ~x580 & ~x627;
assign c6221 =  x344 &  x391;
assign c6223 =  x303 &  x306;
assign c6225 =  x356 & ~x463 & ~x684;
assign c6227 = ~x0 & ~x1 & ~x2 & ~x5 & ~x7 & ~x22 & ~x25 & ~x32 & ~x34 & ~x35 & ~x38 & ~x49 & ~x50 & ~x51 & ~x58 & ~x60 & ~x77 & ~x78 & ~x79 & ~x83 & ~x87 & ~x111 & ~x136 & ~x141 & ~x142 & ~x166 & ~x168 & ~x170 & ~x192 & ~x199 & ~x202 & ~x215 & ~x218 & ~x221 & ~x234 & ~x241 & ~x242 & ~x243 & ~x244 & ~x247 & ~x249 & ~x250 & ~x251 & ~x255 & ~x258 & ~x269 & ~x272 & ~x273 & ~x275 & ~x284 & ~x297 & ~x301 & ~x302 & ~x303 & ~x305 & ~x307 & ~x309 & ~x332 & ~x337 & ~x365 & ~x391 & ~x392 & ~x394 & ~x395 & ~x396 & ~x398 & ~x414 & ~x415 & ~x417 & ~x419 & ~x422 & ~x425 & ~x426 & ~x446 & ~x448 & ~x449 & ~x451 & ~x472 & ~x474 & ~x475 & ~x499 & ~x500 & ~x502 & ~x507 & ~x533 & ~x559 & ~x564 & ~x590 & ~x611 & ~x613 & ~x614 & ~x616 & ~x619 & ~x638 & ~x641 & ~x646 & ~x648 & ~x666 & ~x669 & ~x671 & ~x677 & ~x694 & ~x705 & ~x722 & ~x723 & ~x726 & ~x728 & ~x729 & ~x752 & ~x761 & ~x762 & ~x763 & ~x780 & ~x783;
assign c6229 =  x196;
assign c6231 = ~x405 & ~x462 & ~x464 & ~x548;
assign c6233 =  x154 &  x320 & ~x6 & ~x7 & ~x22 & ~x23 & ~x32 & ~x33 & ~x52 & ~x63 & ~x88 & ~x90 & ~x105 & ~x110 & ~x135 & ~x137 & ~x148 & ~x164 & ~x168 & ~x196 & ~x200 & ~x227 & ~x228 & ~x308 & ~x584 & ~x585 & ~x726 & ~x729 & ~x735 & ~x738 & ~x739 & ~x763 & ~x766;
assign c6235 =  x140;
assign c6237 =  x94 &  x206 & ~x321;
assign c6239 =  x263 &  x290 &  x291 & ~x76 & ~x102 & ~x376 & ~x377;
assign c6241 =  x743 & ~x476 & ~x499 & ~x508 & ~x557 & ~x606 & ~x607 & ~x631 & ~x632;
assign c6243 =  x41 &  x71 &  x125 & ~x159 & ~x203 & ~x444 & ~x640 & ~x643 & ~x677 & ~x760;
assign c6245 = ~x27 & ~x146 & ~x197 & ~x220 & ~x268 & ~x271 & ~x284 & ~x286 & ~x301 & ~x304 & ~x327 & ~x330 & ~x384 & ~x393 & ~x448 & ~x526 & ~x638 & ~x640 & ~x723 & ~x754;
assign c6247 =  x715 & ~x368 & ~x528 & ~x606 & ~x631 & ~x632;
assign c6249 = ~x12 & ~x13 & ~x14 & ~x17 & ~x19 & ~x21 & ~x43 & ~x99 & ~x139 & ~x157 & ~x649 & ~x677 & ~x702 & ~x731 & ~x759 & ~x761 & ~x765;
assign c6251 =  x236 & ~x164 & ~x168 & ~x293 & ~x294 & ~x323 & ~x647 & ~x670 & ~x672 & ~x675 & ~x701 & ~x723 & ~x725 & ~x726 & ~x754 & ~x755 & ~x778;
assign c6253 =  x436 & ~x128 & ~x183 & ~x214 & ~x456 & ~x724;
assign c6255 =  x353 & ~x497 & ~x524 & ~x629 & ~x631;
assign c6257 =  x352 &  x377 & ~x30 & ~x32 & ~x81 & ~x83 & ~x138 & ~x139 & ~x194 & ~x216 & ~x244 & ~x246 & ~x279 & ~x281 & ~x282 & ~x303 & ~x317 & ~x327 & ~x330 & ~x335 & ~x358 & ~x373 & ~x390 & ~x392 & ~x422 & ~x423 & ~x427 & ~x428 & ~x442 & ~x445 & ~x473 & ~x502 & ~x509 & ~x531 & ~x612 & ~x614 & ~x619 & ~x672 & ~x699 & ~x753 & ~x757 & ~x761;
assign c6259 = ~x435 & ~x462 & ~x463 & ~x489 & ~x491;
assign c6261 = ~x17 & ~x43 & ~x44 & ~x72 & ~x129 & ~x420 & ~x687 & ~x714 & ~x716 & ~x717 & ~x745 & ~x773;
assign c6263 =  x84;
assign c6265 = ~x4 & ~x6 & ~x23 & ~x30 & ~x51 & ~x53 & ~x60 & ~x84 & ~x114 & ~x138 & ~x139 & ~x275 & ~x412 & ~x442 & ~x459 & ~x544 & ~x587 & ~x662 & ~x688 & ~x692 & ~x693 & ~x718 & ~x719 & ~x727;
assign c6267 =  x141;
assign c6269 =  x494 &  x521 & ~x17 & ~x53 & ~x73 & ~x221 & ~x245 & ~x258 & ~x364 & ~x476 & ~x478 & ~x643;
assign c6271 =  x175 & ~x100 & ~x155 & ~x182;
assign c6273 =  x438 & ~x388 & ~x631 & ~x632;
assign c6275 =  x743 & ~x110 & ~x139 & ~x163 & ~x215 & ~x234 & ~x261 & ~x272 & ~x299 & ~x327 & ~x391 & ~x419 & ~x456 & ~x528;
assign c6277 =  x342 & ~x577;
assign c6279 =  x139;
assign c6281 =  x349 &  x744 & ~x148 & ~x312 & ~x583;
assign c6283 =  x343 & ~x3 & ~x10 & ~x11 & ~x15 & ~x18 & ~x26 & ~x45 & ~x196 & ~x614 & ~x615 & ~x668 & ~x701 & ~x732 & ~x733 & ~x759 & ~x760 & ~x761;
assign c6285 =  x252;
assign c6287 = ~x97 & ~x355 & ~x525 & ~x527 & ~x529 & ~x625 & ~x716 & ~x717;
assign c6289 = ~x140 & ~x430 & ~x431 & ~x461 & ~x488 & ~x516 & ~x517 & ~x602;
assign c6291 =  x72 &  x127 &  x489 & ~x5 & ~x23 & ~x61 & ~x64 & ~x116 & ~x170 & ~x302 & ~x304 & ~x423 & ~x442 & ~x473 & ~x522 & ~x530 & ~x756;
assign c6293 =  x94 &  x122 &  x206 & ~x16 & ~x138 & ~x559 & ~x566 & ~x642 & ~x703;
assign c6295 =  x196;
assign c6297 =  x95 & ~x12 & ~x47 & ~x157 & ~x184;
assign c6299 =  x319 &  x371 & ~x568 & ~x598 & ~x770;
assign c6301 =  x154 & ~x56 & ~x295 & ~x296 & ~x322 & ~x509 & ~x618 & ~x674;
assign c6303 =  x181 & ~x2 & ~x19 & ~x30 & ~x33 & ~x34 & ~x47 & ~x83 & ~x89 & ~x90 & ~x92 & ~x112 & ~x138 & ~x169 & ~x176 & ~x191 & ~x200 & ~x214 & ~x215 & ~x217 & ~x229 & ~x243 & ~x253 & ~x254 & ~x258 & ~x301 & ~x302 & ~x304 & ~x305 & ~x329 & ~x357 & ~x363 & ~x365 & ~x368 & ~x386 & ~x387 & ~x390 & ~x393 & ~x412 & ~x416 & ~x422 & ~x447 & ~x448 & ~x450 & ~x451 & ~x472 & ~x506 & ~x527 & ~x557 & ~x582 & ~x613 & ~x620 & ~x641 & ~x674 & ~x696 & ~x702 & ~x725 & ~x731 & ~x751 & ~x752 & ~x753 & ~x759;
assign c6305 =  x374 & ~x59 & ~x92 & ~x107 & ~x439 & ~x441 & ~x625 & ~x652 & ~x653 & ~x676 & ~x681 & ~x696 & ~x704 & ~x705 & ~x732;
assign c6307 = ~x1 & ~x28 & ~x280 & ~x545 & ~x547 & ~x573 & ~x574 & ~x575 & ~x600 & ~x632 & ~x644;
assign c6309 =  x411 &  x651 & ~x517;
assign c6311 =  x741 & ~x146 & ~x418 & ~x453 & ~x455 & ~x481 & ~x564 & ~x658 & ~x659;
assign c6313 = ~x28 & ~x30 & ~x31 & ~x35 & ~x52 & ~x107 & ~x111 & ~x165 & ~x193 & ~x309 & ~x397 & ~x420 & ~x421 & ~x424 & ~x439 & ~x440 & ~x448 & ~x465 & ~x466 & ~x467 & ~x468 & ~x472 & ~x493 & ~x494 & ~x495 & ~x504 & ~x520 & ~x521 & ~x522 & ~x523 & ~x524 & ~x530 & ~x533 & ~x547 & ~x549 & ~x552 & ~x553 & ~x671 & ~x679 & ~x699 & ~x705 & ~x707 & ~x709 & ~x737 & ~x759 & ~x783;
assign c6315 =  x112;
assign c6317 =  x466 &  x624 & ~x189 & ~x216 & ~x305 & ~x306 & ~x359 & ~x420 & ~x481 & ~x614;
assign c6319 = ~x26 & ~x35 & ~x52 & ~x197 & ~x518 & ~x521 & ~x544 & ~x547 & ~x549;
assign c6321 =  x415 & ~x528;
assign c6323 =  x700;
assign c6325 =  x745 & ~x78 & ~x554 & ~x580 & ~x607 & ~x632;
assign c6327 =  x265 & ~x1 & ~x4 & ~x27 & ~x35 & ~x51 & ~x52 & ~x82 & ~x133 & ~x169 & ~x221 & ~x552 & ~x553 & ~x578 & ~x579 & ~x615 & ~x654 & ~x681 & ~x682 & ~x683 & ~x709 & ~x712 & ~x734;
assign c6329 =  x80;
assign c6331 =  x464 & ~x3 & ~x24 & ~x26 & ~x27 & ~x50 & ~x57 & ~x59 & ~x60 & ~x61 & ~x80 & ~x85 & ~x90 & ~x92 & ~x106 & ~x108 & ~x113 & ~x114 & ~x115 & ~x116 & ~x139 & ~x142 & ~x143 & ~x146 & ~x162 & ~x164 & ~x166 & ~x168 & ~x169 & ~x171 & ~x173 & ~x174 & ~x191 & ~x195 & ~x196 & ~x214 & ~x217 & ~x227 & ~x242 & ~x248 & ~x251 & ~x253 & ~x256 & ~x259 & ~x271 & ~x272 & ~x273 & ~x278 & ~x283 & ~x286 & ~x300 & ~x302 & ~x303 & ~x305 & ~x311 & ~x312 & ~x340 & ~x364 & ~x366 & ~x390 & ~x392 & ~x393 & ~x413 & ~x417 & ~x446 & ~x447 & ~x452 & ~x504 & ~x505 & ~x506 & ~x535 & ~x558 & ~x561 & ~x587 & ~x591 & ~x611 & ~x613 & ~x619 & ~x644 & ~x645 & ~x646 & ~x650 & ~x670 & ~x671 & ~x672 & ~x675 & ~x676 & ~x678 & ~x701 & ~x727 & ~x731 & ~x733 & ~x734 & ~x751 & ~x754 & ~x756 & ~x758 & ~x779;
assign c6333 =  x754;
assign c6335 =  x757;
assign c6337 =  x87;
assign c6339 =  x111;
assign c6341 =  x299 & ~x463;
assign c6343 =  x432 & ~x47 & ~x61 & ~x86 & ~x112 & ~x113 & ~x141 & ~x146 & ~x169 & ~x242 & ~x243 & ~x244 & ~x270 & ~x273 & ~x274 & ~x276 & ~x310 & ~x327 & ~x340 & ~x419 & ~x507 & ~x617 & ~x643 & ~x649 & ~x674 & ~x683 & ~x756;
assign c6345 =  x204 & ~x292 & ~x294 & ~x321 & ~x703 & ~x749 & ~x773;
assign c6347 =  x436 & ~x69 & ~x470 & ~x475 & ~x499 & ~x554 & ~x559 & ~x569 & ~x597 & ~x626 & ~x653 & ~x681 & ~x745;
assign c6349 =  x120 & ~x73 & ~x101 & ~x182;
assign c6351 =  x139;
assign c6353 =  x491 & ~x7 & ~x111 & ~x267 & ~x272 & ~x280 & ~x281 & ~x300 & ~x327 & ~x328 & ~x388 & ~x394 & ~x445 & ~x504 & ~x618 & ~x647 & ~x723 & ~x731 & ~x759 & ~x761 & ~x762;
assign c6355 = ~x125 & ~x299 & ~x304 & ~x332 & ~x360 & ~x361 & ~x600 & ~x661 & ~x689;
assign c6357 =  x468 & ~x21 & ~x197 & ~x250 & ~x406 & ~x407 & ~x670 & ~x751;
assign c6359 = ~x46 & ~x53 & ~x101 & ~x209 & ~x238 & ~x577;
assign c6361 =  x610 & ~x462;
assign c6363 =  x154 &  x438 & ~x216 & ~x217 & ~x225 & ~x259 & ~x260 & ~x288 & ~x362 & ~x388 & ~x390 & ~x473 & ~x589;
assign c6365 =  x1;
assign c6367 =  x323 & ~x332 & ~x361 & ~x473 & ~x631 & ~x632 & ~x658 & ~x661;
assign c6369 =  x541 & ~x61 & ~x104 & ~x130 & ~x172 & ~x250 & ~x253 & ~x277 & ~x279 & ~x287 & ~x455 & ~x528 & ~x729 & ~x730 & ~x758;
assign c6371 =  x79;
assign c6373 =  x518 & ~x5 & ~x26 & ~x27 & ~x29 & ~x116 & ~x138 & ~x439 & ~x465 & ~x542 & ~x569 & ~x588 & ~x626 & ~x654 & ~x699;
assign c6375 =  x579 & ~x460 & ~x490 & ~x491;
assign c6377 =  x40 &  x410 & ~x203 & ~x277 & ~x305;
assign c6379 =  x359 &  x419;
assign c6381 = ~x6 & ~x11 & ~x23 & ~x27 & ~x29 & ~x30 & ~x31 & ~x50 & ~x54 & ~x59 & ~x60 & ~x61 & ~x78 & ~x85 & ~x87 & ~x111 & ~x113 & ~x138 & ~x140 & ~x141 & ~x170 & ~x193 & ~x279 & ~x358 & ~x364 & ~x392 & ~x420 & ~x477 & ~x503 & ~x528 & ~x532 & ~x542 & ~x552 & ~x558 & ~x579 & ~x584 & ~x612 & ~x614 & ~x626 & ~x627 & ~x634 & ~x635 & ~x643 & ~x655 & ~x670 & ~x671 & ~x675 & ~x684 & ~x701 & ~x703 & ~x728 & ~x729 & ~x730 & ~x754 & ~x756 & ~x758 & ~x760 & ~x761 & ~x779 & ~x782 & ~x783;
assign c6383 =  x218 & ~x153 & ~x302 & ~x443 & ~x445 & ~x499 & ~x527 & ~x529;
assign c6385 =  x742 &  x743 & ~x551 & ~x604 & ~x630;
assign c6387 = ~x18 & ~x31 & ~x102 & ~x156 & ~x183 & ~x184 & ~x225 & ~x333 & ~x693 & ~x704 & ~x718 & ~x734 & ~x772;
assign c6389 = ~x16 & ~x31 & ~x51 & ~x55 & ~x58 & ~x73 & ~x74 & ~x81 & ~x86 & ~x102 & ~x114 & ~x130 & ~x131 & ~x160 & ~x185 & ~x212 & ~x223 & ~x619 & ~x645 & ~x648 & ~x649 & ~x666 & ~x670 & ~x678 & ~x679 & ~x703 & ~x731 & ~x764 & ~x778 & ~x781;
assign c6391 =  x487 &  x514 & ~x76 & ~x140 & ~x255 & ~x340 & ~x365 & ~x394 & ~x523 & ~x576;
assign c6393 =  x168;
assign c6395 =  x775 & ~x602 & ~x631;
assign c6397 =  x651 & ~x599;
assign c6399 =  x180 & ~x28 & ~x56 & ~x57 & ~x65 & ~x88 & ~x115 & ~x251 & ~x577 & ~x579 & ~x605 & ~x606 & ~x607 & ~x625 & ~x681 & ~x772;
assign c6401 =  x544 &  x717 & ~x47 & ~x77 & ~x339 & ~x606;
assign c6403 = ~x18 & ~x56 & ~x99 & ~x102 & ~x109 & ~x128 & ~x156 & ~x252 & ~x714 & ~x743 & ~x759 & ~x768;
assign c6405 =  x283 & ~x367;
assign c6407 =  x518 & ~x7 & ~x73 & ~x130 & ~x646 & ~x668 & ~x719 & ~x744 & ~x745 & ~x750 & ~x768;
assign c6409 =  x699;
assign c6411 = ~x81 & ~x404 & ~x408 & ~x409 & ~x434;
assign c6413 = ~x56 & ~x67 & ~x94 & ~x166 & ~x391 & ~x442 & ~x444 & ~x445 & ~x447 & ~x473 & ~x474 & ~x499 & ~x500 & ~x544 & ~x572 & ~x587 & ~x684 & ~x714;
assign c6415 =  x182 & ~x59 & ~x269 & ~x297 & ~x323 & ~x350 & ~x701;
assign c6417 =  x772 & ~x176 & ~x231 & ~x232 & ~x271 & ~x274 & ~x301 & ~x316 & ~x327 & ~x342 & ~x384 & ~x413 & ~x471;
assign c6419 =  x432 &  x460 &  x716 &  x717 & ~x116 & ~x331 & ~x385 & ~x412 & ~x450;
assign c6421 = ~x4 & ~x46 & ~x101 & ~x128 & ~x139 & ~x184 & ~x186 & ~x211 & ~x213 & ~x455 & ~x670 & ~x676 & ~x699 & ~x723 & ~x724 & ~x780;
assign c6423 = ~x59 & ~x224 & ~x495 & ~x524 & ~x657 & ~x711 & ~x740 & ~x770;
assign c6425 =  x649 & ~x443 & ~x446 & ~x632;
assign c6427 =  x434 & ~x25 & ~x31 & ~x69 & ~x198 & ~x236 & ~x270 & ~x310 & ~x472 & ~x525 & ~x551;
assign c6429 =  x126 &  x209 & ~x131 & ~x135 & ~x159 & ~x350 & ~x504;
assign c6431 = ~x4 & ~x21 & ~x55 & ~x83 & ~x112 & ~x459 & ~x488 & ~x515 & ~x516 & ~x542 & ~x713 & ~x718;
assign c6433 =  x126 &  x154 & ~x268 & ~x269 & ~x294;
assign c6435 =  x439 & ~x4 & ~x76 & ~x220 & ~x375 & ~x390 & ~x404 & ~x405 & ~x431 & ~x533;
assign c6437 =  x84;
assign c6439 =  x374 & ~x12 & ~x16 & ~x26 & ~x47 & ~x48 & ~x52 & ~x73 & ~x75 & ~x139 & ~x140 & ~x336 & ~x643 & ~x668 & ~x669 & ~x673 & ~x696 & ~x697 & ~x698 & ~x721 & ~x732 & ~x765 & ~x781;
assign c6441 = ~x88 & ~x414 & ~x430 & ~x469 & ~x487 & ~x488 & ~x542 & ~x545 & ~x600;
assign c6443 =  x402 &  x430 & ~x253 & ~x412 & ~x439 & ~x496 & ~x626 & ~x731;
assign c6445 = ~x73 & ~x82 & ~x130 & ~x183 & ~x211 & ~x240 & ~x385 & ~x723 & ~x750;
assign c6447 =  x208 &  x491 & ~x0 & ~x21 & ~x32 & ~x51 & ~x53 & ~x56 & ~x62 & ~x78 & ~x84 & ~x86 & ~x107 & ~x116 & ~x144 & ~x145 & ~x196 & ~x197 & ~x214 & ~x220 & ~x223 & ~x228 & ~x243 & ~x245 & ~x246 & ~x247 & ~x248 & ~x254 & ~x255 & ~x274 & ~x276 & ~x279 & ~x281 & ~x300 & ~x304 & ~x306 & ~x307 & ~x333 & ~x335 & ~x362 & ~x391 & ~x392 & ~x422 & ~x449 & ~x478 & ~x613 & ~x642 & ~x669 & ~x670 & ~x672 & ~x697 & ~x727 & ~x753 & ~x783;
assign c6449 = ~x30 & ~x54 & ~x80 & ~x85 & ~x168 & ~x300 & ~x328 & ~x385 & ~x386 & ~x413 & ~x415 & ~x430 & ~x443 & ~x470 & ~x487 & ~x571 & ~x626 & ~x627 & ~x656 & ~x675 & ~x723;
assign c6451 =  x111;
assign c6453 =  x267 & ~x24 & ~x247 & ~x281 & ~x460 & ~x659 & ~x690;
assign c6455 =  x206 & ~x320 & ~x323 & ~x376 & ~x673 & ~x723;
assign c6457 =  x495 & ~x75 & ~x433 & ~x459;
assign c6459 =  x437 &  x465 &  x743 & ~x0 & ~x308 & ~x327 & ~x341 & ~x367 & ~x384 & ~x456 & ~x504 & ~x532 & ~x722 & ~x778;
assign c6461 =  x150 & ~x89 & ~x294 & ~x321 & ~x424 & ~x453 & ~x477 & ~x504 & ~x533 & ~x558 & ~x667 & ~x668 & ~x701 & ~x727;
assign c6463 =  x259 & ~x99 & ~x127 & ~x290;
assign c6465 =  x125 &  x346 & ~x15 & ~x19 & ~x130 & ~x642 & ~x670;
assign c6467 =  x742 & ~x24 & ~x35 & ~x192 & ~x223 & ~x330 & ~x415 & ~x442 & ~x500 & ~x531 & ~x558 & ~x611 & ~x659 & ~x751;
assign c6469 =  x72 & ~x4 & ~x83 & ~x301 & ~x328 & ~x329 & ~x331 & ~x332 & ~x359 & ~x386 & ~x414 & ~x415 & ~x532 & ~x542 & ~x570 & ~x599 & ~x608 & ~x627 & ~x647 & ~x656 & ~x763;
assign c6471 =  x438 &  x466 &  x494 & ~x25 & ~x26 & ~x57 & ~x60 & ~x83 & ~x120 & ~x148 & ~x170 & ~x330 & ~x336 & ~x344 & ~x359 & ~x362 & ~x389 & ~x414 & ~x421 & ~x423 & ~x502 & ~x506 & ~x586 & ~x701 & ~x729;
assign c6473 =  x151 & ~x0 & ~x23 & ~x46 & ~x50 & ~x58 & ~x60 & ~x80 & ~x85 & ~x102 & ~x103 & ~x106 & ~x114 & ~x134 & ~x144 & ~x156 & ~x157 & ~x159 & ~x160 & ~x162 & ~x166 & ~x169 & ~x186 & ~x188 & ~x192 & ~x216 & ~x252 & ~x336 & ~x559 & ~x590 & ~x643 & ~x646 & ~x694 & ~x697 & ~x699 & ~x720 & ~x721 & ~x730 & ~x750 & ~x756 & ~x758 & ~x778 & ~x782;
assign c6475 =  x111;
assign c6477 =  x318 & ~x17 & ~x47 & ~x211 & ~x213 & ~x760;
assign c6479 = ~x98 & ~x126 & ~x235 & ~x277 & ~x660 & ~x689;
assign c6481 =  x741 & ~x160 & ~x244 & ~x426 & ~x454 & ~x529 & ~x657 & ~x693;
assign c6483 = ~x18 & ~x70 & ~x99 & ~x168 & ~x448 & ~x643 & ~x663 & ~x688 & ~x717 & ~x719 & ~x720 & ~x768;
assign c6485 =  x354 &  x410 &  x411 & ~x204 & ~x304;
assign c6487 =  x401 &  x456 & ~x497 & ~x655 & ~x712;
assign c6489 =  x161 & ~x97 & ~x98 & ~x125 & ~x300 & ~x389 & ~x442 & ~x445 & ~x571;
assign c6491 = ~x5 & ~x27 & ~x36 & ~x68 & ~x111 & ~x145 & ~x299 & ~x355 & ~x383 & ~x470 & ~x495 & ~x502 & ~x523 & ~x524 & ~x529 & ~x530 & ~x531 & ~x558 & ~x579 & ~x580 & ~x613 & ~x617 & ~x626 & ~x675 & ~x706 & ~x711 & ~x733 & ~x734 & ~x739 & ~x765;
assign c6493 =  x715 &  x716 & ~x104 & ~x146 & ~x172 & ~x367 & ~x369 & ~x444 & ~x475 & ~x503;
assign c6495 =  x165;
assign c6497 = ~x401 & ~x460 & ~x461 & ~x462 & ~x488 & ~x490 & ~x491 & ~x692 & ~x720 & ~x747;
assign c6499 =  x468 & ~x407 & ~x433;
assign c70 = ~x5 & ~x32 & ~x34 & ~x70 & ~x71 & ~x84 & ~x91 & ~x106 & ~x112 & ~x145 & ~x161 & ~x162 & ~x196 & ~x223 & ~x224 & ~x506 & ~x509 & ~x535 & ~x561 & ~x564 & ~x677 & ~x692 & ~x718 & ~x738 & ~x739 & ~x764 & ~x767;
assign c72 =  x574 &  x764;
assign c74 = ~x18 & ~x20 & ~x50 & ~x83 & ~x85 & ~x483 & ~x511 & ~x523 & ~x524 & ~x539 & ~x540 & ~x551 & ~x556 & ~x568 & ~x570 & ~x580 & ~x581 & ~x583 & ~x587 & ~x589 & ~x597 & ~x615 & ~x702 & ~x731;
assign c76 =  x456 & ~x2 & ~x51 & ~x56 & ~x80 & ~x81 & ~x82 & ~x84 & ~x110 & ~x111 & ~x115 & ~x129 & ~x133 & ~x134 & ~x135 & ~x141 & ~x161 & ~x164 & ~x166 & ~x190 & ~x195 & ~x582 & ~x611 & ~x642 & ~x668 & ~x669 & ~x697 & ~x725 & ~x726 & ~x727 & ~x750 & ~x760 & ~x775 & ~x776 & ~x777 & ~x778 & ~x779 & ~x782;
assign c78 =  x43 &  x400 &  x457 & ~x11;
assign c710 =  x515 & ~x79 & ~x81 & ~x137 & ~x143 & ~x161 & ~x250 & ~x382 & ~x623 & ~x635 & ~x644 & ~x650 & ~x678 & ~x696 & ~x704;
assign c712 =  x518 &  x573 &  x662 & ~x130 & ~x142 & ~x158 & ~x159 & ~x199 & ~x228 & ~x254 & ~x257 & ~x284 & ~x310 & ~x339 & ~x365 & ~x367 & ~x394 & ~x613 & ~x614 & ~x696 & ~x697 & ~x700;
assign c714 =  x286 & ~x5 & ~x87 & ~x224 & ~x392 & ~x502 & ~x510 & ~x527 & ~x530 & ~x537 & ~x538 & ~x558 & ~x576 & ~x591 & ~x619 & ~x650 & ~x698 & ~x702 & ~x734 & ~x757 & ~x758 & ~x761 & ~x773;
assign c716 = ~x4 & ~x452 & ~x474 & ~x506 & ~x562 & ~x566 & ~x575 & ~x576 & ~x579 & ~x607 & ~x635 & ~x644 & ~x660 & ~x661 & ~x665 & ~x666 & ~x674 & ~x678 & ~x702 & ~x718 & ~x723 & ~x732 & ~x749 & ~x755 & ~x761 & ~x774 & ~x776;
assign c718 =  x2;
assign c720 =  x17 &  x252;
assign c722 =  x265 &  x266 & ~x0 & ~x1 & ~x11 & ~x28 & ~x112 & ~x113 & ~x114 & ~x169 & ~x475 & ~x552 & ~x553 & ~x554 & ~x558 & ~x580 & ~x595 & ~x613 & ~x669 & ~x680 & ~x708 & ~x761 & ~x762;
assign c724 =  x352 &  x429 &  x543 & ~x171 & ~x247 & ~x699;
assign c726 =  x189 &  x190 & ~x499 & ~x506 & ~x527 & ~x528 & ~x534 & ~x576 & ~x617 & ~x702 & ~x746;
assign c728 = ~x7 & ~x38 & ~x39 & ~x44 & ~x48 & ~x55 & ~x59 & ~x86 & ~x166 & ~x191 & ~x197 & ~x222 & ~x509 & ~x510 & ~x511 & ~x536 & ~x557 & ~x562 & ~x563 & ~x591 & ~x610 & ~x612 & ~x640 & ~x652 & ~x664 & ~x680 & ~x694 & ~x710 & ~x718 & ~x721 & ~x722 & ~x733 & ~x749 & ~x752 & ~x753;
assign c730 =  x323 &  x482 & ~x4 & ~x9 & ~x10 & ~x30 & ~x31 & ~x57 & ~x81 & ~x82 & ~x84 & ~x88 & ~x89 & ~x106 & ~x109 & ~x111 & ~x113 & ~x115 & ~x133 & ~x135 & ~x138 & ~x139 & ~x140 & ~x142 & ~x165 & ~x168 & ~x169 & ~x170 & ~x171 & ~x189 & ~x190 & ~x192 & ~x194 & ~x195 & ~x196 & ~x224 & ~x252 & ~x253 & ~x280 & ~x281 & ~x641 & ~x668 & ~x699 & ~x726 & ~x727 & ~x729 & ~x754 & ~x757 & ~x760 & ~x774 & ~x775 & ~x777 & ~x783;
assign c732 =  x461 & ~x29 & ~x435 & ~x485 & ~x504 & ~x571 & ~x572 & ~x599 & ~x600 & ~x614 & ~x620 & ~x621 & ~x647 & ~x657 & ~x672 & ~x683 & ~x685 & ~x699 & ~x706 & ~x712 & ~x724 & ~x732 & ~x760 & ~x765 & ~x766;
assign c734 =  x353 & ~x2 & ~x3 & ~x7 & ~x10 & ~x31 & ~x35 & ~x57 & ~x61 & ~x64 & ~x75 & ~x103 & ~x112 & ~x116 & ~x117 & ~x139 & ~x141 & ~x170 & ~x171 & ~x172 & ~x197 & ~x198 & ~x199 & ~x200 & ~x201 & ~x226 & ~x253 & ~x284 & ~x616 & ~x714 & ~x732 & ~x733 & ~x734 & ~x753 & ~x761 & ~x779 & ~x781;
assign c736 =  x508 & ~x25 & ~x114 & ~x129 & ~x196 & ~x201 & ~x245 & ~x284 & ~x310 & ~x312 & ~x364 & ~x595 & ~x677 & ~x757 & ~x777;
assign c738 =  x208 &  x327 & ~x470 & ~x623;
assign c740 =  x83 &  x157;
assign c742 =  x204 &  x233 & ~x19 & ~x27 & ~x50 & ~x416 & ~x432 & ~x467 & ~x477 & ~x507 & ~x535 & ~x561 & ~x633 & ~x673;
assign c744 =  x263 &  x325 &  x510 &  x543 & ~x86 & ~x141 & ~x158 & ~x226 & ~x672 & ~x756;
assign c746 = ~x475 & ~x483 & ~x484 & ~x497 & ~x527 & ~x528 & ~x536 & ~x539 & ~x547 & ~x569 & ~x595 & ~x632 & ~x648 & ~x652 & ~x707 & ~x765;
assign c748 =  x70 &  x72 &  x321 &  x347;
assign c750 =  x251;
assign c752 =  x371 &  x544 & ~x0 & ~x54 & ~x58 & ~x143 & ~x196 & ~x252 & ~x336 & ~x586 & ~x596 & ~x624 & ~x642 & ~x669 & ~x671 & ~x697 & ~x706 & ~x707 & ~x760 & ~x778;
assign c754 =  x444 & ~x24 & ~x26 & ~x77 & ~x82 & ~x84 & ~x107 & ~x108 & ~x132 & ~x134 & ~x135 & ~x159 & ~x161 & ~x166 & ~x187 & ~x188 & ~x189 & ~x191 & ~x194 & ~x221 & ~x249 & ~x279 & ~x307 & ~x565 & ~x587 & ~x613 & ~x615 & ~x620 & ~x622 & ~x637 & ~x640 & ~x641 & ~x666 & ~x668 & ~x669 & ~x694 & ~x697 & ~x702 & ~x723 & ~x728 & ~x751 & ~x753 & ~x754 & ~x755 & ~x757 & ~x759 & ~x778 & ~x782 & ~x783;
assign c756 =  x343 &  x690 & ~x142 & ~x338 & ~x421 & ~x595 & ~x622 & ~x649;
assign c758 =  x66 &  x461 &  x518 & ~x6 & ~x384 & ~x447 & ~x643 & ~x668 & ~x725;
assign c760 =  x210 &  x234 & ~x4 & ~x26 & ~x27 & ~x28 & ~x46 & ~x56 & ~x74 & ~x83 & ~x500 & ~x523 & ~x524 & ~x527 & ~x530 & ~x553 & ~x561 & ~x588 & ~x611 & ~x682 & ~x701 & ~x727;
assign c762 = ~x2 & ~x19 & ~x97 & ~x225 & ~x273 & ~x282 & ~x423 & ~x558 & ~x608 & ~x656 & ~x719 & ~x740 & ~x753 & ~x760;
assign c764 =  x448;
assign c766 =  x486 & ~x0 & ~x9 & ~x25 & ~x28 & ~x30 & ~x31 & ~x33 & ~x34 & ~x35 & ~x50 & ~x51 & ~x83 & ~x84 & ~x85 & ~x166 & ~x167 & ~x170 & ~x252 & ~x568 & ~x595 & ~x596 & ~x622 & ~x623 & ~x624 & ~x641 & ~x644 & ~x652 & ~x653 & ~x673 & ~x678 & ~x700 & ~x706 & ~x725 & ~x726 & ~x727 & ~x730 & ~x733 & ~x734 & ~x735 & ~x760 & ~x761 & ~x762 & ~x777 & ~x779;
assign c768 =  x559;
assign c770 =  x401 &  x486 &  x516 & ~x1 & ~x9 & ~x57 & ~x89 & ~x142 & ~x143 & ~x171 & ~x197 & ~x225 & ~x281 & ~x504 & ~x613 & ~x641 & ~x670 & ~x697 & ~x707 & ~x720 & ~x762;
assign c772 = ~x2 & ~x14 & ~x16 & ~x25 & ~x28 & ~x29 & ~x43 & ~x58 & ~x83 & ~x84 & ~x86 & ~x88 & ~x112 & ~x141 & ~x160 & ~x170 & ~x195 & ~x197 & ~x501 & ~x528 & ~x558 & ~x568 & ~x585 & ~x586 & ~x595 & ~x624 & ~x642 & ~x651 & ~x652 & ~x679 & ~x705 & ~x729 & ~x754 & ~x755 & ~x760;
assign c774 =  x55;
assign c776 = ~x2 & ~x6 & ~x9 & ~x19 & ~x23 & ~x24 & ~x25 & ~x46 & ~x48 & ~x57 & ~x109 & ~x111 & ~x113 & ~x196 & ~x280 & ~x308 & ~x530 & ~x556 & ~x558 & ~x559 & ~x573 & ~x587 & ~x593 & ~x617 & ~x630 & ~x647 & ~x671 & ~x673 & ~x681 & ~x715 & ~x717 & ~x721 & ~x729 & ~x754 & ~x757 & ~x759 & ~x760 & ~x763 & ~x773 & ~x781;
assign c778 =  x474 & ~x13 & ~x111 & ~x171 & ~x172 & ~x174 & ~x192 & ~x198 & ~x217 & ~x226 & ~x244 & ~x246 & ~x277 & ~x637 & ~x755;
assign c780 = ~x50 & ~x56 & ~x113 & ~x396 & ~x423 & ~x447 & ~x512 & ~x530 & ~x537 & ~x555 & ~x556 & ~x557 & ~x564 & ~x566 & ~x569 & ~x588 & ~x589 & ~x591 & ~x620 & ~x625 & ~x632 & ~x644 & ~x647 & ~x650 & ~x653 & ~x660 & ~x681 & ~x698 & ~x703 & ~x716 & ~x717 & ~x728 & ~x730 & ~x735 & ~x737 & ~x764 & ~x765;
assign c782 =  x545 & ~x4 & ~x109 & ~x578 & ~x597 & ~x608 & ~x627 & ~x636 & ~x655 & ~x667 & ~x704 & ~x711 & ~x712 & ~x737 & ~x782;
assign c784 = ~x3 & ~x15 & ~x27 & ~x41 & ~x42 & ~x43 & ~x69 & ~x76 & ~x83 & ~x90 & ~x92 & ~x96 & ~x114 & ~x135 & ~x146 & ~x147 & ~x169 & ~x170 & ~x175 & ~x190 & ~x197 & ~x198 & ~x223 & ~x225 & ~x226 & ~x253 & ~x254 & ~x596 & ~x624 & ~x638 & ~x646 & ~x647 & ~x670 & ~x680 & ~x695 & ~x699 & ~x703 & ~x720 & ~x728 & ~x729 & ~x730 & ~x731 & ~x753 & ~x757 & ~x760 & ~x775 & ~x778;
assign c786 =  x363 &  x417 & ~x310 & ~x529;
assign c788 = ~x32 & ~x54 & ~x140 & ~x141 & ~x169 & ~x381 & ~x383 & ~x384 & ~x511 & ~x568 & ~x580 & ~x581 & ~x582 & ~x583 & ~x584 & ~x593 & ~x594 & ~x610 & ~x613 & ~x614 & ~x638 & ~x651 & ~x652 & ~x656 & ~x678 & ~x701 & ~x710 & ~x728 & ~x734 & ~x736 & ~x740 & ~x783;
assign c790 =  x374 &  x459 & ~x112 & ~x168 & ~x513 & ~x540 & ~x541 & ~x569 & ~x596 & ~x597 & ~x598 & ~x623 & ~x653 & ~x678 & ~x680 & ~x681 & ~x707 & ~x732 & ~x737 & ~x759 & ~x761 & ~x763 & ~x766;
assign c792 = ~x11 & ~x41 & ~x55 & ~x91 & ~x110 & ~x111 & ~x115 & ~x117 & ~x129 & ~x199 & ~x218 & ~x227 & ~x281 & ~x288 & ~x669 & ~x677 & ~x678 & ~x697 & ~x706 & ~x720 & ~x740 & ~x745 & ~x748 & ~x780;
assign c794 =  x290 &  x325 &  x345 &  x346 &  x374 &  x430 & ~x36 & ~x83 & ~x85 & ~x115 & ~x116 & ~x142 & ~x705 & ~x758 & ~x763;
assign c798 =  x538 & ~x3 & ~x4 & ~x23 & ~x25 & ~x27 & ~x31 & ~x57 & ~x60 & ~x102 & ~x103 & ~x105 & ~x113 & ~x129 & ~x135 & ~x138 & ~x139 & ~x196 & ~x198 & ~x280 & ~x286 & ~x312 & ~x313 & ~x392 & ~x422 & ~x587 & ~x726 & ~x754 & ~x775;
assign c7100 = ~x26 & ~x34 & ~x451 & ~x531 & ~x544 & ~x545 & ~x552 & ~x555 & ~x569 & ~x601 & ~x608 & ~x617 & ~x640 & ~x654 & ~x670 & ~x673;
assign c7102 =  x476;
assign c7104 =  x375 &  x383 & ~x31 & ~x144 & ~x170 & ~x174 & ~x196 & ~x282 & ~x641 & ~x746;
assign c7106 =  x378 & ~x2 & ~x3 & ~x92 & ~x140 & ~x147 & ~x160 & ~x164 & ~x173 & ~x199 & ~x255 & ~x257 & ~x280 & ~x555 & ~x586 & ~x641 & ~x674 & ~x687 & ~x714 & ~x742;
assign c7108 =  x292 &  x444 & ~x11 & ~x191 & ~x582 & ~x586 & ~x608 & ~x610 & ~x611 & ~x639 & ~x641 & ~x650 & ~x669 & ~x678 & ~x705 & ~x727 & ~x758;
assign c7110 =  x176 & ~x1 & ~x3 & ~x25 & ~x511 & ~x539 & ~x565 & ~x567 & ~x570 & ~x584 & ~x593 & ~x612 & ~x619 & ~x625 & ~x626 & ~x627 & ~x653 & ~x654 & ~x676 & ~x678 & ~x683 & ~x702 & ~x710 & ~x725 & ~x728 & ~x737 & ~x739 & ~x767;
assign c7112 =  x399 &  x458 &  x515 & ~x132 & ~x540;
assign c7114 =  x204 & ~x55 & ~x452 & ~x478 & ~x492 & ~x506 & ~x507 & ~x509 & ~x538 & ~x563 & ~x585 & ~x592 & ~x593 & ~x605 & ~x637 & ~x662 & ~x673 & ~x693 & ~x748 & ~x760 & ~x781;
assign c7116 = ~x58 & ~x85 & ~x513 & ~x527 & ~x528 & ~x529 & ~x530 & ~x532 & ~x535 & ~x550 & ~x552 & ~x562 & ~x564 & ~x570 & ~x571 & ~x590 & ~x592 & ~x598 & ~x599 & ~x607 & ~x610 & ~x615 & ~x625 & ~x643 & ~x646 & ~x669 & ~x670 & ~x674 & ~x696 & ~x711 & ~x721 & ~x727 & ~x754 & ~x756 & ~x759 & ~x765 & ~x768 & ~x769 & ~x783;
assign c7118 = ~x0 & ~x2 & ~x14 & ~x27 & ~x57 & ~x61 & ~x64 & ~x67 & ~x103 & ~x146 & ~x248 & ~x534 & ~x564 & ~x605 & ~x621 & ~x700 & ~x703 & ~x728 & ~x756 & ~x762;
assign c7120 = ~x57 & ~x351 & ~x380 & ~x391 & ~x419 & ~x446 & ~x454 & ~x470 & ~x472 & ~x495 & ~x500 & ~x511 & ~x525 & ~x528 & ~x567 & ~x594 & ~x595 & ~x637 & ~x650 & ~x673 & ~x729 & ~x732 & ~x759;
assign c7122 = ~x7 & ~x35 & ~x59 & ~x117 & ~x447 & ~x480 & ~x524 & ~x529 & ~x550 & ~x571 & ~x607 & ~x643 & ~x665 & ~x682 & ~x778;
assign c7124 = ~x7 & ~x19 & ~x20 & ~x22 & ~x23 & ~x25 & ~x28 & ~x47 & ~x55 & ~x86 & ~x112 & ~x434 & ~x452 & ~x480 & ~x504 & ~x507 & ~x508 & ~x528 & ~x529 & ~x535 & ~x548 & ~x558 & ~x577 & ~x588 & ~x590 & ~x591 & ~x613 & ~x616 & ~x617 & ~x645 & ~x674 & ~x675 & ~x697 & ~x719 & ~x720 & ~x725 & ~x728 & ~x730 & ~x731 & ~x749 & ~x753 & ~x761 & ~x763 & ~x783;
assign c7126 = ~x4 & ~x27 & ~x196 & ~x353 & ~x474 & ~x475 & ~x500 & ~x501 & ~x524 & ~x528 & ~x530 & ~x571 & ~x580 & ~x581 & ~x583 & ~x644 & ~x666 & ~x674 & ~x675 & ~x676 & ~x684 & ~x685 & ~x701 & ~x728 & ~x757 & ~x767 & ~x772;
assign c7128 =  x600 & ~x130 & ~x131 & ~x160 & ~x161 & ~x171 & ~x188 & ~x199 & ~x202 & ~x230 & ~x255 & ~x257 & ~x283 & ~x301 & ~x312 & ~x313 & ~x332 & ~x340 & ~x422 & ~x448 & ~x761;
assign c7130 = ~x30 & ~x80 & ~x81 & ~x484 & ~x500 & ~x509 & ~x512 & ~x527 & ~x528 & ~x532 & ~x536 & ~x537 & ~x538 & ~x555 & ~x556 & ~x560 & ~x562 & ~x563 & ~x564 & ~x569 & ~x572 & ~x584 & ~x585 & ~x588 & ~x589 & ~x650 & ~x654 & ~x658 & ~x709;
assign c7132 =  x236 & ~x500 & ~x502 & ~x503 & ~x526 & ~x527 & ~x557 & ~x564 & ~x600 & ~x628 & ~x648 & ~x656 & ~x741 & ~x748 & ~x757 & ~x760 & ~x768;
assign c7134 =  x388 &  x389 & ~x53 & ~x198 & ~x332 & ~x705 & ~x778;
assign c7136 =  x420;
assign c7138 =  x615;
assign c7140 =  x412 & ~x232 & ~x255 & ~x258 & ~x312 & ~x365 & ~x497 & ~x698 & ~x780;
assign c7142 =  x466 & ~x6 & ~x7 & ~x24 & ~x25 & ~x32 & ~x33 & ~x37 & ~x47 & ~x50 & ~x55 & ~x57 & ~x65 & ~x68 & ~x77 & ~x82 & ~x91 & ~x105 & ~x119 & ~x133 & ~x135 & ~x138 & ~x139 & ~x147 & ~x226 & ~x253 & ~x254 & ~x645 & ~x704 & ~x706 & ~x719 & ~x721 & ~x735 & ~x746 & ~x761 & ~x769 & ~x775 & ~x779 & ~x780;
assign c7144 =  x783;
assign c7146 =  x508 & ~x171 & ~x199 & ~x226 & ~x227 & ~x255 & ~x256 & ~x257 & ~x258 & ~x301 & ~x302 & ~x338 & ~x339 & ~x622;
assign c7148 = ~x52 & ~x56 & ~x62 & ~x64 & ~x70 & ~x86 & ~x103 & ~x118 & ~x144 & ~x165 & ~x173 & ~x177 & ~x191 & ~x196 & ~x218 & ~x230 & ~x475 & ~x503 & ~x584 & ~x585 & ~x698 & ~x730 & ~x751;
assign c7150 =  x374 &  x429 &  x457 & ~x2 & ~x8 & ~x9 & ~x27 & ~x30 & ~x31 & ~x63 & ~x64 & ~x82 & ~x88 & ~x89 & ~x111 & ~x114 & ~x117 & ~x118 & ~x142 & ~x143 & ~x144 & ~x162 & ~x163 & ~x166 & ~x167 & ~x170 & ~x194 & ~x252 & ~x281 & ~x308 & ~x586 & ~x615 & ~x641 & ~x642 & ~x725 & ~x775 & ~x776;
assign c7152 =  x94 &  x206 &  x289 &  x426 & ~x641;
assign c7154 =  x265 & ~x4 & ~x9 & ~x26 & ~x89 & ~x109 & ~x115 & ~x117 & ~x139 & ~x196 & ~x336 & ~x503 & ~x555 & ~x557 & ~x558 & ~x559 & ~x570 & ~x585 & ~x597 & ~x628 & ~x639 & ~x656 & ~x657 & ~x658 & ~x668 & ~x677 & ~x678 & ~x683 & ~x712 & ~x735 & ~x739 & ~x752 & ~x753 & ~x755 & ~x756;
assign c7156 =  x402 & ~x1 & ~x3 & ~x24 & ~x25 & ~x27 & ~x42 & ~x106 & ~x109 & ~x136 & ~x140 & ~x141 & ~x163 & ~x165 & ~x557 & ~x567 & ~x586 & ~x595 & ~x597 & ~x610 & ~x625 & ~x626 & ~x650 & ~x651 & ~x652 & ~x653 & ~x668 & ~x669 & ~x677 & ~x698 & ~x707 & ~x709 & ~x710 & ~x727 & ~x729 & ~x732 & ~x734 & ~x753 & ~x755 & ~x756 & ~x757 & ~x762 & ~x763 & ~x765 & ~x783;
assign c7158 = ~x4 & ~x5 & ~x19 & ~x29 & ~x32 & ~x54 & ~x113 & ~x335 & ~x390 & ~x391 & ~x417 & ~x418 & ~x445 & ~x448 & ~x460 & ~x469 & ~x470 & ~x475 & ~x478 & ~x488 & ~x495 & ~x499 & ~x524 & ~x528 & ~x530 & ~x532 & ~x535 & ~x546 & ~x552 & ~x554 & ~x560 & ~x561 & ~x562 & ~x581 & ~x583 & ~x584 & ~x587 & ~x613 & ~x618 & ~x619 & ~x647 & ~x671 & ~x674 & ~x697 & ~x702 & ~x758 & ~x782 & ~x783;
assign c7160 =  x408 & ~x1 & ~x3 & ~x17 & ~x25 & ~x26 & ~x30 & ~x31 & ~x89 & ~x101 & ~x102 & ~x115 & ~x116 & ~x130 & ~x132 & ~x158 & ~x172 & ~x196 & ~x197 & ~x198 & ~x200 & ~x201 & ~x225 & ~x228 & ~x229 & ~x254 & ~x255 & ~x279 & ~x280 & ~x285 & ~x308 & ~x311 & ~x336 & ~x338 & ~x340 & ~x365 & ~x366 & ~x392 & ~x394 & ~x420 & ~x423 & ~x447 & ~x448 & ~x477 & ~x504 & ~x505 & ~x560 & ~x642 & ~x699 & ~x727 & ~x728 & ~x754 & ~x758;
assign c7162 = ~x24 & ~x25 & ~x26 & ~x30 & ~x31 & ~x55 & ~x82 & ~x474 & ~x508 & ~x533 & ~x534 & ~x547 & ~x550 & ~x562 & ~x564 & ~x586 & ~x645 & ~x647 & ~x661 & ~x665 & ~x673 & ~x679 & ~x703 & ~x707 & ~x717 & ~x719 & ~x730 & ~x731 & ~x754 & ~x755 & ~x760 & ~x763 & ~x765 & ~x774;
assign c7164 =  x154 &  x155 &  x237 & ~x566 & ~x567;
assign c7166 =  x546 & ~x7 & ~x13 & ~x26 & ~x27 & ~x33 & ~x35 & ~x56 & ~x85 & ~x91 & ~x103 & ~x118 & ~x130 & ~x139 & ~x169 & ~x232 & ~x255 & ~x257 & ~x281 & ~x587 & ~x669 & ~x757;
assign c7168 =  x359 & ~x31 & ~x113 & ~x114 & ~x141 & ~x145 & ~x443 & ~x444 & ~x468 & ~x471 & ~x497 & ~x698 & ~x719 & ~x777;
assign c7170 =  x362 & ~x9 & ~x17 & ~x20 & ~x22 & ~x30 & ~x31 & ~x47 & ~x51 & ~x52 & ~x60 & ~x63 & ~x81 & ~x82 & ~x106 & ~x135 & ~x162 & ~x164 & ~x165 & ~x223 & ~x357 & ~x556 & ~x565 & ~x582 & ~x584 & ~x593 & ~x614 & ~x638 & ~x648 & ~x649 & ~x667 & ~x700 & ~x703 & ~x705 & ~x729 & ~x731 & ~x751 & ~x753 & ~x756 & ~x760 & ~x763 & ~x778 & ~x779;
assign c7172 = ~x455 & ~x457 & ~x468 & ~x475 & ~x486 & ~x498 & ~x501 & ~x509 & ~x516 & ~x529 & ~x536 & ~x557 & ~x564 & ~x566 & ~x589 & ~x594 & ~x619 & ~x627 & ~x641 & ~x646 & ~x672 & ~x680 & ~x682 & ~x707 & ~x756 & ~x759;
assign c7174 =  x270 &  x319 & ~x1 & ~x3 & ~x4 & ~x8 & ~x9 & ~x11 & ~x22 & ~x23 & ~x27 & ~x54 & ~x62 & ~x87 & ~x114 & ~x174 & ~x308 & ~x624 & ~x643 & ~x670 & ~x679 & ~x698 & ~x706 & ~x734 & ~x748 & ~x757 & ~x772 & ~x777 & ~x778 & ~x783;
assign c7176 =  x124 &  x391;
assign c7178 =  x27;
assign c7180 =  x516 & ~x29 & ~x41 & ~x103 & ~x104 & ~x113 & ~x171 & ~x172 & ~x183 & ~x197 & ~x198 & ~x199 & ~x200 & ~x226 & ~x254 & ~x256 & ~x282 & ~x308 & ~x311 & ~x475 & ~x502 & ~x614 & ~x760;
assign c7182 =  x124 &  x502 & ~x313;
assign c7184 =  x280;
assign c7186 =  x238 & ~x31 & ~x50 & ~x53 & ~x70 & ~x79 & ~x83 & ~x136 & ~x164 & ~x352 & ~x509 & ~x565 & ~x591 & ~x594 & ~x622 & ~x644 & ~x647 & ~x665 & ~x672 & ~x673 & ~x674 & ~x697 & ~x702 & ~x723 & ~x749 & ~x750 & ~x764 & ~x782;
assign c7188 = ~x85 & ~x419 & ~x435 & ~x446 & ~x465 & ~x466 & ~x469 & ~x480 & ~x498 & ~x521 & ~x527 & ~x551 & ~x558 & ~x559 & ~x562 & ~x563 & ~x606 & ~x612 & ~x668 & ~x727 & ~x749 & ~x750 & ~x764 & ~x765;
assign c7190 = ~x9 & ~x19 & ~x24 & ~x26 & ~x58 & ~x86 & ~x472 & ~x500 & ~x501 & ~x507 & ~x515 & ~x517 & ~x527 & ~x532 & ~x533 & ~x536 & ~x557 & ~x574 & ~x591 & ~x601 & ~x602 & ~x617 & ~x619 & ~x625 & ~x652 & ~x731 & ~x737 & ~x766;
assign c7192 = ~x2 & ~x7 & ~x12 & ~x21 & ~x36 & ~x37 & ~x71 & ~x78 & ~x87 & ~x117 & ~x142 & ~x143 & ~x169 & ~x171 & ~x189 & ~x216 & ~x222 & ~x223 & ~x225 & ~x226 & ~x567 & ~x586 & ~x596 & ~x613 & ~x615 & ~x620 & ~x622 & ~x625 & ~x637 & ~x641 & ~x672 & ~x673 & ~x677 & ~x701 & ~x721 & ~x722 & ~x756 & ~x767 & ~x774 & ~x775 & ~x776;
assign c7194 =  x518 &  x654 & ~x75 & ~x130 & ~x158 & ~x171 & ~x200 & ~x201 & ~x254 & ~x255 & ~x256 & ~x257 & ~x279 & ~x284 & ~x285 & ~x311 & ~x313 & ~x423 & ~x449;
assign c7196 =  x251;
assign c7198 =  x153 &  x603 &  x722 & ~x555;
assign c7200 =  x122 &  x317 &  x769;
assign c7202 = ~x2 & ~x3 & ~x4 & ~x20 & ~x24 & ~x26 & ~x29 & ~x57 & ~x58 & ~x81 & ~x84 & ~x106 & ~x111 & ~x114 & ~x447 & ~x474 & ~x502 & ~x532 & ~x537 & ~x562 & ~x564 & ~x576 & ~x577 & ~x584 & ~x588 & ~x591 & ~x606 & ~x607 & ~x614 & ~x615 & ~x616 & ~x617 & ~x633 & ~x646 & ~x648 & ~x649 & ~x673 & ~x675 & ~x691 & ~x698 & ~x703 & ~x719 & ~x721 & ~x726 & ~x729 & ~x753 & ~x756 & ~x757 & ~x764 & ~x767;
assign c7204 =  x249 & ~x0 & ~x5 & ~x22 & ~x24 & ~x25 & ~x28 & ~x31 & ~x56 & ~x57 & ~x58 & ~x59 & ~x84 & ~x85 & ~x112 & ~x113 & ~x419 & ~x444 & ~x445 & ~x446 & ~x470 & ~x472 & ~x494 & ~x497 & ~x498 & ~x499 & ~x501 & ~x526 & ~x531 & ~x596 & ~x624 & ~x673 & ~x701 & ~x702 & ~x730 & ~x783;
assign c7206 =  x429 &  x463 & ~x1 & ~x8 & ~x9 & ~x11 & ~x35 & ~x54 & ~x56 & ~x61 & ~x82 & ~x83 & ~x111 & ~x117 & ~x135 & ~x144 & ~x145 & ~x146 & ~x165 & ~x168 & ~x169 & ~x170 & ~x172 & ~x173 & ~x191 & ~x194 & ~x198 & ~x202 & ~x228 & ~x254 & ~x641 & ~x643 & ~x696 & ~x699 & ~x706 & ~x759 & ~x773 & ~x776 & ~x781;
assign c7208 =  x241 &  x361 & ~x327 & ~x475 & ~x503 & ~x530 & ~x553 & ~x555 & ~x642 & ~x705 & ~x753;
assign c7210 =  x352 &  x454 & ~x84 & ~x108 & ~x112 & ~x162 & ~x198 & ~x200 & ~x203 & ~x226 & ~x275 & ~x280 & ~x419 & ~x677 & ~x753 & ~x780;
assign c7212 =  x390 & ~x11 & ~x33 & ~x116 & ~x139 & ~x167 & ~x170 & ~x176 & ~x191 & ~x192 & ~x193 & ~x194 & ~x531 & ~x556 & ~x557 & ~x558 & ~x587 & ~x610 & ~x641 & ~x670 & ~x698 & ~x738 & ~x783;
assign c7214 =  x403 &  x460 & ~x28 & ~x58 & ~x84 & ~x111 & ~x364 & ~x513 & ~x540 & ~x542 & ~x569 & ~x570 & ~x593 & ~x595 & ~x596 & ~x598 & ~x620 & ~x651 & ~x652 & ~x655 & ~x672 & ~x675 & ~x683 & ~x705 & ~x708 & ~x757 & ~x764 & ~x766;
assign c7216 = ~x57 & ~x76 & ~x77 & ~x472 & ~x498 & ~x501 & ~x512 & ~x518 & ~x519 & ~x527 & ~x529 & ~x575 & ~x589 & ~x590 & ~x644 & ~x674 & ~x689 & ~x710;
assign c7218 = ~x24 & ~x31 & ~x32 & ~x115 & ~x408 & ~x419 & ~x447 & ~x479 & ~x495 & ~x498 & ~x502 & ~x504 & ~x554 & ~x556 & ~x611 & ~x641 & ~x646 & ~x668 & ~x682 & ~x698 & ~x701 & ~x709 & ~x727 & ~x783;
assign c7220 =  x643;
assign c7222 = ~x54 & ~x452 & ~x501 & ~x524 & ~x526 & ~x548 & ~x549 & ~x568 & ~x588 & ~x596 & ~x647 & ~x654 & ~x663 & ~x671 & ~x691 & ~x692 & ~x718 & ~x732 & ~x749;
assign c7224 =  x374 &  x408 & ~x10 & ~x108 & ~x134 & ~x201 & ~x742 & ~x761;
assign c7226 =  x179 &  x428 & ~x36 & ~x106 & ~x442 & ~x466 & ~x555 & ~x713 & ~x749 & ~x773 & ~x774;
assign c7228 =  x520 &  x600 &  x692 & ~x113 & ~x274 & ~x280 & ~x449;
assign c7230 =  x233 & ~x457 & ~x472 & ~x496 & ~x514 & ~x599 & ~x675;
assign c7232 =  x294 &  x296 &  x297 & ~x1 & ~x4 & ~x8 & ~x10 & ~x11 & ~x23 & ~x32 & ~x55 & ~x56 & ~x57 & ~x144 & ~x145 & ~x171 & ~x172 & ~x641 & ~x651 & ~x670 & ~x677 & ~x678 & ~x693 & ~x696 & ~x719 & ~x756 & ~x759 & ~x764;
assign c7234 =  x323 &  x628 & ~x132 & ~x144 & ~x172 & ~x186 & ~x255 & ~x286 & ~x311 & ~x312 & ~x338 & ~x340 & ~x422;
assign c7236 = ~x22 & ~x84 & ~x396 & ~x423 & ~x445 & ~x484 & ~x496 & ~x497 & ~x500 & ~x502 & ~x511 & ~x526 & ~x527 & ~x529 & ~x539 & ~x540 & ~x541 & ~x567 & ~x569 & ~x596 & ~x623 & ~x651 & ~x654 & ~x699 & ~x706 & ~x728;
assign c7238 = ~x18 & ~x25 & ~x26 & ~x27 & ~x30 & ~x55 & ~x57 & ~x85 & ~x447 & ~x468 & ~x471 & ~x472 & ~x484 & ~x485 & ~x496 & ~x497 & ~x498 & ~x499 & ~x500 & ~x501 & ~x502 & ~x503 & ~x511 & ~x512 & ~x524 & ~x540 & ~x542 & ~x552 & ~x553 & ~x568 & ~x569 & ~x582 & ~x587 & ~x588 & ~x598 & ~x623 & ~x645 & ~x655 & ~x672 & ~x673 & ~x674 & ~x681 & ~x682 & ~x708 & ~x728 & ~x737 & ~x751 & ~x758 & ~x759 & ~x763 & ~x771;
assign c7240 =  x278 & ~x1 & ~x51 & ~x57 & ~x80 & ~x500 & ~x521 & ~x522 & ~x524 & ~x526 & ~x553 & ~x592 & ~x618 & ~x621 & ~x675 & ~x692 & ~x693 & ~x700 & ~x757 & ~x761 & ~x762 & ~x776;
assign c7242 =  x521 & ~x3 & ~x26 & ~x35 & ~x59 & ~x85 & ~x139 & ~x141 & ~x197 & ~x224 & ~x336 & ~x437 & ~x438 & ~x503 & ~x669 & ~x687 & ~x702 & ~x704 & ~x731 & ~x754 & ~x757 & ~x779;
assign c7244 = ~x508 & ~x513 & ~x516 & ~x524 & ~x525 & ~x527 & ~x531 & ~x536 & ~x541 & ~x543 & ~x553 & ~x554 & ~x555 & ~x570 & ~x573 & ~x583 & ~x600 & ~x640 & ~x655 & ~x657 & ~x669 & ~x701 & ~x703;
assign c7246 =  x180 &  x295 &  x322 &  x345 & ~x27 & ~x53 & ~x55 & ~x83 & ~x84 & ~x89 & ~x90 & ~x111 & ~x117 & ~x143 & ~x555 & ~x556 & ~x669 & ~x758 & ~x760 & ~x761;
assign c7248 = ~x322 & ~x352 & ~x354 & ~x520 & ~x534 & ~x536 & ~x552 & ~x560 & ~x576 & ~x579 & ~x590 & ~x665 & ~x691 & ~x703 & ~x729;
assign c7250 = ~x57 & ~x408 & ~x475 & ~x501 & ~x526 & ~x553 & ~x562 & ~x571 & ~x600 & ~x614 & ~x638 & ~x648 & ~x653 & ~x655 & ~x681 & ~x683 & ~x695 & ~x702 & ~x706 & ~x710 & ~x711 & ~x722 & ~x738 & ~x739 & ~x749 & ~x754;
assign c7252 =  x388 & ~x1 & ~x56 & ~x112 & ~x134 & ~x169 & ~x170 & ~x171 & ~x172 & ~x197 & ~x224 & ~x309 & ~x613 & ~x622 & ~x649 & ~x651 & ~x667 & ~x670 & ~x676 & ~x679 & ~x695 & ~x698 & ~x707 & ~x725 & ~x761 & ~x779;
assign c7254 =  x238 & ~x40 & ~x57 & ~x111 & ~x530 & ~x552 & ~x554 & ~x555 & ~x557 & ~x567 & ~x582 & ~x585 & ~x607 & ~x637 & ~x678 & ~x698 & ~x699 & ~x700 & ~x701 & ~x732 & ~x761;
assign c7256 =  x346 &  x351 & ~x36 & ~x89 & ~x191 & ~x226 & ~x534 & ~x717;
assign c7258 =  x318 &  x373 & ~x5 & ~x88 & ~x130 & ~x159 & ~x212 & ~x252 & ~x313 & ~x334 & ~x367 & ~x506 & ~x728;
assign c7260 =  x472 & ~x20 & ~x49 & ~x169 & ~x190 & ~x198 & ~x199 & ~x204 & ~x226 & ~x227 & ~x231 & ~x252 & ~x254 & ~x255 & ~x256 & ~x257 & ~x280 & ~x283 & ~x284 & ~x304 & ~x311 & ~x342 & ~x368 & ~x369 & ~x695 & ~x699 & ~x752 & ~x777;
assign c7262 =  x80 &  x262 &  x354 &  x603;
assign c7264 =  x29;
assign c7266 = ~x19 & ~x28 & ~x53 & ~x433 & ~x474 & ~x500 & ~x501 & ~x503 & ~x508 & ~x518 & ~x523 & ~x546 & ~x552 & ~x561 & ~x562 & ~x564 & ~x580 & ~x582 & ~x611 & ~x640 & ~x702 & ~x755 & ~x775;
assign c7268 =  x195;
assign c7270 = ~x0 & ~x25 & ~x34 & ~x113 & ~x408 & ~x409 & ~x474 & ~x488 & ~x495 & ~x497 & ~x526 & ~x534 & ~x608 & ~x609 & ~x629 & ~x668 & ~x758;
assign c7272 = ~x2 & ~x3 & ~x4 & ~x6 & ~x8 & ~x9 & ~x10 & ~x12 & ~x13 & ~x20 & ~x22 & ~x24 & ~x25 & ~x27 & ~x29 & ~x33 & ~x35 & ~x38 & ~x39 & ~x43 & ~x44 & ~x50 & ~x51 & ~x55 & ~x56 & ~x57 & ~x59 & ~x62 & ~x63 & ~x78 & ~x79 & ~x81 & ~x83 & ~x86 & ~x87 & ~x90 & ~x91 & ~x105 & ~x106 & ~x108 & ~x109 & ~x110 & ~x112 & ~x115 & ~x117 & ~x138 & ~x139 & ~x140 & ~x143 & ~x168 & ~x170 & ~x190 & ~x219 & ~x560 & ~x561 & ~x562 & ~x564 & ~x586 & ~x589 & ~x591 & ~x592 & ~x610 & ~x611 & ~x612 & ~x618 & ~x619 & ~x635 & ~x638 & ~x639 & ~x645 & ~x662 & ~x664 & ~x667 & ~x670 & ~x671 & ~x674 & ~x676 & ~x689 & ~x690 & ~x692 & ~x693 & ~x694 & ~x696 & ~x697 & ~x700 & ~x706 & ~x719 & ~x726 & ~x727 & ~x728 & ~x729 & ~x732 & ~x734 & ~x737 & ~x738 & ~x746 & ~x747 & ~x749 & ~x751 & ~x752 & ~x753 & ~x754 & ~x759 & ~x760 & ~x761 & ~x763 & ~x765 & ~x766 & ~x767 & ~x768 & ~x769 & ~x774 & ~x776 & ~x778 & ~x779 & ~x780 & ~x781 & ~x782 & ~x783;
assign c7274 =  x379 & ~x2 & ~x3 & ~x17 & ~x30 & ~x31 & ~x44 & ~x45 & ~x57 & ~x58 & ~x71 & ~x87 & ~x105 & ~x114 & ~x132 & ~x160 & ~x189 & ~x197 & ~x199 & ~x224 & ~x254 & ~x257 & ~x272 & ~x311 & ~x313 & ~x393 & ~x448 & ~x705 & ~x723 & ~x753 & ~x760;
assign c7276 =  x380 &  x486 &  x547 & ~x229 & ~x283 & ~x313 & ~x332;
assign c7278 =  x303 & ~x31 & ~x141 & ~x531 & ~x539 & ~x540 & ~x555 & ~x558 & ~x595 & ~x623 & ~x625 & ~x649 & ~x652 & ~x680 & ~x681 & ~x682 & ~x703 & ~x706 & ~x733 & ~x735 & ~x738 & ~x758 & ~x761 & ~x764;
assign c7280 =  x375 &  x382 & ~x41 & ~x83 & ~x84 & ~x87 & ~x168 & ~x439 & ~x440 & ~x673 & ~x728 & ~x758 & ~x762;
assign c7282 = ~x113 & ~x419 & ~x447 & ~x450 & ~x472 & ~x478 & ~x495 & ~x497 & ~x525 & ~x528 & ~x535 & ~x611 & ~x629 & ~x650 & ~x686 & ~x743 & ~x770 & ~x771;
assign c7284 =  x124 &  x304 & ~x7 & ~x84 & ~x113 & ~x532 & ~x556 & ~x624 & ~x651 & ~x730 & ~x759;
assign c7286 =  x335 & ~x526 & ~x624;
assign c7288 =  x312 & ~x21 & ~x49 & ~x50 & ~x59 & ~x509 & ~x535 & ~x537 & ~x538 & ~x552 & ~x563 & ~x564 & ~x565 & ~x566 & ~x580 & ~x581 & ~x582 & ~x583 & ~x592 & ~x593 & ~x595 & ~x596 & ~x608 & ~x610 & ~x614 & ~x617 & ~x623 & ~x624 & ~x639 & ~x651 & ~x666 & ~x667 & ~x677 & ~x701 & ~x702 & ~x703 & ~x720 & ~x721 & ~x728 & ~x749 & ~x755 & ~x762 & ~x766;
assign c7290 =  x296 &  x346 &  x417 & ~x140 & ~x170 & ~x191 & ~x192 & ~x224 & ~x610 & ~x613 & ~x639 & ~x677 & ~x704 & ~x705 & ~x706;
assign c7292 =  x252;
assign c7294 = ~x5 & ~x10 & ~x27 & ~x36 & ~x39 & ~x41 & ~x48 & ~x50 & ~x61 & ~x62 & ~x65 & ~x133 & ~x135 & ~x144 & ~x148 & ~x175 & ~x193 & ~x199 & ~x228 & ~x255 & ~x280 & ~x307 & ~x536 & ~x588 & ~x613 & ~x645 & ~x674 & ~x676 & ~x678 & ~x699 & ~x718 & ~x734 & ~x763 & ~x764 & ~x783;
assign c7296 =  x319 &  x772;
assign c7298 =  x121 &  x125 &  x235 &  x290 & ~x112 & ~x615 & ~x652 & ~x679;
assign c7300 =  x151 &  x188 & ~x499 & ~x573 & ~x574 & ~x602;
assign c7302 =  x320 &  x348 &  x374 &  x425 & ~x10 & ~x35 & ~x61 & ~x197 & ~x558 & ~x586 & ~x730;
assign c7304 =  x430 & ~x3 & ~x17 & ~x33 & ~x141 & ~x144 & ~x146 & ~x204 & ~x232 & ~x253 & ~x254 & ~x281 & ~x282 & ~x708 & ~x782;
assign c7306 =  x414 & ~x110 & ~x111 & ~x163 & ~x355 & ~x356 & ~x497 & ~x498 & ~x668 & ~x731 & ~x741 & ~x759 & ~x770;
assign c7310 =  x233 & ~x379 & ~x447 & ~x537 & ~x551 & ~x552 & ~x566 & ~x595 & ~x679 & ~x744 & ~x749;
assign c7312 = ~x29 & ~x85 & ~x168 & ~x428 & ~x454 & ~x481 & ~x484 & ~x485 & ~x497 & ~x498 & ~x499 & ~x502 & ~x508 & ~x512 & ~x525 & ~x530 & ~x534 & ~x535 & ~x538 & ~x543 & ~x544 & ~x554 & ~x555 & ~x558 & ~x559 & ~x561 & ~x565 & ~x572 & ~x591 & ~x599 & ~x600 & ~x612 & ~x613 & ~x614 & ~x624 & ~x626 & ~x641 & ~x678 & ~x681 & ~x683 & ~x698 & ~x700 & ~x706 & ~x709 & ~x736 & ~x762 & ~x766;
assign c7314 = ~x25 & ~x70 & ~x71 & ~x79 & ~x103 & ~x132 & ~x147 & ~x175 & ~x218 & ~x256 & ~x258 & ~x285 & ~x310 & ~x364 & ~x368 & ~x586 & ~x670 & ~x737 & ~x771 & ~x772;
assign c7316 =  x356 &  x357 & ~x9 & ~x38 & ~x58 & ~x142 & ~x169 & ~x440 & ~x441 & ~x652 & ~x694 & ~x701 & ~x709 & ~x720 & ~x721 & ~x730 & ~x731 & ~x754 & ~x759 & ~x765 & ~x783;
assign c7318 =  x352 &  x357 &  x399 & ~x649;
assign c7320 =  x155 &  x157 & ~x22 & ~x113 & ~x513 & ~x524 & ~x526 & ~x528 & ~x529 & ~x569 & ~x597 & ~x613 & ~x640 & ~x700;
assign c7322 =  x269 &  x291 & ~x1 & ~x31 & ~x33 & ~x34 & ~x60 & ~x62 & ~x83 & ~x108 & ~x114 & ~x137 & ~x139 & ~x256 & ~x556 & ~x557 & ~x584 & ~x587 & ~x611 & ~x643 & ~x652 & ~x695 & ~x725 & ~x751 & ~x756 & ~x770 & ~x771 & ~x777 & ~x783;
assign c7324 =  x429 &  x486 & ~x1 & ~x5 & ~x7 & ~x9 & ~x23 & ~x27 & ~x54 & ~x58 & ~x105 & ~x167 & ~x596 & ~x640 & ~x652 & ~x707 & ~x725 & ~x756 & ~x761 & ~x774 & ~x777 & ~x778 & ~x780;
assign c7326 =  x139;
assign c7328 =  x265 &  x440 & ~x221 & ~x222 & ~x383 & ~x553 & ~x696;
assign c7330 =  x152 & ~x0 & ~x1 & ~x28 & ~x53 & ~x55 & ~x56 & ~x111 & ~x112 & ~x279 & ~x336 & ~x355 & ~x382 & ~x385 & ~x558 & ~x584 & ~x586 & ~x611 & ~x641 & ~x647 & ~x648 & ~x651 & ~x669 & ~x670 & ~x677 & ~x696 & ~x753 & ~x777 & ~x782;
assign c7332 =  x563 & ~x4 & ~x21 & ~x26 & ~x28 & ~x85 & ~x86 & ~x171 & ~x225 & ~x230 & ~x255 & ~x282 & ~x308 & ~x309 & ~x338 & ~x364 & ~x393 & ~x394 & ~x421 & ~x649 & ~x703 & ~x704 & ~x725 & ~x754 & ~x761 & ~x778 & ~x781;
assign c7334 =  x425 &  x572 & ~x22 & ~x26 & ~x53 & ~x106 & ~x139 & ~x142 & ~x168 & ~x169 & ~x170 & ~x222 & ~x223 & ~x226 & ~x615 & ~x624 & ~x651 & ~x696 & ~x703 & ~x728 & ~x731 & ~x753 & ~x782 & ~x783;
assign c7336 =  x326 & ~x58 & ~x89 & ~x108 & ~x116 & ~x142 & ~x170 & ~x171 & ~x173 & ~x216 & ~x254 & ~x281 & ~x617 & ~x637 & ~x667 & ~x669 & ~x671 & ~x695 & ~x700 & ~x702 & ~x703 & ~x718 & ~x721 & ~x731 & ~x737 & ~x747 & ~x749 & ~x750 & ~x755 & ~x763 & ~x765 & ~x773 & ~x775 & ~x783;
assign c7338 =  x570 &  x627 &  x682 &  x683 &  x710 &  x738 & ~x102 & ~x129 & ~x158 & ~x255;
assign c7340 = ~x3 & ~x5 & ~x33 & ~x86 & ~x87 & ~x93 & ~x102 & ~x134 & ~x148 & ~x172 & ~x195 & ~x197 & ~x199 & ~x226 & ~x247 & ~x480 & ~x510 & ~x582 & ~x615 & ~x637 & ~x665 & ~x703 & ~x725 & ~x736 & ~x753 & ~x767 & ~x768;
assign c7342 =  x379 & ~x1 & ~x2 & ~x6 & ~x20 & ~x30 & ~x35 & ~x36 & ~x51 & ~x79 & ~x87 & ~x88 & ~x89 & ~x108 & ~x109 & ~x110 & ~x131 & ~x135 & ~x141 & ~x169 & ~x197 & ~x198 & ~x255 & ~x257 & ~x282 & ~x313 & ~x339 & ~x340 & ~x586 & ~x613 & ~x669 & ~x697 & ~x726 & ~x727 & ~x743 & ~x756 & ~x757 & ~x781;
assign c7344 =  x97 &  x575 & ~x557;
assign c7346 =  x350 &  x525;
assign c7348 =  x452 & ~x147 & ~x197 & ~x201 & ~x225 & ~x227 & ~x243 & ~x253 & ~x254 & ~x284 & ~x623 & ~x637 & ~x639 & ~x723;
assign c7350 =  x409 &  x576 & ~x105 & ~x143 & ~x170 & ~x256 & ~x310 & ~x339 & ~x340 & ~x367 & ~x422 & ~x763;
assign c7352 = ~x5 & ~x42 & ~x49 & ~x51 & ~x55 & ~x58 & ~x83 & ~x91 & ~x92 & ~x134 & ~x162 & ~x168 & ~x197 & ~x254 & ~x275 & ~x563 & ~x588 & ~x641 & ~x667 & ~x669 & ~x696 & ~x700 & ~x717 & ~x736 & ~x737 & ~x781;
assign c7354 =  x236 & ~x0 & ~x502 & ~x513 & ~x538 & ~x569 & ~x570 & ~x591 & ~x592 & ~x599 & ~x618 & ~x620 & ~x635 & ~x648 & ~x663 & ~x664 & ~x672 & ~x680 & ~x708 & ~x734 & ~x736 & ~x749;
assign c7356 =  x301 & ~x384 & ~x531 & ~x581 & ~x600 & ~x610 & ~x628 & ~x657 & ~x696 & ~x703;
assign c7358 =  x408 & ~x17 & ~x28 & ~x57 & ~x87 & ~x145 & ~x170 & ~x198 & ~x199 & ~x227 & ~x230 & ~x280 & ~x282 & ~x285 & ~x339 & ~x367 & ~x699 & ~x744 & ~x767 & ~x770;
assign c7360 =  x402 & ~x6 & ~x8 & ~x25 & ~x35 & ~x37 & ~x38 & ~x89 & ~x117 & ~x171 & ~x198 & ~x201 & ~x254 & ~x255 & ~x256 & ~x280 & ~x282 & ~x614 & ~x673 & ~x687 & ~x726 & ~x731 & ~x733 & ~x734 & ~x745 & ~x755 & ~x759;
assign c7362 =  x289 & ~x3 & ~x23 & ~x24 & ~x47 & ~x57 & ~x112 & ~x483 & ~x503 & ~x509 & ~x511 & ~x525 & ~x527 & ~x541 & ~x553 & ~x556 & ~x590 & ~x596 & ~x650 & ~x651 & ~x654 & ~x674 & ~x757;
assign c7364 = ~x47 & ~x49 & ~x59 & ~x60 & ~x377 & ~x490 & ~x498 & ~x502 & ~x519 & ~x526 & ~x528 & ~x564 & ~x605 & ~x635 & ~x648 & ~x675 & ~x702 & ~x776;
assign c7366 =  x168;
assign c7368 =  x627 &  x710 & ~x26 & ~x27 & ~x31 & ~x85 & ~x87 & ~x103 & ~x112 & ~x113 & ~x114 & ~x157 & ~x169 & ~x170 & ~x198 & ~x366 & ~x421 & ~x446 & ~x448 & ~x641 & ~x669 & ~x761;
assign c7370 =  x461 &  x547 &  x633 & ~x58 & ~x111 & ~x168 & ~x171 & ~x225 & ~x580 & ~x764;
assign c7372 =  x371 &  x486 & ~x0 & ~x7 & ~x28 & ~x29 & ~x31 & ~x60 & ~x78 & ~x81 & ~x85 & ~x107 & ~x111 & ~x112 & ~x139 & ~x511 & ~x595 & ~x672 & ~x675 & ~x694 & ~x697 & ~x728 & ~x729 & ~x731 & ~x752 & ~x755;
assign c7374 = ~x1 & ~x2 & ~x53 & ~x54 & ~x82 & ~x85 & ~x112 & ~x141 & ~x458 & ~x481 & ~x502 & ~x506 & ~x526 & ~x530 & ~x543 & ~x544 & ~x554 & ~x556 & ~x557 & ~x559 & ~x560 & ~x565 & ~x572 & ~x587 & ~x592 & ~x599 & ~x614 & ~x629 & ~x644 & ~x647 & ~x648 & ~x655 & ~x670 & ~x678 & ~x684 & ~x698 & ~x701 & ~x704 & ~x706 & ~x710 & ~x711 & ~x754 & ~x756 & ~x757 & ~x761;
assign c7376 =  x548 & ~x24 & ~x29 & ~x35 & ~x111 & ~x133 & ~x160 & ~x169 & ~x173 & ~x194 & ~x222 & ~x251 & ~x717;
assign c7378 =  x196;
assign c7380 = ~x25 & ~x28 & ~x29 & ~x86 & ~x168 & ~x446 & ~x475 & ~x476 & ~x496 & ~x498 & ~x501 & ~x510 & ~x529 & ~x538 & ~x543 & ~x558 & ~x569 & ~x571 & ~x572 & ~x585 & ~x586 & ~x589 & ~x596 & ~x599 & ~x614 & ~x626 & ~x628 & ~x642 & ~x646 & ~x650 & ~x656 & ~x657 & ~x671 & ~x674 & ~x685 & ~x729 & ~x730 & ~x767 & ~x781;
assign c7382 =  x179 &  x211 & ~x1 & ~x25 & ~x475 & ~x530 & ~x538 & ~x566 & ~x612 & ~x623 & ~x624 & ~x649 & ~x651 & ~x669 & ~x726 & ~x732 & ~x754 & ~x778 & ~x780;
assign c7384 =  x351 &  x517 & ~x1 & ~x70 & ~x88 & ~x141 & ~x170 & ~x226 & ~x253 & ~x393 & ~x615 & ~x668 & ~x673 & ~x752 & ~x772;
assign c7386 = ~x19 & ~x23 & ~x26 & ~x28 & ~x36 & ~x50 & ~x56 & ~x61 & ~x62 & ~x63 & ~x73 & ~x102 & ~x105 & ~x108 & ~x109 & ~x111 & ~x113 & ~x117 & ~x140 & ~x142 & ~x146 & ~x197 & ~x224 & ~x281 & ~x530 & ~x531 & ~x551 & ~x556 & ~x565 & ~x578 & ~x579 & ~x580 & ~x588 & ~x611 & ~x619 & ~x620 & ~x637 & ~x644 & ~x646 & ~x647 & ~x670 & ~x702 & ~x715 & ~x727 & ~x759 & ~x767 & ~x772 & ~x779;
assign c7388 =  x305 & ~x22 & ~x23 & ~x30 & ~x78 & ~x79 & ~x85 & ~x109 & ~x110 & ~x141 & ~x224 & ~x420 & ~x448 & ~x474 & ~x475 & ~x500 & ~x501 & ~x502 & ~x503 & ~x524 & ~x525 & ~x527 & ~x554 & ~x557 & ~x558 & ~x568 & ~x582 & ~x610 & ~x612 & ~x622 & ~x623 & ~x624 & ~x639 & ~x650 & ~x651 & ~x697 & ~x702 & ~x728 & ~x749 & ~x759 & ~x760 & ~x761 & ~x778 & ~x780;
assign c7390 =  x155 &  x220 & ~x501 & ~x520 & ~x527;
assign c7392 =  x16 &  x291 & ~x584 & ~x623;
assign c7394 =  x380 &  x456 &  x457 &  x484 & ~x30 & ~x32 & ~x61 & ~x65 & ~x174 & ~x198;
assign c7396 = ~x8 & ~x9 & ~x19 & ~x20 & ~x24 & ~x28 & ~x30 & ~x32 & ~x35 & ~x36 & ~x56 & ~x59 & ~x60 & ~x63 & ~x80 & ~x84 & ~x89 & ~x90 & ~x106 & ~x109 & ~x111 & ~x113 & ~x140 & ~x141 & ~x142 & ~x170 & ~x197 & ~x198 & ~x225 & ~x561 & ~x630 & ~x632 & ~x672 & ~x674 & ~x687 & ~x701 & ~x719 & ~x725 & ~x728 & ~x732 & ~x734 & ~x742 & ~x743 & ~x745 & ~x748 & ~x749 & ~x750 & ~x753 & ~x756 & ~x757 & ~x759 & ~x760 & ~x761 & ~x762 & ~x772 & ~x775 & ~x776 & ~x777 & ~x778 & ~x783;
assign c7398 =  x296 &  x321 &  x348 &  x373 & ~x7 & ~x8 & ~x10 & ~x84 & ~x110 & ~x136 & ~x144 & ~x162 & ~x191 & ~x194 & ~x195 & ~x197 & ~x224 & ~x559 & ~x586 & ~x614 & ~x641 & ~x671 & ~x696 & ~x704 & ~x723 & ~x728 & ~x729 & ~x734 & ~x735 & ~x751 & ~x752 & ~x753 & ~x755 & ~x783;
assign c7400 =  x418 & ~x35 & ~x53 & ~x85 & ~x109 & ~x221 & ~x222 & ~x336 & ~x414 & ~x586 & ~x637 & ~x700 & ~x732 & ~x766;
assign c7402 = ~x54 & ~x55 & ~x57 & ~x81 & ~x82 & ~x141 & ~x451 & ~x474 & ~x486 & ~x498 & ~x500 & ~x527 & ~x528 & ~x545 & ~x565 & ~x566 & ~x573 & ~x588 & ~x594 & ~x602 & ~x611 & ~x613 & ~x622 & ~x628 & ~x641 & ~x643 & ~x656 & ~x657 & ~x676 & ~x697 & ~x705 & ~x724 & ~x739 & ~x751 & ~x782;
assign c7404 =  x278 & ~x20 & ~x22 & ~x28 & ~x29 & ~x31 & ~x84 & ~x112 & ~x113 & ~x447 & ~x496 & ~x499 & ~x500 & ~x503 & ~x525 & ~x527 & ~x528 & ~x567 & ~x595 & ~x596 & ~x622 & ~x623 & ~x625 & ~x653 & ~x680 & ~x728 & ~x762;
assign c7406 =  x334 & ~x51 & ~x81 & ~x106 & ~x329 & ~x500 & ~x501 & ~x502 & ~x525 & ~x526 & ~x564 & ~x592 & ~x594 & ~x611 & ~x650 & ~x672 & ~x747 & ~x757 & ~x762 & ~x777;
assign c7408 = ~x25 & ~x31 & ~x51 & ~x58 & ~x83 & ~x113 & ~x168 & ~x195 & ~x481 & ~x482 & ~x502 & ~x508 & ~x509 & ~x530 & ~x532 & ~x568 & ~x582 & ~x583 & ~x594 & ~x596 & ~x614 & ~x626 & ~x629 & ~x639 & ~x647 & ~x653 & ~x654 & ~x676 & ~x679 & ~x708 & ~x710 & ~x718 & ~x722 & ~x727 & ~x731 & ~x734 & ~x758 & ~x780;
assign c7410 =  x352 &  x375 & ~x13 & ~x117 & ~x145 & ~x168 & ~x170 & ~x192 & ~x200 & ~x227 & ~x256 & ~x257 & ~x642 & ~x723 & ~x766;
assign c7412 =  x365;
assign c7414 =  x27;
assign c7416 =  x400 &  x514 &  x521 & ~x198 & ~x228;
assign c7418 =  x571 &  x600 & ~x0 & ~x18 & ~x26 & ~x33 & ~x84 & ~x129 & ~x131 & ~x199 & ~x253 & ~x259 & ~x280 & ~x284 & ~x309 & ~x314 & ~x367 & ~x614 & ~x669 & ~x670 & ~x706 & ~x775 & ~x776 & ~x781;
assign c7420 =  x518 & ~x19 & ~x113 & ~x131 & ~x159 & ~x197 & ~x201 & ~x204 & ~x229 & ~x255 & ~x283 & ~x312 & ~x338 & ~x339 & ~x365 & ~x394 & ~x421 & ~x423 & ~x622 & ~x724 & ~x772 & ~x773;
assign c7422 = ~x5 & ~x20 & ~x29 & ~x32 & ~x56 & ~x59 & ~x85 & ~x448 & ~x489 & ~x499 & ~x500 & ~x501 & ~x519 & ~x523 & ~x525 & ~x527 & ~x528 & ~x530 & ~x534 & ~x552 & ~x554 & ~x555 & ~x557 & ~x580 & ~x582 & ~x585 & ~x616 & ~x633 & ~x642 & ~x644 & ~x646 & ~x669 & ~x672 & ~x674 & ~x700 & ~x703 & ~x750 & ~x757 & ~x780 & ~x782 & ~x783;
assign c7424 = ~x113 & ~x391 & ~x448 & ~x462 & ~x498 & ~x505 & ~x527 & ~x534 & ~x551 & ~x576 & ~x589 & ~x590 & ~x597 & ~x645 & ~x661 & ~x729 & ~x746;
assign c7426 = ~x0 & ~x2 & ~x3 & ~x13 & ~x14 & ~x16 & ~x18 & ~x24 & ~x26 & ~x28 & ~x35 & ~x39 & ~x57 & ~x65 & ~x68 & ~x71 & ~x80 & ~x87 & ~x93 & ~x94 & ~x98 & ~x115 & ~x117 & ~x150 & ~x175 & ~x177 & ~x189 & ~x190 & ~x196 & ~x198 & ~x224 & ~x230 & ~x253 & ~x336 & ~x692 & ~x693 & ~x706 & ~x708 & ~x720 & ~x722 & ~x724 & ~x734 & ~x764 & ~x771 & ~x782;
assign c7428 =  x352 &  x509 &  x564 & ~x0 & ~x102 & ~x169 & ~x201 & ~x228 & ~x312 & ~x341 & ~x761;
assign c7430 =  x358 & ~x301 & ~x442 & ~x466 & ~x705 & ~x759;
assign c7432 = ~x418 & ~x445 & ~x447 & ~x465 & ~x466 & ~x467 & ~x469 & ~x472 & ~x474 & ~x494 & ~x496 & ~x499 & ~x500 & ~x522 & ~x542 & ~x552 & ~x555 & ~x556 & ~x558 & ~x580 & ~x599 & ~x626 & ~x653 & ~x654 & ~x655 & ~x681 & ~x682 & ~x765;
assign c7434 =  x17 &  x747;
assign c7436 =  x302 & ~x416 & ~x440 & ~x505 & ~x514 & ~x534 & ~x542 & ~x626 & ~x654;
assign c7438 = ~x0 & ~x2 & ~x10 & ~x21 & ~x28 & ~x30 & ~x51 & ~x58 & ~x77 & ~x82 & ~x83 & ~x86 & ~x107 & ~x108 & ~x112 & ~x224 & ~x279 & ~x530 & ~x531 & ~x558 & ~x559 & ~x560 & ~x579 & ~x580 & ~x581 & ~x584 & ~x585 & ~x586 & ~x594 & ~x595 & ~x596 & ~x597 & ~x607 & ~x609 & ~x610 & ~x612 & ~x613 & ~x614 & ~x622 & ~x623 & ~x624 & ~x625 & ~x636 & ~x637 & ~x638 & ~x641 & ~x642 & ~x644 & ~x650 & ~x651 & ~x652 & ~x653 & ~x654 & ~x665 & ~x666 & ~x667 & ~x668 & ~x672 & ~x673 & ~x674 & ~x679 & ~x680 & ~x681 & ~x682 & ~x683 & ~x693 & ~x696 & ~x697 & ~x700 & ~x702 & ~x706 & ~x708 & ~x709 & ~x710 & ~x722 & ~x723 & ~x724 & ~x726 & ~x727 & ~x728 & ~x729 & ~x732 & ~x733 & ~x736 & ~x740 & ~x750 & ~x751 & ~x752 & ~x756 & ~x759 & ~x761 & ~x763 & ~x765 & ~x766 & ~x777 & ~x780 & ~x781;
assign c7440 =  x490 & ~x27 & ~x58 & ~x83 & ~x102 & ~x111 & ~x156 & ~x158 & ~x168 & ~x185 & ~x200 & ~x222 & ~x225 & ~x226 & ~x227 & ~x255 & ~x283 & ~x284 & ~x309 & ~x339 & ~x587 & ~x613 & ~x614 & ~x616 & ~x724 & ~x752 & ~x775 & ~x780;
assign c7442 =  x184 &  x235 &  x262 & ~x624;
assign c7444 =  x123 &  x249 & ~x54 & ~x56 & ~x82 & ~x495 & ~x496 & ~x503 & ~x527 & ~x529 & ~x532 & ~x538 & ~x552 & ~x555 & ~x564 & ~x583 & ~x594 & ~x615 & ~x622 & ~x645 & ~x670 & ~x672 & ~x698 & ~x706 & ~x734 & ~x757;
assign c7446 = ~x0 & ~x2 & ~x23 & ~x49 & ~x79 & ~x81 & ~x103 & ~x129 & ~x133 & ~x134 & ~x141 & ~x169 & ~x170 & ~x171 & ~x199 & ~x228 & ~x254 & ~x261 & ~x282 & ~x284 & ~x310 & ~x337 & ~x338 & ~x342 & ~x614 & ~x670 & ~x708 & ~x724 & ~x727 & ~x735 & ~x753 & ~x771 & ~x779 & ~x780 & ~x783;
assign c7448 = ~x2 & ~x5 & ~x7 & ~x10 & ~x18 & ~x23 & ~x24 & ~x25 & ~x27 & ~x28 & ~x35 & ~x38 & ~x48 & ~x49 & ~x50 & ~x55 & ~x58 & ~x59 & ~x60 & ~x62 & ~x64 & ~x81 & ~x86 & ~x92 & ~x108 & ~x111 & ~x112 & ~x133 & ~x137 & ~x163 & ~x164 & ~x166 & ~x167 & ~x169 & ~x190 & ~x195 & ~x196 & ~x197 & ~x221 & ~x224 & ~x250 & ~x251 & ~x532 & ~x537 & ~x538 & ~x559 & ~x562 & ~x563 & ~x565 & ~x591 & ~x613 & ~x615 & ~x619 & ~x620 & ~x642 & ~x644 & ~x645 & ~x666 & ~x673 & ~x678 & ~x694 & ~x696 & ~x697 & ~x698 & ~x700 & ~x701 & ~x703 & ~x715 & ~x726 & ~x728 & ~x730 & ~x732 & ~x733 & ~x735 & ~x738 & ~x746 & ~x749 & ~x753 & ~x754 & ~x755 & ~x756 & ~x757 & ~x758 & ~x759 & ~x760 & ~x761 & ~x763 & ~x764 & ~x765 & ~x767 & ~x771 & ~x772 & ~x778 & ~x783;
assign c7450 = ~x0 & ~x21 & ~x26 & ~x29 & ~x57 & ~x68 & ~x80 & ~x115 & ~x120 & ~x133 & ~x136 & ~x137 & ~x175 & ~x188 & ~x189 & ~x230 & ~x257 & ~x475 & ~x502 & ~x530 & ~x531 & ~x555 & ~x586 & ~x669 & ~x677 & ~x719 & ~x720 & ~x756 & ~x760 & ~x768;
assign c7452 =  x238 &  x276 & ~x576 & ~x578 & ~x604 & ~x607 & ~x611 & ~x637 & ~x691 & ~x693 & ~x720 & ~x724 & ~x749 & ~x783;
assign c7454 = ~x24 & ~x54 & ~x55 & ~x89 & ~x435 & ~x474 & ~x475 & ~x492 & ~x493 & ~x498 & ~x499 & ~x531 & ~x553 & ~x579 & ~x599 & ~x617 & ~x618 & ~x634 & ~x637 & ~x646 & ~x665 & ~x668 & ~x694 & ~x696 & ~x726 & ~x727 & ~x748;
assign c7456 =  x520 &  x521 & ~x25 & ~x29 & ~x33 & ~x36 & ~x57 & ~x59 & ~x66 & ~x90 & ~x112 & ~x117 & ~x139 & ~x141 & ~x142 & ~x143 & ~x144 & ~x145 & ~x172 & ~x197 & ~x224 & ~x226 & ~x228 & ~x229 & ~x309 & ~x314 & ~x726 & ~x779;
assign c7458 = ~x4 & ~x78 & ~x79 & ~x85 & ~x86 & ~x168 & ~x446 & ~x473 & ~x477 & ~x478 & ~x495 & ~x496 & ~x498 & ~x500 & ~x556 & ~x601 & ~x629 & ~x674 & ~x688 & ~x702 & ~x743 & ~x762 & ~x773 & ~x774;
assign c7460 = ~x29 & ~x83 & ~x390 & ~x411 & ~x415 & ~x416 & ~x417 & ~x419 & ~x443 & ~x470 & ~x501 & ~x571 & ~x574 & ~x580 & ~x615 & ~x616 & ~x634 & ~x674 & ~x683 & ~x739;
assign c7462 =  x374 & ~x26 & ~x28 & ~x54 & ~x110 & ~x540 & ~x595 & ~x619 & ~x624 & ~x646 & ~x648 & ~x672 & ~x677 & ~x681 & ~x695 & ~x696 & ~x700 & ~x703 & ~x704 & ~x707 & ~x708 & ~x730 & ~x753 & ~x764 & ~x774;
assign c7464 = ~x25 & ~x28 & ~x55 & ~x58 & ~x445 & ~x446 & ~x467 & ~x468 & ~x469 & ~x480 & ~x496 & ~x498 & ~x505 & ~x618 & ~x629 & ~x643 & ~x676 & ~x703 & ~x714 & ~x744 & ~x783;
assign c7466 =  x25;
assign c7468 =  x601 &  x629 &  x716 & ~x31 & ~x33 & ~x57 & ~x85 & ~x188 & ~x218 & ~x307 & ~x614 & ~x651;
assign c7470 =  x408 &  x455 &  x537 &  x601 & ~x132 & ~x228 & ~x254 & ~x395;
assign c7472 =  x213 &  x249 & ~x499 & ~x524 & ~x623;
assign c7474 =  x45 &  x318 &  x456;
assign c7476 =  x122 &  x316 &  x342 & ~x86 & ~x113 & ~x539 & ~x550 & ~x551 & ~x552 & ~x594 & ~x623 & ~x645 & ~x650 & ~x675 & ~x702 & ~x729;
assign c7478 =  x280 &  x323;
assign c7480 =  x573 &  x691 & ~x102 & ~x142 & ~x218 & ~x245 & ~x257;
assign c7482 = ~x25 & ~x59 & ~x140 & ~x323 & ~x532 & ~x537 & ~x539 & ~x549 & ~x555 & ~x561 & ~x577 & ~x579 & ~x589 & ~x605 & ~x618 & ~x625 & ~x636 & ~x647 & ~x663 & ~x679 & ~x682 & ~x690 & ~x708 & ~x728 & ~x737 & ~x747 & ~x757 & ~x775;
assign c7484 = ~x0 & ~x4 & ~x20 & ~x24 & ~x27 & ~x28 & ~x33 & ~x51 & ~x53 & ~x55 & ~x56 & ~x57 & ~x86 & ~x112 & ~x113 & ~x509 & ~x530 & ~x548 & ~x556 & ~x557 & ~x560 & ~x561 & ~x564 & ~x577 & ~x583 & ~x585 & ~x591 & ~x592 & ~x593 & ~x605 & ~x606 & ~x607 & ~x614 & ~x618 & ~x621 & ~x635 & ~x636 & ~x644 & ~x646 & ~x649 & ~x650 & ~x669 & ~x674 & ~x675 & ~x676 & ~x691 & ~x693 & ~x698 & ~x699 & ~x702 & ~x704 & ~x705 & ~x719 & ~x720 & ~x721 & ~x722 & ~x728 & ~x729 & ~x731 & ~x746 & ~x747 & ~x750 & ~x756 & ~x757 & ~x759 & ~x760 & ~x777 & ~x778;
assign c7486 =  x307;
assign c7488 = ~x76 & ~x77 & ~x453 & ~x454 & ~x504 & ~x505 & ~x513 & ~x553 & ~x565 & ~x570 & ~x590 & ~x599 & ~x621 & ~x624 & ~x635 & ~x662 & ~x678 & ~x683 & ~x758 & ~x761;
assign c7490 =  x297 & ~x1 & ~x2 & ~x11 & ~x22 & ~x36 & ~x47 & ~x48 & ~x53 & ~x55 & ~x63 & ~x64 & ~x78 & ~x79 & ~x84 & ~x89 & ~x104 & ~x106 & ~x113 & ~x131 & ~x132 & ~x135 & ~x138 & ~x140 & ~x141 & ~x144 & ~x145 & ~x166 & ~x169 & ~x170 & ~x172 & ~x173 & ~x195 & ~x197 & ~x198 & ~x201 & ~x224 & ~x225 & ~x227 & ~x254 & ~x255 & ~x280 & ~x310 & ~x311 & ~x337 & ~x393 & ~x502 & ~x531 & ~x555 & ~x559 & ~x587 & ~x641 & ~x642 & ~x643 & ~x644 & ~x670 & ~x775 & ~x776;
assign c7492 =  x425 &  x547 & ~x84 & ~x88 & ~x113 & ~x133 & ~x146 & ~x161 & ~x594 & ~x668 & ~x678 & ~x697 & ~x698 & ~x758;
assign c7494 =  x360 & ~x141 & ~x252 & ~x419 & ~x444 & ~x469 & ~x496 & ~x623 & ~x652 & ~x677 & ~x763 & ~x770 & ~x778;
assign c7496 =  x209 &  x286 &  x287 & ~x16 & ~x42 & ~x48 & ~x85 & ~x142 & ~x419 & ~x470 & ~x495 & ~x538 & ~x762;
assign c7498 =  x417 &  x418 & ~x1 & ~x7 & ~x23 & ~x27 & ~x28 & ~x31 & ~x82 & ~x140 & ~x162 & ~x169 & ~x170 & ~x192 & ~x197 & ~x198 & ~x218 & ~x219 & ~x246 & ~x248 & ~x250 & ~x251 & ~x252 & ~x587 & ~x613 & ~x637 & ~x669 & ~x697 & ~x704 & ~x725 & ~x726 & ~x731 & ~x733 & ~x734 & ~x760 & ~x764 & ~x766 & ~x768 & ~x776 & ~x780;
assign c71 = ~x34 & ~x547 & ~x577 & ~x656 & ~x658 & ~x680 & ~x764;
assign c73 = ~x24 & ~x234 & ~x364 & ~x606 & ~x632 & ~x633 & ~x659 & ~x681 & ~x682 & ~x686 & ~x708 & ~x709 & ~x736 & ~x740 & ~x748 & ~x764;
assign c75 = ~x81 & ~x108 & ~x133 & ~x161 & ~x280 & ~x284 & ~x285 & ~x307 & ~x313 & ~x334 & ~x335 & ~x341 & ~x365 & ~x369 & ~x385 & ~x416 & ~x444 & ~x480 & ~x503 & ~x538 & ~x553 & ~x567 & ~x592 & ~x593 & ~x652;
assign c77 = ~x29 & ~x69 & ~x126 & ~x151 & ~x377 & ~x378 & ~x405 & ~x433;
assign c79 = ~x28 & ~x84 & ~x110 & ~x140 & ~x162 & ~x222 & ~x248 & ~x249 & ~x304 & ~x305 & ~x308 & ~x392 & ~x401 & ~x562 & ~x664 & ~x698;
assign c711 = ~x203 & ~x409 & ~x463 & ~x464 & ~x491 & ~x545;
assign c713 =  x183 & ~x110 & ~x136 & ~x141 & ~x161 & ~x194 & ~x219 & ~x248 & ~x280 & ~x337 & ~x361 & ~x362 & ~x391;
assign c715 =  x98 & ~x188 & ~x248 & ~x273 & ~x324 & ~x449 & ~x561;
assign c717 = ~x174 & ~x438 & ~x466 & ~x491 & ~x493 & ~x494 & ~x518 & ~x521 & ~x572 & ~x573 & ~x760;
assign c719 = ~x1 & ~x3 & ~x6 & ~x31 & ~x56 & ~x86 & ~x135 & ~x193 & ~x224 & ~x251 & ~x307 & ~x547 & ~x548 & ~x549 & ~x576 & ~x602 & ~x603 & ~x630 & ~x656 & ~x657 & ~x727 & ~x778;
assign c721 =  x675 & ~x168 & ~x391 & ~x419 & ~x627 & ~x684;
assign c723 = ~x8 & ~x164 & ~x166 & ~x191 & ~x280 & ~x282 & ~x336 & ~x339 & ~x367 & ~x395 & ~x451 & ~x470 & ~x473 & ~x507 & ~x566 & ~x608 & ~x620 & ~x680 & ~x704 & ~x761 & ~x780;
assign c725 =  x622 &  x623 & ~x26 & ~x27 & ~x55 & ~x126 & ~x154 & ~x783;
assign c727 =  x360 & ~x184 & ~x185 & ~x211 & ~x239 & ~x327 & ~x758;
assign c729 =  x43 & ~x79 & ~x190 & ~x221 & ~x251 & ~x363 & ~x391 & ~x510;
assign c731 =  x565 &  x566 &  x593 &  x594 & ~x0 & ~x99 & ~x308 & ~x364 & ~x766 & ~x770;
assign c733 =  x181 &  x741 & ~x55 & ~x82 & ~x83 & ~x190 & ~x222 & ~x305 & ~x501 & ~x702;
assign c735 =  x285 &  x549 & ~x3 & ~x4 & ~x81 & ~x319 & ~x346 & ~x448 & ~x756;
assign c737 =  x604 &  x631 & ~x21 & ~x23 & ~x24 & ~x50 & ~x80 & ~x110 & ~x111 & ~x113 & ~x164 & ~x365 & ~x418 & ~x478 & ~x502 & ~x531 & ~x556 & ~x588 & ~x589 & ~x591 & ~x592 & ~x646 & ~x705 & ~x732 & ~x758 & ~x783;
assign c739 = ~x1 & ~x14 & ~x20 & ~x26 & ~x27 & ~x43 & ~x45 & ~x46 & ~x47 & ~x49 & ~x52 & ~x53 & ~x56 & ~x81 & ~x82 & ~x106 & ~x110 & ~x111 & ~x112 & ~x138 & ~x167 & ~x170 & ~x192 & ~x194 & ~x225 & ~x249 & ~x250 & ~x252 & ~x253 & ~x281 & ~x306 & ~x308 & ~x334 & ~x336 & ~x363 & ~x557 & ~x615 & ~x627 & ~x755 & ~x780;
assign c741 =  x527 &  x555 &  x582 &  x610 & ~x0 & ~x25 & ~x27 & ~x28 & ~x53 & ~x57 & ~x81 & ~x111 & ~x138 & ~x766;
assign c743 =  x556 & ~x0 & ~x27 & ~x28 & ~x574 & ~x601;
assign c745 =  x509 & ~x15 & ~x18 & ~x43 & ~x45 & ~x268 & ~x296 & ~x323 & ~x364 & ~x420 & ~x700 & ~x718 & ~x780 & ~x781;
assign c747 =  x415 &  x443 & ~x0 & ~x54 & ~x409 & ~x410 & ~x438 & ~x465 & ~x466 & ~x493 & ~x699 & ~x756 & ~x783;
assign c749 =  x269 & ~x51 & ~x54 & ~x57 & ~x112 & ~x138 & ~x252 & ~x308 & ~x373 & ~x425 & ~x476 & ~x504 & ~x672 & ~x757;
assign c751 =  x257 &  x538 & ~x224 & ~x420 & ~x690 & ~x691 & ~x718 & ~x719 & ~x746 & ~x747 & ~x762 & ~x772 & ~x775;
assign c753 =  x418 & ~x353 & ~x380 & ~x439 & ~x466 & ~x494 & ~x495;
assign c755 = ~x28 & ~x46 & ~x71 & ~x77 & ~x86 & ~x98 & ~x99 & ~x212 & ~x240 & ~x266;
assign c757 =  x360 &  x416 & ~x2 & ~x4 & ~x115 & ~x365 & ~x412 & ~x774 & ~x776;
assign c759 =  x575 &  x627 & ~x24 & ~x83 & ~x449 & ~x696 & ~x721 & ~x722 & ~x738 & ~x767 & ~x783;
assign c761 = ~x1 & ~x168 & ~x280 & ~x304 & ~x311 & ~x334 & ~x397 & ~x445 & ~x511 & ~x563 & ~x750;
assign c763 =  x556 & ~x322;
assign c765 = ~x19 & ~x71 & ~x127 & ~x209 & ~x237 & ~x417 & ~x445 & ~x473 & ~x474 & ~x475 & ~x503 & ~x558 & ~x560 & ~x561 & ~x643 & ~x729;
assign c767 =  x155 & ~x244 & ~x273 & ~x279 & ~x302 & ~x303 & ~x330 & ~x334 & ~x391 & ~x416 & ~x472 & ~x474 & ~x499 & ~x500 & ~x560;
assign c769 = ~x37 & ~x105 & ~x135 & ~x139 & ~x164 & ~x167 & ~x168 & ~x192 & ~x194 & ~x195 & ~x251 & ~x308 & ~x437 & ~x465 & ~x494 & ~x522 & ~x551 & ~x552;
assign c771 =  x257 & ~x2 & ~x57 & ~x122 & ~x123 & ~x150 & ~x233;
assign c773 = ~x189 & ~x216 & ~x217 & ~x218 & ~x245 & ~x247 & ~x273 & ~x275 & ~x301 & ~x302 & ~x336 & ~x351 & ~x502 & ~x531 & ~x559 & ~x562;
assign c775 =  x668 & ~x24 & ~x26 & ~x307 & ~x363;
assign c777 = ~x1 & ~x26 & ~x207 & ~x233 & ~x376 & ~x430 & ~x431 & ~x512 & ~x513 & ~x531 & ~x761 & ~x778;
assign c779 = ~x56 & ~x381 & ~x435 & ~x462 & ~x489 & ~x653;
assign c781 =  x717 & ~x104 & ~x137 & ~x139 & ~x162 & ~x168 & ~x253 & ~x360 & ~x389 & ~x416 & ~x424 & ~x444 & ~x446 & ~x472 & ~x477 & ~x526 & ~x534 & ~x555 & ~x558 & ~x610 & ~x614 & ~x729;
assign c783 = ~x0 & ~x35 & ~x55 & ~x63 & ~x115 & ~x144 & ~x173 & ~x227 & ~x249 & ~x252 & ~x279 & ~x336 & ~x352 & ~x353 & ~x380 & ~x381 & ~x408 & ~x445 & ~x504;
assign c785 =  x494 &  x575 &  x602 &  x603 & ~x0 & ~x2 & ~x20 & ~x28 & ~x615 & ~x694 & ~x719 & ~x721 & ~x722 & ~x747 & ~x756 & ~x777;
assign c787 = ~x23 & ~x36 & ~x48 & ~x80 & ~x86 & ~x116 & ~x194 & ~x254 & ~x284 & ~x412 & ~x492 & ~x493 & ~x495 & ~x520 & ~x701 & ~x704;
assign c789 = ~x26 & ~x28 & ~x54 & ~x140 & ~x292 & ~x293 & ~x320 & ~x344 & ~x373 & ~x399 & ~x400 & ~x455;
assign c791 =  x496 &  x524 & ~x1 & ~x55 & ~x83 & ~x84 & ~x111 & ~x168 & ~x224 & ~x308 & ~x363 & ~x391 & ~x420 & ~x446 & ~x474 & ~x475 & ~x503 & ~x560 & ~x588 & ~x590 & ~x671 & ~x701 & ~x728 & ~x730 & ~x756 & ~x759;
assign c793 =  x549 &  x576 & ~x15 & ~x26 & ~x27 & ~x111 & ~x422 & ~x555 & ~x695 & ~x722 & ~x750 & ~x758 & ~x778;
assign c795 =  x539 & ~x0 & ~x10 & ~x71 & ~x126 & ~x336 & ~x364 & ~x421 & ~x766 & ~x767 & ~x776;
assign c797 =  x147 & ~x1 & ~x17 & ~x19 & ~x43 & ~x47 & ~x73 & ~x97 & ~x153 & ~x211 & ~x699 & ~x700 & ~x726 & ~x727;
assign c799 = ~x138 & ~x205 & ~x224 & ~x275 & ~x329 & ~x332 & ~x333 & ~x334 & ~x335 & ~x360 & ~x472 & ~x525 & ~x582 & ~x585;
assign c7101 =  x313 & ~x3 & ~x81 & ~x83 & ~x110 & ~x346 & ~x373 & ~x374 & ~x427 & ~x428 & ~x643 & ~x733 & ~x760;
assign c7103 = ~x8 & ~x82 & ~x115 & ~x117 & ~x133 & ~x134 & ~x137 & ~x160 & ~x188 & ~x189 & ~x217 & ~x425 & ~x445 & ~x473 & ~x481 & ~x530 & ~x538;
assign c7105 = ~x162 & ~x188 & ~x190 & ~x193 & ~x219 & ~x225 & ~x227 & ~x246 & ~x253 & ~x274 & ~x361 & ~x389 & ~x420 & ~x508 & ~x511 & ~x534 & ~x538 & ~x539 & ~x592 & ~x670 & ~x726;
assign c7107 =  x568 & ~x1 & ~x3 & ~x4 & ~x26 & ~x51 & ~x53 & ~x54 & ~x58 & ~x252 & ~x336 & ~x455 & ~x482 & ~x504 & ~x588 & ~x671 & ~x699 & ~x700 & ~x761;
assign c7109 = ~x54 & ~x290 & ~x291 & ~x345 & ~x444 & ~x448 & ~x501 & ~x666 & ~x717;
assign c7111 =  x509 & ~x5 & ~x28 & ~x56 & ~x112 & ~x113 & ~x141 & ~x193 & ~x194 & ~x222 & ~x223 & ~x327 & ~x355 & ~x382 & ~x383 & ~x410 & ~x411 & ~x420 & ~x467 & ~x587 & ~x747;
assign c7113 = ~x28 & ~x108 & ~x137 & ~x138 & ~x140 & ~x141 & ~x168 & ~x170 & ~x194 & ~x195 & ~x246 & ~x275 & ~x276 & ~x281 & ~x308 & ~x331 & ~x333 & ~x337 & ~x341 & ~x357 & ~x358 & ~x360 & ~x362 & ~x386 & ~x387 & ~x391 & ~x415 & ~x416 & ~x424 & ~x470 & ~x471 & ~x499 & ~x555 & ~x583 & ~x584 & ~x642 & ~x645 & ~x669 & ~x728 & ~x730;
assign c7115 = ~x24 & ~x27 & ~x109 & ~x139 & ~x147 & ~x164 & ~x194 & ~x462 & ~x489 & ~x573 & ~x629 & ~x780;
assign c7117 =  x548 &  x629 & ~x17 & ~x22 & ~x110 & ~x448 & ~x557 & ~x559 & ~x609 & ~x638 & ~x667 & ~x670 & ~x693 & ~x700 & ~x747 & ~x751;
assign c7119 =  x687 & ~x111 & ~x224 & ~x282 & ~x361 & ~x364 & ~x391 & ~x393 & ~x417 & ~x420 & ~x446 & ~x447 & ~x475 & ~x504 & ~x506 & ~x507 & ~x534 & ~x561 & ~x563 & ~x588 & ~x589 & ~x591 & ~x617 & ~x619 & ~x620 & ~x621 & ~x644 & ~x645 & ~x676 & ~x701 & ~x728 & ~x730 & ~x753 & ~x755 & ~x758 & ~x782 & ~x783;
assign c7121 =  x665 & ~x518 & ~x545 & ~x573;
assign c7123 =  x714 &  x741 & ~x224 & ~x303 & ~x363 & ~x500 & ~x557 & ~x559 & ~x590;
assign c7125 = ~x144 & ~x212 & ~x239 & ~x240 & ~x267 & ~x295 & ~x322 & ~x323 & ~x324 & ~x350 & ~x351 & ~x726 & ~x753 & ~x755 & ~x758 & ~x779 & ~x782;
assign c7127 = ~x25 & ~x80 & ~x108 & ~x347 & ~x373 & ~x399 & ~x401 & ~x427 & ~x428 & ~x454 & ~x480 & ~x481;
assign c7129 = ~x462 & ~x489 & ~x490 & ~x491 & ~x518 & ~x543;
assign c7131 =  x283 & ~x19 & ~x23 & ~x24 & ~x26 & ~x27 & ~x95 & ~x151 & ~x364 & ~x772;
assign c7133 = ~x138 & ~x195 & ~x252 & ~x455 & ~x456 & ~x482 & ~x483 & ~x484 & ~x508 & ~x510 & ~x535 & ~x536 & ~x560;
assign c7135 =  x284 &  x620 & ~x223;
assign c7137 =  x742 & ~x194 & ~x227 & ~x252 & ~x281 & ~x389 & ~x628;
assign c7139 =  x540 & ~x27 & ~x225 & ~x326 & ~x381 & ~x394 & ~x476 & ~x708 & ~x756 & ~x759;
assign c7141 = ~x384 & ~x410 & ~x411 & ~x438 & ~x439 & ~x463 & ~x465 & ~x491 & ~x513 & ~x518 & ~x519 & ~x520 & ~x546;
assign c7143 = ~x14 & ~x84 & ~x347 & ~x373 & ~x427 & ~x481 & ~x507 & ~x509 & ~x587 & ~x589 & ~x616 & ~x618 & ~x669 & ~x726 & ~x729 & ~x752 & ~x776 & ~x778;
assign c7145 = ~x4 & ~x52 & ~x54 & ~x139 & ~x194 & ~x219 & ~x255 & ~x277 & ~x332 & ~x333 & ~x362 & ~x396 & ~x416 & ~x440 & ~x581 & ~x582 & ~x584 & ~x593 & ~x624;
assign c7147 =  x640 & ~x21 & ~x26 & ~x28 & ~x66 & ~x122 & ~x139 & ~x762 & ~x763;
assign c7149 = ~x0 & ~x3 & ~x26 & ~x27 & ~x28 & ~x29 & ~x31 & ~x141 & ~x162 & ~x169 & ~x196 & ~x197 & ~x199 & ~x217 & ~x219 & ~x220 & ~x224 & ~x227 & ~x246 & ~x248 & ~x277 & ~x279 & ~x309 & ~x332 & ~x335 & ~x361 & ~x362 & ~x364 & ~x390 & ~x417 & ~x420 & ~x445 & ~x446 & ~x447 & ~x476 & ~x559 & ~x628 & ~x629;
assign c7151 = ~x2 & ~x14 & ~x57 & ~x185 & ~x212 & ~x267 & ~x296 & ~x322 & ~x352 & ~x587 & ~x616 & ~x759 & ~x779;
assign c7153 = ~x2 & ~x3 & ~x32 & ~x376 & ~x405 & ~x432 & ~x488 & ~x515 & ~x541 & ~x707 & ~x728 & ~x732 & ~x740 & ~x768 & ~x780;
assign c7155 = ~x18 & ~x45 & ~x107 & ~x134 & ~x138 & ~x163 & ~x166 & ~x194 & ~x240 & ~x268 & ~x322 & ~x323 & ~x351 & ~x392 & ~x393 & ~x757;
assign c7157 =  x742 & ~x107 & ~x471 & ~x472 & ~x534;
assign c7159 =  x205 & ~x12 & ~x71 & ~x72 & ~x99 & ~x190 & ~x194 & ~x364 & ~x397 & ~x424 & ~x476 & ~x532;
assign c7161 =  x379 &  x407 &  x434 &  x462 & ~x0 & ~x21 & ~x51 & ~x55 & ~x56 & ~x67 & ~x68 & ~x123 & ~x559 & ~x727 & ~x728 & ~x732;
assign c7163 =  x204 &  x233 & ~x100 & ~x128 & ~x341 & ~x366 & ~x611;
assign c7165 = ~x93 & ~x109 & ~x137 & ~x405 & ~x413 & ~x432 & ~x485 & ~x486;
assign c7167 = ~x3 & ~x8 & ~x86 & ~x161 & ~x163 & ~x190 & ~x219 & ~x222 & ~x275 & ~x336 & ~x361 & ~x388 & ~x389 & ~x390 & ~x447 & ~x500 & ~x529 & ~x531 & ~x562 & ~x587 & ~x593 & ~x638 & ~x647 & ~x650 & ~x652 & ~x665 & ~x731;
assign c7169 = ~x15 & ~x17 & ~x46 & ~x50 & ~x51 & ~x111 & ~x138 & ~x160 & ~x187 & ~x268 & ~x295 & ~x394 & ~x421 & ~x422 & ~x477 & ~x504 & ~x616 & ~x638 & ~x640 & ~x641 & ~x667 & ~x700 & ~x728 & ~x729 & ~x730 & ~x731 & ~x753 & ~x759;
assign c7171 =  x633 &  x660 &  x715 & ~x28 & ~x560 & ~x617 & ~x618 & ~x619 & ~x694 & ~x720;
assign c7173 = ~x28 & ~x234 & ~x463 & ~x491 & ~x519 & ~x547 & ~x574 & ~x600 & ~x601 & ~x756;
assign c7175 = ~x207 & ~x235 & ~x345 & ~x418 & ~x419 & ~x447 & ~x475 & ~x476 & ~x588 & ~x741;
assign c7177 = ~x54 & ~x132 & ~x137 & ~x138 & ~x195 & ~x249 & ~x273 & ~x361 & ~x452 & ~x453 & ~x477 & ~x511;
assign c7179 =  x715 & ~x17 & ~x84 & ~x166 & ~x195 & ~x227 & ~x251 & ~x254 & ~x284 & ~x312 & ~x389 & ~x391 & ~x470 & ~x471 & ~x502 & ~x504 & ~x644 & ~x645 & ~x756 & ~x764;
assign c7181 =  x261 &  x289 & ~x194 & ~x196 & ~x249 & ~x252 & ~x274 & ~x302 & ~x306 & ~x424 & ~x448 & ~x452 & ~x479 & ~x480 & ~x504 & ~x508 & ~x644;
assign c7183 = ~x2 & ~x55 & ~x57 & ~x58 & ~x59 & ~x139 & ~x145 & ~x190 & ~x268 & ~x279 & ~x296 & ~x308 & ~x309 & ~x323 & ~x350 & ~x351 & ~x366 & ~x705 & ~x754 & ~x783;
assign c7185 = ~x3 & ~x138 & ~x228 & ~x456 & ~x475 & ~x479 & ~x484 & ~x505 & ~x532 & ~x562 & ~x563 & ~x619 & ~x647 & ~x703;
assign c7187 = ~x30 & ~x150 & ~x226 & ~x249 & ~x276 & ~x279 & ~x334 & ~x363 & ~x444 & ~x473 & ~x474 & ~x601 & ~x756 & ~x783;
assign c7189 = ~x25 & ~x196 & ~x224 & ~x290 & ~x291 & ~x316 & ~x318 & ~x345 & ~x371 & ~x420 & ~x531 & ~x751 & ~x762 & ~x776;
assign c7191 =  x583 & ~x571 & ~x573;
assign c7193 = ~x26 & ~x35 & ~x55 & ~x63 & ~x140 & ~x189 & ~x190 & ~x221 & ~x278 & ~x281 & ~x361 & ~x362 & ~x445 & ~x513 & ~x514 & ~x584 & ~x671 & ~x727 & ~x752 & ~x755 & ~x782;
assign c7195 = ~x26 & ~x27 & ~x145 & ~x379 & ~x433 & ~x434 & ~x460 & ~x461 & ~x487 & ~x514 & ~x515 & ~x649;
assign c7197 = ~x19 & ~x39 & ~x122 & ~x178 & ~x411 & ~x467 & ~x519 & ~x625 & ~x773;
assign c7199 = ~x14 & ~x24 & ~x30 & ~x48 & ~x73 & ~x75 & ~x112 & ~x137 & ~x166 & ~x323 & ~x365 & ~x393 & ~x679 & ~x702 & ~x725 & ~x739 & ~x765 & ~x780 & ~x781;
assign c7201 =  x87 & ~x391;
assign c7203 =  x257 &  x438 &  x466 &  x493 & ~x390 & ~x755 & ~x783;
assign c7205 = ~x109 & ~x245 & ~x248 & ~x250 & ~x274 & ~x277 & ~x390 & ~x446 & ~x474 & ~x485 & ~x511 & ~x539 & ~x618;
assign c7207 =  x153 & ~x197 & ~x199 & ~x203 & ~x358 & ~x359 & ~x362 & ~x385 & ~x388 & ~x420 & ~x508 & ~x585 & ~x611 & ~x618 & ~x734;
assign c7209 =  x157 &  x185 &  x213 & ~x389 & ~x399 & ~x446;
assign c7211 =  x466 &  x493 & ~x1 & ~x23 & ~x55 & ~x112 & ~x304 & ~x305 & ~x307 & ~x332 & ~x334 & ~x360 & ~x361 & ~x362 & ~x390 & ~x391 & ~x504 & ~x636 & ~x692;
assign c7213 = ~x8 & ~x110 & ~x188 & ~x192 & ~x216 & ~x219 & ~x221 & ~x279 & ~x281 & ~x362 & ~x390 & ~x395 & ~x449 & ~x451 & ~x606 & ~x645 & ~x661 & ~x696 & ~x758 & ~x782;
assign c7215 = ~x135 & ~x136 & ~x169 & ~x278 & ~x303 & ~x305 & ~x331 & ~x359 & ~x360 & ~x361 & ~x362 & ~x389 & ~x393 & ~x417 & ~x419 & ~x445 & ~x448 & ~x449 & ~x560 & ~x610 & ~x635 & ~x638 & ~x690 & ~x692 & ~x694 & ~x722 & ~x723 & ~x747 & ~x761;
assign c7217 =  x458 &  x486 &  x688 & ~x58 & ~x546 & ~x573;
assign c7219 =  x561 & ~x1 & ~x27 & ~x688 & ~x689 & ~x716 & ~x761 & ~x764;
assign c7221 =  x313 &  x566 & ~x0 & ~x7 & ~x17 & ~x44 & ~x111 & ~x775 & ~x777 & ~x782;
assign c7223 = ~x1 & ~x2 & ~x183 & ~x211 & ~x267 & ~x268 & ~x269 & ~x271 & ~x323 & ~x324 & ~x671 & ~x698 & ~x699 & ~x755 & ~x779;
assign c7225 =  x436 & ~x341 & ~x415 & ~x425 & ~x469 & ~x608;
assign c7227 =  x353 &  x436 & ~x362 & ~x418 & ~x446 & ~x458 & ~x474;
assign c7229 = ~x52 & ~x74 & ~x140 & ~x194 & ~x217 & ~x223 & ~x246 & ~x277 & ~x279 & ~x307 & ~x394 & ~x396 & ~x421 & ~x496 & ~x500 & ~x506 & ~x530 & ~x611 & ~x666 & ~x671 & ~x693 & ~x695 & ~x704 & ~x731 & ~x756;
assign c7231 = ~x0 & ~x99 & ~x153 & ~x181 & ~x209 & ~x239 & ~x554 & ~x616;
assign c7233 = ~x28 & ~x56 & ~x84 & ~x140 & ~x141 & ~x165 & ~x168 & ~x217 & ~x224 & ~x246 & ~x248 & ~x251 & ~x273 & ~x275 & ~x276 & ~x278 & ~x328 & ~x330 & ~x331 & ~x332 & ~x336 & ~x360 & ~x385 & ~x389 & ~x390 & ~x391 & ~x416 & ~x421 & ~x442 & ~x443 & ~x444 & ~x472 & ~x473 & ~x475 & ~x499 & ~x502 & ~x504 & ~x558 & ~x671;
assign c7235 = ~x1 & ~x2 & ~x15 & ~x23 & ~x49 & ~x53 & ~x69 & ~x182 & ~x336 & ~x495 & ~x504 & ~x645 & ~x669 & ~x671 & ~x757 & ~x777;
assign c7237 = ~x27 & ~x178 & ~x207 & ~x304 & ~x332 & ~x333 & ~x335 & ~x390 & ~x391 & ~x416 & ~x419 & ~x447 & ~x734;
assign c7239 = ~x23 & ~x27 & ~x55 & ~x81 & ~x110 & ~x139 & ~x167 & ~x436 & ~x463 & ~x464 & ~x517 & ~x518 & ~x543 & ~x727 & ~x765;
assign c7241 = ~x63 & ~x167 & ~x221 & ~x249 & ~x275 & ~x305 & ~x306 & ~x311 & ~x332 & ~x422 & ~x470 & ~x511 & ~x540;
assign c7243 = ~x5 & ~x21 & ~x82 & ~x85 & ~x110 & ~x111 & ~x112 & ~x114 & ~x134 & ~x164 & ~x167 & ~x171 & ~x192 & ~x222 & ~x254 & ~x304 & ~x305 & ~x306 & ~x308 & ~x333 & ~x334 & ~x362 & ~x392 & ~x432 & ~x447 & ~x458 & ~x459 & ~x474 & ~x615 & ~x620 & ~x671 & ~x728;
assign c7245 =  x313 &  x647 & ~x22;
assign c7247 = ~x55 & ~x111 & ~x378 & ~x379 & ~x404 & ~x406 & ~x434 & ~x460 & ~x488 & ~x514 & ~x515 & ~x570 & ~x700 & ~x707 & ~x708 & ~x757 & ~x762;
assign c7249 =  x379 &  x631 & ~x24 & ~x445 & ~x483 & ~x563;
assign c7251 =  x287 & ~x0 & ~x97 & ~x155 & ~x180 & ~x645 & ~x734 & ~x757;
assign c7253 = ~x9 & ~x11 & ~x39 & ~x66 & ~x94 & ~x180 & ~x181 & ~x237 & ~x264;
assign c7255 =  x356 &  x384 &  x413 & ~x21 & ~x111 & ~x112 & ~x115 & ~x142 & ~x224 & ~x334 & ~x362 & ~x446 & ~x560;
assign c7257 = ~x1 & ~x39 & ~x67 & ~x84 & ~x168 & ~x252 & ~x280 & ~x292 & ~x318 & ~x320 & ~x364;
assign c7259 =  x745 &  x772 & ~x138 & ~x248 & ~x253 & ~x418 & ~x555;
assign c7261 = ~x76 & ~x79 & ~x135 & ~x140 & ~x191 & ~x220 & ~x256 & ~x331 & ~x334 & ~x337 & ~x359 & ~x387 & ~x394 & ~x395 & ~x444 & ~x504 & ~x538 & ~x539 & ~x590;
assign c7263 = ~x42 & ~x46 & ~x98 & ~x126 & ~x128 & ~x155 & ~x265 & ~x266 & ~x616 & ~x645;
assign c7265 =  x517 & ~x227 & ~x255 & ~x279 & ~x328 & ~x361 & ~x472 & ~x481 & ~x534 & ~x588 & ~x589 & ~x616 & ~x668 & ~x675;
assign c7267 = ~x101 & ~x106 & ~x137 & ~x347 & ~x402 & ~x425 & ~x428 & ~x536 & ~x619 & ~x646;
assign c7269 = ~x66 & ~x151 & ~x208 & ~x209 & ~x364 & ~x525 & ~x554 & ~x561 & ~x616 & ~x757;
assign c7271 = ~x112 & ~x349 & ~x404 & ~x431 & ~x432 & ~x486 & ~x514 & ~x515 & ~x541 & ~x569 & ~x570 & ~x651 & ~x676 & ~x679 & ~x705 & ~x708 & ~x730;
assign c7273 =  x183 & ~x56 & ~x78 & ~x79 & ~x108 & ~x112 & ~x135 & ~x142 & ~x162 & ~x163 & ~x167 & ~x192 & ~x193 & ~x194 & ~x195 & ~x219 & ~x220 & ~x226 & ~x278 & ~x280 & ~x308 & ~x361 & ~x389 & ~x419 & ~x445 & ~x452;
assign c7275 = ~x0 & ~x25 & ~x52 & ~x139 & ~x378 & ~x404 & ~x405 & ~x432 & ~x456 & ~x459 & ~x512 & ~x513 & ~x672 & ~x699;
assign c7277 = ~x8 & ~x11 & ~x37 & ~x124 & ~x179 & ~x215 & ~x418 & ~x446 & ~x447 & ~x503;
assign c7279 =  x437 & ~x23 & ~x82 & ~x222 & ~x247 & ~x278 & ~x362 & ~x392 & ~x571 & ~x572 & ~x748 & ~x776;
assign c7281 = ~x1 & ~x2 & ~x48 & ~x56 & ~x58 & ~x76 & ~x82 & ~x107 & ~x110 & ~x172 & ~x251 & ~x325 & ~x326 & ~x353 & ~x382 & ~x410 & ~x662 & ~x716 & ~x717 & ~x727 & ~x742 & ~x748 & ~x761;
assign c7283 = ~x110 & ~x223 & ~x376 & ~x377 & ~x448;
assign c7285 = ~x94 & ~x236 & ~x237 & ~x263 & ~x411 & ~x412 & ~x439;
assign c7287 =  x435 &  x461 &  x488 & ~x162 & ~x418 & ~x444 & ~x472 & ~x579 & ~x590 & ~x593 & ~x646 & ~x678 & ~x781;
assign c7289 =  x497 &  x525 &  x580 & ~x224 & ~x533 & ~x559 & ~x589 & ~x618 & ~x671;
assign c7291 = ~x8 & ~x43 & ~x53 & ~x99 & ~x104 & ~x109 & ~x129 & ~x184 & ~x690 & ~x703 & ~x759;
assign c7293 = ~x19 & ~x28 & ~x32 & ~x33 & ~x55 & ~x349 & ~x376 & ~x377 & ~x404 & ~x459 & ~x486 & ~x513 & ~x540 & ~x704 & ~x705 & ~x706 & ~x732 & ~x733 & ~x754;
assign c7295 =  x256 &  x537 & ~x419 & ~x706 & ~x735;
assign c7297 =  x773 & ~x474 & ~x631 & ~x632;
assign c7299 = ~x11 & ~x28 & ~x38 & ~x93 & ~x291 & ~x392 & ~x400 & ~x475 & ~x668;
assign c7301 =  x527 &  x582;
assign c7303 =  x622 & ~x18 & ~x19 & ~x24 & ~x25 & ~x26 & ~x53 & ~x83 & ~x98 & ~x99 & ~x112 & ~x140 & ~x252 & ~x783;
assign c7305 =  x183 & ~x8 & ~x107 & ~x221 & ~x244 & ~x248 & ~x252 & ~x359 & ~x472 & ~x499;
assign c7307 =  x189 & ~x223 & ~x249 & ~x252 & ~x418 & ~x558 & ~x587;
assign c7309 =  x705 & ~x251 & ~x635;
assign c7311 =  x527 & ~x402 & ~x482;
assign c7313 =  x719 & ~x55 & ~x254 & ~x281 & ~x282 & ~x361 & ~x362 & ~x392 & ~x394 & ~x472 & ~x504 & ~x505 & ~x530 & ~x557 & ~x586 & ~x590 & ~x646 & ~x673 & ~x674 & ~x702 & ~x732 & ~x760;
assign c7315 =  x651 &  x679 &  x681 &  x682 & ~x25 & ~x111 & ~x141 & ~x169 & ~x223;
assign c7317 = ~x27 & ~x50 & ~x53 & ~x54 & ~x68 & ~x80 & ~x330 & ~x343 & ~x384 & ~x413 & ~x419 & ~x440 & ~x469;
assign c7319 =  x42 &  x181 & ~x119 & ~x148;
assign c7321 = ~x17 & ~x44 & ~x134 & ~x165 & ~x227 & ~x267 & ~x366 & ~x575;
assign c7323 = ~x1 & ~x140 & ~x235 & ~x244 & ~x262 & ~x290 & ~x318 & ~x571;
assign c7325 =  x155 &  x715 & ~x26 & ~x84 & ~x107 & ~x169 & ~x222 & ~x282 & ~x283 & ~x365 & ~x418 & ~x530 & ~x643 & ~x758 & ~x759;
assign c7327 = ~x37 & ~x81 & ~x83 & ~x112 & ~x127 & ~x128 & ~x155 & ~x183 & ~x267 & ~x336 & ~x365 & ~x588 & ~x707 & ~x767;
assign c7329 = ~x16 & ~x18 & ~x72 & ~x88 & ~x128 & ~x182 & ~x267 & ~x683 & ~x750;
assign c7331 = ~x27 & ~x80 & ~x137 & ~x138 & ~x162 & ~x195 & ~x226 & ~x332 & ~x413 & ~x415 & ~x416 & ~x424 & ~x440 & ~x468 & ~x478 & ~x498 & ~x500 & ~x525 & ~x526 & ~x533 & ~x554 & ~x611 & ~x622 & ~x638 & ~x674 & ~x706 & ~x737;
assign c7333 = ~x27 & ~x84 & ~x112 & ~x140 & ~x173 & ~x195 & ~x223 & ~x438 & ~x464 & ~x465 & ~x466 & ~x492 & ~x518 & ~x519 & ~x520 & ~x521 & ~x548 & ~x574 & ~x575 & ~x602;
assign c7335 = ~x51 & ~x100 & ~x159 & ~x251 & ~x382 & ~x384 & ~x412 & ~x440 & ~x466 & ~x494 & ~x700 & ~x718 & ~x723 & ~x778;
assign c7337 = ~x85 & ~x141 & ~x297 & ~x298 & ~x323 & ~x353 & ~x381 & ~x411 & ~x438 & ~x749 & ~x783;
assign c7339 = ~x23 & ~x25 & ~x26 & ~x27 & ~x54 & ~x85 & ~x111 & ~x140 & ~x165 & ~x166 & ~x167 & ~x168 & ~x169 & ~x196 & ~x197 & ~x199 & ~x202 & ~x227 & ~x252 & ~x308 & ~x400 & ~x401 & ~x428 & ~x504 & ~x588 & ~x616 & ~x618 & ~x644 & ~x672 & ~x673 & ~x700 & ~x728 & ~x754 & ~x781 & ~x783;
assign c7341 =  x639 &  x640 & ~x55 & ~x139 & ~x193 & ~x251;
assign c7343 =  x608 & ~x1 & ~x55 & ~x517 & ~x518 & ~x531 & ~x559;
assign c7345 =  x501 & ~x495 & ~x523 & ~x524 & ~x551 & ~x552 & ~x579 & ~x606;
assign c7347 =  x590 & ~x413 & ~x659 & ~x686 & ~x713;
assign c7349 = ~x13 & ~x37 & ~x96 & ~x151 & ~x154 & ~x155 & ~x335 & ~x337 & ~x420 & ~x558 & ~x586 & ~x614 & ~x615 & ~x616 & ~x644 & ~x755 & ~x759;
assign c7351 = ~x6 & ~x24 & ~x29 & ~x241 & ~x242 & ~x271 & ~x327 & ~x355 & ~x383 & ~x530 & ~x557 & ~x614 & ~x641 & ~x642 & ~x666 & ~x698 & ~x720 & ~x724 & ~x725 & ~x727 & ~x751 & ~x754 & ~x768 & ~x776 & ~x782;
assign c7353 =  x462 & ~x110 & ~x191 & ~x221 & ~x276 & ~x417 & ~x473 & ~x479 & ~x535 & ~x538;
assign c7355 =  x566 & ~x0 & ~x23 & ~x24 & ~x25 & ~x28 & ~x29 & ~x45 & ~x46 & ~x48 & ~x49 & ~x51 & ~x55 & ~x56 & ~x57 & ~x73 & ~x74 & ~x79 & ~x81 & ~x86 & ~x99 & ~x105 & ~x114 & ~x137 & ~x195 & ~x250 & ~x251 & ~x308 & ~x364 & ~x586 & ~x737 & ~x738 & ~x740 & ~x755 & ~x760 & ~x765 & ~x767;
assign c7357 =  x184 & ~x1 & ~x57 & ~x79 & ~x84 & ~x108 & ~x110 & ~x112 & ~x114 & ~x136 & ~x138 & ~x169 & ~x192 & ~x197 & ~x226 & ~x250 & ~x275 & ~x303 & ~x307 & ~x335 & ~x338 & ~x362 & ~x363 & ~x391 & ~x419 & ~x528 & ~x529 & ~x585 & ~x672;
assign c7359 =  x718 &  x773 & ~x283 & ~x311 & ~x338 & ~x617 & ~x701;
assign c7361 =  x156 & ~x26 & ~x53 & ~x55 & ~x233 & ~x250 & ~x280 & ~x281 & ~x306 & ~x335 & ~x391 & ~x418 & ~x446 & ~x475 & ~x476 & ~x559;
assign c7363 = ~x1 & ~x358 & ~x415 & ~x416 & ~x451 & ~x480 & ~x595;
assign c7365 = ~x1 & ~x294 & ~x321 & ~x377 & ~x404 & ~x431 & ~x486 & ~x513 & ~x643 & ~x671 & ~x766;
assign c7367 =  x434 & ~x123 & ~x307 & ~x447 & ~x473 & ~x749 & ~x779;
assign c7369 = ~x24 & ~x109 & ~x113 & ~x135 & ~x137 & ~x141 & ~x199 & ~x228 & ~x247 & ~x250 & ~x311 & ~x332 & ~x333 & ~x364 & ~x388 & ~x417 & ~x419 & ~x424 & ~x470 & ~x471 & ~x476 & ~x527 & ~x529 & ~x538 & ~x554 & ~x557 & ~x558 & ~x616 & ~x643 & ~x734 & ~x782;
assign c7371 = ~x37 & ~x109 & ~x219 & ~x221 & ~x246 & ~x247 & ~x311 & ~x472 & ~x500 & ~x512 & ~x565 & ~x759;
assign c7373 =  x451 &  x479 & ~x575 & ~x602 & ~x628;
assign c7375 =  x537 & ~x17 & ~x28 & ~x269 & ~x296 & ~x297 & ~x324 & ~x325 & ~x351 & ~x643;
assign c7377 =  x480 &  x507 & ~x4 & ~x322 & ~x688 & ~x780 & ~x783;
assign c7379 =  x463 & ~x56 & ~x195 & ~x222 & ~x224 & ~x226 & ~x249 & ~x305 & ~x307 & ~x337 & ~x338 & ~x361 & ~x504 & ~x526 & ~x554 & ~x581 & ~x584 & ~x610 & ~x619 & ~x635 & ~x673;
assign c7381 = ~x0 & ~x6 & ~x10 & ~x168 & ~x351 & ~x378 & ~x405 & ~x407 & ~x433 & ~x435 & ~x461 & ~x490 & ~x517 & ~x542 & ~x755;
assign c7383 = ~x124 & ~x180 & ~x384 & ~x396 & ~x414 & ~x421 & ~x528 & ~x671;
assign c7385 =  x439 &  x495 & ~x4 & ~x51 & ~x52 & ~x55 & ~x56 & ~x58 & ~x59 & ~x111 & ~x140 & ~x224 & ~x252 & ~x280 & ~x335 & ~x363 & ~x391 & ~x418 & ~x419 & ~x473 & ~x501 & ~x506 & ~x531 & ~x672;
assign c7387 = ~x16 & ~x17 & ~x37 & ~x180 & ~x208 & ~x418 & ~x446 & ~x529 & ~x587 & ~x642;
assign c7389 = ~x1 & ~x5 & ~x6 & ~x56 & ~x83 & ~x111 & ~x113 & ~x133 & ~x166 & ~x168 & ~x193 & ~x223 & ~x224 & ~x252 & ~x279 & ~x307 & ~x392 & ~x546 & ~x572 & ~x573 & ~x599 & ~x600 & ~x601 & ~x746 & ~x774;
assign c7391 = ~x4 & ~x33 & ~x55 & ~x109 & ~x136 & ~x273 & ~x274 & ~x276 & ~x302 & ~x304 & ~x330 & ~x332 & ~x384 & ~x385 & ~x396 & ~x416 & ~x445 & ~x450 & ~x471 & ~x500 & ~x558 & ~x564 & ~x582 & ~x583 & ~x611 & ~x645 & ~x677 & ~x726 & ~x730 & ~x776;
assign c7393 =  x576 &  x603 &  x604 & ~x78 & ~x80 & ~x169 & ~x446 & ~x447 & ~x452 & ~x477 & ~x481 & ~x482 & ~x510 & ~x532 & ~x588 & ~x699 & ~x725 & ~x755;
assign c7395 =  x284 & ~x1 & ~x83 & ~x140 & ~x207 & ~x235 & ~x336 & ~x419 & ~x756;
assign c7397 = ~x79 & ~x89 & ~x225 & ~x245 & ~x247 & ~x276 & ~x303 & ~x313 & ~x359 & ~x385 & ~x414 & ~x423 & ~x424 & ~x425 & ~x471 & ~x499 & ~x584 & ~x611 & ~x707;
assign c7399 =  x204 &  x232 & ~x54 & ~x55 & ~x71 & ~x98 & ~x99 & ~x125 & ~x126 & ~x209 & ~x365 & ~x392 & ~x559 & ~x699;
assign c7401 =  x499 &  x554 & ~x27 & ~x573 & ~x587 & ~x756;
assign c7403 =  x437 &  x492 & ~x1 & ~x415 & ~x418 & ~x562 & ~x592;
assign c7405 =  x629 & ~x400 & ~x428 & ~x768;
assign c7407 = ~x0 & ~x3 & ~x14 & ~x15 & ~x17 & ~x27 & ~x124 & ~x126 & ~x152 & ~x153 & ~x180 & ~x181 & ~x364 & ~x420 & ~x532 & ~x583 & ~x616 & ~x728 & ~x775 & ~x783;
assign c7409 = ~x55 & ~x84 & ~x92 & ~x466 & ~x495 & ~x520 & ~x547 & ~x625;
assign c7411 = ~x53 & ~x107 & ~x274 & ~x284 & ~x304 & ~x327 & ~x330 & ~x332 & ~x333 & ~x335 & ~x339 & ~x356 & ~x359 & ~x387 & ~x416 & ~x446 & ~x555 & ~x776;
assign c7413 = ~x127 & ~x378 & ~x406 & ~x433 & ~x544 & ~x572 & ~x626;
assign c7415 = ~x27 & ~x83 & ~x263 & ~x317 & ~x318 & ~x344 & ~x444 & ~x473 & ~x691;
assign c7417 =  x522 &  x577 &  x578 &  x604 & ~x51 & ~x80 & ~x84 & ~x168 & ~x169 & ~x335 & ~x363 & ~x390 & ~x418 & ~x419 & ~x473 & ~x475 & ~x501 & ~x644 & ~x756 & ~x757;
assign c7419 =  x284 &  x564 & ~x18 & ~x448 & ~x588;
assign c7421 =  x555 &  x608 &  x610 &  x636 & ~x168 & ~x196 & ~x559;
assign c7423 =  x243 &  x270 &  x298 & ~x81 & ~x100 & ~x196 & ~x363 & ~x447 & ~x480 & ~x506 & ~x508 & ~x591 & ~x644;
assign c7425 =  x745 &  x772;
assign c7427 = ~x29 & ~x158 & ~x159 & ~x191 & ~x194 & ~x284 & ~x429 & ~x455;
assign c7429 =  x417 &  x473 & ~x27 & ~x382 & ~x439 & ~x467 & ~x523 & ~x616;
assign c7431 = ~x22 & ~x53 & ~x67 & ~x111 & ~x164 & ~x167 & ~x168 & ~x308 & ~x373 & ~x429 & ~x456;
assign c7433 =  x603 & ~x0 & ~x10 & ~x11 & ~x12 & ~x25 & ~x26 & ~x27 & ~x29 & ~x56 & ~x263 & ~x418 & ~x445 & ~x447 & ~x473 & ~x475 & ~x501 & ~x531 & ~x558 & ~x670 & ~x750 & ~x763 & ~x764 & ~x777 & ~x779 & ~x783;
assign c7435 = ~x196 & ~x220 & ~x249 & ~x333 & ~x334 & ~x375 & ~x390 & ~x404 & ~x431 & ~x742 & ~x761 & ~x778;
assign c7437 =  x134 &  x496 &  x524 & ~x24 & ~x53 & ~x447;
assign c7439 =  x556 &  x583 &  x637 & ~x109 & ~x756;
assign c7441 =  x258 & ~x95 & ~x96 & ~x97 & ~x152 & ~x179 & ~x180 & ~x502;
assign c7443 = ~x5 & ~x17 & ~x55 & ~x109 & ~x158 & ~x163 & ~x212 & ~x240 & ~x242 & ~x476 & ~x500 & ~x557 & ~x606 & ~x607 & ~x614 & ~x725 & ~x756 & ~x778;
assign c7445 = ~x14 & ~x42 & ~x45 & ~x129 & ~x155 & ~x182 & ~x211 & ~x212 & ~x239 & ~x267 & ~x420 & ~x559 & ~x616 & ~x620 & ~x646 & ~x673 & ~x699 & ~x704 & ~x726 & ~x758;
assign c7447 = ~x73 & ~x98 & ~x153 & ~x154 & ~x210 & ~x365 & ~x414 & ~x442 & ~x469 & ~x776;
assign c7449 =  x437 & ~x1 & ~x2 & ~x55 & ~x111 & ~x140 & ~x142 & ~x196 & ~x197 & ~x250 & ~x251 & ~x253 & ~x278 & ~x280 & ~x307 & ~x308 & ~x309 & ~x333 & ~x337 & ~x361 & ~x364 & ~x389 & ~x390 & ~x391 & ~x445 & ~x473 & ~x530 & ~x531 & ~x556 & ~x664 & ~x694 & ~x700 & ~x720 & ~x748 & ~x751 & ~x779;
assign c7451 =  x646 & ~x26 & ~x112 & ~x487;
assign c7453 = ~x54 & ~x111 & ~x112 & ~x202 & ~x223 & ~x251 & ~x518 & ~x519 & ~x521 & ~x546 & ~x548 & ~x600 & ~x601 & ~x628;
assign c7455 =  x295 & ~x83 & ~x114 & ~x360 & ~x362 & ~x389 & ~x390 & ~x428 & ~x471 & ~x475 & ~x528 & ~x558 & ~x559 & ~x587;
assign c7457 =  x143 & ~x26 & ~x27 & ~x39 & ~x83 & ~x168 & ~x280 & ~x308;
assign c7459 =  x315 & ~x12 & ~x67 & ~x69 & ~x96 & ~x124 & ~x125 & ~x152 & ~x441 & ~x781;
assign c7461 = ~x2 & ~x84 & ~x137 & ~x151 & ~x179 & ~x402 & ~x513 & ~x726;
assign c7463 = ~x42 & ~x43 & ~x55 & ~x56 & ~x98 & ~x100 & ~x126 & ~x127 & ~x155 & ~x236 & ~x237 & ~x672 & ~x729 & ~x757 & ~x759 & ~x783;
assign c7465 =  x201 &  x229 &  x230 &  x567 & ~x447 & ~x757;
assign c7467 = ~x40 & ~x47 & ~x78 & ~x79 & ~x135 & ~x329 & ~x357 & ~x387 & ~x412 & ~x414 & ~x442 & ~x468 & ~x469 & ~x682 & ~x700 & ~x728 & ~x735 & ~x736 & ~x737 & ~x755;
assign c7469 =  x433 &  x460 & ~x212 & ~x496 & ~x523 & ~x550 & ~x577 & ~x579 & ~x605 & ~x608 & ~x633 & ~x755;
assign c7471 = ~x8 & ~x75 & ~x76 & ~x138 & ~x188 & ~x189 & ~x193 & ~x219 & ~x220 & ~x224 & ~x247 & ~x248 & ~x309 & ~x311 & ~x338 & ~x340 & ~x366 & ~x368 & ~x497 & ~x553 & ~x581 & ~x588 & ~x611 & ~x616 & ~x620 & ~x636 & ~x644 & ~x646 & ~x667 & ~x676 & ~x678 & ~x705 & ~x728 & ~x730 & ~x759 & ~x762 & ~x763 & ~x782;
assign c7473 = ~x25 & ~x42 & ~x44 & ~x45 & ~x103 & ~x155 & ~x184 & ~x210 & ~x239 & ~x589 & ~x592 & ~x613 & ~x615 & ~x645 & ~x752 & ~x756 & ~x760;
assign c7475 = ~x2 & ~x83 & ~x111 & ~x435 & ~x436 & ~x461 & ~x462 & ~x463 & ~x489 & ~x490 & ~x491 & ~x517 & ~x518 & ~x543 & ~x570 & ~x598 & ~x625 & ~x652;
assign c7477 = ~x119 & ~x162 & ~x167 & ~x191 & ~x193 & ~x284 & ~x301 & ~x305 & ~x312 & ~x313 & ~x341 & ~x424 & ~x451 & ~x452 & ~x480 & ~x509 & ~x511;
assign c7479 =  x496 &  x524 &  x552 & ~x2 & ~x24 & ~x83 & ~x84 & ~x85 & ~x112 & ~x140 & ~x168 & ~x252 & ~x280 & ~x308 & ~x336 & ~x391 & ~x418 & ~x446 & ~x447 & ~x448 & ~x474 & ~x475 & ~x476 & ~x504 & ~x671 & ~x755 & ~x756 & ~x758 & ~x761;
assign c7481 =  x634 & ~x9 & ~x548 & ~x627;
assign c7483 =  x285 & ~x28 & ~x66 & ~x180 & ~x392 & ~x699;
assign c7485 =  x649 &  x707 & ~x251;
assign c7487 =  x230 &  x577 &  x604 &  x658 & ~x27 & ~x55 & ~x56 & ~x85 & ~x420 & ~x476 & ~x532 & ~x757;
assign c7489 =  x686 & ~x81 & ~x367 & ~x391 & ~x396 & ~x472 & ~x475 & ~x525 & ~x590 & ~x734;
assign c7491 =  x164 & ~x0 & ~x3 & ~x26 & ~x42 & ~x55 & ~x70 & ~x246 & ~x274 & ~x302 & ~x330 & ~x392 & ~x420;
assign c7493 =  x326 &  x353 & ~x27 & ~x54 & ~x82 & ~x139 & ~x194 & ~x390 & ~x391 & ~x474 & ~x533 & ~x592 & ~x593 & ~x619 & ~x621 & ~x643;
assign c7495 =  x203 & ~x14 & ~x15 & ~x17 & ~x69 & ~x182 & ~x209 & ~x237 & ~x697;
assign c7497 = ~x157 & ~x183 & ~x238 & ~x239 & ~x264 & ~x293 & ~x392 & ~x668 & ~x698 & ~x723 & ~x755;
assign c7499 =  x314 &  x498 &  x526 & ~x0 & ~x26 & ~x27 & ~x55 & ~x308 & ~x337 & ~x364 & ~x420 & ~x588 & ~x777;
assign c80 =  x329 & ~x1 & ~x21 & ~x137 & ~x298 & ~x389 & ~x390 & ~x391 & ~x436 & ~x437 & ~x491 & ~x520;
assign c82 =  x213 &  x241 &  x269 &  x297 &  x409 & ~x2 & ~x26 & ~x28 & ~x31 & ~x52 & ~x53 & ~x54 & ~x55 & ~x60 & ~x77 & ~x80 & ~x83 & ~x84 & ~x85 & ~x105 & ~x106 & ~x107 & ~x108 & ~x133 & ~x134 & ~x139 & ~x168 & ~x171 & ~x190 & ~x192 & ~x197 & ~x198 & ~x222 & ~x224 & ~x246 & ~x250 & ~x251 & ~x275 & ~x277 & ~x302 & ~x303 & ~x330 & ~x359 & ~x366 & ~x660 & ~x757;
assign c84 =  x739 &  x744 & ~x8 & ~x36 & ~x178 & ~x218 & ~x261 & ~x288 & ~x317 & ~x367 & ~x400 & ~x580 & ~x660;
assign c86 =  x488 & ~x23 & ~x50 & ~x52 & ~x53 & ~x59 & ~x63 & ~x86 & ~x91 & ~x116 & ~x118 & ~x143 & ~x145 & ~x148 & ~x161 & ~x162 & ~x164 & ~x170 & ~x174 & ~x176 & ~x193 & ~x198 & ~x202 & ~x217 & ~x252 & ~x257 & ~x284 & ~x308 & ~x310 & ~x317 & ~x337 & ~x340 & ~x364 & ~x427 & ~x456 & ~x474 & ~x479 & ~x481 & ~x502 & ~x531 & ~x533 & ~x551 & ~x555 & ~x562 & ~x563 & ~x578 & ~x579 & ~x584 & ~x670 & ~x697 & ~x725 & ~x729 & ~x730;
assign c88 =  x377 & ~x4 & ~x5 & ~x60 & ~x82 & ~x113 & ~x114 & ~x117 & ~x136 & ~x147 & ~x174 & ~x251 & ~x303 & ~x308 & ~x311 & ~x334 & ~x339 & ~x340 & ~x365 & ~x416 & ~x420 & ~x426 & ~x454 & ~x467 & ~x474 & ~x477 & ~x478 & ~x498 & ~x521 & ~x522 & ~x549 & ~x551 & ~x555 & ~x562 & ~x629 & ~x641 & ~x645 & ~x672 & ~x696 & ~x753 & ~x757;
assign c810 = ~x17 & ~x18 & ~x20 & ~x22 & ~x28 & ~x54 & ~x61 & ~x80 & ~x86 & ~x115 & ~x136 & ~x141 & ~x143 & ~x166 & ~x172 & ~x193 & ~x198 & ~x251 & ~x252 & ~x254 & ~x281 & ~x305 & ~x334 & ~x389 & ~x391 & ~x408 & ~x444 & ~x445 & ~x449 & ~x464 & ~x492 & ~x519 & ~x520 & ~x549 & ~x693 & ~x719 & ~x738 & ~x757 & ~x759 & ~x772 & ~x783;
assign c812 =  x406 & ~x1 & ~x3 & ~x8 & ~x28 & ~x29 & ~x34 & ~x35 & ~x48 & ~x53 & ~x55 & ~x56 & ~x58 & ~x60 & ~x80 & ~x83 & ~x85 & ~x87 & ~x90 & ~x107 & ~x108 & ~x116 & ~x117 & ~x137 & ~x140 & ~x141 & ~x146 & ~x163 & ~x166 & ~x167 & ~x169 & ~x170 & ~x172 & ~x174 & ~x190 & ~x194 & ~x200 & ~x221 & ~x224 & ~x225 & ~x226 & ~x249 & ~x254 & ~x257 & ~x258 & ~x278 & ~x281 & ~x283 & ~x285 & ~x305 & ~x306 & ~x307 & ~x308 & ~x310 & ~x332 & ~x334 & ~x336 & ~x338 & ~x339 & ~x361 & ~x364 & ~x365 & ~x367 & ~x387 & ~x388 & ~x389 & ~x392 & ~x393 & ~x394 & ~x396 & ~x397 & ~x398 & ~x419 & ~x423 & ~x424 & ~x425 & ~x444 & ~x445 & ~x446 & ~x447 & ~x448 & ~x449 & ~x476 & ~x478 & ~x480 & ~x498 & ~x500 & ~x505 & ~x523 & ~x524 & ~x528 & ~x550 & ~x556 & ~x558 & ~x576 & ~x577 & ~x586 & ~x587 & ~x588 & ~x601 & ~x603 & ~x613 & ~x615 & ~x643 & ~x645 & ~x671 & ~x672 & ~x724 & ~x727 & ~x729 & ~x753 & ~x782;
assign c814 =  x738 & ~x58 & ~x109 & ~x164 & ~x219 & ~x247 & ~x333 & ~x364 & ~x414 & ~x415 & ~x441 & ~x444 & ~x449 & ~x502 & ~x606 & ~x607 & ~x633 & ~x655 & ~x683 & ~x782;
assign c816 = ~x3 & ~x6 & ~x49 & ~x77 & ~x85 & ~x100 & ~x103 & ~x156 & ~x170 & ~x228 & ~x251 & ~x296 & ~x297 & ~x314 & ~x335 & ~x339 & ~x354 & ~x382 & ~x474 & ~x476 & ~x532 & ~x550 & ~x551;
assign c818 =  x589 & ~x1 & ~x29 & ~x83 & ~x111 & ~x138 & ~x139 & ~x166 & ~x195 & ~x222 & ~x251 & ~x363 & ~x446 & ~x447 & ~x477 & ~x515;
assign c820 = ~x47 & ~x53 & ~x65 & ~x82 & ~x108 & ~x126 & ~x132 & ~x194 & ~x332 & ~x334 & ~x483 & ~x651 & ~x706 & ~x724 & ~x776;
assign c822 =  x463 &  x488 &  x717 & ~x498 & ~x554;
assign c824 =  x508 & ~x18 & ~x30 & ~x44 & ~x46 & ~x50 & ~x53 & ~x75 & ~x78 & ~x85 & ~x112 & ~x113 & ~x137 & ~x220 & ~x222 & ~x276 & ~x277 & ~x388 & ~x390 & ~x416 & ~x420 & ~x559 & ~x585;
assign c826 = ~x81 & ~x101 & ~x112 & ~x113 & ~x114 & ~x167 & ~x171 & ~x194 & ~x196 & ~x205 & ~x225 & ~x253 & ~x305 & ~x307 & ~x390 & ~x393 & ~x491 & ~x689 & ~x729 & ~x758;
assign c828 = ~x1 & ~x3 & ~x21 & ~x26 & ~x27 & ~x29 & ~x30 & ~x53 & ~x54 & ~x77 & ~x81 & ~x83 & ~x85 & ~x109 & ~x112 & ~x113 & ~x132 & ~x133 & ~x137 & ~x141 & ~x143 & ~x161 & ~x167 & ~x168 & ~x169 & ~x189 & ~x194 & ~x197 & ~x198 & ~x222 & ~x223 & ~x245 & ~x250 & ~x251 & ~x273 & ~x274 & ~x275 & ~x280 & ~x282 & ~x300 & ~x303 & ~x305 & ~x306 & ~x309 & ~x328 & ~x331 & ~x336 & ~x357 & ~x363 & ~x364 & ~x366 & ~x386 & ~x387 & ~x390 & ~x391 & ~x392 & ~x393 & ~x395 & ~x412 & ~x413 & ~x416 & ~x423 & ~x445 & ~x446 & ~x449 & ~x469 & ~x470 & ~x472 & ~x474 & ~x496 & ~x497 & ~x500 & ~x501 & ~x524 & ~x525 & ~x526 & ~x528 & ~x529 & ~x556 & ~x580 & ~x583 & ~x584 & ~x587 & ~x629 & ~x630 & ~x655 & ~x671 & ~x757 & ~x782 & ~x783;
assign c830 =  x374 & ~x1 & ~x26 & ~x45 & ~x46 & ~x82 & ~x84 & ~x85 & ~x89 & ~x142 & ~x167 & ~x170 & ~x171 & ~x196 & ~x226 & ~x252 & ~x309 & ~x336 & ~x362 & ~x363 & ~x419 & ~x422 & ~x447 & ~x474 & ~x475 & ~x493 & ~x548 & ~x549 & ~x574 & ~x575 & ~x755 & ~x777 & ~x778 & ~x783;
assign c832 = ~x23 & ~x24 & ~x42 & ~x50 & ~x139 & ~x166 & ~x219 & ~x220 & ~x222 & ~x249 & ~x250 & ~x277 & ~x331 & ~x359 & ~x387 & ~x388 & ~x457 & ~x596 & ~x730 & ~x735 & ~x743;
assign c834 =  x509 &  x562 &  x622 & ~x80 & ~x137 & ~x365;
assign c836 =  x594 &  x645 & ~x167 & ~x171 & ~x449 & ~x477;
assign c838 =  x450 & ~x277 & ~x360 & ~x401 & ~x429 & ~x486 & ~x707;
assign c840 = ~x1 & ~x25 & ~x28 & ~x55 & ~x56 & ~x57 & ~x77 & ~x80 & ~x83 & ~x84 & ~x87 & ~x108 & ~x110 & ~x111 & ~x114 & ~x131 & ~x137 & ~x139 & ~x140 & ~x142 & ~x143 & ~x161 & ~x165 & ~x166 & ~x195 & ~x197 & ~x198 & ~x216 & ~x217 & ~x221 & ~x224 & ~x245 & ~x248 & ~x249 & ~x250 & ~x275 & ~x303 & ~x307 & ~x332 & ~x334 & ~x335 & ~x336 & ~x337 & ~x359 & ~x363 & ~x392 & ~x395 & ~x413 & ~x414 & ~x415 & ~x441 & ~x446 & ~x447 & ~x468 & ~x469 & ~x470 & ~x471 & ~x472 & ~x474 & ~x496 & ~x500 & ~x504 & ~x528 & ~x559 & ~x579 & ~x583 & ~x584 & ~x588 & ~x605 & ~x611 & ~x616 & ~x627 & ~x628 & ~x631 & ~x669 & ~x672 & ~x700 & ~x728;
assign c842 =  x372 &  x400 &  x540 &  x568 &  x596 & ~x4 & ~x24 & ~x25 & ~x26 & ~x28 & ~x29 & ~x31 & ~x53 & ~x56 & ~x57 & ~x82 & ~x87 & ~x111 & ~x112 & ~x114 & ~x138 & ~x139 & ~x140 & ~x145 & ~x168 & ~x281 & ~x366 & ~x391 & ~x392 & ~x394 & ~x419 & ~x422 & ~x476 & ~x490 & ~x515 & ~x516 & ~x518 & ~x545 & ~x599 & ~x601 & ~x732;
assign c844 = ~x0 & ~x2 & ~x4 & ~x21 & ~x22 & ~x27 & ~x32 & ~x48 & ~x53 & ~x57 & ~x77 & ~x88 & ~x108 & ~x113 & ~x114 & ~x115 & ~x136 & ~x137 & ~x141 & ~x167 & ~x195 & ~x196 & ~x201 & ~x221 & ~x229 & ~x256 & ~x277 & ~x281 & ~x286 & ~x304 & ~x308 & ~x312 & ~x333 & ~x334 & ~x335 & ~x337 & ~x340 & ~x341 & ~x362 & ~x367 & ~x383 & ~x392 & ~x398 & ~x416 & ~x417 & ~x420 & ~x444 & ~x445 & ~x448 & ~x449 & ~x578 & ~x605 & ~x607 & ~x631 & ~x632 & ~x634 & ~x635 & ~x656 & ~x657 & ~x697 & ~x755;
assign c846 =  x573 &  x739 &  x740 &  x742 & ~x243 & ~x454 & ~x509 & ~x538 & ~x593;
assign c848 =  x768 & ~x190 & ~x357 & ~x385 & ~x391 & ~x469 & ~x583 & ~x661 & ~x683 & ~x686;
assign c850 =  x374 &  x430 &  x597 & ~x4 & ~x32 & ~x56 & ~x61 & ~x85 & ~x118 & ~x119 & ~x175 & ~x196 & ~x228 & ~x229 & ~x252 & ~x255 & ~x256 & ~x257 & ~x258 & ~x285 & ~x309 & ~x365 & ~x391 & ~x393 & ~x418 & ~x420 & ~x421 & ~x424 & ~x453 & ~x475 & ~x531;
assign c852 = ~x32 & ~x55 & ~x56 & ~x57 & ~x73 & ~x85 & ~x88 & ~x89 & ~x110 & ~x111 & ~x140 & ~x144 & ~x167 & ~x170 & ~x174 & ~x195 & ~x199 & ~x215 & ~x222 & ~x228 & ~x256 & ~x257 & ~x279 & ~x281 & ~x282 & ~x286 & ~x306 & ~x307 & ~x308 & ~x310 & ~x312 & ~x314 & ~x327 & ~x335 & ~x337 & ~x340 & ~x342 & ~x365 & ~x367 & ~x382 & ~x383 & ~x394 & ~x395 & ~x397 & ~x423 & ~x426 & ~x438 & ~x450 & ~x452 & ~x467 & ~x478 & ~x522 & ~x616 & ~x691 & ~x698 & ~x699 & ~x713 & ~x734 & ~x754 & ~x756 & ~x783;
assign c854 = ~x0 & ~x1 & ~x10 & ~x19 & ~x22 & ~x26 & ~x45 & ~x52 & ~x55 & ~x73 & ~x75 & ~x79 & ~x81 & ~x82 & ~x102 & ~x106 & ~x132 & ~x139 & ~x140 & ~x162 & ~x165 & ~x190 & ~x192 & ~x194 & ~x277 & ~x303 & ~x330 & ~x332 & ~x333 & ~x358 & ~x361 & ~x387 & ~x391 & ~x489 & ~x517 & ~x641 & ~x642 & ~x643 & ~x732 & ~x743 & ~x744 & ~x768 & ~x772;
assign c856 =  x734 & ~x2 & ~x28 & ~x53 & ~x54 & ~x56 & ~x58 & ~x84 & ~x110 & ~x112 & ~x114 & ~x138 & ~x139 & ~x140 & ~x141 & ~x142 & ~x168 & ~x394 & ~x395 & ~x421 & ~x449 & ~x477 & ~x583 & ~x584 & ~x587 & ~x653 & ~x671;
assign c858 =  x512 & ~x1 & ~x23 & ~x24 & ~x27 & ~x28 & ~x30 & ~x51 & ~x81 & ~x84 & ~x88 & ~x109 & ~x111 & ~x115 & ~x117 & ~x135 & ~x139 & ~x140 & ~x141 & ~x144 & ~x170 & ~x193 & ~x194 & ~x223 & ~x247 & ~x276 & ~x277 & ~x336 & ~x387 & ~x418 & ~x420 & ~x422 & ~x423 & ~x480 & ~x529 & ~x532 & ~x534 & ~x559 & ~x629 & ~x630 & ~x656 & ~x670 & ~x684 & ~x729 & ~x755 & ~x782;
assign c860 =  x432 & ~x6 & ~x8 & ~x20 & ~x25 & ~x27 & ~x32 & ~x34 & ~x37 & ~x40 & ~x52 & ~x53 & ~x55 & ~x61 & ~x63 & ~x80 & ~x81 & ~x88 & ~x89 & ~x90 & ~x107 & ~x108 & ~x119 & ~x136 & ~x149 & ~x171 & ~x173 & ~x175 & ~x197 & ~x201 & ~x202 & ~x217 & ~x222 & ~x224 & ~x228 & ~x229 & ~x248 & ~x253 & ~x256 & ~x257 & ~x280 & ~x284 & ~x288 & ~x334 & ~x337 & ~x362 & ~x393 & ~x394 & ~x395 & ~x419 & ~x421 & ~x422 & ~x424 & ~x427 & ~x444 & ~x445 & ~x449 & ~x450 & ~x474 & ~x475 & ~x523 & ~x531 & ~x533 & ~x558 & ~x616 & ~x699 & ~x700 & ~x755 & ~x760;
assign c862 =  x72 &  x128 &  x156 &  x184 &  x212 &  x240 &  x268 & ~x2 & ~x6 & ~x55 & ~x89 & ~x159 & ~x160 & ~x162 & ~x215 & ~x244 & ~x275 & ~x358 & ~x394 & ~x397 & ~x449 & ~x527 & ~x553 & ~x554 & ~x775;
assign c864 =  x247 &  x331 & ~x437 & ~x721;
assign c866 =  x593 &  x706 & ~x22 & ~x23 & ~x25 & ~x27 & ~x84 & ~x85 & ~x141 & ~x142 & ~x169 & ~x171 & ~x198 & ~x226 & ~x280 & ~x336 & ~x625;
assign c868 =  x266 &  x350 &  x378 &  x434 &  x462 & ~x130 & ~x132 & ~x171 & ~x214 & ~x215 & ~x311 & ~x355 & ~x357 & ~x384 & ~x385 & ~x398 & ~x426 & ~x441 & ~x525;
assign c870 = ~x1 & ~x6 & ~x7 & ~x19 & ~x20 & ~x24 & ~x27 & ~x32 & ~x53 & ~x55 & ~x57 & ~x59 & ~x61 & ~x83 & ~x88 & ~x110 & ~x111 & ~x112 & ~x114 & ~x115 & ~x139 & ~x141 & ~x143 & ~x167 & ~x195 & ~x197 & ~x223 & ~x253 & ~x254 & ~x282 & ~x306 & ~x307 & ~x309 & ~x336 & ~x338 & ~x367 & ~x391 & ~x393 & ~x395 & ~x418 & ~x437 & ~x448 & ~x450 & ~x464 & ~x465 & ~x476 & ~x477 & ~x491 & ~x494 & ~x505 & ~x518 & ~x532 & ~x546 & ~x559 & ~x746 & ~x772;
assign c872 = ~x6 & ~x20 & ~x24 & ~x39 & ~x51 & ~x105 & ~x132 & ~x134 & ~x137 & ~x163 & ~x188 & ~x189 & ~x216 & ~x224 & ~x248 & ~x251 & ~x274 & ~x275 & ~x333 & ~x357 & ~x360 & ~x385 & ~x695 & ~x705 & ~x710 & ~x720 & ~x725 & ~x726 & ~x732 & ~x739 & ~x743 & ~x744 & ~x750 & ~x754 & ~x761;
assign c874 =  x429 &  x457 &  x485 &  x653 & ~x26 & ~x29 & ~x58 & ~x60 & ~x88 & ~x110 & ~x138 & ~x140 & ~x196 & ~x280 & ~x335 & ~x392 & ~x517 & ~x545 & ~x548 & ~x744;
assign c876 =  x301 & ~x33 & ~x57 & ~x59 & ~x83 & ~x85 & ~x249 & ~x270 & ~x279 & ~x281 & ~x324 & ~x335 & ~x409 & ~x492 & ~x522;
assign c878 =  x350 &  x489 & ~x25 & ~x84 & ~x163 & ~x164 & ~x166 & ~x192 & ~x198 & ~x219 & ~x221 & ~x226 & ~x246 & ~x247 & ~x249 & ~x276 & ~x278 & ~x301 & ~x304 & ~x331 & ~x389 & ~x391 & ~x395 & ~x441 & ~x444 & ~x445 & ~x451 & ~x471 & ~x499 & ~x532 & ~x551 & ~x555 & ~x556 & ~x578 & ~x580 & ~x627;
assign c880 =  x351 &  x379 &  x435 &  x463 &  x490 &  x517 & ~x0 & ~x23 & ~x28 & ~x51 & ~x52 & ~x55 & ~x79 & ~x80 & ~x84 & ~x111 & ~x112 & ~x113 & ~x114 & ~x132 & ~x137 & ~x160 & ~x163 & ~x164 & ~x189 & ~x190 & ~x193 & ~x197 & ~x199 & ~x218 & ~x219 & ~x220 & ~x223 & ~x224 & ~x245 & ~x247 & ~x248 & ~x250 & ~x255 & ~x274 & ~x277 & ~x281 & ~x301 & ~x308 & ~x309 & ~x311 & ~x337 & ~x359 & ~x368 & ~x387 & ~x390 & ~x391 & ~x393 & ~x394 & ~x414 & ~x416 & ~x420 & ~x442 & ~x443 & ~x445 & ~x450 & ~x452 & ~x454 & ~x468 & ~x471 & ~x478 & ~x480 & ~x482 & ~x497 & ~x498 & ~x505 & ~x507 & ~x524 & ~x527 & ~x530 & ~x533 & ~x534 & ~x551 & ~x553 & ~x555 & ~x581 & ~x588 & ~x614 & ~x615 & ~x669 & ~x673 & ~x697 & ~x725 & ~x728;
assign c882 =  x296 &  x324 & ~x1 & ~x50 & ~x55 & ~x108 & ~x137 & ~x140 & ~x160 & ~x193 & ~x246 & ~x247 & ~x273 & ~x302 & ~x331 & ~x332 & ~x333 & ~x334 & ~x364 & ~x473 & ~x503 & ~x526 & ~x527 & ~x528 & ~x552 & ~x553 & ~x659 & ~x684;
assign c884 = ~x2 & ~x21 & ~x24 & ~x25 & ~x26 & ~x27 & ~x29 & ~x51 & ~x53 & ~x77 & ~x78 & ~x79 & ~x81 & ~x85 & ~x103 & ~x104 & ~x105 & ~x107 & ~x109 & ~x111 & ~x112 & ~x132 & ~x134 & ~x135 & ~x137 & ~x162 & ~x163 & ~x167 & ~x190 & ~x193 & ~x194 & ~x196 & ~x216 & ~x222 & ~x223 & ~x244 & ~x247 & ~x249 & ~x277 & ~x279 & ~x300 & ~x302 & ~x308 & ~x329 & ~x332 & ~x333 & ~x337 & ~x356 & ~x359 & ~x363 & ~x383 & ~x385 & ~x392 & ~x445 & ~x471 & ~x627 & ~x729 & ~x758 & ~x770 & ~x780;
assign c886 =  x240 &  x268 &  x348 &  x625 & ~x117 & ~x173 & ~x777;
assign c888 =  x717 & ~x78 & ~x120 & ~x137 & ~x147 & ~x164 & ~x169 & ~x191 & ~x205 & ~x219 & ~x221 & ~x232 & ~x256 & ~x289 & ~x310 & ~x316 & ~x339 & ~x392 & ~x422 & ~x428 & ~x442 & ~x455 & ~x527 & ~x529 & ~x578 & ~x579 & ~x778;
assign c890 = ~x0 & ~x1 & ~x4 & ~x8 & ~x23 & ~x24 & ~x27 & ~x30 & ~x53 & ~x58 & ~x61 & ~x64 & ~x82 & ~x83 & ~x85 & ~x112 & ~x114 & ~x115 & ~x117 & ~x137 & ~x138 & ~x141 & ~x142 & ~x170 & ~x175 & ~x194 & ~x195 & ~x196 & ~x199 & ~x200 & ~x204 & ~x223 & ~x228 & ~x251 & ~x278 & ~x279 & ~x283 & ~x306 & ~x307 & ~x336 & ~x362 & ~x363 & ~x391 & ~x464 & ~x473 & ~x476 & ~x491 & ~x519 & ~x547 & ~x575 & ~x576 & ~x715 & ~x741 & ~x768 & ~x769;
assign c892 =  x457 & ~x3 & ~x28 & ~x37 & ~x54 & ~x82 & ~x84 & ~x85 & ~x87 & ~x89 & ~x109 & ~x113 & ~x116 & ~x117 & ~x139 & ~x144 & ~x146 & ~x147 & ~x167 & ~x173 & ~x174 & ~x175 & ~x200 & ~x202 & ~x228 & ~x229 & ~x251 & ~x252 & ~x257 & ~x259 & ~x283 & ~x286 & ~x312 & ~x338 & ~x391 & ~x419 & ~x421 & ~x448 & ~x476 & ~x549 & ~x560 & ~x712;
assign c894 =  x179 &  x379 &  x486 & ~x230 & ~x259 & ~x282 & ~x341 & ~x364 & ~x476;
assign c896 =  x377 & ~x86 & ~x248 & ~x330 & ~x364 & ~x372 & ~x397 & ~x466 & ~x473 & ~x574 & ~x600;
assign c898 =  x507 & ~x3 & ~x80 & ~x110 & ~x118 & ~x136 & ~x278 & ~x305 & ~x324 & ~x334 & ~x335 & ~x360 & ~x361 & ~x388;
assign c8100 =  x492 &  x547 & ~x91 & ~x173 & ~x174 & ~x427 & ~x454 & ~x471 & ~x510 & ~x535 & ~x552 & ~x583 & ~x606;
assign c8102 =  x212 &  x296 &  x348 &  x380 & ~x0 & ~x52 & ~x58 & ~x134 & ~x135 & ~x140 & ~x162 & ~x166 & ~x168 & ~x191 & ~x194 & ~x220 & ~x250 & ~x251 & ~x304 & ~x309 & ~x334 & ~x386 & ~x390 & ~x395 & ~x418 & ~x421 & ~x451 & ~x469 & ~x476 & ~x530 & ~x556 & ~x581 & ~x582 & ~x583 & ~x588 & ~x756 & ~x782;
assign c8104 =  x373 & ~x3 & ~x4 & ~x22 & ~x25 & ~x28 & ~x49 & ~x50 & ~x55 & ~x56 & ~x60 & ~x86 & ~x88 & ~x110 & ~x112 & ~x114 & ~x115 & ~x138 & ~x140 & ~x141 & ~x143 & ~x144 & ~x166 & ~x168 & ~x169 & ~x174 & ~x196 & ~x202 & ~x223 & ~x224 & ~x251 & ~x253 & ~x279 & ~x334 & ~x335 & ~x363 & ~x364 & ~x365 & ~x366 & ~x390 & ~x392 & ~x394 & ~x395 & ~x396 & ~x420 & ~x422 & ~x449 & ~x451 & ~x476 & ~x477 & ~x478 & ~x502 & ~x504 & ~x506 & ~x532 & ~x558 & ~x559 & ~x576 & ~x603 & ~x604 & ~x615 & ~x628 & ~x630 & ~x631 & ~x632 & ~x727 & ~x729 & ~x753 & ~x754 & ~x779;
assign c8106 = ~x1 & ~x4 & ~x8 & ~x19 & ~x23 & ~x28 & ~x61 & ~x74 & ~x91 & ~x116 & ~x143 & ~x171 & ~x195 & ~x198 & ~x250 & ~x305 & ~x326 & ~x333 & ~x353 & ~x362 & ~x417 & ~x419 & ~x464 & ~x466 & ~x501 & ~x502 & ~x503 & ~x521 & ~x522 & ~x549 & ~x747;
assign c8108 = ~x1 & ~x16 & ~x43 & ~x53 & ~x78 & ~x81 & ~x105 & ~x106 & ~x109 & ~x133 & ~x136 & ~x138 & ~x161 & ~x164 & ~x189 & ~x192 & ~x218 & ~x219 & ~x226 & ~x246 & ~x250 & ~x273 & ~x276 & ~x303 & ~x304 & ~x305 & ~x307 & ~x329 & ~x331 & ~x332 & ~x357 & ~x358 & ~x385 & ~x403 & ~x657 & ~x738 & ~x762 & ~x765 & ~x766;
assign c8110 =  x469 & ~x22 & ~x85 & ~x167 & ~x173 & ~x281 & ~x334 & ~x338 & ~x354 & ~x435 & ~x437 & ~x491 & ~x521;
assign c8112 =  x427 & ~x2 & ~x25 & ~x33 & ~x34 & ~x55 & ~x60 & ~x62 & ~x83 & ~x85 & ~x110 & ~x115 & ~x116 & ~x118 & ~x140 & ~x142 & ~x166 & ~x169 & ~x172 & ~x196 & ~x198 & ~x199 & ~x223 & ~x225 & ~x226 & ~x279 & ~x337 & ~x351 & ~x363 & ~x377 & ~x379 & ~x391 & ~x405 & ~x421 & ~x433 & ~x460 & ~x461 & ~x463 & ~x488 & ~x517 & ~x544 & ~x545;
assign c8114 = ~x1 & ~x2 & ~x3 & ~x4 & ~x6 & ~x23 & ~x24 & ~x25 & ~x26 & ~x27 & ~x28 & ~x29 & ~x30 & ~x31 & ~x32 & ~x33 & ~x34 & ~x53 & ~x56 & ~x57 & ~x58 & ~x60 & ~x61 & ~x62 & ~x79 & ~x80 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x88 & ~x90 & ~x109 & ~x110 & ~x111 & ~x112 & ~x113 & ~x115 & ~x116 & ~x118 & ~x137 & ~x139 & ~x140 & ~x146 & ~x165 & ~x166 & ~x167 & ~x168 & ~x169 & ~x170 & ~x172 & ~x173 & ~x175 & ~x193 & ~x194 & ~x195 & ~x196 & ~x198 & ~x199 & ~x200 & ~x201 & ~x221 & ~x224 & ~x225 & ~x229 & ~x230 & ~x251 & ~x252 & ~x253 & ~x254 & ~x255 & ~x256 & ~x257 & ~x258 & ~x278 & ~x279 & ~x280 & ~x281 & ~x282 & ~x283 & ~x284 & ~x285 & ~x286 & ~x308 & ~x309 & ~x310 & ~x311 & ~x312 & ~x314 & ~x334 & ~x337 & ~x338 & ~x339 & ~x340 & ~x341 & ~x361 & ~x362 & ~x364 & ~x365 & ~x366 & ~x367 & ~x369 & ~x390 & ~x391 & ~x392 & ~x393 & ~x395 & ~x396 & ~x397 & ~x417 & ~x418 & ~x419 & ~x420 & ~x423 & ~x425 & ~x447 & ~x448 & ~x449 & ~x450 & ~x451 & ~x466 & ~x475 & ~x476 & ~x478 & ~x479 & ~x495 & ~x504 & ~x506 & ~x521 & ~x522 & ~x523 & ~x548 & ~x549 & ~x550 & ~x551 & ~x552 & ~x559 & ~x575 & ~x578 & ~x601 & ~x602 & ~x616 & ~x669 & ~x672 & ~x699 & ~x703 & ~x704 & ~x724 & ~x726 & ~x727 & ~x728 & ~x730 & ~x731 & ~x732 & ~x752 & ~x754 & ~x755 & ~x757 & ~x758 & ~x760 & ~x763 & ~x765 & ~x778 & ~x780 & ~x782 & ~x783;
assign c8116 =  x510 &  x618 &  x706 & ~x365;
assign c8118 =  x520 & ~x342 & ~x454 & ~x581 & ~x605 & ~x607;
assign c8120 =  x185 & ~x3 & ~x4 & ~x118 & ~x166 & ~x364 & ~x365 & ~x396 & ~x450 & ~x465 & ~x477 & ~x547 & ~x548 & ~x572 & ~x573 & ~x778;
assign c8122 =  x748 & ~x77 & ~x107 & ~x114 & ~x115 & ~x163 & ~x188 & ~x218 & ~x246 & ~x423 & ~x630 & ~x654 & ~x655 & ~x656;
assign c8124 =  x302 & ~x33 & ~x54 & ~x57 & ~x61 & ~x84 & ~x86 & ~x89 & ~x197 & ~x391 & ~x417 & ~x465 & ~x519 & ~x522 & ~x749;
assign c8126 =  x735 & ~x255 & ~x422 & ~x424 & ~x452 & ~x560 & ~x629;
assign c8128 = ~x5 & ~x6 & ~x21 & ~x32 & ~x35 & ~x57 & ~x60 & ~x82 & ~x86 & ~x118 & ~x119 & ~x137 & ~x141 & ~x147 & ~x173 & ~x201 & ~x230 & ~x250 & ~x255 & ~x256 & ~x281 & ~x283 & ~x308 & ~x309 & ~x310 & ~x312 & ~x336 & ~x337 & ~x340 & ~x341 & ~x365 & ~x370 & ~x382 & ~x391 & ~x409 & ~x437 & ~x447 & ~x449 & ~x452 & ~x476 & ~x492 & ~x493 & ~x494 & ~x519 & ~x521 & ~x546 & ~x615 & ~x719 & ~x720;
assign c8130 =  x127 &  x155 &  x183 &  x239 &  x267 &  x295 &  x323 &  x351 &  x435 & ~x109 & ~x136 & ~x141 & ~x157 & ~x158 & ~x161 & ~x188 & ~x214 & ~x303 & ~x328 & ~x332 & ~x357 & ~x414 & ~x417 & ~x468 & ~x614;
assign c8132 =  x484 & ~x25 & ~x28 & ~x29 & ~x54 & ~x57 & ~x59 & ~x61 & ~x62 & ~x83 & ~x84 & ~x86 & ~x87 & ~x88 & ~x89 & ~x109 & ~x110 & ~x111 & ~x112 & ~x114 & ~x115 & ~x138 & ~x141 & ~x143 & ~x145 & ~x170 & ~x171 & ~x195 & ~x222 & ~x226 & ~x252 & ~x256 & ~x257 & ~x277 & ~x285 & ~x305 & ~x307 & ~x308 & ~x334 & ~x340 & ~x341 & ~x362 & ~x363 & ~x365 & ~x368 & ~x369 & ~x389 & ~x393 & ~x394 & ~x419 & ~x423 & ~x424 & ~x450 & ~x452 & ~x476 & ~x477 & ~x520 & ~x531 & ~x532 & ~x614 & ~x615 & ~x671 & ~x711 & ~x724 & ~x727 & ~x783;
assign c8134 =  x588 & ~x702;
assign c8136 =  x519 &  x745 & ~x97 & ~x556 & ~x605 & ~x606;
assign c8138 =  x347 & ~x3 & ~x5 & ~x54 & ~x63 & ~x65 & ~x73 & ~x88 & ~x109 & ~x113 & ~x140 & ~x171 & ~x204 & ~x223 & ~x227 & ~x230 & ~x231 & ~x256 & ~x260 & ~x282 & ~x310 & ~x339 & ~x344 & ~x372 & ~x467 & ~x522 & ~x523;
assign c8140 =  x455 &  x539 &  x595 &  x679 & ~x3 & ~x27 & ~x31 & ~x54 & ~x57 & ~x83 & ~x87 & ~x110 & ~x113 & ~x116 & ~x137 & ~x138 & ~x141 & ~x143 & ~x198 & ~x225 & ~x251 & ~x252 & ~x279 & ~x335 & ~x336 & ~x598 & ~x599 & ~x600 & ~x710 & ~x758 & ~x760;
assign c8142 =  x689 & ~x3 & ~x25 & ~x53 & ~x58 & ~x118 & ~x148 & ~x149 & ~x160 & ~x169 & ~x191 & ~x286 & ~x417 & ~x424 & ~x427 & ~x580 & ~x606 & ~x613 & ~x632 & ~x731 & ~x758 & ~x776;
assign c8144 = ~x0 & ~x1 & ~x21 & ~x29 & ~x30 & ~x52 & ~x56 & ~x80 & ~x84 & ~x86 & ~x87 & ~x89 & ~x102 & ~x109 & ~x111 & ~x113 & ~x115 & ~x116 & ~x127 & ~x138 & ~x140 & ~x141 & ~x165 & ~x170 & ~x172 & ~x193 & ~x197 & ~x249 & ~x250 & ~x251 & ~x269 & ~x297 & ~x307 & ~x309 & ~x336 & ~x337 & ~x339 & ~x353 & ~x363 & ~x366 & ~x389 & ~x391 & ~x392 & ~x409 & ~x437 & ~x445 & ~x446 & ~x493 & ~x548 & ~x576;
assign c8146 =  x737 & ~x85 & ~x118 & ~x168 & ~x199 & ~x223 & ~x281 & ~x336 & ~x386 & ~x424 & ~x443 & ~x497 & ~x605 & ~x655 & ~x656 & ~x657 & ~x781;
assign c8148 =  x563 & ~x0 & ~x1 & ~x2 & ~x6 & ~x18 & ~x22 & ~x30 & ~x46 & ~x50 & ~x52 & ~x53 & ~x83 & ~x109 & ~x110 & ~x113 & ~x115 & ~x116 & ~x196 & ~x225 & ~x250 & ~x251 & ~x252 & ~x306 & ~x311 & ~x351 & ~x361 & ~x362 & ~x363 & ~x388 & ~x391 & ~x393 & ~x394 & ~x422 & ~x518 & ~x757;
assign c8150 = ~x79 & ~x107 & ~x135 & ~x138 & ~x157 & ~x165 & ~x170 & ~x198 & ~x220 & ~x242 & ~x270 & ~x297 & ~x325 & ~x333 & ~x354 & ~x362 & ~x409 & ~x447 & ~x493 & ~x718;
assign c8152 =  x690 & ~x161 & ~x189 & ~x413 & ~x553 & ~x578 & ~x629 & ~x630;
assign c8154 =  x434 &  x741 & ~x328 & ~x355 & ~x412 & ~x532 & ~x607 & ~x659 & ~x686;
assign c8156 =  x246 &  x510 & ~x29 & ~x89 & ~x436 & ~x492 & ~x749;
assign c8158 =  x210 &  x267 &  x323 & ~x131 & ~x186 & ~x191 & ~x214 & ~x215 & ~x219 & ~x242 & ~x326 & ~x333 & ~x384 & ~x411 & ~x412 & ~x502;
assign c8160 =  x213 & ~x23 & ~x51 & ~x53 & ~x56 & ~x58 & ~x88 & ~x105 & ~x106 & ~x139 & ~x165 & ~x168 & ~x188 & ~x191 & ~x194 & ~x197 & ~x199 & ~x226 & ~x245 & ~x247 & ~x274 & ~x276 & ~x278 & ~x335 & ~x364 & ~x447 & ~x502 & ~x530 & ~x555 & ~x574 & ~x575 & ~x576;
assign c8162 = ~x15 & ~x18 & ~x19 & ~x26 & ~x28 & ~x29 & ~x30 & ~x31 & ~x43 & ~x45 & ~x50 & ~x53 & ~x72 & ~x77 & ~x78 & ~x102 & ~x103 & ~x104 & ~x105 & ~x106 & ~x107 & ~x108 & ~x115 & ~x129 & ~x130 & ~x131 & ~x132 & ~x134 & ~x136 & ~x137 & ~x139 & ~x158 & ~x159 & ~x167 & ~x170 & ~x171 & ~x189 & ~x191 & ~x192 & ~x216 & ~x217 & ~x219 & ~x220 & ~x221 & ~x244 & ~x246 & ~x248 & ~x249 & ~x251 & ~x271 & ~x272 & ~x273 & ~x276 & ~x278 & ~x279 & ~x300 & ~x303 & ~x305 & ~x329 & ~x330 & ~x331 & ~x332 & ~x357 & ~x358 & ~x359 & ~x362 & ~x363 & ~x384 & ~x387 & ~x388 & ~x389 & ~x390 & ~x412 & ~x414 & ~x415 & ~x416 & ~x417 & ~x440 & ~x442 & ~x443 & ~x476 & ~x584 & ~x585 & ~x616 & ~x726 & ~x758 & ~x783;
assign c8164 = ~x24 & ~x47 & ~x57 & ~x101 & ~x159 & ~x171 & ~x219 & ~x220 & ~x275 & ~x299 & ~x361 & ~x415 & ~x439 & ~x466 & ~x531 & ~x712 & ~x728;
assign c8166 =  x296 & ~x110 & ~x163 & ~x191 & ~x221 & ~x223 & ~x370 & ~x389 & ~x466 & ~x521 & ~x522 & ~x547 & ~x728;
assign c8168 =  x457 &  x569 & ~x3 & ~x25 & ~x30 & ~x32 & ~x34 & ~x58 & ~x82 & ~x84 & ~x139 & ~x146 & ~x171 & ~x173 & ~x195 & ~x202 & ~x223 & ~x224 & ~x225 & ~x227 & ~x231 & ~x251 & ~x253 & ~x256 & ~x257 & ~x284 & ~x308 & ~x309 & ~x335 & ~x337 & ~x364 & ~x365 & ~x392 & ~x393 & ~x449 & ~x478 & ~x516 & ~x683 & ~x755 & ~x759 & ~x780 & ~x783;
assign c8170 =  x507 & ~x15 & ~x16 & ~x29 & ~x51 & ~x77 & ~x79 & ~x81 & ~x137 & ~x223 & ~x248 & ~x277 & ~x279 & ~x306 & ~x388 & ~x389 & ~x695 & ~x699 & ~x701 & ~x717 & ~x728 & ~x734 & ~x774;
assign c8172 = ~x9 & ~x33 & ~x35 & ~x50 & ~x63 & ~x66 & ~x73 & ~x75 & ~x78 & ~x92 & ~x137 & ~x142 & ~x204 & ~x231 & ~x253 & ~x258 & ~x280 & ~x308 & ~x315 & ~x334 & ~x363 & ~x465 & ~x715 & ~x762;
assign c8174 =  x406 &  x462 & ~x25 & ~x35 & ~x49 & ~x58 & ~x59 & ~x60 & ~x63 & ~x64 & ~x80 & ~x83 & ~x88 & ~x132 & ~x141 & ~x146 & ~x147 & ~x148 & ~x164 & ~x176 & ~x188 & ~x195 & ~x224 & ~x225 & ~x231 & ~x233 & ~x251 & ~x256 & ~x260 & ~x261 & ~x287 & ~x316 & ~x317 & ~x337 & ~x361 & ~x368 & ~x370 & ~x372 & ~x390 & ~x398 & ~x400 & ~x422 & ~x425 & ~x445 & ~x450 & ~x497 & ~x554 & ~x699 & ~x724 & ~x750 & ~x761 & ~x777;
assign c8176 = ~x14 & ~x51 & ~x80 & ~x82 & ~x109 & ~x111 & ~x112 & ~x139 & ~x164 & ~x192 & ~x219 & ~x274 & ~x277 & ~x302 & ~x303 & ~x305 & ~x330 & ~x331 & ~x361 & ~x376 & ~x386 & ~x414 & ~x459 & ~x485 & ~x513 & ~x653 & ~x764 & ~x774;
assign c8178 = ~x1 & ~x2 & ~x3 & ~x4 & ~x5 & ~x8 & ~x20 & ~x21 & ~x24 & ~x25 & ~x26 & ~x28 & ~x29 & ~x31 & ~x32 & ~x35 & ~x49 & ~x52 & ~x53 & ~x54 & ~x56 & ~x58 & ~x59 & ~x60 & ~x62 & ~x63 & ~x65 & ~x79 & ~x80 & ~x83 & ~x85 & ~x86 & ~x89 & ~x90 & ~x108 & ~x110 & ~x111 & ~x112 & ~x115 & ~x118 & ~x120 & ~x138 & ~x139 & ~x141 & ~x142 & ~x145 & ~x147 & ~x164 & ~x167 & ~x168 & ~x169 & ~x170 & ~x171 & ~x172 & ~x173 & ~x174 & ~x175 & ~x176 & ~x193 & ~x194 & ~x196 & ~x197 & ~x201 & ~x202 & ~x203 & ~x220 & ~x221 & ~x224 & ~x226 & ~x227 & ~x229 & ~x230 & ~x249 & ~x251 & ~x252 & ~x253 & ~x255 & ~x257 & ~x258 & ~x259 & ~x277 & ~x280 & ~x281 & ~x282 & ~x285 & ~x286 & ~x306 & ~x307 & ~x310 & ~x311 & ~x313 & ~x315 & ~x332 & ~x333 & ~x334 & ~x335 & ~x338 & ~x339 & ~x360 & ~x361 & ~x362 & ~x363 & ~x364 & ~x365 & ~x367 & ~x368 & ~x369 & ~x370 & ~x389 & ~x390 & ~x391 & ~x392 & ~x394 & ~x395 & ~x396 & ~x416 & ~x417 & ~x418 & ~x419 & ~x420 & ~x421 & ~x422 & ~x444 & ~x449 & ~x450 & ~x451 & ~x475 & ~x504 & ~x506 & ~x531 & ~x549 & ~x559 & ~x578 & ~x605 & ~x606 & ~x613 & ~x614 & ~x616 & ~x632 & ~x633 & ~x644 & ~x658 & ~x659 & ~x660 & ~x699 & ~x727 & ~x755 & ~x756 & ~x782 & ~x783;
assign c8180 =  x717 & ~x27 & ~x30 & ~x54 & ~x57 & ~x58 & ~x60 & ~x61 & ~x84 & ~x89 & ~x108 & ~x111 & ~x113 & ~x115 & ~x117 & ~x139 & ~x140 & ~x143 & ~x144 & ~x146 & ~x166 & ~x171 & ~x199 & ~x200 & ~x223 & ~x280 & ~x310 & ~x311 & ~x365 & ~x366 & ~x390 & ~x393 & ~x416 & ~x420 & ~x443 & ~x451 & ~x476 & ~x478 & ~x497 & ~x503 & ~x530 & ~x531 & ~x550 & ~x578 & ~x582 & ~x585 & ~x586 & ~x588 & ~x610 & ~x611 & ~x615 & ~x628 & ~x629 & ~x630 & ~x755;
assign c8182 = ~x0 & ~x25 & ~x51 & ~x52 & ~x53 & ~x61 & ~x62 & ~x81 & ~x83 & ~x84 & ~x111 & ~x138 & ~x141 & ~x163 & ~x166 & ~x169 & ~x172 & ~x190 & ~x192 & ~x193 & ~x199 & ~x222 & ~x223 & ~x224 & ~x225 & ~x246 & ~x252 & ~x254 & ~x273 & ~x274 & ~x276 & ~x301 & ~x302 & ~x332 & ~x334 & ~x336 & ~x337 & ~x357 & ~x360 & ~x361 & ~x363 & ~x386 & ~x391 & ~x440 & ~x448 & ~x470 & ~x496 & ~x498 & ~x520 & ~x525 & ~x528 & ~x534 & ~x546 & ~x553 & ~x558 & ~x559 & ~x571 & ~x572 & ~x573 & ~x585 & ~x726 & ~x755 & ~x760 & ~x777 & ~x781;
assign c8184 = ~x0 & ~x5 & ~x22 & ~x24 & ~x25 & ~x26 & ~x28 & ~x52 & ~x54 & ~x57 & ~x60 & ~x80 & ~x81 & ~x86 & ~x104 & ~x106 & ~x109 & ~x110 & ~x133 & ~x136 & ~x138 & ~x139 & ~x141 & ~x142 & ~x143 & ~x167 & ~x195 & ~x198 & ~x217 & ~x219 & ~x221 & ~x224 & ~x245 & ~x246 & ~x252 & ~x274 & ~x275 & ~x279 & ~x305 & ~x331 & ~x336 & ~x360 & ~x391 & ~x415 & ~x416 & ~x419 & ~x443 & ~x444 & ~x446 & ~x447 & ~x502 & ~x503 & ~x504 & ~x527 & ~x531 & ~x558 & ~x576 & ~x600 & ~x602 & ~x603 & ~x643 & ~x757 & ~x779 & ~x782;
assign c8186 = ~x1 & ~x2 & ~x4 & ~x9 & ~x18 & ~x19 & ~x30 & ~x37 & ~x44 & ~x45 & ~x57 & ~x61 & ~x62 & ~x86 & ~x88 & ~x110 & ~x113 & ~x117 & ~x144 & ~x156 & ~x169 & ~x170 & ~x171 & ~x196 & ~x198 & ~x226 & ~x336 & ~x394 & ~x408 & ~x419 & ~x436 & ~x464 & ~x475 & ~x492 & ~x731 & ~x732 & ~x744 & ~x760 & ~x761 & ~x770;
assign c8188 =  x14 &  x235 &  x431 &  x459 & ~x28 & ~x55 & ~x56 & ~x58 & ~x87 & ~x114 & ~x170 & ~x197 & ~x223 & ~x253 & ~x279 & ~x281 & ~x308 & ~x310 & ~x312 & ~x342 & ~x363 & ~x369 & ~x394 & ~x423 & ~x448 & ~x449 & ~x451 & ~x478 & ~x503 & ~x504 & ~x505 & ~x531 & ~x534 & ~x558 & ~x588;
assign c8190 = ~x0 & ~x12 & ~x13 & ~x16 & ~x47 & ~x57 & ~x83 & ~x107 & ~x109 & ~x110 & ~x165 & ~x171 & ~x247 & ~x278 & ~x331 & ~x358 & ~x401 & ~x485 & ~x673 & ~x680 & ~x691 & ~x707 & ~x708 & ~x709 & ~x736 & ~x767;
assign c8192 =  x573 &  x742 & ~x174 & ~x245 & ~x566 & ~x605 & ~x659;
assign c8194 = ~x19 & ~x34 & ~x50 & ~x87 & ~x135 & ~x136 & ~x165 & ~x192 & ~x193 & ~x221 & ~x276 & ~x305 & ~x323 & ~x360 & ~x387 & ~x388 & ~x407 & ~x434 & ~x463 & ~x491 & ~x679;
assign c8196 = ~x2 & ~x30 & ~x105 & ~x110 & ~x113 & ~x114 & ~x116 & ~x134 & ~x135 & ~x195 & ~x225 & ~x226 & ~x248 & ~x252 & ~x274 & ~x275 & ~x276 & ~x282 & ~x285 & ~x305 & ~x330 & ~x332 & ~x335 & ~x358 & ~x359 & ~x361 & ~x365 & ~x391 & ~x392 & ~x393 & ~x398 & ~x443 & ~x447 & ~x451 & ~x572 & ~x585 & ~x700 & ~x702 & ~x705 & ~x706 & ~x711 & ~x712 & ~x728 & ~x739 & ~x748 & ~x753 & ~x774 & ~x775 & ~x781 & ~x782 & ~x783;
assign c8198 =  x101 &  x129 &  x213 &  x241 & ~x26 & ~x31 & ~x52 & ~x53 & ~x87 & ~x104 & ~x107 & ~x137 & ~x188 & ~x217 & ~x246 & ~x274 & ~x275 & ~x307 & ~x387 & ~x475 & ~x640 & ~x697 & ~x783;
assign c8200 =  x509 &  x534 &  x621 & ~x53 & ~x109 & ~x166 & ~x192 & ~x249 & ~x305;
assign c8202 = ~x23 & ~x24 & ~x25 & ~x55 & ~x58 & ~x104 & ~x109 & ~x115 & ~x136 & ~x141 & ~x171 & ~x172 & ~x194 & ~x227 & ~x246 & ~x248 & ~x256 & ~x281 & ~x303 & ~x311 & ~x313 & ~x333 & ~x361 & ~x391 & ~x418 & ~x438 & ~x443 & ~x446 & ~x451 & ~x465 & ~x475 & ~x493 & ~x505 & ~x528 & ~x548 & ~x561 & ~x576 & ~x601 & ~x602 & ~x646 & ~x698;
assign c8204 =  x539 &  x735 & ~x0 & ~x1 & ~x25 & ~x30 & ~x52 & ~x53 & ~x81 & ~x83 & ~x84 & ~x108 & ~x110 & ~x111 & ~x114 & ~x137 & ~x141 & ~x143 & ~x165 & ~x166 & ~x170 & ~x224 & ~x252 & ~x420 & ~x612;
assign c8206 =  x352 &  x433 & ~x5 & ~x26 & ~x58 & ~x82 & ~x105 & ~x111 & ~x117 & ~x135 & ~x163 & ~x189 & ~x199 & ~x202 & ~x204 & ~x226 & ~x232 & ~x249 & ~x257 & ~x279 & ~x281 & ~x308 & ~x312 & ~x316 & ~x317 & ~x331 & ~x340 & ~x387 & ~x395 & ~x444 & ~x448 & ~x452 & ~x453 & ~x477 & ~x501 & ~x533 & ~x640 & ~x675 & ~x724 & ~x753 & ~x779;
assign c8208 =  x402 &  x652 & ~x4 & ~x27 & ~x32 & ~x57 & ~x58 & ~x59 & ~x61 & ~x82 & ~x86 & ~x90 & ~x111 & ~x115 & ~x117 & ~x138 & ~x142 & ~x145 & ~x146 & ~x168 & ~x195 & ~x223 & ~x226 & ~x254 & ~x280 & ~x281 & ~x282 & ~x308 & ~x310 & ~x312 & ~x340 & ~x391 & ~x397 & ~x421 & ~x425 & ~x448 & ~x521 & ~x588 & ~x750 & ~x760 & ~x762 & ~x779;
assign c8210 =  x396 & ~x164 & ~x278 & ~x360 & ~x387 & ~x458 & ~x485 & ~x541 & ~x729 & ~x764;
assign c8212 =  x747 & ~x86 & ~x87 & ~x110 & ~x134 & ~x167 & ~x189 & ~x198 & ~x224 & ~x250 & ~x362 & ~x366 & ~x387 & ~x388 & ~x394 & ~x395 & ~x470 & ~x506 & ~x555 & ~x581 & ~x606 & ~x633 & ~x644 & ~x656 & ~x728;
assign c8214 = ~x11 & ~x24 & ~x82 & ~x164 & ~x195 & ~x276 & ~x278 & ~x295 & ~x322 & ~x387 & ~x406 & ~x435 & ~x462 & ~x624 & ~x707 & ~x783;
assign c8216 =  x750 & ~x138 & ~x162 & ~x191 & ~x246 & ~x366 & ~x395 & ~x629 & ~x632 & ~x657 & ~x686;
assign c8218 = ~x3 & ~x25 & ~x27 & ~x28 & ~x29 & ~x49 & ~x50 & ~x51 & ~x54 & ~x56 & ~x58 & ~x77 & ~x79 & ~x82 & ~x85 & ~x97 & ~x108 & ~x109 & ~x114 & ~x116 & ~x133 & ~x134 & ~x135 & ~x137 & ~x138 & ~x141 & ~x144 & ~x164 & ~x165 & ~x166 & ~x168 & ~x169 & ~x170 & ~x189 & ~x191 & ~x192 & ~x195 & ~x196 & ~x199 & ~x200 & ~x219 & ~x220 & ~x222 & ~x223 & ~x227 & ~x247 & ~x253 & ~x254 & ~x274 & ~x275 & ~x277 & ~x278 & ~x279 & ~x280 & ~x281 & ~x282 & ~x303 & ~x306 & ~x308 & ~x310 & ~x333 & ~x334 & ~x336 & ~x338 & ~x360 & ~x361 & ~x362 & ~x364 & ~x366 & ~x387 & ~x392 & ~x393 & ~x394 & ~x395 & ~x415 & ~x417 & ~x419 & ~x420 & ~x442 & ~x444 & ~x445 & ~x449 & ~x451 & ~x470 & ~x473 & ~x477 & ~x498 & ~x501 & ~x502 & ~x505 & ~x576 & ~x577 & ~x604 & ~x616 & ~x630 & ~x640 & ~x642 & ~x728 & ~x731 & ~x755 & ~x783;
assign c8220 = ~x11 & ~x17 & ~x42 & ~x53 & ~x57 & ~x109 & ~x176 & ~x348 & ~x387 & ~x460 & ~x516 & ~x528 & ~x767;
assign c8222 =  x616 & ~x83 & ~x138 & ~x573 & ~x702;
assign c8224 = ~x2 & ~x25 & ~x65 & ~x66 & ~x67 & ~x89 & ~x150 & ~x177 & ~x178 & ~x205 & ~x222 & ~x225 & ~x227 & ~x257 & ~x258 & ~x262 & ~x313 & ~x336 & ~x390 & ~x424 & ~x426 & ~x607 & ~x636 & ~x658 & ~x761;
assign c8226 =  x406 & ~x31 & ~x36 & ~x55 & ~x60 & ~x61 & ~x63 & ~x77 & ~x81 & ~x83 & ~x86 & ~x92 & ~x105 & ~x113 & ~x119 & ~x121 & ~x137 & ~x138 & ~x145 & ~x147 & ~x161 & ~x163 & ~x172 & ~x174 & ~x176 & ~x188 & ~x190 & ~x196 & ~x198 & ~x201 & ~x202 & ~x203 & ~x221 & ~x230 & ~x244 & ~x251 & ~x252 & ~x259 & ~x260 & ~x261 & ~x272 & ~x285 & ~x286 & ~x316 & ~x342 & ~x344 & ~x359 & ~x372 & ~x391 & ~x398 & ~x427 & ~x428 & ~x449 & ~x450 & ~x452 & ~x455 & ~x469 & ~x500 & ~x525 & ~x551 & ~x552 & ~x642 & ~x729 & ~x761 & ~x783;
assign c8228 = ~x56 & ~x63 & ~x102 & ~x130 & ~x177 & ~x216 & ~x262 & ~x270 & ~x271 & ~x305 & ~x344 & ~x346 & ~x373 & ~x497 & ~x498 & ~x531 & ~x550 & ~x703 & ~x725;
assign c8230 =  x183 &  x211 &  x239 &  x295 &  x407 & ~x102 & ~x135 & ~x143 & ~x158 & ~x162 & ~x188 & ~x192 & ~x219 & ~x249 & ~x254 & ~x273 & ~x283 & ~x328 & ~x356 & ~x384 & ~x385 & ~x389 & ~x418 & ~x419 & ~x440 & ~x441 & ~x467 & ~x504 & ~x673 & ~x757;
assign c8232 = ~x4 & ~x6 & ~x35 & ~x36 & ~x63 & ~x88 & ~x125 & ~x173 & ~x193 & ~x195 & ~x220 & ~x222 & ~x249 & ~x277 & ~x281 & ~x307 & ~x359 & ~x360 & ~x361 & ~x367 & ~x415 & ~x421 & ~x521 & ~x574 & ~x671 & ~x730 & ~x733 & ~x740 & ~x750 & ~x767 & ~x775;
assign c8234 = ~x23 & ~x34 & ~x53 & ~x55 & ~x58 & ~x62 & ~x75 & ~x77 & ~x78 & ~x86 & ~x101 & ~x111 & ~x114 & ~x120 & ~x164 & ~x166 & ~x193 & ~x197 & ~x221 & ~x222 & ~x251 & ~x259 & ~x280 & ~x364 & ~x417 & ~x445 & ~x446 & ~x476 & ~x477 & ~x519 & ~x547 & ~x548 & ~x743 & ~x770 & ~x783;
assign c8236 =  x545 &  x743 & ~x25 & ~x31 & ~x338 & ~x363 & ~x386 & ~x469 & ~x496 & ~x526 & ~x538 & ~x579 & ~x633 & ~x687;
assign c8238 =  x491 &  x544 & ~x0 & ~x4 & ~x22 & ~x23 & ~x26 & ~x106 & ~x110 & ~x140 & ~x144 & ~x188 & ~x195 & ~x218 & ~x228 & ~x275 & ~x284 & ~x302 & ~x304 & ~x340 & ~x359 & ~x362 & ~x368 & ~x388 & ~x391 & ~x395 & ~x413 & ~x441 & ~x442 & ~x443 & ~x447 & ~x469 & ~x480 & ~x481 & ~x482 & ~x483 & ~x527 & ~x553 & ~x558 & ~x560 & ~x580 & ~x583 & ~x605 & ~x611 & ~x617 & ~x668 & ~x670 & ~x671 & ~x698 & ~x760 & ~x783;
assign c8240 =  x380 & ~x76 & ~x103 & ~x105 & ~x110 & ~x115 & ~x116 & ~x139 & ~x173 & ~x187 & ~x194 & ~x196 & ~x226 & ~x248 & ~x250 & ~x278 & ~x299 & ~x301 & ~x304 & ~x305 & ~x306 & ~x355 & ~x384 & ~x387 & ~x395 & ~x412 & ~x439 & ~x440 & ~x441 & ~x448 & ~x468 & ~x496 & ~x498 & ~x643 & ~x696 & ~x720 & ~x736 & ~x776;
assign c8242 =  x459 &  x624 & ~x3 & ~x27 & ~x55 & ~x81 & ~x82 & ~x87 & ~x91 & ~x113 & ~x114 & ~x116 & ~x138 & ~x140 & ~x147 & ~x165 & ~x166 & ~x175 & ~x193 & ~x195 & ~x197 & ~x198 & ~x227 & ~x230 & ~x256 & ~x258 & ~x282 & ~x283 & ~x285 & ~x309 & ~x310 & ~x311 & ~x336 & ~x338 & ~x366 & ~x367 & ~x392 & ~x394 & ~x397 & ~x422 & ~x426 & ~x453 & ~x474 & ~x475 & ~x476 & ~x522 & ~x560 & ~x588 & ~x643 & ~x779;
assign c8244 =  x743 &  x744 & ~x276 & ~x442 & ~x498 & ~x512 & ~x579 & ~x633 & ~x660 & ~x662 & ~x687;
assign c8246 = ~x23 & ~x24 & ~x26 & ~x140 & ~x219 & ~x245 & ~x246 & ~x331 & ~x385 & ~x392 & ~x461 & ~x488 & ~x515 & ~x571 & ~x572 & ~x584 & ~x656 & ~x710 & ~x780;
assign c8248 = ~x7 & ~x11 & ~x21 & ~x22 & ~x28 & ~x36 & ~x37 & ~x49 & ~x56 & ~x65 & ~x76 & ~x81 & ~x136 & ~x138 & ~x141 & ~x164 & ~x191 & ~x195 & ~x222 & ~x249 & ~x251 & ~x252 & ~x303 & ~x304 & ~x306 & ~x307 & ~x332 & ~x358 & ~x359 & ~x360 & ~x461 & ~x717 & ~x739 & ~x744 & ~x755 & ~x761 & ~x771;
assign c8250 =  x483 &  x592 &  x706 & ~x451 & ~x627;
assign c8252 = ~x2 & ~x6 & ~x23 & ~x25 & ~x32 & ~x48 & ~x49 & ~x53 & ~x57 & ~x58 & ~x59 & ~x81 & ~x92 & ~x103 & ~x113 & ~x114 & ~x119 & ~x120 & ~x121 & ~x131 & ~x143 & ~x159 & ~x160 & ~x163 & ~x166 & ~x167 & ~x171 & ~x175 & ~x176 & ~x177 & ~x188 & ~x194 & ~x196 & ~x199 & ~x202 & ~x205 & ~x206 & ~x215 & ~x222 & ~x223 & ~x233 & ~x234 & ~x249 & ~x252 & ~x260 & ~x261 & ~x278 & ~x279 & ~x281 & ~x286 & ~x287 & ~x289 & ~x306 & ~x307 & ~x315 & ~x317 & ~x334 & ~x336 & ~x362 & ~x371 & ~x372 & ~x373 & ~x393 & ~x411 & ~x412 & ~x421 & ~x440 & ~x449 & ~x474 & ~x522 & ~x523 & ~x524 & ~x560 & ~x587 & ~x671 & ~x728 & ~x733;
assign c8254 =  x518 &  x718 &  x737 & ~x470;
assign c8256 =  x645 & ~x26 & ~x57 & ~x60 & ~x338 & ~x408 & ~x464 & ~x491 & ~x505 & ~x518;
assign c8258 =  x269 &  x353 & ~x22 & ~x25 & ~x26 & ~x30 & ~x50 & ~x52 & ~x79 & ~x105 & ~x109 & ~x110 & ~x135 & ~x137 & ~x138 & ~x162 & ~x192 & ~x194 & ~x219 & ~x221 & ~x222 & ~x248 & ~x274 & ~x280 & ~x302 & ~x334 & ~x364 & ~x391 & ~x419 & ~x498 & ~x525 & ~x551 & ~x556 & ~x582 & ~x603 & ~x629;
assign c8260 =  x733;
assign c8262 =  x375 & ~x2 & ~x28 & ~x29 & ~x30 & ~x56 & ~x82 & ~x83 & ~x85 & ~x88 & ~x111 & ~x114 & ~x119 & ~x137 & ~x140 & ~x142 & ~x148 & ~x167 & ~x168 & ~x171 & ~x174 & ~x175 & ~x176 & ~x196 & ~x201 & ~x203 & ~x204 & ~x221 & ~x228 & ~x231 & ~x250 & ~x256 & ~x257 & ~x259 & ~x260 & ~x278 & ~x279 & ~x287 & ~x335 & ~x362 & ~x364 & ~x390 & ~x391 & ~x419 & ~x446 & ~x447 & ~x448 & ~x501 & ~x503 & ~x504 & ~x549 & ~x558 & ~x560 & ~x577 & ~x587 & ~x602;
assign c8264 =  x454 &  x594 &  x706 & ~x28 & ~x44 & ~x143 & ~x166 & ~x569;
assign c8266 = ~x12 & ~x21 & ~x22 & ~x38 & ~x50 & ~x55 & ~x80 & ~x84 & ~x106 & ~x108 & ~x109 & ~x110 & ~x111 & ~x137 & ~x139 & ~x166 & ~x248 & ~x249 & ~x276 & ~x304 & ~x305 & ~x333 & ~x336 & ~x358 & ~x360 & ~x375 & ~x387 & ~x402 & ~x403 & ~x430 & ~x431 & ~x458 & ~x515 & ~x753 & ~x756 & ~x757 & ~x762 & ~x781;
assign c8268 =  x720 & ~x3 & ~x55 & ~x59 & ~x81 & ~x83 & ~x106 & ~x115 & ~x133 & ~x135 & ~x136 & ~x163 & ~x190 & ~x191 & ~x195 & ~x196 & ~x218 & ~x219 & ~x220 & ~x221 & ~x222 & ~x246 & ~x248 & ~x250 & ~x274 & ~x275 & ~x302 & ~x306 & ~x307 & ~x333 & ~x359 & ~x364 & ~x388 & ~x394 & ~x418 & ~x471 & ~x472 & ~x498 & ~x499 & ~x526 & ~x556 & ~x557 & ~x614 & ~x628 & ~x630;
assign c8270 =  x404 & ~x11 & ~x29 & ~x30 & ~x37 & ~x39 & ~x54 & ~x65 & ~x91 & ~x121 & ~x138 & ~x139 & ~x140 & ~x141 & ~x143 & ~x170 & ~x172 & ~x176 & ~x197 & ~x224 & ~x226 & ~x259 & ~x278 & ~x286 & ~x306 & ~x334 & ~x335 & ~x338 & ~x398 & ~x422 & ~x426 & ~x483 & ~x504 & ~x532 & ~x606;
assign c8272 = ~x16 & ~x30 & ~x52 & ~x79 & ~x105 & ~x107 & ~x111 & ~x131 & ~x135 & ~x139 & ~x162 & ~x164 & ~x166 & ~x167 & ~x192 & ~x217 & ~x219 & ~x220 & ~x246 & ~x277 & ~x301 & ~x305 & ~x331 & ~x333 & ~x357 & ~x358 & ~x361 & ~x386 & ~x387 & ~x420 & ~x489 & ~x683 & ~x739 & ~x742 & ~x752 & ~x753 & ~x754 & ~x761 & ~x767 & ~x772 & ~x773;
assign c8274 =  x480 & ~x305 & ~x355 & ~x361 & ~x403 & ~x542 & ~x543 & ~x750 & ~x758;
assign c8276 =  x454 &  x705 & ~x199 & ~x279 & ~x448 & ~x625 & ~x758;
assign c8278 =  x520 &  x545 &  x547 & ~x25 & ~x86 & ~x217 & ~x286 & ~x305 & ~x328 & ~x329 & ~x369 & ~x426 & ~x443 & ~x472 & ~x580 & ~x590 & ~x604 & ~x606 & ~x616 & ~x726;
assign c8280 =  x295 &  x403 &  x431 & ~x2 & ~x4 & ~x6 & ~x29 & ~x31 & ~x36 & ~x57 & ~x84 & ~x85 & ~x86 & ~x101 & ~x109 & ~x110 & ~x118 & ~x139 & ~x142 & ~x143 & ~x147 & ~x168 & ~x171 & ~x172 & ~x174 & ~x199 & ~x200 & ~x201 & ~x226 & ~x227 & ~x230 & ~x252 & ~x257 & ~x283 & ~x285 & ~x286 & ~x309 & ~x310 & ~x338 & ~x366 & ~x367 & ~x368 & ~x369 & ~x392 & ~x394 & ~x419 & ~x423 & ~x425 & ~x446 & ~x447 & ~x449 & ~x452 & ~x477 & ~x480 & ~x502 & ~x532 & ~x533 & ~x534 & ~x560 & ~x561 & ~x699;
assign c8282 =  x288 &  x372 &  x651 & ~x3 & ~x25 & ~x26 & ~x27 & ~x29 & ~x56 & ~x60 & ~x82 & ~x84 & ~x110 & ~x168 & ~x169 & ~x173 & ~x224 & ~x251 & ~x252 & ~x366 & ~x392 & ~x448 & ~x544 & ~x545 & ~x572 & ~x599 & ~x601 & ~x656;
assign c8284 =  x483 & ~x0 & ~x5 & ~x26 & ~x28 & ~x31 & ~x34 & ~x54 & ~x57 & ~x58 & ~x87 & ~x88 & ~x89 & ~x110 & ~x112 & ~x114 & ~x117 & ~x139 & ~x140 & ~x145 & ~x146 & ~x168 & ~x173 & ~x195 & ~x196 & ~x199 & ~x224 & ~x225 & ~x226 & ~x253 & ~x255 & ~x281 & ~x310 & ~x311 & ~x312 & ~x339 & ~x340 & ~x420 & ~x422 & ~x450 & ~x477 & ~x514 & ~x542 & ~x570 & ~x757 & ~x766;
assign c8286 =  x505 & ~x108 & ~x249 & ~x375 & ~x430 & ~x515;
assign c8288 =  x746 & ~x83 & ~x86 & ~x110 & ~x112 & ~x162 & ~x164 & ~x166 & ~x220 & ~x387 & ~x394 & ~x415 & ~x417 & ~x471 & ~x498 & ~x499 & ~x527 & ~x607 & ~x608 & ~x634 & ~x643 & ~x655 & ~x658 & ~x730;
assign c8290 = ~x12 & ~x14 & ~x23 & ~x25 & ~x27 & ~x39 & ~x40 & ~x51 & ~x79 & ~x81 & ~x82 & ~x105 & ~x110 & ~x111 & ~x133 & ~x162 & ~x165 & ~x190 & ~x192 & ~x196 & ~x218 & ~x219 & ~x221 & ~x246 & ~x247 & ~x274 & ~x275 & ~x302 & ~x303 & ~x305 & ~x331 & ~x332 & ~x357 & ~x359 & ~x385 & ~x386 & ~x547 & ~x643 & ~x670 & ~x683 & ~x699 & ~x727 & ~x753 & ~x754 & ~x761 & ~x766 & ~x782;
assign c8292 =  x401 &  x429 &  x569 & ~x24 & ~x26 & ~x28 & ~x55 & ~x60 & ~x62 & ~x112 & ~x118 & ~x138 & ~x140 & ~x168 & ~x224 & ~x252 & ~x392 & ~x449 & ~x545 & ~x656 & ~x657 & ~x684 & ~x685 & ~x761;
assign c8294 = ~x18 & ~x21 & ~x22 & ~x25 & ~x44 & ~x45 & ~x49 & ~x50 & ~x51 & ~x57 & ~x77 & ~x80 & ~x108 & ~x135 & ~x163 & ~x191 & ~x193 & ~x196 & ~x197 & ~x219 & ~x220 & ~x248 & ~x250 & ~x276 & ~x279 & ~x303 & ~x304 & ~x331 & ~x332 & ~x333 & ~x334 & ~x349 & ~x350 & ~x358 & ~x361 & ~x404 & ~x405 & ~x414 & ~x416 & ~x417 & ~x418 & ~x433 & ~x461 & ~x489 & ~x729 & ~x747 & ~x757 & ~x776;
assign c8296 =  x463 &  x740 & ~x55 & ~x124 & ~x141 & ~x331 & ~x397 & ~x414 & ~x455 & ~x482 & ~x497 & ~x508 & ~x527 & ~x552 & ~x553 & ~x583;
assign c8298 =  x573 &  x740 & ~x68 & ~x384 & ~x442 & ~x454 & ~x589 & ~x611;
assign c8300 = ~x12 & ~x77 & ~x122 & ~x305 & ~x333 & ~x360 & ~x401 & ~x402 & ~x428 & ~x485 & ~x513 & ~x707 & ~x737;
assign c8302 =  x649 & ~x59 & ~x81 & ~x86 & ~x136 & ~x142 & ~x165 & ~x193 & ~x197 & ~x248 & ~x330 & ~x333 & ~x366 & ~x470 & ~x498 & ~x500 & ~x596;
assign c8304 =  x482 &  x537 &  x592 & ~x19 & ~x27 & ~x30 & ~x54 & ~x55 & ~x56 & ~x83 & ~x84 & ~x85 & ~x87 & ~x110 & ~x114 & ~x116 & ~x138 & ~x139 & ~x141 & ~x168 & ~x196 & ~x198 & ~x224 & ~x225 & ~x253 & ~x279 & ~x280 & ~x281 & ~x309 & ~x362 & ~x391 & ~x446 & ~x447 & ~x448 & ~x449 & ~x462 & ~x476 & ~x477 & ~x505 & ~x519 & ~x531 & ~x532 & ~x755;
assign c8306 =  x678 & ~x85 & ~x113 & ~x196 & ~x200 & ~x201 & ~x256 & ~x258 & ~x311 & ~x481 & ~x577 & ~x602 & ~x603 & ~x760;
assign c8308 =  x127 &  x211 &  x379 &  x433 & ~x23 & ~x85 & ~x105 & ~x113 & ~x114 & ~x143 & ~x167 & ~x201 & ~x220 & ~x328 & ~x330 & ~x333 & ~x342 & ~x371 & ~x385 & ~x394 & ~x396 & ~x423 & ~x440 & ~x449 & ~x470 & ~x509 & ~x524 & ~x583 & ~x584 & ~x614 & ~x702 & ~x731 & ~x751 & ~x758 & ~x783;
assign c8310 =  x429 & ~x22 & ~x26 & ~x28 & ~x30 & ~x33 & ~x64 & ~x78 & ~x79 & ~x88 & ~x89 & ~x106 & ~x113 & ~x118 & ~x141 & ~x143 & ~x169 & ~x171 & ~x172 & ~x173 & ~x193 & ~x199 & ~x200 & ~x221 & ~x222 & ~x225 & ~x226 & ~x229 & ~x249 & ~x255 & ~x258 & ~x278 & ~x282 & ~x283 & ~x306 & ~x309 & ~x333 & ~x334 & ~x336 & ~x361 & ~x393 & ~x421 & ~x449 & ~x503 & ~x671 & ~x749 & ~x761 & ~x777 & ~x780 & ~x783;
assign c8312 =  x719 & ~x26 & ~x57 & ~x167 & ~x227 & ~x244 & ~x422 & ~x551 & ~x579 & ~x582 & ~x606 & ~x627 & ~x628 & ~x630 & ~x631;
assign c8314 = ~x82 & ~x163 & ~x192 & ~x218 & ~x219 & ~x276 & ~x294 & ~x305 & ~x322 & ~x350 & ~x359 & ~x360 & ~x378 & ~x406 & ~x434 & ~x513 & ~x569 & ~x625 & ~x690;
assign c8316 =  x379 &  x514 &  x736 & ~x25 & ~x54 & ~x79 & ~x86 & ~x133 & ~x164 & ~x199 & ~x227 & ~x254 & ~x423 & ~x424 & ~x451 & ~x502 & ~x508 & ~x530 & ~x558;
assign c8318 = ~x5 & ~x6 & ~x17 & ~x19 & ~x25 & ~x29 & ~x46 & ~x51 & ~x59 & ~x72 & ~x74 & ~x85 & ~x88 & ~x101 & ~x111 & ~x112 & ~x117 & ~x138 & ~x142 & ~x165 & ~x167 & ~x198 & ~x221 & ~x249 & ~x254 & ~x278 & ~x296 & ~x306 & ~x337 & ~x364 & ~x365 & ~x367 & ~x389 & ~x416 & ~x417 & ~x419 & ~x420 & ~x492 & ~x576 & ~x684 & ~x758;
assign c8320 =  x663 & ~x76 & ~x104 & ~x132 & ~x188 & ~x219 & ~x223 & ~x276 & ~x303 & ~x308 & ~x330 & ~x334 & ~x357 & ~x391 & ~x470 & ~x527 & ~x551 & ~x553 & ~x580 & ~x775;
assign c8322 =  x407 &  x688 &  x689 & ~x131 & ~x221 & ~x242 & ~x299 & ~x362 & ~x384 & ~x525;
assign c8324 =  x720 & ~x0 & ~x22 & ~x29 & ~x56 & ~x80 & ~x82 & ~x83 & ~x84 & ~x104 & ~x111 & ~x141 & ~x161 & ~x162 & ~x164 & ~x165 & ~x168 & ~x169 & ~x190 & ~x194 & ~x197 & ~x198 & ~x218 & ~x219 & ~x220 & ~x245 & ~x247 & ~x253 & ~x274 & ~x279 & ~x280 & ~x302 & ~x303 & ~x306 & ~x308 & ~x332 & ~x335 & ~x337 & ~x338 & ~x359 & ~x361 & ~x363 & ~x366 & ~x389 & ~x390 & ~x391 & ~x393 & ~x394 & ~x416 & ~x419 & ~x420 & ~x446 & ~x447 & ~x449 & ~x450 & ~x470 & ~x471 & ~x474 & ~x475 & ~x477 & ~x502 & ~x504 & ~x527 & ~x528 & ~x529 & ~x531 & ~x555 & ~x558 & ~x560 & ~x585 & ~x629 & ~x631 & ~x642 & ~x756;
assign c8326 = ~x3 & ~x21 & ~x28 & ~x54 & ~x56 & ~x75 & ~x107 & ~x115 & ~x127 & ~x135 & ~x139 & ~x163 & ~x171 & ~x195 & ~x218 & ~x220 & ~x246 & ~x275 & ~x278 & ~x280 & ~x303 & ~x305 & ~x306 & ~x330 & ~x358 & ~x386 & ~x458 & ~x459 & ~x585 & ~x587 & ~x608 & ~x671 & ~x693 & ~x696 & ~x710 & ~x756;
assign c8328 =  x545 &  x546 &  x743 & ~x78 & ~x108 & ~x120 & ~x232 & ~x258 & ~x498 & ~x551 & ~x578;
assign c8330 = ~x3 & ~x4 & ~x5 & ~x6 & ~x24 & ~x27 & ~x28 & ~x31 & ~x32 & ~x52 & ~x54 & ~x55 & ~x56 & ~x89 & ~x90 & ~x101 & ~x107 & ~x113 & ~x118 & ~x137 & ~x139 & ~x141 & ~x145 & ~x146 & ~x173 & ~x194 & ~x226 & ~x251 & ~x310 & ~x311 & ~x335 & ~x366 & ~x408 & ~x418 & ~x436 & ~x447 & ~x547 & ~x604 & ~x630 & ~x633 & ~x732 & ~x758 & ~x760 & ~x763 & ~x770;
assign c8332 =  x511 & ~x0 & ~x1 & ~x2 & ~x3 & ~x4 & ~x23 & ~x24 & ~x25 & ~x26 & ~x28 & ~x29 & ~x30 & ~x31 & ~x34 & ~x53 & ~x54 & ~x55 & ~x57 & ~x59 & ~x62 & ~x83 & ~x85 & ~x86 & ~x88 & ~x89 & ~x110 & ~x114 & ~x115 & ~x117 & ~x118 & ~x140 & ~x142 & ~x143 & ~x144 & ~x165 & ~x168 & ~x169 & ~x170 & ~x171 & ~x173 & ~x193 & ~x194 & ~x195 & ~x197 & ~x198 & ~x200 & ~x201 & ~x223 & ~x229 & ~x250 & ~x251 & ~x252 & ~x254 & ~x255 & ~x256 & ~x277 & ~x279 & ~x280 & ~x281 & ~x282 & ~x283 & ~x305 & ~x309 & ~x310 & ~x312 & ~x334 & ~x337 & ~x363 & ~x364 & ~x365 & ~x393 & ~x394 & ~x395 & ~x420 & ~x421 & ~x423 & ~x424 & ~x446 & ~x447 & ~x449 & ~x450 & ~x451 & ~x476 & ~x478 & ~x502 & ~x503 & ~x505 & ~x517 & ~x518 & ~x529 & ~x530 & ~x531 & ~x543 & ~x544 & ~x557 & ~x558 & ~x559 & ~x560 & ~x586 & ~x587 & ~x614 & ~x643 & ~x644 & ~x731 & ~x755 & ~x756 & ~x759 & ~x783;
assign c8334 =  x400 &  x428 &  x456 &  x679 & ~x0 & ~x1 & ~x2 & ~x3 & ~x24 & ~x27 & ~x29 & ~x31 & ~x56 & ~x58 & ~x60 & ~x61 & ~x82 & ~x83 & ~x84 & ~x85 & ~x88 & ~x89 & ~x114 & ~x116 & ~x138 & ~x139 & ~x140 & ~x141 & ~x143 & ~x145 & ~x168 & ~x169 & ~x170 & ~x171 & ~x172 & ~x196 & ~x197 & ~x224 & ~x225 & ~x226 & ~x252 & ~x253 & ~x254 & ~x281 & ~x364 & ~x365 & ~x420 & ~x423 & ~x448 & ~x517 & ~x572 & ~x573 & ~x628 & ~x699 & ~x726 & ~x760;
assign c8336 = ~x21 & ~x23 & ~x26 & ~x34 & ~x46 & ~x48 & ~x53 & ~x58 & ~x62 & ~x73 & ~x74 & ~x85 & ~x86 & ~x88 & ~x100 & ~x112 & ~x113 & ~x117 & ~x118 & ~x142 & ~x143 & ~x146 & ~x167 & ~x171 & ~x194 & ~x196 & ~x200 & ~x202 & ~x223 & ~x226 & ~x252 & ~x282 & ~x283 & ~x285 & ~x307 & ~x311 & ~x337 & ~x340 & ~x354 & ~x368 & ~x369 & ~x381 & ~x392 & ~x393 & ~x394 & ~x395 & ~x409 & ~x422 & ~x437 & ~x447 & ~x464 & ~x465 & ~x505 & ~x549 & ~x720 & ~x721 & ~x761;
assign c8338 = ~x0 & ~x4 & ~x9 & ~x28 & ~x59 & ~x61 & ~x63 & ~x81 & ~x84 & ~x85 & ~x92 & ~x117 & ~x118 & ~x140 & ~x141 & ~x144 & ~x147 & ~x171 & ~x197 & ~x199 & ~x201 & ~x226 & ~x227 & ~x231 & ~x253 & ~x255 & ~x257 & ~x280 & ~x282 & ~x313 & ~x314 & ~x337 & ~x409 & ~x448 & ~x464 & ~x520 & ~x521 & ~x577 & ~x603 & ~x720 & ~x766 & ~x767;
assign c8340 =  x456 &  x539;
assign c8342 = ~x10 & ~x22 & ~x24 & ~x28 & ~x30 & ~x49 & ~x109 & ~x129 & ~x137 & ~x168 & ~x192 & ~x225 & ~x251 & ~x253 & ~x278 & ~x305 & ~x388 & ~x389 & ~x390 & ~x391 & ~x416 & ~x475 & ~x518 & ~x528 & ~x545 & ~x699 & ~x725 & ~x728 & ~x734 & ~x742 & ~x758 & ~x759 & ~x768 & ~x774;
assign c8344 = ~x0 & ~x18 & ~x31 & ~x47 & ~x49 & ~x53 & ~x59 & ~x73 & ~x106 & ~x108 & ~x135 & ~x138 & ~x160 & ~x165 & ~x189 & ~x217 & ~x220 & ~x224 & ~x244 & ~x251 & ~x272 & ~x275 & ~x301 & ~x303 & ~x336 & ~x357 & ~x384 & ~x387 & ~x432 & ~x459 & ~x460 & ~x488 & ~x516 & ~x572;
assign c8346 =  x267 &  x295 &  x351 &  x407 &  x435 & ~x27 & ~x55 & ~x75 & ~x77 & ~x103 & ~x106 & ~x107 & ~x130 & ~x134 & ~x139 & ~x161 & ~x163 & ~x167 & ~x168 & ~x189 & ~x190 & ~x196 & ~x214 & ~x221 & ~x251 & ~x272 & ~x273 & ~x276 & ~x302 & ~x303 & ~x309 & ~x327 & ~x331 & ~x334 & ~x390 & ~x412 & ~x414 & ~x448 & ~x499 & ~x501 & ~x524 & ~x525 & ~x641 & ~x669 & ~x729 & ~x753 & ~x782;
assign c8348 = ~x17 & ~x21 & ~x24 & ~x30 & ~x49 & ~x53 & ~x70 & ~x74 & ~x82 & ~x84 & ~x105 & ~x110 & ~x131 & ~x137 & ~x138 & ~x139 & ~x189 & ~x190 & ~x217 & ~x220 & ~x246 & ~x303 & ~x332 & ~x337 & ~x358 & ~x359 & ~x386 & ~x570 & ~x641 & ~x642 & ~x710 & ~x725 & ~x738 & ~x759;
assign c8350 =  x768 & ~x0 & ~x83 & ~x104 & ~x109 & ~x133 & ~x138 & ~x158 & ~x159 & ~x163 & ~x168 & ~x186 & ~x188 & ~x189 & ~x190 & ~x199 & ~x200 & ~x215 & ~x218 & ~x244 & ~x249 & ~x253 & ~x270 & ~x271 & ~x273 & ~x281 & ~x298 & ~x299 & ~x305 & ~x328 & ~x332 & ~x355 & ~x356 & ~x357 & ~x383 & ~x384 & ~x412 & ~x425 & ~x439 & ~x442 & ~x468 & ~x499 & ~x559 & ~x615;
assign c8352 =  x16 &  x595 & ~x231;
assign c8354 = ~x1 & ~x3 & ~x26 & ~x110 & ~x111 & ~x137 & ~x142 & ~x169 & ~x190 & ~x191 & ~x217 & ~x220 & ~x247 & ~x250 & ~x279 & ~x307 & ~x329 & ~x364 & ~x388 & ~x441 & ~x458 & ~x516 & ~x729 & ~x737 & ~x738 & ~x765;
assign c8356 = ~x3 & ~x30 & ~x32 & ~x56 & ~x60 & ~x80 & ~x83 & ~x84 & ~x86 & ~x108 & ~x113 & ~x116 & ~x143 & ~x162 & ~x164 & ~x165 & ~x172 & ~x198 & ~x218 & ~x219 & ~x223 & ~x253 & ~x307 & ~x331 & ~x332 & ~x333 & ~x335 & ~x336 & ~x358 & ~x365 & ~x366 & ~x385 & ~x392 & ~x394 & ~x419 & ~x420 & ~x446 & ~x518 & ~x545 & ~x546 & ~x555 & ~x571 & ~x701 & ~x710 & ~x737 & ~x758 & ~x760 & ~x775;
assign c8358 = ~x18 & ~x33 & ~x37 & ~x47 & ~x62 & ~x75 & ~x78 & ~x81 & ~x85 & ~x87 & ~x104 & ~x107 & ~x117 & ~x136 & ~x144 & ~x162 & ~x164 & ~x190 & ~x222 & ~x225 & ~x251 & ~x278 & ~x306 & ~x307 & ~x308 & ~x332 & ~x333 & ~x357 & ~x359 & ~x385 & ~x546 & ~x585 & ~x640 & ~x646 & ~x704 & ~x707 & ~x710 & ~x760 & ~x781;
assign c8360 =  x14 &  x459 & ~x85 & ~x108 & ~x113 & ~x130 & ~x136 & ~x144 & ~x164 & ~x194 & ~x195 & ~x227 & ~x256 & ~x339 & ~x362 & ~x366 & ~x367 & ~x396 & ~x397 & ~x427 & ~x453 & ~x756;
assign c8362 =  x735 & ~x116 & ~x117 & ~x166 & ~x172 & ~x223 & ~x255 & ~x256 & ~x334 & ~x340 & ~x341 & ~x363 & ~x606 & ~x644 & ~x654 & ~x656;
assign c8364 =  x504;
assign c8366 =  x425 &  x506 & ~x81 & ~x167 & ~x279 & ~x418 & ~x461;
assign c8368 = ~x83 & ~x164 & ~x165 & ~x219 & ~x220 & ~x226 & ~x278 & ~x306 & ~x333 & ~x402 & ~x430 & ~x457 & ~x471 & ~x485 & ~x527 & ~x529 & ~x541 & ~x569 & ~x606 & ~x611 & ~x634 & ~x660;
assign c8370 =  x300 &  x440 & ~x3 & ~x5 & ~x23 & ~x26 & ~x29 & ~x30 & ~x31 & ~x32 & ~x60 & ~x84 & ~x85 & ~x88 & ~x89 & ~x197 & ~x335 & ~x336 & ~x365 & ~x366 & ~x391 & ~x520 & ~x521 & ~x587 & ~x756;
assign c8372 =  x216 &  x300 &  x356 & ~x759;
assign c8374 =  x595 & ~x1 & ~x3 & ~x5 & ~x27 & ~x32 & ~x34 & ~x60 & ~x82 & ~x91 & ~x113 & ~x115 & ~x118 & ~x142 & ~x173 & ~x197 & ~x198 & ~x199 & ~x201 & ~x202 & ~x209 & ~x227 & ~x255 & ~x282 & ~x284 & ~x285 & ~x310 & ~x336 & ~x338 & ~x341 & ~x395 & ~x422 & ~x545 & ~x740 & ~x759 & ~x760 & ~x761 & ~x767;
assign c8376 = ~x2 & ~x27 & ~x77 & ~x81 & ~x103 & ~x131 & ~x132 & ~x135 & ~x138 & ~x161 & ~x191 & ~x193 & ~x221 & ~x222 & ~x246 & ~x273 & ~x277 & ~x305 & ~x384 & ~x386 & ~x412 & ~x433 & ~x460 & ~x488 & ~x515 & ~x572 & ~x714 & ~x741;
assign c8378 =  x709 & ~x28 & ~x55 & ~x147 & ~x166 & ~x218 & ~x414 & ~x415 & ~x470 & ~x498 & ~x499 & ~x603 & ~x626;
assign c8380 = ~x22 & ~x24 & ~x27 & ~x32 & ~x35 & ~x45 & ~x48 & ~x62 & ~x63 & ~x73 & ~x77 & ~x80 & ~x81 & ~x99 & ~x109 & ~x136 & ~x139 & ~x142 & ~x165 & ~x166 & ~x169 & ~x194 & ~x221 & ~x251 & ~x252 & ~x276 & ~x277 & ~x278 & ~x280 & ~x297 & ~x304 & ~x324 & ~x325 & ~x360 & ~x363 & ~x380 & ~x388 & ~x389 & ~x408 & ~x417 & ~x419 & ~x444 & ~x445 & ~x464 & ~x475 & ~x491 & ~x492 & ~x520 & ~x754 & ~x782;
assign c8382 =  x462 &  x490 &  x518 &  x743 & ~x24 & ~x26 & ~x28 & ~x52 & ~x56 & ~x59 & ~x60 & ~x86 & ~x138 & ~x160 & ~x166 & ~x171 & ~x192 & ~x250 & ~x274 & ~x275 & ~x279 & ~x281 & ~x303 & ~x331 & ~x334 & ~x359 & ~x364 & ~x392 & ~x393 & ~x414 & ~x445 & ~x451 & ~x452 & ~x453 & ~x454 & ~x475 & ~x498 & ~x499 & ~x510 & ~x527 & ~x529 & ~x531 & ~x534 & ~x535 & ~x536 & ~x554 & ~x556 & ~x580 & ~x581 & ~x584 & ~x605 & ~x612 & ~x632 & ~x670 & ~x672 & ~x727 & ~x729 & ~x730;
assign c8384 =  x317 &  x456 &  x484 &  x512 &  x568 & ~x2 & ~x6 & ~x28 & ~x56 & ~x59 & ~x63 & ~x89 & ~x110 & ~x137 & ~x145 & ~x279 & ~x395 & ~x518 & ~x545 & ~x732;
assign c8386 = ~x3 & ~x21 & ~x24 & ~x29 & ~x33 & ~x55 & ~x60 & ~x61 & ~x78 & ~x106 & ~x107 & ~x112 & ~x125 & ~x136 & ~x137 & ~x138 & ~x141 & ~x146 & ~x166 & ~x173 & ~x192 & ~x193 & ~x223 & ~x224 & ~x246 & ~x281 & ~x308 & ~x337 & ~x339 & ~x366 & ~x452 & ~x472 & ~x501 & ~x605 & ~x611 & ~x630 & ~x656 & ~x671 & ~x684 & ~x688 & ~x697 & ~x728;
assign c8388 =  x15 &  x433 & ~x137 & ~x143 & ~x147 & ~x149 & ~x175 & ~x232 & ~x233 & ~x259 & ~x288 & ~x309 & ~x366 & ~x393 & ~x399 & ~x421 & ~x451 & ~x502 & ~x588;
assign c8390 =  x290 & ~x22 & ~x27 & ~x57 & ~x59 & ~x61 & ~x82 & ~x87 & ~x108 & ~x112 & ~x143 & ~x168 & ~x222 & ~x277 & ~x278 & ~x307 & ~x419 & ~x435 & ~x446 & ~x462 & ~x490 & ~x545 & ~x573 & ~x575 & ~x603 & ~x629 & ~x700 & ~x728 & ~x749;
assign c8392 =  x479 & ~x114 & ~x164 & ~x170 & ~x246 & ~x302 & ~x307 & ~x358 & ~x386 & ~x600;
assign c8394 =  x376 & ~x0 & ~x7 & ~x25 & ~x28 & ~x51 & ~x52 & ~x53 & ~x61 & ~x76 & ~x77 & ~x78 & ~x133 & ~x140 & ~x149 & ~x171 & ~x195 & ~x198 & ~x199 & ~x206 & ~x223 & ~x225 & ~x232 & ~x234 & ~x250 & ~x255 & ~x256 & ~x262 & ~x306 & ~x310 & ~x333 & ~x344 & ~x345 & ~x346 & ~x361 & ~x393 & ~x419 & ~x421 & ~x477 & ~x758;
assign c8396 =  x619 & ~x3 & ~x19 & ~x22 & ~x27 & ~x29 & ~x49 & ~x110 & ~x114 & ~x140 & ~x165 & ~x188 & ~x217 & ~x224 & ~x272 & ~x279 & ~x307 & ~x357 & ~x393 & ~x441 & ~x775;
assign c8398 = ~x18 & ~x30 & ~x35 & ~x53 & ~x60 & ~x64 & ~x75 & ~x79 & ~x90 & ~x140 & ~x144 & ~x155 & ~x167 & ~x168 & ~x195 & ~x198 & ~x199 & ~x252 & ~x278 & ~x279 & ~x324 & ~x335 & ~x417 & ~x434 & ~x448 & ~x462 & ~x504 & ~x759 & ~x771;
assign c8400 = ~x2 & ~x3 & ~x22 & ~x24 & ~x25 & ~x55 & ~x82 & ~x86 & ~x87 & ~x104 & ~x108 & ~x110 & ~x111 & ~x112 & ~x114 & ~x134 & ~x135 & ~x136 & ~x139 & ~x142 & ~x161 & ~x163 & ~x166 & ~x169 & ~x170 & ~x190 & ~x220 & ~x221 & ~x223 & ~x225 & ~x227 & ~x246 & ~x251 & ~x276 & ~x279 & ~x281 & ~x283 & ~x304 & ~x308 & ~x330 & ~x331 & ~x336 & ~x338 & ~x361 & ~x363 & ~x366 & ~x367 & ~x387 & ~x389 & ~x393 & ~x399 & ~x418 & ~x419 & ~x421 & ~x425 & ~x447 & ~x470 & ~x474 & ~x478 & ~x498 & ~x500 & ~x501 & ~x503 & ~x521 & ~x522 & ~x523 & ~x524 & ~x525 & ~x531 & ~x549 & ~x550 & ~x556 & ~x557 & ~x558 & ~x559 & ~x560 & ~x573 & ~x574 & ~x576 & ~x583 & ~x585 & ~x599 & ~x600 & ~x601 & ~x611 & ~x673 & ~x698 & ~x725 & ~x731 & ~x756 & ~x757 & ~x761 & ~x781;
assign c8402 =  x347 &  x457 & ~x27 & ~x30 & ~x86 & ~x113 & ~x114 & ~x175 & ~x201 & ~x256 & ~x343 & ~x369 & ~x393 & ~x453 & ~x454 & ~x747;
assign c8404 =  x511 & ~x34 & ~x56 & ~x62 & ~x82 & ~x84 & ~x85 & ~x86 & ~x89 & ~x110 & ~x115 & ~x142 & ~x169 & ~x200 & ~x201 & ~x281 & ~x335 & ~x396 & ~x423 & ~x448 & ~x450 & ~x515 & ~x518 & ~x519 & ~x543 & ~x547 & ~x600 & ~x602 & ~x759 & ~x768;
assign c8406 =  x343 &  x511 &  x539 & ~x0 & ~x3 & ~x26 & ~x31 & ~x32 & ~x33 & ~x56 & ~x60 & ~x89 & ~x111 & ~x113 & ~x141 & ~x145 & ~x166 & ~x173 & ~x197 & ~x338 & ~x365 & ~x366 & ~x391 & ~x462 & ~x488 & ~x543 & ~x600 & ~x626 & ~x627 & ~x655;
assign c8408 =  x187 & ~x5 & ~x24 & ~x27 & ~x54 & ~x60 & ~x82 & ~x83 & ~x84 & ~x86 & ~x87 & ~x89 & ~x113 & ~x144 & ~x169 & ~x172 & ~x196 & ~x197 & ~x223 & ~x226 & ~x227 & ~x254 & ~x277 & ~x278 & ~x279 & ~x307 & ~x359 & ~x360 & ~x361 & ~x365 & ~x389 & ~x390 & ~x393 & ~x416 & ~x417 & ~x418 & ~x419 & ~x422 & ~x445 & ~x446 & ~x548 & ~x559 & ~x573 & ~x575 & ~x671 & ~x698 & ~x699 & ~x732 & ~x775;
assign c8410 =  x128 &  x184 &  x240 &  x268 &  x296 &  x380 & ~x54 & ~x55 & ~x62 & ~x83 & ~x86 & ~x104 & ~x118 & ~x139 & ~x167 & ~x195 & ~x218 & ~x228 & ~x247 & ~x255 & ~x256 & ~x274 & ~x328 & ~x330 & ~x337 & ~x356 & ~x361 & ~x367 & ~x387 & ~x393 & ~x440 & ~x441 & ~x474 & ~x526 & ~x614 & ~x731 & ~x756;
assign c8412 = ~x1 & ~x6 & ~x7 & ~x27 & ~x30 & ~x33 & ~x34 & ~x36 & ~x54 & ~x59 & ~x78 & ~x81 & ~x83 & ~x88 & ~x90 & ~x108 & ~x118 & ~x137 & ~x138 & ~x139 & ~x143 & ~x166 & ~x167 & ~x192 & ~x196 & ~x201 & ~x202 & ~x203 & ~x231 & ~x249 & ~x256 & ~x281 & ~x282 & ~x286 & ~x303 & ~x307 & ~x311 & ~x313 & ~x314 & ~x335 & ~x338 & ~x366 & ~x370 & ~x388 & ~x392 & ~x394 & ~x398 & ~x419 & ~x425 & ~x426 & ~x445 & ~x447 & ~x452 & ~x473 & ~x530 & ~x532 & ~x534 & ~x549 & ~x551 & ~x552 & ~x556 & ~x560 & ~x562 & ~x577 & ~x589 & ~x603 & ~x604 & ~x619 & ~x628 & ~x629 & ~x642 & ~x644 & ~x671 & ~x672 & ~x723 & ~x725 & ~x728 & ~x754 & ~x761;
assign c8414 = ~x1 & ~x20 & ~x25 & ~x26 & ~x28 & ~x79 & ~x86 & ~x107 & ~x134 & ~x137 & ~x162 & ~x163 & ~x164 & ~x190 & ~x194 & ~x248 & ~x304 & ~x337 & ~x360 & ~x363 & ~x385 & ~x388 & ~x413 & ~x486 & ~x488 & ~x542 & ~x572 & ~x768 & ~x773;
assign c8416 =  x481 & ~x28 & ~x47 & ~x84 & ~x85 & ~x106 & ~x107 & ~x135 & ~x142 & ~x161 & ~x219 & ~x245 & ~x246 & ~x274 & ~x275 & ~x302 & ~x307 & ~x330 & ~x334 & ~x335 & ~x360 & ~x386 & ~x388 & ~x418 & ~x442 & ~x444 & ~x470 & ~x472 & ~x570 & ~x597 & ~x626;
assign c8418 = ~x0 & ~x1 & ~x6 & ~x13 & ~x17 & ~x25 & ~x33 & ~x40 & ~x44 & ~x52 & ~x57 & ~x76 & ~x79 & ~x114 & ~x139 & ~x151 & ~x164 & ~x192 & ~x196 & ~x222 & ~x224 & ~x251 & ~x279 & ~x303 & ~x304 & ~x331 & ~x360 & ~x364 & ~x387 & ~x430 & ~x457 & ~x671 & ~x674 & ~x700 & ~x736 & ~x737 & ~x753 & ~x756 & ~x759 & ~x764 & ~x781;
assign c8420 = ~x0 & ~x15 & ~x52 & ~x71 & ~x77 & ~x78 & ~x85 & ~x87 & ~x105 & ~x110 & ~x135 & ~x137 & ~x138 & ~x139 & ~x141 & ~x162 & ~x163 & ~x195 & ~x220 & ~x247 & ~x249 & ~x278 & ~x279 & ~x305 & ~x332 & ~x357 & ~x359 & ~x384 & ~x487 & ~x616 & ~x643 & ~x670 & ~x690 & ~x711 & ~x731;
assign c8422 =  x212 &  x296 &  x324 &  x436 & ~x48 & ~x105 & ~x166 & ~x189 & ~x214 & ~x242 & ~x249 & ~x270 & ~x271 & ~x298 & ~x327 & ~x356 & ~x415 & ~x441 & ~x442;
assign c8424 =  x451 & ~x52 & ~x135 & ~x191 & ~x303 & ~x306 & ~x332 & ~x414 & ~x695;
assign c8426 =  x483 &  x567 & ~x3 & ~x26 & ~x31 & ~x32 & ~x51 & ~x53 & ~x89 & ~x110 & ~x137 & ~x142 & ~x173 & ~x306 & ~x364 & ~x393 & ~x418 & ~x488 & ~x489 & ~x544 & ~x732 & ~x757 & ~x774;
assign c8428 =  x505 & ~x337 & ~x402 & ~x430 & ~x514 & ~x569;
assign c8430 =  x120 &  x399 & ~x15 & ~x179 & ~x206 & ~x226 & ~x520 & ~x543;
assign c8432 =  x322 &  x378 &  x486 & ~x54 & ~x79 & ~x83 & ~x88 & ~x89 & ~x137 & ~x140 & ~x144 & ~x165 & ~x168 & ~x217 & ~x222 & ~x225 & ~x258 & ~x285 & ~x308 & ~x336 & ~x363 & ~x365 & ~x393 & ~x415 & ~x421 & ~x423 & ~x424 & ~x426 & ~x452 & ~x499 & ~x505 & ~x526 & ~x530 & ~x558 & ~x755 & ~x756;
assign c8434 =  x15 &  x405 & ~x48 & ~x59 & ~x92 & ~x117 & ~x118 & ~x138 & ~x168 & ~x173 & ~x175 & ~x189 & ~x224 & ~x257 & ~x259 & ~x277 & ~x287 & ~x341 & ~x371 & ~x397 & ~x472 & ~x506 & ~x560 & ~x561 & ~x700;
assign c8436 =  x590 & ~x53 & ~x80 & ~x165 & ~x192 & ~x277 & ~x280 & ~x281 & ~x308 & ~x333 & ~x361 & ~x363 & ~x392 & ~x418 & ~x420 & ~x444 & ~x445 & ~x446 & ~x730 & ~x748;
assign c8438 = ~x50 & ~x52 & ~x85 & ~x108 & ~x110 & ~x112 & ~x134 & ~x136 & ~x137 & ~x164 & ~x166 & ~x168 & ~x172 & ~x218 & ~x222 & ~x230 & ~x249 & ~x259 & ~x280 & ~x282 & ~x286 & ~x306 & ~x309 & ~x311 & ~x334 & ~x359 & ~x361 & ~x365 & ~x388 & ~x392 & ~x394 & ~x395 & ~x419 & ~x423 & ~x426 & ~x448 & ~x477 & ~x501 & ~x605 & ~x608 & ~x633 & ~x658 & ~x659 & ~x669 & ~x671 & ~x683 & ~x699 & ~x727 & ~x781 & ~x783;
assign c8440 =  x428 &  x652 & ~x1 & ~x2 & ~x24 & ~x25 & ~x31 & ~x55 & ~x60 & ~x82 & ~x83 & ~x85 & ~x87 & ~x112 & ~x113 & ~x114 & ~x115 & ~x116 & ~x141 & ~x143 & ~x145 & ~x170 & ~x197 & ~x198 & ~x223 & ~x224 & ~x225 & ~x252 & ~x281 & ~x308 & ~x309 & ~x393 & ~x420 & ~x492 & ~x516 & ~x545 & ~x548 & ~x572 & ~x600 & ~x628 & ~x657 & ~x699 & ~x755 & ~x759 & ~x760;
assign c8442 =  x463 &  x517 &  x743 & ~x58 & ~x86 & ~x109 & ~x113 & ~x135 & ~x144 & ~x165 & ~x170 & ~x197 & ~x220 & ~x222 & ~x246 & ~x249 & ~x278 & ~x285 & ~x391 & ~x414 & ~x427 & ~x443 & ~x470 & ~x479 & ~x481 & ~x508 & ~x527 & ~x531 & ~x534 & ~x552 & ~x553 & ~x562 & ~x589 & ~x606 & ~x608 & ~x632 & ~x633;
assign c8444 =  x406 &  x434 & ~x53 & ~x114 & ~x115 & ~x140 & ~x142 & ~x166 & ~x172 & ~x173 & ~x196 & ~x199 & ~x224 & ~x228 & ~x247 & ~x258 & ~x275 & ~x277 & ~x278 & ~x303 & ~x306 & ~x311 & ~x334 & ~x341 & ~x359 & ~x392 & ~x394 & ~x397 & ~x424 & ~x426 & ~x448 & ~x453 & ~x500 & ~x561 & ~x590 & ~x605 & ~x607 & ~x632 & ~x635 & ~x657 & ~x658 & ~x729;
assign c8446 =  x351 &  x465 &  x709 &  x737 & ~x277 & ~x524;
assign c8448 =  x480 & ~x44 & ~x47 & ~x56 & ~x82 & ~x106 & ~x137 & ~x165 & ~x166 & ~x170 & ~x220 & ~x276 & ~x281 & ~x307 & ~x360 & ~x361 & ~x387 & ~x420 & ~x445 & ~x569 & ~x783;
assign c8450 =  x616;
assign c8452 =  x564 & ~x24 & ~x25 & ~x48 & ~x49 & ~x51 & ~x77 & ~x78 & ~x85 & ~x105 & ~x106 & ~x108 & ~x109 & ~x133 & ~x135 & ~x136 & ~x137 & ~x139 & ~x161 & ~x166 & ~x190 & ~x192 & ~x219 & ~x223 & ~x247 & ~x248 & ~x302 & ~x307 & ~x330 & ~x332 & ~x360 & ~x499 & ~x541 & ~x570 & ~x626 & ~x783;
assign c8454 =  x456 &  x708 & ~x1 & ~x3 & ~x4 & ~x26 & ~x27 & ~x30 & ~x54 & ~x56 & ~x59 & ~x82 & ~x85 & ~x86 & ~x110 & ~x112 & ~x113 & ~x115 & ~x140 & ~x144 & ~x146 & ~x166 & ~x168 & ~x170 & ~x172 & ~x173 & ~x195 & ~x196 & ~x197 & ~x200 & ~x201 & ~x226 & ~x227 & ~x228 & ~x252 & ~x280 & ~x364 & ~x420 & ~x421 & ~x423 & ~x450 & ~x601;
assign c8456 =  x463 &  x516 & ~x6 & ~x22 & ~x23 & ~x26 & ~x32 & ~x49 & ~x58 & ~x77 & ~x78 & ~x80 & ~x85 & ~x108 & ~x109 & ~x111 & ~x112 & ~x117 & ~x135 & ~x137 & ~x141 & ~x167 & ~x170 & ~x172 & ~x174 & ~x175 & ~x191 & ~x195 & ~x196 & ~x197 & ~x198 & ~x200 & ~x219 & ~x222 & ~x228 & ~x230 & ~x246 & ~x247 & ~x248 & ~x255 & ~x256 & ~x278 & ~x284 & ~x305 & ~x309 & ~x312 & ~x333 & ~x334 & ~x367 & ~x386 & ~x387 & ~x416 & ~x417 & ~x418 & ~x419 & ~x420 & ~x426 & ~x445 & ~x449 & ~x451 & ~x472 & ~x480 & ~x500 & ~x504 & ~x510 & ~x527 & ~x530 & ~x537 & ~x550 & ~x551 & ~x552 & ~x554 & ~x556 & ~x558 & ~x560 & ~x563 & ~x577 & ~x578 & ~x579 & ~x580 & ~x581 & ~x582 & ~x583 & ~x591 & ~x610 & ~x611 & ~x618 & ~x619 & ~x668 & ~x672 & ~x695 & ~x727 & ~x757 & ~x783;
assign c8458 = ~x3 & ~x5 & ~x26 & ~x38 & ~x54 & ~x56 & ~x58 & ~x59 & ~x61 & ~x72 & ~x73 & ~x82 & ~x84 & ~x99 & ~x114 & ~x117 & ~x143 & ~x144 & ~x155 & ~x168 & ~x169 & ~x173 & ~x174 & ~x224 & ~x284 & ~x307 & ~x308 & ~x309 & ~x336 & ~x337 & ~x342 & ~x369 & ~x465 & ~x476 & ~x520 & ~x548 & ~x604 & ~x759;
assign c8460 =  x407 &  x435 & ~x0 & ~x3 & ~x6 & ~x19 & ~x23 & ~x25 & ~x26 & ~x50 & ~x52 & ~x55 & ~x80 & ~x83 & ~x85 & ~x87 & ~x106 & ~x110 & ~x130 & ~x131 & ~x133 & ~x136 & ~x137 & ~x138 & ~x139 & ~x142 & ~x159 & ~x160 & ~x161 & ~x162 & ~x164 & ~x168 & ~x170 & ~x187 & ~x188 & ~x189 & ~x190 & ~x191 & ~x193 & ~x197 & ~x214 & ~x216 & ~x217 & ~x219 & ~x220 & ~x225 & ~x243 & ~x249 & ~x270 & ~x271 & ~x272 & ~x273 & ~x275 & ~x280 & ~x281 & ~x298 & ~x302 & ~x305 & ~x307 & ~x326 & ~x328 & ~x357 & ~x384 & ~x385 & ~x387 & ~x391 & ~x412 & ~x441 & ~x446 & ~x502 & ~x530 & ~x553 & ~x613 & ~x668 & ~x697 & ~x698 & ~x726 & ~x759 & ~x780 & ~x781 & ~x783;
assign c8462 =  x539 & ~x1 & ~x22 & ~x31 & ~x56 & ~x77 & ~x107 & ~x137 & ~x165 & ~x166 & ~x192 & ~x220 & ~x221 & ~x282 & ~x307 & ~x333 & ~x363 & ~x365 & ~x389 & ~x416 & ~x491 & ~x546 & ~x548 & ~x642 & ~x643 & ~x746 & ~x769;
assign c8464 =  x745 & ~x51 & ~x52 & ~x80 & ~x146 & ~x163 & ~x165 & ~x168 & ~x170 & ~x196 & ~x197 & ~x231 & ~x253 & ~x254 & ~x277 & ~x281 & ~x316 & ~x332 & ~x360 & ~x361 & ~x365 & ~x387 & ~x417 & ~x473 & ~x474 & ~x484 & ~x525 & ~x527 & ~x528 & ~x530 & ~x539 & ~x581 & ~x588 & ~x605 & ~x606 & ~x612 & ~x632 & ~x640 & ~x675 & ~x702 & ~x752 & ~x753 & ~x758 & ~x783;
assign c8466 = ~x8 & ~x20 & ~x25 & ~x28 & ~x35 & ~x89 & ~x90 & ~x104 & ~x106 & ~x132 & ~x135 & ~x136 & ~x137 & ~x140 & ~x162 & ~x170 & ~x222 & ~x252 & ~x302 & ~x304 & ~x305 & ~x333 & ~x339 & ~x363 & ~x393 & ~x419 & ~x443 & ~x503 & ~x521 & ~x573 & ~x670 & ~x698 & ~x739 & ~x766 & ~x774 & ~x776;
assign c8468 =  x635 & ~x7 & ~x74 & ~x130 & ~x163 & ~x165 & ~x193 & ~x384 & ~x386 & ~x413 & ~x418 & ~x446 & ~x470 & ~x473 & ~x497 & ~x498 & ~x524 & ~x555 & ~x774 & ~x775;
assign c8470 =  x240 &  x352 &  x380 & ~x47 & ~x60 & ~x104 & ~x115 & ~x131 & ~x139 & ~x141 & ~x159 & ~x160 & ~x163 & ~x170 & ~x216 & ~x217 & ~x223 & ~x245 & ~x256 & ~x272 & ~x329 & ~x331 & ~x357 & ~x363 & ~x385 & ~x414 & ~x443 & ~x444 & ~x467 & ~x468 & ~x560 & ~x701 & ~x760;
assign c8472 =  x126 &  x154 &  x210 &  x322 &  x378 &  x406 &  x460 & ~x189 & ~x195 & ~x247 & ~x273 & ~x340 & ~x357 & ~x469 & ~x475 & ~x584;
assign c8474 =  x397 & ~x19 & ~x48 & ~x168 & ~x304 & ~x387 & ~x433 & ~x489 & ~x722 & ~x745 & ~x779;
assign c8476 =  x263 &  x453 &  x507 &  x562 & ~x80;
assign c8478 =  x454 &  x509 & ~x0 & ~x17 & ~x21 & ~x26 & ~x28 & ~x51 & ~x52 & ~x53 & ~x78 & ~x80 & ~x83 & ~x106 & ~x109 & ~x135 & ~x136 & ~x164 & ~x192 & ~x194 & ~x219 & ~x246 & ~x274 & ~x275 & ~x276 & ~x277 & ~x302 & ~x330 & ~x332 & ~x364 & ~x387 & ~x389 & ~x414 & ~x418 & ~x599;
assign c8480 = ~x0 & ~x3 & ~x7 & ~x8 & ~x23 & ~x34 & ~x54 & ~x56 & ~x57 & ~x62 & ~x82 & ~x89 & ~x90 & ~x91 & ~x109 & ~x114 & ~x116 & ~x118 & ~x145 & ~x166 & ~x168 & ~x170 & ~x173 & ~x174 & ~x195 & ~x222 & ~x224 & ~x257 & ~x258 & ~x259 & ~x278 & ~x283 & ~x285 & ~x286 & ~x314 & ~x339 & ~x341 & ~x368 & ~x394 & ~x410 & ~x422 & ~x437 & ~x448 & ~x450 & ~x451 & ~x464 & ~x465 & ~x474 & ~x478 & ~x493 & ~x519 & ~x573 & ~x642 & ~x760 & ~x762 & ~x767 & ~x779 & ~x783;
assign c8482 =  x320 &  x351 &  x458 & ~x34 & ~x106 & ~x163 & ~x193 & ~x220 & ~x225 & ~x341 & ~x343 & ~x369 & ~x504 & ~x532;
assign c8484 =  x538 & ~x55 & ~x56 & ~x71 & ~x73 & ~x110 & ~x167 & ~x275 & ~x279 & ~x361 & ~x443 & ~x712 & ~x717 & ~x738;
assign c8486 =  x207 &  x486 & ~x82 & ~x110 & ~x137 & ~x138 & ~x147 & ~x201 & ~x251 & ~x313 & ~x395 & ~x478 & ~x685;
assign c8488 = ~x16 & ~x18 & ~x19 & ~x21 & ~x44 & ~x48 & ~x49 & ~x52 & ~x72 & ~x74 & ~x79 & ~x80 & ~x84 & ~x101 & ~x106 & ~x108 & ~x112 & ~x113 & ~x114 & ~x129 & ~x135 & ~x136 & ~x137 & ~x142 & ~x158 & ~x164 & ~x167 & ~x188 & ~x191 & ~x194 & ~x216 & ~x223 & ~x243 & ~x244 & ~x247 & ~x248 & ~x249 & ~x250 & ~x251 & ~x275 & ~x276 & ~x278 & ~x299 & ~x300 & ~x302 & ~x303 & ~x304 & ~x329 & ~x332 & ~x333 & ~x355 & ~x356 & ~x383 & ~x387 & ~x390 & ~x411 & ~x419 & ~x439 & ~x530 & ~x555 & ~x579 & ~x581 & ~x724 & ~x730 & ~x749 & ~x754 & ~x758 & ~x762 & ~x779;
assign c8490 =  x660 &  x661 & ~x191 & ~x247 & ~x361 & ~x550 & ~x553 & ~x601;
assign c8492 =  x482 &  x565 &  x594 &  x650 & ~x1 & ~x27 & ~x30 & ~x32 & ~x43 & ~x84 & ~x125 & ~x152 & ~x170 & ~x179 & ~x199 & ~x225 & ~x282 & ~x364 & ~x365 & ~x489 & ~x542 & ~x731;
assign c8494 = ~x1 & ~x7 & ~x24 & ~x73 & ~x74 & ~x79 & ~x87 & ~x112 & ~x114 & ~x118 & ~x171 & ~x172 & ~x196 & ~x200 & ~x250 & ~x278 & ~x306 & ~x334 & ~x336 & ~x391 & ~x420 & ~x462 & ~x463 & ~x476 & ~x490 & ~x491 & ~x504 & ~x546 & ~x741 & ~x742 & ~x764;
assign c8496 =  x546 &  x739 &  x743 & ~x104 & ~x145 & ~x193 & ~x218 & ~x244 & ~x301 & ~x391 & ~x414 & ~x447 & ~x470 & ~x508 & ~x610 & ~x620 & ~x783;
assign c8498 =  x343 & ~x24 & ~x50 & ~x51 & ~x61 & ~x89 & ~x109 & ~x111 & ~x123 & ~x124 & ~x144 & ~x167 & ~x206 & ~x251 & ~x252 & ~x277 & ~x359 & ~x360 & ~x433 & ~x460 & ~x485 & ~x757;
assign c81 =  x363;
assign c83 = ~x1 & ~x20 & ~x54 & ~x114 & ~x163 & ~x215 & ~x217 & ~x253 & ~x307 & ~x334 & ~x360 & ~x361 & ~x393 & ~x449 & ~x475 & ~x519 & ~x630 & ~x641 & ~x647 & ~x660 & ~x672 & ~x723 & ~x777 & ~x781 & ~x782 & ~x783;
assign c85 =  x419;
assign c87 =  x184 & ~x419 & ~x424 & ~x475 & ~x624 & ~x682 & ~x735 & ~x738;
assign c89 =  x518 & ~x389 & ~x589 & ~x644 & ~x742 & ~x743 & ~x769 & ~x770;
assign c811 = ~x59 & ~x193 & ~x197 & ~x210 & ~x211 & ~x334 & ~x375 & ~x477 & ~x531 & ~x561 & ~x585 & ~x613 & ~x614 & ~x615 & ~x616 & ~x617 & ~x619 & ~x620 & ~x675 & ~x697 & ~x698 & ~x700 & ~x724 & ~x731 & ~x753 & ~x758;
assign c813 =  x192 & ~x359 & ~x417;
assign c815 = ~x145 & ~x173 & ~x197 & ~x254 & ~x510 & ~x532 & ~x569 & ~x626 & ~x653 & ~x710;
assign c817 = ~x2 & ~x28 & ~x56 & ~x87 & ~x98 & ~x112 & ~x197 & ~x252 & ~x304 & ~x332 & ~x339 & ~x365 & ~x366 & ~x367 & ~x368 & ~x451 & ~x505 & ~x507 & ~x516 & ~x591 & ~x643 & ~x645 & ~x646 & ~x647 & ~x665 & ~x670 & ~x672 & ~x699 & ~x724 & ~x729;
assign c819 =  x256 &  x311 & ~x425;
assign c821 =  x200 & ~x634;
assign c823 = ~x25 & ~x51 & ~x55 & ~x83 & ~x98 & ~x99 & ~x100 & ~x137 & ~x420 & ~x450 & ~x452 & ~x476 & ~x508 & ~x563 & ~x592 & ~x616 & ~x618 & ~x641 & ~x698 & ~x735 & ~x736 & ~x754 & ~x763 & ~x766;
assign c825 =  x548 &  x549 & ~x18 & ~x310 & ~x533 & ~x719 & ~x774;
assign c827 = ~x2 & ~x110 & ~x169 & ~x228 & ~x252 & ~x477 & ~x500 & ~x501 & ~x504 & ~x560 & ~x561 & ~x569 & ~x595 & ~x624 & ~x625 & ~x626 & ~x650 & ~x651 & ~x652 & ~x670 & ~x679 & ~x727 & ~x735 & ~x760;
assign c829 =  x285 & ~x371 & ~x398;
assign c831 =  x656 &  x684 & ~x16 & ~x368 & ~x386 & ~x561 & ~x563 & ~x607 & ~x618 & ~x619 & ~x635 & ~x729;
assign c833 = ~x308 & ~x351 & ~x480 & ~x530 & ~x564 & ~x592 & ~x653 & ~x737 & ~x752 & ~x764 & ~x766;
assign c835 = ~x57 & ~x166 & ~x223 & ~x394 & ~x439 & ~x468 & ~x477 & ~x496 & ~x504 & ~x526 & ~x532 & ~x542 & ~x596 & ~x623 & ~x625 & ~x679 & ~x681 & ~x708 & ~x740 & ~x761;
assign c837 =  x268 & ~x57 & ~x152 & ~x207 & ~x317 & ~x344 & ~x408 & ~x503;
assign c839 =  x338;
assign c841 =  x381 & ~x14 & ~x43 & ~x214 & ~x390 & ~x720 & ~x764;
assign c843 = ~x28 & ~x38 & ~x50 & ~x51 & ~x58 & ~x108 & ~x354 & ~x379 & ~x505 & ~x529 & ~x612 & ~x639 & ~x647 & ~x674 & ~x737;
assign c845 =  x345 & ~x187 & ~x505 & ~x512 & ~x513 & ~x561 & ~x590;
assign c847 =  x239 &  x657 &  x685 & ~x566 & ~x567;
assign c849 =  x469 &  x578;
assign c851 =  x96 & ~x216 & ~x242 & ~x585 & ~x647 & ~x662 & ~x674 & ~x701 & ~x720 & ~x761;
assign c853 =  x70 & ~x102 & ~x104 & ~x131 & ~x229 & ~x374 & ~x376 & ~x588 & ~x618 & ~x645 & ~x648 & ~x703;
assign c855 = ~x18 & ~x47 & ~x55 & ~x78 & ~x168 & ~x200 & ~x267 & ~x332 & ~x547 & ~x582 & ~x585 & ~x648 & ~x649 & ~x667 & ~x782;
assign c857 = ~x0 & ~x81 & ~x82 & ~x114 & ~x141 & ~x164 & ~x173 & ~x200 & ~x218 & ~x307 & ~x445 & ~x474 & ~x484 & ~x505 & ~x508 & ~x536 & ~x616 & ~x619 & ~x633 & ~x644 & ~x645 & ~x649 & ~x717 & ~x745 & ~x779;
assign c859 =  x205 &  x206 &  x207 & ~x20 & ~x32 & ~x47 & ~x73 & ~x166 & ~x252 & ~x614 & ~x647 & ~x673 & ~x728 & ~x730 & ~x756 & ~x758;
assign c861 =  x414 & ~x161 & ~x218 & ~x219 & ~x248 & ~x363 & ~x449 & ~x751;
assign c863 =  x100 & ~x65 & ~x66 & ~x352 & ~x506 & ~x588;
assign c865 = ~x20 & ~x55 & ~x118 & ~x166 & ~x195 & ~x223 & ~x256 & ~x363 & ~x367 & ~x390 & ~x420 & ~x449 & ~x450 & ~x479 & ~x529 & ~x598 & ~x625 & ~x653 & ~x679 & ~x682 & ~x738;
assign c867 = ~x425 & ~x443 & ~x480 & ~x570 & ~x596 & ~x626 & ~x654 & ~x682 & ~x706 & ~x707 & ~x736;
assign c869 =  x199;
assign c871 =  x656 & ~x9 & ~x54 & ~x55 & ~x77 & ~x145 & ~x256 & ~x313 & ~x530 & ~x534 & ~x560 & ~x635 & ~x643 & ~x644 & ~x701 & ~x727 & ~x732 & ~x758 & ~x761 & ~x781;
assign c873 =  x360 &  x396;
assign c875 =  x116;
assign c877 = ~x2 & ~x143 & ~x163 & ~x192 & ~x336 & ~x363 & ~x447 & ~x449 & ~x485 & ~x505 & ~x531 & ~x563 & ~x591 & ~x617 & ~x675 & ~x688 & ~x717 & ~x723 & ~x751 & ~x772 & ~x774 & ~x783;
assign c879 =  x362;
assign c881 =  x98 &  x627 &  x655 & ~x329 & ~x607;
assign c883 =  x182 & ~x17 & ~x287 & ~x458 & ~x459 & ~x732 & ~x750;
assign c885 =  x404 & ~x71 & ~x536 & ~x562 & ~x591 & ~x617 & ~x646 & ~x764 & ~x766;
assign c887 =  x356 & ~x5 & ~x17 & ~x72 & ~x188 & ~x189 & ~x215 & ~x217 & ~x251 & ~x253 & ~x335 & ~x700 & ~x730 & ~x754 & ~x757 & ~x781;
assign c889 =  x455 & ~x541 & ~x569 & ~x595 & ~x596 & ~x622 & ~x623 & ~x677 & ~x678 & ~x707 & ~x732 & ~x733 & ~x735 & ~x783;
assign c891 =  x134 & ~x274 & ~x301;
assign c893 =  x127 & ~x431 & ~x434 & ~x532 & ~x535 & ~x669;
assign c895 = ~x81 & ~x107 & ~x339 & ~x511 & ~x541 & ~x566 & ~x567 & ~x624 & ~x649 & ~x675 & ~x722 & ~x727 & ~x744 & ~x753;
assign c897 = ~x6 & ~x56 & ~x165 & ~x168 & ~x187 & ~x214 & ~x216 & ~x222 & ~x253 & ~x254 & ~x392 & ~x473 & ~x476 & ~x507 & ~x531 & ~x532 & ~x533 & ~x557 & ~x563 & ~x588 & ~x589 & ~x592 & ~x601 & ~x602 & ~x619 & ~x629 & ~x637 & ~x639 & ~x646 & ~x647 & ~x665 & ~x666 & ~x673 & ~x692 & ~x701 & ~x702 & ~x722 & ~x749 & ~x751;
assign c899 =  x238 &  x242 & ~x223 & ~x326;
assign c8101 =  x655 &  x683 &  x684 &  x712 &  x741 & ~x5 & ~x82 & ~x107 & ~x311 & ~x706 & ~x760;
assign c8103 = ~x0 & ~x18 & ~x19 & ~x20 & ~x24 & ~x25 & ~x29 & ~x32 & ~x35 & ~x51 & ~x54 & ~x58 & ~x79 & ~x83 & ~x86 & ~x89 & ~x113 & ~x140 & ~x141 & ~x143 & ~x170 & ~x172 & ~x195 & ~x196 & ~x197 & ~x218 & ~x219 & ~x250 & ~x277 & ~x283 & ~x304 & ~x306 & ~x308 & ~x309 & ~x332 & ~x394 & ~x414 & ~x422 & ~x450 & ~x476 & ~x479 & ~x505 & ~x506 & ~x529 & ~x555 & ~x557 & ~x560 & ~x562 & ~x584 & ~x585 & ~x586 & ~x590 & ~x611 & ~x614 & ~x615 & ~x618 & ~x619 & ~x620 & ~x639 & ~x642 & ~x645 & ~x648 & ~x667 & ~x669 & ~x671 & ~x676 & ~x695 & ~x712 & ~x724 & ~x726 & ~x729 & ~x739 & ~x740 & ~x752 & ~x767 & ~x768 & ~x769 & ~x779 & ~x781;
assign c8105 =  x175 & ~x42 & ~x453 & ~x735;
assign c8107 =  x206 &  x546 &  x601 & ~x15 & ~x55;
assign c8109 = ~x51 & ~x115 & ~x200 & ~x368 & ~x403 & ~x431 & ~x433 & ~x477 & ~x479 & ~x505 & ~x508 & ~x528 & ~x535 & ~x536 & ~x561 & ~x563 & ~x646 & ~x667 & ~x669 & ~x671 & ~x675 & ~x728 & ~x729;
assign c8111 =  x522 & ~x26 & ~x457 & ~x505 & ~x534 & ~x561 & ~x562 & ~x747 & ~x753;
assign c8113 =  x335;
assign c8115 =  x175 & ~x14 & ~x266 & ~x369;
assign c8117 = ~x2 & ~x4 & ~x5 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x26 & ~x28 & ~x29 & ~x30 & ~x31 & ~x33 & ~x34 & ~x52 & ~x53 & ~x55 & ~x56 & ~x57 & ~x58 & ~x59 & ~x80 & ~x82 & ~x83 & ~x84 & ~x86 & ~x88 & ~x110 & ~x111 & ~x112 & ~x113 & ~x114 & ~x115 & ~x116 & ~x137 & ~x138 & ~x140 & ~x142 & ~x143 & ~x165 & ~x166 & ~x167 & ~x168 & ~x170 & ~x171 & ~x172 & ~x196 & ~x222 & ~x223 & ~x224 & ~x250 & ~x253 & ~x277 & ~x280 & ~x307 & ~x308 & ~x309 & ~x332 & ~x333 & ~x335 & ~x338 & ~x360 & ~x361 & ~x362 & ~x363 & ~x364 & ~x365 & ~x367 & ~x389 & ~x391 & ~x393 & ~x394 & ~x417 & ~x419 & ~x420 & ~x421 & ~x422 & ~x446 & ~x449 & ~x450 & ~x475 & ~x476 & ~x477 & ~x478 & ~x502 & ~x503 & ~x504 & ~x505 & ~x506 & ~x529 & ~x530 & ~x531 & ~x532 & ~x533 & ~x558 & ~x559 & ~x560 & ~x561 & ~x562 & ~x586 & ~x588 & ~x590 & ~x600 & ~x614 & ~x615 & ~x616 & ~x617 & ~x618 & ~x627 & ~x642 & ~x643 & ~x644 & ~x645 & ~x646 & ~x669 & ~x670 & ~x671 & ~x673 & ~x674 & ~x687 & ~x697 & ~x698 & ~x699 & ~x700 & ~x701 & ~x726 & ~x727 & ~x728 & ~x737 & ~x738 & ~x752 & ~x753 & ~x754 & ~x756 & ~x763 & ~x780;
assign c8119 = ~x342 & ~x365 & ~x457 & ~x477 & ~x486 & ~x515 & ~x536 & ~x537 & ~x540 & ~x567;
assign c8121 = ~x1 & ~x6 & ~x135 & ~x197 & ~x308 & ~x337 & ~x477 & ~x514 & ~x568 & ~x569 & ~x594 & ~x598 & ~x600 & ~x623 & ~x643 & ~x649 & ~x727 & ~x731 & ~x732;
assign c8123 =  x445;
assign c8125 =  x284 & ~x95 & ~x425;
assign c8127 =  x245 & ~x328 & ~x329;
assign c8129 =  x363;
assign c8131 =  x260 &  x487 & ~x346 & ~x374 & ~x764;
assign c8133 = ~x0 & ~x2 & ~x24 & ~x25 & ~x28 & ~x30 & ~x31 & ~x53 & ~x54 & ~x55 & ~x59 & ~x61 & ~x80 & ~x84 & ~x85 & ~x86 & ~x87 & ~x88 & ~x109 & ~x114 & ~x138 & ~x140 & ~x141 & ~x143 & ~x169 & ~x170 & ~x224 & ~x252 & ~x309 & ~x310 & ~x316 & ~x337 & ~x364 & ~x365 & ~x367 & ~x388 & ~x389 & ~x390 & ~x393 & ~x416 & ~x420 & ~x421 & ~x431 & ~x432 & ~x433 & ~x445 & ~x447 & ~x449 & ~x459 & ~x460 & ~x461 & ~x462 & ~x473 & ~x476 & ~x477 & ~x501 & ~x503 & ~x504 & ~x505 & ~x529 & ~x531 & ~x533 & ~x560 & ~x561 & ~x590 & ~x615 & ~x617 & ~x641 & ~x644 & ~x645 & ~x670 & ~x672 & ~x697 & ~x726 & ~x727 & ~x730 & ~x753 & ~x754 & ~x755 & ~x757 & ~x781 & ~x783;
assign c8135 = ~x20 & ~x58 & ~x102 & ~x132 & ~x134 & ~x138 & ~x171 & ~x211 & ~x213 & ~x214 & ~x280 & ~x476 & ~x478 & ~x556 & ~x604 & ~x674 & ~x675 & ~x676 & ~x694 & ~x704 & ~x733 & ~x760 & ~x764;
assign c8137 =  x384 & ~x130 & ~x245 & ~x560 & ~x621 & ~x649;
assign c8139 =  x136;
assign c8141 =  x712 & ~x16 & ~x102 & ~x251 & ~x336 & ~x533 & ~x601 & ~x640 & ~x663 & ~x666 & ~x700 & ~x722;
assign c8143 = ~x213 & ~x269 & ~x396 & ~x561 & ~x564 & ~x582 & ~x592 & ~x601 & ~x731 & ~x755;
assign c8145 =  x171 & ~x693;
assign c8147 =  x68 &  x353 & ~x241;
assign c8149 =  x352 &  x467 & ~x445 & ~x475 & ~x720;
assign c8151 = ~x24 & ~x31 & ~x52 & ~x86 & ~x110 & ~x195 & ~x220 & ~x248 & ~x366 & ~x368 & ~x477 & ~x479 & ~x483 & ~x487 & ~x489 & ~x506 & ~x511 & ~x643 & ~x699 & ~x721 & ~x780;
assign c8153 =  x501 &  x572;
assign c8155 = ~x9 & ~x52 & ~x55 & ~x112 & ~x203 & ~x281 & ~x336 & ~x367 & ~x451 & ~x478 & ~x570 & ~x595 & ~x596 & ~x598 & ~x623 & ~x672 & ~x727 & ~x750 & ~x756 & ~x770;
assign c8157 = ~x1 & ~x33 & ~x56 & ~x58 & ~x84 & ~x141 & ~x171 & ~x172 & ~x249 & ~x280 & ~x420 & ~x455 & ~x483 & ~x485 & ~x488 & ~x489 & ~x562 & ~x592 & ~x614 & ~x669 & ~x699 & ~x702 & ~x759 & ~x782 & ~x783;
assign c8159 =  x263 &  x491 &  x575 & ~x614;
assign c8161 =  x359 & ~x135 & ~x191;
assign c8163 =  x241 & ~x292 & ~x344 & ~x374 & ~x402 & ~x436;
assign c8165 =  x370 & ~x28 & ~x55 & ~x73 & ~x110 & ~x111 & ~x140 & ~x144 & ~x165 & ~x195 & ~x227 & ~x255 & ~x282 & ~x309 & ~x310 & ~x312 & ~x338 & ~x364 & ~x450 & ~x501 & ~x504 & ~x505 & ~x506 & ~x533 & ~x561 & ~x562 & ~x586 & ~x589 & ~x613 & ~x616 & ~x617 & ~x618 & ~x643 & ~x645 & ~x646 & ~x647 & ~x671 & ~x674 & ~x702 & ~x756 & ~x758;
assign c8167 =  x278;
assign c8169 =  x96 & ~x214 & ~x279 & ~x396 & ~x556 & ~x603 & ~x611 & ~x647 & ~x696 & ~x698;
assign c8171 = ~x0 & ~x2 & ~x6 & ~x27 & ~x57 & ~x82 & ~x113 & ~x114 & ~x115 & ~x170 & ~x249 & ~x305 & ~x366 & ~x388 & ~x391 & ~x415 & ~x417 & ~x419 & ~x442 & ~x446 & ~x448 & ~x504 & ~x528 & ~x533 & ~x534 & ~x559 & ~x573 & ~x588 & ~x633 & ~x643 & ~x645 & ~x661 & ~x662 & ~x663 & ~x664 & ~x720 & ~x724 & ~x752 & ~x763 & ~x764 & ~x781;
assign c8173 = ~x58 & ~x250 & ~x340 & ~x498 & ~x533 & ~x563 & ~x582 & ~x583 & ~x626 & ~x646 & ~x653 & ~x670 & ~x674 & ~x681 & ~x682 & ~x708 & ~x709 & ~x710 & ~x726 & ~x735 & ~x754 & ~x781;
assign c8175 =  x575 &  x603 &  x632 & ~x565;
assign c8177 = ~x19 & ~x20 & ~x53 & ~x163 & ~x442 & ~x492 & ~x499 & ~x578 & ~x580 & ~x582 & ~x681 & ~x725 & ~x736 & ~x758 & ~x779;
assign c8179 =  x329 & ~x25 & ~x43 & ~x110 & ~x162 & ~x188 & ~x189 & ~x191 & ~x392 & ~x763;
assign c8181 =  x173 &  x650 & ~x509;
assign c8183 =  x334;
assign c8185 = ~x2 & ~x21 & ~x54 & ~x111 & ~x136 & ~x138 & ~x306 & ~x450 & ~x473 & ~x504 & ~x506 & ~x533 & ~x559 & ~x560 & ~x571 & ~x598 & ~x625 & ~x626 & ~x651 & ~x652 & ~x706 & ~x707 & ~x709 & ~x726 & ~x733 & ~x734 & ~x735 & ~x736 & ~x753 & ~x754 & ~x761 & ~x764;
assign c8187 =  x711 & ~x26 & ~x28 & ~x114 & ~x166 & ~x215 & ~x391 & ~x562 & ~x675 & ~x690 & ~x692 & ~x703 & ~x720 & ~x776;
assign c8189 =  x602 &  x630 &  x657 & ~x769;
assign c8191 = ~x1 & ~x29 & ~x200 & ~x212 & ~x213 & ~x309 & ~x312 & ~x339 & ~x421 & ~x505 & ~x622 & ~x629 & ~x707 & ~x733;
assign c8193 =  x87;
assign c8195 =  x417 & ~x247;
assign c8197 =  x577 & ~x17 & ~x112 & ~x485 & ~x536;
assign c8199 =  x574 & ~x484 & ~x538 & ~x744;
assign c8201 =  x298 & ~x159 & ~x401 & ~x430 & ~x432 & ~x533 & ~x588 & ~x749;
assign c8203 =  x386 & ~x105 & ~x161 & ~x162 & ~x752 & ~x778;
assign c8205 =  x327 & ~x17 & ~x28 & ~x216 & ~x225 & ~x243 & ~x250 & ~x252 & ~x419 & ~x698 & ~x699 & ~x728 & ~x748 & ~x752 & ~x753 & ~x756;
assign c8207 =  x418;
assign c8209 =  x138;
assign c8211 = ~x4 & ~x110 & ~x227 & ~x252 & ~x453 & ~x487 & ~x489 & ~x539 & ~x540 & ~x568;
assign c8213 = ~x7 & ~x34 & ~x82 & ~x161 & ~x173 & ~x192 & ~x196 & ~x220 & ~x308 & ~x339 & ~x365 & ~x416 & ~x449 & ~x451 & ~x477 & ~x535 & ~x558 & ~x561 & ~x619 & ~x666 & ~x674 & ~x716 & ~x725 & ~x773;
assign c8215 =  x367;
assign c8217 = ~x252 & ~x440 & ~x468 & ~x526 & ~x551 & ~x570 & ~x580 & ~x651 & ~x670 & ~x696 & ~x704 & ~x726 & ~x727 & ~x733 & ~x772;
assign c8219 = ~x1 & ~x9 & ~x25 & ~x29 & ~x85 & ~x138 & ~x169 & ~x225 & ~x278 & ~x280 & ~x283 & ~x304 & ~x305 & ~x332 & ~x333 & ~x338 & ~x345 & ~x360 & ~x363 & ~x374 & ~x394 & ~x395 & ~x402 & ~x420 & ~x421 & ~x450 & ~x478 & ~x479 & ~x503 & ~x504 & ~x520 & ~x530 & ~x560 & ~x588 & ~x590 & ~x591 & ~x604 & ~x612 & ~x616 & ~x618 & ~x644 & ~x647 & ~x702 & ~x704 & ~x726 & ~x729 & ~x754 & ~x756;
assign c8221 =  x660 & ~x516 & ~x537 & ~x538 & ~x566 & ~x568;
assign c8223 =  x199;
assign c8225 = ~x10 & ~x19 & ~x57 & ~x201 & ~x254 & ~x352 & ~x354 & ~x368 & ~x395 & ~x556 & ~x611 & ~x648 & ~x721;
assign c8227 = ~x53 & ~x112 & ~x192 & ~x200 & ~x201 & ~x216 & ~x225 & ~x249 & ~x276 & ~x307 & ~x311 & ~x447 & ~x475 & ~x502 & ~x505 & ~x528 & ~x530 & ~x573 & ~x601 & ~x614 & ~x619 & ~x636 & ~x645 & ~x647 & ~x698 & ~x720 & ~x729 & ~x731 & ~x776 & ~x783;
assign c8229 =  x445 & ~x650;
assign c8231 = ~x10 & ~x91 & ~x102 & ~x132 & ~x134 & ~x135 & ~x540 & ~x541 & ~x552 & ~x594 & ~x595 & ~x621 & ~x623 & ~x625 & ~x650 & ~x675 & ~x679 & ~x695 & ~x704 & ~x705 & ~x727 & ~x772;
assign c8233 =  x467 & ~x26 & ~x225 & ~x419 & ~x429 & ~x533 & ~x644 & ~x719;
assign c8235 =  x462;
assign c8237 =  x390;
assign c8239 =  x245 & ~x306 & ~x445 & ~x477 & ~x478 & ~x501 & ~x505 & ~x531 & ~x532 & ~x618 & ~x647 & ~x698 & ~x760;
assign c8241 =  x109;
assign c8243 =  x712 & ~x159 & ~x546 & ~x674;
assign c8245 =  x473 & ~x219 & ~x292 & ~x293 & ~x608;
assign c8247 = ~x0 & ~x1 & ~x194 & ~x221 & ~x228 & ~x254 & ~x325 & ~x326 & ~x394 & ~x419 & ~x449 & ~x477 & ~x576 & ~x583 & ~x668 & ~x707 & ~x766 & ~x781;
assign c8249 =  x288 &  x515 & ~x374;
assign c8251 =  x554 &  x582;
assign c8253 =  x126 & ~x257 & ~x431 & ~x432 & ~x479;
assign c8255 =  x361;
assign c8257 =  x215 &  x548 & ~x75;
assign c8259 =  x630 &  x686 & ~x92 & ~x633;
assign c8261 =  x361;
assign c8263 =  x127 &  x545 & ~x492;
assign c8265 =  x573 &  x628 & ~x697 & ~x741;
assign c8267 = ~x28 & ~x82 & ~x262 & ~x290 & ~x345 & ~x394 & ~x407 & ~x428 & ~x456 & ~x484 & ~x489 & ~x504 & ~x505 & ~x533 & ~x641 & ~x700 & ~x726;
assign c8269 = ~x24 & ~x108 & ~x280 & ~x281 & ~x284 & ~x403 & ~x405 & ~x420 & ~x458 & ~x461 & ~x475 & ~x476 & ~x531 & ~x533 & ~x534 & ~x559 & ~x619 & ~x669 & ~x674 & ~x755;
assign c8271 =  x521 &  x550 & ~x59 & ~x74 & ~x85 & ~x334 & ~x335 & ~x362 & ~x532 & ~x561 & ~x589;
assign c8273 = ~x79 & ~x168 & ~x184 & ~x186 & ~x212 & ~x216 & ~x244 & ~x273 & ~x294 & ~x301 & ~x392 & ~x420 & ~x667 & ~x669 & ~x673 & ~x697 & ~x700 & ~x701 & ~x724 & ~x725 & ~x731 & ~x759 & ~x780;
assign c8275 =  x362 &  x391;
assign c8277 =  x425 & ~x4 & ~x32 & ~x88 & ~x307 & ~x390 & ~x400 & ~x418 & ~x447 & ~x448 & ~x474 & ~x478 & ~x503 & ~x504 & ~x533 & ~x560 & ~x562 & ~x590 & ~x618 & ~x645 & ~x646 & ~x698 & ~x728 & ~x782;
assign c8279 =  x391;
assign c8281 =  x200;
assign c8283 =  x367 &  x395 & ~x598;
assign c8285 = ~x21 & ~x23 & ~x48 & ~x85 & ~x186 & ~x187 & ~x331 & ~x503 & ~x504 & ~x537 & ~x546 & ~x565 & ~x603 & ~x617 & ~x621 & ~x663 & ~x670 & ~x672 & ~x701;
assign c8287 =  x573 &  x656 & ~x330 & ~x479;
assign c8289 =  x387 &  x446 & ~x293;
assign c8291 = ~x9 & ~x11 & ~x65 & ~x133 & ~x192 & ~x219 & ~x223 & ~x468 & ~x493 & ~x541 & ~x567 & ~x620 & ~x622 & ~x625 & ~x669;
assign c8293 =  x500 &  x501 &  x529;
assign c8295 =  x171;
assign c8297 =  x487 &  x597 & ~x373;
assign c8299 = ~x59 & ~x60 & ~x140 & ~x164 & ~x166 & ~x192 & ~x195 & ~x249 & ~x308 & ~x320 & ~x321 & ~x350 & ~x367 & ~x446 & ~x449 & ~x450 & ~x451 & ~x476 & ~x505 & ~x529 & ~x530 & ~x532 & ~x588 & ~x591 & ~x616 & ~x641 & ~x643 & ~x647 & ~x670 & ~x672 & ~x674 & ~x698 & ~x699 & ~x701 & ~x726 & ~x780 & ~x781;
assign c8301 =  x363;
assign c8303 =  x372 &  x628 & ~x131 & ~x161;
assign c8305 =  x396 &  x611 & ~x482;
assign c8307 = ~x57 & ~x197 & ~x219 & ~x246 & ~x275 & ~x298 & ~x324 & ~x325 & ~x327 & ~x351 & ~x364 & ~x524 & ~x643 & ~x674 & ~x704 & ~x706 & ~x707 & ~x729 & ~x734 & ~x735;
assign c8309 = ~x112 & ~x195 & ~x224 & ~x347 & ~x348 & ~x349 & ~x421 & ~x423 & ~x451 & ~x452 & ~x531 & ~x586 & ~x615 & ~x671 & ~x701 & ~x708 & ~x736;
assign c8311 = ~x1 & ~x9 & ~x14 & ~x22 & ~x26 & ~x32 & ~x44 & ~x52 & ~x55 & ~x57 & ~x61 & ~x73 & ~x77 & ~x104 & ~x112 & ~x113 & ~x114 & ~x115 & ~x135 & ~x136 & ~x139 & ~x146 & ~x147 & ~x160 & ~x161 & ~x162 & ~x163 & ~x169 & ~x170 & ~x188 & ~x195 & ~x219 & ~x220 & ~x221 & ~x222 & ~x252 & ~x276 & ~x279 & ~x280 & ~x306 & ~x307 & ~x335 & ~x363 & ~x392 & ~x531 & ~x532 & ~x559 & ~x586 & ~x587 & ~x588 & ~x617 & ~x619 & ~x647 & ~x670 & ~x671 & ~x673 & ~x698 & ~x702 & ~x703 & ~x724 & ~x727 & ~x730 & ~x752 & ~x755 & ~x777;
assign c8313 =  x260 & ~x81 & ~x85 & ~x281 & ~x345 & ~x400 & ~x448 & ~x477 & ~x506 & ~x645 & ~x726;
assign c8315 =  x97 &  x99 & ~x403;
assign c8317 =  x118 & ~x70 & ~x592;
assign c8319 =  x79 & ~x274;
assign c8321 = ~x4 & ~x15 & ~x23 & ~x83 & ~x135 & ~x163 & ~x167 & ~x196 & ~x222 & ~x304 & ~x333 & ~x367 & ~x381 & ~x419 & ~x435 & ~x448 & ~x506 & ~x563 & ~x583 & ~x620 & ~x647 & ~x668 & ~x672 & ~x702 & ~x728 & ~x729 & ~x752;
assign c8323 =  x629 &  x658 & ~x534 & ~x606;
assign c8325 =  x76 & ~x344;
assign c8327 =  x183 &  x186 & ~x24 & ~x58 & ~x298 & ~x560 & ~x783;
assign c8329 = ~x22 & ~x23 & ~x52 & ~x55 & ~x60 & ~x111 & ~x112 & ~x166 & ~x198 & ~x304 & ~x333 & ~x361 & ~x449 & ~x503 & ~x504 & ~x505 & ~x533 & ~x559 & ~x561 & ~x586 & ~x589 & ~x605 & ~x616 & ~x644 & ~x688 & ~x689 & ~x700 & ~x716 & ~x724 & ~x726 & ~x728 & ~x744 & ~x745 & ~x746 & ~x748 & ~x749 & ~x753 & ~x755 & ~x763 & ~x781;
assign c8331 = ~x27 & ~x32 & ~x56 & ~x352 & ~x479 & ~x505 & ~x508 & ~x562 & ~x563 & ~x587 & ~x618 & ~x626 & ~x653 & ~x679 & ~x707;
assign c8333 =  x365 &  x366;
assign c8335 =  x203 & ~x28 & ~x55 & ~x223 & ~x316 & ~x336 & ~x344 & ~x345 & ~x390 & ~x446 & ~x473 & ~x615 & ~x700 & ~x774 & ~x783;
assign c8337 =  x177 &  x179 &  x180 & ~x590 & ~x704 & ~x756;
assign c8339 = ~x1 & ~x55 & ~x56 & ~x79 & ~x110 & ~x135 & ~x251 & ~x374 & ~x375 & ~x377 & ~x388 & ~x392 & ~x421 & ~x445 & ~x454 & ~x503 & ~x504 & ~x505 & ~x645;
assign c8341 =  x207 & ~x80 & ~x193 & ~x216 & ~x361 & ~x431 & ~x449 & ~x457 & ~x481 & ~x533 & ~x535;
assign c8343 = ~x51 & ~x54 & ~x108 & ~x165 & ~x172 & ~x198 & ~x254 & ~x278 & ~x279 & ~x337 & ~x346 & ~x361 & ~x363 & ~x391 & ~x392 & ~x420 & ~x450 & ~x477 & ~x490 & ~x505 & ~x555 & ~x556 & ~x557 & ~x562 & ~x588 & ~x589 & ~x590 & ~x614 & ~x616 & ~x617 & ~x631 & ~x640 & ~x645 & ~x646 & ~x673 & ~x674 & ~x700 & ~x701 & ~x726 & ~x727 & ~x728 & ~x729 & ~x753 & ~x754 & ~x764 & ~x766 & ~x781;
assign c8345 = ~x4 & ~x50 & ~x54 & ~x85 & ~x116 & ~x143 & ~x171 & ~x192 & ~x221 & ~x244 & ~x330 & ~x335 & ~x364 & ~x365 & ~x366 & ~x368 & ~x394 & ~x416 & ~x451 & ~x452 & ~x499 & ~x506 & ~x532 & ~x533 & ~x536 & ~x547 & ~x556 & ~x589 & ~x593 & ~x616 & ~x618 & ~x619 & ~x631 & ~x640 & ~x644 & ~x645 & ~x646 & ~x665 & ~x668 & ~x694 & ~x704 & ~x735 & ~x779;
assign c8347 = ~x3 & ~x4 & ~x24 & ~x28 & ~x29 & ~x31 & ~x55 & ~x58 & ~x111 & ~x112 & ~x168 & ~x307 & ~x334 & ~x336 & ~x363 & ~x391 & ~x392 & ~x393 & ~x419 & ~x424 & ~x446 & ~x447 & ~x448 & ~x452 & ~x476 & ~x477 & ~x480 & ~x503 & ~x504 & ~x559 & ~x599 & ~x616 & ~x627 & ~x644 & ~x653 & ~x654 & ~x680 & ~x681 & ~x707 & ~x708 & ~x727 & ~x762 & ~x778 & ~x780 & ~x782 & ~x783;
assign c8349 =  x606 & ~x225 & ~x347 & ~x509 & ~x728 & ~x778;
assign c8351 = ~x169 & ~x171 & ~x191 & ~x195 & ~x276 & ~x416 & ~x450 & ~x477 & ~x479 & ~x508 & ~x570 & ~x618 & ~x625 & ~x671 & ~x681 & ~x707 & ~x728;
assign c8353 = ~x359;
assign c8355 = ~x3 & ~x28 & ~x29 & ~x48 & ~x79 & ~x269 & ~x275 & ~x365 & ~x423 & ~x470 & ~x498 & ~x504 & ~x506 & ~x507 & ~x509 & ~x528 & ~x529 & ~x534 & ~x555 & ~x589 & ~x592 & ~x593 & ~x602 & ~x619 & ~x649 & ~x674 & ~x675 & ~x676 & ~x699 & ~x703 & ~x727 & ~x734 & ~x759 & ~x778 & ~x780;
assign c8357 =  x237 &  x686 & ~x680 & ~x708;
assign c8359 =  x118 & ~x533 & ~x641 & ~x749;
assign c8361 =  x230 & ~x344 & ~x399 & ~x418 & ~x561 & ~x645;
assign c8363 =  x301 & ~x107 & ~x411 & ~x413;
assign c8365 =  x651 & ~x152 & ~x262 & ~x317 & ~x344 & ~x345 & ~x455 & ~x587;
assign c8367 =  x303 &  x419;
assign c8369 =  x632 & ~x117 & ~x566 & ~x596 & ~x758;
assign c8371 =  x87;
assign c8373 =  x344 & ~x57 & ~x104 & ~x338 & ~x364 & ~x368 & ~x476 & ~x624 & ~x651 & ~x671 & ~x679 & ~x733 & ~x734 & ~x735 & ~x736;
assign c8375 =  x212 & ~x0 & ~x3 & ~x30 & ~x31 & ~x61 & ~x84 & ~x86 & ~x111 & ~x137 & ~x142 & ~x166 & ~x197 & ~x226 & ~x250 & ~x254 & ~x277 & ~x280 & ~x282 & ~x310 & ~x317 & ~x334 & ~x335 & ~x394 & ~x400 & ~x436 & ~x447 & ~x474 & ~x476 & ~x502 & ~x503 & ~x505 & ~x531 & ~x586 & ~x699 & ~x758 & ~x781;
assign c8377 =  x300 & ~x18 & ~x439 & ~x505 & ~x619;
assign c8379 =  x96 &  x408 & ~x721;
assign c8381 =  x184 &  x573;
assign c8383 = ~x32 & ~x144 & ~x227 & ~x229 & ~x275 & ~x338 & ~x418 & ~x430 & ~x431 & ~x432 & ~x485 & ~x507 & ~x561 & ~x646 & ~x667;
assign c8385 = ~x6 & ~x55 & ~x112 & ~x159 & ~x376 & ~x418 & ~x449 & ~x547 & ~x561 & ~x589 & ~x592 & ~x700 & ~x734;
assign c8387 =  x711 & ~x1 & ~x130 & ~x170 & ~x362 & ~x365 & ~x460 & ~x475 & ~x476 & ~x488 & ~x558 & ~x585 & ~x591 & ~x648 & ~x675 & ~x702;
assign c8389 =  x547 &  x603 & ~x60 & ~x450 & ~x673 & ~x747;
assign c8391 =  x89 &  x119;
assign c8393 =  x759;
assign c8395 =  x205 & ~x344 & ~x602 & ~x719;
assign c8397 =  x240 &  x327 & ~x344 & ~x345;
assign c8399 =  x267 & ~x403 & ~x404 & ~x536 & ~x538 & ~x562 & ~x722 & ~x726 & ~x735;
assign c8401 = ~x32 & ~x81 & ~x83 & ~x196 & ~x226 & ~x241 & ~x250 & ~x281 & ~x330 & ~x363 & ~x388 & ~x419 & ~x476 & ~x503 & ~x532 & ~x561 & ~x589 & ~x623 & ~x624 & ~x625 & ~x644 & ~x652 & ~x678 & ~x679 & ~x681 & ~x707 & ~x734 & ~x760 & ~x761 & ~x763 & ~x779;
assign c8403 = ~x20 & ~x28 & ~x77 & ~x84 & ~x163 & ~x169 & ~x192 & ~x212 & ~x218 & ~x476 & ~x497 & ~x554 & ~x575 & ~x606 & ~x609 & ~x633 & ~x660 & ~x700 & ~x727 & ~x732 & ~x735 & ~x755;
assign c8405 = ~x0 & ~x16 & ~x17 & ~x22 & ~x23 & ~x24 & ~x45 & ~x62 & ~x73 & ~x103 & ~x106 & ~x113 & ~x137 & ~x143 & ~x145 & ~x174 & ~x196 & ~x198 & ~x216 & ~x225 & ~x282 & ~x310 & ~x336 & ~x391 & ~x393 & ~x415 & ~x417 & ~x422 & ~x446 & ~x449 & ~x478 & ~x502 & ~x503 & ~x531 & ~x560 & ~x601 & ~x619 & ~x637 & ~x649 & ~x663 & ~x724 & ~x729 & ~x750;
assign c8407 =  x386 & ~x132 & ~x246;
assign c8409 =  x549 & ~x17 & ~x71 & ~x141 & ~x533 & ~x561 & ~x590 & ~x719;
assign c8411 =  x296 &  x610 & ~x656;
assign c8413 = ~x34 & ~x49 & ~x143 & ~x320 & ~x321 & ~x394 & ~x449 & ~x451 & ~x506 & ~x568 & ~x641 & ~x645 & ~x668 & ~x768;
assign c8415 =  x273 &  x274 & ~x95 & ~x105;
assign c8417 = ~x284 & ~x360 & ~x406 & ~x416 & ~x427 & ~x450 & ~x478 & ~x500 & ~x529 & ~x575 & ~x661 & ~x668 & ~x766;
assign c8419 =  x361 & ~x650;
assign c8421 = ~x5 & ~x6 & ~x27 & ~x31 & ~x83 & ~x86 & ~x167 & ~x170 & ~x224 & ~x254 & ~x282 & ~x333 & ~x370 & ~x394 & ~x419 & ~x420 & ~x450 & ~x529 & ~x561 & ~x586 & ~x612 & ~x614 & ~x615 & ~x644 & ~x672 & ~x681 & ~x697 & ~x707 & ~x764 & ~x782;
assign c8423 = ~x58 & ~x158 & ~x267 & ~x273 & ~x419 & ~x600 & ~x673 & ~x674 & ~x681 & ~x729 & ~x737 & ~x753;
assign c8425 =  x520 &  x581;
assign c8427 = ~x108 & ~x109 & ~x141 & ~x200 & ~x201 & ~x276 & ~x373 & ~x377 & ~x387 & ~x421 & ~x432 & ~x505 & ~x508 & ~x555 & ~x699;
assign c8429 =  x89 & ~x561;
assign c8431 =  x603 &  x633;
assign c8433 = ~x3 & ~x59 & ~x111 & ~x138 & ~x144 & ~x165 & ~x168 & ~x225 & ~x310 & ~x336 & ~x360 & ~x361 & ~x365 & ~x422 & ~x451 & ~x477 & ~x478 & ~x479 & ~x535 & ~x557 & ~x562 & ~x563 & ~x613 & ~x616 & ~x619 & ~x626 & ~x627 & ~x641 & ~x655 & ~x668 & ~x670 & ~x681 & ~x737 & ~x757 & ~x763 & ~x764 & ~x780 & ~x783;
assign c8435 =  x285 & ~x453 & ~x481 & ~x764;
assign c8437 = ~x2 & ~x24 & ~x28 & ~x31 & ~x58 & ~x82 & ~x86 & ~x89 & ~x112 & ~x113 & ~x118 & ~x135 & ~x140 & ~x169 & ~x248 & ~x277 & ~x280 & ~x281 & ~x312 & ~x341 & ~x359 & ~x365 & ~x390 & ~x395 & ~x396 & ~x415 & ~x445 & ~x446 & ~x475 & ~x478 & ~x502 & ~x507 & ~x508 & ~x512 & ~x527 & ~x535 & ~x536 & ~x554 & ~x563 & ~x582 & ~x585 & ~x588 & ~x590 & ~x612 & ~x639 & ~x641 & ~x649 & ~x666 & ~x670 & ~x677 & ~x751 & ~x752 & ~x772;
assign c8439 =  x317 &  x573 & ~x702;
assign c8441 =  x175 & ~x504 & ~x507 & ~x535 & ~x591 & ~x617 & ~x735;
assign c8443 = ~x29 & ~x32 & ~x55 & ~x113 & ~x151 & ~x197 & ~x206 & ~x207 & ~x262 & ~x289 & ~x344 & ~x372 & ~x417 & ~x447 & ~x488 & ~x503 & ~x572 & ~x602 & ~x630 & ~x655 & ~x672 & ~x711 & ~x782 & ~x783;
assign c8445 =  x501 & ~x623 & ~x624;
assign c8447 =  x685 &  x714 & ~x652 & ~x705;
assign c8449 =  x258 & ~x289 & ~x316 & ~x399 & ~x427;
assign c8451 = ~x20 & ~x31 & ~x81 & ~x111 & ~x173 & ~x189 & ~x195 & ~x198 & ~x221 & ~x255 & ~x256 & ~x362 & ~x378 & ~x379 & ~x389 & ~x406 & ~x418 & ~x450 & ~x500 & ~x507 & ~x534 & ~x585 & ~x589 & ~x619 & ~x643 & ~x672 & ~x676 & ~x731 & ~x732;
assign c8453 =  x519 &  x579 & ~x1 & ~x3 & ~x4 & ~x18 & ~x20 & ~x26 & ~x32 & ~x54 & ~x55 & ~x58 & ~x59 & ~x85 & ~x87 & ~x111 & ~x112 & ~x115 & ~x116 & ~x141 & ~x142 & ~x198 & ~x224 & ~x253 & ~x281 & ~x282 & ~x283 & ~x305 & ~x309 & ~x333 & ~x336 & ~x337 & ~x338 & ~x362 & ~x363 & ~x365 & ~x366 & ~x389 & ~x421 & ~x422 & ~x448 & ~x449 & ~x450 & ~x473 & ~x476 & ~x477 & ~x478 & ~x503 & ~x504 & ~x505 & ~x531 & ~x533 & ~x560 & ~x561 & ~x588 & ~x617 & ~x698 & ~x699 & ~x707 & ~x727 & ~x734 & ~x736 & ~x738 & ~x755 & ~x756 & ~x757 & ~x781 & ~x783;
assign c8455 =  x357 & ~x161 & ~x188 & ~x216 & ~x217 & ~x218 & ~x246 & ~x752;
assign c8457 = ~x18 & ~x528 & ~x597 & ~x651 & ~x653 & ~x703 & ~x706 & ~x749 & ~x750;
assign c8459 =  x411 & ~x15 & ~x196 & ~x215 & ~x216 & ~x665;
assign c8461 = ~x10 & ~x53 & ~x109 & ~x166 & ~x310 & ~x395 & ~x422 & ~x424 & ~x459 & ~x512 & ~x639 & ~x717 & ~x726 & ~x745;
assign c8463 =  x396 & ~x6 & ~x25 & ~x29 & ~x32 & ~x55 & ~x84 & ~x85 & ~x111 & ~x114 & ~x169 & ~x227 & ~x280 & ~x306 & ~x308 & ~x363 & ~x418 & ~x447 & ~x449 & ~x476 & ~x502 & ~x505 & ~x531 & ~x532 & ~x533 & ~x560 & ~x561 & ~x586 & ~x587 & ~x588 & ~x589 & ~x615 & ~x616 & ~x671 & ~x673 & ~x726;
assign c8465 =  x713 & ~x23 & ~x46 & ~x51 & ~x72 & ~x78 & ~x79 & ~x82 & ~x83 & ~x84 & ~x110 & ~x166 & ~x171 & ~x187 & ~x362 & ~x364 & ~x420 & ~x422 & ~x446 & ~x503 & ~x505 & ~x528 & ~x530 & ~x533 & ~x562 & ~x588 & ~x614 & ~x616 & ~x635 & ~x641 & ~x663 & ~x664 & ~x666 & ~x700 & ~x702 & ~x730 & ~x732 & ~x733 & ~x762 & ~x763 & ~x781;
assign c8467 = ~x9 & ~x55 & ~x197 & ~x241 & ~x267 & ~x532 & ~x555 & ~x586 & ~x621;
assign c8469 = ~x2 & ~x5 & ~x16 & ~x17 & ~x18 & ~x77 & ~x134 & ~x135 & ~x170 & ~x225 & ~x226 & ~x282 & ~x308 & ~x360 & ~x361 & ~x368 & ~x418 & ~x424 & ~x425 & ~x461 & ~x462 & ~x474 & ~x476 & ~x508 & ~x531 & ~x532 & ~x559 & ~x590 & ~x669 & ~x674 & ~x698 & ~x700 & ~x726 & ~x727 & ~x781;
assign c8471 =  x279;
assign c8473 = ~x121 & ~x159 & ~x187 & ~x476 & ~x512 & ~x540 & ~x562 & ~x567 & ~x591 & ~x594 & ~x614 & ~x673 & ~x674 & ~x697 & ~x744;
assign c8475 =  x204 & ~x372 & ~x427 & ~x504 & ~x549;
assign c8477 =  x118 &  x145 &  x161;
assign c8479 =  x606 & ~x446 & ~x485 & ~x505 & ~x590 & ~x645;
assign c8481 =  x466 & ~x280 & ~x444 & ~x536 & ~x574 & ~x665 & ~x692 & ~x722;
assign c8483 = ~x12 & ~x21 & ~x35 & ~x269 & ~x270 & ~x368 & ~x383 & ~x420 & ~x582 & ~x583 & ~x585 & ~x603 & ~x640 & ~x722;
assign c8485 =  x203 & ~x42 & ~x123 & ~x344 & ~x399 & ~x530 & ~x561 & ~x576 & ~x617 & ~x630 & ~x657 & ~x672 & ~x753;
assign c8487 = ~x17 & ~x19 & ~x104 & ~x375 & ~x735;
assign c8489 = ~x104 & ~x407 & ~x431 & ~x432 & ~x477 & ~x481 & ~x482 & ~x504 & ~x673;
assign c8491 =  x198;
assign c8493 =  x573 &  x600 & ~x132 & ~x476 & ~x767;
assign c8495 =  x97 &  x126 &  x711 &  x740 & ~x46 & ~x533;
assign c8497 =  x119 & ~x9 & ~x182 & ~x704;
assign c8499 = ~x536 & ~x565 & ~x570 & ~x596 & ~x620 & ~x626 & ~x653 & ~x706 & ~x722 & ~x751 & ~x779;
assign c90 =  x273 & ~x46 & ~x104 & ~x105 & ~x130 & ~x153 & ~x363 & ~x385 & ~x390 & ~x420 & ~x422 & ~x440 & ~x450 & ~x470 & ~x477 & ~x526 & ~x560 & ~x701 & ~x702;
assign c92 = ~x10 & ~x21 & ~x26 & ~x51 & ~x54 & ~x55 & ~x72 & ~x76 & ~x101 & ~x109 & ~x137 & ~x140 & ~x165 & ~x186 & ~x190 & ~x192 & ~x212 & ~x218 & ~x242 & ~x245 & ~x246 & ~x269 & ~x281 & ~x295 & ~x334 & ~x362 & ~x380 & ~x503 & ~x557 & ~x610 & ~x611 & ~x636 & ~x639 & ~x640 & ~x641 & ~x642 & ~x673 & ~x675 & ~x726 & ~x751 & ~x760;
assign c94 = ~x43 & ~x46 & ~x50 & ~x56 & ~x105 & ~x130 & ~x183 & ~x185 & ~x211 & ~x344 & ~x364 & ~x367 & ~x397 & ~x398 & ~x415 & ~x421 & ~x441 & ~x446 & ~x468 & ~x499 & ~x505 & ~x528 & ~x533 & ~x618 & ~x696 & ~x763;
assign c96 =  x266 &  x295 &  x352 & ~x359 & ~x444 & ~x500 & ~x708 & ~x756 & ~x770;
assign c98 = ~x0 & ~x18 & ~x76 & ~x79 & ~x111 & ~x185 & ~x290 & ~x317 & ~x344 & ~x345 & ~x392 & ~x421 & ~x440 & ~x447 & ~x451 & ~x452 & ~x476 & ~x506 & ~x701 & ~x702;
assign c910 =  x207 &  x713 &  x717 & ~x55 & ~x139 & ~x279 & ~x281 & ~x285 & ~x311 & ~x314 & ~x337 & ~x342 & ~x447 & ~x449 & ~x502 & ~x530 & ~x531 & ~x579 & ~x580 & ~x581 & ~x583 & ~x586 & ~x593 & ~x607 & ~x614 & ~x618 & ~x620 & ~x621 & ~x644 & ~x645 & ~x646 & ~x647 & ~x648 & ~x675 & ~x676 & ~x701 & ~x729;
assign c912 =  x293 &  x294 &  x322 &  x323 &  x350 &  x351 & ~x21 & ~x26 & ~x27 & ~x280 & ~x336 & ~x360 & ~x361 & ~x364 & ~x390 & ~x391 & ~x392 & ~x416 & ~x417 & ~x419 & ~x420 & ~x444 & ~x445 & ~x446 & ~x447 & ~x448 & ~x473 & ~x474 & ~x500 & ~x501 & ~x504 & ~x529 & ~x530 & ~x531 & ~x559 & ~x586 & ~x587 & ~x615 & ~x735 & ~x736 & ~x757 & ~x763;
assign c914 = ~x12 & ~x84 & ~x126 & ~x127 & ~x139 & ~x153 & ~x154 & ~x155 & ~x182 & ~x336 & ~x371 & ~x393 & ~x398 & ~x399 & ~x417 & ~x418 & ~x421 & ~x423 & ~x445 & ~x503 & ~x504 & ~x505 & ~x506 & ~x507 & ~x532 & ~x562 & ~x586 & ~x589 & ~x590 & ~x673 & ~x730 & ~x756 & ~x763 & ~x782;
assign c916 = ~x2 & ~x10 & ~x11 & ~x13 & ~x14 & ~x21 & ~x22 & ~x26 & ~x39 & ~x40 & ~x76 & ~x101 & ~x122 & ~x336 & ~x369 & ~x475 & ~x497 & ~x500 & ~x503 & ~x524 & ~x526 & ~x556 & ~x557 & ~x612 & ~x613 & ~x614 & ~x642 & ~x696 & ~x723 & ~x728 & ~x730 & ~x731 & ~x756 & ~x759 & ~x779 & ~x782;
assign c918 =  x741 &  x742 & ~x98 & ~x493 & ~x524 & ~x525 & ~x530 & ~x553 & ~x554 & ~x604 & ~x637 & ~x639 & ~x761 & ~x779 & ~x780;
assign c920 =  x496 & ~x273 & ~x280 & ~x301 & ~x318 & ~x362 & ~x388 & ~x391 & ~x419 & ~x448 & ~x529 & ~x530 & ~x534 & ~x561 & ~x635 & ~x663 & ~x692;
assign c922 =  x466 &  x637 & ~x470 & ~x526 & ~x527 & ~x555 & ~x583 & ~x698 & ~x774 & ~x775;
assign c924 =  x302 & ~x74 & ~x99 & ~x107 & ~x128 & ~x131 & ~x132 & ~x133 & ~x156 & ~x157 & ~x159 & ~x160 & ~x162 & ~x163 & ~x184 & ~x185 & ~x417 & ~x418 & ~x423 & ~x443 & ~x446 & ~x469 & ~x470 & ~x471 & ~x472 & ~x473 & ~x475 & ~x502 & ~x528 & ~x558 & ~x614 & ~x616 & ~x642 & ~x672 & ~x673 & ~x698 & ~x725;
assign c926 =  x744 & ~x525 & ~x540 & ~x568 & ~x580 & ~x610 & ~x633 & ~x658 & ~x661;
assign c928 =  x461 & ~x42 & ~x44 & ~x158 & ~x338 & ~x339 & ~x415 & ~x417 & ~x439 & ~x440 & ~x444 & ~x466 & ~x469 & ~x474 & ~x497 & ~x645 & ~x674 & ~x703;
assign c930 =  x497 &  x583 &  x640 &  x697 & ~x637 & ~x665;
assign c932 =  x110 & ~x277;
assign c934 = ~x70 & ~x204 & ~x245 & ~x396 & ~x447 & ~x576 & ~x579 & ~x639;
assign c936 = ~x5 & ~x7 & ~x19 & ~x22 & ~x24 & ~x27 & ~x28 & ~x47 & ~x48 & ~x50 & ~x52 & ~x56 & ~x77 & ~x78 & ~x80 & ~x81 & ~x83 & ~x84 & ~x104 & ~x106 & ~x111 & ~x112 & ~x131 & ~x133 & ~x134 & ~x136 & ~x156 & ~x159 & ~x162 & ~x163 & ~x184 & ~x185 & ~x186 & ~x187 & ~x189 & ~x208 & ~x209 & ~x223 & ~x236 & ~x237 & ~x265 & ~x266 & ~x307 & ~x420 & ~x476 & ~x477 & ~x498 & ~x500 & ~x501 & ~x504 & ~x505 & ~x526 & ~x527 & ~x528 & ~x533 & ~x555 & ~x581 & ~x583 & ~x587 & ~x588 & ~x589 & ~x617 & ~x644 & ~x673 & ~x700 & ~x702 & ~x725 & ~x726 & ~x727 & ~x729 & ~x757 & ~x758 & ~x759 & ~x781;
assign c938 =  x205 &  x386 &  x741 &  x743 & ~x106 & ~x140 & ~x213 & ~x503 & ~x554;
assign c940 = ~x2 & ~x126 & ~x133 & ~x155 & ~x167 & ~x184 & ~x308 & ~x343 & ~x367 & ~x394 & ~x419 & ~x440 & ~x441 & ~x444 & ~x468 & ~x470 & ~x471 & ~x473 & ~x498 & ~x499 & ~x550 & ~x563 & ~x588 & ~x589 & ~x670 & ~x699 & ~x729 & ~x754 & ~x765;
assign c942 = ~x21 & ~x23 & ~x48 & ~x132 & ~x135 & ~x161 & ~x162 & ~x186 & ~x237 & ~x266 & ~x283 & ~x294 & ~x296 & ~x475 & ~x551 & ~x554 & ~x578 & ~x579 & ~x580 & ~x581 & ~x593 & ~x607 & ~x611 & ~x612 & ~x620 & ~x643 & ~x648 & ~x669 & ~x674 & ~x675 & ~x704 & ~x760;
assign c944 =  x621 & ~x35 & ~x36 & ~x234 & ~x262 & ~x263 & ~x330 & ~x335 & ~x391 & ~x393 & ~x420 & ~x531 & ~x534 & ~x717 & ~x756 & ~x763;
assign c946 =  x519 &  x744 & ~x28 & ~x189 & ~x250 & ~x514 & ~x542 & ~x596 & ~x666 & ~x725 & ~x758;
assign c948 =  x464 & ~x0 & ~x167 & ~x280 & ~x308 & ~x388 & ~x391 & ~x446 & ~x448 & ~x502 & ~x503 & ~x504 & ~x530 & ~x532 & ~x558 & ~x559 & ~x597 & ~x605 & ~x615 & ~x625 & ~x652 & ~x659 & ~x662 & ~x707 & ~x733 & ~x734 & ~x756;
assign c950 =  x78 & ~x25 & ~x151 & ~x219 & ~x246 & ~x249 & ~x276 & ~x277 & ~x303 & ~x305 & ~x476;
assign c952 = ~x26 & ~x67 & ~x81 & ~x94 & ~x134 & ~x151 & ~x213 & ~x237 & ~x391 & ~x393 & ~x563 & ~x589 & ~x619 & ~x646 & ~x669 & ~x672 & ~x730;
assign c954 =  x467 &  x524 & ~x300 & ~x307 & ~x330 & ~x358 & ~x448 & ~x499 & ~x532 & ~x556 & ~x586 & ~x635 & ~x661 & ~x691 & ~x718;
assign c956 =  x442 & ~x2 & ~x161 & ~x218 & ~x246 & ~x247 & ~x252 & ~x275 & ~x276 & ~x277 & ~x304 & ~x305 & ~x307 & ~x334 & ~x504 & ~x552 & ~x553 & ~x578 & ~x580 & ~x581 & ~x603 & ~x609 & ~x615 & ~x635 & ~x638;
assign c958 =  x378 &  x406 & ~x2 & ~x15 & ~x16 & ~x17 & ~x22 & ~x23 & ~x29 & ~x30 & ~x41 & ~x42 & ~x43 & ~x53 & ~x54 & ~x56 & ~x69 & ~x82 & ~x111 & ~x306 & ~x332 & ~x333 & ~x334 & ~x335 & ~x360 & ~x361 & ~x362 & ~x388 & ~x391 & ~x392 & ~x416 & ~x417 & ~x418 & ~x420 & ~x445 & ~x446 & ~x447 & ~x448 & ~x473 & ~x475 & ~x502 & ~x503 & ~x504 & ~x505 & ~x531 & ~x558 & ~x588 & ~x615 & ~x681 & ~x756;
assign c960 =  x234 &  x289 & ~x132 & ~x190 & ~x242 & ~x246 & ~x312 & ~x484 & ~x559 & ~x610 & ~x619 & ~x644;
assign c962 = ~x165 & ~x167 & ~x189 & ~x226 & ~x243 & ~x375 & ~x429 & ~x458 & ~x502 & ~x566 & ~x586 & ~x649 & ~x669;
assign c964 =  x238 &  x295 & ~x25 & ~x28 & ~x359 & ~x360 & ~x391 & ~x444 & ~x446 & ~x560 & ~x614 & ~x689 & ~x736 & ~x742 & ~x747;
assign c966 =  x273 & ~x359 & ~x363 & ~x384 & ~x414 & ~x415 & ~x451 & ~x670 & ~x674 & ~x761;
assign c968 = ~x26 & ~x69 & ~x152 & ~x279 & ~x390 & ~x415 & ~x445 & ~x529 & ~x530 & ~x551 & ~x558 & ~x573 & ~x577 & ~x578 & ~x600 & ~x604 & ~x608 & ~x635 & ~x637 & ~x665;
assign c970 =  x293 & ~x2 & ~x26 & ~x53 & ~x223 & ~x252 & ~x319 & ~x401 & ~x445 & ~x446 & ~x447 & ~x529 & ~x615 & ~x680 & ~x707 & ~x709;
assign c972 =  x268 &  x382 &  x439 &  x524 &  x581 & ~x358 & ~x635 & ~x691;
assign c974 = ~x132 & ~x159 & ~x165 & ~x184 & ~x191 & ~x223 & ~x266 & ~x280 & ~x293 & ~x294 & ~x295 & ~x308 & ~x352 & ~x508 & ~x581 & ~x585 & ~x613 & ~x616 & ~x642 & ~x647 & ~x674 & ~x730;
assign c976 =  x508 & ~x390 & ~x446 & ~x602 & ~x633 & ~x663 & ~x679 & ~x705 & ~x719;
assign c978 =  x137 &  x295 & ~x304;
assign c980 =  x322 &  x350 &  x378 &  x715 & ~x0 & ~x28 & ~x155 & ~x280 & ~x364 & ~x391 & ~x473 & ~x495 & ~x496 & ~x500 & ~x522 & ~x523 & ~x524 & ~x525 & ~x550 & ~x552 & ~x559 & ~x560 & ~x562 & ~x613 & ~x615 & ~x618 & ~x647 & ~x674;
assign c982 =  x238 & ~x0 & ~x55 & ~x84 & ~x85 & ~x280 & ~x304 & ~x317 & ~x336 & ~x344 & ~x445 & ~x473 & ~x474 & ~x502 & ~x531 & ~x596 & ~x603 & ~x624 & ~x651 & ~x653 & ~x681 & ~x707 & ~x734 & ~x735 & ~x762;
assign c984 =  x413 &  x739 &  x741 &  x743 & ~x191 & ~x193 & ~x221 & ~x566 & ~x581 & ~x582 & ~x605;
assign c986 = ~x2 & ~x7 & ~x27 & ~x54 & ~x55 & ~x59 & ~x60 & ~x80 & ~x130 & ~x336 & ~x365 & ~x441 & ~x443 & ~x477 & ~x500 & ~x502 & ~x506 & ~x507 & ~x558 & ~x561 & ~x562 & ~x564 & ~x587 & ~x645 & ~x717 & ~x718 & ~x740 & ~x741 & ~x743 & ~x745 & ~x766 & ~x773 & ~x774;
assign c988 = ~x30 & ~x49 & ~x80 & ~x81 & ~x137 & ~x163 & ~x167 & ~x186 & ~x190 & ~x191 & ~x238 & ~x245 & ~x251 & ~x278 & ~x297 & ~x428 & ~x454 & ~x475 & ~x500 & ~x537 & ~x551 & ~x560 & ~x563 & ~x580 & ~x581 & ~x582 & ~x584 & ~x585 & ~x590 & ~x591 & ~x592 & ~x617 & ~x643 & ~x703 & ~x761;
assign c990 = ~x27 & ~x28 & ~x65 & ~x93 & ~x151 & ~x152 & ~x179 & ~x208 & ~x237 & ~x393 & ~x420 & ~x452 & ~x473 & ~x507 & ~x532 & ~x533 & ~x535 & ~x561 & ~x674 & ~x729 & ~x737 & ~x756 & ~x757 & ~x764 & ~x770 & ~x774 & ~x778;
assign c992 =  x435 &  x744 & ~x17 & ~x28 & ~x77 & ~x139 & ~x165 & ~x187 & ~x402 & ~x420 & ~x456 & ~x476 & ~x482 & ~x510 & ~x529 & ~x538 & ~x551 & ~x554 & ~x556 & ~x590 & ~x607 & ~x614 & ~x616 & ~x635 & ~x639 & ~x645 & ~x703 & ~x734;
assign c994 = ~x76 & ~x156 & ~x183 & ~x223 & ~x311 & ~x428 & ~x469 & ~x473 & ~x498 & ~x508 & ~x509 & ~x522 & ~x524 & ~x550 & ~x731 & ~x759 & ~x774;
assign c996 = ~x18 & ~x71 & ~x72 & ~x124 & ~x153 & ~x262 & ~x320 & ~x365 & ~x398 & ~x415 & ~x445 & ~x473 & ~x478 & ~x500 & ~x561;
assign c998 =  x357 & ~x187 & ~x190 & ~x192 & ~x215 & ~x240 & ~x244 & ~x426 & ~x445 & ~x473 & ~x475 & ~x496 & ~x498 & ~x503 & ~x525 & ~x526;
assign c9100 =  x59 & ~x9 & ~x528 & ~x557 & ~x585 & ~x607 & ~x635;
assign c9102 =  x145 &  x459 & ~x43 & ~x336 & ~x364 & ~x366 & ~x450 & ~x451 & ~x452 & ~x473 & ~x474 & ~x475 & ~x503 & ~x504 & ~x532 & ~x533 & ~x534 & ~x559 & ~x562 & ~x590 & ~x616 & ~x617 & ~x644 & ~x646 & ~x670 & ~x701 & ~x754 & ~x757;
assign c9104 =  x324 & ~x29 & ~x31 & ~x329 & ~x330 & ~x332 & ~x336 & ~x357 & ~x362 & ~x416 & ~x473 & ~x529 & ~x530 & ~x532 & ~x713 & ~x714 & ~x737 & ~x738 & ~x741 & ~x744 & ~x745 & ~x768 & ~x774;
assign c9106 =  x468 &  x469 &  x583 & ~x608 & ~x665 & ~x722;
assign c9108 =  x351 & ~x28 & ~x35 & ~x62 & ~x98 & ~x125 & ~x167 & ~x196 & ~x388 & ~x390 & ~x391 & ~x417 & ~x418 & ~x448 & ~x475 & ~x587 & ~x709 & ~x741 & ~x744 & ~x746 & ~x774;
assign c9110 = ~x79 & ~x99 & ~x110 & ~x127 & ~x444 & ~x452 & ~x454 & ~x499 & ~x522 & ~x555 & ~x616 & ~x732 & ~x754;
assign c9112 =  x632 & ~x9 & ~x14 & ~x22 & ~x156 & ~x157 & ~x481 & ~x563 & ~x742 & ~x772 & ~x775;
assign c9114 =  x481 & ~x304 & ~x391 & ~x475 & ~x552 & ~x560 & ~x603 & ~x609 & ~x627 & ~x665 & ~x695;
assign c9116 =  x207 & ~x26 & ~x30 & ~x47 & ~x74 & ~x160 & ~x162 & ~x195 & ~x222 & ~x310 & ~x431 & ~x446 & ~x449 & ~x511 & ~x512 & ~x552 & ~x558 & ~x580 & ~x582 & ~x621 & ~x675 & ~x704 & ~x757;
assign c9118 = ~x21 & ~x34 & ~x50 & ~x51 & ~x53 & ~x75 & ~x80 & ~x104 & ~x132 & ~x185 & ~x186 & ~x212 & ~x367 & ~x369 & ~x446 & ~x592 & ~x675 & ~x709 & ~x737 & ~x765 & ~x771 & ~x774 & ~x781;
assign c9120 = ~x155 & ~x156 & ~x388 & ~x426 & ~x452 & ~x473 & ~x492 & ~x494 & ~x505 & ~x520 & ~x533 & ~x550 & ~x648;
assign c9122 = ~x275 & ~x308 & ~x333 & ~x334 & ~x361 & ~x504 & ~x531 & ~x559 & ~x571 & ~x579 & ~x588 & ~x627 & ~x633 & ~x634 & ~x657 & ~x662 & ~x686 & ~x714 & ~x720 & ~x737 & ~x749 & ~x763 & ~x765;
assign c9124 = ~x12 & ~x21 & ~x22 & ~x47 & ~x49 & ~x68 & ~x71 & ~x78 & ~x139 & ~x157 & ~x360 & ~x385 & ~x415 & ~x416 & ~x445 & ~x447 & ~x476 & ~x500 & ~x502 & ~x530 & ~x585 & ~x588 & ~x680 & ~x706 & ~x707 & ~x733 & ~x737 & ~x738 & ~x766 & ~x783;
assign c9126 =  x107 &  x239 &  x267 & ~x276;
assign c9128 =  x332 & ~x17 & ~x134 & ~x136 & ~x138 & ~x218 & ~x243 & ~x442 & ~x470 & ~x473 & ~x532 & ~x558 & ~x559 & ~x646;
assign c9130 =  x211 &  x313 & ~x60 & ~x168 & ~x225 & ~x234 & ~x245 & ~x262 & ~x318 & ~x417 & ~x478 & ~x504 & ~x534 & ~x560 & ~x561 & ~x662;
assign c9132 =  x742 & ~x160 & ~x309 & ~x457 & ~x604 & ~x606 & ~x608 & ~x632;
assign c9134 =  x201 & ~x20 & ~x25 & ~x45 & ~x48 & ~x92 & ~x135 & ~x136 & ~x161 & ~x189 & ~x192 & ~x243 & ~x395 & ~x509 & ~x620 & ~x696 & ~x700 & ~x732;
assign c9136 =  x137 & ~x151 & ~x219 & ~x248 & ~x277 & ~x279 & ~x305 & ~x447 & ~x679;
assign c9138 =  x436 & ~x5 & ~x29 & ~x189 & ~x233 & ~x415 & ~x417 & ~x472 & ~x502 & ~x679 & ~x683;
assign c9140 =  x234 &  x489 & ~x194 & ~x471 & ~x503 & ~x610 & ~x729;
assign c9142 =  x206 &  x742 &  x743 & ~x53 & ~x84 & ~x132 & ~x135 & ~x139 & ~x157 & ~x186 & ~x196 & ~x238 & ~x239 & ~x257 & ~x284 & ~x501 & ~x502 & ~x528 & ~x530 & ~x532 & ~x558 & ~x582 & ~x583 & ~x607 & ~x610 & ~x613 & ~x615 & ~x632 & ~x633 & ~x640 & ~x698 & ~x699 & ~x729 & ~x757 & ~x779;
assign c9144 =  x411 & ~x34 & ~x159 & ~x290 & ~x318;
assign c9146 =  x122 &  x149 & ~x56 & ~x130 & ~x131 & ~x135 & ~x156 & ~x185 & ~x212 & ~x529 & ~x556 & ~x606 & ~x607 & ~x618 & ~x673 & ~x760;
assign c9148 = ~x162 & ~x252 & ~x429 & ~x443 & ~x484 & ~x510 & ~x511 & ~x552 & ~x649 & ~x679 & ~x706;
assign c9150 =  x652 & ~x256 & ~x338 & ~x498 & ~x523 & ~x553 & ~x578 & ~x583 & ~x619 & ~x646 & ~x647 & ~x701 & ~x759;
assign c9152 =  x136 &  x293 & ~x274 & ~x303 & ~x331 & ~x416;
assign c9154 =  x87 & ~x309 & ~x576;
assign c9156 =  x199 & ~x176 & ~x232 & ~x260 & ~x473 & ~x477 & ~x505 & ~x530;
assign c9158 = ~x75 & ~x157 & ~x158 & ~x280 & ~x374 & ~x401 & ~x429 & ~x509 & ~x511 & ~x524 & ~x567 & ~x579 & ~x607 & ~x706;
assign c9160 =  x414 &  x741 & ~x133 & ~x241 & ~x249 & ~x510 & ~x524 & ~x550 & ~x552 & ~x553 & ~x554 & ~x580 & ~x607 & ~x634 & ~x636 & ~x666;
assign c9162 =  x146 &  x324 & ~x26 & ~x179 & ~x390 & ~x477 & ~x547 & ~x759;
assign c9164 = ~x45 & ~x47 & ~x72 & ~x131 & ~x132 & ~x182 & ~x443 & ~x453 & ~x496 & ~x499 & ~x534 & ~x559 & ~x642 & ~x669 & ~x671 & ~x702 & ~x704 & ~x713 & ~x724 & ~x781;
assign c9166 =  x379 & ~x2 & ~x7 & ~x25 & ~x26 & ~x29 & ~x32 & ~x53 & ~x70 & ~x71 & ~x97 & ~x262 & ~x291 & ~x363 & ~x416 & ~x472 & ~x473 & ~x502 & ~x503 & ~x507 & ~x530 & ~x534 & ~x559 & ~x561 & ~x589 & ~x737 & ~x764;
assign c9168 =  x433 & ~x2 & ~x12 & ~x13 & ~x52 & ~x56 & ~x70 & ~x71 & ~x413 & ~x416 & ~x418 & ~x420 & ~x444 & ~x449 & ~x470 & ~x504 & ~x507 & ~x526 & ~x588 & ~x643 & ~x672 & ~x674 & ~x731 & ~x736 & ~x766 & ~x767 & ~x782;
assign c9170 =  x87 & ~x449 & ~x603;
assign c9172 =  x468 & ~x245 & ~x303 & ~x360 & ~x417 & ~x445 & ~x446 & ~x474 & ~x505 & ~x588 & ~x626 & ~x635 & ~x661 & ~x691 & ~x707 & ~x735 & ~x763;
assign c9174 = ~x124 & ~x129 & ~x207 & ~x216 & ~x234 & ~x235 & ~x392 & ~x446 & ~x472 & ~x499 & ~x505 & ~x527 & ~x532 & ~x556 & ~x585 & ~x670 & ~x682 & ~x697 & ~x699 & ~x763 & ~x772;
assign c9176 = ~x18 & ~x25 & ~x31 & ~x55 & ~x112 & ~x168 & ~x386 & ~x443 & ~x444 & ~x446 & ~x447 & ~x474 & ~x500 & ~x504 & ~x529 & ~x556 & ~x560 & ~x614 & ~x642 & ~x681 & ~x709 & ~x712 & ~x716 & ~x717 & ~x742 & ~x747 & ~x765 & ~x766 & ~x769 & ~x770 & ~x774;
assign c9178 = ~x15 & ~x25 & ~x40 & ~x44 & ~x66 & ~x68 & ~x106 & ~x120 & ~x122 & ~x124 & ~x177 & ~x336 & ~x417 & ~x418 & ~x449 & ~x476 & ~x532 & ~x667 & ~x696 & ~x697 & ~x752 & ~x757 & ~x775;
assign c9180 = ~x2 & ~x123 & ~x234 & ~x444 & ~x479 & ~x504 & ~x505 & ~x506 & ~x507 & ~x531 & ~x532 & ~x534 & ~x558 & ~x559 & ~x560 & ~x682 & ~x691 & ~x712 & ~x713 & ~x715 & ~x717 & ~x729 & ~x737 & ~x739 & ~x740 & ~x741 & ~x744 & ~x757 & ~x764 & ~x765 & ~x776;
assign c9182 = ~x33 & ~x163 & ~x239 & ~x402 & ~x415 & ~x450 & ~x455 & ~x508 & ~x522 & ~x530 & ~x552 & ~x556 & ~x647 & ~x751;
assign c9184 = ~x2 & ~x26 & ~x75 & ~x132 & ~x162 & ~x189 & ~x214 & ~x402 & ~x429 & ~x458 & ~x485 & ~x525 & ~x594 & ~x596 & ~x616 & ~x620 & ~x623 & ~x699 & ~x706 & ~x709 & ~x768;
assign c9186 =  x352 & ~x70 & ~x445 & ~x561 & ~x585 & ~x654 & ~x662 & ~x709 & ~x710 & ~x719 & ~x736 & ~x747 & ~x772 & ~x775;
assign c9188 =  x410 & ~x109 & ~x443 & ~x449 & ~x470 & ~x501 & ~x503 & ~x556 & ~x584 & ~x585 & ~x605 & ~x680 & ~x706 & ~x737 & ~x762;
assign c9190 =  x498 & ~x3 & ~x28 & ~x84 & ~x224 & ~x278 & ~x303 & ~x331 & ~x332 & ~x333 & ~x335 & ~x359 & ~x360 & ~x361 & ~x362 & ~x390 & ~x447 & ~x475 & ~x529 & ~x530 & ~x558 & ~x559 & ~x580 & ~x608 & ~x636 & ~x637 & ~x664 & ~x692 & ~x722 & ~x723 & ~x751;
assign c9192 =  x438 &  x466 &  x637 & ~x441 & ~x470 & ~x499 & ~x527 & ~x556 & ~x606;
assign c9194 = ~x12 & ~x13 & ~x17 & ~x55 & ~x67 & ~x74 & ~x94 & ~x120 & ~x176 & ~x280 & ~x475 & ~x503 & ~x531 & ~x551 & ~x609 & ~x729 & ~x751 & ~x756;
assign c9196 = ~x38 & ~x39 & ~x53 & ~x58 & ~x365 & ~x392 & ~x415 & ~x446 & ~x447 & ~x477 & ~x505 & ~x532 & ~x534 & ~x560 & ~x562 & ~x563 & ~x588 & ~x670 & ~x671 & ~x700 & ~x708 & ~x740 & ~x741 & ~x742 & ~x743 & ~x746 & ~x756 & ~x759 & ~x762 & ~x765 & ~x771 & ~x772 & ~x775 & ~x776 & ~x778 & ~x783;
assign c9198 = ~x135 & ~x186 & ~x242 & ~x243 & ~x430 & ~x454 & ~x456 & ~x475 & ~x484 & ~x526 & ~x537 & ~x538 & ~x552 & ~x555 & ~x557 & ~x586 & ~x591 & ~x677 & ~x703 & ~x763 & ~x765;
assign c9200 =  x212 & ~x111 & ~x168 & ~x206 & ~x252 & ~x331 & ~x359 & ~x361 & ~x387 & ~x388 & ~x392 & ~x417 & ~x477 & ~x504 & ~x531 & ~x579 & ~x662 & ~x664 & ~x720 & ~x736;
assign c9202 = ~x13 & ~x65 & ~x66 & ~x148 & ~x177 & ~x391 & ~x416 & ~x473 & ~x505 & ~x551 & ~x578 & ~x579 & ~x604 & ~x608 & ~x613 & ~x614 & ~x637 & ~x728 & ~x733 & ~x756;
assign c9204 =  x206 &  x414 &  x741 &  x742 & ~x20 & ~x31 & ~x49 & ~x138 & ~x214 & ~x218 & ~x219 & ~x501 & ~x525 & ~x528 & ~x529 & ~x530 & ~x552 & ~x556 & ~x579 & ~x580 & ~x583 & ~x611 & ~x636 & ~x642 & ~x648 & ~x672 & ~x676 & ~x702 & ~x755 & ~x781;
assign c9206 = ~x21 & ~x22 & ~x55 & ~x106 & ~x168 & ~x183 & ~x210 & ~x220 & ~x245 & ~x427 & ~x454 & ~x480 & ~x501 & ~x527 & ~x551 & ~x556 & ~x558 & ~x590 & ~x605 & ~x613 & ~x619 & ~x729 & ~x751;
assign c9208 = ~x16 & ~x26 & ~x66 & ~x122 & ~x132 & ~x148 & ~x149 & ~x175 & ~x203 & ~x204 & ~x205 & ~x231 & ~x232 & ~x330 & ~x387 & ~x388 & ~x392 & ~x415 & ~x418 & ~x445 & ~x446 & ~x447 & ~x473 & ~x474 & ~x477 & ~x502 & ~x587 & ~x615 & ~x643 & ~x750 & ~x757 & ~x758 & ~x763;
assign c9210 = ~x53 & ~x130 & ~x157 & ~x182 & ~x184 & ~x211 & ~x283 & ~x339 & ~x367 & ~x374 & ~x402 & ~x428 & ~x472 & ~x480 & ~x483 & ~x498 & ~x563 & ~x586 & ~x592 & ~x614 & ~x615 & ~x616 & ~x672 & ~x701 & ~x702 & ~x707 & ~x727 & ~x733 & ~x764;
assign c9212 = ~x5 & ~x108 & ~x153 & ~x181 & ~x223 & ~x244 & ~x366 & ~x418 & ~x446 & ~x471 & ~x472 & ~x477 & ~x529 & ~x531 & ~x608 & ~x614 & ~x615 & ~x662 & ~x693;
assign c9214 =  x412 &  x526 & ~x0 & ~x3 & ~x26 & ~x280 & ~x444 & ~x445 & ~x472 & ~x474 & ~x532 & ~x559 & ~x608 & ~x635 & ~x654 & ~x655 & ~x691 & ~x693 & ~x721;
assign c9216 =  x220 &  x325 & ~x52 & ~x179 & ~x335 & ~x359;
assign c9218 =  x744 &  x745 & ~x46 & ~x55 & ~x111 & ~x138 & ~x195 & ~x222 & ~x420 & ~x485 & ~x539 & ~x566 & ~x580 & ~x611 & ~x620 & ~x633 & ~x645 & ~x672 & ~x705 & ~x756;
assign c9220 =  x302 & ~x24 & ~x44 & ~x45 & ~x49 & ~x76 & ~x78 & ~x105 & ~x107 & ~x130 & ~x132 & ~x133 & ~x136 & ~x159 & ~x191 & ~x195 & ~x416 & ~x417 & ~x418 & ~x441 & ~x442 & ~x444 & ~x445 & ~x449 & ~x470 & ~x472 & ~x473 & ~x477 & ~x498 & ~x502 & ~x505 & ~x586 & ~x590 & ~x645 & ~x701 & ~x728 & ~x730 & ~x755 & ~x783;
assign c9222 = ~x16 & ~x20 & ~x21 & ~x43 & ~x49 & ~x75 & ~x97 & ~x125 & ~x127 & ~x153 & ~x309 & ~x367 & ~x395 & ~x410 & ~x415 & ~x440 & ~x497 & ~x499 & ~x505 & ~x528 & ~x535 & ~x555 & ~x561 & ~x562 & ~x583 & ~x586 & ~x615 & ~x646 & ~x667 & ~x670 & ~x697 & ~x701 & ~x728 & ~x729;
assign c9224 =  x211 &  x496 & ~x302 & ~x362 & ~x445 & ~x587 & ~x596 & ~x635 & ~x707;
assign c9226 =  x295 &  x323 &  x466 & ~x3 & ~x27 & ~x359 & ~x360 & ~x387 & ~x388 & ~x391 & ~x415 & ~x476 & ~x503 & ~x530 & ~x532 & ~x557 & ~x559 & ~x587 & ~x662 & ~x683 & ~x737 & ~x738 & ~x765;
assign c9228 =  x432 &  x460 & ~x29 & ~x45 & ~x181 & ~x443 & ~x470 & ~x472 & ~x478 & ~x499 & ~x556 & ~x557 & ~x561 & ~x563 & ~x590 & ~x615 & ~x616 & ~x701 & ~x726 & ~x755 & ~x764 & ~x773 & ~x775 & ~x783;
assign c9230 = ~x9 & ~x10 & ~x18 & ~x21 & ~x35 & ~x37 & ~x44 & ~x49 & ~x51 & ~x65 & ~x108 & ~x132 & ~x160 & ~x183 & ~x211 & ~x239 & ~x392 & ~x393 & ~x481 & ~x535 & ~x562 & ~x564 & ~x588 & ~x592 & ~x617 & ~x620 & ~x647 & ~x674 & ~x700 & ~x738 & ~x754 & ~x774 & ~x776;
assign c9232 =  x239 & ~x2 & ~x71 & ~x178 & ~x224 & ~x234 & ~x306 & ~x334 & ~x336 & ~x359 & ~x388 & ~x418 & ~x501 & ~x505 & ~x529 & ~x587 & ~x604 & ~x671;
assign c9234 =  x708 & ~x13 & ~x159 & ~x336 & ~x577 & ~x631 & ~x753;
assign c9236 =  x268 &  x382 &  x468 & ~x317 & ~x663;
assign c9238 = ~x47 & ~x109 & ~x214 & ~x346 & ~x347 & ~x374 & ~x402 & ~x428 & ~x446 & ~x553 & ~x579 & ~x639 & ~x731;
assign c9240 =  x109 & ~x151 & ~x152 & ~x219 & ~x248 & ~x249 & ~x276 & ~x277 & ~x278 & ~x304 & ~x343 & ~x361;
assign c9242 = ~x7 & ~x10 & ~x18 & ~x36 & ~x63 & ~x79 & ~x97 & ~x182 & ~x336 & ~x365 & ~x367 & ~x447 & ~x450 & ~x470 & ~x471 & ~x503 & ~x504 & ~x506 & ~x534 & ~x562 & ~x590 & ~x709 & ~x738 & ~x762 & ~x771 & ~x772 & ~x774;
assign c9244 = ~x26 & ~x54 & ~x55 & ~x79 & ~x99 & ~x100 & ~x109 & ~x125 & ~x127 & ~x136 & ~x139 & ~x152 & ~x184 & ~x262 & ~x291 & ~x338 & ~x364 & ~x395 & ~x421 & ~x480 & ~x500 & ~x535 & ~x583 & ~x587 & ~x673 & ~x697 & ~x725 & ~x781 & ~x782;
assign c9246 = ~x74 & ~x157 & ~x186 & ~x428 & ~x500 & ~x526 & ~x552 & ~x576 & ~x605 & ~x729;
assign c9248 =  x385 & ~x57 & ~x304 & ~x306 & ~x333 & ~x334 & ~x419 & ~x420 & ~x447 & ~x572 & ~x580 & ~x600 & ~x608 & ~x609 & ~x627 & ~x629 & ~x634 & ~x658 & ~x659 & ~x666 & ~x693 & ~x722;
assign c9250 = ~x71 & ~x183 & ~x372 & ~x417 & ~x443 & ~x466 & ~x667;
assign c9252 = ~x3 & ~x24 & ~x25 & ~x26 & ~x28 & ~x31 & ~x59 & ~x83 & ~x85 & ~x113 & ~x224 & ~x254 & ~x305 & ~x307 & ~x308 & ~x334 & ~x361 & ~x362 & ~x363 & ~x389 & ~x390 & ~x391 & ~x416 & ~x418 & ~x420 & ~x445 & ~x447 & ~x448 & ~x472 & ~x474 & ~x501 & ~x502 & ~x503 & ~x504 & ~x515 & ~x558 & ~x559 & ~x569 & ~x570 & ~x587 & ~x597 & ~x605 & ~x606 & ~x624 & ~x633 & ~x634 & ~x635 & ~x664 & ~x679 & ~x692 & ~x734 & ~x761;
assign c9254 =  x739 &  x744 & ~x231 & ~x353 & ~x607 & ~x699;
assign c9256 = ~x0 & ~x6 & ~x34 & ~x87 & ~x112 & ~x197 & ~x280 & ~x317 & ~x334 & ~x362 & ~x389 & ~x421 & ~x448 & ~x504 & ~x515 & ~x551 & ~x602 & ~x631 & ~x665 & ~x722 & ~x735 & ~x736 & ~x763;
assign c9258 = ~x9 & ~x15 & ~x16 & ~x41 & ~x42 & ~x70 & ~x71 & ~x72 & ~x84 & ~x101 & ~x152 & ~x153 & ~x223 & ~x309 & ~x392 & ~x419 & ~x420 & ~x421 & ~x472 & ~x477 & ~x498 & ~x505 & ~x524 & ~x547 & ~x556 & ~x557 & ~x583 & ~x584 & ~x611 & ~x613 & ~x615 & ~x616 & ~x640 & ~x644 & ~x671 & ~x697 & ~x701 & ~x754 & ~x755 & ~x780;
assign c9260 =  x355 & ~x76 & ~x158 & ~x215 & ~x397 & ~x416 & ~x442 & ~x445 & ~x469 & ~x498 & ~x500 & ~x616 & ~x729 & ~x758;
assign c9262 = ~x2 & ~x64 & ~x90 & ~x98 & ~x140 & ~x152 & ~x262 & ~x418 & ~x419 & ~x473 & ~x533 & ~x585 & ~x681 & ~x682 & ~x735 & ~x772 & ~x775;
assign c9264 =  x294 & ~x17 & ~x18 & ~x26 & ~x46 & ~x55 & ~x71 & ~x74 & ~x76 & ~x112 & ~x126 & ~x334 & ~x335 & ~x360 & ~x361 & ~x363 & ~x387 & ~x415 & ~x416 & ~x444 & ~x446 & ~x475 & ~x502 & ~x528 & ~x561 & ~x699 & ~x737 & ~x753 & ~x757 & ~x759 & ~x782 & ~x783;
assign c9266 = ~x93 & ~x133 & ~x212 & ~x391 & ~x415 & ~x449 & ~x450 & ~x565;
assign c9268 = ~x72 & ~x185 & ~x186 & ~x373 & ~x400 & ~x455 & ~x482 & ~x522 & ~x523 & ~x526 & ~x548 & ~x670;
assign c9270 =  x519 & ~x133 & ~x162 & ~x271 & ~x280 & ~x298 & ~x430 & ~x431 & ~x446 & ~x457 & ~x512 & ~x530 & ~x539 & ~x559 & ~x606 & ~x705 & ~x734;
assign c9272 = ~x0 & ~x13 & ~x47 & ~x51 & ~x52 & ~x55 & ~x102 & ~x103 & ~x131 & ~x134 & ~x158 & ~x161 & ~x163 & ~x164 & ~x168 & ~x186 & ~x187 & ~x190 & ~x191 & ~x194 & ~x195 & ~x215 & ~x222 & ~x223 & ~x238 & ~x248 & ~x266 & ~x276 & ~x282 & ~x296 & ~x308 & ~x309 & ~x312 & ~x364 & ~x528 & ~x582 & ~x586 & ~x589 & ~x638 & ~x667 & ~x697 & ~x701 & ~x722 & ~x727 & ~x774 & ~x775 & ~x778 & ~x781;
assign c9274 = ~x55 & ~x83 & ~x244 & ~x252 & ~x305 & ~x307 & ~x308 & ~x336 & ~x358 & ~x392 & ~x447 & ~x477 & ~x500 & ~x502 & ~x504 & ~x558 & ~x587 & ~x626 & ~x633 & ~x680 & ~x681 & ~x686 & ~x708 & ~x711 & ~x712 & ~x714 & ~x716 & ~x741 & ~x757;
assign c9276 =  x275 & ~x73 & ~x78 & ~x82 & ~x105 & ~x109 & ~x186 & ~x360 & ~x385 & ~x390 & ~x413 & ~x416 & ~x417 & ~x471 & ~x532;
assign c9278 =  x438 & ~x24 & ~x27 & ~x55 & ~x139 & ~x223 & ~x281 & ~x301 & ~x307 & ~x331 & ~x333 & ~x476 & ~x477 & ~x528 & ~x532 & ~x562 & ~x586 & ~x606 & ~x627 & ~x630 & ~x634 & ~x661 & ~x662 & ~x670 & ~x689 & ~x691;
assign c9280 = ~x13 & ~x15 & ~x21 & ~x98 & ~x127 & ~x128 & ~x153 & ~x155 & ~x168 & ~x182 & ~x336 & ~x392 & ~x395 & ~x420 & ~x426 & ~x441 & ~x443 & ~x452 & ~x473 & ~x500 & ~x526 & ~x620 & ~x732;
assign c9282 =  x623 & ~x212 & ~x251 & ~x280 & ~x523 & ~x527 & ~x547 & ~x548 & ~x549 & ~x552 & ~x555 & ~x584 & ~x603 & ~x610 & ~x645 & ~x696;
assign c9284 = ~x48 & ~x74 & ~x223 & ~x259 & ~x279 & ~x287 & ~x308 & ~x314 & ~x342 & ~x579 & ~x586 & ~x594 & ~x603 & ~x604 & ~x605 & ~x607 & ~x632 & ~x661 & ~x733 & ~x783;
assign c9286 = ~x77 & ~x100 & ~x153 & ~x154 & ~x372 & ~x425 & ~x471 & ~x475 & ~x497 & ~x507 & ~x564 & ~x590 & ~x763 & ~x764 & ~x781;
assign c9288 =  x744 & ~x104 & ~x107 & ~x210 & ~x229 & ~x401 & ~x501 & ~x508 & ~x581;
assign c9290 = ~x12 & ~x80 & ~x111 & ~x195 & ~x392 & ~x402 & ~x429 & ~x483 & ~x508 & ~x525 & ~x527 & ~x540 & ~x579 & ~x623 & ~x676 & ~x724 & ~x735 & ~x760;
assign c9292 = ~x3 & ~x31 & ~x196 & ~x206 & ~x217 & ~x233 & ~x302 & ~x331 & ~x389 & ~x418 & ~x487 & ~x504 & ~x515 & ~x530 & ~x558 & ~x615 & ~x625 & ~x651 & ~x652 & ~x690 & ~x775;
assign c9294 =  x382 & ~x43 & ~x45 & ~x47 & ~x208 & ~x215 & ~x500 & ~x523 & ~x552 & ~x702 & ~x781;
assign c9296 = ~x5 & ~x179 & ~x217 & ~x234 & ~x246 & ~x275 & ~x316 & ~x331 & ~x364 & ~x416 & ~x445 & ~x473 & ~x559 & ~x560 & ~x570 & ~x573 & ~x574 & ~x597 & ~x599 & ~x615 & ~x652 & ~x679 & ~x681 & ~x706 & ~x708;
assign c9298 = ~x5 & ~x7 & ~x31 & ~x57 & ~x60 & ~x86 & ~x112 & ~x252 & ~x305 & ~x333 & ~x361 & ~x363 & ~x389 & ~x417 & ~x419 & ~x445 & ~x446 & ~x447 & ~x459 & ~x474 & ~x487 & ~x513 & ~x540 & ~x597 & ~x606 & ~x623 & ~x625 & ~x633 & ~x662 & ~x677 & ~x679 & ~x704 & ~x706 & ~x759;
assign c9300 =  x212 &  x440 & ~x234 & ~x417 & ~x579 & ~x607 & ~x662 & ~x708 & ~x735;
assign c9302 =  x739 &  x769 & ~x326 & ~x352 & ~x532 & ~x606;
assign c9304 =  x144 &  x404 & ~x27 & ~x43 & ~x414 & ~x417 & ~x443 & ~x477 & ~x529 & ~x586;
assign c9306 =  x262 &  x289 &  x743 & ~x51 & ~x241 & ~x475 & ~x552 & ~x609 & ~x635 & ~x669 & ~x673;
assign c9308 =  x125 &  x519 & ~x46 & ~x83 & ~x85 & ~x134 & ~x161 & ~x164 & ~x167 & ~x222 & ~x258 & ~x266 & ~x272 & ~x278 & ~x280 & ~x285 & ~x296 & ~x298 & ~x310 & ~x313 & ~x324 & ~x338 & ~x340 & ~x448 & ~x501 & ~x580 & ~x582 & ~x593 & ~x611 & ~x620 & ~x646 & ~x647 & ~x648 & ~x697 & ~x698 & ~x703 & ~x782;
assign c9310 = ~x2 & ~x6 & ~x14 & ~x31 & ~x56 & ~x79 & ~x81 & ~x83 & ~x108 & ~x131 & ~x136 & ~x141 & ~x162 & ~x163 & ~x166 & ~x191 & ~x195 & ~x197 & ~x198 & ~x212 & ~x213 & ~x218 & ~x219 & ~x225 & ~x226 & ~x237 & ~x249 & ~x250 & ~x256 & ~x283 & ~x295 & ~x335 & ~x337 & ~x475 & ~x500 & ~x501 & ~x524 & ~x531 & ~x553 & ~x557 & ~x558 & ~x580 & ~x582 & ~x585 & ~x609 & ~x612 & ~x613 & ~x615 & ~x619 & ~x620 & ~x645 & ~x668 & ~x670 & ~x693 & ~x694 & ~x726 & ~x780 & ~x782;
assign c9312 =  x738 &  x740 & ~x213 & ~x214 & ~x215 & ~x216 & ~x257 & ~x266 & ~x268 & ~x279 & ~x295 & ~x529 & ~x553 & ~x577 & ~x580 & ~x584 & ~x604 & ~x617 & ~x728 & ~x731 & ~x732;
assign c9314 =  x381 &  x495 &  x695 & ~x692;
assign c9316 =  x324 & ~x28 & ~x140 & ~x170 & ~x223 & ~x234 & ~x262 & ~x357 & ~x362 & ~x393 & ~x415 & ~x416 & ~x420 & ~x421 & ~x441 & ~x445 & ~x475 & ~x527 & ~x531 & ~x556 & ~x587 & ~x641 & ~x643 & ~x698 & ~x700 & ~x707 & ~x709 & ~x735 & ~x764 & ~x783;
assign c9318 = ~x15 & ~x100 & ~x107 & ~x152 & ~x180 & ~x210 & ~x239 & ~x263 & ~x295 & ~x421 & ~x450 & ~x479 & ~x526 & ~x533 & ~x563 & ~x589 & ~x702 & ~x728 & ~x756 & ~x777;
assign c9320 = ~x1 & ~x3 & ~x18 & ~x29 & ~x55 & ~x59 & ~x87 & ~x364 & ~x431 & ~x446 & ~x472 & ~x486 & ~x513 & ~x531 & ~x540 & ~x550 & ~x559 & ~x569 & ~x578 & ~x595 & ~x607 & ~x624 & ~x635 & ~x661 & ~x664;
assign c9322 =  x415 & ~x26 & ~x80 & ~x107 & ~x164 & ~x190 & ~x223 & ~x272 & ~x273 & ~x274 & ~x295 & ~x296 & ~x298 & ~x558 & ~x583 & ~x592 & ~x609;
assign c9324 =  x303 & ~x24 & ~x27 & ~x49 & ~x77 & ~x83 & ~x105 & ~x106 & ~x108 & ~x109 & ~x161 & ~x162 & ~x166 & ~x167 & ~x189 & ~x367 & ~x391 & ~x422 & ~x423 & ~x442 & ~x443 & ~x445 & ~x446 & ~x447 & ~x449 & ~x471 & ~x501 & ~x502 & ~x530 & ~x560 & ~x587 & ~x614 & ~x615 & ~x616 & ~x644 & ~x645 & ~x672 & ~x675 & ~x699 & ~x702 & ~x728;
assign c9326 =  x467 & ~x7 & ~x8 & ~x10 & ~x191 & ~x308 & ~x361 & ~x447 & ~x474 & ~x587 & ~x626 & ~x634 & ~x662 & ~x664 & ~x692;
assign c9328 = ~x8 & ~x21 & ~x44 & ~x45 & ~x48 & ~x51 & ~x53 & ~x68 & ~x78 & ~x80 & ~x94 & ~x136 & ~x156 & ~x183 & ~x212 & ~x241 & ~x425 & ~x499 & ~x562 & ~x640 & ~x759;
assign c9330 = ~x25 & ~x26 & ~x71 & ~x152 & ~x164 & ~x179 & ~x187 & ~x235 & ~x243 & ~x265 & ~x292 & ~x426 & ~x448 & ~x472 & ~x474 & ~x507 & ~x533 & ~x535 & ~x640 & ~x699 & ~x728 & ~x764;
assign c9332 = ~x153 & ~x154 & ~x284 & ~x313 & ~x342 & ~x492 & ~x495 & ~x498 & ~x523 & ~x551 & ~x554 & ~x579 & ~x605 & ~x607 & ~x612 & ~x615 & ~x753;
assign c9334 =  x246 &  x379 & ~x24 & ~x51 & ~x101 & ~x103 & ~x106 & ~x390 & ~x413 & ~x414 & ~x415 & ~x443 & ~x448 & ~x470 & ~x471 & ~x532 & ~x561 & ~x587 & ~x644 & ~x671;
assign c9336 =  x97 & ~x4 & ~x18 & ~x79 & ~x106 & ~x141 & ~x162 & ~x163 & ~x221 & ~x429 & ~x456 & ~x458 & ~x511 & ~x558 & ~x580 & ~x610 & ~x621;
assign c9338 = ~x9 & ~x78 & ~x84 & ~x105 & ~x245 & ~x246 & ~x248 & ~x251 & ~x267 & ~x273 & ~x296 & ~x339 & ~x429 & ~x458 & ~x528 & ~x530 & ~x534 & ~x538 & ~x539 & ~x554 & ~x555 & ~x566 & ~x581 & ~x612 & ~x614 & ~x622 & ~x645 & ~x648 & ~x672 & ~x678 & ~x697 & ~x704 & ~x732 & ~x760;
assign c9340 =  x487 & ~x83 & ~x307 & ~x359 & ~x360 & ~x473 & ~x562 & ~x713 & ~x714 & ~x716 & ~x736 & ~x746;
assign c9342 =  x263 & ~x163 & ~x192 & ~x267 & ~x309 & ~x325 & ~x457 & ~x458 & ~x511 & ~x532 & ~x539 & ~x554 & ~x566 & ~x608;
assign c9344 = ~x32 & ~x46 & ~x250 & ~x251 & ~x270 & ~x419 & ~x450 & ~x456 & ~x473 & ~x484 & ~x500 & ~x553 & ~x564 & ~x566 & ~x579 & ~x641 & ~x734 & ~x759 & ~x760;
assign c9346 =  x525 &  x611 &  x696 & ~x636;
assign c9348 =  x566 &  x676 & ~x54 & ~x273 & ~x290 & ~x534 & ~x559 & ~x589 & ~x680 & ~x690;
assign c9350 = ~x197 & ~x279 & ~x282 & ~x291 & ~x303 & ~x308 & ~x318 & ~x336 & ~x362 & ~x392 & ~x393 & ~x420 & ~x473 & ~x506 & ~x561 & ~x627 & ~x654 & ~x659 & ~x661 & ~x682 & ~x689 & ~x709 & ~x711 & ~x739 & ~x741 & ~x766;
assign c9352 =  x485 & ~x22 & ~x28 & ~x55 & ~x56 & ~x83 & ~x126 & ~x252 & ~x308 & ~x317 & ~x386 & ~x391 & ~x445 & ~x474 & ~x500 & ~x501 & ~x529 & ~x557 & ~x558 & ~x585 & ~x586 & ~x590 & ~x640 & ~x701 & ~x726 & ~x728 & ~x758 & ~x774;
assign c9354 =  x429 &  x457 & ~x26 & ~x71 & ~x124 & ~x151 & ~x251 & ~x306 & ~x334 & ~x363 & ~x364 & ~x395 & ~x396 & ~x421 & ~x422 & ~x452 & ~x476 & ~x477 & ~x478 & ~x479 & ~x503 & ~x506 & ~x529 & ~x557 & ~x559 & ~x561 & ~x612 & ~x613 & ~x615 & ~x617 & ~x618 & ~x642 & ~x645 & ~x699 & ~x702 & ~x728 & ~x756 & ~x758 & ~x782;
assign c9356 =  x414 &  x490 & ~x107 & ~x222 & ~x240 & ~x511 & ~x537 & ~x580 & ~x581 & ~x584;
assign c9358 =  x549 & ~x28 & ~x29 & ~x51 & ~x106 & ~x308 & ~x413 & ~x442 & ~x480 & ~x591 & ~x618 & ~x682 & ~x737 & ~x738 & ~x739 & ~x770;
assign c9360 =  x711 & ~x47 & ~x73 & ~x99 & ~x101 & ~x282 & ~x310 & ~x311 & ~x334 & ~x337 & ~x523 & ~x524 & ~x526 & ~x529 & ~x549 & ~x557 & ~x558 & ~x603 & ~x609 & ~x618 & ~x633 & ~x641 & ~x726;
assign c9362 =  x323 & ~x31 & ~x32 & ~x53 & ~x55 & ~x57 & ~x336 & ~x358 & ~x361 & ~x364 & ~x415 & ~x417 & ~x444 & ~x474 & ~x503 & ~x533 & ~x558 & ~x559 & ~x560 & ~x681 & ~x687 & ~x688 & ~x689 & ~x708 & ~x711 & ~x736 & ~x739 & ~x740 & ~x741 & ~x775;
assign c9364 =  x377 &  x405 & ~x2 & ~x16 & ~x55 & ~x73 & ~x84 & ~x140 & ~x141 & ~x252 & ~x280 & ~x302 & ~x331 & ~x332 & ~x333 & ~x360 & ~x361 & ~x362 & ~x364 & ~x389 & ~x390 & ~x418 & ~x419 & ~x446 & ~x447 & ~x474 & ~x475 & ~x502 & ~x503 & ~x505 & ~x571 & ~x663 & ~x692 & ~x737 & ~x777;
assign c9366 =  x172 & ~x25 & ~x105 & ~x122 & ~x177 & ~x473 & ~x502 & ~x587 & ~x678;
assign c9368 = ~x49 & ~x77 & ~x134 & ~x136 & ~x270 & ~x367 & ~x376 & ~x427 & ~x479 & ~x498 & ~x509 & ~x560 & ~x586 & ~x709 & ~x729 & ~x764;
assign c9370 = ~x12 & ~x14 & ~x22 & ~x23 & ~x46 & ~x51 & ~x54 & ~x79 & ~x82 & ~x102 & ~x103 & ~x104 & ~x111 & ~x129 & ~x132 & ~x158 & ~x209 & ~x211 & ~x420 & ~x443 & ~x448 & ~x452 & ~x472 & ~x480 & ~x481 & ~x508 & ~x527 & ~x529 & ~x555 & ~x558 & ~x562 & ~x592 & ~x646 & ~x672 & ~x673 & ~x725 & ~x727 & ~x728 & ~x733 & ~x758 & ~x761 & ~x781;
assign c9372 =  x356 &  x434 & ~x0 & ~x161 & ~x223 & ~x445 & ~x504 & ~x511 & ~x579 & ~x632 & ~x782 & ~x783;
assign c9374 = ~x2 & ~x4 & ~x27 & ~x55 & ~x56 & ~x60 & ~x83 & ~x140 & ~x168 & ~x251 & ~x252 & ~x334 & ~x344 & ~x361 & ~x417 & ~x418 & ~x449 & ~x460 & ~x488 & ~x503 & ~x504 & ~x516 & ~x532 & ~x570 & ~x578 & ~x606 & ~x635 & ~x665 & ~x694 & ~x722;
assign c9376 =  x462 &  x715 &  x747 & ~x133 & ~x342 & ~x529 & ~x593 & ~x620 & ~x706 & ~x734;
assign c9378 =  x263 & ~x243 & ~x251 & ~x283 & ~x284 & ~x286 & ~x294 & ~x312 & ~x324 & ~x567 & ~x578 & ~x580 & ~x593 & ~x608 & ~x615 & ~x619 & ~x637 & ~x648 & ~x667 & ~x695 & ~x762;
assign c9380 =  x494 & ~x27 & ~x28 & ~x29 & ~x54 & ~x84 & ~x130 & ~x138 & ~x140 & ~x250 & ~x251 & ~x252 & ~x308 & ~x332 & ~x333 & ~x335 & ~x336 & ~x337 & ~x356 & ~x359 & ~x364 & ~x392 & ~x419 & ~x421 & ~x449 & ~x501 & ~x503 & ~x527 & ~x528 & ~x531 & ~x556 & ~x558 & ~x585 & ~x612 & ~x633 & ~x640 & ~x669 & ~x670 & ~x671 & ~x688 & ~x690 & ~x782;
assign c9382 = ~x54 & ~x82 & ~x98 & ~x111 & ~x135 & ~x163 & ~x192 & ~x234 & ~x291 & ~x319 & ~x364 & ~x365 & ~x392 & ~x476 & ~x477 & ~x500 & ~x505 & ~x525 & ~x555 & ~x639 & ~x701 & ~x702 & ~x725 & ~x728 & ~x730 & ~x738 & ~x764 & ~x768;
assign c9384 =  x88 & ~x421 & ~x582 & ~x602 & ~x609;
assign c9386 =  x358 & ~x163 & ~x187 & ~x191 & ~x217 & ~x241 & ~x242 & ~x268 & ~x364 & ~x475 & ~x510 & ~x524 & ~x590 & ~x761;
assign c9388 = ~x278 & ~x281 & ~x388 & ~x390 & ~x449 & ~x474 & ~x554 & ~x605 & ~x632 & ~x652 & ~x653 & ~x662 & ~x682 & ~x712 & ~x713 & ~x726 & ~x735 & ~x772;
assign c9390 = ~x21 & ~x27 & ~x99 & ~x308 & ~x309 & ~x310 & ~x337 & ~x357 & ~x358 & ~x391 & ~x394 & ~x416 & ~x419 & ~x420 & ~x421 & ~x442 & ~x443 & ~x444 & ~x449 & ~x476 & ~x477 & ~x479 & ~x532 & ~x535 & ~x584 & ~x585 & ~x586 & ~x617 & ~x717 & ~x727 & ~x741 & ~x744 & ~x769 & ~x774 & ~x776;
assign c9392 =  x351 & ~x69 & ~x72 & ~x96 & ~x126 & ~x386 & ~x418 & ~x473 & ~x503 & ~x534 & ~x617 & ~x739 & ~x743 & ~x745 & ~x757 & ~x774;
assign c9394 =  x376 &  x432 & ~x100 & ~x280 & ~x337 & ~x342 & ~x392 & ~x397 & ~x466 & ~x532 & ~x673 & ~x674;
assign c9396 =  x465 & ~x55 & ~x231 & ~x363 & ~x391 & ~x476 & ~x485 & ~x502 & ~x503 & ~x512 & ~x549 & ~x567 & ~x576 & ~x594 & ~x622 & ~x643 & ~x707 & ~x762;
assign c9398 =  x740 & ~x70 & ~x99 & ~x155 & ~x156 & ~x523 & ~x524 & ~x576 & ~x578 & ~x606 & ~x637 & ~x659 & ~x759;
assign c9400 =  x238 &  x266 &  x427 & ~x37 & ~x301 & ~x303 & ~x304 & ~x305 & ~x330 & ~x331 & ~x358 & ~x387 & ~x448 & ~x472 & ~x473 & ~x474 & ~x500;
assign c9402 =  x480 & ~x56 & ~x86 & ~x217 & ~x247 & ~x248 & ~x276 & ~x304 & ~x305 & ~x333 & ~x363 & ~x502 & ~x559 & ~x579 & ~x587 & ~x633 & ~x634 & ~x635 & ~x636 & ~x664 & ~x721;
assign c9404 =  x708 &  x738 &  x740 &  x741 &  x742 & ~x46 & ~x134 & ~x136 & ~x187 & ~x214 & ~x252 & ~x503 & ~x550 & ~x551 & ~x577 & ~x579 & ~x581 & ~x583 & ~x586 & ~x607 & ~x609 & ~x633 & ~x638 & ~x781;
assign c9406 =  x142 & ~x19 & ~x50 & ~x131 & ~x473 & ~x534 & ~x560 & ~x588 & ~x589 & ~x616 & ~x644 & ~x646 & ~x729 & ~x731 & ~x757 & ~x761;
assign c9408 = ~x4 & ~x27 & ~x140 & ~x235 & ~x252 & ~x275 & ~x279 & ~x280 & ~x310 & ~x335 & ~x390 & ~x391 & ~x449 & ~x475 & ~x531 & ~x533 & ~x580 & ~x600 & ~x628 & ~x633 & ~x634 & ~x657 & ~x658 & ~x662 & ~x691 & ~x711 & ~x720;
assign c9410 =  x545 &  x716 & ~x0 & ~x80 & ~x133 & ~x162 & ~x164 & ~x167 & ~x191 & ~x196 & ~x475 & ~x502 & ~x539 & ~x557 & ~x580 & ~x585 & ~x613 & ~x632 & ~x636 & ~x647 & ~x648 & ~x727;
assign c9412 =  x495 & ~x54 & ~x196 & ~x273 & ~x300 & ~x306 & ~x478 & ~x505 & ~x563 & ~x681 & ~x689 & ~x736 & ~x738 & ~x781;
assign c9414 = ~x210 & ~x399 & ~x442 & ~x453 & ~x464 & ~x471 & ~x479 & ~x505 & ~x521 & ~x646 & ~x701 & ~x775;
assign c9416 = ~x74 & ~x310 & ~x370 & ~x393 & ~x395 & ~x419 & ~x424 & ~x443 & ~x467 & ~x471 & ~x494 & ~x496 & ~x527 & ~x550 & ~x551 & ~x575 & ~x576 & ~x580 & ~x589 & ~x620 & ~x735 & ~x781;
assign c9418 =  x146 & ~x106 & ~x137 & ~x151 & ~x163 & ~x181 & ~x208 & ~x420 & ~x421 & ~x479 & ~x506 & ~x526 & ~x528 & ~x529 & ~x563 & ~x617 & ~x618 & ~x674 & ~x701 & ~x727 & ~x758;
assign c9420 =  x137 &  x591 & ~x246 & ~x275 & ~x276 & ~x304;
assign c9422 =  x466 &  x609 & ~x441 & ~x498 & ~x555 & ~x556 & ~x640 & ~x662;
assign c9424 =  x494 &  x548 & ~x22 & ~x82 & ~x317 & ~x346 & ~x653 & ~x661 & ~x686 & ~x738;
assign c9426 =  x325 &  x352 & ~x16 & ~x43 & ~x44 & ~x48 & ~x70 & ~x76 & ~x78 & ~x101 & ~x103 & ~x157 & ~x184 & ~x413 & ~x414 & ~x441 & ~x442 & ~x443 & ~x446 & ~x471 & ~x473 & ~x498 & ~x505 & ~x646 & ~x701;
assign c9428 = ~x44 & ~x79 & ~x100 & ~x127 & ~x132 & ~x167 & ~x198 & ~x309 & ~x312 & ~x345 & ~x363 & ~x373 & ~x399 & ~x400 & ~x444 & ~x553 & ~x584 & ~x590 & ~x592 & ~x616 & ~x731 & ~x781;
assign c9430 =  x490 &  x545 &  x713 &  x716 & ~x21 & ~x26 & ~x45 & ~x138 & ~x162 & ~x167 & ~x191 & ~x193 & ~x223 & ~x448 & ~x502 & ~x530 & ~x531 & ~x539 & ~x592 & ~x608 & ~x618 & ~x619 & ~x648 & ~x676 & ~x734 & ~x753;
assign c9432 = ~x12 & ~x13 & ~x41 & ~x49 & ~x71 & ~x106 & ~x364 & ~x367 & ~x427 & ~x497 & ~x499 & ~x522 & ~x563 & ~x588 & ~x734 & ~x761;
assign c9434 = ~x31 & ~x57 & ~x130 & ~x159 & ~x272 & ~x279 & ~x301 & ~x336 & ~x445 & ~x447 & ~x448 & ~x473 & ~x500 & ~x528 & ~x533 & ~x585 & ~x615 & ~x644 & ~x672 & ~x681 & ~x685 & ~x686 & ~x698 & ~x712 & ~x728 & ~x744 & ~x745 & ~x764 & ~x775;
assign c9436 =  x238 &  x295 &  x410 & ~x388 & ~x446 & ~x683 & ~x717 & ~x746;
assign c9438 =  x491 & ~x46 & ~x160 & ~x166 & ~x215 & ~x216 & ~x402 & ~x430 & ~x483 & ~x511 & ~x528 & ~x552 & ~x553 & ~x556 & ~x565 & ~x579 & ~x590 & ~x612 & ~x622 & ~x623 & ~x640 & ~x673 & ~x675 & ~x733 & ~x754;
assign c9440 = ~x3 & ~x7 & ~x21 & ~x34 & ~x51 & ~x72 & ~x98 & ~x125 & ~x126 & ~x161 & ~x236 & ~x251 & ~x290 & ~x366 & ~x563 & ~x564 & ~x587 & ~x620 & ~x766 & ~x782;
assign c9442 =  x211 & ~x16 & ~x17 & ~x26 & ~x113 & ~x196 & ~x278 & ~x305 & ~x334 & ~x360 & ~x362 & ~x364 & ~x445 & ~x475 & ~x502 & ~x531 & ~x569 & ~x587 & ~x597 & ~x605 & ~x624 & ~x632 & ~x633 & ~x634 & ~x660 & ~x661 & ~x679 & ~x707 & ~x734 & ~x761;
assign c9444 =  x405 & ~x28 & ~x52 & ~x308 & ~x360 & ~x361 & ~x390 & ~x392 & ~x393 & ~x416 & ~x419 & ~x447 & ~x475 & ~x502 & ~x506 & ~x531 & ~x534 & ~x559 & ~x588 & ~x616 & ~x710 & ~x711 & ~x728 & ~x737 & ~x741 & ~x742 & ~x743 & ~x744 & ~x746 & ~x767 & ~x773 & ~x774;
assign c9446 =  x164 &  x240 & ~x178 & ~x304 & ~x333 & ~x361 & ~x388;
assign c9448 =  x359 & ~x20 & ~x27 & ~x108 & ~x139 & ~x140 & ~x164 & ~x189 & ~x213 & ~x218 & ~x242 & ~x270 & ~x296 & ~x445 & ~x468 & ~x469 & ~x471 & ~x498 & ~x502 & ~x615 & ~x674 & ~x700 & ~x731 & ~x783;
assign c9450 = ~x1 & ~x48 & ~x85 & ~x108 & ~x159 & ~x167 & ~x187 & ~x216 & ~x223 & ~x268 & ~x270 & ~x293 & ~x294 & ~x297 & ~x314 & ~x341 & ~x368 & ~x420 & ~x501 & ~x528 & ~x530 & ~x532 & ~x559 & ~x588 & ~x593 & ~x643 & ~x644 & ~x649 & ~x668 & ~x704 & ~x727 & ~x756;
assign c9452 =  x184 & ~x305 & ~x487 & ~x541 & ~x579 & ~x604 & ~x624 & ~x632 & ~x634 & ~x655;
assign c9454 = ~x6 & ~x19 & ~x23 & ~x67 & ~x79 & ~x133 & ~x150 & ~x152 & ~x211 & ~x364 & ~x421 & ~x562 & ~x584 & ~x724 & ~x772 & ~x774;
assign c9456 = ~x23 & ~x24 & ~x39 & ~x83 & ~x108 & ~x126 & ~x134 & ~x137 & ~x156 & ~x159 & ~x162 & ~x163 & ~x181 & ~x241 & ~x268 & ~x269 & ~x297 & ~x419 & ~x477 & ~x504 & ~x505 & ~x506 & ~x525 & ~x526 & ~x556 & ~x585 & ~x586 & ~x587 & ~x592 & ~x645 & ~x697 & ~x755 & ~x757;
assign c9458 =  x701 & ~x304 & ~x333 & ~x445 & ~x559 & ~x607 & ~x634 & ~x635 & ~x692 & ~x706 & ~x707 & ~x735;
assign c9460 =  x411 & ~x0 & ~x326 & ~x456 & ~x471 & ~x483 & ~x528 & ~x553 & ~x557;
assign c9462 =  x741 & ~x192 & ~x216 & ~x267 & ~x300 & ~x306 & ~x381 & ~x458 & ~x556 & ~x578 & ~x583 & ~x592;
assign c9464 = ~x6 & ~x25 & ~x71 & ~x77 & ~x100 & ~x125 & ~x126 & ~x131 & ~x152 & ~x153 & ~x183 & ~x184 & ~x365 & ~x418 & ~x444 & ~x471 & ~x498 & ~x507 & ~x525 & ~x590 & ~x593 & ~x645 & ~x702 & ~x765 & ~x781 & ~x783;
assign c9466 =  x441 & ~x16 & ~x161 & ~x189 & ~x220 & ~x246 & ~x247 & ~x248 & ~x277 & ~x281 & ~x293 & ~x305 & ~x306 & ~x309 & ~x310 & ~x336 & ~x504 & ~x550 & ~x606 & ~x607 & ~x609 & ~x635 & ~x664 & ~x694 & ~x695 & ~x756;
assign c9468 = ~x4 & ~x27 & ~x49 & ~x74 & ~x105 & ~x107 & ~x108 & ~x136 & ~x157 & ~x160 & ~x161 & ~x186 & ~x210 & ~x310 & ~x343 & ~x362 & ~x366 & ~x391 & ~x394 & ~x396 & ~x453 & ~x530 & ~x536 & ~x585 & ~x586 & ~x589 & ~x590 & ~x591 & ~x611 & ~x614 & ~x674 & ~x754 & ~x763;
assign c9470 =  x81 & ~x98 & ~x259;
assign c9472 =  x488 &  x516 &  x544 & ~x28 & ~x52 & ~x55 & ~x128 & ~x208 & ~x502 & ~x554 & ~x561 & ~x616 & ~x618 & ~x639 & ~x727;
assign c9474 = ~x8 & ~x55 & ~x140 & ~x216 & ~x363 & ~x416 & ~x532 & ~x586 & ~x597 & ~x599 & ~x633 & ~x656 & ~x659 & ~x747;
assign c9476 = ~x4 & ~x73 & ~x77 & ~x82 & ~x103 & ~x105 & ~x106 & ~x126 & ~x131 & ~x136 & ~x155 & ~x184 & ~x370 & ~x495 & ~x534 & ~x582 & ~x583 & ~x723 & ~x750 & ~x756 & ~x779;
assign c9478 =  x715 & ~x105 & ~x167 & ~x374 & ~x455 & ~x576;
assign c9480 = ~x103 & ~x178 & ~x262 & ~x417 & ~x421 & ~x448 & ~x474 & ~x506 & ~x507 & ~x563 & ~x588 & ~x644 & ~x672 & ~x681 & ~x737 & ~x739 & ~x742 & ~x745 & ~x746 & ~x768;
assign c9482 =  x407 & ~x7 & ~x79 & ~x137 & ~x182 & ~x186 & ~x187 & ~x209 & ~x211 & ~x213 & ~x216 & ~x239 & ~x444 & ~x470 & ~x471 & ~x472 & ~x481 & ~x499 & ~x644 & ~x724;
assign c9484 =  x582 &  x610 & ~x252 & ~x472 & ~x500 & ~x585 & ~x625 & ~x636 & ~x662 & ~x693;
assign c9486 =  x143 &  x349 & ~x418 & ~x446 & ~x447 & ~x473 & ~x474 & ~x475 & ~x477 & ~x501 & ~x503 & ~x504 & ~x706 & ~x707 & ~x728;
assign c9488 = ~x74 & ~x108 & ~x339 & ~x346 & ~x483 & ~x565 & ~x593 & ~x607 & ~x636 & ~x708;
assign c9490 =  x331 & ~x1 & ~x16 & ~x24 & ~x51 & ~x76 & ~x79 & ~x81 & ~x107 & ~x109 & ~x110 & ~x111 & ~x112 & ~x133 & ~x138 & ~x160 & ~x162 & ~x165 & ~x186 & ~x187 & ~x188 & ~x189 & ~x192 & ~x193 & ~x194 & ~x241 & ~x364 & ~x392 & ~x421 & ~x442 & ~x443 & ~x446 & ~x447 & ~x469 & ~x471 & ~x472 & ~x474 & ~x501 & ~x532 & ~x560 & ~x590 & ~x617 & ~x644 & ~x646 & ~x647 & ~x672 & ~x673 & ~x674 & ~x675 & ~x700 & ~x701 & ~x702 & ~x727 & ~x728 & ~x730 & ~x756 & ~x764 & ~x781 & ~x783;
assign c9492 =  x377 & ~x21 & ~x55 & ~x335 & ~x346 & ~x358 & ~x363 & ~x392 & ~x417 & ~x419 & ~x444 & ~x448 & ~x474 & ~x503 & ~x534 & ~x560 & ~x663 & ~x690;
assign c9494 =  x137 & ~x178 & ~x275 & ~x276 & ~x304 & ~x363 & ~x628;
assign c9496 =  x323 &  x351 &  x379 &  x485 & ~x26 & ~x206 & ~x234 & ~x262 & ~x473 & ~x532;
assign c9498 = ~x124 & ~x261 & ~x303 & ~x304 & ~x360 & ~x392 & ~x417 & ~x418 & ~x444 & ~x473 & ~x501 & ~x502 & ~x504 & ~x531 & ~x608 & ~x643 & ~x692 & ~x693 & ~x707 & ~x714 & ~x749;
assign c91 = ~x92 & ~x229 & ~x230 & ~x231 & ~x256 & ~x258 & ~x260 & ~x281 & ~x288 & ~x312 & ~x333 & ~x358 & ~x372 & ~x398 & ~x399 & ~x424 & ~x444 & ~x470 & ~x484;
assign c93 =  x582 & ~x25 & ~x56 & ~x103 & ~x113 & ~x167 & ~x223 & ~x225 & ~x249;
assign c95 =  x294 & ~x50 & ~x115 & ~x177 & ~x230 & ~x258 & ~x634 & ~x690;
assign c97 =  x408 &  x457 & ~x88 & ~x143 & ~x191 & ~x201 & ~x494 & ~x508;
assign c99 = ~x30 & ~x31 & ~x82 & ~x139 & ~x223 & ~x236 & ~x436 & ~x492 & ~x575 & ~x738;
assign c911 = ~x356 & ~x357 & ~x693 & ~x694 & ~x750;
assign c913 =  x505 & ~x742;
assign c915 =  x292 & ~x3 & ~x80 & ~x108 & ~x138 & ~x154 & ~x242 & ~x304 & ~x388 & ~x668;
assign c917 = ~x17 & ~x19 & ~x25 & ~x33 & ~x114 & ~x143 & ~x165 & ~x193 & ~x195 & ~x220 & ~x250 & ~x255 & ~x515 & ~x516 & ~x518 & ~x559 & ~x704;
assign c919 = ~x22 & ~x81 & ~x82 & ~x84 & ~x167 & ~x250 & ~x379 & ~x406 & ~x445 & ~x462 & ~x545 & ~x546 & ~x572 & ~x573 & ~x603 & ~x658;
assign c921 =  x607 & ~x408;
assign c923 =  x554 & ~x213 & ~x668;
assign c925 =  x661 & ~x15 & ~x23 & ~x58 & ~x140 & ~x144 & ~x166 & ~x170 & ~x192 & ~x224 & ~x225 & ~x249 & ~x251 & ~x252 & ~x280 & ~x305 & ~x361 & ~x390 & ~x391 & ~x420 & ~x447 & ~x474 & ~x476 & ~x501 & ~x504 & ~x558 & ~x560 & ~x585 & ~x586 & ~x616 & ~x783;
assign c927 = ~x27 & ~x34 & ~x140 & ~x168 & ~x169 & ~x382 & ~x410 & ~x432 & ~x439 & ~x466 & ~x495;
assign c929 =  x307;
assign c931 =  x322 &  x349 & ~x142 & ~x227 & ~x303 & ~x313 & ~x329 & ~x498;
assign c933 =  x241 &  x361;
assign c935 = ~x24 & ~x33 & ~x47 & ~x80 & ~x89 & ~x106 & ~x118 & ~x131 & ~x143 & ~x144 & ~x187 & ~x199 & ~x201 & ~x217 & ~x218 & ~x220 & ~x231 & ~x232 & ~x244 & ~x256 & ~x260 & ~x271 & ~x300 & ~x302 & ~x308 & ~x315 & ~x356 & ~x358 & ~x360 & ~x365 & ~x370 & ~x387 & ~x388 & ~x414 & ~x415 & ~x418 & ~x419 & ~x422 & ~x442 & ~x443 & ~x444 & ~x451 & ~x478 & ~x498 & ~x501 & ~x508 & ~x554 & ~x564 & ~x590 & ~x617 & ~x618 & ~x619 & ~x643 & ~x669 & ~x696 & ~x698 & ~x723;
assign c937 =  x67 &  x182 & ~x369 & ~x416 & ~x480 & ~x504 & ~x535;
assign c939 =  x184 & ~x57 & ~x77 & ~x106 & ~x107 & ~x108 & ~x114 & ~x136 & ~x163 & ~x191 & ~x198 & ~x199 & ~x290 & ~x727 & ~x777;
assign c941 =  x342 &  x370 &  x426 & ~x3 & ~x20 & ~x29 & ~x56 & ~x57 & ~x82 & ~x86 & ~x168 & ~x475 & ~x503 & ~x584 & ~x613 & ~x642 & ~x670 & ~x699 & ~x701 & ~x704 & ~x725 & ~x752 & ~x756;
assign c943 = ~x19 & ~x22 & ~x24 & ~x27 & ~x28 & ~x52 & ~x54 & ~x55 & ~x81 & ~x82 & ~x83 & ~x85 & ~x110 & ~x112 & ~x113 & ~x139 & ~x141 & ~x167 & ~x168 & ~x195 & ~x221 & ~x224 & ~x242 & ~x250 & ~x251 & ~x307 & ~x335 & ~x392 & ~x410 & ~x438 & ~x439 & ~x449 & ~x468 & ~x494 & ~x496 & ~x644 & ~x687 & ~x754 & ~x755 & ~x756 & ~x783;
assign c945 =  x216 & ~x321 & ~x431;
assign c947 = ~x26 & ~x114 & ~x188 & ~x190 & ~x201 & ~x218 & ~x222 & ~x226 & ~x229 & ~x233 & ~x250 & ~x261 & ~x272 & ~x301 & ~x303 & ~x366 & ~x470 & ~x497 & ~x509 & ~x536 & ~x560 & ~x561 & ~x618 & ~x637 & ~x644 & ~x690 & ~x692 & ~x753 & ~x756 & ~x777 & ~x782;
assign c949 =  x272 & ~x53 & ~x195 & ~x406 & ~x561 & ~x755;
assign c951 =  x264 & ~x24 & ~x110 & ~x167 & ~x196 & ~x224 & ~x335 & ~x349 & ~x350 & ~x474 & ~x507 & ~x535 & ~x546 & ~x756;
assign c953 = ~x3 & ~x24 & ~x56 & ~x85 & ~x236 & ~x271 & ~x272 & ~x328 & ~x355 & ~x383 & ~x385 & ~x394 & ~x411 & ~x412 & ~x413 & ~x440 & ~x469 & ~x503 & ~x588 & ~x595 & ~x670 & ~x673 & ~x755 & ~x756 & ~x760 & ~x783;
assign c955 = ~x20 & ~x23 & ~x31 & ~x75 & ~x76 & ~x81 & ~x86 & ~x105 & ~x141 & ~x167 & ~x170 & ~x253 & ~x606 & ~x673 & ~x679 & ~x688 & ~x699 & ~x703 & ~x704 & ~x707 & ~x716 & ~x727 & ~x729 & ~x744 & ~x751 & ~x753 & ~x760 & ~x761 & ~x780 & ~x782;
assign c957 =  x528 & ~x187 & ~x214;
assign c959 = ~x35 & ~x92 & ~x112 & ~x113 & ~x114 & ~x115 & ~x119 & ~x148 & ~x172 & ~x173 & ~x176 & ~x590 & ~x603 & ~x604 & ~x709 & ~x731;
assign c961 =  x187 & ~x320 & ~x321 & ~x526 & ~x588;
assign c963 =  x317 &  x379 & ~x26 & ~x110 & ~x138 & ~x192 & ~x196 & ~x199 & ~x246 & ~x276 & ~x359 & ~x360 & ~x361 & ~x370;
assign c965 =  x408 &  x460 & ~x243 & ~x274 & ~x299 & ~x327 & ~x386 & ~x387;
assign c967 =  x464 & ~x115 & ~x342 & ~x537 & ~x564 & ~x636 & ~x689 & ~x690 & ~x697 & ~x746 & ~x747;
assign c969 = ~x55 & ~x58 & ~x84 & ~x85 & ~x87 & ~x335 & ~x391 & ~x439 & ~x465 & ~x467 & ~x494 & ~x504 & ~x541 & ~x542 & ~x551 & ~x570 & ~x682 & ~x738 & ~x755 & ~x758;
assign c971 =  x570 & ~x87 & ~x443 & ~x444 & ~x460 & ~x484;
assign c973 =  x302 & ~x408 & ~x740;
assign c975 = ~x19 & ~x29 & ~x54 & ~x56 & ~x57 & ~x81 & ~x110 & ~x138 & ~x140 & ~x165 & ~x489 & ~x519 & ~x573 & ~x574 & ~x575 & ~x603 & ~x629 & ~x657 & ~x658 & ~x715 & ~x741;
assign c977 =  x186 & ~x28 & ~x31 & ~x113 & ~x118 & ~x141 & ~x143 & ~x168 & ~x498 & ~x531 & ~x728;
assign c979 =  x262 &  x379 & ~x23 & ~x52 & ~x86 & ~x115 & ~x128 & ~x138 & ~x141 & ~x142 & ~x170 & ~x196 & ~x198 & ~x249 & ~x279 & ~x333 & ~x361 & ~x365 & ~x448 & ~x531 & ~x533 & ~x615 & ~x644 & ~x668 & ~x672 & ~x675 & ~x692 & ~x697 & ~x724 & ~x749 & ~x751;
assign c981 = ~x15 & ~x29 & ~x56 & ~x58 & ~x208 & ~x410 & ~x411 & ~x439 & ~x458 & ~x461 & ~x499 & ~x776;
assign c983 =  x231 & ~x0 & ~x26 & ~x382 & ~x724 & ~x729 & ~x730 & ~x746 & ~x747 & ~x757 & ~x758 & ~x774 & ~x776 & ~x777;
assign c985 =  x561;
assign c987 =  x238 &  x516 & ~x230;
assign c989 =  x130 & ~x52 & ~x442 & ~x471 & ~x472 & ~x486 & ~x499 & ~x525 & ~x751;
assign c991 =  x605 & ~x348 & ~x432;
assign c993 =  x233 &  x258 & ~x1 & ~x29 & ~x58 & ~x83 & ~x672 & ~x673 & ~x741 & ~x742 & ~x769;
assign c995 =  x549 & ~x24 & ~x27 & ~x56 & ~x58 & ~x168 & ~x224 & ~x449 & ~x476 & ~x531 & ~x554 & ~x583 & ~x584 & ~x586 & ~x587 & ~x608 & ~x609 & ~x610 & ~x611 & ~x612 & ~x613 & ~x615 & ~x638 & ~x639 & ~x640 & ~x641 & ~x643 & ~x644 & ~x665 & ~x666 & ~x667 & ~x669 & ~x671 & ~x672 & ~x673 & ~x692 & ~x696 & ~x698 & ~x701 & ~x719 & ~x721 & ~x725 & ~x726 & ~x731 & ~x747 & ~x748 & ~x749 & ~x750 & ~x751 & ~x758 & ~x763 & ~x776 & ~x777 & ~x778 & ~x783;
assign c997 =  x330 & ~x81 & ~x82 & ~x109 & ~x113 & ~x224 & ~x362 & ~x391 & ~x435 & ~x476 & ~x504 & ~x559 & ~x588 & ~x643 & ~x671;
assign c999 = ~x5 & ~x65 & ~x86 & ~x93 & ~x142 & ~x150 & ~x171 & ~x257 & ~x310 & ~x343 & ~x385 & ~x426 & ~x442 & ~x456 & ~x497 & ~x510 & ~x701;
assign c9101 = ~x1 & ~x5 & ~x32 & ~x46 & ~x49 & ~x50 & ~x61 & ~x75 & ~x76 & ~x81 & ~x82 & ~x107 & ~x111 & ~x115 & ~x118 & ~x131 & ~x133 & ~x135 & ~x146 & ~x171 & ~x198 & ~x229 & ~x247 & ~x280 & ~x284 & ~x307 & ~x311 & ~x312 & ~x338 & ~x339 & ~x359 & ~x388 & ~x396 & ~x417 & ~x448 & ~x450 & ~x478 & ~x528 & ~x601 & ~x602 & ~x605 & ~x615 & ~x617 & ~x629 & ~x631 & ~x645 & ~x658 & ~x660 & ~x667 & ~x698 & ~x731 & ~x757 & ~x758 & ~x779 & ~x782;
assign c9103 = ~x0 & ~x5 & ~x6 & ~x24 & ~x30 & ~x32 & ~x34 & ~x39 & ~x61 & ~x62 & ~x336 & ~x364 & ~x527 & ~x529 & ~x530 & ~x555 & ~x558 & ~x559 & ~x581 & ~x582 & ~x583 & ~x584 & ~x611 & ~x613 & ~x617 & ~x623 & ~x635 & ~x637 & ~x638 & ~x639 & ~x640 & ~x641 & ~x642 & ~x646 & ~x650 & ~x662 & ~x663 & ~x664 & ~x668 & ~x669 & ~x671 & ~x675 & ~x679 & ~x680 & ~x690 & ~x692 & ~x693 & ~x695 & ~x703 & ~x707 & ~x708 & ~x718 & ~x719 & ~x724 & ~x725 & ~x726 & ~x728 & ~x731 & ~x732 & ~x735 & ~x745 & ~x748 & ~x750 & ~x752 & ~x761 & ~x765 & ~x773 & ~x775 & ~x776 & ~x778 & ~x781 & ~x783;
assign c9105 =  x235 & ~x52 & ~x88 & ~x91 & ~x143 & ~x169 & ~x196 & ~x422 & ~x447 & ~x477 & ~x480 & ~x502 & ~x531 & ~x532 & ~x668 & ~x690 & ~x746 & ~x753 & ~x754 & ~x758 & ~x774 & ~x775 & ~x780;
assign c9107 = ~x1 & ~x23 & ~x79 & ~x80 & ~x82 & ~x85 & ~x108 & ~x138 & ~x141 & ~x142 & ~x169 & ~x252 & ~x455 & ~x483 & ~x558 & ~x614 & ~x641 & ~x642 & ~x644 & ~x646 & ~x668 & ~x669 & ~x696 & ~x702 & ~x716 & ~x729 & ~x731 & ~x743 & ~x752 & ~x756 & ~x758 & ~x782;
assign c9109 =  x449;
assign c9111 = ~x6 & ~x23 & ~x30 & ~x49 & ~x56 & ~x58 & ~x87 & ~x117 & ~x118 & ~x140 & ~x189 & ~x195 & ~x215 & ~x217 & ~x243 & ~x247 & ~x251 & ~x271 & ~x272 & ~x274 & ~x310 & ~x355 & ~x383 & ~x386 & ~x411 & ~x414 & ~x471 & ~x472 & ~x502 & ~x526 & ~x556 & ~x558 & ~x612 & ~x673 & ~x731;
assign c9113 =  x535 & ~x41 & ~x182 & ~x702;
assign c9115 = ~x2 & ~x5 & ~x6 & ~x15 & ~x17 & ~x19 & ~x20 & ~x23 & ~x25 & ~x27 & ~x28 & ~x30 & ~x31 & ~x34 & ~x48 & ~x49 & ~x50 & ~x51 & ~x52 & ~x53 & ~x54 & ~x55 & ~x56 & ~x57 & ~x77 & ~x81 & ~x82 & ~x85 & ~x88 & ~x100 & ~x103 & ~x105 & ~x107 & ~x111 & ~x136 & ~x137 & ~x141 & ~x142 & ~x143 & ~x144 & ~x161 & ~x164 & ~x166 & ~x167 & ~x170 & ~x190 & ~x192 & ~x195 & ~x217 & ~x218 & ~x219 & ~x222 & ~x226 & ~x246 & ~x248 & ~x252 & ~x253 & ~x275 & ~x279 & ~x280 & ~x281 & ~x305 & ~x306 & ~x310 & ~x334 & ~x335 & ~x337 & ~x361 & ~x362 & ~x365 & ~x367 & ~x388 & ~x390 & ~x391 & ~x393 & ~x394 & ~x417 & ~x420 & ~x444 & ~x447 & ~x448 & ~x474 & ~x476 & ~x502 & ~x504 & ~x533 & ~x560 & ~x584 & ~x644 & ~x671 & ~x699 & ~x720 & ~x721 & ~x727 & ~x756 & ~x758 & ~x767 & ~x779;
assign c9117 =  x360 & ~x717 & ~x718 & ~x746;
assign c9119 =  x397 & ~x0 & ~x20 & ~x49 & ~x51 & ~x52 & ~x141 & ~x322 & ~x323 & ~x698 & ~x735 & ~x751 & ~x753;
assign c9121 =  x126 &  x267 & ~x61 & ~x87 & ~x112 & ~x228 & ~x533 & ~x641 & ~x642;
assign c9123 =  x449;
assign c9125 = ~x18 & ~x22 & ~x23 & ~x31 & ~x52 & ~x81 & ~x110 & ~x113 & ~x134 & ~x136 & ~x167 & ~x196 & ~x491 & ~x503 & ~x519 & ~x575 & ~x602 & ~x630 & ~x659 & ~x709 & ~x755 & ~x769 & ~x783;
assign c9127 =  x602 & ~x0 & ~x23 & ~x25 & ~x27 & ~x83 & ~x85 & ~x86 & ~x111 & ~x112 & ~x113 & ~x195 & ~x252 & ~x393 & ~x469 & ~x497 & ~x502 & ~x531 & ~x557 & ~x560 & ~x581 & ~x582 & ~x583 & ~x608 & ~x636 & ~x639 & ~x645 & ~x646 & ~x664 & ~x665 & ~x720 & ~x724 & ~x730 & ~x731 & ~x748 & ~x751 & ~x758 & ~x776 & ~x783;
assign c9129 = ~x23 & ~x230 & ~x242 & ~x298 & ~x302 & ~x328 & ~x354 & ~x370 & ~x384 & ~x411 & ~x424 & ~x427 & ~x440 & ~x441 & ~x496 & ~x497 & ~x509 & ~x532 & ~x563 & ~x594;
assign c9131 =  x323 & ~x5 & ~x36 & ~x50 & ~x54 & ~x58 & ~x89 & ~x93 & ~x113 & ~x171 & ~x257 & ~x481 & ~x508 & ~x776;
assign c9133 = ~x33 & ~x87 & ~x89 & ~x139 & ~x520 & ~x530 & ~x577 & ~x684 & ~x712 & ~x731 & ~x756;
assign c9135 =  x205 &  x547 &  x603 & ~x196 & ~x308 & ~x335 & ~x748 & ~x750;
assign c9137 =  x633 & ~x0 & ~x27 & ~x53 & ~x56 & ~x57 & ~x83 & ~x85 & ~x113 & ~x196 & ~x224 & ~x253 & ~x307 & ~x335 & ~x362 & ~x363 & ~x364 & ~x390 & ~x418 & ~x497 & ~x498 & ~x499 & ~x501 & ~x502 & ~x503 & ~x530 & ~x532 & ~x544 & ~x553 & ~x558 & ~x559 & ~x561 & ~x626 & ~x754;
assign c9139 = ~x24 & ~x27 & ~x50 & ~x56 & ~x83 & ~x85 & ~x89 & ~x111 & ~x112 & ~x144 & ~x193 & ~x198 & ~x199 & ~x249 & ~x304 & ~x447 & ~x452 & ~x463 & ~x472 & ~x489 & ~x559 & ~x588 & ~x601;
assign c9141 =  x126 &  x154 &  x182 &  x266 &  x294 & ~x31 & ~x45 & ~x61 & ~x88 & ~x106 & ~x117 & ~x142 & ~x171 & ~x224 & ~x335 & ~x363 & ~x391 & ~x415 & ~x422 & ~x499 & ~x671 & ~x699 & ~x753;
assign c9143 = ~x1 & ~x14 & ~x26 & ~x29 & ~x30 & ~x32 & ~x57 & ~x58 & ~x83 & ~x86 & ~x111 & ~x114 & ~x115 & ~x140 & ~x141 & ~x142 & ~x167 & ~x196 & ~x553 & ~x555 & ~x584 & ~x598 & ~x608 & ~x609 & ~x614 & ~x615 & ~x616 & ~x625 & ~x637 & ~x641 & ~x643 & ~x645 & ~x646 & ~x668 & ~x674 & ~x690 & ~x695 & ~x696 & ~x698 & ~x700 & ~x703 & ~x708 & ~x718 & ~x724 & ~x726 & ~x731 & ~x735 & ~x748 & ~x752 & ~x761 & ~x775 & ~x781 & ~x783;
assign c9145 =  x714 & ~x29 & ~x47 & ~x60 & ~x87 & ~x114 & ~x115 & ~x117 & ~x118 & ~x132 & ~x145 & ~x146 & ~x199 & ~x200 & ~x201 & ~x219 & ~x220 & ~x243 & ~x250 & ~x256 & ~x275 & ~x277 & ~x283 & ~x302 & ~x303 & ~x304 & ~x305 & ~x330 & ~x331 & ~x357 & ~x385 & ~x397 & ~x413 & ~x414 & ~x425 & ~x442 & ~x453 & ~x480 & ~x507 & ~x509 & ~x527 & ~x668;
assign c9147 =  x298 &  x444;
assign c9149 =  x589 &  x677;
assign c9151 = ~x1 & ~x4 & ~x5 & ~x16 & ~x23 & ~x26 & ~x27 & ~x29 & ~x31 & ~x34 & ~x51 & ~x56 & ~x59 & ~x62 & ~x63 & ~x75 & ~x78 & ~x79 & ~x80 & ~x81 & ~x83 & ~x84 & ~x87 & ~x91 & ~x115 & ~x118 & ~x119 & ~x133 & ~x134 & ~x136 & ~x140 & ~x161 & ~x163 & ~x166 & ~x167 & ~x193 & ~x196 & ~x197 & ~x199 & ~x201 & ~x220 & ~x223 & ~x226 & ~x245 & ~x249 & ~x250 & ~x251 & ~x272 & ~x273 & ~x274 & ~x275 & ~x281 & ~x304 & ~x305 & ~x306 & ~x310 & ~x311 & ~x312 & ~x330 & ~x331 & ~x332 & ~x333 & ~x359 & ~x362 & ~x367 & ~x387 & ~x388 & ~x415 & ~x416 & ~x417 & ~x420 & ~x423 & ~x442 & ~x444 & ~x445 & ~x446 & ~x448 & ~x449 & ~x471 & ~x473 & ~x475 & ~x499 & ~x503 & ~x506 & ~x509 & ~x534 & ~x537 & ~x556 & ~x560 & ~x561 & ~x563 & ~x565 & ~x584 & ~x591 & ~x612 & ~x617 & ~x622 & ~x640 & ~x645 & ~x646 & ~x662 & ~x665 & ~x667 & ~x669 & ~x673 & ~x675 & ~x676 & ~x678 & ~x692 & ~x704 & ~x705 & ~x706 & ~x723 & ~x726 & ~x730 & ~x734 & ~x751 & ~x752 & ~x753 & ~x755 & ~x760 & ~x761 & ~x778 & ~x779;
assign c9153 =  x747 & ~x53 & ~x108 & ~x222 & ~x252 & ~x255 & ~x304 & ~x333 & ~x359 & ~x415 & ~x418 & ~x493;
assign c9155 =  x314 &  x317 &  x341 & ~x78 & ~x783;
assign c9157 =  x277 &  x360;
assign c9159 = ~x81 & ~x82 & ~x86 & ~x109 & ~x112 & ~x135 & ~x197 & ~x252 & ~x323 & ~x448 & ~x689 & ~x717 & ~x718 & ~x742 & ~x745 & ~x769;
assign c9161 = ~x1 & ~x16 & ~x17 & ~x20 & ~x24 & ~x26 & ~x29 & ~x50 & ~x51 & ~x54 & ~x57 & ~x78 & ~x81 & ~x82 & ~x83 & ~x107 & ~x108 & ~x109 & ~x110 & ~x112 & ~x114 & ~x137 & ~x138 & ~x139 & ~x141 & ~x164 & ~x165 & ~x166 & ~x191 & ~x192 & ~x193 & ~x196 & ~x220 & ~x221 & ~x223 & ~x224 & ~x248 & ~x249 & ~x250 & ~x251 & ~x277 & ~x280 & ~x305 & ~x364 & ~x438 & ~x743 & ~x744 & ~x745 & ~x771 & ~x783;
assign c9163 = ~x1 & ~x2 & ~x4 & ~x24 & ~x51 & ~x54 & ~x57 & ~x58 & ~x82 & ~x83 & ~x114 & ~x141 & ~x168 & ~x170 & ~x182 & ~x197 & ~x198 & ~x208 & ~x249 & ~x307 & ~x345 & ~x433 & ~x448 & ~x715;
assign c9165 =  x541 &  x542 & ~x117 & ~x230 & ~x651;
assign c9167 = ~x3 & ~x4 & ~x22 & ~x24 & ~x25 & ~x27 & ~x31 & ~x32 & ~x78 & ~x79 & ~x81 & ~x112 & ~x139 & ~x167 & ~x448 & ~x552 & ~x559 & ~x581 & ~x582 & ~x606 & ~x608 & ~x609 & ~x610 & ~x611 & ~x637 & ~x641 & ~x643 & ~x645 & ~x651 & ~x662 & ~x666 & ~x673 & ~x690 & ~x701 & ~x704 & ~x706 & ~x708 & ~x718 & ~x720 & ~x725 & ~x730 & ~x732 & ~x734 & ~x746 & ~x747 & ~x748 & ~x754 & ~x756 & ~x759 & ~x772 & ~x775;
assign c9169 = ~x3 & ~x19 & ~x23 & ~x25 & ~x29 & ~x57 & ~x82 & ~x85 & ~x86 & ~x196 & ~x350 & ~x351 & ~x365 & ~x390 & ~x405 & ~x421 & ~x505 & ~x557 & ~x679 & ~x680 & ~x681 & ~x708 & ~x709 & ~x736 & ~x737 & ~x763 & ~x765;
assign c9171 =  x322 &  x349 & ~x86 & ~x87 & ~x106 & ~x118 & ~x119 & ~x131 & ~x162 & ~x171 & ~x174 & ~x225 & ~x228;
assign c9173 =  x211 & ~x1 & ~x20 & ~x53 & ~x56 & ~x80 & ~x81 & ~x103 & ~x104 & ~x110 & ~x131 & ~x134 & ~x137 & ~x141 & ~x144 & ~x161 & ~x165 & ~x189 & ~x192 & ~x195 & ~x198 & ~x199 & ~x200 & ~x229 & ~x255 & ~x420 & ~x529 & ~x727 & ~x757 & ~x782;
assign c9175 =  x556;
assign c9177 =  x456 & ~x171 & ~x244 & ~x360 & ~x444 & ~x537 & ~x546 & ~x549 & ~x697 & ~x781;
assign c9179 =  x288 &  x456 &  x457 & ~x735;
assign c9181 =  x181 &  x435 & ~x145 & ~x189 & ~x227 & ~x301 & ~x330 & ~x387;
assign c9183 =  x306 & ~x582 & ~x692 & ~x718 & ~x723;
assign c9185 =  x473;
assign c9187 =  x314 & ~x24 & ~x25 & ~x31 & ~x41 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x59 & ~x83 & ~x88 & ~x111 & ~x127 & ~x130 & ~x154 & ~x280 & ~x524 & ~x525 & ~x552 & ~x553 & ~x768 & ~x781;
assign c9189 =  x71 & ~x468 & ~x527 & ~x611 & ~x654;
assign c9191 =  x606 & ~x23 & ~x57 & ~x140 & ~x170 & ~x220 & ~x221 & ~x224 & ~x226 & ~x250 & ~x252 & ~x253 & ~x280 & ~x307 & ~x308 & ~x334 & ~x335 & ~x390 & ~x476 & ~x506 & ~x560 & ~x727 & ~x754 & ~x777 & ~x781 & ~x782;
assign c9193 =  x524 & ~x240 & ~x431;
assign c9195 =  x379 & ~x245 & ~x302 & ~x330 & ~x384 & ~x413 & ~x468 & ~x493 & ~x496 & ~x552 & ~x582 & ~x607 & ~x676;
assign c9197 =  x546 & ~x39 & ~x55 & ~x83 & ~x252 & ~x555 & ~x634 & ~x665 & ~x720 & ~x742 & ~x753;
assign c9199 = ~x110 & ~x137 & ~x138 & ~x165 & ~x170 & ~x195 & ~x222 & ~x249 & ~x250 & ~x251 & ~x696 & ~x697 & ~x726 & ~x727;
assign c9201 =  x249 & ~x301 & ~x638 & ~x720 & ~x748 & ~x749;
assign c9203 =  x528 & ~x78 & ~x81;
assign c9205 =  x557 & ~x357;
assign c9207 =  x287 &  x399 &  x427 & ~x650 & ~x725;
assign c9209 = ~x3 & ~x24 & ~x83 & ~x84 & ~x112 & ~x167 & ~x195 & ~x252 & ~x267 & ~x305 & ~x307 & ~x322 & ~x359 & ~x364 & ~x375 & ~x377 & ~x388 & ~x389 & ~x391 & ~x414 & ~x448 & ~x472 & ~x588 & ~x643 & ~x729 & ~x754;
assign c9211 =  x292 &  x488 & ~x89 & ~x136 & ~x146 & ~x175 & ~x177 & ~x646;
assign c9213 =  x429 & ~x19 & ~x88 & ~x138 & ~x168 & ~x194 & ~x494 & ~x496 & ~x653 & ~x709;
assign c9215 = ~x0 & ~x31 & ~x53 & ~x57 & ~x58 & ~x59 & ~x112 & ~x113 & ~x141 & ~x168 & ~x224 & ~x437 & ~x465 & ~x485 & ~x486 & ~x501 & ~x531 & ~x541 & ~x556 & ~x558 & ~x730 & ~x745 & ~x757;
assign c9217 = ~x0 & ~x2 & ~x3 & ~x7 & ~x8 & ~x23 & ~x26 & ~x28 & ~x29 & ~x31 & ~x51 & ~x54 & ~x56 & ~x58 & ~x59 & ~x60 & ~x84 & ~x85 & ~x110 & ~x114 & ~x390 & ~x419 & ~x420 & ~x445 & ~x447 & ~x471 & ~x472 & ~x475 & ~x498 & ~x499 & ~x500 & ~x503 & ~x504 & ~x526 & ~x529 & ~x530 & ~x531 & ~x553 & ~x557 & ~x558 & ~x568 & ~x569 & ~x582 & ~x583 & ~x584 & ~x587 & ~x595 & ~x609 & ~x610 & ~x612 & ~x613 & ~x614 & ~x615 & ~x616 & ~x617 & ~x623 & ~x635 & ~x636 & ~x639 & ~x640 & ~x641 & ~x644 & ~x645 & ~x646 & ~x649 & ~x650 & ~x664 & ~x665 & ~x666 & ~x672 & ~x673 & ~x674 & ~x675 & ~x676 & ~x677 & ~x678 & ~x691 & ~x692 & ~x693 & ~x694 & ~x695 & ~x696 & ~x698 & ~x699 & ~x700 & ~x703 & ~x719 & ~x721 & ~x722 & ~x723 & ~x724 & ~x726 & ~x727 & ~x728 & ~x729 & ~x731 & ~x732 & ~x733 & ~x734 & ~x746 & ~x747 & ~x748 & ~x751 & ~x752 & ~x753 & ~x754 & ~x757 & ~x758 & ~x759 & ~x763 & ~x776 & ~x777 & ~x778 & ~x780 & ~x781 & ~x782 & ~x783;
assign c9219 = ~x1 & ~x3 & ~x5 & ~x17 & ~x18 & ~x23 & ~x27 & ~x31 & ~x57 & ~x58 & ~x59 & ~x86 & ~x87 & ~x100 & ~x111 & ~x113 & ~x114 & ~x196 & ~x364 & ~x475 & ~x529 & ~x531 & ~x552 & ~x556 & ~x557 & ~x580 & ~x581 & ~x582 & ~x583 & ~x588 & ~x609 & ~x611 & ~x613 & ~x635 & ~x636 & ~x638 & ~x639 & ~x642 & ~x643 & ~x645 & ~x646 & ~x650 & ~x662 & ~x664 & ~x666 & ~x667 & ~x670 & ~x671 & ~x674 & ~x676 & ~x678 & ~x679 & ~x691 & ~x692 & ~x695 & ~x696 & ~x700 & ~x701 & ~x705 & ~x706 & ~x721 & ~x722 & ~x725 & ~x726 & ~x727 & ~x730 & ~x732 & ~x734 & ~x744 & ~x747 & ~x748 & ~x749 & ~x750 & ~x753 & ~x758 & ~x759 & ~x774 & ~x775 & ~x777 & ~x778 & ~x779 & ~x780 & ~x782;
assign c9221 = ~x6 & ~x19 & ~x59 & ~x63 & ~x82 & ~x86 & ~x135 & ~x148 & ~x164 & ~x169 & ~x176 & ~x191 & ~x199 & ~x201 & ~x204 & ~x205 & ~x219 & ~x226 & ~x228 & ~x252 & ~x255 & ~x283 & ~x338 & ~x446 & ~x561 & ~x562 & ~x603 & ~x730 & ~x756;
assign c9223 = ~x0 & ~x22 & ~x23 & ~x29 & ~x81 & ~x138 & ~x195 & ~x252 & ~x281 & ~x385 & ~x412 & ~x467 & ~x468 & ~x505 & ~x720 & ~x721 & ~x751 & ~x779;
assign c9225 = ~x37 & ~x269 & ~x380 & ~x381 & ~x409 & ~x528 & ~x742;
assign c9227 =  x93 &  x289 & ~x24 & ~x85 & ~x196 & ~x477 & ~x749;
assign c9229 =  x547 & ~x0 & ~x25 & ~x28 & ~x58 & ~x586 & ~x634 & ~x645 & ~x670 & ~x676 & ~x677 & ~x699 & ~x700 & ~x703 & ~x705 & ~x723 & ~x724 & ~x731 & ~x732 & ~x733 & ~x742 & ~x752 & ~x753 & ~x756 & ~x779 & ~x781 & ~x782;
assign c9231 =  x158 & ~x30 & ~x391 & ~x561 & ~x672 & ~x750 & ~x759;
assign c9233 = ~x1 & ~x51 & ~x81 & ~x83 & ~x110 & ~x112 & ~x137 & ~x138 & ~x139 & ~x167 & ~x278 & ~x349 & ~x417 & ~x445 & ~x448 & ~x450 & ~x475 & ~x516 & ~x542 & ~x644 & ~x697 & ~x755 & ~x782;
assign c9235 = ~x51 & ~x53 & ~x324 & ~x351 & ~x406 & ~x432 & ~x710 & ~x737 & ~x755 & ~x764;
assign c9237 = ~x3 & ~x50 & ~x51 & ~x78 & ~x109 & ~x114 & ~x138 & ~x145 & ~x149 & ~x172 & ~x200 & ~x327 & ~x414 & ~x522 & ~x652;
assign c9239 = ~x87 & ~x111 & ~x114 & ~x118 & ~x138 & ~x179 & ~x228 & ~x287 & ~x426 & ~x454 & ~x482 & ~x661;
assign c9241 = ~x12 & ~x29 & ~x168 & ~x320 & ~x321 & ~x347 & ~x349 & ~x374 & ~x375 & ~x377 & ~x474 & ~x542 & ~x571 & ~x726;
assign c9243 = ~x19 & ~x49 & ~x77 & ~x78 & ~x81 & ~x113 & ~x170 & ~x173 & ~x193 & ~x605 & ~x644 & ~x687 & ~x715 & ~x744 & ~x750 & ~x770;
assign c9245 =  x151 &  x152 &  x715 &  x743 & ~x278 & ~x331 & ~x358 & ~x387 & ~x471 & ~x680;
assign c9247 =  x237 &  x571 & ~x117 & ~x173 & ~x201 & ~x229 & ~x301;
assign c9249 = ~x25 & ~x26 & ~x29 & ~x30 & ~x55 & ~x110 & ~x195 & ~x348 & ~x418 & ~x463 & ~x474 & ~x502 & ~x571 & ~x574 & ~x575 & ~x599 & ~x603 & ~x656 & ~x727 & ~x782;
assign c9251 =  x633 & ~x141 & ~x252 & ~x505 & ~x555 & ~x618 & ~x637 & ~x641 & ~x749 & ~x759;
assign c9253 =  x473;
assign c9255 =  x237 &  x543 &  x569;
assign c9257 = ~x1 & ~x2 & ~x24 & ~x27 & ~x30 & ~x56 & ~x58 & ~x61 & ~x82 & ~x85 & ~x86 & ~x110 & ~x111 & ~x114 & ~x138 & ~x140 & ~x167 & ~x168 & ~x222 & ~x224 & ~x336 & ~x353 & ~x382 & ~x409 & ~x410 & ~x438 & ~x474 & ~x476 & ~x493 & ~x521 & ~x755 & ~x757;
assign c9259 = ~x0 & ~x1 & ~x29 & ~x58 & ~x141 & ~x378 & ~x379 & ~x405 & ~x407 & ~x547 & ~x574 & ~x575 & ~x644 & ~x768;
assign c9261 = ~x30 & ~x51 & ~x57 & ~x80 & ~x81 & ~x82 & ~x106 & ~x112 & ~x114 & ~x136 & ~x141 & ~x162 & ~x193 & ~x195 & ~x223 & ~x308 & ~x378 & ~x379 & ~x415 & ~x416 & ~x671 & ~x710 & ~x740;
assign c9263 =  x353 &  x521 & ~x406 & ~x730;
assign c9265 = ~x32 & ~x114 & ~x115 & ~x147 & ~x148 & ~x170 & ~x176 & ~x198 & ~x200 & ~x201 & ~x204 & ~x225 & ~x227 & ~x229 & ~x231 & ~x233 & ~x256 & ~x257 & ~x258 & ~x260 & ~x760;
assign c9267 =  x348 & ~x90 & ~x165 & ~x234 & ~x303 & ~x593;
assign c9269 =  x656 & ~x358 & ~x375 & ~x376 & ~x415 & ~x441 & ~x442 & ~x587;
assign c9271 = ~x3 & ~x27 & ~x30 & ~x83 & ~x140 & ~x296 & ~x351 & ~x444 & ~x462 & ~x471 & ~x498 & ~x499 & ~x527 & ~x769;
assign c9273 =  x236 &  x515 & ~x3 & ~x60 & ~x112 & ~x115 & ~x131 & ~x132 & ~x141 & ~x199 & ~x652 & ~x680;
assign c9275 =  x596 &  x598 & ~x276 & ~x332 & ~x364 & ~x444;
assign c9277 = ~x29 & ~x53 & ~x54 & ~x58 & ~x110 & ~x111 & ~x138 & ~x170 & ~x249 & ~x278 & ~x305 & ~x459 & ~x460 & ~x461 & ~x462 & ~x469 & ~x500 & ~x746 & ~x748 & ~x753 & ~x758 & ~x777;
assign c9279 = ~x1 & ~x58 & ~x148 & ~x231 & ~x232 & ~x288 & ~x328 & ~x442 & ~x590 & ~x662 & ~x680 & ~x721;
assign c9281 =  x324 & ~x5 & ~x26 & ~x49 & ~x87 & ~x88 & ~x115 & ~x170 & ~x526 & ~x582 & ~x584 & ~x587 & ~x609 & ~x613 & ~x614 & ~x636 & ~x637 & ~x640 & ~x642 & ~x643 & ~x647 & ~x663 & ~x665 & ~x675 & ~x690 & ~x691 & ~x719 & ~x730 & ~x757 & ~x760 & ~x776 & ~x778 & ~x780;
assign c9283 =  x247 & ~x28 & ~x433 & ~x755;
assign c9285 =  x125 &  x293 &  x543 & ~x90 & ~x145 & ~x201;
assign c9287 =  x159 & ~x23 & ~x294;
assign c9289 =  x743 & ~x147 & ~x272 & ~x287 & ~x311 & ~x383 & ~x427 & ~x441 & ~x450 & ~x479 & ~x482 & ~x497;
assign c9291 = ~x2 & ~x16 & ~x29 & ~x41 & ~x85 & ~x111 & ~x182 & ~x195 & ~x196 & ~x209 & ~x308 & ~x310 & ~x387 & ~x406 & ~x653 & ~x779;
assign c9293 = ~x1 & ~x56 & ~x168 & ~x296 & ~x323 & ~x394 & ~x406 & ~x416 & ~x417 & ~x421 & ~x433 & ~x434 & ~x444 & ~x461 & ~x653 & ~x680 & ~x681;
assign c9295 = ~x114 & ~x427 & ~x559 & ~x671 & ~x692 & ~x700 & ~x716 & ~x755 & ~x756 & ~x773;
assign c9297 =  x214 &  x388;
assign c9299 = ~x1 & ~x2 & ~x26 & ~x27 & ~x28 & ~x31 & ~x81 & ~x82 & ~x110 & ~x111 & ~x113 & ~x136 & ~x139 & ~x164 & ~x166 & ~x192 & ~x221 & ~x224 & ~x249 & ~x251 & ~x253 & ~x307 & ~x361 & ~x362 & ~x391 & ~x445 & ~x446 & ~x447 & ~x448 & ~x474 & ~x476 & ~x504 & ~x518 & ~x529 & ~x544 & ~x545 & ~x547 & ~x558 & ~x560 & ~x573 & ~x574 & ~x601 & ~x602 & ~x603 & ~x615 & ~x660 & ~x672 & ~x726 & ~x753 & ~x755;
assign c9301 =  x444 & ~x766;
assign c9303 = ~x2 & ~x5 & ~x54 & ~x78 & ~x82 & ~x85 & ~x90 & ~x108 & ~x114 & ~x115 & ~x136 & ~x145 & ~x193 & ~x198 & ~x220 & ~x281 & ~x448 & ~x449 & ~x506 & ~x545 & ~x546 & ~x547 & ~x572 & ~x575 & ~x601 & ~x603 & ~x728 & ~x755;
assign c9305 = ~x42 & ~x209 & ~x405 & ~x406 & ~x415 & ~x517 & ~x542 & ~x544;
assign c9307 =  x260 &  x288 &  x344 & ~x85 & ~x114 & ~x196 & ~x437;
assign c9309 = ~x2 & ~x28 & ~x32 & ~x55 & ~x87 & ~x170 & ~x251 & ~x338 & ~x364 & ~x418 & ~x434 & ~x435 & ~x442 & ~x444 & ~x461 & ~x474 & ~x601 & ~x628 & ~x629 & ~x672 & ~x699 & ~x750;
assign c9311 = ~x3 & ~x29 & ~x32 & ~x54 & ~x84 & ~x110 & ~x112 & ~x166 & ~x298 & ~x354 & ~x383 & ~x410 & ~x438 & ~x466 & ~x493 & ~x494 & ~x504 & ~x523 & ~x532 & ~x550 & ~x578 & ~x615 & ~x728 & ~x763;
assign c9313 =  x244 & ~x13 & ~x41 & ~x349 & ~x405 & ~x507;
assign c9315 = ~x33 & ~x53 & ~x192 & ~x216 & ~x218 & ~x257 & ~x299 & ~x327 & ~x360 & ~x385 & ~x441 & ~x453 & ~x481 & ~x503 & ~x549 & ~x661 & ~x762;
assign c9317 =  x241 & ~x23 & ~x56 & ~x137 & ~x139 & ~x197 & ~x426 & ~x428 & ~x444 & ~x471 & ~x482;
assign c9319 = ~x87 & ~x91 & ~x205 & ~x231 & ~x256 & ~x315 & ~x645 & ~x661 & ~x673 & ~x718;
assign c9321 =  x406 &  x407 &  x431 & ~x62 & ~x171 & ~x217 & ~x596;
assign c9323 =  x603 &  x681 & ~x748;
assign c9325 =  x444 & ~x467;
assign c9327 =  x524 & ~x0 & ~x23 & ~x30 & ~x55 & ~x111 & ~x168 & ~x336 & ~x447 & ~x501 & ~x502 & ~x504 & ~x531 & ~x556 & ~x557 & ~x583 & ~x584 & ~x588 & ~x610 & ~x612 & ~x614 & ~x615 & ~x638 & ~x639 & ~x642 & ~x644 & ~x670 & ~x693 & ~x697 & ~x699 & ~x701 & ~x729 & ~x749 & ~x750 & ~x759 & ~x762 & ~x777 & ~x780;
assign c9329 =  x665 & ~x79 & ~x198 & ~x220 & ~x278 & ~x335;
assign c9331 =  x513 &  x514 &  x515 & ~x4 & ~x59 & ~x75 & ~x88 & ~x143 & ~x145 & ~x161 & ~x174 & ~x198 & ~x199 & ~x200 & ~x274 & ~x303 & ~x332;
assign c9333 =  x343 &  x371 &  x455 & ~x85 & ~x611 & ~x612 & ~x636 & ~x638 & ~x668 & ~x672 & ~x692 & ~x694 & ~x696 & ~x727 & ~x735;
assign c9335 = ~x39 & ~x54 & ~x58 & ~x382 & ~x384 & ~x608 & ~x661 & ~x741 & ~x783;
assign c9337 =  x577 & ~x83 & ~x363 & ~x418 & ~x421 & ~x500 & ~x505 & ~x526 & ~x527 & ~x541 & ~x696 & ~x699 & ~x725 & ~x726 & ~x748 & ~x752 & ~x756;
assign c9339 =  x541 &  x542 & ~x2 & ~x19 & ~x24 & ~x49 & ~x56 & ~x59 & ~x77 & ~x87 & ~x113 & ~x114 & ~x117 & ~x118 & ~x141 & ~x142 & ~x144 & ~x145 & ~x167 & ~x168 & ~x169 & ~x170 & ~x172 & ~x191 & ~x192 & ~x195 & ~x200 & ~x201 & ~x253 & ~x255 & ~x280 & ~x332 & ~x335 & ~x336 & ~x388 & ~x392 & ~x446 & ~x473 & ~x475 & ~x476 & ~x557 & ~x601 & ~x729;
assign c9341 =  x444 & ~x169 & ~x587;
assign c9343 =  x100 &  x212 &  x268 & ~x25 & ~x426;
assign c9345 = ~x30 & ~x52 & ~x81 & ~x109 & ~x113 & ~x320 & ~x327 & ~x355 & ~x356 & ~x383 & ~x411 & ~x416 & ~x494;
assign c9347 = ~x23 & ~x63 & ~x64 & ~x87 & ~x119 & ~x121 & ~x139 & ~x140 & ~x143 & ~x145 & ~x161 & ~x175 & ~x192 & ~x201 & ~x202 & ~x252 & ~x255 & ~x257 & ~x258 & ~x259 & ~x274 & ~x283 & ~x304 & ~x340 & ~x391 & ~x395 & ~x397 & ~x424 & ~x425 & ~x452 & ~x455 & ~x479 & ~x480 & ~x499 & ~x506 & ~x535 & ~x557 & ~x560 & ~x561 & ~x611 & ~x643 & ~x673 & ~x703 & ~x728 & ~x732 & ~x751 & ~x757 & ~x780 & ~x783;
assign c9349 =  x189 & ~x25 & ~x26 & ~x31 & ~x296;
assign c9351 =  x634 & ~x4 & ~x30 & ~x53 & ~x80 & ~x81 & ~x135 & ~x195 & ~x222 & ~x225 & ~x226 & ~x248 & ~x249 & ~x250 & ~x253 & ~x306 & ~x307 & ~x308 & ~x333 & ~x336 & ~x361 & ~x363 & ~x389 & ~x392 & ~x393 & ~x532 & ~x557 & ~x588;
assign c9353 = ~x27 & ~x85 & ~x86 & ~x410 & ~x466 & ~x541 & ~x607 & ~x642 & ~x645 & ~x742 & ~x782;
assign c9355 = ~x26 & ~x34 & ~x85 & ~x92 & ~x118 & ~x120 & ~x159 & ~x171 & ~x177 & ~x201 & ~x226 & ~x311 & ~x468 & ~x529 & ~x537 & ~x568 & ~x661;
assign c9357 = ~x3 & ~x6 & ~x8 & ~x36 & ~x53 & ~x55 & ~x58 & ~x60 & ~x77 & ~x78 & ~x80 & ~x84 & ~x87 & ~x88 & ~x92 & ~x103 & ~x111 & ~x112 & ~x113 & ~x131 & ~x132 & ~x133 & ~x138 & ~x140 & ~x141 & ~x159 & ~x162 & ~x165 & ~x168 & ~x170 & ~x173 & ~x201 & ~x218 & ~x220 & ~x225 & ~x227 & ~x229 & ~x230 & ~x251 & ~x254 & ~x259 & ~x280 & ~x311 & ~x337 & ~x342 & ~x357 & ~x360 & ~x385 & ~x394 & ~x471 & ~x474 & ~x476 & ~x499 & ~x503 & ~x508 & ~x529 & ~x532 & ~x533 & ~x534 & ~x555 & ~x562 & ~x584 & ~x590 & ~x611 & ~x618 & ~x639 & ~x643 & ~x666 & ~x668 & ~x669 & ~x670 & ~x671 & ~x701 & ~x702 & ~x724 & ~x725 & ~x730 & ~x753 & ~x755 & ~x780 & ~x781;
assign c9359 =  x621 & ~x21 & ~x22 & ~x24 & ~x25 & ~x27 & ~x51 & ~x52 & ~x55 & ~x57 & ~x78 & ~x79 & ~x80 & ~x82 & ~x83 & ~x84 & ~x106 & ~x107 & ~x108 & ~x109 & ~x113 & ~x134 & ~x135 & ~x136 & ~x137 & ~x138 & ~x140 & ~x164 & ~x165 & ~x166 & ~x167 & ~x191 & ~x193 & ~x195 & ~x220 & ~x221 & ~x222 & ~x248 & ~x250 & ~x275 & ~x277 & ~x278 & ~x279 & ~x305 & ~x306 & ~x335 & ~x363 & ~x417 & ~x474 & ~x475 & ~x531 & ~x532 & ~x756 & ~x779 & ~x781 & ~x782;
assign c9361 =  x127 &  x155 &  x239 &  x378 & ~x78 & ~x106 & ~x199;
assign c9363 =  x315 &  x371 &  x400 & ~x28 & ~x30 & ~x140 & ~x252 & ~x498 & ~x524 & ~x526 & ~x553 & ~x671 & ~x779;
assign c9365 =  x317 &  x512 & ~x89 & ~x199;
assign c9367 =  x502;
assign c9369 =  x620 & ~x22 & ~x114 & ~x165 & ~x248 & ~x436;
assign c9371 =  x607 &  x608;
assign c9373 =  x324 & ~x0 & ~x3 & ~x31 & ~x32 & ~x57 & ~x59 & ~x62 & ~x88 & ~x115 & ~x116 & ~x166 & ~x169 & ~x196 & ~x222 & ~x226 & ~x245 & ~x247 & ~x304 & ~x305 & ~x365 & ~x419 & ~x425 & ~x445 & ~x447 & ~x474 & ~x506 & ~x509 & ~x510 & ~x618 & ~x700 & ~x701;
assign c9375 =  x610 & ~x27 & ~x52 & ~x137 & ~x138 & ~x139 & ~x140 & ~x165 & ~x170 & ~x194 & ~x220 & ~x277 & ~x753;
assign c9377 =  x92 &  x287 & ~x55 & ~x696 & ~x721 & ~x724 & ~x750 & ~x751 & ~x757 & ~x775;
assign c9379 =  x555 & ~x51 & ~x82 & ~x136 & ~x192 & ~x277 & ~x335 & ~x670;
assign c9381 =  x178 &  x205 &  x549 & ~x505 & ~x669;
assign c9383 = ~x1 & ~x2 & ~x4 & ~x24 & ~x26 & ~x27 & ~x29 & ~x30 & ~x32 & ~x52 & ~x53 & ~x56 & ~x58 & ~x63 & ~x82 & ~x83 & ~x86 & ~x113 & ~x114 & ~x252 & ~x308 & ~x314 & ~x336 & ~x418 & ~x419 & ~x423 & ~x444 & ~x446 & ~x447 & ~x448 & ~x451 & ~x452 & ~x473 & ~x476 & ~x477 & ~x479 & ~x499 & ~x500 & ~x501 & ~x502 & ~x505 & ~x506 & ~x508 & ~x525 & ~x529 & ~x530 & ~x531 & ~x532 & ~x533 & ~x534 & ~x535 & ~x556 & ~x557 & ~x558 & ~x563 & ~x569 & ~x582 & ~x583 & ~x584 & ~x586 & ~x587 & ~x588 & ~x589 & ~x591 & ~x595 & ~x611 & ~x615 & ~x616 & ~x618 & ~x620 & ~x637 & ~x638 & ~x639 & ~x640 & ~x643 & ~x645 & ~x647 & ~x651 & ~x667 & ~x669 & ~x670 & ~x672 & ~x673 & ~x674 & ~x676 & ~x679 & ~x692 & ~x693 & ~x696 & ~x698 & ~x701 & ~x702 & ~x703 & ~x707 & ~x708 & ~x709 & ~x720 & ~x721 & ~x722 & ~x723 & ~x725 & ~x731 & ~x732 & ~x736 & ~x748 & ~x749 & ~x750 & ~x755 & ~x757 & ~x761 & ~x762 & ~x778 & ~x783;
assign c9385 =  x526 & ~x24 & ~x52 & ~x56 & ~x85 & ~x138 & ~x222 & ~x252 & ~x640 & ~x643 & ~x669 & ~x698 & ~x724 & ~x727 & ~x775 & ~x780;
assign c9387 =  x298 & ~x23 & ~x27 & ~x28 & ~x50 & ~x53 & ~x54 & ~x56 & ~x81 & ~x82 & ~x108 & ~x110 & ~x112 & ~x114 & ~x137 & ~x141 & ~x163 & ~x165 & ~x167 & ~x170 & ~x193 & ~x196 & ~x221 & ~x223 & ~x249 & ~x276 & ~x305 & ~x308 & ~x333 & ~x334 & ~x335 & ~x336 & ~x390 & ~x391 & ~x433 & ~x447;
assign c9389 = ~x23 & ~x25 & ~x27 & ~x52 & ~x56 & ~x126 & ~x139 & ~x140 & ~x221 & ~x462 & ~x475 & ~x490 & ~x545 & ~x574 & ~x575 & ~x603 & ~x631 & ~x657 & ~x687 & ~x688 & ~x768;
assign c9391 = ~x30 & ~x51 & ~x53 & ~x85 & ~x92 & ~x122 & ~x135 & ~x145 & ~x191 & ~x200 & ~x221 & ~x223 & ~x249 & ~x308 & ~x331 & ~x335 & ~x500 & ~x519 & ~x534 & ~x558 & ~x759;
assign c9393 =  x187;
assign c9395 =  x361 & ~x721 & ~x765;
assign c9397 =  x212 & ~x3 & ~x49 & ~x77 & ~x81 & ~x166 & ~x469 & ~x497 & ~x559 & ~x627 & ~x653;
assign c9399 =  x530;
assign c9401 =  x210 & ~x23 & ~x85 & ~x86 & ~x113 & ~x116 & ~x387 & ~x397 & ~x398 & ~x415 & ~x421 & ~x442 & ~x473 & ~x482 & ~x500 & ~x507 & ~x531 & ~x534 & ~x617 & ~x699 & ~x759 & ~x781;
assign c9403 =  x269 & ~x3 & ~x21 & ~x27 & ~x30 & ~x32 & ~x34 & ~x51 & ~x54 & ~x56 & ~x58 & ~x80 & ~x86 & ~x108 & ~x109 & ~x110 & ~x112 & ~x134 & ~x135 & ~x138 & ~x140 & ~x142 & ~x143 & ~x162 & ~x165 & ~x169 & ~x190 & ~x191 & ~x192 & ~x196 & ~x247 & ~x276 & ~x310 & ~x391 & ~x418 & ~x445 & ~x701 & ~x726 & ~x728 & ~x729 & ~x752;
assign c9405 =  x182 & ~x31 & ~x232 & ~x252 & ~x261 & ~x285 & ~x308 & ~x451 & ~x480 & ~x535;
assign c9407 =  x325 & ~x24 & ~x28 & ~x57 & ~x82 & ~x87 & ~x114 & ~x141 & ~x168 & ~x250 & ~x252 & ~x279 & ~x342 & ~x370 & ~x454 & ~x482 & ~x484 & ~x505 & ~x537 & ~x561 & ~x586 & ~x644 & ~x670 & ~x701;
assign c9409 =  x550 &  x713 & ~x196 & ~x489;
assign c9411 = ~x0 & ~x1 & ~x2 & ~x3 & ~x4 & ~x5 & ~x6 & ~x15 & ~x16 & ~x17 & ~x19 & ~x20 & ~x21 & ~x22 & ~x23 & ~x24 & ~x25 & ~x26 & ~x27 & ~x28 & ~x29 & ~x30 & ~x31 & ~x32 & ~x33 & ~x34 & ~x42 & ~x45 & ~x48 & ~x49 & ~x50 & ~x51 & ~x52 & ~x53 & ~x54 & ~x55 & ~x56 & ~x57 & ~x58 & ~x59 & ~x60 & ~x61 & ~x73 & ~x74 & ~x76 & ~x77 & ~x78 & ~x80 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x86 & ~x87 & ~x88 & ~x89 & ~x101 & ~x103 & ~x104 & ~x105 & ~x106 & ~x107 & ~x108 & ~x109 & ~x110 & ~x111 & ~x112 & ~x113 & ~x114 & ~x115 & ~x116 & ~x117 & ~x130 & ~x131 & ~x132 & ~x133 & ~x134 & ~x135 & ~x136 & ~x137 & ~x138 & ~x139 & ~x141 & ~x142 & ~x143 & ~x144 & ~x160 & ~x161 & ~x162 & ~x163 & ~x165 & ~x166 & ~x167 & ~x168 & ~x169 & ~x170 & ~x171 & ~x172 & ~x173 & ~x187 & ~x189 & ~x190 & ~x191 & ~x192 & ~x193 & ~x194 & ~x195 & ~x196 & ~x197 & ~x198 & ~x199 & ~x200 & ~x201 & ~x216 & ~x217 & ~x218 & ~x219 & ~x220 & ~x221 & ~x222 & ~x223 & ~x224 & ~x225 & ~x226 & ~x227 & ~x228 & ~x245 & ~x246 & ~x248 & ~x249 & ~x250 & ~x251 & ~x252 & ~x253 & ~x254 & ~x256 & ~x274 & ~x276 & ~x277 & ~x278 & ~x279 & ~x280 & ~x281 & ~x282 & ~x283 & ~x302 & ~x303 & ~x304 & ~x305 & ~x306 & ~x307 & ~x308 & ~x309 & ~x310 & ~x311 & ~x312 & ~x329 & ~x330 & ~x331 & ~x332 & ~x333 & ~x334 & ~x335 & ~x336 & ~x337 & ~x338 & ~x359 & ~x360 & ~x361 & ~x362 & ~x363 & ~x364 & ~x365 & ~x366 & ~x368 & ~x385 & ~x387 & ~x388 & ~x389 & ~x390 & ~x391 & ~x392 & ~x393 & ~x394 & ~x414 & ~x415 & ~x416 & ~x417 & ~x418 & ~x419 & ~x420 & ~x421 & ~x422 & ~x423 & ~x442 & ~x443 & ~x444 & ~x445 & ~x446 & ~x447 & ~x448 & ~x449 & ~x450 & ~x471 & ~x472 & ~x473 & ~x474 & ~x475 & ~x476 & ~x477 & ~x478 & ~x479 & ~x480 & ~x498 & ~x500 & ~x501 & ~x502 & ~x503 & ~x504 & ~x506 & ~x526 & ~x527 & ~x528 & ~x529 & ~x530 & ~x531 & ~x532 & ~x533 & ~x534 & ~x535 & ~x555 & ~x558 & ~x559 & ~x560 & ~x561 & ~x585 & ~x586 & ~x587 & ~x588 & ~x613 & ~x614 & ~x615 & ~x616 & ~x617 & ~x640 & ~x642 & ~x643 & ~x644 & ~x645 & ~x669 & ~x671 & ~x672 & ~x673 & ~x699 & ~x700 & ~x702 & ~x726 & ~x727 & ~x728 & ~x729 & ~x730 & ~x731 & ~x753 & ~x754 & ~x756 & ~x757 & ~x758 & ~x759 & ~x781 & ~x782 & ~x783;
assign c9413 =  x267 &  x708 & ~x110 & ~x142;
assign c9415 =  x445;
assign c9417 = ~x332 & ~x346 & ~x349 & ~x374 & ~x413 & ~x414 & ~x440 & ~x722 & ~x724 & ~x728 & ~x735 & ~x748 & ~x749 & ~x750 & ~x752 & ~x777 & ~x782;
assign c9419 = ~x34 & ~x59 & ~x64 & ~x83 & ~x91 & ~x111 & ~x148 & ~x171 & ~x174 & ~x176 & ~x190 & ~x201 & ~x204 & ~x229 & ~x230 & ~x231 & ~x257 & ~x259 & ~x284 & ~x287 & ~x342 & ~x369 & ~x390 & ~x394 & ~x452 & ~x507 & ~x562 & ~x663 & ~x692;
assign c9421 =  x306 & ~x328 & ~x694;
assign c9423 =  x352 & ~x3 & ~x4 & ~x23 & ~x24 & ~x26 & ~x28 & ~x29 & ~x31 & ~x47 & ~x48 & ~x50 & ~x51 & ~x54 & ~x55 & ~x56 & ~x58 & ~x75 & ~x78 & ~x79 & ~x81 & ~x86 & ~x88 & ~x101 & ~x103 & ~x104 & ~x106 & ~x107 & ~x111 & ~x112 & ~x113 & ~x114 & ~x115 & ~x116 & ~x130 & ~x131 & ~x132 & ~x133 & ~x135 & ~x137 & ~x139 & ~x140 & ~x141 & ~x142 & ~x144 & ~x163 & ~x164 & ~x165 & ~x168 & ~x171 & ~x191 & ~x192 & ~x193 & ~x194 & ~x196 & ~x199 & ~x216 & ~x218 & ~x220 & ~x222 & ~x224 & ~x246 & ~x247 & ~x248 & ~x255 & ~x274 & ~x275 & ~x277 & ~x279 & ~x280 & ~x303 & ~x304 & ~x306 & ~x309 & ~x331 & ~x333 & ~x334 & ~x335 & ~x336 & ~x338 & ~x361 & ~x364 & ~x388 & ~x389 & ~x392 & ~x419 & ~x420 & ~x473 & ~x474 & ~x475 & ~x532 & ~x588 & ~x645 & ~x702 & ~x725 & ~x726 & ~x729 & ~x752 & ~x753 & ~x755 & ~x757 & ~x758 & ~x779 & ~x781;
assign c9425 =  x295 & ~x83 & ~x123 & ~x161 & ~x192 & ~x219 & ~x221 & ~x301 & ~x560 & ~x614 & ~x671 & ~x754 & ~x781;
assign c9427 = ~x5 & ~x30 & ~x61 & ~x314 & ~x359 & ~x370 & ~x391 & ~x398 & ~x405 & ~x406 & ~x426 & ~x444 & ~x471 & ~x502 & ~x509 & ~x665;
assign c9429 =  x232 & ~x377 & ~x386 & ~x391 & ~x413 & ~x416 & ~x423;
assign c9431 = ~x3 & ~x79 & ~x80 & ~x103 & ~x104 & ~x118 & ~x133 & ~x143 & ~x167 & ~x171 & ~x299 & ~x300 & ~x332 & ~x339 & ~x603 & ~x608 & ~x631 & ~x632 & ~x634 & ~x681 & ~x701 & ~x708 & ~x734 & ~x782;
assign c9433 =  x73 &  x213 & ~x611;
assign c9435 = ~x54 & ~x56 & ~x141 & ~x287 & ~x313 & ~x343 & ~x372 & ~x394 & ~x482 & ~x484 & ~x485 & ~x501 & ~x512 & ~x513 & ~x644 & ~x661 & ~x719 & ~x720 & ~x725 & ~x749;
assign c9437 = ~x30 & ~x36 & ~x47 & ~x82 & ~x85 & ~x86 & ~x105 & ~x106 & ~x108 & ~x135 & ~x136 & ~x144 & ~x161 & ~x165 & ~x191 & ~x195 & ~x216 & ~x225 & ~x230 & ~x231 & ~x245 & ~x248 & ~x251 & ~x252 & ~x273 & ~x283 & ~x306 & ~x308 & ~x311 & ~x312 & ~x327 & ~x336 & ~x357 & ~x358 & ~x385 & ~x389 & ~x391 & ~x415 & ~x442 & ~x443 & ~x453 & ~x472 & ~x480 & ~x499 & ~x502 & ~x505 & ~x532 & ~x730 & ~x731 & ~x752;
assign c9439 =  x516 &  x688 & ~x61 & ~x145 & ~x173 & ~x200 & ~x247 & ~x358 & ~x387;
assign c9441 = ~x26 & ~x57 & ~x91 & ~x106 & ~x107 & ~x144 & ~x163 & ~x197 & ~x203 & ~x219 & ~x233 & ~x282 & ~x303 & ~x305 & ~x366 & ~x471 & ~x503 & ~x602 & ~x603 & ~x606 & ~x759;
assign c9443 =  x305 & ~x611 & ~x637 & ~x638 & ~x665 & ~x693;
assign c9445 =  x99 & ~x23 & ~x60 & ~x87 & ~x197 & ~x279 & ~x386 & ~x388 & ~x469 & ~x496 & ~x508 & ~x525 & ~x527 & ~x614;
assign c9447 =  x133 & ~x267 & ~x485;
assign c9449 = ~x25 & ~x55 & ~x140 & ~x168 & ~x280 & ~x347 & ~x366 & ~x391 & ~x441 & ~x487 & ~x489 & ~x496 & ~x698 & ~x726 & ~x754;
assign c9451 = ~x0 & ~x5 & ~x16 & ~x28 & ~x43 & ~x54 & ~x61 & ~x78 & ~x84 & ~x112 & ~x115 & ~x117 & ~x138 & ~x141 & ~x164 & ~x165 & ~x171 & ~x221 & ~x250 & ~x252 & ~x270 & ~x271 & ~x272 & ~x304 & ~x305 & ~x306 & ~x334 & ~x337 & ~x475 & ~x502 & ~x545 & ~x547 & ~x640 & ~x646 & ~x697 & ~x728 & ~x754 & ~x758 & ~x762;
assign c9453 =  x636 & ~x194 & ~x222 & ~x278 & ~x279 & ~x280 & ~x334 & ~x361 & ~x750 & ~x751 & ~x779;
assign c9455 = ~x110 & ~x111 & ~x114 & ~x371 & ~x399 & ~x403 & ~x422 & ~x454 & ~x503 & ~x510 & ~x533 & ~x699 & ~x716 & ~x728 & ~x771;
assign c9457 =  x533 & ~x766;
assign c9459 = ~x24 & ~x26 & ~x27 & ~x55 & ~x56 & ~x58 & ~x59 & ~x83 & ~x84 & ~x85 & ~x111 & ~x113 & ~x463 & ~x464 & ~x475 & ~x492 & ~x531 & ~x547 & ~x548 & ~x575 & ~x603 & ~x631 & ~x681 & ~x700 & ~x739 & ~x757 & ~x766 & ~x767 & ~x783;
assign c9461 =  x314 &  x371 &  x398 &  x399 & ~x466;
assign c9463 =  x267 & ~x53 & ~x114 & ~x115 & ~x137 & ~x143 & ~x166 & ~x191 & ~x197 & ~x456 & ~x560 & ~x701 & ~x754 & ~x771 & ~x780;
assign c9465 =  x635 &  x663 & ~x53 & ~x109 & ~x113 & ~x137 & ~x140 & ~x142 & ~x169 & ~x193 & ~x196 & ~x197 & ~x251 & ~x254;
assign c9467 = ~x28 & ~x168 & ~x267 & ~x322 & ~x337 & ~x390 & ~x404 & ~x405 & ~x431 & ~x459 & ~x460 & ~x700 & ~x767 & ~x782;
assign c9469 =  x348 & ~x1 & ~x5 & ~x24 & ~x25 & ~x27 & ~x28 & ~x31 & ~x33 & ~x48 & ~x52 & ~x59 & ~x74 & ~x75 & ~x83 & ~x88 & ~x90 & ~x102 & ~x103 & ~x106 & ~x115 & ~x133 & ~x134 & ~x136 & ~x137 & ~x139 & ~x140 & ~x142 & ~x145 & ~x159 & ~x172 & ~x191 & ~x192 & ~x198 & ~x199 & ~x202 & ~x221 & ~x224 & ~x226 & ~x244 & ~x248 & ~x251 & ~x274 & ~x276 & ~x278 & ~x303 & ~x304 & ~x305 & ~x338 & ~x340 & ~x367 & ~x386 & ~x387 & ~x388 & ~x389 & ~x394 & ~x395 & ~x420 & ~x444 & ~x477 & ~x478 & ~x480 & ~x507 & ~x508 & ~x532 & ~x535 & ~x557 & ~x589 & ~x618 & ~x755 & ~x756;
assign c9471 = ~x101 & ~x214 & ~x242 & ~x270 & ~x357 & ~x397 & ~x411 & ~x441 & ~x479 & ~x482 & ~x603;
assign c9473 =  x152 & ~x80 & ~x81 & ~x143 & ~x421 & ~x473 & ~x546 & ~x547 & ~x600;
assign c9475 = ~x50 & ~x51 & ~x58 & ~x78 & ~x105 & ~x108 & ~x117 & ~x144 & ~x161 & ~x171 & ~x173 & ~x229 & ~x272 & ~x506 & ~x549 & ~x574 & ~x577 & ~x604 & ~x611 & ~x631 & ~x634 & ~x680;
assign c9477 = ~x295 & ~x324 & ~x351 & ~x464 & ~x519 & ~x543;
assign c9479 =  x121 & ~x646 & ~x664 & ~x670 & ~x695 & ~x698 & ~x720 & ~x721 & ~x734 & ~x746 & ~x747 & ~x749 & ~x751 & ~x752 & ~x755 & ~x757 & ~x758;
assign c9481 = ~x1 & ~x17 & ~x24 & ~x31 & ~x71 & ~x79 & ~x85 & ~x86 & ~x87 & ~x105 & ~x110 & ~x113 & ~x170 & ~x252 & ~x277 & ~x309 & ~x323 & ~x333 & ~x366 & ~x373 & ~x417 & ~x420 & ~x450 & ~x586 & ~x754 & ~x768;
assign c9483 = ~x30 & ~x47 & ~x87 & ~x89 & ~x105 & ~x134 & ~x135 & ~x145 & ~x152 & ~x159 & ~x164 & ~x171 & ~x173 & ~x190 & ~x193 & ~x198 & ~x199 & ~x301 & ~x780;
assign c9485 =  x184 & ~x23 & ~x27 & ~x29 & ~x30 & ~x56 & ~x82 & ~x140 & ~x371 & ~x397 & ~x416 & ~x446 & ~x452 & ~x453 & ~x454 & ~x474 & ~x481 & ~x700 & ~x781;
assign c9487 =  x370 &  x398 &  x426 & ~x98 & ~x242 & ~x678;
assign c9489 =  x45 & ~x120 & ~x348 & ~x486;
assign c9491 =  x264 & ~x0 & ~x30 & ~x80 & ~x108 & ~x111 & ~x168 & ~x226 & ~x254 & ~x306 & ~x349 & ~x350 & ~x471 & ~x501 & ~x507 & ~x535 & ~x755 & ~x756;
assign c9493 =  x73 & ~x309 & ~x385;
assign c9495 =  x312 & ~x81 & ~x82 & ~x224 & ~x408 & ~x433;
assign c9497 = ~x8 & ~x31 & ~x53 & ~x409 & ~x437 & ~x464 & ~x489 & ~x493 & ~x520 & ~x521 & ~x766;
assign c9499 =  x567 &  x595 & ~x324;

endmodule