module tm( x0,x1,x2,x3,x4,x5,x6,x7,x8,x9,x10,x11,x12,x13,x14,x15,x16,x17,x18,x19,x20,x21,x22,x23,x24,x25,x26,x27,x28,x29,x30,x31,x32,x33,x34,x35,x36,x37,x38,x39,x40,x41,x42,x43,x44,x45,x46,x47,x48,x49,x50,x51,x52,x53,x54,x55,x56,x57,x58,x59,x60,x61,x62,x63,x64,x65,x66,x67,x68,x69,x70,x71,x72,x73,x74,x75,x76,x77,x78,x79,x80,x81,x82,x83,x84,x85,x86,x87,x88,x89,x90,x91,x92,x93,x94,x95,x96,x97,x98,x99,x100,x101,x102,x103,x104,x105,x106,x107,x108,x109,x110,x111,x112,x113,x114,x115,x116,x117,x118,x119,x120,x121,x122,x123,x124,x125,x126,x127,x128,x129,x130,x131,x132,x133,x134,x135,x136,x137,x138,x139,x140,x141,x142,x143,x144,x145,x146,x147,x148,x149,x150,x151,x152,x153,x154,x155,x156,x157,x158,x159,x160,x161,x162,x163,x164,x165,x166,x167,x168,x169,x170,x171,x172,x173,x174,x175,x176,x177,x178,x179,x180,x181,x182,x183,x184,x185,x186,x187,x188,x189,x190,x191,x192,x193,x194,x195,x196,x197,x198,x199,x200,x201,x202,x203,x204,x205,x206,x207,x208,x209,x210,x211,x212,x213,x214,x215,x216,x217,x218,x219,x220,x221,x222,x223,x224,x225,x226,x227,x228,x229,x230,x231,x232,x233,x234,x235,x236,x237,x238,x239,x240,x241,x242,x243,x244,x245,x246,x247,x248,x249,x250,x251,x252,x253,x254,x255,x256,x257,x258,x259,x260,x261,x262,x263,x264,x265,x266,x267,x268,x269,x270,x271,x272,x273,x274,x275,x276,x277,x278,x279,x280,x281,x282,x283,x284,x285,x286,x287,x288,x289,x290,x291,x292,x293,x294,x295,x296,x297,x298,x299,x300,x301,x302,x303,x304,x305,x306,x307,x308,x309,x310,x311,x312,x313,x314,x315,x316,x317,x318,x319,x320,x321,x322,x323,c1254,c0560,c1172,c0443,c1566,c1460,c1588,c1280,c1577,c1159,c0173,c1373,c130,c1271,c1426,c1423,c169,c1197,c1470,c0231,c0242,c0206,c0284,c0485,c1495,c0439,c1578,c0316,c033,c0338,c1104,c1276,c1556,c0562,c0469,c0572,c154,c014,c0130,c0423,c0131,c187,c1391,c097,c088,c0182,c179,c1177,c0565,c0526,c0548,c1182,c1573,c1480,c0273,c136,c0203,c0126,c0496,c1274,c0493,c1251,c1505,c1560,c0156,c0544,c1387,c1435,c0483,c0208,c0567,c1264,c1394,c0481,c1440,c1576,c1481,c095,c0115,c0505,c0262,c0547,c1102,c135,c1581,c0110,c09,c185,c0277,c0291,c1528,c1108,c1382,c193,c144,c0459,c0527,c0365,c1113,c1357,c0204,c0234,c0410,c0159,c0399,c1220,c1562,c1401,c0444,c0116,c1356,c1354,c1595,c1317,c0205,c0337,c0364,c1138,c0592,c0350,c0180,c1257,c1329,c0289,c021,c196,c0335,c1393,c1273,c1451,c0134,c0224,c1530,c0343,c1170,c0557,c0490,c0128,c1477,c0161,c1375,c0144,c0461,c1244,c1115,c0569,c0430,c1390,c1389,c177,c1285,c0595,c0452,c1313,c1455,c082,c1561,c1352,c1240,c1359,c047,c0556,c1453,c1221,c0402,c1307,c1133,c0422,c1157,c0373,c1139,c0523,c0340,c1281,c0346,c019,c0293,c0323,c1164,c1342,c1124,c1410,c0228,c0475,c0396,c1272,c1123,c0453,c1315,c1433,c0362,c0207,c020,c142,c1210,c0164,c114,c1494,c1325,c0491,c0448,c1176,c1223,c0146,c0278,c0458,c1100,c125,c0122,c085,c178,c1370,c057,c1169,c0319,c0286,c0468,c0516,c0209,c1484,c1506,c1259,c098,c0441,c1184,c1550,c1568,c1424,c0139,c1186,c0584,c0473,c065,c176,c0106,c1542,c1118,c1181,c1472,c1537,c1473,c1127,c1487,c0219,c0158,c0237,c18,c1296,c1203,c0514,c198,c1405,c0247,c1485,c1567,c0541,c16,c0359,c1112,c110,c1166,c1348,c197,c069,c1450,c0433,c0446,c059,c1585,c0260,c1142,c1427,c1597,c1187,c016,c1199,c0412,c063,c1458,c1361,c1366,c018,c186,c1103,c1572,c1589,c1217,c078,c0288,c0290,c1336,c1462,c139,c1582,c1156,c091,c0489,c127,c08,c0425,c160,c1409,c1431,c1493,c1551,c0332,c0409,c1490,c0268,c0258,c1143,c0141,c0357,c1149,c0306,c1403,c056,c1583,c0303,c1587,c066,c0507,c184,c1237,c1422,c0255,c1362,c00,c1498,c0368,c0371,c1419,c183,c0404,c046,c180,c1488,c129,c037,c19,c1529,c1299,c0581,c1541,c0176,c0460,c0317,c148,c1564,c1479,c1309,c0213,c0521,c0154,c0244,c1209,c0401,c1231,c1492,c1260,c1128,c0384,c0271,c1368,c199,c0326,c0484,c0598,c1412,c0478,c1324,c1253,c0480,c128,c1126,c1552,c162,c0358,c1467,c1464,c1226,c194,c149,c0202,c0539,c0543,c0295,c1243,c1141,c1442,c173,c0440,c0225,c1160,c0536,c060,c0442,c029,c1500,c1167,c1267,c0499,c0486,c0554,c096,c0349,c0381,c140,c1286,c0117,c0152,c0166,c0416,c1318,c0127,c0217,c1183,c182,c0573,c0570,c1507,c0515,c0511,c0179,c0533,c0298,c1413,c04,c0472,c1534,c1547,c0162,c011,c0467,c081,c1398,c1219,c0347,c0575,c1386,c159,c137,c0148,c0568,c077,c165,c0451,c0197,c0502,c1486,c071,c1596,c0385,c0125,c1563,c1591,c1311,c0108,c1255,c0253,c025,c1346,c0477,c1289,c0354,c0531,c0160,c1117,c1445,c0417,c158,c0553,c157,c076,c111,c0574,c0545,c0456,c1408,c0353,c1555,c1465,c0342,c118,c1165,c0307,c0590,c1206,c053,c0263,c0324,c1543,c1283,c1469,c1147,c1208,c0339,c171,c1175,c0427,c0438,c0360,c1351,c1457,c0518,c0378,c1153,c1436,c1163,c036,c073,c0397,c0103,c0487,c039,c0457,c1101,c0375,c1353,c1459,c1234,c0114,c0200,c07,c0285,c1122,c0445,c0328,c0394,c122,c0194,c0227,c167,c1151,c0420,c1508,c11,c0129,c0538,c0509,c1238,c0413,c0415,c1111,c0281,c092,c152,c1499,c0157,c0563,c1407,c1202,c074,c1252,c1345,c0257,c190,c0239,c0411,c1476,c1198,c1168,c0226,c1288,c0382,c0177,c1132,c0153,c05,c0546,c1235,c1570,c1593,c0230,c1554,c044,c1385,c0535,c0185,c022,c072,c0591,c0344,c0132,c0232,c1590,c1188,c1355,c1383,c1193,c1228,c062,c0418,c1497,c034,c0240,c0193,c0261,c1270,c0503,c1449,c1247,c094,c1200,c166,c0336,c1162,c0169,c1278,c1392,c1178,c145,c02,c1416,c0550,c026,c1524,c0241,c0351,c1207,c1399,c1429,c01,c1279,c0571,c1310,c1349,c0308,c0313,c1146,c1192,c1224,c0149,c1502,c1292,c1293,c1214,c0549,c0426,c1190,c0388,c0434,c1434,c1107,c1579,c0333,c0264,c0348,c0579,c06,c1430,c1265,c040,c1300,c0530,c0168,c0107,c1438,c1452,c1548,c0165,c1250,c1179,c0294,c0431,c0120,c1420,c1205,c0250,c1526,c0407,c0133,c043,c121,c1417,c1191,c1491,c1535,c174,c028,c1599,c0501,c012,c1131,c151,c1303,c1371,c0525,c1249,c146,c0498,c0561,c0424,c1114,c0379,c113,c1565,c0455,c0589,c0100,c0198,c172,c1444,c0566,c0214,c068,c0196,c116,c1195,c1475,c1148,c156,c1538,c1531,c0189,c1376,c195,c1261,c1363,c1174,c058,c0513,c1268,c0529,c133,c1135,c112,c0155,c0462,c0296,c0292,c1482,c0534,c1109,c1580,c0474,c1246,c0540,c0245,c1521,c0147,c1461,c1374,c0356,c084,c0386,c0135,c150,c1532,c161,c1327,c0184,c0283,c1212,c0421,c0435,c0576,c0450,c0520,c1194,c0594,c0597,c1504,c0265,c0138,c0593,c0512,c1294,c1343,c1216,c1245,c1395,c1236,c1338,c0118,c015,c0140,c0183,c03,c1322,c1134,c1364,c061,c0287,c0398,c0243,c1189,c1574,c1367,c1312,c0429,c1125,c075,c052,c1155,c1379,c1308,c0587,c1544,c0508,c0437,c0192,c0406,c0471,c1277,c1145,c0248,c0464,c0408,c0275,c1432,c0220,c1592,c1347,c1468,c032,c049,c1263,c1204,c086,c143,c1341,c0121,c0270,c1384,c1522,c1443,c0201,c0235,c0389,c0510,c0367,c1333,c1350,c1397,c0136,c1402,c12,c0238,c1594,c0470,c1518,c1284,c189,c079,c0476,c1161,c0187,c0327,c0387,c10,c1150,c1489,c1512,c1171,c1400,c0272,c1425,c1137,c0274,c048,c1509,c115,c045,c0330,c0580,c1287,c087,c070,c0400,c0150,c0119,c1242,c1306,c1414,c035,c1304,c1540,c1229,c1513,c1258,c1337,c141,c0370,c1319,c0376,c1569,c181,c1330,c123,c1471,c1144,c1421,c1586,c0123,c14,c1523,c0178,c0331,c1339,c0211,c0414,c0552,c0267,c1130,c1290,c1514,c1557,c1533,c1316,c0341,c1515,c1227,c175,c1331,c1428,c0256,c0345,c0532,c1369,c1332,c0186,c0403,c0311,c1314,c1388,c1437,c1344,c132,c1404,c1335,c0102,c1116,c027,c0105,c0583,c0558,c1291,c1483,c0352,c1106,c1525,c0428,c0251,c0463,c0174,c0419,c0304,c1456,c164,c170,c054,c089,c0301,c1553,c1232,c0266,c1380,c0586,c0555,c013,c0221,c0392,c1448,c0218,c031,c0195,c0494,c1323,c1282,c1381,c0318,c1520,c0504,c0190,c1519,c024,c1154,c0297,c017,c055,c038,c0151,c0391,c083,c0577,c1152,c147,c1211,c1269,c1501,c099,c1396,c1545,c0322,c0537,c0374,c0145,c120,c1158,c0212,c0143,c1510,c0334,c0111,c0223,c0355,c023,c153,c1120,c0432,c093,c0578,c0113,c0361,c0312,c1503,c1546,c1446,c0393,c1340,c1119,c0390,c0259,c1358,c15,c050,c0142,c0363,c0395,c1262,c0181,c0124,c17,c0320,c1230,c041,c134,c1527,c0321,c1539,c0405,c0599,c1233,c0488,c0310,c0236,c0369,c1320,c0377,c0582,c1466,c1275,c1295,c0522,c1511,c1110,c1239,c0191,c0495,c0249,c0137,c0559,c080,c1321,c0482,c1365,c1196,c0112,c030,c0172,c0454,c0325,c0542,c1297,c1439,c0436,c0276,c168,c1136,c1406,c1478,c0500,c1378,c0517,c188,c1180,c090,c0170,c1218,c1185,c191,c1121,c1213,c0216,c0588,c1305,c0280,c0528,c0305,c0519,c163,c0104,c192,c0282,c1372,c1215,c0465,c051,c0329,c1256,c0269,c0524,c0163,c0551,c1377,c0254,c1140,c0233,c1201,c1496,c0564,c1454,c0167,c1598,c138,c0380,c0302,c1302,c0497,c1298,c1517,c155,c131,c1173,c0188,c0215,c0101,c0309,c124,c117,c0492,c1575,c0109,c0252,c1558,c0300,c0506,c0246,c0229,c0585,c1301,c1571,c0366,c1326,c0479,c1241,c1536,c0383,c1129,c1418,c1225,c0466,c067,c1222,c1415,c0175,c0596,c0315,c010,c0199,c0447,c13,c1411,c1105,c1463,c1516,c0279,c0299,c126,c119,c0210,c0314,c0222,c1328,c1447,c1334,c1360,c1474,c1549,c0372,c064,c042,c0171,c0449,c1559,c1248,c1266,c1584,c1441 );

input x0;
input x1;
input x2;
input x3;
input x4;
input x5;
input x6;
input x7;
input x8;
input x9;
input x10;
input x11;
input x12;
input x13;
input x14;
input x15;
input x16;
input x17;
input x18;
input x19;
input x20;
input x21;
input x22;
input x23;
input x24;
input x25;
input x26;
input x27;
input x28;
input x29;
input x30;
input x31;
input x32;
input x33;
input x34;
input x35;
input x36;
input x37;
input x38;
input x39;
input x40;
input x41;
input x42;
input x43;
input x44;
input x45;
input x46;
input x47;
input x48;
input x49;
input x50;
input x51;
input x52;
input x53;
input x54;
input x55;
input x56;
input x57;
input x58;
input x59;
input x60;
input x61;
input x62;
input x63;
input x64;
input x65;
input x66;
input x67;
input x68;
input x69;
input x70;
input x71;
input x72;
input x73;
input x74;
input x75;
input x76;
input x77;
input x78;
input x79;
input x80;
input x81;
input x82;
input x83;
input x84;
input x85;
input x86;
input x87;
input x88;
input x89;
input x90;
input x91;
input x92;
input x93;
input x94;
input x95;
input x96;
input x97;
input x98;
input x99;
input x100;
input x101;
input x102;
input x103;
input x104;
input x105;
input x106;
input x107;
input x108;
input x109;
input x110;
input x111;
input x112;
input x113;
input x114;
input x115;
input x116;
input x117;
input x118;
input x119;
input x120;
input x121;
input x122;
input x123;
input x124;
input x125;
input x126;
input x127;
input x128;
input x129;
input x130;
input x131;
input x132;
input x133;
input x134;
input x135;
input x136;
input x137;
input x138;
input x139;
input x140;
input x141;
input x142;
input x143;
input x144;
input x145;
input x146;
input x147;
input x148;
input x149;
input x150;
input x151;
input x152;
input x153;
input x154;
input x155;
input x156;
input x157;
input x158;
input x159;
input x160;
input x161;
input x162;
input x163;
input x164;
input x165;
input x166;
input x167;
input x168;
input x169;
input x170;
input x171;
input x172;
input x173;
input x174;
input x175;
input x176;
input x177;
input x178;
input x179;
input x180;
input x181;
input x182;
input x183;
input x184;
input x185;
input x186;
input x187;
input x188;
input x189;
input x190;
input x191;
input x192;
input x193;
input x194;
input x195;
input x196;
input x197;
input x198;
input x199;
input x200;
input x201;
input x202;
input x203;
input x204;
input x205;
input x206;
input x207;
input x208;
input x209;
input x210;
input x211;
input x212;
input x213;
input x214;
input x215;
input x216;
input x217;
input x218;
input x219;
input x220;
input x221;
input x222;
input x223;
input x224;
input x225;
input x226;
input x227;
input x228;
input x229;
input x230;
input x231;
input x232;
input x233;
input x234;
input x235;
input x236;
input x237;
input x238;
input x239;
input x240;
input x241;
input x242;
input x243;
input x244;
input x245;
input x246;
input x247;
input x248;
input x249;
input x250;
input x251;
input x252;
input x253;
input x254;
input x255;
input x256;
input x257;
input x258;
input x259;
input x260;
input x261;
input x262;
input x263;
input x264;
input x265;
input x266;
input x267;
input x268;
input x269;
input x270;
input x271;
input x272;
input x273;
input x274;
input x275;
input x276;
input x277;
input x278;
input x279;
input x280;
input x281;
input x282;
input x283;
input x284;
input x285;
input x286;
input x287;
input x288;
input x289;
input x290;
input x291;
input x292;
input x293;
input x294;
input x295;
input x296;
input x297;
input x298;
input x299;
input x300;
input x301;
input x302;
input x303;
input x304;
input x305;
input x306;
input x307;
input x308;
input x309;
input x310;
input x311;
input x312;
input x313;
input x314;
input x315;
input x316;
input x317;
input x318;
input x319;
input x320;
input x321;
input x322;
input x323;
output c1254;
output c0560;
output c1172;
output c0443;
output c1566;
output c1460;
output c1588;
output c1280;
output c1577;
output c1159;
output c0173;
output c1373;
output c130;
output c1271;
output c1426;
output c1423;
output c169;
output c1197;
output c1470;
output c0231;
output c0242;
output c0206;
output c0284;
output c0485;
output c1495;
output c0439;
output c1578;
output c0316;
output c033;
output c0338;
output c1104;
output c1276;
output c1556;
output c0562;
output c0469;
output c0572;
output c154;
output c014;
output c0130;
output c0423;
output c0131;
output c187;
output c1391;
output c097;
output c088;
output c0182;
output c179;
output c1177;
output c0565;
output c0526;
output c0548;
output c1182;
output c1573;
output c1480;
output c0273;
output c136;
output c0203;
output c0126;
output c0496;
output c1274;
output c0493;
output c1251;
output c1505;
output c1560;
output c0156;
output c0544;
output c1387;
output c1435;
output c0483;
output c0208;
output c0567;
output c1264;
output c1394;
output c0481;
output c1440;
output c1576;
output c1481;
output c095;
output c0115;
output c0505;
output c0262;
output c0547;
output c1102;
output c135;
output c1581;
output c0110;
output c09;
output c185;
output c0277;
output c0291;
output c1528;
output c1108;
output c1382;
output c193;
output c144;
output c0459;
output c0527;
output c0365;
output c1113;
output c1357;
output c0204;
output c0234;
output c0410;
output c0159;
output c0399;
output c1220;
output c1562;
output c1401;
output c0444;
output c0116;
output c1356;
output c1354;
output c1595;
output c1317;
output c0205;
output c0337;
output c0364;
output c1138;
output c0592;
output c0350;
output c0180;
output c1257;
output c1329;
output c0289;
output c021;
output c196;
output c0335;
output c1393;
output c1273;
output c1451;
output c0134;
output c0224;
output c1530;
output c0343;
output c1170;
output c0557;
output c0490;
output c0128;
output c1477;
output c0161;
output c1375;
output c0144;
output c0461;
output c1244;
output c1115;
output c0569;
output c0430;
output c1390;
output c1389;
output c177;
output c1285;
output c0595;
output c0452;
output c1313;
output c1455;
output c082;
output c1561;
output c1352;
output c1240;
output c1359;
output c047;
output c0556;
output c1453;
output c1221;
output c0402;
output c1307;
output c1133;
output c0422;
output c1157;
output c0373;
output c1139;
output c0523;
output c0340;
output c1281;
output c0346;
output c019;
output c0293;
output c0323;
output c1164;
output c1342;
output c1124;
output c1410;
output c0228;
output c0475;
output c0396;
output c1272;
output c1123;
output c0453;
output c1315;
output c1433;
output c0362;
output c0207;
output c020;
output c142;
output c1210;
output c0164;
output c114;
output c1494;
output c1325;
output c0491;
output c0448;
output c1176;
output c1223;
output c0146;
output c0278;
output c0458;
output c1100;
output c125;
output c0122;
output c085;
output c178;
output c1370;
output c057;
output c1169;
output c0319;
output c0286;
output c0468;
output c0516;
output c0209;
output c1484;
output c1506;
output c1259;
output c098;
output c0441;
output c1184;
output c1550;
output c1568;
output c1424;
output c0139;
output c1186;
output c0584;
output c0473;
output c065;
output c176;
output c0106;
output c1542;
output c1118;
output c1181;
output c1472;
output c1537;
output c1473;
output c1127;
output c1487;
output c0219;
output c0158;
output c0237;
output c18;
output c1296;
output c1203;
output c0514;
output c198;
output c1405;
output c0247;
output c1485;
output c1567;
output c0541;
output c16;
output c0359;
output c1112;
output c110;
output c1166;
output c1348;
output c197;
output c069;
output c1450;
output c0433;
output c0446;
output c059;
output c1585;
output c0260;
output c1142;
output c1427;
output c1597;
output c1187;
output c016;
output c1199;
output c0412;
output c063;
output c1458;
output c1361;
output c1366;
output c018;
output c186;
output c1103;
output c1572;
output c1589;
output c1217;
output c078;
output c0288;
output c0290;
output c1336;
output c1462;
output c139;
output c1582;
output c1156;
output c091;
output c0489;
output c127;
output c08;
output c0425;
output c160;
output c1409;
output c1431;
output c1493;
output c1551;
output c0332;
output c0409;
output c1490;
output c0268;
output c0258;
output c1143;
output c0141;
output c0357;
output c1149;
output c0306;
output c1403;
output c056;
output c1583;
output c0303;
output c1587;
output c066;
output c0507;
output c184;
output c1237;
output c1422;
output c0255;
output c1362;
output c00;
output c1498;
output c0368;
output c0371;
output c1419;
output c183;
output c0404;
output c046;
output c180;
output c1488;
output c129;
output c037;
output c19;
output c1529;
output c1299;
output c0581;
output c1541;
output c0176;
output c0460;
output c0317;
output c148;
output c1564;
output c1479;
output c1309;
output c0213;
output c0521;
output c0154;
output c0244;
output c1209;
output c0401;
output c1231;
output c1492;
output c1260;
output c1128;
output c0384;
output c0271;
output c1368;
output c199;
output c0326;
output c0484;
output c0598;
output c1412;
output c0478;
output c1324;
output c1253;
output c0480;
output c128;
output c1126;
output c1552;
output c162;
output c0358;
output c1467;
output c1464;
output c1226;
output c194;
output c149;
output c0202;
output c0539;
output c0543;
output c0295;
output c1243;
output c1141;
output c1442;
output c173;
output c0440;
output c0225;
output c1160;
output c0536;
output c060;
output c0442;
output c029;
output c1500;
output c1167;
output c1267;
output c0499;
output c0486;
output c0554;
output c096;
output c0349;
output c0381;
output c140;
output c1286;
output c0117;
output c0152;
output c0166;
output c0416;
output c1318;
output c0127;
output c0217;
output c1183;
output c182;
output c0573;
output c0570;
output c1507;
output c0515;
output c0511;
output c0179;
output c0533;
output c0298;
output c1413;
output c04;
output c0472;
output c1534;
output c1547;
output c0162;
output c011;
output c0467;
output c081;
output c1398;
output c1219;
output c0347;
output c0575;
output c1386;
output c159;
output c137;
output c0148;
output c0568;
output c077;
output c165;
output c0451;
output c0197;
output c0502;
output c1486;
output c071;
output c1596;
output c0385;
output c0125;
output c1563;
output c1591;
output c1311;
output c0108;
output c1255;
output c0253;
output c025;
output c1346;
output c0477;
output c1289;
output c0354;
output c0531;
output c0160;
output c1117;
output c1445;
output c0417;
output c158;
output c0553;
output c157;
output c076;
output c111;
output c0574;
output c0545;
output c0456;
output c1408;
output c0353;
output c1555;
output c1465;
output c0342;
output c118;
output c1165;
output c0307;
output c0590;
output c1206;
output c053;
output c0263;
output c0324;
output c1543;
output c1283;
output c1469;
output c1147;
output c1208;
output c0339;
output c171;
output c1175;
output c0427;
output c0438;
output c0360;
output c1351;
output c1457;
output c0518;
output c0378;
output c1153;
output c1436;
output c1163;
output c036;
output c073;
output c0397;
output c0103;
output c0487;
output c039;
output c0457;
output c1101;
output c0375;
output c1353;
output c1459;
output c1234;
output c0114;
output c0200;
output c07;
output c0285;
output c1122;
output c0445;
output c0328;
output c0394;
output c122;
output c0194;
output c0227;
output c167;
output c1151;
output c0420;
output c1508;
output c11;
output c0129;
output c0538;
output c0509;
output c1238;
output c0413;
output c0415;
output c1111;
output c0281;
output c092;
output c152;
output c1499;
output c0157;
output c0563;
output c1407;
output c1202;
output c074;
output c1252;
output c1345;
output c0257;
output c190;
output c0239;
output c0411;
output c1476;
output c1198;
output c1168;
output c0226;
output c1288;
output c0382;
output c0177;
output c1132;
output c0153;
output c05;
output c0546;
output c1235;
output c1570;
output c1593;
output c0230;
output c1554;
output c044;
output c1385;
output c0535;
output c0185;
output c022;
output c072;
output c0591;
output c0344;
output c0132;
output c0232;
output c1590;
output c1188;
output c1355;
output c1383;
output c1193;
output c1228;
output c062;
output c0418;
output c1497;
output c034;
output c0240;
output c0193;
output c0261;
output c1270;
output c0503;
output c1449;
output c1247;
output c094;
output c1200;
output c166;
output c0336;
output c1162;
output c0169;
output c1278;
output c1392;
output c1178;
output c145;
output c02;
output c1416;
output c0550;
output c026;
output c1524;
output c0241;
output c0351;
output c1207;
output c1399;
output c1429;
output c01;
output c1279;
output c0571;
output c1310;
output c1349;
output c0308;
output c0313;
output c1146;
output c1192;
output c1224;
output c0149;
output c1502;
output c1292;
output c1293;
output c1214;
output c0549;
output c0426;
output c1190;
output c0388;
output c0434;
output c1434;
output c1107;
output c1579;
output c0333;
output c0264;
output c0348;
output c0579;
output c06;
output c1430;
output c1265;
output c040;
output c1300;
output c0530;
output c0168;
output c0107;
output c1438;
output c1452;
output c1548;
output c0165;
output c1250;
output c1179;
output c0294;
output c0431;
output c0120;
output c1420;
output c1205;
output c0250;
output c1526;
output c0407;
output c0133;
output c043;
output c121;
output c1417;
output c1191;
output c1491;
output c1535;
output c174;
output c028;
output c1599;
output c0501;
output c012;
output c1131;
output c151;
output c1303;
output c1371;
output c0525;
output c1249;
output c146;
output c0498;
output c0561;
output c0424;
output c1114;
output c0379;
output c113;
output c1565;
output c0455;
output c0589;
output c0100;
output c0198;
output c172;
output c1444;
output c0566;
output c0214;
output c068;
output c0196;
output c116;
output c1195;
output c1475;
output c1148;
output c156;
output c1538;
output c1531;
output c0189;
output c1376;
output c195;
output c1261;
output c1363;
output c1174;
output c058;
output c0513;
output c1268;
output c0529;
output c133;
output c1135;
output c112;
output c0155;
output c0462;
output c0296;
output c0292;
output c1482;
output c0534;
output c1109;
output c1580;
output c0474;
output c1246;
output c0540;
output c0245;
output c1521;
output c0147;
output c1461;
output c1374;
output c0356;
output c084;
output c0386;
output c0135;
output c150;
output c1532;
output c161;
output c1327;
output c0184;
output c0283;
output c1212;
output c0421;
output c0435;
output c0576;
output c0450;
output c0520;
output c1194;
output c0594;
output c0597;
output c1504;
output c0265;
output c0138;
output c0593;
output c0512;
output c1294;
output c1343;
output c1216;
output c1245;
output c1395;
output c1236;
output c1338;
output c0118;
output c015;
output c0140;
output c0183;
output c03;
output c1322;
output c1134;
output c1364;
output c061;
output c0287;
output c0398;
output c0243;
output c1189;
output c1574;
output c1367;
output c1312;
output c0429;
output c1125;
output c075;
output c052;
output c1155;
output c1379;
output c1308;
output c0587;
output c1544;
output c0508;
output c0437;
output c0192;
output c0406;
output c0471;
output c1277;
output c1145;
output c0248;
output c0464;
output c0408;
output c0275;
output c1432;
output c0220;
output c1592;
output c1347;
output c1468;
output c032;
output c049;
output c1263;
output c1204;
output c086;
output c143;
output c1341;
output c0121;
output c0270;
output c1384;
output c1522;
output c1443;
output c0201;
output c0235;
output c0389;
output c0510;
output c0367;
output c1333;
output c1350;
output c1397;
output c0136;
output c1402;
output c12;
output c0238;
output c1594;
output c0470;
output c1518;
output c1284;
output c189;
output c079;
output c0476;
output c1161;
output c0187;
output c0327;
output c0387;
output c10;
output c1150;
output c1489;
output c1512;
output c1171;
output c1400;
output c0272;
output c1425;
output c1137;
output c0274;
output c048;
output c1509;
output c115;
output c045;
output c0330;
output c0580;
output c1287;
output c087;
output c070;
output c0400;
output c0150;
output c0119;
output c1242;
output c1306;
output c1414;
output c035;
output c1304;
output c1540;
output c1229;
output c1513;
output c1258;
output c1337;
output c141;
output c0370;
output c1319;
output c0376;
output c1569;
output c181;
output c1330;
output c123;
output c1471;
output c1144;
output c1421;
output c1586;
output c0123;
output c14;
output c1523;
output c0178;
output c0331;
output c1339;
output c0211;
output c0414;
output c0552;
output c0267;
output c1130;
output c1290;
output c1514;
output c1557;
output c1533;
output c1316;
output c0341;
output c1515;
output c1227;
output c175;
output c1331;
output c1428;
output c0256;
output c0345;
output c0532;
output c1369;
output c1332;
output c0186;
output c0403;
output c0311;
output c1314;
output c1388;
output c1437;
output c1344;
output c132;
output c1404;
output c1335;
output c0102;
output c1116;
output c027;
output c0105;
output c0583;
output c0558;
output c1291;
output c1483;
output c0352;
output c1106;
output c1525;
output c0428;
output c0251;
output c0463;
output c0174;
output c0419;
output c0304;
output c1456;
output c164;
output c170;
output c054;
output c089;
output c0301;
output c1553;
output c1232;
output c0266;
output c1380;
output c0586;
output c0555;
output c013;
output c0221;
output c0392;
output c1448;
output c0218;
output c031;
output c0195;
output c0494;
output c1323;
output c1282;
output c1381;
output c0318;
output c1520;
output c0504;
output c0190;
output c1519;
output c024;
output c1154;
output c0297;
output c017;
output c055;
output c038;
output c0151;
output c0391;
output c083;
output c0577;
output c1152;
output c147;
output c1211;
output c1269;
output c1501;
output c099;
output c1396;
output c1545;
output c0322;
output c0537;
output c0374;
output c0145;
output c120;
output c1158;
output c0212;
output c0143;
output c1510;
output c0334;
output c0111;
output c0223;
output c0355;
output c023;
output c153;
output c1120;
output c0432;
output c093;
output c0578;
output c0113;
output c0361;
output c0312;
output c1503;
output c1546;
output c1446;
output c0393;
output c1340;
output c1119;
output c0390;
output c0259;
output c1358;
output c15;
output c050;
output c0142;
output c0363;
output c0395;
output c1262;
output c0181;
output c0124;
output c17;
output c0320;
output c1230;
output c041;
output c134;
output c1527;
output c0321;
output c1539;
output c0405;
output c0599;
output c1233;
output c0488;
output c0310;
output c0236;
output c0369;
output c1320;
output c0377;
output c0582;
output c1466;
output c1275;
output c1295;
output c0522;
output c1511;
output c1110;
output c1239;
output c0191;
output c0495;
output c0249;
output c0137;
output c0559;
output c080;
output c1321;
output c0482;
output c1365;
output c1196;
output c0112;
output c030;
output c0172;
output c0454;
output c0325;
output c0542;
output c1297;
output c1439;
output c0436;
output c0276;
output c168;
output c1136;
output c1406;
output c1478;
output c0500;
output c1378;
output c0517;
output c188;
output c1180;
output c090;
output c0170;
output c1218;
output c1185;
output c191;
output c1121;
output c1213;
output c0216;
output c0588;
output c1305;
output c0280;
output c0528;
output c0305;
output c0519;
output c163;
output c0104;
output c192;
output c0282;
output c1372;
output c1215;
output c0465;
output c051;
output c0329;
output c1256;
output c0269;
output c0524;
output c0163;
output c0551;
output c1377;
output c0254;
output c1140;
output c0233;
output c1201;
output c1496;
output c0564;
output c1454;
output c0167;
output c1598;
output c138;
output c0380;
output c0302;
output c1302;
output c0497;
output c1298;
output c1517;
output c155;
output c131;
output c1173;
output c0188;
output c0215;
output c0101;
output c0309;
output c124;
output c117;
output c0492;
output c1575;
output c0109;
output c0252;
output c1558;
output c0300;
output c0506;
output c0246;
output c0229;
output c0585;
output c1301;
output c1571;
output c0366;
output c1326;
output c0479;
output c1241;
output c1536;
output c0383;
output c1129;
output c1418;
output c1225;
output c0466;
output c067;
output c1222;
output c1415;
output c0175;
output c0596;
output c0315;
output c010;
output c0199;
output c0447;
output c13;
output c1411;
output c1105;
output c1463;
output c1516;
output c0279;
output c0299;
output c126;
output c119;
output c0210;
output c0314;
output c0222;
output c1328;
output c1447;
output c1334;
output c1360;
output c1474;
output c1549;
output c0372;
output c064;
output c042;
output c0171;
output c0449;
output c1559;
output c1248;
output c1266;
output c1584;
output c1441;

assign c00 = ~x4 & ~x22 & ~x60 & ~x154;
assign c02 =  x25 &  x92 &  x240 &  x258 & ~x223;
assign c04 =  x285 &  x289 &  x312 & ~x174;
assign c06 =  x96 &  x155 &  x319 & ~x219;
assign c08 =  x12 &  x225 &  x277 & ~x220;
assign c010 =  x292 & ~x242 & ~x261;
assign c012 =  x151 &  x277 &  x296 & ~x288;
assign c014 =  x191 &  x231 & ~x63 & ~x71;
assign c016 =  x264 & ~x154;
assign c018 =  x133 &  x321 &  x322 & ~x302;
assign c020 =  x68 & ~x295 & ~x313 & ~x317 & ~x319;
assign c022 =  x150 &  x240 &  x269 &  x312;
assign c024 = ~x99 & ~x147 & ~x295 & ~x318;
assign c026 =  x43 & ~x100 & ~x133 & ~x257;
assign c028 =  x49 &  x148 & ~x270;
assign c030 = ~x102 & ~x193 & ~x281;
assign c032 =  x103 &  x312 & ~x302;
assign c034 = ~x6 & ~x37 & ~x60 & ~x168 & ~x220;
assign c036 =  x55 & ~x214 & ~x236 & ~x237;
assign c038 =  x263 & ~x30 & ~x39 & ~x174 & ~x199;
assign c040 =  x287 &  x317 & ~x203;
assign c042 =  x110 &  x319 & ~x126;
assign c044 =  x139 &  x150 & ~x192;
assign c046 =  x264 & ~x96 & ~x106 & ~x107;
assign c048 =  x82 &  x212 &  x226;
assign c050 =  x159 &  x168 & ~x75;
assign c052 =  x68 &  x87 & ~x8 & ~x268;
assign c054 =  x230 &  x257 & ~x308;
assign c056 =  x31 &  x101 &  x193 &  x266 &  x269;
assign c058 =  x95 &  x135 &  x203 & ~x132;
assign c060 =  x65 &  x182 & ~x197;
assign c062 =  x143 &  x229 & ~x185;
assign c064 =  x142 & ~x108 & ~x157 & ~x309;
assign c066 =  x78 &  x186 &  x235 & ~x156;
assign c068 = ~x93 & ~x148 & ~x223;
assign c070 =  x321 & ~x153 & ~x246;
assign c072 =  x64 &  x226 & ~x79;
assign c074 = ~x121 & ~x161 & ~x316;
assign c076 =  x83 &  x268 &  x293 &  x316;
assign c078 =  x25 & ~x105 & ~x180 & ~x262;
assign c080 =  x38 &  x94 & ~x14;
assign c082 =  x96 &  x258 & ~x39 & ~x64;
assign c084 =  x203 &  x222 & ~x214;
assign c086 =  x23 &  x101 &  x112 &  x303;
assign c088 =  x285 & ~x84 & ~x291;
assign c090 =  x89 & ~x54 & ~x166;
assign c092 =  x51 &  x133 & ~x248;
assign c094 =  x264 &  x277 & ~x107 & ~x127;
assign c096 =  x115 &  x142 &  x144 & ~x319;
assign c098 =  x24 &  x51 &  x78 &  x96 & ~x21 & ~x43 & ~x142;
assign c0100 =  x57 & ~x152 & ~x265 & ~x287;
assign c0102 =  x15 &  x303 & ~x295 & ~x309;
assign c0104 =  x96 &  x258 &  x315 & ~x48;
assign c0106 =  x132 &  x244 & ~x202 & ~x259;
assign c0108 =  x15 &  x307 & ~x10;
assign c0110 =  x43 &  x89 & ~x99 & ~x136;
assign c0112 =  x20 &  x128 & ~x162 & ~x189 & ~x192;
assign c0114 =  x25 & ~x105 & ~x274;
assign c0116 =  x47 &  x240 &  x269 & ~x105;
assign c0118 =  x259 & ~x19 & ~x113;
assign c0120 =  x93 & ~x183;
assign c0122 = ~x45 & ~x102 & ~x154 & ~x157 & ~x194;
assign c0124 =  x133 &  x308 & ~x275;
assign c0126 =  x285 & ~x291;
assign c0128 =  x62 & ~x270 & ~x300;
assign c0130 =  x157 &  x161 &  x266 &  x305;
assign c0132 =  x51 &  x78 &  x262 &  x290 & ~x264;
assign c0134 =  x16 &  x52 &  x84 & ~x49;
assign c0136 =  x12 & ~x159 & ~x274 & ~x303;
assign c0138 =  x128 &  x256 &  x294;
assign c0140 =  x182 & ~x36 & ~x127 & ~x228 & ~x266;
assign c0142 =  x67 &  x206 &  x240 &  x287 & ~x142;
assign c0144 =  x42 &  x188 & ~x120;
assign c0146 =  x76 &  x247 &  x264 &  x305 &  x316;
assign c0148 =  x38 &  x200 &  x245 &  x267 & ~x153;
assign c0150 =  x39 &  x187 & ~x262 & ~x288;
assign c0152 =  x25 &  x110 &  x164 &  x200 &  x272 & ~x112;
assign c0154 =  x76 &  x96 &  x319 & ~x176 & ~x204;
assign c0156 =  x26 &  x79 &  x106;
assign c0158 =  x26 & ~x86 & ~x116 & ~x224;
assign c0160 = ~x128 & ~x312 & ~x315;
assign c0162 =  x94 &  x240 & ~x111 & ~x165;
assign c0164 =  x96 &  x150 & ~x12 & ~x275;
assign c0166 =  x123 & ~x12 & ~x64;
assign c0168 =  x81 &  x112 & ~x115 & ~x230 & ~x244;
assign c0170 =  x103 &  x106 &  x132 &  x242 &  x256 &  x294;
assign c0172 =  x102 & ~x13 & ~x95 & ~x100;
assign c0174 =  x101 &  x133 &  x157 &  x158 &  x161;
assign c0176 =  x290 & ~x111 & ~x264;
assign c0178 =  x101 &  x236 &  x266 & ~x212;
assign c0180 =  x52 &  x240 & ~x36 & ~x198 & ~x301;
assign c0182 =  x236 &  x303 & ~x105 & ~x133;
assign c0184 =  x190 & ~x157 & ~x169 & ~x319;
assign c0186 = ~x273 & ~x309 & ~x321 & ~x323;
assign c0188 =  x103 &  x267 &  x285 &  x312;
assign c0190 =  x21 &  x142 &  x241 &  x250 & ~x300;
assign c0192 =  x188 &  x231 &  x277;
assign c0194 =  x71 &  x313 & ~x138 & ~x191;
assign c0196 =  x186 &  x242 &  x276 &  x303;
assign c0198 = ~x35 & ~x44 & ~x89 & ~x108;
assign c0200 =  x264 &  x321 & ~x109 & ~x118;
assign c0202 =  x122 & ~x201 & ~x317 & ~x323;
assign c0204 =  x101 &  x122 &  x134;
assign c0206 =  x96 &  x200 &  x253 &  x258 &  x271 & ~x247;
assign c0208 =  x214 & ~x154 & ~x230 & ~x289;
assign c0210 =  x102 &  x238;
assign c0212 =  x25 &  x187 &  x321 & ~x81;
assign c0214 =  x195 &  x268 &  x294;
assign c0216 =  x64 &  x321 & ~x306;
assign c0218 =  x166 & ~x46 & ~x174 & ~x233;
assign c0220 =  x123 &  x315 &  x316;
assign c0222 =  x162 &  x285 &  x312 & ~x318;
assign c0224 = ~x107 & ~x192 & ~x268 & ~x300 & ~x319 & ~x321;
assign c0226 =  x95 &  x131 & ~x263;
assign c0228 =  x33 &  x102 &  x276 &  x316;
assign c0230 =  x249 &  x289 & ~x291 & ~x322;
assign c0232 =  x92 &  x254 & ~x88;
assign c0234 =  x236 &  x300 & ~x149 & ~x261;
assign c0236 =  x267 & ~x39 & ~x48 & ~x122;
assign c0238 =  x68 &  x257 & ~x66 & ~x290 & ~x318;
assign c0240 =  x114 &  x140 & ~x35 & ~x44 & ~x171;
assign c0242 =  x240 & ~x20 & ~x119 & ~x140;
assign c0244 = ~x96 & ~x103 & ~x105 & ~x262;
assign c0246 =  x116 &  x121 &  x132 & ~x115;
assign c0248 =  x137 &  x240 & ~x145;
assign c0250 = ~x96 & ~x105 & ~x154 & ~x224 & ~x269;
assign c0252 = ~x34 & ~x157 & ~x168 & ~x269 & ~x293;
assign c0254 =  x103 &  x105 &  x106 &  x132 &  x294;
assign c0256 =  x77 & ~x291 & ~x309 & ~x321;
assign c0258 =  x56 &  x106 &  x128 &  x267;
assign c0260 =  x262 & ~x164 & ~x166 & ~x223;
assign c0262 =  x123 & ~x129 & ~x304;
assign c0264 =  x150 &  x240 &  x263 & ~x111;
assign c0266 =  x86 &  x297 & ~x9 & ~x67;
assign c0268 =  x226 & ~x85 & ~x129 & ~x228 & ~x263;
assign c0270 =  x7 & ~x123 & ~x251;
assign c0272 =  x322 & ~x5 & ~x28 & ~x307;
assign c0274 =  x307 & ~x138 & ~x323;
assign c0276 =  x92 &  x169 &  x213 &  x292 & ~x284;
assign c0278 =  x18 &  x168 &  x186;
assign c0280 =  x25 &  x187 & ~x23 & ~x105;
assign c0282 =  x22 & ~x118;
assign c0284 = ~x217 & ~x224 & ~x248;
assign c0286 =  x37 & ~x240 & ~x292 & ~x296;
assign c0288 =  x223 &  x285 & ~x271;
assign c0290 =  x226 &  x253 & ~x51;
assign c0292 = ~x169 & ~x260 & ~x279;
assign c0294 =  x24 &  x241 &  x312 & ~x136 & ~x172;
assign c0296 =  x234 & ~x4 & ~x17;
assign c0298 =  x240 & ~x8 & ~x34 & ~x99;
assign c0300 =  x96 &  x213 &  x315;
assign c0302 =  x184 &  x310;
assign c0304 =  x243 & ~x58 & ~x219 & ~x220 & ~x236;
assign c0306 =  x199 & ~x1 & ~x134;
assign c0308 =  x262 & ~x129 & ~x318;
assign c0310 =  x49 & ~x32 & ~x38 & ~x311;
assign c0312 =  x11 & ~x174 & ~x291;
assign c0314 =  x185 &  x306 & ~x160 & ~x320;
assign c0316 = ~x80 & ~x150 & ~x301;
assign c0318 =  x194 & ~x134 & ~x191 & ~x288 & ~x316;
assign c0320 = ~x24 & ~x128 & ~x267 & ~x268;
assign c0322 =  x184 &  x285 &  x312 & ~x230;
assign c0324 =  x154 &  x312;
assign c0326 =  x121 &  x317 & ~x3 & ~x280;
assign c0328 =  x102 &  x321 & ~x68 & ~x203 & ~x262;
assign c0330 =  x168 &  x311 & ~x246;
assign c0332 =  x154 & ~x138 & ~x228 & ~x237;
assign c0334 =  x123 &  x159 &  x312 & ~x21 & ~x115;
assign c0336 =  x178 & ~x0 & ~x27 & ~x150;
assign c0338 =  x151 &  x187 & ~x18 & ~x100 & ~x127;
assign c0340 =  x24 &  x56 &  x245 & ~x174;
assign c0342 =  x43 & ~x134 & ~x261 & ~x268 & ~x300;
assign c0344 =  x11 &  x200 & ~x287;
assign c0346 =  x38 &  x42 &  x101 &  x105;
assign c0348 =  x130 & ~x219;
assign c0350 =  x18 &  x159 &  x240 & ~x194;
assign c0352 =  x24 &  x101 &  x144;
assign c0354 = ~x128 & ~x269 & ~x315 & ~x316 & ~x321;
assign c0356 =  x25 & ~x255;
assign c0358 = ~x4 & ~x14 & ~x101 & ~x167 & ~x224;
assign c0360 =  x64 & ~x160 & ~x278;
assign c0362 =  x146 &  x208 & ~x130 & ~x189 & ~x264;
assign c0364 =  x18 & ~x157 & ~x316;
assign c0366 =  x105 &  x166 & ~x93 & ~x250;
assign c0368 = ~x6 & ~x9 & ~x212 & ~x217;
assign c0370 =  x241 &  x295 & ~x31 & ~x222;
assign c0372 =  x106 &  x209 & ~x5 & ~x75;
assign c0374 =  x160 &  x315;
assign c0376 =  x49 &  x110;
assign c0378 = ~x76 & ~x159 & ~x245;
assign c0380 =  x71 &  x80 &  x143 &  x160 &  x215 & ~x220;
assign c0382 =  x26 &  x102 & ~x99 & ~x318;
assign c0384 =  x96 &  x166 & ~x113;
assign c0386 = ~x14 & ~x22 & ~x157 & ~x314;
assign c0388 =  x203 & ~x0 & ~x164 & ~x223;
assign c0390 =  x33 &  x114 &  x240 &  x314;
assign c0392 = ~x8 & ~x205;
assign c0394 = ~x67 & ~x94 & ~x154 & ~x256 & ~x316;
assign c0396 =  x24 &  x47 &  x51 & ~x217;
assign c0398 =  x283 &  x316;
assign c0400 =  x107 & ~x144 & ~x148 & ~x286;
assign c0402 =  x6 & ~x99 & ~x105;
assign c0404 =  x47 &  x74 &  x182 &  x236 &  x308 &  x312;
assign c0406 = ~x1 & ~x5 & ~x101 & ~x128 & ~x263 & ~x316;
assign c0408 =  x183 & ~x33 & ~x167 & ~x195;
assign c0410 =  x20 &  x80 & ~x217;
assign c0412 =  x137 &  x294 & ~x86 & ~x275;
assign c0414 =  x49 &  x215 &  x290;
assign c0416 =  x256 & ~x217;
assign c0418 =  x5 &  x94 &  x101 & ~x203;
assign c0420 =  x52 &  x84 & ~x103 & ~x253;
assign c0422 =  x96 &  x101 &  x123 & ~x30;
assign c0424 =  x46 &  x243 & ~x4 & ~x205 & ~x256;
assign c0426 =  x106 & ~x115 & ~x255 & ~x277;
assign c0428 =  x63 &  x290 & ~x64;
assign c0430 =  x5 &  x211 &  x293;
assign c0432 =  x22 &  x102 & ~x297;
assign c0434 =  x24 &  x74 & ~x126 & ~x304;
assign c0436 =  x56 &  x163 &  x191 &  x224;
assign c0438 =  x294 &  x323 & ~x84;
assign c0440 =  x239 & ~x277 & ~x319;
assign c0442 =  x43 &  x52 & ~x132 & ~x288;
assign c0444 =  x40 &  x184 & ~x54;
assign c0446 =  x315 &  x321 & ~x177;
assign c0448 =  x173 & ~x99 & ~x126 & ~x153 & ~x233;
assign c0450 =  x15 &  x114 &  x128 &  x249 &  x276 &  x303;
assign c0452 =  x25 & ~x100 & ~x131 & ~x224;
assign c0454 =  x262 &  x266 &  x297;
assign c0456 =  x60 &  x71 &  x155 &  x316;
assign c0458 =  x152 & ~x152 & ~x211;
assign c0460 =  x69 &  x222 & ~x300;
assign c0462 = ~x0 & ~x18 & ~x125 & ~x162 & ~x220 & ~x252;
assign c0464 =  x69 &  x314 &  x321 & ~x271;
assign c0466 =  x106 &  x267 &  x315;
assign c0468 = ~x18 & ~x24 & ~x46 & ~x131 & ~x262;
assign c0470 = ~x163 & ~x167 & ~x319 & ~x321;
assign c0472 = ~x33 & ~x83 & ~x195 & ~x224 & ~x227;
assign c0474 =  x20 &  x75 & ~x125 & ~x260 & ~x266;
assign c0476 = ~x36 & ~x126 & ~x199;
assign c0478 =  x151 & ~x103 & ~x105 & ~x127 & ~x154;
assign c0480 = ~x4 & ~x128 & ~x161 & ~x314;
assign c0482 =  x15 &  x40 &  x316;
assign c0484 =  x47 & ~x68 & ~x201 & ~x248;
assign c0486 =  x102 & ~x3 & ~x230;
assign c0488 =  x66 &  x96 &  x119 &  x123 & ~x192;
assign c0490 =  x16 &  x214 & ~x19 & ~x103 & ~x127;
assign c0492 =  x93 & ~x280;
assign c0494 = ~x134 & ~x167 & ~x207 & ~x256 & ~x260;
assign c0496 =  x23 &  x226 & ~x211;
assign c0498 =  x141 & ~x296 & ~x318 & ~x319;
assign c0500 =  x55 & ~x119 & ~x288;
assign c0502 =  x132 &  x261 & ~x167;
assign c0504 = ~x0 & ~x6 & ~x60 & ~x163 & ~x220 & ~x221;
assign c0506 =  x118 & ~x94 & ~x148 & ~x315;
assign c0508 =  x221 & ~x92 & ~x133;
assign c0510 =  x177 &  x312 & ~x199 & ~x226;
assign c0512 =  x72 &  x128 &  x148;
assign c0514 =  x40 &  x87 &  x283 & ~x3;
assign c0516 =  x94 & ~x140 & ~x237;
assign c0518 =  x80 &  x184 &  x269;
assign c0520 =  x24 &  x101 &  x292 & ~x8;
assign c0522 =  x111 &  x238 & ~x284;
assign c0524 =  x294 & ~x140 & ~x309;
assign c0526 = ~x77 & ~x113 & ~x279 & ~x287;
assign c0528 =  x67 &  x241 &  x258;
assign c0530 =  x148 &  x202 &  x215 &  x320;
assign c0532 =  x262 & ~x138 & ~x192 & ~x223;
assign c0534 =  x218 & ~x48 & ~x142;
assign c0536 =  x21 & ~x8 & ~x219 & ~x228 & ~x300;
assign c0538 =  x80 &  x158 & ~x48;
assign c0540 =  x20 &  x184 & ~x3;
assign c0542 =  x15 &  x94 &  x158;
assign c0544 =  x128 & ~x48 & ~x251;
assign c0546 =  x24 &  x51 &  x95 &  x213 &  x303 &  x312;
assign c0548 = ~x105 & ~x150 & ~x163 & ~x224;
assign c0550 =  x158 &  x160 & ~x212;
assign c0552 =  x194 & ~x160 & ~x296 & ~x319 & ~x322;
assign c0554 =  x99 & ~x228 & ~x301;
assign c0556 = ~x37 & ~x81 & ~x137 & ~x192 & ~x301;
assign c0558 =  x289 & ~x39 & ~x203 & ~x248;
assign c0560 =  x315 & ~x305;
assign c0562 =  x152 &  x206 &  x245 &  x260 & ~x3;
assign c0564 =  x11 &  x52 & ~x297;
assign c0566 = ~x146 & ~x151 & ~x160 & ~x241 & ~x290 & ~x300 & ~x313 & ~x317;
assign c0568 =  x97 &  x263 &  x312 & ~x117;
assign c0570 =  x148 &  x289 &  x312;
assign c0572 =  x200 & ~x135 & ~x291 & ~x318;
assign c0574 =  x7 &  x12 &  x291 & ~x307;
assign c0576 = ~x31 & ~x56 & ~x222 & ~x269 & ~x294;
assign c0578 =  x13 & ~x255;
assign c0580 =  x250 & ~x106 & ~x132 & ~x134 & ~x154 & ~x294;
assign c0582 =  x21 & ~x130 & ~x262;
assign c0584 =  x97 & ~x99 & ~x313;
assign c0586 =  x128 &  x263 & ~x30 & ~x271;
assign c0588 =  x24 &  x76 &  x312;
assign c0590 =  x307 &  x311 & ~x318 & ~x319;
assign c0592 =  x132 & ~x156 & ~x210;
assign c0594 =  x173 & ~x219 & ~x306 & ~x316;
assign c0596 =  x43 &  x209 & ~x18 & ~x311;
assign c0598 =  x159 &  x200 &  x245 & ~x210;
assign c01 =  x297 & ~x231 & ~x240 & ~x241 & ~x303 & ~x312 & ~x313;
assign c03 =  x107 &  x264 &  x284;
assign c05 =  x154 &  x155 &  x212 &  x284 &  x289 &  x290 &  x316;
assign c07 =  x90 &  x228 &  x300 & ~x281;
assign c09 =  x269 & ~x186 & ~x258 & ~x263;
assign c011 =  x63 &  x147 &  x282 &  x283;
assign c013 =  x1 &  x2 &  x147 &  x217;
assign c015 =  x108 & ~x47 & ~x74 & ~x146 & ~x182 & ~x183 & ~x209;
assign c017 =  x71 &  x138 &  x205 &  x206 &  x273 &  x278;
assign c019 =  x146 &  x209 &  x280 &  x281 & ~x90 & ~x292;
assign c021 =  x237 &  x238 &  x309 &  x310 & ~x42 & ~x177;
assign c023 =  x70 &  x142 &  x278 & ~x271 & ~x297;
assign c025 =  x66 &  x111 &  x201 &  x266 &  x273;
assign c027 =  x199 &  x240 &  x291;
assign c029 =  x221 &  x292 & ~x278;
assign c031 =  x1 &  x192 & ~x168 & ~x195;
assign c033 =  x32 &  x63 &  x135 &  x167 &  x198 &  x224;
assign c035 =  x28 & ~x158 & ~x311;
assign c037 =  x254 & ~x40 & ~x112 & ~x121 & ~x319;
assign c039 =  x47 &  x182 & ~x122 & ~x294;
assign c041 =  x70 &  x183 &  x187 &  x277 & ~x64;
assign c043 =  x5 &  x12 &  x84 &  x181;
assign c045 = ~x159 & ~x233 & ~x234 & ~x294 & ~x297 & ~x305;
assign c047 =  x18 &  x55 &  x90 &  x190 & ~x196;
assign c049 =  x144 &  x299 & ~x316;
assign c051 =  x36 &  x108 &  x171 &  x243 &  x251 & ~x195;
assign c053 =  x43 & ~x92 & ~x271 & ~x272;
assign c055 =  x1 &  x2 &  x29 & ~x97;
assign c057 =  x162 & ~x67 & ~x68 & ~x76 & ~x139 & ~x140 & ~x148;
assign c059 =  x140 & ~x43 & ~x250 & ~x261;
assign c061 =  x167 &  x183 & ~x50 & ~x185;
assign c063 = ~x18 & ~x46 & ~x90 & ~x181 & ~x209 & ~x281;
assign c065 =  x75 &  x282 &  x283 & ~x42;
assign c067 =  x5 &  x12 &  x13 & ~x58 & ~x193;
assign c069 =  x50 & ~x44 & ~x126 & ~x179 & ~x261;
assign c071 =  x48 &  x120 &  x183 &  x205 &  x255 & ~x198 & ~x270;
assign c073 =  x84 & ~x67 & ~x148 & ~x202 & ~x203;
assign c075 =  x77 &  x130 &  x212 &  x230 &  x302;
assign c077 =  x287 & ~x155 & ~x289 & ~x290 & ~x316;
assign c079 =  x35 &  x44 &  x162 &  x170 &  x194;
assign c081 =  x262 &  x263 &  x289 & ~x276;
assign c083 =  x117 & ~x78 & ~x150 & ~x213 & ~x214 & ~x285;
assign c085 =  x66 &  x151 &  x202 &  x273 &  x274;
assign c087 =  x9 &  x17 &  x26 & ~x69;
assign c089 =  x147 &  x234 &  x306 & ~x260;
assign c091 =  x108 &  x109 &  x244 & ~x67 & ~x68;
assign c093 =  x122 &  x248 &  x257 & ~x235 & ~x298;
assign c095 =  x23 &  x95 & ~x39 & ~x111 & ~x174 & ~x200 & ~x246 & ~x272;
assign c097 = ~x155 & ~x238 & ~x290 & ~x302 & ~x316;
assign c099 =  x195 & ~x79 & ~x258 & ~x259;
assign c0101 =  x156 &  x217 &  x225 &  x297;
assign c0103 =  x0 &  x1 &  x26 &  x99;
assign c0105 =  x10 &  x20 &  x92 &  x279;
assign c0107 =  x237 &  x309 &  x319 & ~x72 & ~x207;
assign c0109 =  x219 & ~x58;
assign c0111 =  x55 &  x56 &  x190 &  x191 &  x218 &  x309;
assign c0113 =  x27 &  x116 &  x162 & ~x61;
assign c0115 = ~x228 & ~x229 & ~x273 & ~x297 & ~x301;
assign c0117 =  x259 & ~x233 & ~x242 & ~x305 & ~x306 & ~x314 & ~x315;
assign c0119 =  x79 &  x151 &  x152 &  x286 & ~x20 & ~x92;
assign c0121 =  x7 &  x232 &  x304 & ~x192;
assign c0123 =  x5 &  x73 &  x85 &  x145 &  x208;
assign c0125 =  x127 &  x128 & ~x15 & ~x87;
assign c0127 =  x33 &  x60 &  x194 &  x195 & ~x139;
assign c0129 =  x240 &  x312 &  x313 & ~x229 & ~x238 & ~x301 & ~x310;
assign c0131 =  x37 &  x109 &  x172 &  x243 &  x244 &  x268;
assign c0133 =  x178 &  x249 &  x250 & ~x37 & ~x64 & ~x109;
assign c0135 =  x37 &  x65 &  x109 &  x259 & ~x5;
assign c0137 =  x74 &  x75 &  x146 &  x147 &  x209 &  x282 &  x305;
assign c0139 =  x143 &  x168 & ~x234 & ~x306 & ~x315;
assign c0141 =  x238 &  x310 & ~x127 & ~x128 & ~x262 & ~x263;
assign c0143 =  x0 &  x1 &  x17 & ~x143;
assign c0145 =  x34 &  x61 &  x169 &  x195 & ~x220;
assign c0147 = ~x96 & ~x173 & ~x174 & ~x246;
assign c0149 =  x10 &  x82 &  x322 & ~x44;
assign c0151 =  x119 &  x145 &  x146 & ~x108 & ~x243;
assign c0153 =  x242 &  x314 & ~x54 & ~x189 & ~x312;
assign c0155 =  x66 &  x100 &  x101 &  x138 &  x273;
assign c0157 =  x209 &  x281 & ~x52 & ~x149 & ~x284;
assign c0159 =  x41 & ~x10 & ~x231;
assign c0161 =  x226 &  x234 &  x306 & ~x173;
assign c0163 =  x42 &  x68 &  x140 &  x160;
assign c0165 =  x64 &  x135 &  x161 &  x198 &  x199;
assign c0167 =  x64 &  x68 &  x140 &  x275 &  x285;
assign c0169 =  x64 &  x109 &  x110 &  x136 & ~x239;
assign c0171 =  x68 &  x279 & ~x37 & ~x38 & ~x173;
assign c0173 = ~x67 & ~x69 & ~x140 & ~x203 & ~x276;
assign c0175 =  x157 &  x292 & ~x145 & ~x285;
assign c0177 =  x278 & ~x3 & ~x12 & ~x13 & ~x84;
assign c0179 =  x220 &  x221 &  x230 &  x279;
assign c0181 =  x127 &  x153 &  x154 &  x262 &  x288 &  x315;
assign c0183 =  x43 &  x52 &  x115 &  x187 &  x250 &  x261;
assign c0185 =  x48 &  x49 &  x120 &  x156 &  x183 &  x255 &  x264;
assign c0187 =  x23 &  x95 &  x216 &  x288;
assign c0189 = ~x133 & ~x151 & ~x217 & ~x286;
assign c0191 =  x38 &  x110 &  x173 &  x245 & ~x238 & ~x310 & ~x319;
assign c0193 = ~x47 & ~x48 & ~x119 & ~x120 & ~x146 & ~x182 & ~x183 & ~x209 & ~x254 & ~x255;
assign c0195 =  x70 &  x205 &  x277 & ~x199 & ~x227 & ~x298 & ~x299;
assign c0197 = ~x51 & ~x132 & ~x267 & ~x294 & ~x322;
assign c0199 =  x268 & ~x232 & ~x237 & ~x304;
assign c0201 =  x174 &  x246 &  x286 &  x314;
assign c0203 =  x43 &  x68 &  x100 &  x101 &  x115 &  x178 &  x250;
assign c0205 =  x46 &  x47 &  x118 &  x207 & ~x35;
assign c0207 =  x77 &  x129 &  x149 &  x212 &  x264 &  x284 &  x285;
assign c0209 =  x228 &  x300 & ~x71 & ~x179 & ~x206;
assign c0211 =  x93 &  x217 &  x288;
assign c0213 =  x219 & ~x157 & ~x222;
assign c0215 =  x75 &  x147 & ~x114 & ~x243;
assign c0217 =  x49 &  x121 & ~x26 & ~x52 & ~x98 & ~x124 & ~x259;
assign c0219 =  x219 &  x228 &  x238 &  x239 &  x301 &  x311;
assign c0221 = ~x17 & ~x27 & ~x30 & ~x62 & ~x171;
assign c0223 = ~x33 & ~x44 & ~x179 & ~x237;
assign c0225 =  x154 &  x291 & ~x108 & ~x243;
assign c0227 =  x49 &  x121 &  x122 &  x256 & ~x260;
assign c0229 =  x312 & ~x182 & ~x289;
assign c0231 =  x73 &  x145 &  x207 &  x280 & ~x242 & ~x314;
assign c0233 =  x154 &  x155 & ~x45 & ~x46 & ~x181;
assign c0235 = ~x18 & ~x216 & ~x224 & ~x225 & ~x226 & ~x297;
assign c0237 =  x216 & ~x145 & ~x236 & ~x308;
assign c0239 =  x27 &  x30 &  x31 &  x39 &  x174;
assign c0241 =  x172 &  x244 &  x252 & ~x204;
assign c0243 =  x218 & ~x9 & ~x26 & ~x81 & ~x89 & ~x98;
assign c0245 =  x232 & ~x226 & ~x317;
assign c0247 =  x241 &  x313 & ~x317;
assign c0249 =  x1 &  x57 &  x91 &  x192;
assign c0251 =  x12 &  x13 &  x84 &  x85 &  x111 & ~x51;
assign c0253 =  x63 &  x135 &  x198 &  x207 &  x270 &  x279 & ~x315;
assign c0255 =  x71 &  x143 &  x178 &  x277 &  x278 & ~x36;
assign c0257 =  x44 &  x179 & ~x96 & ~x303;
assign c0259 =  x5 &  x13 &  x21 &  x48 &  x120;
assign c0261 = ~x13 & ~x21 & ~x48 & ~x85 & ~x161;
assign c0263 =  x6 &  x118 &  x253 & ~x67 & ~x202;
assign c0265 =  x318 & ~x61 & ~x321 & ~x322;
assign c0267 =  x269 & ~x101 & ~x147;
assign c0269 =  x171 &  x243 &  x286 & ~x236;
assign c0271 =  x142 &  x178 &  x214 &  x250 & ~x110 & ~x173;
assign c0273 = ~x16 & ~x50 & ~x51 & ~x288;
assign c0275 =  x224 &  x233 &  x234 &  x305 &  x306 & ~x163;
assign c0277 =  x139 &  x174 &  x246 &  x247 & ~x22 & ~x94;
assign c0279 =  x232 &  x304 & ~x111 & ~x175 & ~x247;
assign c0281 =  x9 &  x18 &  x81 &  x90 &  x98 &  x99;
assign c0283 =  x51 &  x258 & ~x128 & ~x311;
assign c0285 =  x248 &  x249 &  x253 &  x294;
assign c0287 =  x48 &  x120 &  x309 &  x319;
assign c0289 =  x66 &  x139 &  x202 &  x273 &  x274 & ~x240;
assign c0291 =  x146 &  x209 &  x226 &  x235 &  x280 &  x281 &  x298 &  x307;
assign c0293 =  x238 &  x310 &  x319 & ~x175 & ~x176 & ~x248;
assign c0295 =  x64 &  x65 &  x135 &  x137 &  x270 &  x271;
assign c0297 =  x125 &  x188 &  x260 &  x310 &  x318;
assign c0299 =  x291 & ~x83 & ~x96;
assign c0301 = ~x20 & ~x128 & ~x154 & ~x155 & ~x262 & ~x263;
assign c0303 =  x135 & ~x127 & ~x128 & ~x155 & ~x262 & ~x263 & ~x290;
assign c0305 =  x14 & ~x88 & ~x161;
assign c0307 =  x156 & ~x98 & ~x102 & ~x216;
assign c0309 =  x34 &  x232 &  x304 &  x319;
assign c0311 =  x170 & ~x42 & ~x69 & ~x177 & ~x213;
assign c0313 =  x77 &  x149 &  x158 &  x212 &  x265 &  x266 &  x284 & ~x182;
assign c0315 =  x194 &  x223 &  x270;
assign c0317 =  x321 & ~x21 & ~x22 & ~x85 & ~x93 & ~x102;
assign c0319 =  x62 &  x197 & ~x231 & ~x303;
assign c0321 =  x60 &  x127 &  x155 &  x272;
assign c0323 =  x153 &  x207 &  x218 &  x279 &  x288;
assign c0325 =  x196 &  x237 &  x309 &  x319;
assign c0327 =  x151 &  x204 & ~x216 & ~x274;
assign c0329 =  x141 &  x242 &  x276 &  x318;
assign c0331 =  x45 &  x86 & ~x79 & ~x214;
assign c0333 =  x63 &  x143 & ~x209 & ~x282;
assign c0335 =  x91 &  x110 &  x245 & ~x213;
assign c0337 =  x53 & ~x49 & ~x50 & ~x122 & ~x185;
assign c0339 =  x42 &  x86 &  x207 & ~x4 & ~x35;
assign c0341 =  x249 &  x271 & ~x27 & ~x116 & ~x179 & ~x251;
assign c0343 =  x43 &  x48 &  x49 &  x115 &  x120 &  x250 &  x255;
assign c0345 =  x212 &  x264 &  x297;
assign c0347 =  x130 &  x153 &  x219 &  x288;
assign c0349 =  x114 &  x115 &  x186 &  x249 &  x250 & ~x171;
assign c0351 =  x55 &  x219 & ~x61;
assign c0353 =  x60 &  x288 & ~x172;
assign c0355 =  x284 &  x313 & ~x177;
assign c0357 =  x233 &  x234 &  x305 &  x306 & ~x31 & ~x166;
assign c0359 =  x203 & ~x45 & ~x180 & ~x188 & ~x252 & ~x260;
assign c0361 = ~x29 & ~x100 & ~x165 & ~x217;
assign c0363 =  x122 &  x130 &  x131 &  x185 &  x257 &  x266 & ~x119;
assign c0365 =  x115 &  x116 & ~x135;
assign c0367 =  x219 &  x220 &  x229 &  x230 &  x302;
assign c0369 =  x259 &  x288 & ~x31;
assign c0371 =  x93 & ~x87 & ~x88;
assign c0373 = ~x42 & ~x157 & ~x240;
assign c0375 =  x48 &  x120 &  x240 &  x255 & ~x202 & ~x274;
assign c0377 =  x294 &  x322 & ~x155;
assign c0379 =  x5 &  x21 &  x84 &  x93 & ~x287;
assign c0381 =  x54 &  x189 &  x298 &  x322;
assign c0383 =  x128 &  x155 &  x263 &  x290 & ~x319;
assign c0385 =  x39 &  x40 &  x111 &  x112 &  x174 &  x175 &  x246 &  x247 & ~x19;
assign c0387 =  x107 &  x129 &  x189 &  x264;
assign c0389 =  x155 &  x290 & ~x161 & ~x200 & ~x296;
assign c0391 =  x238 &  x239 &  x310 &  x311 &  x318 &  x319;
assign c0393 =  x29 &  x146 &  x164 &  x281 &  x307;
assign c0395 =  x156 &  x205 & ~x137 & ~x199 & ~x271 & ~x300;
assign c0397 =  x53 &  x81 &  x125 & ~x42;
assign c0399 =  x102 &  x262 & ~x96;
assign c0401 =  x165 &  x228 &  x238 &  x301 & ~x69 & ~x204;
assign c0403 =  x242 &  x314 & ~x59 & ~x189 & ~x198;
assign c0405 =  x13 &  x85 & ~x19 & ~x91 & ~x227 & ~x299;
assign c0407 =  x113 &  x176 & ~x230 & ~x301;
assign c0409 =  x296 & ~x154 & ~x242 & ~x314;
assign c0411 =  x53 &  x77 &  x125 &  x149 &  x212 &  x260 &  x284;
assign c0413 =  x67 &  x68 &  x140 &  x203 &  x275 &  x291;
assign c0415 =  x319 & ~x42 & ~x270;
assign c0417 = ~x43 & ~x115 & ~x132 & ~x250 & ~x267;
assign c0419 = ~x195 & ~x223 & ~x224 & ~x275 & ~x297;
assign c0421 =  x108 &  x125 &  x136 &  x271;
assign c0423 =  x61 & ~x11 & ~x83 & ~x237 & ~x309;
assign c0425 = ~x240 & ~x248 & ~x303 & ~x312;
assign c0427 =  x41 &  x49 &  x121 & ~x29 & ~x200 & ~x245;
assign c0429 =  x158 &  x293 & ~x72 & ~x144 & ~x271;
assign c0431 =  x52 &  x124 &  x213 &  x275 &  x285;
assign c0433 =  x127 &  x145 &  x154 &  x155 & ~x260;
assign c0435 =  x320 & ~x65 & ~x110;
assign c0437 =  x286 & ~x307 & ~x308 & ~x316;
assign c0439 =  x118 & ~x122 & ~x257 & ~x258;
assign c0441 =  x28 &  x55 &  x190 &  x191 &  x218 &  x322;
assign c0443 =  x14 &  x52 &  x86 &  x222;
assign c0445 =  x40 &  x112 &  x175 &  x176 &  x247 &  x248 & ~x21 & ~x93;
assign c0447 =  x132 &  x159 &  x294 &  x322 & ~x49 & ~x121 & ~x184 & ~x256;
assign c0449 =  x100 &  x114 &  x115 &  x249 &  x250;
assign c0451 =  x70 &  x112 &  x142 &  x178 &  x179 &  x277;
assign c0453 =  x17 &  x26 &  x29 &  x81 &  x89 &  x98 &  x164;
assign c0455 =  x233 &  x234 &  x288 & ~x245;
assign c0457 =  x69 &  x141 &  x276 &  x291 & ~x272;
assign c0459 =  x75 &  x111 &  x138 &  x174 &  x210 &  x245 &  x273 &  x282;
assign c0461 = ~x7 & ~x10 & ~x18 & ~x19 & ~x82 & ~x90 & ~x91;
assign c0463 =  x84 &  x131 &  x159 &  x266 &  x294;
assign c0465 =  x39 &  x40 &  x48 &  x49 &  x111 &  x112 &  x183;
assign c0467 =  x32 &  x36 &  x77 &  x108 &  x171;
assign c0469 =  x29 &  x164 &  x285 & ~x33 & ~x168;
assign c0471 =  x259 & ~x4 & ~x13 & ~x21;
assign c0473 =  x82 &  x211 & ~x197;
assign c0475 =  x211 &  x273 &  x283 & ~x141 & ~x249;
assign c0477 = ~x16 & ~x88 & ~x231 & ~x303 & ~x319;
assign c0479 =  x77 &  x149 &  x212 &  x284 & ~x167 & ~x206;
assign c0481 =  x82 &  x142 &  x277 & ~x45;
assign c0483 =  x79 &  x105 &  x120 &  x214;
assign c0485 =  x192 &  x247 & ~x20;
assign c0487 =  x3 &  x29 &  x55 &  x56 &  x164 &  x165 &  x190;
assign c0489 =  x42 &  x144 &  x176 &  x177 &  x207 &  x248 &  x249 &  x279;
assign c0491 =  x71 &  x143 &  x206 &  x278 & ~x263 & ~x316;
assign c0493 =  x67 &  x139 &  x140 & ~x44 & ~x179;
assign c0495 =  x36 &  x37 & ~x173;
assign c0497 = ~x105 & ~x222 & ~x276;
assign c0499 = ~x33 & ~x168 & ~x177 & ~x178 & ~x195;
assign c0501 =  x29 &  x165 & ~x68 & ~x69 & ~x203;
assign c0503 =  x180 &  x252 &  x253 & ~x19;
assign c0505 = ~x78 & ~x141 & ~x142 & ~x204 & ~x205 & ~x277;
assign c0507 = ~x78 & ~x150 & ~x151 & ~x212 & ~x213 & ~x285 & ~x286;
assign c0509 =  x129 &  x234 &  x264 &  x280;
assign c0511 =  x126 & ~x67 & ~x76 & ~x148 & ~x202 & ~x274;
assign c0513 =  x132 &  x133 &  x267 &  x268 &  x295 &  x302;
assign c0515 =  x193 & ~x21 & ~x323;
assign c0517 =  x128 &  x254 &  x263 & ~x242 & ~x314;
assign c0519 = ~x79 & ~x188 & ~x214;
assign c0521 =  x81 & ~x47 & ~x118 & ~x181 & ~x182 & ~x253;
assign c0523 =  x45 &  x95 & ~x17 & ~x89;
assign c0525 =  x158 &  x228 & ~x215;
assign c0527 =  x73 &  x145 &  x207 &  x208 &  x279 & ~x238 & ~x301 & ~x310;
assign c0529 =  x29 &  x191 & ~x33 & ~x168;
assign c0531 =  x64 &  x125 & ~x94;
assign c0533 = ~x21 & ~x48 & ~x93 & ~x105;
assign c0535 =  x59 &  x86 &  x194 &  x224 &  x225 &  x297;
assign c0537 =  x267 &  x295 & ~x157 & ~x211 & ~x283 & ~x292;
assign c0539 =  x41 &  x42 &  x113 &  x176 & ~x11 & ~x38 & ~x83 & ~x173;
assign c0541 =  x3 &  x51 & ~x272;
assign c0543 =  x3 &  x4 &  x233 &  x242 &  x305;
assign c0545 =  x42 &  x69 &  x114 &  x177 &  x207 &  x249 & ~x238;
assign c0547 =  x119 &  x145 &  x254 &  x264;
assign c0549 =  x46 &  x118 &  x181 &  x254 & ~x241 & ~x242;
assign c0551 =  x99 &  x264 & ~x116;
assign c0553 =  x265 & ~x224 & ~x234 & ~x306;
assign c0555 = ~x17 & ~x36 & ~x81 & ~x89 & ~x98 & ~x108 & ~x116 & ~x125;
assign c0557 =  x38 & ~x69 & ~x204 & ~x306;
assign c0559 =  x85 &  x94 & ~x25 & ~x97 & ~x123;
assign c0561 =  x156 &  x157 &  x292 & ~x321;
assign c0563 =  x69 &  x122 &  x140 &  x185 &  x204 &  x232;
assign c0565 =  x94 & ~x12 & ~x316;
assign c0567 =  x59 &  x194 &  x215 &  x287 & ~x284;
assign c0569 =  x224 & ~x29 & ~x231;
assign c0571 =  x93 &  x158 &  x293 &  x311 &  x320;
assign c0573 =  x48 &  x120 &  x154 &  x155 &  x183 &  x289;
assign c0575 =  x263 &  x289 &  x297 & ~x256;
assign c0577 = ~x144 & ~x207 & ~x225 & ~x234 & ~x297 & ~x307;
assign c0579 =  x262 & ~x76 & ~x98 & ~x148 & ~x157;
assign c0581 =  x3 &  x131 &  x217;
assign c0583 =  x17 &  x52 &  x89 &  x127;
assign c0585 =  x215 & ~x228 & ~x229 & ~x238 & ~x239 & ~x300 & ~x301 & ~x310 & ~x311;
assign c0587 =  x79 &  x214 &  x242 &  x286 &  x313 &  x314;
assign c0589 = ~x73 & ~x280 & ~x312;
assign c0591 =  x161 &  x296 &  x319 & ~x76;
assign c0593 =  x0 &  x73 &  x145 &  x208 &  x280 &  x307;
assign c0595 =  x0 &  x25 &  x97 &  x322;
assign c0597 =  x55 &  x68 &  x140 &  x190 &  x203 &  x275 &  x276;
assign c0599 =  x9 &  x29 &  x89 &  x200;
assign c10 =  x69 &  x141 &  x204 & ~x26 & ~x89 & ~x98 & ~x173;
assign c12 =  x18 &  x90 & ~x44 & ~x116 & ~x179 & ~x251;
assign c14 =  x194 &  x207 & ~x238;
assign c16 =  x66 &  x138 &  x201 &  x211 &  x273 &  x283 & ~x141;
assign c18 =  x5 &  x48 &  x120 & ~x257;
assign c110 =  x131 & ~x118 & ~x127 & ~x128 & ~x262 & ~x263;
assign c112 =  x41 &  x120 &  x183 & ~x102;
assign c114 =  x111 &  x120 &  x147 &  x148 &  x183 &  x255 &  x282;
assign c116 =  x237 &  x305 &  x309 &  x318;
assign c118 =  x48 &  x120 &  x315 &  x318;
assign c120 =  x118 &  x127 &  x165 &  x253;
assign c122 =  x242 &  x314 & ~x107 & ~x224;
assign c124 =  x28 &  x55 &  x163 &  x164 &  x190 &  x218 &  x322;
assign c126 =  x52 &  x53 &  x187 &  x188 &  x288;
assign c128 = ~x7 & ~x34 & ~x96 & ~x169;
assign c130 =  x72 &  x101 &  x207 & ~x310;
assign c132 =  x228 &  x229 &  x238 &  x301 &  x310 &  x311;
assign c134 =  x224 & ~x289 & ~x290 & ~x316;
assign c136 =  x252 & ~x50 & ~x122 & ~x150;
assign c138 =  x197 & ~x21 & ~x240;
assign c140 =  x36 &  x108 &  x167 &  x171 &  x172 &  x243;
assign c142 =  x105 &  x184 &  x256 & ~x102;
assign c144 =  x233 &  x305 &  x306 & ~x128;
assign c146 =  x30 &  x165 &  x315 & ~x72;
assign c148 = ~x10 & ~x28 & ~x29 & ~x56 & ~x92 & ~x164 & ~x191 & ~x217;
assign c150 =  x21 &  x34 &  x84 &  x93 & ~x192;
assign c152 =  x210 &  x282 & ~x207 & ~x213;
assign c154 =  x154 &  x290 & ~x90;
assign c156 = ~x43 & ~x44 & ~x115 & ~x178 & ~x238;
assign c158 =  x233 &  x305 & ~x51 & ~x227;
assign c160 =  x98 &  x107 &  x284 & ~x253;
assign c162 =  x17 &  x27 &  x89 & ~x22;
assign c164 =  x141 &  x249 &  x276 & ~x231;
assign c166 =  x178 &  x250 & ~x65 & ~x110 & ~x137 & ~x199 & ~x200;
assign c168 =  x234 &  x235 &  x306 &  x307 & ~x31 & ~x166;
assign c170 = ~x17 & ~x26 & ~x81 & ~x90 & ~x98 & ~x303;
assign c172 =  x66 &  x273 &  x274 &  x283 & ~x42;
assign c174 =  x75 &  x76 &  x111 &  x147 &  x183 &  x210 &  x282;
assign c176 =  x3 &  x4 &  x12 &  x84 &  x238;
assign c178 =  x45 &  x117 &  x118 &  x180 & ~x79 & ~x151;
assign c180 =  x64 &  x77 &  x212 &  x317;
assign c182 =  x30 &  x125 &  x165 & ~x42 & ~x69;
assign c184 =  x288 &  x306 &  x315 & ~x132;
assign c186 = ~x55 & ~x63 & ~x189 & ~x198 & ~x216 & ~x225 & ~x270;
assign c188 =  x241 &  x286 & ~x290;
assign c190 =  x275 &  x291 & ~x151 & ~x286;
assign c192 =  x242 &  x314 & ~x64 & ~x72 & ~x271;
assign c194 =  x29 &  x154 &  x174 &  x289;
assign c196 =  x95 &  x206 &  x207 &  x248 &  x278 &  x279;
assign c198 =  x167 & ~x23 & ~x301;
assign c1100 =  x3 &  x4 &  x21 &  x48 &  x93;
assign c1102 =  x50 &  x122 &  x175 &  x185 &  x248 &  x257 & ~x110;
assign c1104 =  x55 &  x302 & ~x247;
assign c1106 =  x9 &  x18 &  x81 &  x98 & ~x47 & ~x119;
assign c1108 = ~x115 & ~x178 & ~x186 & ~x187 & ~x250 & ~x258;
assign c1110 =  x66 &  x164 &  x201 &  x273 & ~x72 & ~x207;
assign c1112 =  x73 &  x145 &  x160 &  x185 &  x208 &  x280 &  x295;
assign c1114 =  x88 &  x161 &  x194;
assign c1116 =  x48 &  x120 &  x131 & ~x225;
assign c1118 =  x0 & ~x156 & ~x157 & ~x283;
assign c1120 = ~x147 & ~x234 & ~x235 & ~x297 & ~x307;
assign c1122 =  x124 &  x212 & ~x13 & ~x84 & ~x85;
assign c1124 =  x129 &  x155 &  x156 &  x264 &  x289 &  x290 &  x291;
assign c1126 =  x162 &  x214 & ~x67 & ~x76;
assign c1128 =  x127 &  x128 &  x154 &  x263 &  x289 & ~x312;
assign c1130 =  x274 & ~x146 & ~x183 & ~x209 & ~x255;
assign c1132 =  x229 &  x301 & ~x168 & ~x241;
assign c1134 =  x200 & ~x168 & ~x203;
assign c1136 =  x42 &  x177 & ~x21 & ~x26 & ~x93 & ~x98;
assign c1138 =  x49 &  x256 & ~x298 & ~x322;
assign c1140 =  x309 & ~x42 & ~x198 & ~x270;
assign c1142 =  x100 &  x142 & ~x13;
assign c1144 =  x73 &  x145 &  x154 &  x208 &  x280 &  x289 & ~x287;
assign c1146 =  x18 & ~x61 & ~x170 & ~x196;
assign c1148 =  x224 &  x225 &  x297 & ~x126 & ~x261;
assign c1150 =  x18 &  x90 &  x191 &  x300;
assign c1152 =  x86 &  x295 & ~x308;
assign c1154 =  x0 &  x9 &  x17 &  x81 &  x89 & ~x24;
assign c1156 =  x29 &  x100 &  x164 &  x217 &  x218;
assign c1158 =  x30 &  x101 &  x190;
assign c1160 =  x83 &  x255 & ~x26 & ~x102;
assign c1162 =  x43 &  x250 &  x261 & ~x147;
assign c1164 =  x71 &  x143 &  x206 &  x278 & ~x77 & ~x315;
assign c1166 =  x236 & ~x78 & ~x150 & ~x187 & ~x213 & ~x285;
assign c1168 =  x65 &  x272 & ~x24 & ~x25 & ~x96;
assign c1170 =  x7 &  x150 &  x285 &  x319;
assign c1172 =  x81 & ~x78 & ~x123 & ~x213;
assign c1174 =  x2 &  x51 &  x258 & ~x33;
assign c1176 =  x34 &  x169 &  x216 &  x217;
assign c1178 =  x1 & ~x177 & ~x247;
assign c1180 =  x68 &  x203 &  x223 &  x297 &  x306;
assign c1182 =  x45 &  x77 &  x108 &  x117 &  x149 &  x212 &  x284;
assign c1184 =  x156 &  x239 &  x302 & ~x252;
assign c1186 =  x3 &  x156 &  x240 &  x291;
assign c1188 =  x1 &  x86 &  x98;
assign c1190 = ~x172 & ~x240 & ~x312;
assign c1192 =  x14 &  x22 &  x86 & ~x80 & ~x152 & ~x215;
assign c1194 =  x168 &  x248 & ~x234 & ~x306;
assign c1196 =  x41 &  x143 &  x176 &  x278 & ~x11 & ~x83;
assign c1198 =  x60 &  x194 &  x198 &  x270 &  x271;
assign c1200 =  x51 &  x122 & ~x116 & ~x125 & ~x188 & ~x251 & ~x260;
assign c1202 = ~x78 & ~x79 & ~x211 & ~x212;
assign c1204 =  x181 &  x253 & ~x26 & ~x225;
assign c1206 =  x285 & ~x19 & ~x76 & ~x91 & ~x148;
assign c1208 =  x229 &  x302 &  x310 &  x311 &  x319;
assign c1210 =  x57 &  x192 &  x201 & ~x303;
assign c1212 = ~x6 & ~x7 & ~x237 & ~x238 & ~x300 & ~x309;
assign c1214 =  x52 &  x120 &  x128 &  x129 &  x264;
assign c1216 = ~x25 & ~x26 & ~x89 & ~x97 & ~x98 & ~x226;
assign c1218 = ~x47 & ~x193 & ~x216 & ~x225;
assign c1220 =  x54 &  x55 &  x189 &  x190 &  x199 &  x227;
assign c1222 =  x14 &  x284 & ~x287;
assign c1224 = ~x7 & ~x38 & ~x39 & ~x173 & ~x174 & ~x246;
assign c1226 =  x28 & ~x22 & ~x46;
assign c1228 =  x28 &  x219 & ~x148;
assign c1230 =  x314 & ~x23 & ~x102;
assign c1232 =  x8 &  x237 &  x238 &  x310 &  x319;
assign c1234 =  x13 &  x21 &  x93 & ~x152;
assign c1236 =  x57 &  x65 &  x147 &  x192;
assign c1238 =  x131 &  x266 &  x317 & ~x152;
assign c1240 =  x95 & ~x73 & ~x74 & ~x146 & ~x182 & ~x209 & ~x254 & ~x281;
assign c1242 =  x111 &  x158 & ~x145 & ~x280;
assign c1244 =  x23 &  x95 & ~x111 & ~x241;
assign c1246 =  x10 &  x19 & ~x242 & ~x314;
assign c1248 = ~x75 & ~x147 & ~x154 & ~x234 & ~x282;
assign c1250 =  x131 &  x158 &  x239 &  x284 &  x293 &  x311 &  x320;
assign c1252 =  x48 &  x49 &  x207 &  x255 &  x264;
assign c1254 =  x124 &  x132 &  x221 &  x267;
assign c1256 =  x107 &  x133 &  x134 &  x268 &  x284;
assign c1258 =  x227 &  x298 &  x299 & ~x238 & ~x310;
assign c1260 =  x9 &  x17 &  x26 &  x89 & ~x204;
assign c1262 =  x279 & ~x26 & ~x53 & ~x98 & ~x125;
assign c1264 = ~x46 & ~x207 & ~x224 & ~x225;
assign c1266 =  x76 &  x148 &  x211 &  x283 & ~x128 & ~x155 & ~x290;
assign c1268 =  x120 &  x183 & ~x87;
assign c1270 =  x30 &  x39 &  x40 &  x111 &  x165 &  x174 &  x175 &  x246;
assign c1272 =  x6 &  x34 &  x169 &  x196 &  x223 & ~x54;
assign c1274 =  x65 &  x136 &  x137 &  x272 & ~x321;
assign c1276 =  x22 &  x59 &  x94 &  x194 &  x198 &  x270;
assign c1278 =  x63 &  x72 &  x198 &  x207 &  x270 &  x279 & ~x242 & ~x314;
assign c1280 =  x42 &  x207 & ~x31 & ~x35 & ~x170;
assign c1282 =  x123 & ~x239 & ~x311 & ~x316;
assign c1284 =  x140 &  x203 &  x230 &  x290 & ~x278;
assign c1286 =  x55 &  x190 &  x217 &  x241 &  x313;
assign c1288 =  x267 & ~x42 & ~x240;
assign c1290 =  x203 &  x275 & ~x12 & ~x84 & ~x261;
assign c1292 =  x68 &  x106 &  x139 &  x140 &  x203 &  x275;
assign c1294 =  x154 &  x155 & ~x159 & ~x293;
assign c1296 =  x6 &  x128 &  x154 &  x155 &  x262 &  x263 &  x289;
assign c1298 = ~x8 & ~x35 & ~x39 & ~x166;
assign c1300 =  x245 &  x322 & ~x177;
assign c1302 =  x238 &  x310 & ~x42 & ~x177 & ~x186 & ~x249;
assign c1304 =  x46 & ~x39 & ~x116 & ~x179 & ~x188;
assign c1306 =  x99 &  x207 &  x226 &  x279;
assign c1308 =  x224 &  x225 &  x234 &  x297 & ~x163;
assign c1310 =  x144 & ~x100 & ~x101 & ~x290;
assign c1312 =  x82 &  x98 & ~x114;
assign c1314 =  x118 &  x181 &  x253 & ~x230 & ~x238 & ~x314;
assign c1316 = ~x18 & ~x90 & ~x99 & ~x102 & ~x107 & ~x129;
assign c1318 =  x71 &  x143 &  x278 & ~x17 & ~x186;
assign c1320 =  x40 &  x112 &  x247 & ~x20 & ~x291;
assign c1322 =  x54 &  x314 &  x318;
assign c1324 =  x109 &  x228 &  x244 &  x300 &  x301;
assign c1326 =  x9 &  x81 &  x82 & ~x20;
assign c1328 =  x73 &  x74 &  x136 &  x145 &  x146 &  x208 &  x209 &  x271 &  x280 &  x281;
assign c1330 =  x223 & ~x76 & ~x148 & ~x157 & ~x256;
assign c1332 =  x63 &  x135 &  x160 & ~x305;
assign c1334 =  x39 & ~x9 & ~x17 & ~x18 & ~x26 & ~x81 & ~x89 & ~x90 & ~x98 & ~x107;
assign c1336 =  x61 &  x152 & ~x27 & ~x163;
assign c1338 =  x36 &  x116 &  x171 &  x179 &  x251 & ~x223;
assign c1340 =  x168 &  x169 & ~x65 & ~x137 & ~x173 & ~x200 & ~x245 & ~x272;
assign c1342 =  x70 &  x111 &  x112 &  x142 &  x178 &  x247;
assign c1344 =  x191 & ~x25 & ~x26 & ~x97 & ~x98;
assign c1346 =  x20 &  x120 & ~x90 & ~x95;
assign c1348 =  x138 &  x211 &  x283 & ~x51;
assign c1350 = ~x12 & ~x25 & ~x89 & ~x111;
assign c1352 = ~x4 & ~x13 & ~x21 & ~x49 & ~x84;
assign c1354 = ~x154 & ~x155 & ~x214 & ~x289 & ~x290 & ~x316;
assign c1356 =  x127 &  x128 & ~x158;
assign c1358 = ~x141 & ~x204 & ~x231 & ~x276 & ~x303 & ~x308;
assign c1360 =  x206 &  x278 & ~x78 & ~x150 & ~x232;
assign c1362 =  x33 &  x48 &  x183 & ~x283;
assign c1364 =  x48 &  x242 &  x282 & ~x198;
assign c1366 =  x130 & ~x133 & ~x151;
assign c1368 =  x14 &  x22 &  x77 &  x86 &  x212;
assign c1370 = ~x133 & ~x156 & ~x213;
assign c1372 =  x223 &  x224 &  x225 &  x233 &  x234 &  x297 &  x306;
assign c1374 =  x37 &  x172 & ~x312;
assign c1376 =  x296 & ~x184 & ~x205;
assign c1378 =  x17 &  x192 &  x277;
assign c1380 =  x57 &  x192 &  x193 & ~x65;
assign c1382 =  x89 &  x218 &  x288;
assign c1384 =  x128 &  x263 & ~x35 & ~x313;
assign c1386 = ~x225 & ~x228 & ~x238 & ~x297 & ~x300 & ~x301 & ~x310 & ~x311;
assign c1388 =  x27 &  x162 &  x220 & ~x60;
assign c1390 =  x23 &  x86 & ~x44 & ~x111 & ~x179;
assign c1392 =  x0 &  x3 &  x39 &  x111 &  x246;
assign c1394 = ~x19 & ~x47 & ~x48 & ~x91 & ~x119 & ~x182 & ~x254;
assign c1396 =  x79 &  x115 &  x154 &  x178 &  x214 &  x250 &  x286;
assign c1398 =  x49 &  x112 &  x115 &  x121 &  x178 &  x250;
assign c1400 =  x222 &  x223 & ~x29 & ~x56 & ~x57 & ~x164;
assign c1402 =  x43 &  x250 & ~x17 & ~x64 & ~x89;
assign c1404 =  x279 & ~x18 & ~x81 & ~x90 & ~x313;
assign c1406 =  x42 &  x115 &  x147 &  x177 &  x183;
assign c1408 =  x31 &  x54 &  x174 &  x189;
assign c1410 =  x111 &  x174 &  x246 & ~x68 & ~x94;
assign c1412 =  x44 &  x127 &  x178 &  x179 &  x250;
assign c1414 =  x285 & ~x19 & ~x236 & ~x308;
assign c1416 =  x41 &  x113 &  x135 &  x136 &  x198 &  x207;
assign c1418 =  x77 &  x217 &  x264;
assign c1420 =  x74 &  x234 &  x282 &  x306;
assign c1422 =  x6 & ~x238 & ~x239 & ~x310 & ~x311 & ~x319;
assign c1424 =  x59 &  x194 &  x224 &  x270 &  x271;
assign c1426 =  x100 & ~x40 & ~x49 & ~x112 & ~x121 & ~x175 & ~x184 & ~x247 & ~x256;
assign c1428 =  x69 & ~x82 & ~x83 & ~x108 & ~x109;
assign c1430 =  x5 &  x85 & ~x54 & ~x189;
assign c1432 =  x224 & ~x231 & ~x241 & ~x303;
assign c1434 =  x35 &  x304 & ~x109 & ~x244;
assign c1436 =  x77 &  x130 &  x149 &  x150 &  x212 &  x284;
assign c1438 =  x68 &  x254 & ~x12 & ~x84 & ~x310;
assign c1440 =  x38 &  x110 &  x173 &  x245 & ~x234 & ~x242 & ~x306 & ~x314 & ~x315;
assign c1442 =  x99 &  x217 &  x288;
assign c1444 =  x64 &  x136 & ~x13 & ~x21 & ~x84 & ~x93;
assign c1446 =  x315 & ~x137 & ~x138 & ~x173 & ~x272 & ~x273;
assign c1448 =  x63 &  x102 &  x129 &  x135 &  x264;
assign c1450 = ~x73 & ~x208 & ~x226 & ~x234 & ~x235 & ~x298 & ~x306;
assign c1452 =  x26 &  x107 &  x189 &  x216;
assign c1454 =  x74 &  x75 &  x282 & ~x103 & ~x130;
assign c1456 =  x60 & ~x11 & ~x29 & ~x38 & ~x83 & ~x164;
assign c1458 =  x223 &  x233 &  x305 & ~x56 & ~x163;
assign c1460 =  x145 &  x146 &  x280 & ~x80 & ~x188 & ~x215;
assign c1462 = ~x30 & ~x222 & ~x237 & ~x299;
assign c1464 =  x23 &  x25 &  x129 &  x264;
assign c1466 =  x70 &  x119 &  x120 &  x205 & ~x64;
assign c1468 =  x126 &  x127 &  x153 &  x261 &  x279 &  x288;
assign c1470 =  x84 &  x85 &  x112 & ~x81;
assign c1472 = ~x20 & ~x21 & ~x46 & ~x47 & ~x92 & ~x118 & ~x119;
assign c1474 =  x55 &  x149 &  x190 &  x241;
assign c1476 =  x103 & ~x29 & ~x96;
assign c1478 =  x12 &  x21 &  x84 &  x93 &  x233 &  x305;
assign c1480 =  x239 &  x311 &  x318 & ~x139;
assign c1482 = ~x127 & ~x128 & ~x154 & ~x155 & ~x262 & ~x263 & ~x289 & ~x290 & ~x316 & ~x317;
assign c1484 =  x170 &  x178 &  x179 & ~x82;
assign c1486 =  x252 & ~x59 & ~x157 & ~x292;
assign c1488 =  x127 &  x262 &  x263 & ~x96;
assign c1490 =  x192 & ~x33 & ~x60 & ~x61 & ~x168 & ~x196;
assign c1492 =  x91 & ~x240 & ~x303;
assign c1494 =  x182 &  x253 & ~x24 & ~x96;
assign c1496 =  x232 &  x292 & ~x268;
assign c1498 =  x48 &  x115 &  x319;
assign c1500 =  x175 &  x194 & ~x13;
assign c1502 =  x14 &  x21 &  x86 &  x93 & ~x96;
assign c1504 =  x125 &  x243 &  x260 & ~x233 & ~x305;
assign c1506 =  x283 & ~x72 & ~x207 & ~x252;
assign c1508 =  x53 &  x212 &  x219;
assign c1510 = ~x15 & ~x115 & ~x250 & ~x322;
assign c1512 =  x107 &  x270 & ~x9;
assign c1514 =  x132 & ~x107 & ~x153 & ~x288;
assign c1516 =  x164 & ~x47 & ~x73 & ~x208 & ~x209;
assign c1518 =  x55 &  x163 &  x190 &  x219 & ~x195;
assign c1520 =  x2 &  x122 &  x322;
assign c1522 =  x122 & ~x100 & ~x101 & ~x182;
assign c1524 =  x55 &  x103 &  x190 &  x275;
assign c1526 =  x118 &  x182 &  x253 &  x254;
assign c1528 = ~x48 & ~x105 & ~x272;
assign c1530 =  x246 & ~x30 & ~x190 & ~x191;
assign c1532 =  x3 &  x82 &  x108;
assign c1534 =  x114 &  x118 &  x119 &  x254 & ~x53 & ~x125 & ~x260;
assign c1536 =  x65 &  x137 & ~x212 & ~x224 & ~x225 & ~x297;
assign c1538 =  x305 & ~x134 & ~x160 & ~x268 & ~x269 & ~x295;
assign c1540 =  x42 & ~x27 & ~x39 & ~x44 & ~x162 & ~x319;
assign c1542 =  x81 &  x99 & ~x105;
assign c1544 =  x107 & ~x20 & ~x92 & ~x101;
assign c1546 =  x5 &  x12 &  x13 &  x21 &  x48 &  x84;
assign c1548 =  x215 &  x287 & ~x238 & ~x239 & ~x310 & ~x311 & ~x320;
assign c1550 =  x52 &  x53 &  x116 &  x124 &  x125 &  x188 &  x260 & ~x141;
assign c1552 =  x157 &  x205 &  x242 &  x314 & ~x271;
assign c1554 =  x78 & ~x179 & ~x184 & ~x256;
assign c1556 =  x71 &  x143 & ~x12 & ~x84 & ~x319;
assign c1558 =  x153 &  x288 & ~x91 & ~x96;
assign c1560 =  x14 &  x22 &  x46 &  x94 &  x118 &  x253;
assign c1562 =  x113 &  x176 &  x248 & ~x118 & ~x200;
assign c1564 =  x150 & ~x22 & ~x23 & ~x216;
assign c1566 =  x0 &  x17 &  x89 &  x203 &  x302;
assign c1568 =  x42 &  x99 &  x114 & ~x11;
assign c1570 =  x70 &  x142 &  x205 &  x277 & ~x128 & ~x262 & ~x263;
assign c1572 =  x117 & ~x132 & ~x165;
assign c1574 =  x14 &  x90 &  x225;
assign c1576 =  x108 &  x125 &  x260 & ~x49;
assign c1578 =  x51 &  x52 &  x123 &  x124 &  x187 &  x259 & ~x40 & ~x196;
assign c1580 =  x96 &  x142 &  x277 & ~x18 & ~x26 & ~x98;
assign c1582 =  x29 &  x82 &  x129;
assign c1584 =  x5 & ~x128 & ~x154 & ~x289;
assign c1586 =  x122 &  x140 &  x159 &  x203 &  x275;
assign c1588 =  x33 & ~x302 & ~x310 & ~x320;
assign c1590 =  x229 &  x230 &  x302 & ~x61 & ~x196;
assign c1592 =  x156 &  x263 & ~x300 & ~x301;
assign c1594 =  x291 & ~x12 & ~x92;
assign c1596 =  x0 &  x1 &  x9 &  x89 &  x228;
assign c1598 =  x51 &  x123 &  x186 &  x288 & ~x85;
assign c11 =  x79 &  x133 & ~x253 & ~x282;
assign c13 =  x2 &  x166 & ~x202 & ~x243;
assign c15 =  x101 &  x123 & ~x138;
assign c17 =  x240 &  x289 & ~x304;
assign c19 =  x16 & ~x99 & ~x105 & ~x262;
assign c111 =  x256 &  x308 & ~x277;
assign c113 =  x83 &  x148 &  x267 & ~x48;
assign c115 =  x96 &  x123 &  x267 & ~x93 & ~x115;
assign c117 =  x26 &  x227 & ~x138;
assign c119 =  x306 & ~x318 & ~x320;
assign c121 =  x76 &  x213 & ~x116;
assign c123 =  x46 &  x98 &  x118 &  x201;
assign c125 =  x78 &  x87 &  x103;
assign c127 =  x51 & ~x136 & ~x212 & ~x300;
assign c129 =  x88 &  x227 & ~x105;
assign c131 =  x240 &  x314 & ~x39;
assign c133 =  x103 &  x132 &  x290 & ~x275;
assign c135 =  x52 &  x193 & ~x105;
assign c137 =  x123 &  x148 &  x224 &  x314;
assign c139 =  x168 &  x269 &  x312 &  x316;
assign c141 =  x110 &  x227 & ~x126 & ~x140 & ~x207;
assign c143 =  x38 & ~x86 & ~x100 & ~x130;
assign c145 =  x160 &  x209 & ~x73 & ~x244;
assign c147 =  x50 & ~x94 & ~x164 & ~x166 & ~x192 & ~x202;
assign c149 =  x208 &  x229 & ~x44 & ~x116;
assign c151 =  x93 & ~x105 & ~x265;
assign c153 =  x60 &  x71 &  x294 & ~x0 & ~x52;
assign c155 =  x71 &  x80 & ~x0 & ~x129 & ~x286;
assign c157 =  x124 & ~x220 & ~x311;
assign c159 =  x140 &  x199 &  x248 & ~x268;
assign c161 = ~x0 & ~x18 & ~x106 & ~x163 & ~x192 & ~x310;
assign c163 =  x101 &  x177 &  x289 & ~x318;
assign c165 =  x258 & ~x12 & ~x184;
assign c167 =  x5 &  x15 &  x33 &  x94 &  x242;
assign c169 = ~x4 & ~x263 & ~x269 & ~x296;
assign c171 =  x87 &  x128 & ~x226;
assign c173 = ~x83 & ~x228 & ~x291;
assign c175 =  x91 &  x229 & ~x84 & ~x304;
assign c177 =  x161 &  x168 &  x316;
assign c179 =  x103 &  x132 &  x294;
assign c181 =  x209 &  x272 &  x290;
assign c183 =  x132 & ~x57 & ~x75 & ~x282;
assign c185 =  x70 & ~x162 & ~x220 & ~x269;
assign c187 =  x131 &  x132 &  x176 & ~x84;
assign c189 =  x190 &  x208 & ~x228;
assign c191 =  x6 &  x221 & ~x100;
assign c193 =  x141 &  x255 & ~x55 & ~x58 & ~x293 & ~x320;
assign c195 =  x190 & ~x49 & ~x211;
assign c197 = ~x148 & ~x251 & ~x270 & ~x282;
assign c199 =  x160 & ~x12 & ~x146 & ~x280;
assign c1101 =  x185 &  x275 & ~x304 & ~x321 & ~x323;
assign c1103 =  x243 & ~x1 & ~x151 & ~x220;
assign c1105 =  x26 &  x294 &  x320 & ~x39;
assign c1107 = ~x152 & ~x157 & ~x260 & ~x265 & ~x316;
assign c1109 =  x80 &  x106 &  x206;
assign c1111 =  x269 &  x312 &  x316 & ~x280;
assign c1113 =  x24 &  x101 & ~x30;
assign c1115 =  x21 &  x52 & ~x127;
assign c1117 = ~x78 & ~x128 & ~x294 & ~x312;
assign c1119 =  x114 &  x235 & ~x64 & ~x198 & ~x296;
assign c1121 =  x157 &  x312 &  x315;
assign c1123 =  x123 &  x144 &  x315 & ~x255;
assign c1125 =  x141 &  x247 &  x315;
assign c1127 =  x155 & ~x86 & ~x275;
assign c1129 =  x184 &  x222 & ~x43;
assign c1131 =  x33 &  x315 &  x322 & ~x68 & ~x248;
assign c1133 = ~x54 & ~x162 & ~x220 & ~x259;
assign c1135 = ~x28 & ~x102 & ~x321;
assign c1137 =  x105 &  x323 & ~x21;
assign c1139 =  x16 &  x79 & ~x103 & ~x154;
assign c1141 = ~x76 & ~x133;
assign c1143 =  x63 & ~x89 & ~x192 & ~x201 & ~x219;
assign c1145 = ~x57 & ~x169 & ~x219 & ~x227 & ~x283;
assign c1147 =  x76 &  x133 & ~x41 & ~x140 & ~x250;
assign c1149 =  x67 & ~x147 & ~x174;
assign c1151 =  x20 &  x303 & ~x64 & ~x264;
assign c1153 =  x307 & ~x156 & ~x291 & ~x318 & ~x319;
assign c1155 =  x97 &  x290 &  x315;
assign c1157 =  x78 &  x103 &  x213 &  x312 &  x323;
assign c1159 =  x217 &  x244 & ~x11 & ~x160;
assign c1161 = ~x76 & ~x134 & ~x285 & ~x301;
assign c1163 = ~x13 & ~x85 & ~x125 & ~x151 & ~x218;
assign c1165 =  x113 & ~x65 & ~x191 & ~x220 & ~x268;
assign c1167 =  x187 &  x227 & ~x145 & ~x288;
assign c1169 = ~x38 & ~x150 & ~x151 & ~x201;
assign c1171 =  x76 &  x308 & ~x257;
assign c1173 =  x106 &  x132 & ~x99 & ~x151;
assign c1175 =  x148 &  x215 &  x312 &  x316;
assign c1177 =  x96 &  x258;
assign c1179 =  x204 &  x276 & ~x1 & ~x27 & ~x28 & ~x57 & ~x162 & ~x192;
assign c1181 = ~x45 & ~x60 & ~x169 & ~x289;
assign c1183 =  x173 &  x245 & ~x111 & ~x255;
assign c1185 =  x25 & ~x100;
assign c1187 =  x38 &  x209 & ~x262;
assign c1189 =  x22 &  x195 & ~x84;
assign c1191 =  x158 &  x292 &  x294 & ~x84;
assign c1193 =  x173 & ~x237 & ~x290;
assign c1195 =  x267 & ~x64 & ~x99;
assign c1197 =  x316 & ~x300;
assign c1199 =  x56 &  x245 & ~x143;
assign c1201 =  x193 &  x269 & ~x99;
assign c1203 =  x195 &  x264 & ~x105 & ~x154;
assign c1205 = ~x12 & ~x138 & ~x255;
assign c1207 =  x290 & ~x130 & ~x261;
assign c1209 =  x3 &  x65 & ~x72 & ~x287;
assign c1211 =  x71 &  x175 &  x188 &  x247 & ~x271;
assign c1213 = ~x134 & ~x173 & ~x192 & ~x223 & ~x311;
assign c1215 =  x33 &  x64 & ~x241 & ~x300;
assign c1217 =  x107 &  x323 & ~x217;
assign c1219 =  x14 &  x15 &  x24 &  x101 &  x123;
assign c1221 =  x25 & ~x132;
assign c1223 =  x87 &  x269 & ~x81 & ~x270;
assign c1225 =  x97 &  x200 &  x320 & ~x131;
assign c1227 =  x159 &  x267 & ~x4 & ~x32 & ~x242;
assign c1229 =  x281 & ~x28 & ~x64 & ~x197;
assign c1231 =  x20 &  x242 &  x279;
assign c1233 =  x200 & ~x53 & ~x139 & ~x144;
assign c1235 =  x314 & ~x306;
assign c1237 = ~x21 & ~x57 & ~x120;
assign c1239 = ~x157 & ~x247 & ~x278 & ~x296 & ~x323;
assign c1241 =  x315 & ~x2 & ~x153 & ~x164;
assign c1243 =  x52 &  x303 & ~x82 & ~x194;
assign c1245 =  x47 & ~x64 & ~x162 & ~x217 & ~x226;
assign c1247 =  x148 &  x188 &  x294;
assign c1249 =  x1 &  x85 &  x159;
assign c1251 =  x47 &  x159 & ~x129;
assign c1253 =  x103 &  x105 & ~x93;
assign c1255 = ~x140 & ~x217 & ~x284 & ~x298;
assign c1257 = ~x215 & ~x233 & ~x256;
assign c1259 =  x57 &  x303 & ~x100 & ~x280;
assign c1261 =  x285 & ~x156 & ~x253;
assign c1263 = ~x193 & ~x264;
assign c1265 =  x84 & ~x37 & ~x109 & ~x268;
assign c1267 =  x11 &  x128 &  x245;
assign c1269 =  x58 &  x273 & ~x127 & ~x280;
assign c1271 =  x17 &  x321 & ~x212;
assign c1273 =  x78 &  x213 & ~x84 & ~x273 & ~x280 & ~x297;
assign c1275 =  x71 &  x80 &  x87 &  x131;
assign c1277 =  x20 &  x112;
assign c1279 =  x90 &  x131 &  x269 & ~x199;
assign c1281 =  x5 &  x67 &  x166 &  x197 & ~x2;
assign c1283 =  x41 &  x282 &  x286 & ~x27;
assign c1285 =  x80 &  x276 & ~x219;
assign c1287 = ~x1 & ~x168 & ~x192 & ~x195;
assign c1289 =  x53 & ~x244;
assign c1291 = ~x146 & ~x187 & ~x269;
assign c1293 =  x141 &  x234;
assign c1295 =  x140 &  x203 & ~x155 & ~x156;
assign c1297 =  x280 & ~x296 & ~x310 & ~x321;
assign c1299 =  x96 &  x123 &  x154 &  x263 &  x290 & ~x111;
assign c1301 =  x11 &  x38 &  x110 &  x311 & ~x255;
assign c1303 =  x69 & ~x126 & ~x260 & ~x279;
assign c1305 =  x265 &  x269 &  x293 &  x321;
assign c1307 = ~x106 & ~x219 & ~x229 & ~x287;
assign c1309 =  x97 &  x310 & ~x271;
assign c1311 =  x78 &  x258 & ~x39 & ~x99 & ~x156;
assign c1313 =  x47 &  x74 & ~x72 & ~x148 & ~x153;
assign c1315 =  x7 &  x115 & ~x24 & ~x100 & ~x105;
assign c1317 =  x64 &  x172 & ~x313;
assign c1319 =  x151 &  x186 &  x312 & ~x34;
assign c1321 =  x290 &  x323 & ~x118;
assign c1323 =  x56 &  x106 &  x247 & ~x300;
assign c1325 =  x18 &  x40 &  x211 &  x315 &  x321;
assign c1327 =  x11 & ~x73 & ~x91 & ~x154 & ~x253;
assign c1329 =  x141 & ~x28 & ~x126 & ~x217 & ~x311;
assign c1331 = ~x24 & ~x90 & ~x107 & ~x127 & ~x301;
assign c1333 =  x77 & ~x281 & ~x286 & ~x300;
assign c1335 = ~x6 & ~x78 & ~x159 & ~x220 & ~x283;
assign c1337 =  x51 &  x150 & ~x136 & ~x226;
assign c1339 =  x276 & ~x148 & ~x292 & ~x320;
assign c1341 =  x101 &  x285 &  x312 & ~x68;
assign c1343 =  x5 &  x256 &  x263 &  x312;
assign c1345 =  x162 &  x285 & ~x210 & ~x291;
assign c1347 =  x102 &  x121 &  x159 &  x294 & ~x122;
assign c1349 =  x38 &  x268 & ~x203 & ~x282;
assign c1351 =  x52 & ~x19 & ~x258;
assign c1353 =  x257 & ~x35 & ~x201 & ~x236;
assign c1355 =  x182 & ~x5 & ~x41 & ~x217;
assign c1357 =  x312 & ~x68 & ~x147 & ~x284;
assign c1359 =  x148 &  x307;
assign c1361 = ~x46 & ~x111;
assign c1363 =  x10 &  x102 &  x167;
assign c1365 =  x214 & ~x54 & ~x104 & ~x153;
assign c1367 = ~x181 & ~x257 & ~x262 & ~x266;
assign c1369 =  x265 &  x269 &  x312 &  x316;
assign c1371 =  x5 &  x148 &  x152;
assign c1373 =  x271 & ~x151 & ~x160 & ~x209;
assign c1375 =  x21 &  x129 & ~x99 & ~x100 & ~x262;
assign c1377 =  x320 & ~x93 & ~x153;
assign c1379 =  x218 & ~x151 & ~x219;
assign c1381 =  x122 & ~x33 & ~x279 & ~x319;
assign c1383 =  x51 &  x168 &  x256;
assign c1385 =  x40 &  x78 &  x134 &  x265 &  x312;
assign c1387 =  x68 &  x122 & ~x129 & ~x259;
assign c1389 =  x82 & ~x292 & ~x322;
assign c1391 =  x52 &  x102 &  x321 & ~x297;
assign c1393 =  x208 &  x239 & ~x130 & ~x316;
assign c1395 =  x154 &  x222 &  x289 & ~x237 & ~x259;
assign c1397 =  x106 & ~x47 & ~x210 & ~x281;
assign c1399 =  x24 &  x96 &  x240 &  x258 & ~x84 & ~x246;
assign c1401 =  x13 &  x15 &  x60 & ~x118;
assign c1403 =  x154 & ~x155;
assign c1405 = ~x11 & ~x137 & ~x189 & ~x304;
assign c1407 = ~x6 & ~x56 & ~x65 & ~x168 & ~x191 & ~x227;
assign c1409 =  x24 & ~x18 & ~x97 & ~x193 & ~x219;
assign c1411 =  x79 &  x250 & ~x105 & ~x262;
assign c1413 =  x15 &  x211 &  x317 & ~x68;
assign c1415 =  x261 & ~x295 & ~x318 & ~x320 & ~x322 & ~x323;
assign c1417 =  x229 & ~x126 & ~x248 & ~x265;
assign c1419 = ~x146 & ~x241 & ~x291 & ~x318;
assign c1421 =  x155 &  x240 & ~x105 & ~x266;
assign c1423 =  x140 &  x142 & ~x6;
assign c1425 =  x58 &  x67 &  x76 &  x242;
assign c1427 =  x21 & ~x10 & ~x37 & ~x267 & ~x268;
assign c1429 =  x281 &  x317 & ~x96;
assign c1431 =  x241 &  x254 & ~x309;
assign c1433 = ~x39 & ~x273 & ~x313;
assign c1435 =  x203 & ~x308 & ~x313 & ~x321 & ~x323;
assign c1437 =  x267 & ~x8 & ~x22 & ~x188;
assign c1439 =  x186 & ~x11 & ~x39;
assign c1441 =  x46 &  x181 &  x271 & ~x268;
assign c1443 =  x36 &  x293 & ~x84;
assign c1445 =  x118 &  x122 & ~x319 & ~x321;
assign c1447 =  x101 &  x123 &  x128 &  x177 &  x249 &  x289;
assign c1449 =  x94 &  x98 &  x175 &  x272;
assign c1451 =  x56 &  x315 & ~x39 & ~x126;
assign c1453 =  x244 & ~x134 & ~x256 & ~x316;
assign c1455 = ~x129 & ~x263 & ~x308;
assign c1457 =  x30 & ~x36 & ~x49 & ~x139;
assign c1459 =  x44 &  x98 & ~x70;
assign c1461 = ~x73 & ~x91 & ~x113 & ~x118 & ~x167;
assign c1463 =  x278 &  x296 &  x316 &  x322 & ~x30;
assign c1465 =  x184 & ~x12 & ~x48 & ~x100;
assign c1467 =  x200 &  x245 & ~x207 & ~x261;
assign c1469 =  x53 & ~x144 & ~x153;
assign c1471 =  x101 &  x133 &  x157 &  x269;
assign c1473 =  x16 &  x38 &  x133;
assign c1475 =  x50 &  x69 & ~x264;
assign c1477 = ~x1 & ~x5 & ~x124 & ~x316;
assign c1479 =  x67 &  x315 &  x316 &  x323;
assign c1481 =  x199 & ~x152 & ~x166 & ~x296;
assign c1483 =  x236 & ~x39 & ~x212;
assign c1485 =  x276 &  x307 & ~x295 & ~x320 & ~x322;
assign c1487 =  x190 & ~x47 & ~x175;
assign c1489 =  x91 &  x172 & ~x156 & ~x264;
assign c1491 = ~x193 & ~x265 & ~x269 & ~x315 & ~x316;
assign c1493 =  x179 &  x183 & ~x5 & ~x193 & ~x194;
assign c1495 =  x87 &  x93 &  x231 & ~x295;
assign c1497 =  x73 &  x128 &  x132 & ~x3;
assign c1499 =  x132 &  x245 & ~x113 & ~x181;
assign c1501 =  x25 &  x79 &  x321 & ~x280;
assign c1503 =  x95 &  x265 &  x303;
assign c1505 =  x22 &  x69 & ~x156;
assign c1507 =  x74 &  x292 & ~x255;
assign c1509 =  x25 &  x259 & ~x99 & ~x318;
assign c1511 =  x15 &  x71 &  x263;
assign c1513 =  x132 & ~x75 & ~x317;
assign c1515 = ~x2 & ~x27 & ~x64 & ~x220 & ~x227;
assign c1517 =  x101 &  x143 &  x157 &  x161 &  x316;
assign c1519 =  x132 &  x196 & ~x75 & ~x120;
assign c1521 =  x150 & ~x115 & ~x277;
assign c1523 =  x50 &  x105 &  x224 &  x231;
assign c1525 =  x184 &  x285;
assign c1527 =  x175 &  x209 & ~x39;
assign c1529 =  x136 & ~x90 & ~x108;
assign c1531 =  x102 &  x155 &  x287 &  x312;
assign c1533 =  x33 &  x106 &  x267 & ~x286;
assign c1535 =  x66 &  x214 & ~x86 & ~x159;
assign c1537 = ~x133 & ~x223 & ~x316;
assign c1539 =  x185 & ~x123 & ~x254;
assign c1541 =  x28 &  x150 & ~x288 & ~x318;
assign c1543 =  x151 & ~x255 & ~x300;
assign c1545 =  x160 &  x171 & ~x112;
assign c1547 =  x203 & ~x4 & ~x5 & ~x134;
assign c1549 =  x290 & ~x36 & ~x192 & ~x218 & ~x251;
assign c1551 =  x150 &  x186 &  x236 &  x312 & ~x153;
assign c1553 =  x123 & ~x3 & ~x115;
assign c1555 =  x105 &  x159 &  x311 & ~x286;
assign c1557 =  x92 &  x182 &  x254 &  x281 & ~x95;
assign c1559 =  x225 &  x302 & ~x228 & ~x320;
assign c1561 =  x75 & ~x77 & ~x102 & ~x153 & ~x157 & ~x266;
assign c1563 =  x11 & ~x107 & ~x145 & ~x289;
assign c1565 =  x184 &  x285 & ~x230 & ~x271;
assign c1567 =  x40 &  x120 & ~x0 & ~x1 & ~x220;
assign c1569 =  x42 &  x47 &  x265 &  x316;
assign c1571 =  x12 &  x151 &  x200 & ~x262;
assign c1573 =  x52 &  x303 & ~x105;
assign c1575 = ~x228 & ~x259 & ~x290 & ~x319;
assign c1577 =  x122 &  x170;
assign c1579 =  x71 &  x242 & ~x7 & ~x111 & ~x230;
assign c1581 =  x159 &  x168 & ~x291;
assign c1583 =  x65 &  x106 &  x289 & ~x217;
assign c1585 =  x21 &  x151 &  x236 &  x286 &  x290;
assign c1587 =  x121 &  x128 &  x312;
assign c1589 =  x52 & ~x0 & ~x19 & ~x220;
assign c1591 =  x2 &  x5 &  x164 & ~x322;
assign c1593 =  x106 &  x132 &  x159 & ~x115 & ~x255;
assign c1595 =  x21 &  x87 & ~x125 & ~x228;
assign c1597 =  x227 &  x250 & ~x53;
assign c1599 = ~x128 & ~x157 & ~x265 & ~x316;

endmodule