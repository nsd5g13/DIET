module tm( x0,x1,x2,x3,x4,x5,x6,x7,x8,x9,x10,x11,x12,x13,x14,x15,x16,x17,x18,x19,x20,x21,x22,x23,x24,x25,x26,x27,x28,x29,x30,x31,x32,x33,x34,x35,x36,x37,x38,x39,x40,x41,x42,x43,x44,x45,x46,x47,x48,x49,x50,x51,x52,x53,x54,x55,x56,x57,x58,x59,x60,x61,x62,x63,x64,x65,x66,x67,x68,x69,x70,x71,x72,x73,x74,x75,x76,x77,x78,x79,x80,x81,x82,x83,x84,x85,x86,x87,x88,x89,x90,x91,x92,x93,x94,x95,x96,x97,x98,x99,x100,x101,x102,x103,x104,x105,x106,x107,x108,x109,x110,x111,x112,x113,x114,x115,x116,x117,x118,x119,x120,x121,x122,x123,x124,x125,x126,x127,x128,x129,x130,x131,x132,x133,x134,x135,x136,x137,x138,x139,x140,x141,x142,x143,x144,x145,x146,x147,x148,x149,x150,x151,x152,x153,x154,x155,x156,x157,x158,x159,x160,x161,x162,x163,x164,x165,x166,x167,x168,x169,x170,x171,x172,x173,x174,x175,x176,x177,x178,x179,x180,x181,x182,x183,x184,x185,x186,x187,x188,x189,x190,x191,x192,x193,x194,x195,x196,x197,x198,x199,x200,x201,x202,x203,x204,x205,x206,x207,x208,x209,x210,x211,x212,x213,x214,x215,x216,x217,x218,x219,x220,x221,x222,x223,x224,x225,x226,x227,x228,x229,x230,x231,x232,x233,x234,x235,x236,x237,x238,x239,x240,x241,x242,x243,x244,x245,x246,x247,x248,x249,x250,x251,x252,x253,x254,x255,x256,x257,x258,x259,x260,x261,x262,x263,x264,x265,x266,x267,x268,x269,x270,x271,x272,x273,x274,x275,x276,x277,x278,x279,x280,x281,x282,x283,x284,x285,x286,x287,x288,x289,x290,x291,x292,x293,x294,x295,x296,x297,x298,x299,x300,x301,x302,x303,x304,x305,x306,x307,x308,x309,x310,x311,x312,x313,x314,x315,x316,x317,x318,x319,x320,x321,x322,x323,x324,x325,x326,x327,x328,x329,x330,x331,x332,x333,x334,x335,x336,x337,x338,x339,x340,x341,x342,x343,x344,x345,x346,x347,x348,x349,x350,x351,x352,x353,x354,x355,x356,x357,x358,x359,x360,x361,x362,x363,x364,x365,x366,x367,x368,x369,x370,x371,x372,x373,x374,x375,x376,x377,x378,x379,x380,x381,x382,x383,x384,x385,x386,x387,x388,x389,x390,x391,x392,x393,x394,x395,x396,x397,x398,x399,x400,x401,x402,x403,x404,x405,x406,x407,x408,x409,x410,x411,x412,x413,x414,x415,x416,x417,x418,x419,x420,x421,x422,x423,x424,x425,x426,x427,x428,x429,x430,x431,x432,x433,x434,x435,x436,x437,x438,x439,x440,x441,x442,x443,x444,x445,x446,x447,x448,x449,x450,x451,x452,x453,x454,x455,x456,x457,x458,x459,x460,x461,x462,x463,x464,x465,x466,x467,x468,x469,x470,x471,x472,x473,x474,x475,x476,x477,x478,x479,x480,x481,x482,x483,x484,x485,x486,x487,x488,x489,x490,x491,x492,x493,x494,x495,x496,x497,x498,x499,x500,x501,x502,x503,x504,x505,x506,x507,x508,x509,x510,x511,x512,x513,x514,x515,x516,x517,x518,x519,x520,x521,x522,x523,x524,x525,x526,x527,x528,x529,x530,x531,x532,x533,x534,x535,x536,x537,x538,x539,x540,x541,x542,x543,x544,x545,x546,x547,x548,x549,x550,x551,x552,x553,x554,x555,x556,x557,x558,x559,x560,x561,x562,x563,x564,x565,x566,x567,x568,x569,x570,x571,x572,x573,x574,x575,x576,x577,x578,x579,x580,x581,x582,x583,x584,x585,x586,x587,x588,x589,x590,x591,x592,x593,x594,x595,x596,x597,x598,x599,x600,x601,x602,x603,x604,x605,x606,x607,x608,x609,x610,x611,x612,x613,x614,x615,x616,x617,x618,x619,x620,x621,x622,x623,x624,x625,x626,x627,x628,x629,x630,x631,x632,x633,x634,x635,x636,x637,x638,x639,x640,x641,x642,x643,x644,x645,x646,x647,x648,x649,x650,x651,x652,x653,x654,x655,x656,x657,x658,x659,x660,x661,x662,x663,x664,x665,x666,x667,x668,x669,x670,x671,x672,x673,x674,x675,x676,x677,x678,x679,x680,x681,x682,x683,x684,x685,x686,x687,x688,x689,x690,x691,x692,x693,x694,x695,x696,x697,x698,x699,x700,x701,x702,x703,x704,x705,x706,x707,x708,x709,x710,x711,x712,x713,x714,x715,x716,x717,x718,x719,x720,x721,x722,x723,x724,x725,x726,x727,x728,x729,x730,x731,x732,x733,x734,x735,x736,x737,x738,x739,x740,x741,x742,x743,x744,x745,x746,x747,x748,x749,x750,x751,x752,x753,x754,x755,x756,x757,x758,x759,x760,x761,x762,x763,x764,x765,x766,x767,x768,x769,x770,x771,x772,x773,x774,x775,x776,x777,x778,x779,x780,x781,x782,x783,c38,c6296,c8194,c0144,c7168,c3161,c623,c08,c050,c753,c239,c062,c3123,c962,c177,c2209,c9294,c93,c392,c4137,c5193,c122,c0170,c1199,c1279,c0290,c3163,c35,c2213,c0161,c4237,c8277,c875,c199,c139,c6208,c3271,c0201,c6271,c4182,c0209,c0193,c387,c7243,c924,c7108,c3117,c91,c9199,c6105,c957,c5244,c7221,c932,c9119,c8202,c771,c1121,c9156,c685,c470,c378,c180,c6174,c295,c365,c137,c5253,c9158,c5278,c179,c0231,c4145,c946,c5225,c5246,c9265,c626,c4129,c0124,c2216,c6278,c447,c2174,c5243,c6128,c5223,c255,c6195,c190,c469,c95,c2183,c4271,c357,c664,c791,c9120,c3233,c2166,c9219,c938,c785,c4115,c2223,c651,c899,c0135,c0224,c6298,c0154,c1239,c4242,c0292,c9128,c920,c484,c4204,c8104,c0293,c2221,c5129,c0277,c5281,c5292,c5265,c7244,c836,c960,c191,c874,c9148,c1264,c8119,c7130,c0270,c6215,c0133,c2181,c9297,c7270,c935,c0178,c0299,c3159,c5115,c8191,c816,c114,c6149,c450,c4222,c27,c1293,c210,c1186,c344,c5286,c9125,c4235,c377,c6224,c6205,c8195,c070,c7235,c3142,c5119,c1195,c5255,c2142,c4206,c8295,c5170,c2292,c6135,c321,c5240,c2180,c4134,c554,c1242,c1193,c252,c3126,c481,c214,c5111,c1252,c2293,c493,c218,c5126,c620,c0197,c2191,c1166,c7203,c8156,c788,c937,c956,c2111,c7163,c3147,c9208,c1269,c2201,c4223,c318,c545,c832,c3152,c4226,c3241,c0166,c3208,c1180,c2154,c970,c358,c3209,c0137,c5175,c9177,c1271,c811,c1203,c548,c6147,c8243,c0216,c9124,c349,c1236,c4107,c7214,c7266,c864,c9201,c656,c1161,c4266,c645,c7134,c0284,c7264,c3243,c9190,c2207,c5264,c683,c9269,c9204,c5155,c77,c2187,c076,c0297,c1245,c1174,c3128,c7157,c910,c166,c953,c8267,c896,c1140,c13,c87,c272,c1155,c427,c611,c0229,c6189,c4126,c559,c297,c8111,c9252,c0127,c212,c262,c8248,c016,c23,c66,c674,c939,c977,c0234,c9135,c2297,c591,c3193,c087,c7268,c7180,c9205,c9150,c1154,c12,c3279,c216,c690,c715,c9292,c6153,c368,c3212,c5237,c9253,c115,c5251,c519,c5168,c211,c0245,c6265,c347,c615,c693,c0276,c3182,c170,c0149,c142,c3215,c4207,c3127,c2149,c464,c538,c446,c9145,c933,c7138,c0184,c9175,c7121,c2215,c442,c931,c0174,c7247,c39,c7155,c348,c088,c116,c598,c3291,c4211,c52,c5232,c9151,c0195,c023,c661,c512,c747,c5146,c1226,c2259,c054,c1200,c4148,c6130,c677,c6273,c725,c98,c46,c7286,c9105,c3216,c9164,c25,c217,c2169,c1232,c9154,c4247,c1144,c1251,c1257,c9107,c335,c7145,c057,c533,c927,c0114,c0132,c737,c4273,c440,c589,c792,c4289,c8219,c8291,c3148,c9237,c6113,c7105,c813,c0217,c4109,c90,c6252,c394,c520,c7225,c43,c0122,c3282,c7147,c327,c6248,c369,c165,c4205,c9243,c892,c6158,c3111,c0176,c3295,c6173,c528,c232,c9100,c071,c0177,c9216,c7154,c3281,c547,c793,c0222,c6125,c6241,c624,c3229,c680,c8160,c1230,c5201,c1142,c526,c126,c7280,c861,c4239,c7279,c5142,c7184,c8174,c8176,c734,c7287,c820,c9165,c280,c279,c8161,c2122,c6170,c19,c3139,c185,c2281,c4270,c2152,c3177,c5171,c0238,c035,c0117,c722,c8221,c73,c879,c150,c7102,c6276,c0131,c6254,c948,c058,c0215,c2283,c2200,c3236,c5271,c873,c8270,c3140,c492,c2222,c4298,c68,c0196,c969,c483,c5176,c5295,c8288,c1281,c997,c192,c018,c3294,c0283,c455,c2123,c189,c4128,c668,c8100,c173,c479,c638,c0241,c4119,c3115,c6259,c9121,c866,c521,c1106,c544,c1233,c3156,c8263,c422,c2134,c3245,c64,c3119,c0136,c0103,c7255,c048,c5274,c88,c419,c1178,c6151,c460,c9236,c6101,c2116,c0112,c5268,c4161,c0107,c6238,c0260,c5140,c5279,c621,c7110,c356,c8276,c3114,c678,c2178,c7164,c2238,c5150,c7124,c1116,c313,c8183,c3183,c2240,c4261,c220,c2228,c4249,c7173,c6201,c3172,c375,c259,c1295,c3132,c1219,c3213,c373,c1130,c1192,c3157,c3259,c1262,c1225,c1229,c55,c9281,c8196,c8150,c4293,c75,c7201,c867,c473,c8149,c4216,c119,c8290,c986,c3125,c4106,c4178,c786,c6227,c9256,c4102,c0115,c9191,c8224,c171,c3200,c0298,c5294,c583,c9167,c0249,c557,c8264,c0218,c1113,c660,c7211,c649,c629,c0203,c857,c6137,c6178,c6166,c719,c594,c2140,c964,c2263,c1127,c9123,c2220,c5218,c6292,c934,c6243,c1198,c0169,c3274,c1266,c5269,c420,c7188,c7238,c2161,c8118,c7234,c9147,c5164,c8292,c4127,c5215,c0274,c7114,c4123,c288,c4156,c686,c6262,c9171,c371,c353,c031,c9106,c145,c4164,c745,c9162,c3278,c5160,c4187,c748,c2232,c841,c752,c153,c2163,c625,c835,c9229,c8182,c186,c1253,c240,c458,c4238,c5187,c643,c6275,c2112,c4160,c4253,c7149,c9133,c4152,c3260,c1176,c1115,c2120,c246,c6213,c887,c9101,c0205,c333,c4248,c397,c731,c049,c517,c494,c7156,c3155,c7171,c783,c8192,c799,c720,c770,c6132,c6206,c4256,c399,c7289,c083,c9186,c7198,c815,c3251,c159,c3230,c711,c4179,c3110,c9169,c3254,c4263,c773,c2273,c8102,c848,c7116,c8293,c5195,c268,c1104,c7195,c3219,c4218,c069,c081,c099,c549,c9280,c8170,c5254,c2282,c6180,c5296,c020,c9264,c7151,c2237,c024,c4283,c558,c3131,c477,c5154,c80,c8259,c6266,c2179,c3227,c8130,c543,c7290,c579,c2264,c8143,c7166,c973,c6294,c5216,c6285,c486,c7144,c336,c7159,c891,c41,c3138,c2102,c7174,c689,c3146,c673,c9235,c2299,c981,c0199,c6237,c1181,c5169,c8272,c182,c2212,c5267,c6255,c254,c1128,c9267,c0232,c30,c4241,c633,c8113,c6263,c337,c6235,c9117,c034,c2241,c396,c3253,c6157,c6165,c1249,c5167,c4284,c111,c3108,c8175,c4291,c7228,c4171,c8289,c9221,c5152,c7263,c541,c679,c4282,c7237,c154,c155,c4221,c1159,c249,c0227,c81,c138,c9157,c0183,c8145,c498,c2151,c4153,c444,c9132,c315,c1184,c0272,c172,c5159,c2195,c6297,c6247,c499,c0247,c6299,c6286,c0106,c143,c1231,c9104,c2211,c0273,c671,c2136,c7250,c030,c247,c665,c3255,c3112,c0138,c619,c4259,c0286,c733,c8140,c5219,c1214,c9295,c6245,c9131,c5231,c3202,c2162,c6162,c6225,c052,c2214,c7249,c453,c919,c610,c293,c413,c8137,c465,c8299,c5228,c4147,c4138,c1123,c2156,c8231,c817,c918,c075,c5127,c2295,c1119,c4112,c4194,c175,c7104,c5257,c6172,c740,c6161,c147,c667,c366,c1276,c4117,c515,c7131,c0243,c090,c2114,c345,c244,c5189,c7197,c1172,c290,c7275,c0179,c2141,c121,c4170,c5108,c6202,c2204,c3218,c0146,c07,c1216,c213,c9217,c7119,c6244,c8114,c555,c1109,c1124,c1107,c5105,c56,c0110,c157,c4210,c9255,c550,c716,c0160,c124,c0189,c4130,c915,c044,c697,c917,c5172,c5113,c194,c4254,c8255,c669,c2198,c1133,c530,c127,c627,c1145,c219,c4236,c954,c9140,c146,c3250,c830,c2131,c2286,c0240,c993,c0155,c1175,c0214,c5181,c5182,c637,c3101,c0248,c6123,c0256,c6164,c8116,c8144,c0268,c0120,c2266,c8257,c7260,c652,c8126,c6230,c3194,c7127,c2298,c094,c1118,c5128,c0172,c432,c0237,c1135,c476,c7132,c6214,c881,c2121,c3228,c721,c7293,c3120,c040,c7191,c3199,c0202,c1164,c1153,c224,c4143,c926,c940,c342,c6216,c376,c6109,c0167,c1138,c790,c6145,c4240,c4118,c6148,c9178,c1179,c9245,c4177,c4183,c242,c974,c043,c529,c237,c6119,c1265,c2280,c0263,c6269,c883,c8153,c292,c221,c5266,c270,c514,c7175,c0295,c7224,c046,c1210,c24,c2185,c4243,c983,c8136,c0198,c9298,c324,c0145,c4281,c7122,c2160,c9149,c144,c7152,c478,c765,c9161,c360,c4195,c4142,c34,c0171,c36,c5125,c2106,c5226,c518,c5143,c681,c243,c0221,c15,c32,c4209,c0244,c9142,c3289,c578,c818,c4113,c72,c3268,c911,c958,c9289,c8208,c8148,c5206,c769,c7209,c8132,c540,c1220,c1131,c9274,c3258,c9166,c631,c837,c8251,c1147,c6155,c5145,c4120,c1280,c381,c9283,c3105,c754,c0228,c825,c812,c2203,c980,c2235,c380,c343,c5134,c7259,c846,c3256,c971,c1137,c3221,c4122,c8262,c066,c3210,c6199,c1171,c2250,c463,c9138,c1187,c7192,c8239,c3252,c9254,c1260,c9110,c372,c9278,c1268,c364,c70,c7143,c4192,c7113,c346,c061,c5280,c0280,c0212,c7186,c264,c2239,c9272,c0140,c4220,c5258,c6184,c1148,c231,c7278,c095,c8268,c8278,c666,c3187,c5220,c876,c76,c2197,c856,c736,c9215,c233,c1146,c074,c0251,c1177,c2157,c7253,c1163,c5208,c5165,c7298,c4144,c9134,c0123,c9129,c9143,c4163,c2253,c7129,c8162,c2147,c467,c439,c1258,c225,c3106,c4100,c889,c7182,c1191,c4133,c131,c7190,c859,c9260,c0164,c7161,c642,c0143,c9240,c743,c2272,c4234,c296,c1223,c2247,c1125,c2242,c8186,c9282,c762,c4186,c9109,c5249,c852,c979,c445,c810,c8236,c8253,c0121,c0192,c0258,c0287,c9168,c6120,c8154,c6293,c289,c6127,c0296,c4151,c8207,c4279,c62,c222,c2189,c695,c0291,c065,c3238,c4146,c7125,c2171,c749,c3224,c5166,c9118,c4228,c398,c064,c9182,c9287,c3235,c8280,c9238,c894,c7126,c6168,c0102,c4154,c7123,c947,c291,c4136,c1235,c33,c226,c2133,c6144,c655,c9266,c2125,c9247,c078,c0134,c729,c4175,c1103,c1156,c9258,c532,c516,c8178,c5141,c1273,c9211,c7218,c314,c634,c6289,c978,c4131,c6134,c923,c0211,c4285,c0111,c7106,c5112,c9159,c1110,c688,c1102,c267,c067,c4196,c0101,c1267,c1143,c7254,c17,c780,c8169,c5212,c2269,c1227,c4229,c18,c0225,c497,c0142,c4258,c524,c390,c3263,c0152,c437,c5173,c767,c276,c855,c2182,c014,c6188,c367,c041,c776,c4286,c8227,c1286,c449,c09,c1275,c5221,c278,c6219,c755,c843,c113,c036,c5118,c7208,c1222,c8283,c6114,c0226,c2285,c9218,c9176,c187,c3287,c941,c6112,c4295,c3284,c2210,c2206,c9249,c990,c5276,c845,c886,c534,c4245,c196,c4246,c3270,c71,c6287,c880,c8237,c3249,c8205,c5184,c258,c3116,c6102,c7282,c0104,c0266,c3141,c7236,c7148,c539,c184,c1136,c482,c8139,c3207,c22,c0180,c7294,c819,c417,c618,c6256,c6196,c582,c6250,c5131,c6186,c6274,c3267,c9226,c316,c4201,c7137,c4250,c00,c8181,c647,c3129,c5136,c5290,c6159,c9170,c6231,c1277,c3121,c7283,c350,c0210,c263,c1228,c4165,c1168,c8198,c4184,c132,c2275,c9126,c6221,c7269,c1196,c860,c9185,c9116,c3286,c8211,c5291,c2288,c3100,c1162,c698,c5248,c0252,c0153,c4185,c692,c7162,c7295,c8287,c3197,c936,c6110,c847,c9299,c7140,c271,c1201,c5234,c125,c3166,c310,c027,c3292,c3220,c5229,c8133,c013,c338,c21,c355,c794,c5110,c4230,c564,c2100,c751,c8275,c7142,c862,c0255,c8146,c2265,c4124,c063,c1120,c4267,c8177,c53,c97,c423,c5297,c330,c4125,c83,c3165,c37,c193,c58,c1182,c7272,c0246,c8134,c227,c4168,c7248,c7167,c8163,c4290,c628,c967,c3266,c3143,c3276,c895,c332,c2153,c8206,c0162,c4104,c6209,c03,c2257,c6220,c9137,c2193,c0250,c7141,c0109,c4174,c4188,c0129,c913,c0191,c322,c1204,c1255,c632,c912,c925,c5210,c527,c635,c8244,c0168,c084,c3188,c0150,c452,c8123,c42,c340,c188,c566,c1207,c433,c5147,c7187,c8220,c942,c7265,c3298,c2262,c7220,c5288,c485,c531,c388,c9244,c176,c6290,c6222,c0118,c759,c587,c5217,c7165,c839,c230,c011,c149,c7150,c05,c160,c1297,c730,c4297,c5289,c8138,c174,c5148,c9228,c3160,c1259,c4294,c148,c8274,c250,c575,c436,c1209,c2158,c3186,c4141,c6116,c7292,c4166,c8103,c7262,c0116,c982,c2117,c3265,c2196,c968,c9261,c0259,c441,c096,c2105,c3150,c471,c9285,c3240,c727,c2256,c7232,c872,c039,c9293,c248,c976,c513,c898,c2287,c5144,c8115,c010,c9277,c5250,c5287,c3102,c2254,c552,c7256,c617,c7189,c2137,c9263,c914,c6118,c6100,c2103,c916,c4110,c7245,c161,c012,c4202,c1274,c1185,c1285,c3167,c7251,c8223,c1183,c6133,c50,c7100,c0281,c7281,c1298,c7273,c9233,c943,c370,c4274,c6291,c468,c5299,c699,c2227,c238,c6131,c298,c140,c5121,c8249,c5163,c8155,c9248,c2155,c3162,c2172,c2258,c1160,c5256,c654,c8109,c9181,c1173,c3133,c3164,c63,c576,c9127,c8188,c134,c0288,c6260,c6194,c7230,c9202,c312,c797,c0139,c5203,c047,c472,c2276,c7233,c9196,c0108,c8128,c9197,c2104,c1288,c3154,c2101,c586,c5157,c2251,c6198,c774,c5197,c2148,c6111,c1294,c945,c6267,c8213,c54,c4108,c117,c5191,c828,c823,c3223,c3170,c284,c5102,c8110,c2233,c9173,c2278,c1100,c3214,c2268,c9207,c991,c4149,c1194,c457,c5137,c2289,c7206,c8166,c5239,c3118,c568,c2224,c2236,c294,c8281,c9225,c14,c1287,c994,c29,c6179,c1212,c283,c5233,c5200,c893,c756,c0105,c3239,c051,c7101,c8141,c487,c6268,c3124,c764,c5263,c865,c5270,c630,c6284,c6207,c261,c5101,c3109,c3169,c4116,c3225,c82,c8229,c6264,c9189,c525,c5238,c7146,c60,c3226,c5282,c6171,c431,c2108,c650,c4140,c4200,c4169,c746,c684,c2294,c5259,c6177,c4276,c556,c7242,c826,c320,c4198,c9246,c0148,c8185,c098,c0128,c8250,c329,c592,c9241,c253,c884,c2249,c391,c5120,c141,c8180,c4203,c7229,c8168,c584,c9122,c3201,c085,c653,c0158,c952,c6258,c8233,c74,c384,c4280,c6277,c1218,c5213,c7103,c3217,c8142,c8105,c0100,c0230,c5107,c3174,c972,c6163,c7226,c2145,c868,c2139,c1296,c04,c659,c168,c9270,c5178,c285,c6108,c5222,c7202,c8218,c9155,c4132,c6234,c3293,c4193,c7240,c3261,c425,c4231,c5214,c723,c4213,c0253,c2150,c5180,c6129,c6136,c49,c490,c4219,c8120,c8273,c1206,c3184,c5186,c772,c164,c8258,c4268,c0194,c4255,c0257,c395,c06,c572,c1197,c2234,c5199,c5224,c636,c9113,c9193,c033,c6200,c4225,c7285,c7291,c4150,c658,c092,c662,c032,c178,c5177,c026,c0275,c045,c1272,c1105,c8158,c9276,c8129,c2138,c888,c0119,c5161,c5117,c323,c4208,c871,c6169,c8247,c7223,c2167,c5285,c5284,c7176,c2129,c286,c1282,c929,c6239,c6279,c7277,c1150,c6272,c7169,c0165,c5207,c47,c325,c1299,c491,c5179,c2128,c028,c612,c3269,c0289,c1290,c5283,c2205,c120,c9206,c4232,c7133,c8245,c163,c789,c0186,c0157,c5156,c4159,c1134,c1217,c6228,c827,c428,c5241,c646,c448,c574,c766,c8260,c3299,c6190,c5293,c299,c6106,c1224,c3153,c6261,c26,c6142,c6223,c7241,c079,c1132,c6233,c2277,c8122,c9188,c158,c4251,c712,c260,c577,c1170,c3190,c6288,c3103,c474,c9296,c275,c1284,c6183,c897,c6193,c738,c84,c5260,c169,c5116,c2252,c495,c1202,c2110,c3203,c2245,c596,c2130,c9251,c824,c8157,c710,c742,c844,c4139,c7111,c7207,c687,c334,c3297,c724,c416,c5100,c6257,c2119,c5190,c3242,c9290,c0207,c1111,c4180,c6126,c1261,c8187,c3113,c8107,c877,c3137,c1278,c060,c5103,c616,c0147,c537,c7216,c2192,c0188,c8193,c8173,c999,c4199,c5109,c6154,c412,c7297,c7177,c435,c475,c8112,c0204,c8214,c426,c99,c6156,c029,c4189,c9112,c8199,c0265,c7213,c9146,c4277,c3205,c3272,c7120,c0219,c8204,c2132,c1112,c4260,c3206,c9102,c265,c257,c2217,c331,c3180,c0262,c5261,c2248,c9179,c2168,c9200,c1213,c0254,c7185,c6182,c3196,c2229,c8285,c622,c985,c7200,c8209,c7204,c9174,c955,c1248,c8203,c480,c2199,c9214,c5183,c3237,c663,c9108,c3168,c9195,c714,c2113,c7118,c9286,c2271,c0151,c2118,c718,c7212,c9130,c6218,c9223,c31,c96,c311,c277,c6167,c561,c760,c6253,c0175,c0190,c1247,c5236,c0264,c833,c1221,c9239,c682,c0113,c156,c966,c8200,c8164,c571,c5132,c0173,c251,c2159,c4217,c732,c691,c7109,c461,c7135,c2260,c1151,c056,c4292,c726,c9139,c6204,c3273,c8106,c11,c6103,c8125,c1246,c8254,c7227,c8201,c4296,c5204,c8286,c3104,c40,c6141,c133,c45,c2226,c717,c5298,c7246,c8127,c281,c2270,c0213,c8167,c086,c3264,c5272,c1291,c454,c9222,c2146,c6121,c5245,c3191,c1114,c7210,c4233,c8242,c588,c6249,c019,c0271,c7299,c79,c849,c1117,c198,c570,c2246,c778,c3232,c0126,c9141,c3248,c563,c542,c10,c0130,c2190,c928,c930,c8265,c362,c3145,c8246,c5211,c8222,c8226,c9288,c6146,c6210,c2107,c3192,c328,c9220,c7271,c2135,c597,c7219,c675,c8294,c1270,c4288,c4157,c5209,c838,c9172,c7160,c7172,c374,c963,c4257,c511,c768,c2231,c4252,c569,c01,c042,c885,c9187,c585,c496,c162,c7170,c183,c8279,c3189,c9257,c949,c829,c2255,c3122,c1141,c8269,c950,c5192,c0159,c0141,c6191,c9209,c1205,c462,c8190,c4101,c8284,c9227,c0278,c48,c6143,c443,c4299,c3244,c110,c9103,c082,c269,c6212,c9184,c2230,c266,c5275,c763,c0285,c4181,c7222,c3246,c5198,c560,c5124,c0163,c5174,c421,c9203,c1256,c438,c567,c744,c3158,c3176,c89,c7267,c8282,c352,c4191,c0233,c6203,c735,c488,c8117,c4172,c782,c215,c5138,c7217,c713,c0187,c7288,c5135,c236,c6251,c1254,c595,c9213,c0208,c1241,c2244,c94,c961,c0239,c739,c181,c44,c6236,c3234,c599,c3231,c3277,c9250,c798,c7296,c7139,c5104,c0223,c135,c3195,c025,c089,c1243,c644,c363,c229,c093,c5130,c8228,c3211,c5133,c640,c613,c9144,c3283,c750,c8235,c6181,c015,c359,c672,c8225,c696,c7136,c9275,c822,c6152,c4173,c7128,c2175,c9232,c4244,c758,c3135,c2218,c430,c535,c28,c3181,c67,c4197,c670,c995,c339,c5196,c9136,c1263,c6197,c5277,c2176,c3136,c038,c351,c4121,c5205,c4190,c562,c7179,c424,c1167,c2170,c2184,c5188,c389,c3175,c1240,c411,c7257,c8296,c4114,c241,c1190,c4111,c4269,c097,c536,c5106,c456,c1169,c4155,c57,c6138,c152,c6270,c922,c0269,c361,c6140,c78,c580,c0279,c0182,c0181,c3173,c3134,c590,c20,c1189,c3257,c4287,c414,c9262,c6115,c1238,c8165,c2144,c944,c5194,c1158,c6295,c741,c2124,c2208,c2284,c3280,c5252,c3107,c6281,c989,c2177,c0156,c9115,c386,c7199,c8179,c6240,c2290,c9230,c8232,c130,c6187,c6232,c2164,c9234,c840,c6122,c834,c987,c055,c234,c1122,c223,c0220,c123,c5153,c6283,c8108,c4272,c9242,c7196,c992,c965,c2188,c6282,c9111,c2225,c7276,c0206,c5185,c4167,c7112,c1139,c8215,c0125,c8152,c7231,c4212,c112,c1188,c9183,c195,c6229,c8266,c8151,c2126,c5273,c415,c8121,c996,c282,c86,c3171,c382,c6242,c16,c2127,c51,c65,c2173,c451,c2261,c9180,c9212,c85,c851,c4224,c6107,c8159,c9114,c853,c546,c385,c6192,c0294,c0235,c459,c8212,c4103,c3130,c8297,c8172,c3204,c9194,c0267,c1283,c1244,c1215,c777,c383,c167,c4265,c869,c2243,c8184,c287,c7274,c1129,c69,c017,c7117,c2202,c1149,c7115,c814,c5162,c779,c6217,c2143,c4264,c8216,c1234,c1211,c2291,c3151,c489,c858,c4214,c6280,c882,c7205,c8189,c0236,c379,c6150,c5122,c4135,c7158,c878,c068,c0185,c1152,c3222,c5158,c795,c9268,c197,c319,c988,c1250,c393,c2219,c1292,c8147,c9198,c1237,c2165,c053,c256,c3179,c5151,c9271,c796,c92,c129,c5149,c418,c676,c614,c7181,c9192,c4162,c4215,c8131,c7252,c3275,c0261,c8238,c5202,c890,c5139,c581,c434,c9273,c6246,c3198,c551,c3144,c02,c565,c073,c8171,c4275,c136,c61,c7183,c8217,c1157,c326,c3185,c757,c7107,c5262,c573,c3285,c7261,c4262,c7194,c466,c9163,c2115,c5114,c228,c523,c5235,c761,c787,c59,c5247,c9279,c5230,c021,c317,c354,c2274,c6226,c522,c7239,c3290,c4278,c341,c0242,c151,c728,c7153,c639,c3149,c037,c2267,c091,c9224,c6185,c0200,c1108,c7258,c8256,c274,c8252,c9210,c553,c648,c850,c7284,c0282,c842,c5123,c781,c998,c8101,c784,c9231,c3296,c2109,c245,c022,c8261,c273,c1101,c2186,c6104,c3262,c959,c2194,c2296,c3288,c128,c870,c8135,c921,c6117,c831,c8298,c8271,c6139,c694,c1289,c072,c3247,c8210,c8234,c410,c7178,c6176,c775,c059,c080,c118,c1165,c4227,c510,c9152,c641,c593,c984,c6211,c854,c1208,c1126,c6124,c8124,c8197,c975,c5242,c6160,c4158,c8240,c9153,c7193,c7215,c9259,c077,c2279,c3178,c4105,c9160,c429,c6175,c9284,c8230,c863,c235,c821,c951,c9291,c5227,c4176,c8241,c657 );

input x0;
input x1;
input x2;
input x3;
input x4;
input x5;
input x6;
input x7;
input x8;
input x9;
input x10;
input x11;
input x12;
input x13;
input x14;
input x15;
input x16;
input x17;
input x18;
input x19;
input x20;
input x21;
input x22;
input x23;
input x24;
input x25;
input x26;
input x27;
input x28;
input x29;
input x30;
input x31;
input x32;
input x33;
input x34;
input x35;
input x36;
input x37;
input x38;
input x39;
input x40;
input x41;
input x42;
input x43;
input x44;
input x45;
input x46;
input x47;
input x48;
input x49;
input x50;
input x51;
input x52;
input x53;
input x54;
input x55;
input x56;
input x57;
input x58;
input x59;
input x60;
input x61;
input x62;
input x63;
input x64;
input x65;
input x66;
input x67;
input x68;
input x69;
input x70;
input x71;
input x72;
input x73;
input x74;
input x75;
input x76;
input x77;
input x78;
input x79;
input x80;
input x81;
input x82;
input x83;
input x84;
input x85;
input x86;
input x87;
input x88;
input x89;
input x90;
input x91;
input x92;
input x93;
input x94;
input x95;
input x96;
input x97;
input x98;
input x99;
input x100;
input x101;
input x102;
input x103;
input x104;
input x105;
input x106;
input x107;
input x108;
input x109;
input x110;
input x111;
input x112;
input x113;
input x114;
input x115;
input x116;
input x117;
input x118;
input x119;
input x120;
input x121;
input x122;
input x123;
input x124;
input x125;
input x126;
input x127;
input x128;
input x129;
input x130;
input x131;
input x132;
input x133;
input x134;
input x135;
input x136;
input x137;
input x138;
input x139;
input x140;
input x141;
input x142;
input x143;
input x144;
input x145;
input x146;
input x147;
input x148;
input x149;
input x150;
input x151;
input x152;
input x153;
input x154;
input x155;
input x156;
input x157;
input x158;
input x159;
input x160;
input x161;
input x162;
input x163;
input x164;
input x165;
input x166;
input x167;
input x168;
input x169;
input x170;
input x171;
input x172;
input x173;
input x174;
input x175;
input x176;
input x177;
input x178;
input x179;
input x180;
input x181;
input x182;
input x183;
input x184;
input x185;
input x186;
input x187;
input x188;
input x189;
input x190;
input x191;
input x192;
input x193;
input x194;
input x195;
input x196;
input x197;
input x198;
input x199;
input x200;
input x201;
input x202;
input x203;
input x204;
input x205;
input x206;
input x207;
input x208;
input x209;
input x210;
input x211;
input x212;
input x213;
input x214;
input x215;
input x216;
input x217;
input x218;
input x219;
input x220;
input x221;
input x222;
input x223;
input x224;
input x225;
input x226;
input x227;
input x228;
input x229;
input x230;
input x231;
input x232;
input x233;
input x234;
input x235;
input x236;
input x237;
input x238;
input x239;
input x240;
input x241;
input x242;
input x243;
input x244;
input x245;
input x246;
input x247;
input x248;
input x249;
input x250;
input x251;
input x252;
input x253;
input x254;
input x255;
input x256;
input x257;
input x258;
input x259;
input x260;
input x261;
input x262;
input x263;
input x264;
input x265;
input x266;
input x267;
input x268;
input x269;
input x270;
input x271;
input x272;
input x273;
input x274;
input x275;
input x276;
input x277;
input x278;
input x279;
input x280;
input x281;
input x282;
input x283;
input x284;
input x285;
input x286;
input x287;
input x288;
input x289;
input x290;
input x291;
input x292;
input x293;
input x294;
input x295;
input x296;
input x297;
input x298;
input x299;
input x300;
input x301;
input x302;
input x303;
input x304;
input x305;
input x306;
input x307;
input x308;
input x309;
input x310;
input x311;
input x312;
input x313;
input x314;
input x315;
input x316;
input x317;
input x318;
input x319;
input x320;
input x321;
input x322;
input x323;
input x324;
input x325;
input x326;
input x327;
input x328;
input x329;
input x330;
input x331;
input x332;
input x333;
input x334;
input x335;
input x336;
input x337;
input x338;
input x339;
input x340;
input x341;
input x342;
input x343;
input x344;
input x345;
input x346;
input x347;
input x348;
input x349;
input x350;
input x351;
input x352;
input x353;
input x354;
input x355;
input x356;
input x357;
input x358;
input x359;
input x360;
input x361;
input x362;
input x363;
input x364;
input x365;
input x366;
input x367;
input x368;
input x369;
input x370;
input x371;
input x372;
input x373;
input x374;
input x375;
input x376;
input x377;
input x378;
input x379;
input x380;
input x381;
input x382;
input x383;
input x384;
input x385;
input x386;
input x387;
input x388;
input x389;
input x390;
input x391;
input x392;
input x393;
input x394;
input x395;
input x396;
input x397;
input x398;
input x399;
input x400;
input x401;
input x402;
input x403;
input x404;
input x405;
input x406;
input x407;
input x408;
input x409;
input x410;
input x411;
input x412;
input x413;
input x414;
input x415;
input x416;
input x417;
input x418;
input x419;
input x420;
input x421;
input x422;
input x423;
input x424;
input x425;
input x426;
input x427;
input x428;
input x429;
input x430;
input x431;
input x432;
input x433;
input x434;
input x435;
input x436;
input x437;
input x438;
input x439;
input x440;
input x441;
input x442;
input x443;
input x444;
input x445;
input x446;
input x447;
input x448;
input x449;
input x450;
input x451;
input x452;
input x453;
input x454;
input x455;
input x456;
input x457;
input x458;
input x459;
input x460;
input x461;
input x462;
input x463;
input x464;
input x465;
input x466;
input x467;
input x468;
input x469;
input x470;
input x471;
input x472;
input x473;
input x474;
input x475;
input x476;
input x477;
input x478;
input x479;
input x480;
input x481;
input x482;
input x483;
input x484;
input x485;
input x486;
input x487;
input x488;
input x489;
input x490;
input x491;
input x492;
input x493;
input x494;
input x495;
input x496;
input x497;
input x498;
input x499;
input x500;
input x501;
input x502;
input x503;
input x504;
input x505;
input x506;
input x507;
input x508;
input x509;
input x510;
input x511;
input x512;
input x513;
input x514;
input x515;
input x516;
input x517;
input x518;
input x519;
input x520;
input x521;
input x522;
input x523;
input x524;
input x525;
input x526;
input x527;
input x528;
input x529;
input x530;
input x531;
input x532;
input x533;
input x534;
input x535;
input x536;
input x537;
input x538;
input x539;
input x540;
input x541;
input x542;
input x543;
input x544;
input x545;
input x546;
input x547;
input x548;
input x549;
input x550;
input x551;
input x552;
input x553;
input x554;
input x555;
input x556;
input x557;
input x558;
input x559;
input x560;
input x561;
input x562;
input x563;
input x564;
input x565;
input x566;
input x567;
input x568;
input x569;
input x570;
input x571;
input x572;
input x573;
input x574;
input x575;
input x576;
input x577;
input x578;
input x579;
input x580;
input x581;
input x582;
input x583;
input x584;
input x585;
input x586;
input x587;
input x588;
input x589;
input x590;
input x591;
input x592;
input x593;
input x594;
input x595;
input x596;
input x597;
input x598;
input x599;
input x600;
input x601;
input x602;
input x603;
input x604;
input x605;
input x606;
input x607;
input x608;
input x609;
input x610;
input x611;
input x612;
input x613;
input x614;
input x615;
input x616;
input x617;
input x618;
input x619;
input x620;
input x621;
input x622;
input x623;
input x624;
input x625;
input x626;
input x627;
input x628;
input x629;
input x630;
input x631;
input x632;
input x633;
input x634;
input x635;
input x636;
input x637;
input x638;
input x639;
input x640;
input x641;
input x642;
input x643;
input x644;
input x645;
input x646;
input x647;
input x648;
input x649;
input x650;
input x651;
input x652;
input x653;
input x654;
input x655;
input x656;
input x657;
input x658;
input x659;
input x660;
input x661;
input x662;
input x663;
input x664;
input x665;
input x666;
input x667;
input x668;
input x669;
input x670;
input x671;
input x672;
input x673;
input x674;
input x675;
input x676;
input x677;
input x678;
input x679;
input x680;
input x681;
input x682;
input x683;
input x684;
input x685;
input x686;
input x687;
input x688;
input x689;
input x690;
input x691;
input x692;
input x693;
input x694;
input x695;
input x696;
input x697;
input x698;
input x699;
input x700;
input x701;
input x702;
input x703;
input x704;
input x705;
input x706;
input x707;
input x708;
input x709;
input x710;
input x711;
input x712;
input x713;
input x714;
input x715;
input x716;
input x717;
input x718;
input x719;
input x720;
input x721;
input x722;
input x723;
input x724;
input x725;
input x726;
input x727;
input x728;
input x729;
input x730;
input x731;
input x732;
input x733;
input x734;
input x735;
input x736;
input x737;
input x738;
input x739;
input x740;
input x741;
input x742;
input x743;
input x744;
input x745;
input x746;
input x747;
input x748;
input x749;
input x750;
input x751;
input x752;
input x753;
input x754;
input x755;
input x756;
input x757;
input x758;
input x759;
input x760;
input x761;
input x762;
input x763;
input x764;
input x765;
input x766;
input x767;
input x768;
input x769;
input x770;
input x771;
input x772;
input x773;
input x774;
input x775;
input x776;
input x777;
input x778;
input x779;
input x780;
input x781;
input x782;
input x783;
output c38;
output c6296;
output c8194;
output c0144;
output c7168;
output c3161;
output c623;
output c08;
output c050;
output c753;
output c239;
output c062;
output c3123;
output c962;
output c177;
output c2209;
output c9294;
output c93;
output c392;
output c4137;
output c5193;
output c122;
output c0170;
output c1199;
output c1279;
output c0290;
output c3163;
output c35;
output c2213;
output c0161;
output c4237;
output c8277;
output c875;
output c199;
output c139;
output c6208;
output c3271;
output c0201;
output c6271;
output c4182;
output c0209;
output c0193;
output c387;
output c7243;
output c924;
output c7108;
output c3117;
output c91;
output c9199;
output c6105;
output c957;
output c5244;
output c7221;
output c932;
output c9119;
output c8202;
output c771;
output c1121;
output c9156;
output c685;
output c470;
output c378;
output c180;
output c6174;
output c295;
output c365;
output c137;
output c5253;
output c9158;
output c5278;
output c179;
output c0231;
output c4145;
output c946;
output c5225;
output c5246;
output c9265;
output c626;
output c4129;
output c0124;
output c2216;
output c6278;
output c447;
output c2174;
output c5243;
output c6128;
output c5223;
output c255;
output c6195;
output c190;
output c469;
output c95;
output c2183;
output c4271;
output c357;
output c664;
output c791;
output c9120;
output c3233;
output c2166;
output c9219;
output c938;
output c785;
output c4115;
output c2223;
output c651;
output c899;
output c0135;
output c0224;
output c6298;
output c0154;
output c1239;
output c4242;
output c0292;
output c9128;
output c920;
output c484;
output c4204;
output c8104;
output c0293;
output c2221;
output c5129;
output c0277;
output c5281;
output c5292;
output c5265;
output c7244;
output c836;
output c960;
output c191;
output c874;
output c9148;
output c1264;
output c8119;
output c7130;
output c0270;
output c6215;
output c0133;
output c2181;
output c9297;
output c7270;
output c935;
output c0178;
output c0299;
output c3159;
output c5115;
output c8191;
output c816;
output c114;
output c6149;
output c450;
output c4222;
output c27;
output c1293;
output c210;
output c1186;
output c344;
output c5286;
output c9125;
output c4235;
output c377;
output c6224;
output c6205;
output c8195;
output c070;
output c7235;
output c3142;
output c5119;
output c1195;
output c5255;
output c2142;
output c4206;
output c8295;
output c5170;
output c2292;
output c6135;
output c321;
output c5240;
output c2180;
output c4134;
output c554;
output c1242;
output c1193;
output c252;
output c3126;
output c481;
output c214;
output c5111;
output c1252;
output c2293;
output c493;
output c218;
output c5126;
output c620;
output c0197;
output c2191;
output c1166;
output c7203;
output c8156;
output c788;
output c937;
output c956;
output c2111;
output c7163;
output c3147;
output c9208;
output c1269;
output c2201;
output c4223;
output c318;
output c545;
output c832;
output c3152;
output c4226;
output c3241;
output c0166;
output c3208;
output c1180;
output c2154;
output c970;
output c358;
output c3209;
output c0137;
output c5175;
output c9177;
output c1271;
output c811;
output c1203;
output c548;
output c6147;
output c8243;
output c0216;
output c9124;
output c349;
output c1236;
output c4107;
output c7214;
output c7266;
output c864;
output c9201;
output c656;
output c1161;
output c4266;
output c645;
output c7134;
output c0284;
output c7264;
output c3243;
output c9190;
output c2207;
output c5264;
output c683;
output c9269;
output c9204;
output c5155;
output c77;
output c2187;
output c076;
output c0297;
output c1245;
output c1174;
output c3128;
output c7157;
output c910;
output c166;
output c953;
output c8267;
output c896;
output c1140;
output c13;
output c87;
output c272;
output c1155;
output c427;
output c611;
output c0229;
output c6189;
output c4126;
output c559;
output c297;
output c8111;
output c9252;
output c0127;
output c212;
output c262;
output c8248;
output c016;
output c23;
output c66;
output c674;
output c939;
output c977;
output c0234;
output c9135;
output c2297;
output c591;
output c3193;
output c087;
output c7268;
output c7180;
output c9205;
output c9150;
output c1154;
output c12;
output c3279;
output c216;
output c690;
output c715;
output c9292;
output c6153;
output c368;
output c3212;
output c5237;
output c9253;
output c115;
output c5251;
output c519;
output c5168;
output c211;
output c0245;
output c6265;
output c347;
output c615;
output c693;
output c0276;
output c3182;
output c170;
output c0149;
output c142;
output c3215;
output c4207;
output c3127;
output c2149;
output c464;
output c538;
output c446;
output c9145;
output c933;
output c7138;
output c0184;
output c9175;
output c7121;
output c2215;
output c442;
output c931;
output c0174;
output c7247;
output c39;
output c7155;
output c348;
output c088;
output c116;
output c598;
output c3291;
output c4211;
output c52;
output c5232;
output c9151;
output c0195;
output c023;
output c661;
output c512;
output c747;
output c5146;
output c1226;
output c2259;
output c054;
output c1200;
output c4148;
output c6130;
output c677;
output c6273;
output c725;
output c98;
output c46;
output c7286;
output c9105;
output c3216;
output c9164;
output c25;
output c217;
output c2169;
output c1232;
output c9154;
output c4247;
output c1144;
output c1251;
output c1257;
output c9107;
output c335;
output c7145;
output c057;
output c533;
output c927;
output c0114;
output c0132;
output c737;
output c4273;
output c440;
output c589;
output c792;
output c4289;
output c8219;
output c8291;
output c3148;
output c9237;
output c6113;
output c7105;
output c813;
output c0217;
output c4109;
output c90;
output c6252;
output c394;
output c520;
output c7225;
output c43;
output c0122;
output c3282;
output c7147;
output c327;
output c6248;
output c369;
output c165;
output c4205;
output c9243;
output c892;
output c6158;
output c3111;
output c0176;
output c3295;
output c6173;
output c528;
output c232;
output c9100;
output c071;
output c0177;
output c9216;
output c7154;
output c3281;
output c547;
output c793;
output c0222;
output c6125;
output c6241;
output c624;
output c3229;
output c680;
output c8160;
output c1230;
output c5201;
output c1142;
output c526;
output c126;
output c7280;
output c861;
output c4239;
output c7279;
output c5142;
output c7184;
output c8174;
output c8176;
output c734;
output c7287;
output c820;
output c9165;
output c280;
output c279;
output c8161;
output c2122;
output c6170;
output c19;
output c3139;
output c185;
output c2281;
output c4270;
output c2152;
output c3177;
output c5171;
output c0238;
output c035;
output c0117;
output c722;
output c8221;
output c73;
output c879;
output c150;
output c7102;
output c6276;
output c0131;
output c6254;
output c948;
output c058;
output c0215;
output c2283;
output c2200;
output c3236;
output c5271;
output c873;
output c8270;
output c3140;
output c492;
output c2222;
output c4298;
output c68;
output c0196;
output c969;
output c483;
output c5176;
output c5295;
output c8288;
output c1281;
output c997;
output c192;
output c018;
output c3294;
output c0283;
output c455;
output c2123;
output c189;
output c4128;
output c668;
output c8100;
output c173;
output c479;
output c638;
output c0241;
output c4119;
output c3115;
output c6259;
output c9121;
output c866;
output c521;
output c1106;
output c544;
output c1233;
output c3156;
output c8263;
output c422;
output c2134;
output c3245;
output c64;
output c3119;
output c0136;
output c0103;
output c7255;
output c048;
output c5274;
output c88;
output c419;
output c1178;
output c6151;
output c460;
output c9236;
output c6101;
output c2116;
output c0112;
output c5268;
output c4161;
output c0107;
output c6238;
output c0260;
output c5140;
output c5279;
output c621;
output c7110;
output c356;
output c8276;
output c3114;
output c678;
output c2178;
output c7164;
output c2238;
output c5150;
output c7124;
output c1116;
output c313;
output c8183;
output c3183;
output c2240;
output c4261;
output c220;
output c2228;
output c4249;
output c7173;
output c6201;
output c3172;
output c375;
output c259;
output c1295;
output c3132;
output c1219;
output c3213;
output c373;
output c1130;
output c1192;
output c3157;
output c3259;
output c1262;
output c1225;
output c1229;
output c55;
output c9281;
output c8196;
output c8150;
output c4293;
output c75;
output c7201;
output c867;
output c473;
output c8149;
output c4216;
output c119;
output c8290;
output c986;
output c3125;
output c4106;
output c4178;
output c786;
output c6227;
output c9256;
output c4102;
output c0115;
output c9191;
output c8224;
output c171;
output c3200;
output c0298;
output c5294;
output c583;
output c9167;
output c0249;
output c557;
output c8264;
output c0218;
output c1113;
output c660;
output c7211;
output c649;
output c629;
output c0203;
output c857;
output c6137;
output c6178;
output c6166;
output c719;
output c594;
output c2140;
output c964;
output c2263;
output c1127;
output c9123;
output c2220;
output c5218;
output c6292;
output c934;
output c6243;
output c1198;
output c0169;
output c3274;
output c1266;
output c5269;
output c420;
output c7188;
output c7238;
output c2161;
output c8118;
output c7234;
output c9147;
output c5164;
output c8292;
output c4127;
output c5215;
output c0274;
output c7114;
output c4123;
output c288;
output c4156;
output c686;
output c6262;
output c9171;
output c371;
output c353;
output c031;
output c9106;
output c145;
output c4164;
output c745;
output c9162;
output c3278;
output c5160;
output c4187;
output c748;
output c2232;
output c841;
output c752;
output c153;
output c2163;
output c625;
output c835;
output c9229;
output c8182;
output c186;
output c1253;
output c240;
output c458;
output c4238;
output c5187;
output c643;
output c6275;
output c2112;
output c4160;
output c4253;
output c7149;
output c9133;
output c4152;
output c3260;
output c1176;
output c1115;
output c2120;
output c246;
output c6213;
output c887;
output c9101;
output c0205;
output c333;
output c4248;
output c397;
output c731;
output c049;
output c517;
output c494;
output c7156;
output c3155;
output c7171;
output c783;
output c8192;
output c799;
output c720;
output c770;
output c6132;
output c6206;
output c4256;
output c399;
output c7289;
output c083;
output c9186;
output c7198;
output c815;
output c3251;
output c159;
output c3230;
output c711;
output c4179;
output c3110;
output c9169;
output c3254;
output c4263;
output c773;
output c2273;
output c8102;
output c848;
output c7116;
output c8293;
output c5195;
output c268;
output c1104;
output c7195;
output c3219;
output c4218;
output c069;
output c081;
output c099;
output c549;
output c9280;
output c8170;
output c5254;
output c2282;
output c6180;
output c5296;
output c020;
output c9264;
output c7151;
output c2237;
output c024;
output c4283;
output c558;
output c3131;
output c477;
output c5154;
output c80;
output c8259;
output c6266;
output c2179;
output c3227;
output c8130;
output c543;
output c7290;
output c579;
output c2264;
output c8143;
output c7166;
output c973;
output c6294;
output c5216;
output c6285;
output c486;
output c7144;
output c336;
output c7159;
output c891;
output c41;
output c3138;
output c2102;
output c7174;
output c689;
output c3146;
output c673;
output c9235;
output c2299;
output c981;
output c0199;
output c6237;
output c1181;
output c5169;
output c8272;
output c182;
output c2212;
output c5267;
output c6255;
output c254;
output c1128;
output c9267;
output c0232;
output c30;
output c4241;
output c633;
output c8113;
output c6263;
output c337;
output c6235;
output c9117;
output c034;
output c2241;
output c396;
output c3253;
output c6157;
output c6165;
output c1249;
output c5167;
output c4284;
output c111;
output c3108;
output c8175;
output c4291;
output c7228;
output c4171;
output c8289;
output c9221;
output c5152;
output c7263;
output c541;
output c679;
output c4282;
output c7237;
output c154;
output c155;
output c4221;
output c1159;
output c249;
output c0227;
output c81;
output c138;
output c9157;
output c0183;
output c8145;
output c498;
output c2151;
output c4153;
output c444;
output c9132;
output c315;
output c1184;
output c0272;
output c172;
output c5159;
output c2195;
output c6297;
output c6247;
output c499;
output c0247;
output c6299;
output c6286;
output c0106;
output c143;
output c1231;
output c9104;
output c2211;
output c0273;
output c671;
output c2136;
output c7250;
output c030;
output c247;
output c665;
output c3255;
output c3112;
output c0138;
output c619;
output c4259;
output c0286;
output c733;
output c8140;
output c5219;
output c1214;
output c9295;
output c6245;
output c9131;
output c5231;
output c3202;
output c2162;
output c6162;
output c6225;
output c052;
output c2214;
output c7249;
output c453;
output c919;
output c610;
output c293;
output c413;
output c8137;
output c465;
output c8299;
output c5228;
output c4147;
output c4138;
output c1123;
output c2156;
output c8231;
output c817;
output c918;
output c075;
output c5127;
output c2295;
output c1119;
output c4112;
output c4194;
output c175;
output c7104;
output c5257;
output c6172;
output c740;
output c6161;
output c147;
output c667;
output c366;
output c1276;
output c4117;
output c515;
output c7131;
output c0243;
output c090;
output c2114;
output c345;
output c244;
output c5189;
output c7197;
output c1172;
output c290;
output c7275;
output c0179;
output c2141;
output c121;
output c4170;
output c5108;
output c6202;
output c2204;
output c3218;
output c0146;
output c07;
output c1216;
output c213;
output c9217;
output c7119;
output c6244;
output c8114;
output c555;
output c1109;
output c1124;
output c1107;
output c5105;
output c56;
output c0110;
output c157;
output c4210;
output c9255;
output c550;
output c716;
output c0160;
output c124;
output c0189;
output c4130;
output c915;
output c044;
output c697;
output c917;
output c5172;
output c5113;
output c194;
output c4254;
output c8255;
output c669;
output c2198;
output c1133;
output c530;
output c127;
output c627;
output c1145;
output c219;
output c4236;
output c954;
output c9140;
output c146;
output c3250;
output c830;
output c2131;
output c2286;
output c0240;
output c993;
output c0155;
output c1175;
output c0214;
output c5181;
output c5182;
output c637;
output c3101;
output c0248;
output c6123;
output c0256;
output c6164;
output c8116;
output c8144;
output c0268;
output c0120;
output c2266;
output c8257;
output c7260;
output c652;
output c8126;
output c6230;
output c3194;
output c7127;
output c2298;
output c094;
output c1118;
output c5128;
output c0172;
output c432;
output c0237;
output c1135;
output c476;
output c7132;
output c6214;
output c881;
output c2121;
output c3228;
output c721;
output c7293;
output c3120;
output c040;
output c7191;
output c3199;
output c0202;
output c1164;
output c1153;
output c224;
output c4143;
output c926;
output c940;
output c342;
output c6216;
output c376;
output c6109;
output c0167;
output c1138;
output c790;
output c6145;
output c4240;
output c4118;
output c6148;
output c9178;
output c1179;
output c9245;
output c4177;
output c4183;
output c242;
output c974;
output c043;
output c529;
output c237;
output c6119;
output c1265;
output c2280;
output c0263;
output c6269;
output c883;
output c8153;
output c292;
output c221;
output c5266;
output c270;
output c514;
output c7175;
output c0295;
output c7224;
output c046;
output c1210;
output c24;
output c2185;
output c4243;
output c983;
output c8136;
output c0198;
output c9298;
output c324;
output c0145;
output c4281;
output c7122;
output c2160;
output c9149;
output c144;
output c7152;
output c478;
output c765;
output c9161;
output c360;
output c4195;
output c4142;
output c34;
output c0171;
output c36;
output c5125;
output c2106;
output c5226;
output c518;
output c5143;
output c681;
output c243;
output c0221;
output c15;
output c32;
output c4209;
output c0244;
output c9142;
output c3289;
output c578;
output c818;
output c4113;
output c72;
output c3268;
output c911;
output c958;
output c9289;
output c8208;
output c8148;
output c5206;
output c769;
output c7209;
output c8132;
output c540;
output c1220;
output c1131;
output c9274;
output c3258;
output c9166;
output c631;
output c837;
output c8251;
output c1147;
output c6155;
output c5145;
output c4120;
output c1280;
output c381;
output c9283;
output c3105;
output c754;
output c0228;
output c825;
output c812;
output c2203;
output c980;
output c2235;
output c380;
output c343;
output c5134;
output c7259;
output c846;
output c3256;
output c971;
output c1137;
output c3221;
output c4122;
output c8262;
output c066;
output c3210;
output c6199;
output c1171;
output c2250;
output c463;
output c9138;
output c1187;
output c7192;
output c8239;
output c3252;
output c9254;
output c1260;
output c9110;
output c372;
output c9278;
output c1268;
output c364;
output c70;
output c7143;
output c4192;
output c7113;
output c346;
output c061;
output c5280;
output c0280;
output c0212;
output c7186;
output c264;
output c2239;
output c9272;
output c0140;
output c4220;
output c5258;
output c6184;
output c1148;
output c231;
output c7278;
output c095;
output c8268;
output c8278;
output c666;
output c3187;
output c5220;
output c876;
output c76;
output c2197;
output c856;
output c736;
output c9215;
output c233;
output c1146;
output c074;
output c0251;
output c1177;
output c2157;
output c7253;
output c1163;
output c5208;
output c5165;
output c7298;
output c4144;
output c9134;
output c0123;
output c9129;
output c9143;
output c4163;
output c2253;
output c7129;
output c8162;
output c2147;
output c467;
output c439;
output c1258;
output c225;
output c3106;
output c4100;
output c889;
output c7182;
output c1191;
output c4133;
output c131;
output c7190;
output c859;
output c9260;
output c0164;
output c7161;
output c642;
output c0143;
output c9240;
output c743;
output c2272;
output c4234;
output c296;
output c1223;
output c2247;
output c1125;
output c2242;
output c8186;
output c9282;
output c762;
output c4186;
output c9109;
output c5249;
output c852;
output c979;
output c445;
output c810;
output c8236;
output c8253;
output c0121;
output c0192;
output c0258;
output c0287;
output c9168;
output c6120;
output c8154;
output c6293;
output c289;
output c6127;
output c0296;
output c4151;
output c8207;
output c4279;
output c62;
output c222;
output c2189;
output c695;
output c0291;
output c065;
output c3238;
output c4146;
output c7125;
output c2171;
output c749;
output c3224;
output c5166;
output c9118;
output c4228;
output c398;
output c064;
output c9182;
output c9287;
output c3235;
output c8280;
output c9238;
output c894;
output c7126;
output c6168;
output c0102;
output c4154;
output c7123;
output c947;
output c291;
output c4136;
output c1235;
output c33;
output c226;
output c2133;
output c6144;
output c655;
output c9266;
output c2125;
output c9247;
output c078;
output c0134;
output c729;
output c4175;
output c1103;
output c1156;
output c9258;
output c532;
output c516;
output c8178;
output c5141;
output c1273;
output c9211;
output c7218;
output c314;
output c634;
output c6289;
output c978;
output c4131;
output c6134;
output c923;
output c0211;
output c4285;
output c0111;
output c7106;
output c5112;
output c9159;
output c1110;
output c688;
output c1102;
output c267;
output c067;
output c4196;
output c0101;
output c1267;
output c1143;
output c7254;
output c17;
output c780;
output c8169;
output c5212;
output c2269;
output c1227;
output c4229;
output c18;
output c0225;
output c497;
output c0142;
output c4258;
output c524;
output c390;
output c3263;
output c0152;
output c437;
output c5173;
output c767;
output c276;
output c855;
output c2182;
output c014;
output c6188;
output c367;
output c041;
output c776;
output c4286;
output c8227;
output c1286;
output c449;
output c09;
output c1275;
output c5221;
output c278;
output c6219;
output c755;
output c843;
output c113;
output c036;
output c5118;
output c7208;
output c1222;
output c8283;
output c6114;
output c0226;
output c2285;
output c9218;
output c9176;
output c187;
output c3287;
output c941;
output c6112;
output c4295;
output c3284;
output c2210;
output c2206;
output c9249;
output c990;
output c5276;
output c845;
output c886;
output c534;
output c4245;
output c196;
output c4246;
output c3270;
output c71;
output c6287;
output c880;
output c8237;
output c3249;
output c8205;
output c5184;
output c258;
output c3116;
output c6102;
output c7282;
output c0104;
output c0266;
output c3141;
output c7236;
output c7148;
output c539;
output c184;
output c1136;
output c482;
output c8139;
output c3207;
output c22;
output c0180;
output c7294;
output c819;
output c417;
output c618;
output c6256;
output c6196;
output c582;
output c6250;
output c5131;
output c6186;
output c6274;
output c3267;
output c9226;
output c316;
output c4201;
output c7137;
output c4250;
output c00;
output c8181;
output c647;
output c3129;
output c5136;
output c5290;
output c6159;
output c9170;
output c6231;
output c1277;
output c3121;
output c7283;
output c350;
output c0210;
output c263;
output c1228;
output c4165;
output c1168;
output c8198;
output c4184;
output c132;
output c2275;
output c9126;
output c6221;
output c7269;
output c1196;
output c860;
output c9185;
output c9116;
output c3286;
output c8211;
output c5291;
output c2288;
output c3100;
output c1162;
output c698;
output c5248;
output c0252;
output c0153;
output c4185;
output c692;
output c7162;
output c7295;
output c8287;
output c3197;
output c936;
output c6110;
output c847;
output c9299;
output c7140;
output c271;
output c1201;
output c5234;
output c125;
output c3166;
output c310;
output c027;
output c3292;
output c3220;
output c5229;
output c8133;
output c013;
output c338;
output c21;
output c355;
output c794;
output c5110;
output c4230;
output c564;
output c2100;
output c751;
output c8275;
output c7142;
output c862;
output c0255;
output c8146;
output c2265;
output c4124;
output c063;
output c1120;
output c4267;
output c8177;
output c53;
output c97;
output c423;
output c5297;
output c330;
output c4125;
output c83;
output c3165;
output c37;
output c193;
output c58;
output c1182;
output c7272;
output c0246;
output c8134;
output c227;
output c4168;
output c7248;
output c7167;
output c8163;
output c4290;
output c628;
output c967;
output c3266;
output c3143;
output c3276;
output c895;
output c332;
output c2153;
output c8206;
output c0162;
output c4104;
output c6209;
output c03;
output c2257;
output c6220;
output c9137;
output c2193;
output c0250;
output c7141;
output c0109;
output c4174;
output c4188;
output c0129;
output c913;
output c0191;
output c322;
output c1204;
output c1255;
output c632;
output c912;
output c925;
output c5210;
output c527;
output c635;
output c8244;
output c0168;
output c084;
output c3188;
output c0150;
output c452;
output c8123;
output c42;
output c340;
output c188;
output c566;
output c1207;
output c433;
output c5147;
output c7187;
output c8220;
output c942;
output c7265;
output c3298;
output c2262;
output c7220;
output c5288;
output c485;
output c531;
output c388;
output c9244;
output c176;
output c6290;
output c6222;
output c0118;
output c759;
output c587;
output c5217;
output c7165;
output c839;
output c230;
output c011;
output c149;
output c7150;
output c05;
output c160;
output c1297;
output c730;
output c4297;
output c5289;
output c8138;
output c174;
output c5148;
output c9228;
output c3160;
output c1259;
output c4294;
output c148;
output c8274;
output c250;
output c575;
output c436;
output c1209;
output c2158;
output c3186;
output c4141;
output c6116;
output c7292;
output c4166;
output c8103;
output c7262;
output c0116;
output c982;
output c2117;
output c3265;
output c2196;
output c968;
output c9261;
output c0259;
output c441;
output c096;
output c2105;
output c3150;
output c471;
output c9285;
output c3240;
output c727;
output c2256;
output c7232;
output c872;
output c039;
output c9293;
output c248;
output c976;
output c513;
output c898;
output c2287;
output c5144;
output c8115;
output c010;
output c9277;
output c5250;
output c5287;
output c3102;
output c2254;
output c552;
output c7256;
output c617;
output c7189;
output c2137;
output c9263;
output c914;
output c6118;
output c6100;
output c2103;
output c916;
output c4110;
output c7245;
output c161;
output c012;
output c4202;
output c1274;
output c1185;
output c1285;
output c3167;
output c7251;
output c8223;
output c1183;
output c6133;
output c50;
output c7100;
output c0281;
output c7281;
output c1298;
output c7273;
output c9233;
output c943;
output c370;
output c4274;
output c6291;
output c468;
output c5299;
output c699;
output c2227;
output c238;
output c6131;
output c298;
output c140;
output c5121;
output c8249;
output c5163;
output c8155;
output c9248;
output c2155;
output c3162;
output c2172;
output c2258;
output c1160;
output c5256;
output c654;
output c8109;
output c9181;
output c1173;
output c3133;
output c3164;
output c63;
output c576;
output c9127;
output c8188;
output c134;
output c0288;
output c6260;
output c6194;
output c7230;
output c9202;
output c312;
output c797;
output c0139;
output c5203;
output c047;
output c472;
output c2276;
output c7233;
output c9196;
output c0108;
output c8128;
output c9197;
output c2104;
output c1288;
output c3154;
output c2101;
output c586;
output c5157;
output c2251;
output c6198;
output c774;
output c5197;
output c2148;
output c6111;
output c1294;
output c945;
output c6267;
output c8213;
output c54;
output c4108;
output c117;
output c5191;
output c828;
output c823;
output c3223;
output c3170;
output c284;
output c5102;
output c8110;
output c2233;
output c9173;
output c2278;
output c1100;
output c3214;
output c2268;
output c9207;
output c991;
output c4149;
output c1194;
output c457;
output c5137;
output c2289;
output c7206;
output c8166;
output c5239;
output c3118;
output c568;
output c2224;
output c2236;
output c294;
output c8281;
output c9225;
output c14;
output c1287;
output c994;
output c29;
output c6179;
output c1212;
output c283;
output c5233;
output c5200;
output c893;
output c756;
output c0105;
output c3239;
output c051;
output c7101;
output c8141;
output c487;
output c6268;
output c3124;
output c764;
output c5263;
output c865;
output c5270;
output c630;
output c6284;
output c6207;
output c261;
output c5101;
output c3109;
output c3169;
output c4116;
output c3225;
output c82;
output c8229;
output c6264;
output c9189;
output c525;
output c5238;
output c7146;
output c60;
output c3226;
output c5282;
output c6171;
output c431;
output c2108;
output c650;
output c4140;
output c4200;
output c4169;
output c746;
output c684;
output c2294;
output c5259;
output c6177;
output c4276;
output c556;
output c7242;
output c826;
output c320;
output c4198;
output c9246;
output c0148;
output c8185;
output c098;
output c0128;
output c8250;
output c329;
output c592;
output c9241;
output c253;
output c884;
output c2249;
output c391;
output c5120;
output c141;
output c8180;
output c4203;
output c7229;
output c8168;
output c584;
output c9122;
output c3201;
output c085;
output c653;
output c0158;
output c952;
output c6258;
output c8233;
output c74;
output c384;
output c4280;
output c6277;
output c1218;
output c5213;
output c7103;
output c3217;
output c8142;
output c8105;
output c0100;
output c0230;
output c5107;
output c3174;
output c972;
output c6163;
output c7226;
output c2145;
output c868;
output c2139;
output c1296;
output c04;
output c659;
output c168;
output c9270;
output c5178;
output c285;
output c6108;
output c5222;
output c7202;
output c8218;
output c9155;
output c4132;
output c6234;
output c3293;
output c4193;
output c7240;
output c3261;
output c425;
output c4231;
output c5214;
output c723;
output c4213;
output c0253;
output c2150;
output c5180;
output c6129;
output c6136;
output c49;
output c490;
output c4219;
output c8120;
output c8273;
output c1206;
output c3184;
output c5186;
output c772;
output c164;
output c8258;
output c4268;
output c0194;
output c4255;
output c0257;
output c395;
output c06;
output c572;
output c1197;
output c2234;
output c5199;
output c5224;
output c636;
output c9113;
output c9193;
output c033;
output c6200;
output c4225;
output c7285;
output c7291;
output c4150;
output c658;
output c092;
output c662;
output c032;
output c178;
output c5177;
output c026;
output c0275;
output c045;
output c1272;
output c1105;
output c8158;
output c9276;
output c8129;
output c2138;
output c888;
output c0119;
output c5161;
output c5117;
output c323;
output c4208;
output c871;
output c6169;
output c8247;
output c7223;
output c2167;
output c5285;
output c5284;
output c7176;
output c2129;
output c286;
output c1282;
output c929;
output c6239;
output c6279;
output c7277;
output c1150;
output c6272;
output c7169;
output c0165;
output c5207;
output c47;
output c325;
output c1299;
output c491;
output c5179;
output c2128;
output c028;
output c612;
output c3269;
output c0289;
output c1290;
output c5283;
output c2205;
output c120;
output c9206;
output c4232;
output c7133;
output c8245;
output c163;
output c789;
output c0186;
output c0157;
output c5156;
output c4159;
output c1134;
output c1217;
output c6228;
output c827;
output c428;
output c5241;
output c646;
output c448;
output c574;
output c766;
output c8260;
output c3299;
output c6190;
output c5293;
output c299;
output c6106;
output c1224;
output c3153;
output c6261;
output c26;
output c6142;
output c6223;
output c7241;
output c079;
output c1132;
output c6233;
output c2277;
output c8122;
output c9188;
output c158;
output c4251;
output c712;
output c260;
output c577;
output c1170;
output c3190;
output c6288;
output c3103;
output c474;
output c9296;
output c275;
output c1284;
output c6183;
output c897;
output c6193;
output c738;
output c84;
output c5260;
output c169;
output c5116;
output c2252;
output c495;
output c1202;
output c2110;
output c3203;
output c2245;
output c596;
output c2130;
output c9251;
output c824;
output c8157;
output c710;
output c742;
output c844;
output c4139;
output c7111;
output c7207;
output c687;
output c334;
output c3297;
output c724;
output c416;
output c5100;
output c6257;
output c2119;
output c5190;
output c3242;
output c9290;
output c0207;
output c1111;
output c4180;
output c6126;
output c1261;
output c8187;
output c3113;
output c8107;
output c877;
output c3137;
output c1278;
output c060;
output c5103;
output c616;
output c0147;
output c537;
output c7216;
output c2192;
output c0188;
output c8193;
output c8173;
output c999;
output c4199;
output c5109;
output c6154;
output c412;
output c7297;
output c7177;
output c435;
output c475;
output c8112;
output c0204;
output c8214;
output c426;
output c99;
output c6156;
output c029;
output c4189;
output c9112;
output c8199;
output c0265;
output c7213;
output c9146;
output c4277;
output c3205;
output c3272;
output c7120;
output c0219;
output c8204;
output c2132;
output c1112;
output c4260;
output c3206;
output c9102;
output c265;
output c257;
output c2217;
output c331;
output c3180;
output c0262;
output c5261;
output c2248;
output c9179;
output c2168;
output c9200;
output c1213;
output c0254;
output c7185;
output c6182;
output c3196;
output c2229;
output c8285;
output c622;
output c985;
output c7200;
output c8209;
output c7204;
output c9174;
output c955;
output c1248;
output c8203;
output c480;
output c2199;
output c9214;
output c5183;
output c3237;
output c663;
output c9108;
output c3168;
output c9195;
output c714;
output c2113;
output c7118;
output c9286;
output c2271;
output c0151;
output c2118;
output c718;
output c7212;
output c9130;
output c6218;
output c9223;
output c31;
output c96;
output c311;
output c277;
output c6167;
output c561;
output c760;
output c6253;
output c0175;
output c0190;
output c1247;
output c5236;
output c0264;
output c833;
output c1221;
output c9239;
output c682;
output c0113;
output c156;
output c966;
output c8200;
output c8164;
output c571;
output c5132;
output c0173;
output c251;
output c2159;
output c4217;
output c732;
output c691;
output c7109;
output c461;
output c7135;
output c2260;
output c1151;
output c056;
output c4292;
output c726;
output c9139;
output c6204;
output c3273;
output c8106;
output c11;
output c6103;
output c8125;
output c1246;
output c8254;
output c7227;
output c8201;
output c4296;
output c5204;
output c8286;
output c3104;
output c40;
output c6141;
output c133;
output c45;
output c2226;
output c717;
output c5298;
output c7246;
output c8127;
output c281;
output c2270;
output c0213;
output c8167;
output c086;
output c3264;
output c5272;
output c1291;
output c454;
output c9222;
output c2146;
output c6121;
output c5245;
output c3191;
output c1114;
output c7210;
output c4233;
output c8242;
output c588;
output c6249;
output c019;
output c0271;
output c7299;
output c79;
output c849;
output c1117;
output c198;
output c570;
output c2246;
output c778;
output c3232;
output c0126;
output c9141;
output c3248;
output c563;
output c542;
output c10;
output c0130;
output c2190;
output c928;
output c930;
output c8265;
output c362;
output c3145;
output c8246;
output c5211;
output c8222;
output c8226;
output c9288;
output c6146;
output c6210;
output c2107;
output c3192;
output c328;
output c9220;
output c7271;
output c2135;
output c597;
output c7219;
output c675;
output c8294;
output c1270;
output c4288;
output c4157;
output c5209;
output c838;
output c9172;
output c7160;
output c7172;
output c374;
output c963;
output c4257;
output c511;
output c768;
output c2231;
output c4252;
output c569;
output c01;
output c042;
output c885;
output c9187;
output c585;
output c496;
output c162;
output c7170;
output c183;
output c8279;
output c3189;
output c9257;
output c949;
output c829;
output c2255;
output c3122;
output c1141;
output c8269;
output c950;
output c5192;
output c0159;
output c0141;
output c6191;
output c9209;
output c1205;
output c462;
output c8190;
output c4101;
output c8284;
output c9227;
output c0278;
output c48;
output c6143;
output c443;
output c4299;
output c3244;
output c110;
output c9103;
output c082;
output c269;
output c6212;
output c9184;
output c2230;
output c266;
output c5275;
output c763;
output c0285;
output c4181;
output c7222;
output c3246;
output c5198;
output c560;
output c5124;
output c0163;
output c5174;
output c421;
output c9203;
output c1256;
output c438;
output c567;
output c744;
output c3158;
output c3176;
output c89;
output c7267;
output c8282;
output c352;
output c4191;
output c0233;
output c6203;
output c735;
output c488;
output c8117;
output c4172;
output c782;
output c215;
output c5138;
output c7217;
output c713;
output c0187;
output c7288;
output c5135;
output c236;
output c6251;
output c1254;
output c595;
output c9213;
output c0208;
output c1241;
output c2244;
output c94;
output c961;
output c0239;
output c739;
output c181;
output c44;
output c6236;
output c3234;
output c599;
output c3231;
output c3277;
output c9250;
output c798;
output c7296;
output c7139;
output c5104;
output c0223;
output c135;
output c3195;
output c025;
output c089;
output c1243;
output c644;
output c363;
output c229;
output c093;
output c5130;
output c8228;
output c3211;
output c5133;
output c640;
output c613;
output c9144;
output c3283;
output c750;
output c8235;
output c6181;
output c015;
output c359;
output c672;
output c8225;
output c696;
output c7136;
output c9275;
output c822;
output c6152;
output c4173;
output c7128;
output c2175;
output c9232;
output c4244;
output c758;
output c3135;
output c2218;
output c430;
output c535;
output c28;
output c3181;
output c67;
output c4197;
output c670;
output c995;
output c339;
output c5196;
output c9136;
output c1263;
output c6197;
output c5277;
output c2176;
output c3136;
output c038;
output c351;
output c4121;
output c5205;
output c4190;
output c562;
output c7179;
output c424;
output c1167;
output c2170;
output c2184;
output c5188;
output c389;
output c3175;
output c1240;
output c411;
output c7257;
output c8296;
output c4114;
output c241;
output c1190;
output c4111;
output c4269;
output c097;
output c536;
output c5106;
output c456;
output c1169;
output c4155;
output c57;
output c6138;
output c152;
output c6270;
output c922;
output c0269;
output c361;
output c6140;
output c78;
output c580;
output c0279;
output c0182;
output c0181;
output c3173;
output c3134;
output c590;
output c20;
output c1189;
output c3257;
output c4287;
output c414;
output c9262;
output c6115;
output c1238;
output c8165;
output c2144;
output c944;
output c5194;
output c1158;
output c6295;
output c741;
output c2124;
output c2208;
output c2284;
output c3280;
output c5252;
output c3107;
output c6281;
output c989;
output c2177;
output c0156;
output c9115;
output c386;
output c7199;
output c8179;
output c6240;
output c2290;
output c9230;
output c8232;
output c130;
output c6187;
output c6232;
output c2164;
output c9234;
output c840;
output c6122;
output c834;
output c987;
output c055;
output c234;
output c1122;
output c223;
output c0220;
output c123;
output c5153;
output c6283;
output c8108;
output c4272;
output c9242;
output c7196;
output c992;
output c965;
output c2188;
output c6282;
output c9111;
output c2225;
output c7276;
output c0206;
output c5185;
output c4167;
output c7112;
output c1139;
output c8215;
output c0125;
output c8152;
output c7231;
output c4212;
output c112;
output c1188;
output c9183;
output c195;
output c6229;
output c8266;
output c8151;
output c2126;
output c5273;
output c415;
output c8121;
output c996;
output c282;
output c86;
output c3171;
output c382;
output c6242;
output c16;
output c2127;
output c51;
output c65;
output c2173;
output c451;
output c2261;
output c9180;
output c9212;
output c85;
output c851;
output c4224;
output c6107;
output c8159;
output c9114;
output c853;
output c546;
output c385;
output c6192;
output c0294;
output c0235;
output c459;
output c8212;
output c4103;
output c3130;
output c8297;
output c8172;
output c3204;
output c9194;
output c0267;
output c1283;
output c1244;
output c1215;
output c777;
output c383;
output c167;
output c4265;
output c869;
output c2243;
output c8184;
output c287;
output c7274;
output c1129;
output c69;
output c017;
output c7117;
output c2202;
output c1149;
output c7115;
output c814;
output c5162;
output c779;
output c6217;
output c2143;
output c4264;
output c8216;
output c1234;
output c1211;
output c2291;
output c3151;
output c489;
output c858;
output c4214;
output c6280;
output c882;
output c7205;
output c8189;
output c0236;
output c379;
output c6150;
output c5122;
output c4135;
output c7158;
output c878;
output c068;
output c0185;
output c1152;
output c3222;
output c5158;
output c795;
output c9268;
output c197;
output c319;
output c988;
output c1250;
output c393;
output c2219;
output c1292;
output c8147;
output c9198;
output c1237;
output c2165;
output c053;
output c256;
output c3179;
output c5151;
output c9271;
output c796;
output c92;
output c129;
output c5149;
output c418;
output c676;
output c614;
output c7181;
output c9192;
output c4162;
output c4215;
output c8131;
output c7252;
output c3275;
output c0261;
output c8238;
output c5202;
output c890;
output c5139;
output c581;
output c434;
output c9273;
output c6246;
output c3198;
output c551;
output c3144;
output c02;
output c565;
output c073;
output c8171;
output c4275;
output c136;
output c61;
output c7183;
output c8217;
output c1157;
output c326;
output c3185;
output c757;
output c7107;
output c5262;
output c573;
output c3285;
output c7261;
output c4262;
output c7194;
output c466;
output c9163;
output c2115;
output c5114;
output c228;
output c523;
output c5235;
output c761;
output c787;
output c59;
output c5247;
output c9279;
output c5230;
output c021;
output c317;
output c354;
output c2274;
output c6226;
output c522;
output c7239;
output c3290;
output c4278;
output c341;
output c0242;
output c151;
output c728;
output c7153;
output c639;
output c3149;
output c037;
output c2267;
output c091;
output c9224;
output c6185;
output c0200;
output c1108;
output c7258;
output c8256;
output c274;
output c8252;
output c9210;
output c553;
output c648;
output c850;
output c7284;
output c0282;
output c842;
output c5123;
output c781;
output c998;
output c8101;
output c784;
output c9231;
output c3296;
output c2109;
output c245;
output c022;
output c8261;
output c273;
output c1101;
output c2186;
output c6104;
output c3262;
output c959;
output c2194;
output c2296;
output c3288;
output c128;
output c870;
output c8135;
output c921;
output c6117;
output c831;
output c8298;
output c8271;
output c6139;
output c694;
output c1289;
output c072;
output c3247;
output c8210;
output c8234;
output c410;
output c7178;
output c6176;
output c775;
output c059;
output c080;
output c118;
output c1165;
output c4227;
output c510;
output c9152;
output c641;
output c593;
output c984;
output c6211;
output c854;
output c1208;
output c1126;
output c6124;
output c8124;
output c8197;
output c975;
output c5242;
output c6160;
output c4158;
output c8240;
output c9153;
output c7193;
output c7215;
output c9259;
output c077;
output c2279;
output c3178;
output c4105;
output c9160;
output c429;
output c6175;
output c9284;
output c8230;
output c863;
output c235;
output c821;
output c951;
output c9291;
output c5227;
output c4176;
output c8241;
output c657;

assign c00 =  x184 &  x601 & ~x29 & ~x86 & ~x88 & ~x97 & ~x102 & ~x111 & ~x113 & ~x136 & ~x168 & ~x190 & ~x194 & ~x249 & ~x278 & ~x286 & ~x305 & ~x310 & ~x336 & ~x359 & ~x386 & ~x417 & ~x422 & ~x423 & ~x450 & ~x475 & ~x496 & ~x504 & ~x510 & ~x527 & ~x589 & ~x612 & ~x613 & ~x617 & ~x621 & ~x634 & ~x666 & ~x680 & ~x681 & ~x683 & ~x699 & ~x700 & ~x704 & ~x713 & ~x716 & ~x736 & ~x737 & ~x759 & ~x767 & ~x774 & ~x783;
assign c02 =  x537 & ~x18 & ~x53 & ~x94 & ~x98 & ~x129 & ~x154 & ~x251 & ~x277 & ~x409 & ~x432 & ~x447 & ~x460 & ~x514 & ~x558 & ~x615 & ~x643 & ~x665 & ~x678 & ~x723 & ~x726 & ~x754;
assign c04 =  x401 &  x512 &  x625 & ~x229 & ~x308 & ~x563 & ~x644 & ~x674 & ~x700 & ~x774;
assign c06 =  x369 &  x414 &  x425 &  x453 & ~x20 & ~x81 & ~x256 & ~x403 & ~x408 & ~x410 & ~x411 & ~x421 & ~x423 & ~x431 & ~x434 & ~x563 & ~x691 & ~x692 & ~x697 & ~x716 & ~x721;
assign c08 =  x187 &  x385 &  x399 & ~x3 & ~x6 & ~x7 & ~x10 & ~x16 & ~x17 & ~x23 & ~x33 & ~x38 & ~x44 & ~x69 & ~x82 & ~x86 & ~x89 & ~x90 & ~x93 & ~x106 & ~x112 & ~x119 & ~x121 & ~x147 & ~x148 & ~x164 & ~x172 & ~x174 & ~x175 & ~x202 & ~x204 & ~x227 & ~x256 & ~x258 & ~x278 & ~x308 & ~x312 & ~x338 & ~x363 & ~x366 & ~x378 & ~x417 & ~x430 & ~x448 & ~x449 & ~x459 & ~x474 & ~x499 & ~x557 & ~x607 & ~x639 & ~x640 & ~x648 & ~x661 & ~x662 & ~x667 & ~x668 & ~x670 & ~x686 & ~x705 & ~x708 & ~x713 & ~x714 & ~x721 & ~x726 & ~x754 & ~x758 & ~x769 & ~x772 & ~x783;
assign c010 =  x154 &  x262 & ~x17 & ~x46 & ~x53 & ~x55 & ~x61 & ~x62 & ~x78 & ~x84 & ~x93 & ~x114 & ~x116 & ~x136 & ~x139 & ~x200 & ~x220 & ~x222 & ~x223 & ~x281 & ~x305 & ~x334 & ~x349 & ~x364 & ~x366 & ~x396 & ~x405 & ~x476 & ~x502 & ~x506 & ~x507 & ~x557 & ~x590 & ~x614 & ~x620 & ~x621 & ~x692 & ~x722 & ~x729 & ~x763 & ~x765;
assign c012 =  x416 &  x444 &  x483 & ~x97 & ~x352 & ~x353 & ~x354 & ~x381 & ~x383 & ~x408 & ~x409 & ~x433 & ~x436 & ~x438 & ~x439 & ~x440 & ~x459 & ~x460 & ~x461 & ~x462 & ~x464 & ~x465 & ~x466 & ~x467 & ~x489 & ~x490 & ~x491 & ~x780;
assign c014 =  x239 &  x267 &  x386 &  x414 &  x442 & ~x7 & ~x81 & ~x96 & ~x103 & ~x150 & ~x166 & ~x336 & ~x364 & ~x408 & ~x410 & ~x434 & ~x437 & ~x449 & ~x462 & ~x465 & ~x640 & ~x662 & ~x693 & ~x746;
assign c016 =  x471 &  x499 & ~x0 & ~x10 & ~x22 & ~x24 & ~x33 & ~x36 & ~x38 & ~x44 & ~x66 & ~x69 & ~x70 & ~x71 & ~x87 & ~x91 & ~x99 & ~x106 & ~x109 & ~x112 & ~x117 & ~x140 & ~x143 & ~x144 & ~x193 & ~x198 & ~x225 & ~x228 & ~x254 & ~x279 & ~x281 & ~x307 & ~x311 & ~x334 & ~x346 & ~x347 & ~x362 & ~x375 & ~x376 & ~x380 & ~x381 & ~x390 & ~x394 & ~x403 & ~x404 & ~x408 & ~x409 & ~x410 & ~x418 & ~x432 & ~x434 & ~x438 & ~x439 & ~x463 & ~x464 & ~x476 & ~x491 & ~x492 & ~x494 & ~x558 & ~x560 & ~x561 & ~x586 & ~x588 & ~x612 & ~x618 & ~x619 & ~x642 & ~x643 & ~x647 & ~x665 & ~x675 & ~x677 & ~x695 & ~x698 & ~x699 & ~x709 & ~x711 & ~x712 & ~x715 & ~x722 & ~x731 & ~x738 & ~x740 & ~x750 & ~x757 & ~x760 & ~x762 & ~x773 & ~x775 & ~x783;
assign c018 =  x331 &  x482 &  x539 & ~x7 & ~x8 & ~x17 & ~x18 & ~x26 & ~x30 & ~x42 & ~x65 & ~x85 & ~x94 & ~x98 & ~x103 & ~x112 & ~x115 & ~x141 & ~x142 & ~x169 & ~x171 & ~x196 & ~x222 & ~x255 & ~x279 & ~x283 & ~x309 & ~x327 & ~x338 & ~x355 & ~x356 & ~x382 & ~x383 & ~x390 & ~x410 & ~x411 & ~x436 & ~x476 & ~x477 & ~x506 & ~x558 & ~x560 & ~x587 & ~x592 & ~x616 & ~x645 & ~x664 & ~x668 & ~x669 & ~x691 & ~x695 & ~x699 & ~x715 & ~x718 & ~x720 & ~x728 & ~x735 & ~x738 & ~x740 & ~x741 & ~x742 & ~x745 & ~x748 & ~x749 & ~x757 & ~x770 & ~x775 & ~x780;
assign c020 = ~x1 & ~x3 & ~x7 & ~x8 & ~x11 & ~x23 & ~x24 & ~x25 & ~x29 & ~x33 & ~x35 & ~x36 & ~x38 & ~x47 & ~x49 & ~x51 & ~x52 & ~x55 & ~x61 & ~x63 & ~x69 & ~x72 & ~x80 & ~x83 & ~x87 & ~x94 & ~x99 & ~x113 & ~x132 & ~x137 & ~x138 & ~x141 & ~x165 & ~x169 & ~x170 & ~x172 & ~x193 & ~x220 & ~x221 & ~x225 & ~x251 & ~x253 & ~x257 & ~x278 & ~x279 & ~x283 & ~x321 & ~x341 & ~x348 & ~x368 & ~x376 & ~x377 & ~x418 & ~x432 & ~x446 & ~x461 & ~x508 & ~x517 & ~x534 & ~x547 & ~x561 & ~x563 & ~x586 & ~x588 & ~x616 & ~x619 & ~x623 & ~x640 & ~x643 & ~x651 & ~x667 & ~x673 & ~x680 & ~x681 & ~x695 & ~x701 & ~x706 & ~x719 & ~x720 & ~x726 & ~x733 & ~x735 & ~x738 & ~x743 & ~x744 & ~x745 & ~x764 & ~x769 & ~x774 & ~x778 & ~x782;
assign c022 =  x669;
assign c024 =  x236 &  x289 &  x316 &  x317 &  x371 &  x399 &  x427 & ~x3 & ~x4 & ~x6 & ~x7 & ~x10 & ~x11 & ~x17 & ~x19 & ~x22 & ~x28 & ~x31 & ~x36 & ~x37 & ~x38 & ~x45 & ~x48 & ~x50 & ~x52 & ~x55 & ~x56 & ~x57 & ~x58 & ~x62 & ~x64 & ~x65 & ~x66 & ~x67 & ~x68 & ~x71 & ~x73 & ~x74 & ~x76 & ~x82 & ~x84 & ~x85 & ~x92 & ~x94 & ~x97 & ~x107 & ~x111 & ~x116 & ~x117 & ~x120 & ~x121 & ~x134 & ~x136 & ~x137 & ~x143 & ~x145 & ~x146 & ~x163 & ~x164 & ~x165 & ~x166 & ~x168 & ~x171 & ~x191 & ~x192 & ~x193 & ~x195 & ~x197 & ~x220 & ~x221 & ~x226 & ~x227 & ~x249 & ~x252 & ~x253 & ~x255 & ~x277 & ~x278 & ~x279 & ~x282 & ~x305 & ~x306 & ~x308 & ~x309 & ~x311 & ~x334 & ~x337 & ~x338 & ~x339 & ~x340 & ~x362 & ~x363 & ~x364 & ~x365 & ~x368 & ~x375 & ~x390 & ~x394 & ~x395 & ~x396 & ~x408 & ~x419 & ~x421 & ~x436 & ~x437 & ~x447 & ~x449 & ~x475 & ~x478 & ~x502 & ~x504 & ~x505 & ~x506 & ~x507 & ~x535 & ~x559 & ~x586 & ~x616 & ~x619 & ~x639 & ~x643 & ~x645 & ~x646 & ~x647 & ~x670 & ~x675 & ~x679 & ~x694 & ~x697 & ~x700 & ~x701 & ~x704 & ~x705 & ~x709 & ~x711 & ~x716 & ~x717 & ~x718 & ~x720 & ~x721 & ~x722 & ~x725 & ~x726 & ~x728 & ~x730 & ~x733 & ~x737 & ~x738 & ~x740 & ~x743 & ~x745 & ~x746 & ~x747 & ~x749 & ~x750 & ~x752 & ~x756 & ~x767 & ~x768 & ~x769 & ~x771 & ~x773 & ~x777 & ~x780 & ~x781 & ~x782;
assign c026 =  x329 & ~x32 & ~x48 & ~x59 & ~x89 & ~x123 & ~x139 & ~x141 & ~x149 & ~x150 & ~x171 & ~x204 & ~x451 & ~x488 & ~x507 & ~x562 & ~x607 & ~x644 & ~x663 & ~x698 & ~x736 & ~x747 & ~x760;
assign c028 =  x348 &  x354 &  x382 &  x431 &  x459 & ~x5 & ~x13 & ~x26 & ~x62 & ~x76 & ~x79 & ~x81 & ~x93 & ~x110 & ~x111 & ~x132 & ~x134 & ~x165 & ~x220 & ~x276 & ~x309 & ~x311 & ~x330 & ~x366 & ~x369 & ~x414 & ~x426 & ~x434 & ~x451 & ~x471 & ~x503 & ~x531 & ~x536 & ~x537 & ~x538 & ~x620 & ~x642 & ~x651 & ~x665 & ~x668 & ~x690 & ~x726 & ~x734 & ~x760 & ~x771 & ~x772 & ~x777;
assign c030 =  x290 &  x401 &  x429 &  x467 &  x485 &  x628 &  x630 & ~x12 & ~x15 & ~x29 & ~x71 & ~x81 & ~x85 & ~x120 & ~x142 & ~x163 & ~x170 & ~x171 & ~x173 & ~x175 & ~x196 & ~x199 & ~x249 & ~x277 & ~x278 & ~x281 & ~x313 & ~x472 & ~x479 & ~x481 & ~x554 & ~x583 & ~x610 & ~x612 & ~x636 & ~x645 & ~x662 & ~x664 & ~x665 & ~x689 & ~x714 & ~x723 & ~x725 & ~x744 & ~x760 & ~x766 & ~x767 & ~x768 & ~x776;
assign c032 =  x64 &  x108;
assign c034 =  x773;
assign c036 = ~x6 & ~x7 & ~x9 & ~x13 & ~x14 & ~x15 & ~x18 & ~x21 & ~x23 & ~x24 & ~x25 & ~x26 & ~x27 & ~x28 & ~x31 & ~x34 & ~x35 & ~x36 & ~x37 & ~x39 & ~x40 & ~x41 & ~x43 & ~x45 & ~x46 & ~x49 & ~x52 & ~x53 & ~x54 & ~x55 & ~x56 & ~x57 & ~x59 & ~x60 & ~x61 & ~x63 & ~x65 & ~x66 & ~x67 & ~x69 & ~x70 & ~x71 & ~x74 & ~x75 & ~x78 & ~x79 & ~x81 & ~x83 & ~x86 & ~x87 & ~x88 & ~x90 & ~x91 & ~x92 & ~x93 & ~x105 & ~x107 & ~x111 & ~x113 & ~x114 & ~x115 & ~x118 & ~x119 & ~x120 & ~x122 & ~x134 & ~x135 & ~x139 & ~x140 & ~x142 & ~x143 & ~x146 & ~x162 & ~x165 & ~x168 & ~x169 & ~x170 & ~x173 & ~x174 & ~x192 & ~x193 & ~x194 & ~x195 & ~x197 & ~x199 & ~x200 & ~x203 & ~x221 & ~x222 & ~x223 & ~x225 & ~x249 & ~x252 & ~x253 & ~x279 & ~x280 & ~x281 & ~x306 & ~x307 & ~x308 & ~x309 & ~x310 & ~x312 & ~x313 & ~x338 & ~x340 & ~x341 & ~x363 & ~x364 & ~x365 & ~x366 & ~x367 & ~x368 & ~x377 & ~x378 & ~x379 & ~x391 & ~x392 & ~x394 & ~x405 & ~x407 & ~x419 & ~x433 & ~x434 & ~x436 & ~x437 & ~x446 & ~x447 & ~x448 & ~x450 & ~x451 & ~x452 & ~x463 & ~x475 & ~x476 & ~x477 & ~x478 & ~x489 & ~x504 & ~x505 & ~x506 & ~x529 & ~x530 & ~x534 & ~x536 & ~x560 & ~x561 & ~x562 & ~x563 & ~x564 & ~x584 & ~x585 & ~x587 & ~x588 & ~x589 & ~x590 & ~x592 & ~x610 & ~x612 & ~x617 & ~x618 & ~x635 & ~x638 & ~x639 & ~x641 & ~x643 & ~x644 & ~x645 & ~x648 & ~x649 & ~x661 & ~x663 & ~x666 & ~x671 & ~x673 & ~x674 & ~x677 & ~x686 & ~x691 & ~x692 & ~x693 & ~x694 & ~x697 & ~x699 & ~x702 & ~x703 & ~x704 & ~x705 & ~x706 & ~x707 & ~x708 & ~x709 & ~x710 & ~x711 & ~x712 & ~x713 & ~x714 & ~x716 & ~x717 & ~x718 & ~x723 & ~x725 & ~x726 & ~x728 & ~x729 & ~x730 & ~x731 & ~x734 & ~x735 & ~x738 & ~x742 & ~x744 & ~x745 & ~x746 & ~x749 & ~x750 & ~x751 & ~x754 & ~x755 & ~x756 & ~x757 & ~x759 & ~x761 & ~x763 & ~x765 & ~x768 & ~x771 & ~x772 & ~x773 & ~x776 & ~x778 & ~x779 & ~x780 & ~x783;
assign c038 =  x262 &  x290 &  x370 &  x398 &  x442 &  x470 & ~x408 & ~x432 & ~x434;
assign c040 =  x156 & ~x28 & ~x51 & ~x84 & ~x101 & ~x102 & ~x110 & ~x123 & ~x134 & ~x165 & ~x221 & ~x230 & ~x256 & ~x304 & ~x323 & ~x337 & ~x339 & ~x394 & ~x423 & ~x433 & ~x517 & ~x588 & ~x612 & ~x621 & ~x640 & ~x642 & ~x677 & ~x706 & ~x715 & ~x740 & ~x744 & ~x746 & ~x750 & ~x759 & ~x761 & ~x772 & ~x780;
assign c042 = ~x10 & ~x21 & ~x22 & ~x35 & ~x37 & ~x40 & ~x54 & ~x56 & ~x60 & ~x61 & ~x62 & ~x66 & ~x68 & ~x69 & ~x70 & ~x75 & ~x86 & ~x93 & ~x106 & ~x107 & ~x135 & ~x142 & ~x148 & ~x163 & ~x174 & ~x192 & ~x195 & ~x197 & ~x251 & ~x254 & ~x277 & ~x278 & ~x283 & ~x284 & ~x306 & ~x308 & ~x324 & ~x335 & ~x337 & ~x434 & ~x437 & ~x445 & ~x461 & ~x463 & ~x472 & ~x476 & ~x491 & ~x500 & ~x501 & ~x518 & ~x526 & ~x559 & ~x563 & ~x582 & ~x590 & ~x615 & ~x636 & ~x642 & ~x643 & ~x668 & ~x678 & ~x705 & ~x706 & ~x708 & ~x711 & ~x712 & ~x717 & ~x724 & ~x726 & ~x740 & ~x753 & ~x762 & ~x763 & ~x774 & ~x775 & ~x776 & ~x777;
assign c044 = ~x4 & ~x9 & ~x19 & ~x20 & ~x21 & ~x22 & ~x23 & ~x39 & ~x45 & ~x49 & ~x54 & ~x58 & ~x66 & ~x67 & ~x69 & ~x70 & ~x83 & ~x89 & ~x92 & ~x103 & ~x106 & ~x108 & ~x113 & ~x117 & ~x130 & ~x131 & ~x133 & ~x139 & ~x141 & ~x142 & ~x160 & ~x194 & ~x200 & ~x245 & ~x247 & ~x250 & ~x276 & ~x304 & ~x310 & ~x322 & ~x333 & ~x334 & ~x350 & ~x377 & ~x390 & ~x404 & ~x432 & ~x435 & ~x445 & ~x450 & ~x461 & ~x463 & ~x474 & ~x493 & ~x501 & ~x529 & ~x534 & ~x557 & ~x558 & ~x562 & ~x586 & ~x587 & ~x589 & ~x592 & ~x611 & ~x614 & ~x617 & ~x620 & ~x642 & ~x672 & ~x674 & ~x679 & ~x690 & ~x696 & ~x700 & ~x703 & ~x707 & ~x713 & ~x714 & ~x715 & ~x718 & ~x728 & ~x730 & ~x736 & ~x738 & ~x755 & ~x756 & ~x762 & ~x768 & ~x772 & ~x778 & ~x779 & ~x783;
assign c046 =  x426 &  x482 & ~x16 & ~x20 & ~x28 & ~x34 & ~x45 & ~x46 & ~x54 & ~x60 & ~x61 & ~x65 & ~x68 & ~x73 & ~x81 & ~x110 & ~x138 & ~x141 & ~x142 & ~x164 & ~x173 & ~x174 & ~x201 & ~x222 & ~x223 & ~x224 & ~x227 & ~x278 & ~x284 & ~x305 & ~x307 & ~x309 & ~x349 & ~x363 & ~x364 & ~x380 & ~x391 & ~x404 & ~x407 & ~x422 & ~x433 & ~x449 & ~x479 & ~x502 & ~x504 & ~x507 & ~x530 & ~x534 & ~x557 & ~x559 & ~x578 & ~x579 & ~x589 & ~x631 & ~x633 & ~x643 & ~x666 & ~x676 & ~x713 & ~x721 & ~x743 & ~x745 & ~x746 & ~x756 & ~x765 & ~x767 & ~x776;
assign c048 =  x245 &  x441 & ~x75 & ~x81 & ~x88 & ~x109 & ~x115 & ~x147 & ~x166 & ~x172 & ~x175 & ~x231 & ~x339 & ~x354 & ~x394 & ~x417 & ~x501 & ~x532 & ~x583 & ~x585 & ~x610 & ~x634 & ~x641 & ~x688 & ~x691 & ~x700 & ~x739 & ~x752 & ~x754 & ~x769 & ~x778;
assign c050 =  x400 & ~x7 & ~x12 & ~x17 & ~x18 & ~x31 & ~x36 & ~x54 & ~x61 & ~x62 & ~x63 & ~x69 & ~x70 & ~x77 & ~x79 & ~x82 & ~x88 & ~x93 & ~x98 & ~x107 & ~x108 & ~x119 & ~x145 & ~x146 & ~x169 & ~x171 & ~x173 & ~x177 & ~x198 & ~x205 & ~x224 & ~x251 & ~x255 & ~x258 & ~x277 & ~x283 & ~x286 & ~x314 & ~x335 & ~x339 & ~x362 & ~x364 & ~x366 & ~x367 & ~x389 & ~x391 & ~x395 & ~x409 & ~x431 & ~x445 & ~x447 & ~x449 & ~x450 & ~x459 & ~x504 & ~x529 & ~x531 & ~x532 & ~x534 & ~x557 & ~x580 & ~x581 & ~x585 & ~x588 & ~x610 & ~x618 & ~x634 & ~x640 & ~x641 & ~x642 & ~x647 & ~x665 & ~x668 & ~x671 & ~x688 & ~x693 & ~x696 & ~x702 & ~x703 & ~x708 & ~x709 & ~x710 & ~x713 & ~x714 & ~x720 & ~x722 & ~x723 & ~x726 & ~x730 & ~x731 & ~x733 & ~x738 & ~x742 & ~x744 & ~x746 & ~x748 & ~x749 & ~x766 & ~x767 & ~x769 & ~x770 & ~x782;
assign c052 =  x76 &  x444 &  x620;
assign c054 =  x210 & ~x0 & ~x1 & ~x9 & ~x10 & ~x14 & ~x24 & ~x30 & ~x38 & ~x39 & ~x41 & ~x45 & ~x48 & ~x51 & ~x53 & ~x66 & ~x67 & ~x70 & ~x71 & ~x73 & ~x76 & ~x79 & ~x101 & ~x103 & ~x109 & ~x111 & ~x113 & ~x115 & ~x117 & ~x118 & ~x120 & ~x122 & ~x127 & ~x131 & ~x132 & ~x134 & ~x138 & ~x146 & ~x147 & ~x163 & ~x164 & ~x175 & ~x176 & ~x192 & ~x193 & ~x194 & ~x198 & ~x202 & ~x203 & ~x221 & ~x228 & ~x249 & ~x256 & ~x277 & ~x278 & ~x282 & ~x311 & ~x313 & ~x333 & ~x339 & ~x362 & ~x366 & ~x367 & ~x393 & ~x394 & ~x409 & ~x421 & ~x437 & ~x446 & ~x448 & ~x465 & ~x473 & ~x476 & ~x491 & ~x493 & ~x529 & ~x532 & ~x534 & ~x545 & ~x556 & ~x559 & ~x561 & ~x583 & ~x589 & ~x615 & ~x616 & ~x664 & ~x666 & ~x668 & ~x670 & ~x671 & ~x674 & ~x675 & ~x692 & ~x696 & ~x697 & ~x702 & ~x704 & ~x712 & ~x713 & ~x716 & ~x720 & ~x721 & ~x730 & ~x744 & ~x750 & ~x752 & ~x758 & ~x762 & ~x767;
assign c056 =  x217 &  x374 &  x428 &  x596 & ~x29 & ~x66 & ~x67 & ~x75 & ~x108 & ~x672;
assign c058 =  x629 & ~x3 & ~x5 & ~x9 & ~x13 & ~x16 & ~x17 & ~x20 & ~x21 & ~x23 & ~x26 & ~x27 & ~x28 & ~x31 & ~x36 & ~x38 & ~x39 & ~x42 & ~x43 & ~x48 & ~x51 & ~x59 & ~x66 & ~x67 & ~x70 & ~x87 & ~x89 & ~x92 & ~x102 & ~x105 & ~x117 & ~x119 & ~x130 & ~x131 & ~x137 & ~x138 & ~x140 & ~x141 & ~x142 & ~x143 & ~x145 & ~x159 & ~x161 & ~x164 & ~x166 & ~x167 & ~x168 & ~x170 & ~x171 & ~x188 & ~x190 & ~x194 & ~x196 & ~x197 & ~x198 & ~x220 & ~x221 & ~x224 & ~x249 & ~x250 & ~x252 & ~x277 & ~x280 & ~x307 & ~x308 & ~x310 & ~x320 & ~x339 & ~x348 & ~x361 & ~x362 & ~x363 & ~x365 & ~x366 & ~x367 & ~x376 & ~x377 & ~x404 & ~x406 & ~x416 & ~x420 & ~x433 & ~x434 & ~x435 & ~x445 & ~x447 & ~x461 & ~x462 & ~x464 & ~x473 & ~x474 & ~x488 & ~x490 & ~x491 & ~x502 & ~x506 & ~x518 & ~x519 & ~x520 & ~x530 & ~x532 & ~x583 & ~x587 & ~x589 & ~x592 & ~x613 & ~x614 & ~x621 & ~x644 & ~x645 & ~x647 & ~x667 & ~x677 & ~x691 & ~x694 & ~x695 & ~x697 & ~x700 & ~x703 & ~x704 & ~x705 & ~x706 & ~x707 & ~x708 & ~x710 & ~x718 & ~x719 & ~x723 & ~x727 & ~x731 & ~x736 & ~x739 & ~x740 & ~x741 & ~x743 & ~x744 & ~x746 & ~x747 & ~x750 & ~x753 & ~x755 & ~x761 & ~x768 & ~x782 & ~x783;
assign c060 =  x213 & ~x0 & ~x4 & ~x16 & ~x21 & ~x23 & ~x53 & ~x59 & ~x60 & ~x63 & ~x72 & ~x80 & ~x86 & ~x88 & ~x92 & ~x93 & ~x97 & ~x99 & ~x111 & ~x122 & ~x123 & ~x140 & ~x142 & ~x143 & ~x148 & ~x149 & ~x150 & ~x165 & ~x168 & ~x169 & ~x190 & ~x199 & ~x228 & ~x231 & ~x250 & ~x251 & ~x255 & ~x259 & ~x261 & ~x274 & ~x277 & ~x278 & ~x280 & ~x307 & ~x311 & ~x333 & ~x343 & ~x358 & ~x369 & ~x389 & ~x391 & ~x474 & ~x477 & ~x502 & ~x523 & ~x534 & ~x535 & ~x551 & ~x552 & ~x559 & ~x587 & ~x588 & ~x613 & ~x614 & ~x616 & ~x619 & ~x650 & ~x664 & ~x669 & ~x675 & ~x679 & ~x680 & ~x687 & ~x703 & ~x704 & ~x709 & ~x710 & ~x711 & ~x719 & ~x725 & ~x748 & ~x751 & ~x753 & ~x759 & ~x778 & ~x782;
assign c062 =  x317 &  x429 &  x513 &  x570 &  x628 & ~x6 & ~x9 & ~x10 & ~x48 & ~x76 & ~x86 & ~x87 & ~x142 & ~x162 & ~x189 & ~x230 & ~x304 & ~x305 & ~x309 & ~x391 & ~x393 & ~x425 & ~x448 & ~x489 & ~x508 & ~x538 & ~x564 & ~x587 & ~x618 & ~x652 & ~x669 & ~x697 & ~x710 & ~x719 & ~x722 & ~x757 & ~x766 & ~x771;
assign c064 =  x154 &  x180 &  x234 &  x316 &  x344 &  x483 &  x598 &  x628 &  x630 &  x631 & ~x10 & ~x11 & ~x15 & ~x29 & ~x30 & ~x33 & ~x66 & ~x70 & ~x74 & ~x76 & ~x78 & ~x82 & ~x85 & ~x93 & ~x98 & ~x99 & ~x100 & ~x116 & ~x117 & ~x133 & ~x136 & ~x169 & ~x170 & ~x192 & ~x198 & ~x202 & ~x228 & ~x252 & ~x255 & ~x256 & ~x257 & ~x277 & ~x284 & ~x285 & ~x307 & ~x313 & ~x335 & ~x362 & ~x367 & ~x394 & ~x421 & ~x451 & ~x475 & ~x502 & ~x504 & ~x505 & ~x531 & ~x561 & ~x615 & ~x617 & ~x618 & ~x619 & ~x646 & ~x677 & ~x694 & ~x695 & ~x707 & ~x715 & ~x722 & ~x727 & ~x729 & ~x732 & ~x734 & ~x767 & ~x768 & ~x770 & ~x772;
assign c066 =  x265 &  x326 &  x515 &  x543 &  x544 &  x551 & ~x46 & ~x58 & ~x98 & ~x132 & ~x146 & ~x424 & ~x446 & ~x452 & ~x636 & ~x664 & ~x701 & ~x767 & ~x783;
assign c068 = ~x11 & ~x14 & ~x23 & ~x42 & ~x68 & ~x71 & ~x101 & ~x106 & ~x109 & ~x116 & ~x121 & ~x129 & ~x191 & ~x194 & ~x196 & ~x230 & ~x256 & ~x276 & ~x322 & ~x343 & ~x378 & ~x387 & ~x419 & ~x420 & ~x504 & ~x517 & ~x518 & ~x533 & ~x559 & ~x590 & ~x613 & ~x618 & ~x648 & ~x651 & ~x680 & ~x694 & ~x707 & ~x715 & ~x721 & ~x727 & ~x728 & ~x747 & ~x756 & ~x757 & ~x770;
assign c070 =  x647;
assign c072 = ~x9 & ~x21 & ~x34 & ~x38 & ~x39 & ~x49 & ~x54 & ~x63 & ~x81 & ~x90 & ~x97 & ~x103 & ~x115 & ~x116 & ~x118 & ~x134 & ~x137 & ~x141 & ~x144 & ~x162 & ~x166 & ~x170 & ~x172 & ~x197 & ~x246 & ~x253 & ~x255 & ~x265 & ~x279 & ~x284 & ~x324 & ~x337 & ~x352 & ~x379 & ~x388 & ~x390 & ~x407 & ~x408 & ~x418 & ~x420 & ~x434 & ~x463 & ~x474 & ~x489 & ~x501 & ~x502 & ~x503 & ~x507 & ~x530 & ~x560 & ~x591 & ~x615 & ~x616 & ~x620 & ~x643 & ~x668 & ~x670 & ~x671 & ~x695 & ~x698 & ~x699 & ~x700 & ~x702 & ~x714 & ~x720 & ~x723 & ~x726 & ~x729 & ~x739 & ~x744 & ~x756 & ~x757 & ~x760 & ~x767 & ~x778 & ~x781 & ~x783;
assign c074 =  x188 &  x246 &  x330 &  x413 & ~x22 & ~x27 & ~x28 & ~x47 & ~x117 & ~x120 & ~x505 & ~x634 & ~x709 & ~x715 & ~x754;
assign c076 =  x215 &  x485 & ~x76 & ~x84 & ~x106 & ~x117 & ~x136 & ~x146 & ~x192 & ~x227 & ~x419 & ~x504 & ~x560 & ~x583 & ~x586 & ~x709 & ~x714 & ~x721 & ~x722 & ~x732 & ~x743 & ~x775;
assign c078 =  x355 &  x457 & ~x94 & ~x117 & ~x153 & ~x447 & ~x582 & ~x688 & ~x781;
assign c080 =  x571 & ~x5 & ~x6 & ~x7 & ~x8 & ~x10 & ~x12 & ~x13 & ~x14 & ~x19 & ~x21 & ~x23 & ~x25 & ~x27 & ~x29 & ~x30 & ~x34 & ~x37 & ~x38 & ~x43 & ~x51 & ~x54 & ~x58 & ~x59 & ~x62 & ~x66 & ~x72 & ~x77 & ~x79 & ~x82 & ~x92 & ~x93 & ~x98 & ~x102 & ~x109 & ~x115 & ~x117 & ~x119 & ~x121 & ~x124 & ~x131 & ~x133 & ~x137 & ~x142 & ~x144 & ~x150 & ~x159 & ~x161 & ~x166 & ~x167 & ~x169 & ~x170 & ~x172 & ~x187 & ~x189 & ~x190 & ~x192 & ~x195 & ~x200 & ~x203 & ~x217 & ~x221 & ~x224 & ~x228 & ~x244 & ~x247 & ~x256 & ~x276 & ~x277 & ~x282 & ~x285 & ~x305 & ~x307 & ~x309 & ~x311 & ~x332 & ~x334 & ~x335 & ~x336 & ~x339 & ~x360 & ~x361 & ~x363 & ~x364 & ~x365 & ~x369 & ~x390 & ~x392 & ~x406 & ~x419 & ~x420 & ~x434 & ~x451 & ~x506 & ~x531 & ~x558 & ~x582 & ~x583 & ~x584 & ~x585 & ~x586 & ~x588 & ~x593 & ~x609 & ~x610 & ~x616 & ~x617 & ~x618 & ~x620 & ~x637 & ~x641 & ~x642 & ~x643 & ~x651 & ~x653 & ~x664 & ~x669 & ~x672 & ~x679 & ~x680 & ~x682 & ~x692 & ~x694 & ~x697 & ~x698 & ~x704 & ~x709 & ~x712 & ~x713 & ~x715 & ~x718 & ~x723 & ~x724 & ~x730 & ~x731 & ~x733 & ~x734 & ~x736 & ~x743 & ~x745 & ~x747 & ~x758 & ~x760 & ~x761 & ~x766 & ~x767 & ~x768 & ~x773 & ~x774 & ~x776 & ~x779 & ~x781 & ~x783;
assign c082 =  x272 &  x328 &  x402 & ~x37 & ~x89 & ~x147 & ~x170 & ~x258 & ~x360 & ~x420 & ~x444 & ~x502 & ~x504 & ~x581 & ~x639 & ~x690 & ~x698 & ~x707 & ~x724 & ~x730 & ~x737 & ~x738;
assign c084 =  x359 &  x415 & ~x1 & ~x4 & ~x5 & ~x7 & ~x9 & ~x11 & ~x12 & ~x13 & ~x14 & ~x17 & ~x18 & ~x19 & ~x21 & ~x22 & ~x24 & ~x25 & ~x26 & ~x28 & ~x29 & ~x31 & ~x32 & ~x33 & ~x34 & ~x38 & ~x40 & ~x45 & ~x47 & ~x48 & ~x49 & ~x51 & ~x52 & ~x53 & ~x55 & ~x56 & ~x58 & ~x61 & ~x62 & ~x64 & ~x66 & ~x68 & ~x70 & ~x71 & ~x72 & ~x74 & ~x75 & ~x77 & ~x79 & ~x80 & ~x81 & ~x83 & ~x85 & ~x93 & ~x94 & ~x96 & ~x97 & ~x98 & ~x99 & ~x102 & ~x104 & ~x106 & ~x107 & ~x108 & ~x109 & ~x111 & ~x112 & ~x113 & ~x114 & ~x115 & ~x117 & ~x122 & ~x123 & ~x127 & ~x136 & ~x137 & ~x138 & ~x139 & ~x140 & ~x142 & ~x143 & ~x147 & ~x148 & ~x165 & ~x169 & ~x170 & ~x173 & ~x174 & ~x176 & ~x192 & ~x194 & ~x195 & ~x196 & ~x199 & ~x200 & ~x201 & ~x202 & ~x221 & ~x222 & ~x224 & ~x226 & ~x227 & ~x228 & ~x249 & ~x250 & ~x251 & ~x252 & ~x256 & ~x277 & ~x278 & ~x280 & ~x281 & ~x282 & ~x283 & ~x305 & ~x312 & ~x334 & ~x340 & ~x361 & ~x362 & ~x365 & ~x366 & ~x367 & ~x390 & ~x392 & ~x393 & ~x394 & ~x395 & ~x409 & ~x410 & ~x411 & ~x417 & ~x418 & ~x420 & ~x421 & ~x423 & ~x436 & ~x446 & ~x448 & ~x449 & ~x450 & ~x451 & ~x475 & ~x476 & ~x479 & ~x502 & ~x503 & ~x504 & ~x529 & ~x531 & ~x532 & ~x533 & ~x535 & ~x557 & ~x558 & ~x559 & ~x560 & ~x562 & ~x564 & ~x588 & ~x589 & ~x590 & ~x591 & ~x592 & ~x611 & ~x614 & ~x615 & ~x617 & ~x618 & ~x620 & ~x638 & ~x639 & ~x640 & ~x641 & ~x643 & ~x645 & ~x664 & ~x665 & ~x669 & ~x670 & ~x672 & ~x673 & ~x674 & ~x676 & ~x677 & ~x688 & ~x691 & ~x692 & ~x693 & ~x695 & ~x697 & ~x698 & ~x699 & ~x703 & ~x713 & ~x714 & ~x715 & ~x719 & ~x720 & ~x721 & ~x723 & ~x726 & ~x728 & ~x730 & ~x731 & ~x732 & ~x734 & ~x735 & ~x738 & ~x742 & ~x743 & ~x747 & ~x750 & ~x751 & ~x755 & ~x760 & ~x761 & ~x764 & ~x765 & ~x766 & ~x767 & ~x770 & ~x773 & ~x774 & ~x775 & ~x776 & ~x779 & ~x780;
assign c086 = ~x10 & ~x21 & ~x75 & ~x101 & ~x119 & ~x120 & ~x138 & ~x167 & ~x173 & ~x178 & ~x205 & ~x259 & ~x309 & ~x407 & ~x417 & ~x426 & ~x427 & ~x451 & ~x490 & ~x511 & ~x551 & ~x581 & ~x614 & ~x623 & ~x634 & ~x649 & ~x673 & ~x677 & ~x688 & ~x710 & ~x721 & ~x731 & ~x734 & ~x735 & ~x754 & ~x759 & ~x778;
assign c088 =  x238 &  x239 &  x241 &  x265 &  x266 &  x267 &  x268 &  x270 &  x345 &  x412 &  x428 &  x429 &  x440 &  x457 &  x468 & ~x0 & ~x6 & ~x22 & ~x27 & ~x28 & ~x30 & ~x40 & ~x45 & ~x55 & ~x57 & ~x76 & ~x77 & ~x83 & ~x85 & ~x94 & ~x101 & ~x106 & ~x107 & ~x142 & ~x165 & ~x171 & ~x195 & ~x198 & ~x199 & ~x225 & ~x229 & ~x249 & ~x252 & ~x256 & ~x278 & ~x279 & ~x284 & ~x336 & ~x365 & ~x396 & ~x418 & ~x420 & ~x449 & ~x477 & ~x504 & ~x558 & ~x561 & ~x585 & ~x614 & ~x644 & ~x647 & ~x666 & ~x667 & ~x670 & ~x672 & ~x695 & ~x704 & ~x722 & ~x723 & ~x742 & ~x749 & ~x761 & ~x762 & ~x763 & ~x772;
assign c090 =  x236 &  x262 &  x317 &  x455 & ~x17 & ~x22 & ~x30 & ~x39 & ~x44 & ~x48 & ~x69 & ~x82 & ~x89 & ~x91 & ~x96 & ~x98 & ~x99 & ~x105 & ~x111 & ~x119 & ~x123 & ~x124 & ~x135 & ~x136 & ~x137 & ~x140 & ~x146 & ~x164 & ~x171 & ~x191 & ~x195 & ~x227 & ~x282 & ~x306 & ~x309 & ~x334 & ~x335 & ~x338 & ~x375 & ~x395 & ~x404 & ~x405 & ~x406 & ~x408 & ~x434 & ~x436 & ~x463 & ~x464 & ~x507 & ~x530 & ~x535 & ~x558 & ~x589 & ~x647 & ~x673 & ~x694 & ~x716 & ~x718 & ~x720 & ~x736 & ~x738 & ~x743 & ~x751 & ~x755 & ~x756 & ~x757 & ~x764 & ~x765 & ~x766 & ~x776 & ~x781;
assign c092 =  x570 &  x630 &  x631 & ~x9 & ~x40 & ~x45 & ~x57 & ~x69 & ~x71 & ~x76 & ~x93 & ~x94 & ~x98 & ~x106 & ~x115 & ~x136 & ~x162 & ~x173 & ~x196 & ~x197 & ~x226 & ~x332 & ~x353 & ~x362 & ~x381 & ~x389 & ~x394 & ~x408 & ~x423 & ~x436 & ~x446 & ~x462 & ~x464 & ~x490 & ~x491 & ~x518 & ~x519 & ~x530 & ~x537 & ~x558 & ~x562 & ~x587 & ~x590 & ~x593 & ~x618 & ~x708 & ~x728 & ~x745 & ~x749 & ~x752 & ~x765 & ~x775;
assign c094 =  x287 &  x288 &  x315 &  x316 &  x370 &  x371 &  x398 &  x416 & ~x77 & ~x408 & ~x437 & ~x465;
assign c096 = ~x30 & ~x36 & ~x44 & ~x45 & ~x67 & ~x80 & ~x90 & ~x95 & ~x110 & ~x115 & ~x119 & ~x150 & ~x196 & ~x207 & ~x225 & ~x227 & ~x229 & ~x256 & ~x260 & ~x277 & ~x278 & ~x369 & ~x433 & ~x449 & ~x478 & ~x517 & ~x526 & ~x533 & ~x556 & ~x558 & ~x620 & ~x633 & ~x669 & ~x687 & ~x743;
assign c098 = ~x7 & ~x11 & ~x16 & ~x24 & ~x38 & ~x40 & ~x46 & ~x47 & ~x54 & ~x62 & ~x69 & ~x85 & ~x92 & ~x98 & ~x107 & ~x113 & ~x122 & ~x132 & ~x138 & ~x150 & ~x170 & ~x189 & ~x198 & ~x205 & ~x217 & ~x218 & ~x227 & ~x274 & ~x275 & ~x281 & ~x306 & ~x313 & ~x332 & ~x338 & ~x358 & ~x368 & ~x379 & ~x386 & ~x391 & ~x393 & ~x406 & ~x407 & ~x415 & ~x417 & ~x423 & ~x435 & ~x441 & ~x447 & ~x450 & ~x453 & ~x471 & ~x472 & ~x474 & ~x481 & ~x508 & ~x510 & ~x526 & ~x529 & ~x532 & ~x536 & ~x538 & ~x555 & ~x557 & ~x563 & ~x565 & ~x590 & ~x592 & ~x593 & ~x611 & ~x621 & ~x636 & ~x670 & ~x677 & ~x678 & ~x688 & ~x701 & ~x703 & ~x717 & ~x718 & ~x729 & ~x741 & ~x744 & ~x757 & ~x779;
assign c0100 =  x597 & ~x54 & ~x88 & ~x351 & ~x379 & ~x394 & ~x460 & ~x488 & ~x515 & ~x607 & ~x631 & ~x669;
assign c0102 =  x210 &  x269 &  x487 & ~x1 & ~x6 & ~x14 & ~x29 & ~x43 & ~x46 & ~x53 & ~x56 & ~x58 & ~x80 & ~x86 & ~x98 & ~x99 & ~x105 & ~x115 & ~x120 & ~x133 & ~x141 & ~x147 & ~x162 & ~x170 & ~x173 & ~x189 & ~x195 & ~x202 & ~x219 & ~x226 & ~x245 & ~x249 & ~x253 & ~x258 & ~x278 & ~x279 & ~x283 & ~x301 & ~x305 & ~x314 & ~x331 & ~x334 & ~x366 & ~x415 & ~x422 & ~x434 & ~x446 & ~x451 & ~x453 & ~x479 & ~x527 & ~x529 & ~x537 & ~x538 & ~x560 & ~x561 & ~x563 & ~x567 & ~x612 & ~x617 & ~x623 & ~x624 & ~x641 & ~x644 & ~x664 & ~x665 & ~x678 & ~x704 & ~x706 & ~x707 & ~x708 & ~x716 & ~x717 & ~x727 & ~x738 & ~x748 & ~x749 & ~x752 & ~x754 & ~x756 & ~x764 & ~x778;
assign c0104 =  x430 & ~x101 & ~x190 & ~x371 & ~x378 & ~x407 & ~x420 & ~x473 & ~x490 & ~x534 & ~x539 & ~x558 & ~x563 & ~x692 & ~x736 & ~x753;
assign c0106 =  x315 &  x397 &  x498 & ~x253 & ~x364 & ~x406 & ~x407 & ~x410 & ~x432 & ~x437 & ~x465 & ~x466 & ~x491;
assign c0108 =  x370 &  x398 & ~x0 & ~x1 & ~x2 & ~x3 & ~x4 & ~x5 & ~x7 & ~x8 & ~x9 & ~x10 & ~x11 & ~x12 & ~x13 & ~x14 & ~x15 & ~x16 & ~x18 & ~x19 & ~x21 & ~x22 & ~x23 & ~x24 & ~x27 & ~x29 & ~x30 & ~x32 & ~x35 & ~x36 & ~x37 & ~x38 & ~x39 & ~x40 & ~x41 & ~x42 & ~x43 & ~x44 & ~x45 & ~x46 & ~x47 & ~x48 & ~x49 & ~x50 & ~x51 & ~x52 & ~x53 & ~x55 & ~x56 & ~x58 & ~x59 & ~x60 & ~x61 & ~x62 & ~x63 & ~x64 & ~x65 & ~x66 & ~x68 & ~x69 & ~x70 & ~x71 & ~x72 & ~x74 & ~x75 & ~x76 & ~x77 & ~x78 & ~x79 & ~x80 & ~x82 & ~x84 & ~x86 & ~x88 & ~x89 & ~x90 & ~x91 & ~x92 & ~x93 & ~x94 & ~x95 & ~x96 & ~x97 & ~x98 & ~x100 & ~x101 & ~x102 & ~x103 & ~x104 & ~x105 & ~x106 & ~x109 & ~x110 & ~x112 & ~x113 & ~x114 & ~x115 & ~x116 & ~x117 & ~x119 & ~x120 & ~x121 & ~x131 & ~x134 & ~x135 & ~x136 & ~x137 & ~x138 & ~x139 & ~x140 & ~x144 & ~x146 & ~x147 & ~x148 & ~x164 & ~x165 & ~x166 & ~x167 & ~x168 & ~x171 & ~x172 & ~x173 & ~x174 & ~x192 & ~x193 & ~x194 & ~x195 & ~x196 & ~x197 & ~x198 & ~x199 & ~x200 & ~x201 & ~x202 & ~x220 & ~x221 & ~x222 & ~x223 & ~x225 & ~x226 & ~x227 & ~x228 & ~x229 & ~x250 & ~x251 & ~x253 & ~x254 & ~x256 & ~x276 & ~x277 & ~x278 & ~x279 & ~x281 & ~x282 & ~x283 & ~x284 & ~x305 & ~x307 & ~x309 & ~x310 & ~x311 & ~x312 & ~x333 & ~x336 & ~x337 & ~x338 & ~x339 & ~x340 & ~x361 & ~x364 & ~x365 & ~x366 & ~x367 & ~x368 & ~x375 & ~x391 & ~x392 & ~x394 & ~x395 & ~x396 & ~x402 & ~x406 & ~x407 & ~x408 & ~x419 & ~x421 & ~x423 & ~x432 & ~x436 & ~x446 & ~x448 & ~x450 & ~x451 & ~x474 & ~x475 & ~x476 & ~x477 & ~x479 & ~x502 & ~x503 & ~x504 & ~x507 & ~x532 & ~x534 & ~x535 & ~x558 & ~x561 & ~x562 & ~x563 & ~x585 & ~x587 & ~x588 & ~x589 & ~x591 & ~x611 & ~x612 & ~x613 & ~x614 & ~x615 & ~x616 & ~x619 & ~x620 & ~x621 & ~x639 & ~x640 & ~x641 & ~x642 & ~x643 & ~x644 & ~x645 & ~x646 & ~x647 & ~x648 & ~x649 & ~x665 & ~x667 & ~x668 & ~x669 & ~x670 & ~x671 & ~x672 & ~x674 & ~x675 & ~x676 & ~x677 & ~x678 & ~x679 & ~x680 & ~x681 & ~x690 & ~x691 & ~x692 & ~x693 & ~x695 & ~x696 & ~x697 & ~x698 & ~x699 & ~x701 & ~x704 & ~x705 & ~x706 & ~x707 & ~x709 & ~x710 & ~x711 & ~x712 & ~x713 & ~x714 & ~x716 & ~x717 & ~x718 & ~x719 & ~x720 & ~x721 & ~x722 & ~x723 & ~x724 & ~x725 & ~x726 & ~x727 & ~x730 & ~x731 & ~x732 & ~x733 & ~x734 & ~x735 & ~x737 & ~x738 & ~x739 & ~x741 & ~x743 & ~x744 & ~x745 & ~x746 & ~x747 & ~x748 & ~x749 & ~x750 & ~x751 & ~x752 & ~x755 & ~x756 & ~x757 & ~x758 & ~x760 & ~x761 & ~x764 & ~x765 & ~x766 & ~x768 & ~x769 & ~x770 & ~x772 & ~x773 & ~x774 & ~x775 & ~x777 & ~x778 & ~x780 & ~x782 & ~x783;
assign c0110 =  x386 & ~x1 & ~x9 & ~x16 & ~x18 & ~x19 & ~x34 & ~x45 & ~x47 & ~x49 & ~x50 & ~x58 & ~x73 & ~x75 & ~x79 & ~x99 & ~x104 & ~x106 & ~x107 & ~x119 & ~x141 & ~x145 & ~x161 & ~x165 & ~x168 & ~x192 & ~x256 & ~x282 & ~x283 & ~x320 & ~x333 & ~x335 & ~x339 & ~x348 & ~x349 & ~x354 & ~x363 & ~x376 & ~x381 & ~x389 & ~x403 & ~x405 & ~x410 & ~x431 & ~x432 & ~x435 & ~x438 & ~x448 & ~x451 & ~x464 & ~x465 & ~x474 & ~x491 & ~x494 & ~x504 & ~x505 & ~x533 & ~x612 & ~x614 & ~x644 & ~x702 & ~x703 & ~x710 & ~x718 & ~x721 & ~x736 & ~x740 & ~x751 & ~x763 & ~x771;
assign c0112 =  x213 &  x270 & ~x0 & ~x4 & ~x5 & ~x19 & ~x31 & ~x35 & ~x71 & ~x94 & ~x100 & ~x114 & ~x123 & ~x136 & ~x154 & ~x163 & ~x172 & ~x175 & ~x208 & ~x248 & ~x255 & ~x259 & ~x306 & ~x339 & ~x364 & ~x396 & ~x423 & ~x446 & ~x447 & ~x461 & ~x501 & ~x507 & ~x531 & ~x560 & ~x585 & ~x636 & ~x637 & ~x661 & ~x671 & ~x687 & ~x694 & ~x703 & ~x717 & ~x736 & ~x737 & ~x753 & ~x759;
assign c0114 =  x264 &  x319 &  x344 &  x357 &  x373 &  x428 & ~x490;
assign c0116 =  x331 &  x359 & ~x0 & ~x5 & ~x11 & ~x12 & ~x19 & ~x26 & ~x34 & ~x39 & ~x41 & ~x44 & ~x47 & ~x70 & ~x72 & ~x74 & ~x75 & ~x81 & ~x84 & ~x85 & ~x90 & ~x104 & ~x107 & ~x114 & ~x118 & ~x123 & ~x126 & ~x134 & ~x136 & ~x166 & ~x169 & ~x170 & ~x172 & ~x196 & ~x197 & ~x198 & ~x204 & ~x256 & ~x326 & ~x327 & ~x334 & ~x336 & ~x354 & ~x355 & ~x361 & ~x365 & ~x393 & ~x394 & ~x395 & ~x418 & ~x450 & ~x476 & ~x504 & ~x590 & ~x616 & ~x638 & ~x666 & ~x667 & ~x676 & ~x677 & ~x688 & ~x695 & ~x697 & ~x698 & ~x705 & ~x708 & ~x709 & ~x712 & ~x718 & ~x720 & ~x721 & ~x725 & ~x727 & ~x728 & ~x731 & ~x732 & ~x736 & ~x738 & ~x745 & ~x746 & ~x750 & ~x752 & ~x756 & ~x762;
assign c0118 =  x315 &  x342 &  x343 &  x372 &  x399 &  x415 &  x471 &  x527;
assign c0120 =  x212 & ~x2 & ~x3 & ~x6 & ~x7 & ~x8 & ~x12 & ~x13 & ~x15 & ~x16 & ~x18 & ~x21 & ~x22 & ~x29 & ~x30 & ~x32 & ~x35 & ~x36 & ~x38 & ~x40 & ~x48 & ~x50 & ~x51 & ~x57 & ~x59 & ~x64 & ~x65 & ~x68 & ~x70 & ~x72 & ~x73 & ~x74 & ~x75 & ~x77 & ~x78 & ~x79 & ~x84 & ~x88 & ~x92 & ~x99 & ~x100 & ~x101 & ~x102 & ~x104 & ~x108 & ~x109 & ~x112 & ~x113 & ~x115 & ~x118 & ~x119 & ~x121 & ~x127 & ~x128 & ~x130 & ~x132 & ~x142 & ~x164 & ~x165 & ~x166 & ~x168 & ~x171 & ~x192 & ~x193 & ~x195 & ~x197 & ~x199 & ~x201 & ~x222 & ~x226 & ~x227 & ~x228 & ~x249 & ~x250 & ~x251 & ~x252 & ~x253 & ~x254 & ~x255 & ~x277 & ~x279 & ~x283 & ~x307 & ~x309 & ~x311 & ~x335 & ~x337 & ~x338 & ~x339 & ~x351 & ~x352 & ~x363 & ~x365 & ~x366 & ~x367 & ~x393 & ~x405 & ~x407 & ~x409 & ~x410 & ~x419 & ~x434 & ~x450 & ~x461 & ~x462 & ~x463 & ~x464 & ~x465 & ~x478 & ~x488 & ~x489 & ~x490 & ~x492 & ~x502 & ~x503 & ~x505 & ~x517 & ~x529 & ~x530 & ~x531 & ~x534 & ~x557 & ~x562 & ~x591 & ~x615 & ~x616 & ~x617 & ~x618 & ~x643 & ~x648 & ~x666 & ~x669 & ~x674 & ~x676 & ~x692 & ~x693 & ~x694 & ~x698 & ~x700 & ~x701 & ~x710 & ~x711 & ~x718 & ~x719 & ~x720 & ~x721 & ~x723 & ~x727 & ~x729 & ~x730 & ~x731 & ~x733 & ~x734 & ~x740 & ~x745 & ~x747 & ~x752 & ~x754 & ~x755 & ~x756 & ~x762 & ~x766 & ~x770 & ~x772 & ~x774 & ~x778 & ~x780 & ~x783;
assign c0122 =  x25;
assign c0124 =  x766;
assign c0126 =  x212 &  x291 &  x412 &  x467 & ~x1 & ~x40 & ~x45 & ~x83 & ~x88 & ~x103 & ~x149 & ~x259 & ~x281 & ~x315 & ~x337 & ~x352 & ~x365 & ~x473 & ~x474 & ~x555 & ~x608 & ~x749 & ~x768;
assign c0128 =  x186 &  x215 &  x273 &  x357 &  x413 &  x441 &  x468 &  x496 &  x523 &  x626 & ~x4 & ~x18 & ~x19 & ~x111 & ~x136 & ~x141 & ~x145 & ~x167 & ~x168 & ~x170 & ~x227 & ~x276 & ~x310 & ~x390 & ~x391 & ~x451 & ~x506 & ~x530 & ~x531 & ~x608 & ~x609 & ~x636 & ~x646 & ~x649 & ~x669 & ~x709 & ~x733 & ~x734 & ~x765 & ~x782;
assign c0130 =  x571 & ~x0 & ~x3 & ~x6 & ~x12 & ~x14 & ~x16 & ~x18 & ~x26 & ~x27 & ~x29 & ~x42 & ~x45 & ~x46 & ~x51 & ~x54 & ~x55 & ~x56 & ~x60 & ~x75 & ~x78 & ~x89 & ~x91 & ~x95 & ~x99 & ~x101 & ~x103 & ~x119 & ~x135 & ~x145 & ~x146 & ~x147 & ~x149 & ~x161 & ~x165 & ~x168 & ~x170 & ~x171 & ~x173 & ~x190 & ~x193 & ~x194 & ~x195 & ~x202 & ~x231 & ~x254 & ~x259 & ~x274 & ~x283 & ~x303 & ~x309 & ~x313 & ~x336 & ~x340 & ~x350 & ~x389 & ~x416 & ~x423 & ~x473 & ~x500 & ~x501 & ~x529 & ~x530 & ~x554 & ~x566 & ~x582 & ~x588 & ~x591 & ~x615 & ~x622 & ~x640 & ~x647 & ~x650 & ~x664 & ~x670 & ~x682 & ~x688 & ~x706 & ~x707 & ~x714 & ~x720 & ~x731 & ~x736 & ~x749 & ~x753 & ~x755 & ~x757 & ~x758 & ~x765 & ~x775 & ~x777 & ~x778 & ~x780 & ~x783;
assign c0132 = ~x54 & ~x66 & ~x100 & ~x110 & ~x169 & ~x202 & ~x203 & ~x257 & ~x287 & ~x314 & ~x334 & ~x361 & ~x365 & ~x390 & ~x391 & ~x408 & ~x426 & ~x435 & ~x452 & ~x482 & ~x491 & ~x526 & ~x527 & ~x538 & ~x564 & ~x567 & ~x590 & ~x592 & ~x593 & ~x621 & ~x665 & ~x691 & ~x693 & ~x706 & ~x713 & ~x731 & ~x737 & ~x749 & ~x751 & ~x773;
assign c0134 =  x186 &  x293 &  x347 &  x540 & ~x0 & ~x3 & ~x6 & ~x75 & ~x84 & ~x90 & ~x105 & ~x109 & ~x121 & ~x151 & ~x194 & ~x197 & ~x204 & ~x227 & ~x258 & ~x306 & ~x309 & ~x339 & ~x390 & ~x395 & ~x445 & ~x498 & ~x523 & ~x527 & ~x528 & ~x531 & ~x555 & ~x563 & ~x579 & ~x591 & ~x604 & ~x605 & ~x606 & ~x610 & ~x632 & ~x644 & ~x646 & ~x668 & ~x686 & ~x707 & ~x711 & ~x720 & ~x721 & ~x738 & ~x760 & ~x776 & ~x779;
assign c0136 =  x429 &  x630 & ~x11 & ~x29 & ~x73 & ~x86 & ~x108 & ~x109 & ~x134 & ~x163 & ~x191 & ~x196 & ~x197 & ~x199 & ~x251 & ~x275 & ~x278 & ~x366 & ~x376 & ~x379 & ~x394 & ~x433 & ~x450 & ~x463 & ~x474 & ~x479 & ~x518 & ~x530 & ~x589 & ~x641 & ~x643 & ~x695 & ~x712 & ~x714 & ~x720 & ~x739 & ~x748 & ~x778;
assign c0138 =  x214 & ~x1 & ~x7 & ~x11 & ~x12 & ~x14 & ~x21 & ~x22 & ~x27 & ~x31 & ~x36 & ~x41 & ~x43 & ~x45 & ~x46 & ~x48 & ~x50 & ~x54 & ~x56 & ~x57 & ~x58 & ~x68 & ~x74 & ~x75 & ~x77 & ~x80 & ~x82 & ~x83 & ~x87 & ~x89 & ~x101 & ~x103 & ~x104 & ~x119 & ~x120 & ~x121 & ~x132 & ~x133 & ~x134 & ~x141 & ~x144 & ~x145 & ~x147 & ~x162 & ~x163 & ~x166 & ~x170 & ~x174 & ~x191 & ~x196 & ~x197 & ~x221 & ~x224 & ~x250 & ~x252 & ~x253 & ~x255 & ~x257 & ~x279 & ~x281 & ~x282 & ~x308 & ~x311 & ~x312 & ~x333 & ~x335 & ~x336 & ~x354 & ~x355 & ~x362 & ~x364 & ~x365 & ~x382 & ~x383 & ~x390 & ~x391 & ~x394 & ~x410 & ~x417 & ~x418 & ~x420 & ~x421 & ~x438 & ~x446 & ~x447 & ~x464 & ~x465 & ~x474 & ~x487 & ~x491 & ~x492 & ~x501 & ~x506 & ~x530 & ~x557 & ~x559 & ~x560 & ~x561 & ~x586 & ~x587 & ~x589 & ~x591 & ~x614 & ~x615 & ~x617 & ~x619 & ~x640 & ~x641 & ~x642 & ~x645 & ~x646 & ~x647 & ~x668 & ~x669 & ~x673 & ~x675 & ~x696 & ~x697 & ~x701 & ~x703 & ~x704 & ~x716 & ~x728 & ~x730 & ~x732 & ~x738 & ~x740 & ~x741 & ~x743 & ~x747 & ~x755 & ~x757 & ~x760 & ~x761 & ~x764 & ~x765 & ~x766 & ~x768 & ~x772 & ~x773 & ~x774 & ~x775 & ~x776 & ~x779 & ~x782;
assign c0140 =  x245 &  x246 &  x357 &  x510 & ~x150 & ~x175 & ~x203;
assign c0142 =  x430 & ~x17 & ~x41 & ~x57 & ~x65 & ~x391 & ~x405 & ~x406 & ~x447 & ~x461 & ~x489 & ~x523 & ~x557 & ~x616 & ~x618;
assign c0144 = ~x3 & ~x5 & ~x6 & ~x12 & ~x26 & ~x27 & ~x29 & ~x33 & ~x36 & ~x38 & ~x39 & ~x41 & ~x46 & ~x48 & ~x57 & ~x60 & ~x65 & ~x69 & ~x76 & ~x84 & ~x87 & ~x89 & ~x114 & ~x117 & ~x129 & ~x137 & ~x140 & ~x144 & ~x166 & ~x171 & ~x200 & ~x221 & ~x225 & ~x226 & ~x247 & ~x253 & ~x276 & ~x284 & ~x303 & ~x308 & ~x310 & ~x319 & ~x320 & ~x337 & ~x347 & ~x349 & ~x350 & ~x361 & ~x365 & ~x366 & ~x367 & ~x377 & ~x391 & ~x419 & ~x420 & ~x432 & ~x466 & ~x477 & ~x491 & ~x492 & ~x493 & ~x506 & ~x508 & ~x519 & ~x532 & ~x533 & ~x562 & ~x563 & ~x593 & ~x594 & ~x619 & ~x640 & ~x641 & ~x643 & ~x652 & ~x667 & ~x672 & ~x692 & ~x699 & ~x700 & ~x710 & ~x711 & ~x712 & ~x717 & ~x721 & ~x726 & ~x729 & ~x737 & ~x738 & ~x741 & ~x744 & ~x745 & ~x749 & ~x750 & ~x752 & ~x757 & ~x758 & ~x773 & ~x775 & ~x779 & ~x780 & ~x782;
assign c0146 =  x327 &  x348 &  x411 &  x430 & ~x63 & ~x146 & ~x196 & ~x247 & ~x250 & ~x288 & ~x390 & ~x449 & ~x501;
assign c0148 =  x327 &  x383 &  x429 & ~x24 & ~x29 & ~x49 & ~x58 & ~x59 & ~x72 & ~x96 & ~x105 & ~x122 & ~x144 & ~x199 & ~x230 & ~x231 & ~x248 & ~x259 & ~x314 & ~x336 & ~x367 & ~x391 & ~x393 & ~x414 & ~x425 & ~x470 & ~x554 & ~x561 & ~x589 & ~x609 & ~x634 & ~x636 & ~x642 & ~x644 & ~x661 & ~x663 & ~x669 & ~x670 & ~x676 & ~x696 & ~x697 & ~x708 & ~x711 & ~x724 & ~x739 & ~x741 & ~x749 & ~x769;
assign c0150 =  x184 &  x238 &  x628 & ~x1 & ~x9 & ~x10 & ~x12 & ~x24 & ~x31 & ~x40 & ~x54 & ~x55 & ~x64 & ~x81 & ~x119 & ~x121 & ~x131 & ~x163 & ~x164 & ~x166 & ~x168 & ~x169 & ~x174 & ~x222 & ~x224 & ~x249 & ~x254 & ~x334 & ~x360 & ~x394 & ~x416 & ~x476 & ~x561 & ~x583 & ~x584 & ~x589 & ~x591 & ~x619 & ~x621 & ~x622 & ~x665 & ~x666 & ~x667 & ~x669 & ~x697 & ~x703 & ~x710 & ~x711 & ~x713 & ~x730 & ~x760 & ~x783;
assign c0152 =  x262 &  x358 &  x386 &  x397 &  x481;
assign c0154 =  x21;
assign c0156 = ~x4 & ~x9 & ~x10 & ~x31 & ~x36 & ~x41 & ~x42 & ~x52 & ~x54 & ~x60 & ~x63 & ~x69 & ~x82 & ~x83 & ~x85 & ~x86 & ~x91 & ~x103 & ~x108 & ~x109 & ~x116 & ~x131 & ~x142 & ~x157 & ~x170 & ~x189 & ~x192 & ~x195 & ~x199 & ~x222 & ~x224 & ~x247 & ~x248 & ~x251 & ~x257 & ~x277 & ~x308 & ~x315 & ~x340 & ~x350 & ~x365 & ~x366 & ~x387 & ~x392 & ~x393 & ~x395 & ~x396 & ~x422 & ~x424 & ~x433 & ~x436 & ~x448 & ~x450 & ~x490 & ~x528 & ~x529 & ~x533 & ~x536 & ~x585 & ~x586 & ~x591 & ~x611 & ~x614 & ~x616 & ~x623 & ~x646 & ~x653 & ~x666 & ~x674 & ~x679 & ~x689 & ~x703 & ~x705 & ~x712 & ~x721 & ~x732 & ~x746 & ~x747 & ~x750 & ~x770 & ~x775 & ~x776 & ~x779;
assign c0158 =  x371 &  x385 &  x399 &  x454 &  x482 &  x483 &  x510 &  x539 &  x567 & ~x3 & ~x22 & ~x36 & ~x55 & ~x65 & ~x68 & ~x78 & ~x101 & ~x103 & ~x109 & ~x118 & ~x124 & ~x132 & ~x146 & ~x165 & ~x166 & ~x171 & ~x174 & ~x192 & ~x250 & ~x251 & ~x257 & ~x283 & ~x284 & ~x307 & ~x312 & ~x340 & ~x364 & ~x367 & ~x388 & ~x448 & ~x449 & ~x475 & ~x530 & ~x563 & ~x639 & ~x666 & ~x694 & ~x702 & ~x704 & ~x716 & ~x729 & ~x744 & ~x746 & ~x755 & ~x760 & ~x763 & ~x781;
assign c0160 =  x538 &  x566 &  x595 & ~x8 & ~x93 & ~x94 & ~x97 & ~x113 & ~x116 & ~x118 & ~x126 & ~x166 & ~x175 & ~x179 & ~x279 & ~x313 & ~x338 & ~x396 & ~x408 & ~x435 & ~x462 & ~x516 & ~x562 & ~x563 & ~x615 & ~x665 & ~x696 & ~x705 & ~x706 & ~x732;
assign c0162 =  x241 &  x427 &  x569 & ~x0 & ~x10 & ~x11 & ~x17 & ~x31 & ~x34 & ~x43 & ~x48 & ~x58 & ~x60 & ~x61 & ~x67 & ~x68 & ~x69 & ~x71 & ~x74 & ~x92 & ~x93 & ~x95 & ~x102 & ~x106 & ~x122 & ~x137 & ~x142 & ~x160 & ~x163 & ~x171 & ~x173 & ~x174 & ~x175 & ~x201 & ~x202 & ~x223 & ~x229 & ~x230 & ~x255 & ~x257 & ~x277 & ~x280 & ~x310 & ~x335 & ~x364 & ~x422 & ~x472 & ~x473 & ~x474 & ~x478 & ~x504 & ~x507 & ~x535 & ~x556 & ~x558 & ~x559 & ~x563 & ~x584 & ~x611 & ~x642 & ~x643 & ~x644 & ~x663 & ~x673 & ~x675 & ~x677 & ~x678 & ~x699 & ~x703 & ~x709 & ~x712 & ~x714 & ~x724 & ~x730 & ~x731 & ~x733 & ~x737 & ~x740 & ~x744 & ~x745 & ~x750 & ~x757 & ~x762 & ~x765 & ~x770 & ~x776 & ~x780;
assign c0164 =  x456 &  x484 & ~x6 & ~x10 & ~x12 & ~x13 & ~x15 & ~x16 & ~x19 & ~x22 & ~x29 & ~x41 & ~x42 & ~x48 & ~x49 & ~x50 & ~x54 & ~x56 & ~x57 & ~x62 & ~x67 & ~x68 & ~x69 & ~x72 & ~x75 & ~x79 & ~x84 & ~x85 & ~x95 & ~x107 & ~x115 & ~x118 & ~x130 & ~x135 & ~x136 & ~x137 & ~x145 & ~x169 & ~x170 & ~x220 & ~x223 & ~x227 & ~x228 & ~x247 & ~x253 & ~x254 & ~x255 & ~x256 & ~x277 & ~x281 & ~x283 & ~x307 & ~x311 & ~x335 & ~x339 & ~x348 & ~x375 & ~x381 & ~x395 & ~x403 & ~x408 & ~x409 & ~x410 & ~x420 & ~x421 & ~x422 & ~x436 & ~x445 & ~x447 & ~x451 & ~x475 & ~x480 & ~x504 & ~x565 & ~x585 & ~x591 & ~x592 & ~x617 & ~x618 & ~x620 & ~x642 & ~x646 & ~x667 & ~x669 & ~x670 & ~x677 & ~x697 & ~x703 & ~x711 & ~x721 & ~x723 & ~x725 & ~x728 & ~x729 & ~x736 & ~x742 & ~x745 & ~x746 & ~x750 & ~x755 & ~x762 & ~x764 & ~x766 & ~x767 & ~x768 & ~x771 & ~x772 & ~x776 & ~x779;
assign c0166 =  x484 &  x541 & ~x2 & ~x7 & ~x8 & ~x10 & ~x19 & ~x22 & ~x23 & ~x30 & ~x31 & ~x35 & ~x38 & ~x39 & ~x44 & ~x48 & ~x51 & ~x52 & ~x54 & ~x56 & ~x57 & ~x62 & ~x65 & ~x68 & ~x69 & ~x80 & ~x83 & ~x84 & ~x87 & ~x88 & ~x92 & ~x93 & ~x99 & ~x103 & ~x105 & ~x113 & ~x116 & ~x117 & ~x137 & ~x140 & ~x142 & ~x143 & ~x168 & ~x169 & ~x191 & ~x198 & ~x221 & ~x224 & ~x250 & ~x277 & ~x280 & ~x281 & ~x283 & ~x305 & ~x307 & ~x311 & ~x321 & ~x322 & ~x337 & ~x349 & ~x350 & ~x363 & ~x364 & ~x376 & ~x378 & ~x393 & ~x396 & ~x405 & ~x406 & ~x419 & ~x420 & ~x423 & ~x432 & ~x450 & ~x460 & ~x461 & ~x464 & ~x476 & ~x479 & ~x491 & ~x502 & ~x504 & ~x506 & ~x508 & ~x516 & ~x530 & ~x534 & ~x557 & ~x558 & ~x588 & ~x589 & ~x618 & ~x620 & ~x622 & ~x643 & ~x644 & ~x645 & ~x646 & ~x650 & ~x651 & ~x652 & ~x653 & ~x668 & ~x670 & ~x671 & ~x674 & ~x681 & ~x682 & ~x694 & ~x698 & ~x700 & ~x703 & ~x710 & ~x711 & ~x714 & ~x715 & ~x716 & ~x717 & ~x720 & ~x726 & ~x727 & ~x731 & ~x735 & ~x736 & ~x737 & ~x738 & ~x739 & ~x740 & ~x741 & ~x742 & ~x745 & ~x746 & ~x760 & ~x762 & ~x764 & ~x768 & ~x770 & ~x774 & ~x775 & ~x778;
assign c0168 =  x364;
assign c0170 =  x657 & ~x17 & ~x41 & ~x42 & ~x71 & ~x72 & ~x77 & ~x82 & ~x87 & ~x89 & ~x107 & ~x110 & ~x139 & ~x140 & ~x144 & ~x148 & ~x171 & ~x174 & ~x194 & ~x201 & ~x220 & ~x229 & ~x230 & ~x285 & ~x322 & ~x335 & ~x419 & ~x434 & ~x490 & ~x518 & ~x530 & ~x563 & ~x588 & ~x665 & ~x671 & ~x711 & ~x742 & ~x756 & ~x757 & ~x761 & ~x773 & ~x774;
assign c0172 =  x239 &  x302 &  x427 & ~x24 & ~x28 & ~x67 & ~x72 & ~x84 & ~x108 & ~x111 & ~x125 & ~x166 & ~x176 & ~x177 & ~x196 & ~x231 & ~x333 & ~x338 & ~x340 & ~x502 & ~x560 & ~x589 & ~x615 & ~x631 & ~x642 & ~x658 & ~x682 & ~x683 & ~x692 & ~x694 & ~x715 & ~x717 & ~x727 & ~x730 & ~x732 & ~x754 & ~x764;
assign c0174 =  x454 &  x652 & ~x7 & ~x150 & ~x461 & ~x543;
assign c0176 = ~x4 & ~x18 & ~x19 & ~x40 & ~x46 & ~x48 & ~x50 & ~x52 & ~x53 & ~x76 & ~x77 & ~x82 & ~x89 & ~x90 & ~x101 & ~x108 & ~x119 & ~x137 & ~x141 & ~x162 & ~x168 & ~x169 & ~x176 & ~x197 & ~x199 & ~x201 & ~x219 & ~x226 & ~x231 & ~x276 & ~x278 & ~x281 & ~x294 & ~x321 & ~x332 & ~x334 & ~x335 & ~x338 & ~x340 & ~x349 & ~x361 & ~x366 & ~x377 & ~x448 & ~x451 & ~x472 & ~x473 & ~x503 & ~x519 & ~x547 & ~x560 & ~x585 & ~x586 & ~x645 & ~x651 & ~x667 & ~x671 & ~x673 & ~x678 & ~x696 & ~x697 & ~x704 & ~x707 & ~x714 & ~x720 & ~x730 & ~x742 & ~x748 & ~x759 & ~x763 & ~x782;
assign c0178 =  x520 & ~x20 & ~x28 & ~x32 & ~x36 & ~x79 & ~x116 & ~x123 & ~x144 & ~x181 & ~x192 & ~x195 & ~x252 & ~x364 & ~x379 & ~x419 & ~x462 & ~x579 & ~x636 & ~x660 & ~x686 & ~x691 & ~x699 & ~x718 & ~x726 & ~x738 & ~x748 & ~x756 & ~x776;
assign c0180 =  x454 & ~x2 & ~x6 & ~x9 & ~x12 & ~x13 & ~x22 & ~x27 & ~x29 & ~x31 & ~x32 & ~x35 & ~x38 & ~x39 & ~x48 & ~x50 & ~x51 & ~x59 & ~x60 & ~x65 & ~x72 & ~x75 & ~x77 & ~x78 & ~x80 & ~x84 & ~x93 & ~x94 & ~x96 & ~x97 & ~x100 & ~x101 & ~x103 & ~x106 & ~x114 & ~x116 & ~x119 & ~x124 & ~x126 & ~x129 & ~x131 & ~x138 & ~x140 & ~x145 & ~x146 & ~x148 & ~x150 & ~x153 & ~x165 & ~x166 & ~x167 & ~x168 & ~x173 & ~x175 & ~x177 & ~x178 & ~x180 & ~x195 & ~x202 & ~x222 & ~x226 & ~x231 & ~x256 & ~x257 & ~x258 & ~x279 & ~x281 & ~x282 & ~x285 & ~x305 & ~x309 & ~x310 & ~x311 & ~x362 & ~x363 & ~x367 & ~x393 & ~x409 & ~x420 & ~x421 & ~x450 & ~x460 & ~x487 & ~x501 & ~x529 & ~x556 & ~x559 & ~x560 & ~x562 & ~x582 & ~x583 & ~x584 & ~x589 & ~x590 & ~x608 & ~x634 & ~x635 & ~x636 & ~x639 & ~x663 & ~x664 & ~x668 & ~x671 & ~x672 & ~x673 & ~x675 & ~x690 & ~x696 & ~x704 & ~x706 & ~x709 & ~x711 & ~x712 & ~x713 & ~x717 & ~x723 & ~x726 & ~x736 & ~x738 & ~x744 & ~x752 & ~x756 & ~x760 & ~x769 & ~x770 & ~x772 & ~x779 & ~x782;
assign c0182 =  x272 &  x373 &  x384 &  x412 &  x455 &  x569 & ~x2 & ~x12 & ~x29 & ~x31 & ~x52 & ~x66 & ~x107 & ~x117 & ~x139 & ~x147 & ~x193 & ~x196 & ~x200 & ~x223 & ~x305 & ~x364 & ~x368 & ~x532 & ~x708 & ~x710 & ~x754 & ~x762 & ~x765 & ~x782;
assign c0184 =  x293 & ~x9 & ~x168 & ~x192 & ~x288 & ~x380 & ~x533 & ~x605 & ~x660 & ~x710 & ~x711 & ~x725 & ~x735;
assign c0186 =  x385 &  x413 & ~x0 & ~x2 & ~x6 & ~x9 & ~x10 & ~x12 & ~x13 & ~x17 & ~x20 & ~x22 & ~x23 & ~x25 & ~x26 & ~x29 & ~x31 & ~x39 & ~x44 & ~x49 & ~x55 & ~x62 & ~x65 & ~x66 & ~x67 & ~x71 & ~x74 & ~x78 & ~x87 & ~x89 & ~x90 & ~x91 & ~x93 & ~x107 & ~x112 & ~x113 & ~x136 & ~x137 & ~x138 & ~x139 & ~x143 & ~x146 & ~x147 & ~x167 & ~x171 & ~x191 & ~x192 & ~x195 & ~x201 & ~x225 & ~x250 & ~x252 & ~x278 & ~x279 & ~x284 & ~x304 & ~x307 & ~x333 & ~x336 & ~x337 & ~x339 & ~x348 & ~x364 & ~x391 & ~x392 & ~x404 & ~x409 & ~x410 & ~x416 & ~x419 & ~x422 & ~x423 & ~x432 & ~x437 & ~x477 & ~x491 & ~x500 & ~x502 & ~x503 & ~x504 & ~x505 & ~x506 & ~x530 & ~x531 & ~x557 & ~x584 & ~x590 & ~x591 & ~x611 & ~x612 & ~x613 & ~x618 & ~x638 & ~x644 & ~x647 & ~x665 & ~x693 & ~x701 & ~x703 & ~x709 & ~x713 & ~x715 & ~x716 & ~x719 & ~x729 & ~x732 & ~x733 & ~x735 & ~x737 & ~x738 & ~x739 & ~x741 & ~x742 & ~x744 & ~x746 & ~x752 & ~x756 & ~x759 & ~x763 & ~x768 & ~x769 & ~x771 & ~x775 & ~x778 & ~x780;
assign c0188 =  x522 &  x627 & ~x58 & ~x69 & ~x71 & ~x114 & ~x118 & ~x149 & ~x165 & ~x226 & ~x250 & ~x306 & ~x337 & ~x349 & ~x377 & ~x405 & ~x417 & ~x460 & ~x463 & ~x587 & ~x690 & ~x691 & ~x712 & ~x714 & ~x737 & ~x763 & ~x765;
assign c0190 =  x369 &  x444;
assign c0192 =  x207 &  x412 &  x570 &  x599 & ~x0 & ~x19 & ~x40 & ~x52 & ~x55 & ~x68 & ~x102 & ~x103 & ~x114 & ~x120 & ~x132 & ~x147 & ~x160 & ~x168 & ~x197 & ~x202 & ~x219 & ~x229 & ~x248 & ~x366 & ~x390 & ~x415 & ~x421 & ~x448 & ~x461 & ~x476 & ~x530 & ~x583 & ~x584 & ~x594 & ~x640 & ~x641 & ~x642 & ~x643 & ~x648 & ~x665 & ~x674 & ~x708 & ~x710 & ~x716 & ~x719 & ~x733 & ~x744 & ~x751 & ~x757 & ~x764 & ~x766;
assign c0194 =  x442 & ~x6 & ~x8 & ~x9 & ~x11 & ~x12 & ~x16 & ~x18 & ~x21 & ~x22 & ~x31 & ~x32 & ~x33 & ~x34 & ~x36 & ~x38 & ~x39 & ~x41 & ~x42 & ~x43 & ~x46 & ~x49 & ~x51 & ~x52 & ~x55 & ~x56 & ~x57 & ~x58 & ~x63 & ~x65 & ~x66 & ~x67 & ~x68 & ~x70 & ~x72 & ~x73 & ~x74 & ~x76 & ~x77 & ~x83 & ~x86 & ~x87 & ~x88 & ~x91 & ~x93 & ~x95 & ~x96 & ~x97 & ~x98 & ~x100 & ~x101 & ~x105 & ~x106 & ~x107 & ~x109 & ~x110 & ~x114 & ~x117 & ~x118 & ~x119 & ~x130 & ~x131 & ~x135 & ~x138 & ~x142 & ~x145 & ~x148 & ~x163 & ~x164 & ~x172 & ~x191 & ~x192 & ~x194 & ~x197 & ~x200 & ~x223 & ~x225 & ~x226 & ~x249 & ~x250 & ~x252 & ~x254 & ~x282 & ~x283 & ~x307 & ~x309 & ~x310 & ~x377 & ~x391 & ~x392 & ~x393 & ~x404 & ~x405 & ~x406 & ~x418 & ~x420 & ~x421 & ~x422 & ~x423 & ~x434 & ~x436 & ~x464 & ~x475 & ~x477 & ~x478 & ~x532 & ~x534 & ~x556 & ~x561 & ~x590 & ~x610 & ~x613 & ~x616 & ~x621 & ~x637 & ~x640 & ~x641 & ~x643 & ~x663 & ~x664 & ~x671 & ~x674 & ~x676 & ~x677 & ~x688 & ~x690 & ~x693 & ~x694 & ~x695 & ~x696 & ~x699 & ~x701 & ~x702 & ~x703 & ~x704 & ~x707 & ~x708 & ~x713 & ~x715 & ~x716 & ~x717 & ~x720 & ~x725 & ~x726 & ~x727 & ~x728 & ~x729 & ~x730 & ~x732 & ~x739 & ~x740 & ~x741 & ~x745 & ~x750 & ~x751 & ~x753 & ~x757 & ~x759 & ~x760 & ~x764 & ~x770 & ~x778 & ~x779 & ~x782;
assign c0196 =  x330 &  x399 &  x414;
assign c0198 =  x456 &  x485 &  x512 &  x629 & ~x3 & ~x38 & ~x39 & ~x45 & ~x62 & ~x88 & ~x89 & ~x96 & ~x97 & ~x103 & ~x108 & ~x110 & ~x111 & ~x112 & ~x138 & ~x167 & ~x199 & ~x225 & ~x308 & ~x309 & ~x340 & ~x369 & ~x420 & ~x421 & ~x436 & ~x463 & ~x503 & ~x516 & ~x531 & ~x558 & ~x721 & ~x733 & ~x738 & ~x743 & ~x747 & ~x765 & ~x772 & ~x779 & ~x782;
assign c0200 =  x65;
assign c0202 =  x624 & ~x149 & ~x179 & ~x180 & ~x204 & ~x341 & ~x378 & ~x515;
assign c0204 =  x346 &  x514 & ~x7 & ~x20 & ~x130 & ~x131 & ~x134 & ~x139 & ~x145 & ~x172 & ~x201 & ~x222 & ~x281 & ~x357 & ~x427 & ~x483 & ~x502 & ~x531 & ~x539 & ~x590 & ~x623 & ~x647 & ~x710 & ~x751;
assign c0206 =  x268 &  x403 &  x431 &  x514 & ~x3 & ~x10 & ~x22 & ~x27 & ~x28 & ~x56 & ~x57 & ~x60 & ~x63 & ~x66 & ~x67 & ~x70 & ~x74 & ~x85 & ~x102 & ~x110 & ~x116 & ~x136 & ~x145 & ~x162 & ~x167 & ~x222 & ~x231 & ~x247 & ~x251 & ~x256 & ~x280 & ~x284 & ~x396 & ~x417 & ~x422 & ~x448 & ~x450 & ~x451 & ~x461 & ~x501 & ~x562 & ~x586 & ~x610 & ~x637 & ~x642 & ~x645 & ~x646 & ~x688 & ~x690 & ~x695 & ~x699 & ~x704 & ~x708 & ~x711 & ~x714 & ~x718 & ~x719 & ~x722 & ~x744 & ~x747 & ~x748 & ~x756 & ~x758 & ~x765 & ~x771 & ~x783;
assign c0208 =  x345 &  x485 &  x577 &  x655 & ~x258 & ~x453;
assign c0210 =  x238 & ~x13 & ~x16 & ~x18 & ~x21 & ~x23 & ~x24 & ~x26 & ~x29 & ~x33 & ~x36 & ~x42 & ~x46 & ~x51 & ~x52 & ~x53 & ~x56 & ~x59 & ~x64 & ~x65 & ~x67 & ~x70 & ~x71 & ~x79 & ~x88 & ~x89 & ~x93 & ~x95 & ~x97 & ~x98 & ~x100 & ~x102 & ~x103 & ~x104 & ~x105 & ~x106 & ~x107 & ~x109 & ~x110 & ~x114 & ~x116 & ~x117 & ~x119 & ~x124 & ~x125 & ~x127 & ~x129 & ~x130 & ~x133 & ~x135 & ~x137 & ~x139 & ~x142 & ~x145 & ~x162 & ~x164 & ~x169 & ~x170 & ~x172 & ~x190 & ~x192 & ~x193 & ~x194 & ~x195 & ~x197 & ~x198 & ~x200 & ~x228 & ~x247 & ~x250 & ~x251 & ~x253 & ~x278 & ~x281 & ~x284 & ~x311 & ~x312 & ~x333 & ~x334 & ~x335 & ~x338 & ~x360 & ~x366 & ~x381 & ~x389 & ~x391 & ~x392 & ~x408 & ~x409 & ~x418 & ~x419 & ~x420 & ~x447 & ~x450 & ~x451 & ~x474 & ~x477 & ~x479 & ~x503 & ~x504 & ~x506 & ~x518 & ~x531 & ~x533 & ~x556 & ~x557 & ~x561 & ~x562 & ~x583 & ~x589 & ~x590 & ~x610 & ~x614 & ~x616 & ~x620 & ~x639 & ~x643 & ~x647 & ~x665 & ~x666 & ~x668 & ~x669 & ~x675 & ~x689 & ~x690 & ~x692 & ~x694 & ~x697 & ~x699 & ~x705 & ~x709 & ~x710 & ~x714 & ~x717 & ~x718 & ~x719 & ~x720 & ~x721 & ~x722 & ~x730 & ~x732 & ~x737 & ~x740 & ~x742 & ~x743 & ~x745 & ~x746 & ~x747 & ~x748 & ~x750 & ~x752 & ~x755 & ~x757 & ~x768 & ~x769 & ~x775 & ~x776 & ~x777 & ~x778 & ~x782 & ~x783;
assign c0212 =  x321 &  x411 & ~x0 & ~x126 & ~x173 & ~x179 & ~x337 & ~x366 & ~x392 & ~x396 & ~x664 & ~x714 & ~x729 & ~x737 & ~x742 & ~x757 & ~x777;
assign c0214 =  x616;
assign c0216 =  x493 & ~x7 & ~x11 & ~x13 & ~x14 & ~x16 & ~x23 & ~x25 & ~x26 & ~x30 & ~x37 & ~x44 & ~x49 & ~x51 & ~x60 & ~x65 & ~x66 & ~x67 & ~x72 & ~x75 & ~x76 & ~x77 & ~x78 & ~x82 & ~x94 & ~x95 & ~x99 & ~x101 & ~x107 & ~x109 & ~x113 & ~x115 & ~x123 & ~x124 & ~x136 & ~x141 & ~x143 & ~x146 & ~x149 & ~x166 & ~x171 & ~x173 & ~x174 & ~x176 & ~x177 & ~x192 & ~x197 & ~x199 & ~x200 & ~x221 & ~x225 & ~x226 & ~x227 & ~x230 & ~x250 & ~x254 & ~x256 & ~x260 & ~x261 & ~x277 & ~x288 & ~x289 & ~x306 & ~x308 & ~x314 & ~x331 & ~x337 & ~x340 & ~x362 & ~x363 & ~x364 & ~x367 & ~x371 & ~x387 & ~x394 & ~x396 & ~x418 & ~x422 & ~x443 & ~x453 & ~x471 & ~x478 & ~x499 & ~x505 & ~x507 & ~x525 & ~x528 & ~x529 & ~x536 & ~x555 & ~x559 & ~x580 & ~x582 & ~x584 & ~x586 & ~x592 & ~x606 & ~x613 & ~x615 & ~x617 & ~x619 & ~x620 & ~x633 & ~x634 & ~x636 & ~x637 & ~x641 & ~x642 & ~x644 & ~x645 & ~x660 & ~x664 & ~x666 & ~x667 & ~x669 & ~x677 & ~x693 & ~x706 & ~x710 & ~x712 & ~x714 & ~x718 & ~x719 & ~x729 & ~x734 & ~x738 & ~x743 & ~x746 & ~x750 & ~x755 & ~x762 & ~x765 & ~x770 & ~x773 & ~x779 & ~x783;
assign c0218 =  x342 &  x369 &  x386 &  x397 &  x414 &  x482 & ~x436;
assign c0220 =  x375 &  x404 &  x432 &  x437 & ~x368 & ~x406 & ~x441 & ~x497 & ~x502 & ~x553 & ~x567 & ~x682;
assign c0222 =  x748;
assign c0224 =  x186 & ~x4 & ~x9 & ~x12 & ~x36 & ~x78 & ~x125 & ~x143 & ~x175 & ~x201 & ~x253 & ~x312 & ~x325 & ~x337 & ~x380 & ~x407 & ~x408 & ~x435 & ~x527 & ~x545 & ~x583 & ~x612 & ~x636 & ~x643 & ~x646 & ~x662 & ~x673 & ~x702 & ~x707 & ~x728 & ~x742;
assign c0226 =  x217 &  x302 &  x399 &  x454 &  x566 & ~x54 & ~x423 & ~x608 & ~x669;
assign c0228 =  x213 &  x355 &  x438 &  x627 & ~x26 & ~x76 & ~x91 & ~x121 & ~x124 & ~x140 & ~x164 & ~x168 & ~x177 & ~x192 & ~x204 & ~x234 & ~x256 & ~x285 & ~x288 & ~x340 & ~x418 & ~x442 & ~x447 & ~x479 & ~x501 & ~x505 & ~x528 & ~x535 & ~x537 & ~x580 & ~x588 & ~x660 & ~x689 & ~x694 & ~x716 & ~x723 & ~x735 & ~x749 & ~x764 & ~x767;
assign c0230 = ~x1 & ~x10 & ~x12 & ~x13 & ~x14 & ~x18 & ~x19 & ~x20 & ~x23 & ~x25 & ~x31 & ~x34 & ~x38 & ~x42 & ~x47 & ~x48 & ~x50 & ~x51 & ~x54 & ~x55 & ~x56 & ~x57 & ~x59 & ~x60 & ~x61 & ~x62 & ~x65 & ~x67 & ~x68 & ~x70 & ~x71 & ~x75 & ~x80 & ~x84 & ~x86 & ~x87 & ~x88 & ~x89 & ~x106 & ~x108 & ~x109 & ~x110 & ~x113 & ~x116 & ~x119 & ~x120 & ~x136 & ~x138 & ~x140 & ~x141 & ~x145 & ~x146 & ~x148 & ~x166 & ~x168 & ~x174 & ~x192 & ~x194 & ~x195 & ~x197 & ~x199 & ~x200 & ~x201 & ~x203 & ~x221 & ~x222 & ~x225 & ~x226 & ~x227 & ~x250 & ~x277 & ~x279 & ~x280 & ~x305 & ~x306 & ~x308 & ~x310 & ~x323 & ~x324 & ~x338 & ~x350 & ~x351 & ~x352 & ~x353 & ~x364 & ~x366 & ~x368 & ~x378 & ~x379 & ~x380 & ~x381 & ~x395 & ~x407 & ~x409 & ~x418 & ~x422 & ~x432 & ~x433 & ~x434 & ~x447 & ~x451 & ~x460 & ~x461 & ~x462 & ~x463 & ~x464 & ~x473 & ~x477 & ~x488 & ~x489 & ~x490 & ~x501 & ~x505 & ~x506 & ~x517 & ~x531 & ~x533 & ~x534 & ~x557 & ~x560 & ~x561 & ~x562 & ~x583 & ~x586 & ~x587 & ~x590 & ~x611 & ~x614 & ~x617 & ~x619 & ~x620 & ~x621 & ~x637 & ~x638 & ~x641 & ~x642 & ~x645 & ~x646 & ~x648 & ~x663 & ~x668 & ~x671 & ~x674 & ~x675 & ~x676 & ~x677 & ~x690 & ~x691 & ~x693 & ~x694 & ~x696 & ~x697 & ~x700 & ~x701 & ~x702 & ~x704 & ~x706 & ~x707 & ~x708 & ~x709 & ~x710 & ~x712 & ~x713 & ~x714 & ~x716 & ~x717 & ~x718 & ~x719 & ~x720 & ~x721 & ~x722 & ~x723 & ~x727 & ~x731 & ~x732 & ~x733 & ~x735 & ~x740 & ~x742 & ~x746 & ~x749 & ~x753 & ~x754 & ~x755 & ~x757 & ~x759 & ~x762 & ~x763 & ~x764 & ~x765 & ~x766 & ~x772 & ~x773 & ~x775 & ~x781 & ~x782 & ~x783;
assign c0232 =  x626 & ~x50 & ~x53 & ~x87 & ~x89 & ~x249 & ~x338 & ~x378 & ~x516 & ~x524 & ~x552 & ~x561 & ~x605 & ~x632 & ~x671 & ~x680 & ~x740;
assign c0234 =  x356 &  x629 &  x632 & ~x28 & ~x45 & ~x49 & ~x54 & ~x65 & ~x72 & ~x76 & ~x78 & ~x119 & ~x138 & ~x159 & ~x246 & ~x275 & ~x283 & ~x311 & ~x338 & ~x387 & ~x389 & ~x448 & ~x463 & ~x503 & ~x557 & ~x562 & ~x584 & ~x585 & ~x586 & ~x642 & ~x666 & ~x673 & ~x676 & ~x731 & ~x770;
assign c0236 =  x3;
assign c0238 =  x557;
assign c0240 =  x627 & ~x28 & ~x29 & ~x41 & ~x59 & ~x114 & ~x115 & ~x152 & ~x163 & ~x165 & ~x167 & ~x200 & ~x229 & ~x260 & ~x306 & ~x311 & ~x336 & ~x337 & ~x419 & ~x462 & ~x524 & ~x557 & ~x558 & ~x641 & ~x647 & ~x662 & ~x669 & ~x677 & ~x701 & ~x709 & ~x713 & ~x716 & ~x730 & ~x745;
assign c0242 =  x328 &  x384 &  x412 &  x429 &  x457 &  x484 & ~x1 & ~x2 & ~x6 & ~x7 & ~x16 & ~x18 & ~x20 & ~x23 & ~x25 & ~x27 & ~x34 & ~x43 & ~x49 & ~x50 & ~x52 & ~x59 & ~x65 & ~x72 & ~x73 & ~x74 & ~x80 & ~x82 & ~x96 & ~x98 & ~x105 & ~x106 & ~x111 & ~x112 & ~x114 & ~x117 & ~x120 & ~x134 & ~x135 & ~x138 & ~x143 & ~x144 & ~x146 & ~x162 & ~x173 & ~x175 & ~x191 & ~x196 & ~x200 & ~x226 & ~x276 & ~x277 & ~x278 & ~x280 & ~x283 & ~x284 & ~x304 & ~x306 & ~x334 & ~x335 & ~x362 & ~x363 & ~x389 & ~x390 & ~x393 & ~x417 & ~x420 & ~x446 & ~x447 & ~x451 & ~x473 & ~x476 & ~x477 & ~x501 & ~x508 & ~x534 & ~x536 & ~x537 & ~x556 & ~x561 & ~x563 & ~x583 & ~x587 & ~x588 & ~x589 & ~x615 & ~x617 & ~x618 & ~x619 & ~x620 & ~x642 & ~x647 & ~x648 & ~x649 & ~x666 & ~x669 & ~x671 & ~x677 & ~x689 & ~x695 & ~x700 & ~x701 & ~x709 & ~x710 & ~x711 & ~x713 & ~x717 & ~x724 & ~x732 & ~x734 & ~x736 & ~x739 & ~x741 & ~x743 & ~x745 & ~x749 & ~x765 & ~x766 & ~x768 & ~x769 & ~x773 & ~x776 & ~x781;
assign c0244 = ~x0 & ~x3 & ~x6 & ~x12 & ~x21 & ~x22 & ~x35 & ~x36 & ~x66 & ~x75 & ~x88 & ~x94 & ~x99 & ~x102 & ~x104 & ~x113 & ~x117 & ~x136 & ~x144 & ~x147 & ~x149 & ~x151 & ~x161 & ~x166 & ~x217 & ~x222 & ~x229 & ~x230 & ~x251 & ~x279 & ~x301 & ~x341 & ~x357 & ~x362 & ~x367 & ~x390 & ~x395 & ~x406 & ~x415 & ~x445 & ~x447 & ~x497 & ~x502 & ~x534 & ~x553 & ~x579 & ~x594 & ~x609 & ~x611 & ~x635 & ~x640 & ~x647 & ~x648 & ~x650 & ~x660 & ~x662 & ~x674 & ~x679 & ~x693 & ~x704 & ~x714 & ~x717 & ~x739 & ~x742 & ~x750;
assign c0246 =  x245 &  x347 &  x429 &  x596 & ~x139 & ~x176 & ~x361 & ~x683;
assign c0248 =  x348 &  x512 & ~x11 & ~x452 & ~x475 & ~x579 & ~x605 & ~x619;
assign c0250 =  x218 &  x330 &  x537 & ~x179 & ~x606;
assign c0252 =  x243 &  x328 &  x356 &  x457 &  x569 & ~x1 & ~x16 & ~x21 & ~x28 & ~x32 & ~x33 & ~x48 & ~x54 & ~x56 & ~x76 & ~x83 & ~x102 & ~x109 & ~x114 & ~x119 & ~x140 & ~x143 & ~x164 & ~x166 & ~x172 & ~x173 & ~x199 & ~x201 & ~x223 & ~x227 & ~x251 & ~x252 & ~x256 & ~x303 & ~x305 & ~x332 & ~x333 & ~x340 & ~x392 & ~x393 & ~x394 & ~x419 & ~x422 & ~x445 & ~x531 & ~x555 & ~x560 & ~x589 & ~x609 & ~x639 & ~x643 & ~x645 & ~x646 & ~x665 & ~x667 & ~x676 & ~x693 & ~x703 & ~x705 & ~x709 & ~x720 & ~x723 & ~x726 & ~x728 & ~x729 & ~x731 & ~x737 & ~x743 & ~x744 & ~x750 & ~x751 & ~x754 & ~x755 & ~x783;
assign c0254 =  x295 & ~x16 & ~x48 & ~x53 & ~x57 & ~x91 & ~x94 & ~x95 & ~x106 & ~x112 & ~x125 & ~x138 & ~x170 & ~x175 & ~x222 & ~x224 & ~x234 & ~x344 & ~x366 & ~x420 & ~x451 & ~x471 & ~x523 & ~x551 & ~x558 & ~x634 & ~x648 & ~x676 & ~x714 & ~x734;
assign c0256 =  x400 &  x569 & ~x29 & ~x30 & ~x125 & ~x226 & ~x338 & ~x497 & ~x580 & ~x608 & ~x637 & ~x657 & ~x669 & ~x683 & ~x697 & ~x700 & ~x718 & ~x733 & ~x743;
assign c0258 =  x330 &  x427 &  x565;
assign c0260 =  x189 &  x246 &  x302 &  x330 &  x358 &  x386;
assign c0262 = ~x1 & ~x7 & ~x12 & ~x13 & ~x14 & ~x15 & ~x21 & ~x27 & ~x28 & ~x32 & ~x34 & ~x36 & ~x37 & ~x38 & ~x42 & ~x43 & ~x45 & ~x51 & ~x52 & ~x55 & ~x60 & ~x74 & ~x75 & ~x78 & ~x80 & ~x87 & ~x91 & ~x96 & ~x103 & ~x110 & ~x112 & ~x118 & ~x138 & ~x165 & ~x167 & ~x171 & ~x174 & ~x193 & ~x196 & ~x199 & ~x201 & ~x222 & ~x224 & ~x228 & ~x252 & ~x255 & ~x256 & ~x279 & ~x298 & ~x311 & ~x325 & ~x326 & ~x334 & ~x336 & ~x340 & ~x376 & ~x391 & ~x394 & ~x395 & ~x408 & ~x409 & ~x410 & ~x411 & ~x422 & ~x432 & ~x436 & ~x437 & ~x447 & ~x459 & ~x462 & ~x463 & ~x464 & ~x465 & ~x487 & ~x489 & ~x490 & ~x491 & ~x492 & ~x506 & ~x515 & ~x516 & ~x519 & ~x529 & ~x531 & ~x532 & ~x543 & ~x544 & ~x558 & ~x561 & ~x583 & ~x586 & ~x613 & ~x615 & ~x618 & ~x620 & ~x639 & ~x647 & ~x667 & ~x691 & ~x693 & ~x699 & ~x700 & ~x709 & ~x711 & ~x712 & ~x713 & ~x716 & ~x718 & ~x719 & ~x724 & ~x726 & ~x729 & ~x730 & ~x734 & ~x743 & ~x745 & ~x749 & ~x750 & ~x755 & ~x762 & ~x763 & ~x765 & ~x769 & ~x771 & ~x778 & ~x780 & ~x783;
assign c0264 =  x644;
assign c0266 = ~x18 & ~x38 & ~x50 & ~x51 & ~x80 & ~x138 & ~x139 & ~x166 & ~x167 & ~x221 & ~x223 & ~x228 & ~x255 & ~x267 & ~x279 & ~x294 & ~x320 & ~x321 & ~x322 & ~x335 & ~x339 & ~x349 & ~x352 & ~x353 & ~x381 & ~x393 & ~x403 & ~x408 & ~x423 & ~x437 & ~x438 & ~x464 & ~x465 & ~x473 & ~x489 & ~x490 & ~x491 & ~x493 & ~x520 & ~x547 & ~x548 & ~x589 & ~x614 & ~x620 & ~x701 & ~x711 & ~x714 & ~x716 & ~x724 & ~x727 & ~x728 & ~x765 & ~x766 & ~x774;
assign c0268 = ~x4 & ~x5 & ~x20 & ~x25 & ~x28 & ~x29 & ~x32 & ~x42 & ~x53 & ~x55 & ~x59 & ~x61 & ~x65 & ~x67 & ~x69 & ~x71 & ~x74 & ~x76 & ~x80 & ~x81 & ~x83 & ~x89 & ~x90 & ~x92 & ~x95 & ~x100 & ~x104 & ~x105 & ~x107 & ~x113 & ~x115 & ~x118 & ~x121 & ~x138 & ~x139 & ~x140 & ~x144 & ~x150 & ~x165 & ~x167 & ~x170 & ~x200 & ~x201 & ~x202 & ~x220 & ~x222 & ~x224 & ~x229 & ~x232 & ~x249 & ~x251 & ~x253 & ~x257 & ~x258 & ~x277 & ~x281 & ~x282 & ~x284 & ~x286 & ~x306 & ~x311 & ~x332 & ~x336 & ~x353 & ~x365 & ~x390 & ~x407 & ~x419 & ~x443 & ~x446 & ~x451 & ~x476 & ~x477 & ~x499 & ~x500 & ~x501 & ~x505 & ~x528 & ~x529 & ~x532 & ~x534 & ~x552 & ~x553 & ~x580 & ~x583 & ~x584 & ~x586 & ~x587 & ~x608 & ~x610 & ~x620 & ~x635 & ~x642 & ~x643 & ~x645 & ~x648 & ~x649 & ~x660 & ~x666 & ~x672 & ~x677 & ~x687 & ~x691 & ~x695 & ~x698 & ~x701 & ~x707 & ~x713 & ~x716 & ~x721 & ~x737 & ~x746 & ~x748 & ~x750 & ~x753 & ~x759 & ~x763 & ~x764 & ~x765 & ~x767 & ~x776 & ~x778 & ~x779 & ~x780 & ~x783;
assign c0270 =  x272 &  x328 &  x356 &  x440 & ~x9 & ~x21 & ~x30 & ~x34 & ~x51 & ~x62 & ~x66 & ~x73 & ~x74 & ~x105 & ~x115 & ~x134 & ~x147 & ~x168 & ~x197 & ~x246 & ~x258 & ~x277 & ~x278 & ~x365 & ~x388 & ~x552 & ~x555 & ~x637 & ~x689 & ~x697 & ~x715 & ~x734 & ~x758;
assign c0272 =  x324 &  x357 &  x399 &  x400 &  x413 &  x427 &  x441 &  x482 &  x484 &  x512;
assign c0274 =  x181 & ~x6 & ~x9 & ~x37 & ~x48 & ~x53 & ~x54 & ~x58 & ~x101 & ~x109 & ~x119 & ~x140 & ~x167 & ~x169 & ~x170 & ~x175 & ~x192 & ~x193 & ~x274 & ~x305 & ~x310 & ~x334 & ~x351 & ~x363 & ~x421 & ~x425 & ~x435 & ~x462 & ~x478 & ~x491 & ~x505 & ~x531 & ~x565 & ~x567 & ~x592 & ~x613 & ~x642 & ~x647 & ~x650 & ~x651 & ~x670 & ~x672 & ~x679 & ~x690 & ~x696 & ~x697 & ~x707 & ~x713 & ~x724 & ~x744 & ~x752 & ~x762 & ~x779;
assign c0276 =  x239 &  x266 &  x295 &  x357 &  x511 & ~x12 & ~x14 & ~x21 & ~x35 & ~x37 & ~x42 & ~x57 & ~x71 & ~x77 & ~x84 & ~x89 & ~x94 & ~x100 & ~x102 & ~x104 & ~x105 & ~x107 & ~x115 & ~x134 & ~x135 & ~x140 & ~x143 & ~x149 & ~x165 & ~x202 & ~x222 & ~x257 & ~x276 & ~x277 & ~x282 & ~x307 & ~x310 & ~x311 & ~x334 & ~x337 & ~x338 & ~x362 & ~x419 & ~x447 & ~x474 & ~x475 & ~x507 & ~x533 & ~x534 & ~x558 & ~x585 & ~x641 & ~x642 & ~x646 & ~x662 & ~x665 & ~x666 & ~x688 & ~x693 & ~x694 & ~x703 & ~x708 & ~x713 & ~x715 & ~x717 & ~x718 & ~x723 & ~x741 & ~x758 & ~x769 & ~x770;
assign c0278 = ~x17 & ~x38 & ~x39 & ~x42 & ~x53 & ~x69 & ~x79 & ~x88 & ~x93 & ~x192 & ~x255 & ~x274 & ~x282 & ~x324 & ~x379 & ~x380 & ~x396 & ~x475 & ~x481 & ~x490 & ~x505 & ~x555 & ~x641 & ~x732 & ~x734 & ~x743 & ~x783;
assign c0280 =  x315 &  x427 &  x470 &  x498 &  x553 & ~x2 & ~x4 & ~x18 & ~x22 & ~x27 & ~x44 & ~x52 & ~x53 & ~x54 & ~x58 & ~x63 & ~x70 & ~x71 & ~x89 & ~x94 & ~x104 & ~x109 & ~x118 & ~x119 & ~x134 & ~x163 & ~x166 & ~x223 & ~x253 & ~x254 & ~x279 & ~x333 & ~x339 & ~x377 & ~x391 & ~x405 & ~x407 & ~x420 & ~x422 & ~x463 & ~x501 & ~x502 & ~x558 & ~x617 & ~x639 & ~x642 & ~x674 & ~x676 & ~x693 & ~x694 & ~x703 & ~x717 & ~x718 & ~x720 & ~x729 & ~x740 & ~x742 & ~x746 & ~x752 & ~x756 & ~x764 & ~x773 & ~x774;
assign c0282 =  x211 &  x239 &  x240 &  x241 &  x415 & ~x0 & ~x2 & ~x9 & ~x10 & ~x20 & ~x21 & ~x29 & ~x34 & ~x35 & ~x66 & ~x68 & ~x70 & ~x74 & ~x91 & ~x92 & ~x96 & ~x116 & ~x118 & ~x119 & ~x126 & ~x143 & ~x170 & ~x221 & ~x250 & ~x367 & ~x393 & ~x395 & ~x409 & ~x421 & ~x436 & ~x437 & ~x447 & ~x461 & ~x462 & ~x464 & ~x465 & ~x466 & ~x477 & ~x488 & ~x506 & ~x561 & ~x645 & ~x668 & ~x670 & ~x698 & ~x707 & ~x717 & ~x721 & ~x736 & ~x748 & ~x749 & ~x750 & ~x753 & ~x764 & ~x778;
assign c0284 =  x331 &  x387 &  x415 & ~x0 & ~x2 & ~x25 & ~x29 & ~x63 & ~x94 & ~x97 & ~x108 & ~x114 & ~x115 & ~x121 & ~x123 & ~x124 & ~x137 & ~x165 & ~x177 & ~x252 & ~x309 & ~x326 & ~x327 & ~x333 & ~x336 & ~x354 & ~x355 & ~x394 & ~x408 & ~x421 & ~x436 & ~x437 & ~x464 & ~x531 & ~x612 & ~x613 & ~x639 & ~x673 & ~x697 & ~x716 & ~x731 & ~x773;
assign c0286 =  x288 &  x399 &  x427 &  x484 &  x512 &  x569 &  x598 &  x627 &  x657 & ~x0 & ~x6 & ~x10 & ~x11 & ~x13 & ~x14 & ~x22 & ~x27 & ~x32 & ~x34 & ~x36 & ~x41 & ~x42 & ~x50 & ~x51 & ~x55 & ~x64 & ~x70 & ~x71 & ~x74 & ~x78 & ~x80 & ~x82 & ~x83 & ~x94 & ~x96 & ~x97 & ~x99 & ~x108 & ~x113 & ~x134 & ~x136 & ~x145 & ~x164 & ~x167 & ~x170 & ~x193 & ~x221 & ~x222 & ~x254 & ~x255 & ~x256 & ~x279 & ~x284 & ~x308 & ~x309 & ~x312 & ~x335 & ~x336 & ~x337 & ~x362 & ~x368 & ~x392 & ~x394 & ~x395 & ~x396 & ~x421 & ~x446 & ~x451 & ~x462 & ~x473 & ~x475 & ~x479 & ~x503 & ~x504 & ~x530 & ~x532 & ~x535 & ~x557 & ~x562 & ~x584 & ~x587 & ~x588 & ~x590 & ~x591 & ~x592 & ~x616 & ~x617 & ~x618 & ~x645 & ~x646 & ~x650 & ~x665 & ~x673 & ~x677 & ~x693 & ~x708 & ~x716 & ~x719 & ~x723 & ~x725 & ~x731 & ~x732 & ~x733 & ~x737 & ~x739 & ~x740 & ~x743 & ~x745 & ~x746 & ~x750 & ~x752 & ~x759 & ~x767 & ~x768 & ~x770 & ~x773 & ~x776 & ~x778 & ~x781 & ~x782 & ~x783;
assign c0288 =  x358 & ~x0 & ~x8 & ~x17 & ~x20 & ~x23 & ~x24 & ~x25 & ~x31 & ~x32 & ~x37 & ~x38 & ~x39 & ~x41 & ~x47 & ~x50 & ~x53 & ~x54 & ~x62 & ~x65 & ~x66 & ~x68 & ~x76 & ~x78 & ~x81 & ~x82 & ~x87 & ~x89 & ~x96 & ~x105 & ~x111 & ~x120 & ~x125 & ~x132 & ~x136 & ~x137 & ~x139 & ~x148 & ~x162 & ~x165 & ~x167 & ~x170 & ~x193 & ~x196 & ~x221 & ~x225 & ~x228 & ~x249 & ~x250 & ~x252 & ~x279 & ~x281 & ~x282 & ~x284 & ~x306 & ~x333 & ~x335 & ~x350 & ~x352 & ~x361 & ~x381 & ~x395 & ~x406 & ~x407 & ~x410 & ~x411 & ~x433 & ~x434 & ~x448 & ~x449 & ~x461 & ~x502 & ~x504 & ~x531 & ~x557 & ~x558 & ~x585 & ~x612 & ~x614 & ~x615 & ~x619 & ~x620 & ~x641 & ~x646 & ~x647 & ~x665 & ~x666 & ~x667 & ~x672 & ~x673 & ~x693 & ~x694 & ~x705 & ~x710 & ~x714 & ~x715 & ~x724 & ~x725 & ~x730 & ~x737 & ~x738 & ~x742 & ~x745 & ~x746 & ~x748 & ~x757 & ~x761 & ~x772 & ~x773 & ~x779 & ~x781;
assign c0290 =  x154 &  x629 & ~x2 & ~x6 & ~x10 & ~x18 & ~x32 & ~x51 & ~x58 & ~x61 & ~x62 & ~x67 & ~x88 & ~x92 & ~x102 & ~x103 & ~x111 & ~x118 & ~x119 & ~x120 & ~x144 & ~x164 & ~x172 & ~x190 & ~x192 & ~x198 & ~x277 & ~x293 & ~x308 & ~x320 & ~x375 & ~x390 & ~x403 & ~x421 & ~x473 & ~x475 & ~x519 & ~x520 & ~x546 & ~x586 & ~x640 & ~x641 & ~x708 & ~x729 & ~x734 & ~x740 & ~x751 & ~x771 & ~x783;
assign c0292 =  x244 &  x357 &  x371 &  x385 &  x482 &  x510 &  x597 & ~x5 & ~x6 & ~x31 & ~x52 & ~x66 & ~x75 & ~x136 & ~x194 & ~x224 & ~x476 & ~x533 & ~x676 & ~x738 & ~x747;
assign c0294 =  x270 &  x357 &  x455 & ~x0 & ~x1 & ~x5 & ~x7 & ~x11 & ~x12 & ~x14 & ~x22 & ~x24 & ~x36 & ~x48 & ~x61 & ~x65 & ~x66 & ~x70 & ~x75 & ~x78 & ~x84 & ~x89 & ~x90 & ~x96 & ~x101 & ~x102 & ~x103 & ~x111 & ~x115 & ~x117 & ~x132 & ~x135 & ~x170 & ~x221 & ~x223 & ~x224 & ~x227 & ~x228 & ~x279 & ~x305 & ~x312 & ~x336 & ~x338 & ~x362 & ~x389 & ~x394 & ~x407 & ~x420 & ~x424 & ~x434 & ~x446 & ~x451 & ~x474 & ~x477 & ~x479 & ~x507 & ~x533 & ~x536 & ~x557 & ~x584 & ~x589 & ~x612 & ~x614 & ~x616 & ~x617 & ~x618 & ~x619 & ~x638 & ~x645 & ~x667 & ~x668 & ~x676 & ~x677 & ~x680 & ~x691 & ~x692 & ~x694 & ~x698 & ~x702 & ~x706 & ~x707 & ~x711 & ~x716 & ~x717 & ~x719 & ~x720 & ~x722 & ~x723 & ~x726 & ~x731 & ~x751 & ~x755 & ~x756 & ~x759 & ~x762 & ~x765 & ~x768 & ~x771 & ~x773 & ~x782;
assign c0296 =  x628 &  x698 & ~x26 & ~x134 & ~x168 & ~x190 & ~x363 & ~x612 & ~x677;
assign c0298 =  x453 & ~x5 & ~x15 & ~x21 & ~x25 & ~x26 & ~x28 & ~x29 & ~x31 & ~x37 & ~x57 & ~x64 & ~x73 & ~x78 & ~x90 & ~x93 & ~x95 & ~x96 & ~x109 & ~x110 & ~x112 & ~x117 & ~x123 & ~x134 & ~x142 & ~x148 & ~x163 & ~x168 & ~x172 & ~x200 & ~x226 & ~x250 & ~x251 & ~x280 & ~x308 & ~x333 & ~x363 & ~x382 & ~x405 & ~x408 & ~x410 & ~x411 & ~x422 & ~x431 & ~x434 & ~x436 & ~x437 & ~x438 & ~x447 & ~x451 & ~x459 & ~x461 & ~x463 & ~x477 & ~x488 & ~x502 & ~x504 & ~x506 & ~x531 & ~x556 & ~x559 & ~x562 & ~x583 & ~x612 & ~x637 & ~x641 & ~x666 & ~x676 & ~x685 & ~x686 & ~x689 & ~x691 & ~x694 & ~x698 & ~x700 & ~x703 & ~x706 & ~x716 & ~x717 & ~x718 & ~x730 & ~x732 & ~x743 & ~x745 & ~x748 & ~x750 & ~x752 & ~x756 & ~x765 & ~x768 & ~x769 & ~x775 & ~x778;
assign c01 =  x719;
assign c03 =  x489 &  x519 & ~x12 & ~x29 & ~x35 & ~x36 & ~x45 & ~x54 & ~x68 & ~x71 & ~x117 & ~x171 & ~x174 & ~x197 & ~x229 & ~x231 & ~x250 & ~x256 & ~x260 & ~x287 & ~x328 & ~x330 & ~x334 & ~x475 & ~x503 & ~x505 & ~x584 & ~x614 & ~x617 & ~x704 & ~x719 & ~x730 & ~x768;
assign c05 =  x529;
assign c07 = ~x156 & ~x235 & ~x571 & ~x596;
assign c09 = ~x1 & ~x3 & ~x9 & ~x13 & ~x16 & ~x18 & ~x19 & ~x20 & ~x24 & ~x28 & ~x31 & ~x32 & ~x33 & ~x35 & ~x36 & ~x39 & ~x51 & ~x54 & ~x64 & ~x70 & ~x73 & ~x79 & ~x82 & ~x89 & ~x109 & ~x110 & ~x138 & ~x140 & ~x142 & ~x143 & ~x144 & ~x164 & ~x165 & ~x166 & ~x170 & ~x194 & ~x199 & ~x226 & ~x252 & ~x254 & ~x255 & ~x256 & ~x275 & ~x280 & ~x282 & ~x283 & ~x285 & ~x286 & ~x287 & ~x304 & ~x306 & ~x307 & ~x311 & ~x313 & ~x314 & ~x330 & ~x332 & ~x343 & ~x360 & ~x362 & ~x363 & ~x367 & ~x368 & ~x369 & ~x370 & ~x371 & ~x389 & ~x395 & ~x397 & ~x398 & ~x399 & ~x400 & ~x415 & ~x420 & ~x422 & ~x424 & ~x426 & ~x428 & ~x429 & ~x430 & ~x431 & ~x432 & ~x445 & ~x456 & ~x457 & ~x458 & ~x459 & ~x460 & ~x472 & ~x477 & ~x503 & ~x529 & ~x530 & ~x534 & ~x557 & ~x587 & ~x589 & ~x613 & ~x638 & ~x639 & ~x641 & ~x646 & ~x648 & ~x665 & ~x675 & ~x676 & ~x688 & ~x689 & ~x692 & ~x693 & ~x695 & ~x696 & ~x697 & ~x699 & ~x700 & ~x702 & ~x704 & ~x706 & ~x710 & ~x712 & ~x713 & ~x714 & ~x715 & ~x716 & ~x718 & ~x724 & ~x727 & ~x730 & ~x731 & ~x735 & ~x737 & ~x738 & ~x739 & ~x744 & ~x747 & ~x748 & ~x755 & ~x759 & ~x760 & ~x765 & ~x768 & ~x770 & ~x771 & ~x773 & ~x775 & ~x780 & ~x782 & ~x783;
assign c011 = ~x2 & ~x5 & ~x7 & ~x8 & ~x12 & ~x13 & ~x15 & ~x16 & ~x19 & ~x20 & ~x21 & ~x24 & ~x25 & ~x26 & ~x37 & ~x38 & ~x40 & ~x41 & ~x44 & ~x46 & ~x48 & ~x53 & ~x55 & ~x58 & ~x59 & ~x62 & ~x65 & ~x68 & ~x70 & ~x71 & ~x73 & ~x77 & ~x78 & ~x79 & ~x83 & ~x85 & ~x89 & ~x97 & ~x98 & ~x99 & ~x102 & ~x105 & ~x114 & ~x116 & ~x139 & ~x144 & ~x163 & ~x164 & ~x170 & ~x171 & ~x190 & ~x196 & ~x197 & ~x222 & ~x223 & ~x224 & ~x225 & ~x252 & ~x254 & ~x280 & ~x307 & ~x308 & ~x309 & ~x310 & ~x334 & ~x338 & ~x360 & ~x362 & ~x363 & ~x366 & ~x367 & ~x389 & ~x394 & ~x396 & ~x423 & ~x424 & ~x445 & ~x446 & ~x449 & ~x450 & ~x451 & ~x452 & ~x476 & ~x477 & ~x479 & ~x480 & ~x483 & ~x484 & ~x485 & ~x486 & ~x487 & ~x502 & ~x503 & ~x508 & ~x509 & ~x510 & ~x529 & ~x558 & ~x561 & ~x562 & ~x584 & ~x586 & ~x588 & ~x590 & ~x591 & ~x617 & ~x618 & ~x619 & ~x641 & ~x642 & ~x643 & ~x665 & ~x675 & ~x676 & ~x687 & ~x688 & ~x689 & ~x693 & ~x696 & ~x698 & ~x700 & ~x701 & ~x705 & ~x724 & ~x725 & ~x726 & ~x728 & ~x729 & ~x731 & ~x739 & ~x741 & ~x743 & ~x747 & ~x749 & ~x750 & ~x751 & ~x752 & ~x753 & ~x754 & ~x756 & ~x759 & ~x762 & ~x763 & ~x764 & ~x765 & ~x766 & ~x768 & ~x769 & ~x771 & ~x772 & ~x775 & ~x776 & ~x779 & ~x783;
assign c013 =  x460 & ~x47 & ~x63 & ~x319 & ~x345 & ~x707;
assign c015 =  x408 &  x409 & ~x297 & ~x298;
assign c017 = ~x16 & ~x55 & ~x73 & ~x84 & ~x193 & ~x304 & ~x316 & ~x331 & ~x346 & ~x372 & ~x421 & ~x443 & ~x558 & ~x632 & ~x652 & ~x655 & ~x656 & ~x682 & ~x697 & ~x704;
assign c019 = ~x48 & ~x74 & ~x76 & ~x178 & ~x206 & ~x207 & ~x233 & ~x254 & ~x278 & ~x281 & ~x335 & ~x385 & ~x388 & ~x409 & ~x410 & ~x413 & ~x414 & ~x437 & ~x473 & ~x525 & ~x719 & ~x761 & ~x762 & ~x778 & ~x782;
assign c021 =  x434 & ~x30 & ~x542;
assign c023 = ~x25 & ~x36 & ~x49 & ~x139 & ~x154 & ~x156 & ~x333 & ~x360 & ~x388 & ~x499 & ~x500 & ~x515 & ~x542 & ~x567 & ~x569 & ~x593 & ~x594 & ~x616 & ~x623 & ~x750;
assign c025 =  x349 &  x350 &  x351 & ~x9 & ~x29 & ~x45 & ~x116 & ~x194 & ~x225 & ~x250 & ~x273 & ~x300 & ~x422 & ~x424 & ~x464 & ~x536 & ~x593 & ~x620 & ~x678 & ~x767 & ~x780;
assign c027 =  x351 &  x377 & ~x13 & ~x24 & ~x34 & ~x172 & ~x196 & ~x226 & ~x284 & ~x304 & ~x329 & ~x331 & ~x359 & ~x480 & ~x544 & ~x546 & ~x699 & ~x709 & ~x757;
assign c029 = ~x10 & ~x15 & ~x22 & ~x55 & ~x58 & ~x59 & ~x60 & ~x63 & ~x66 & ~x80 & ~x85 & ~x106 & ~x108 & ~x113 & ~x117 & ~x136 & ~x146 & ~x147 & ~x167 & ~x170 & ~x192 & ~x221 & ~x226 & ~x244 & ~x246 & ~x249 & ~x270 & ~x271 & ~x278 & ~x285 & ~x297 & ~x298 & ~x299 & ~x301 & ~x302 & ~x303 & ~x311 & ~x331 & ~x332 & ~x366 & ~x367 & ~x394 & ~x420 & ~x445 & ~x449 & ~x452 & ~x475 & ~x480 & ~x532 & ~x556 & ~x564 & ~x566 & ~x594 & ~x595 & ~x613 & ~x618 & ~x620 & ~x622 & ~x640 & ~x643 & ~x648 & ~x664 & ~x667 & ~x669 & ~x670 & ~x671 & ~x673 & ~x677 & ~x693 & ~x716 & ~x728 & ~x735 & ~x739 & ~x746 & ~x749 & ~x750 & ~x754 & ~x762 & ~x766 & ~x767 & ~x768 & ~x774;
assign c031 =  x432 &  x433 &  x434 &  x435 &  x436 & ~x1 & ~x2 & ~x3 & ~x8 & ~x9 & ~x18 & ~x20 & ~x22 & ~x27 & ~x28 & ~x29 & ~x30 & ~x31 & ~x33 & ~x35 & ~x37 & ~x38 & ~x39 & ~x41 & ~x42 & ~x43 & ~x44 & ~x48 & ~x49 & ~x50 & ~x52 & ~x53 & ~x54 & ~x56 & ~x58 & ~x63 & ~x67 & ~x70 & ~x71 & ~x73 & ~x76 & ~x79 & ~x80 & ~x84 & ~x85 & ~x87 & ~x93 & ~x105 & ~x108 & ~x113 & ~x120 & ~x134 & ~x138 & ~x144 & ~x165 & ~x169 & ~x170 & ~x197 & ~x198 & ~x200 & ~x201 & ~x251 & ~x252 & ~x253 & ~x256 & ~x279 & ~x280 & ~x282 & ~x308 & ~x333 & ~x335 & ~x338 & ~x340 & ~x361 & ~x364 & ~x365 & ~x367 & ~x391 & ~x395 & ~x396 & ~x419 & ~x420 & ~x421 & ~x422 & ~x423 & ~x448 & ~x451 & ~x473 & ~x474 & ~x502 & ~x505 & ~x529 & ~x531 & ~x532 & ~x534 & ~x558 & ~x560 & ~x563 & ~x585 & ~x587 & ~x614 & ~x616 & ~x617 & ~x620 & ~x643 & ~x644 & ~x649 & ~x664 & ~x666 & ~x668 & ~x669 & ~x670 & ~x671 & ~x675 & ~x676 & ~x689 & ~x692 & ~x693 & ~x696 & ~x701 & ~x705 & ~x718 & ~x722 & ~x723 & ~x727 & ~x728 & ~x730 & ~x731 & ~x734 & ~x738 & ~x743 & ~x745 & ~x748 & ~x749 & ~x753 & ~x759 & ~x763 & ~x765 & ~x767 & ~x770 & ~x771 & ~x773 & ~x774 & ~x781 & ~x782 & ~x783;
assign c033 =  x350 &  x378 &  x380 &  x406 & ~x274;
assign c035 =  x458 &  x459 &  x463 & ~x51 & ~x69 & ~x135 & ~x164 & ~x280 & ~x448 & ~x505 & ~x562 & ~x696 & ~x743 & ~x744 & ~x779;
assign c037 = ~x0 & ~x1 & ~x36 & ~x84 & ~x95 & ~x96 & ~x134 & ~x135 & ~x152 & ~x167 & ~x222 & ~x226 & ~x305 & ~x331 & ~x338 & ~x362 & ~x365 & ~x366 & ~x387 & ~x389 & ~x444 & ~x449 & ~x534 & ~x542 & ~x543 & ~x567 & ~x568 & ~x569 & ~x571 & ~x645 & ~x699 & ~x723 & ~x724 & ~x777;
assign c039 =  x242 &  x244 & ~x17 & ~x27 & ~x39 & ~x62 & ~x63 & ~x87 & ~x92 & ~x96 & ~x97 & ~x128 & ~x129 & ~x143 & ~x197 & ~x201 & ~x397 & ~x417 & ~x418 & ~x421 & ~x442 & ~x456 & ~x471 & ~x485 & ~x557 & ~x560 & ~x610 & ~x618 & ~x668 & ~x701 & ~x723 & ~x729 & ~x743 & ~x768;
assign c041 =  x460 & ~x78 & ~x167 & ~x324 & ~x631 & ~x739;
assign c043 = ~x5 & ~x6 & ~x10 & ~x27 & ~x51 & ~x70 & ~x79 & ~x140 & ~x200 & ~x224 & ~x240 & ~x241 & ~x242 & ~x243 & ~x282 & ~x417 & ~x536 & ~x539 & ~x560 & ~x561 & ~x618 & ~x677 & ~x686 & ~x702 & ~x759 & ~x770;
assign c045 =  x348 &  x350 & ~x44 & ~x199 & ~x240 & ~x268 & ~x312 & ~x420 & ~x492 & ~x529 & ~x561 & ~x644 & ~x669 & ~x674 & ~x720 & ~x724 & ~x740 & ~x744 & ~x767;
assign c047 = ~x4 & ~x9 & ~x10 & ~x15 & ~x18 & ~x30 & ~x31 & ~x32 & ~x37 & ~x41 & ~x44 & ~x53 & ~x64 & ~x139 & ~x171 & ~x190 & ~x195 & ~x198 & ~x224 & ~x246 & ~x247 & ~x248 & ~x249 & ~x254 & ~x259 & ~x271 & ~x272 & ~x273 & ~x298 & ~x303 & ~x304 & ~x325 & ~x331 & ~x332 & ~x389 & ~x416 & ~x417 & ~x420 & ~x421 & ~x452 & ~x480 & ~x508 & ~x560 & ~x588 & ~x619 & ~x640 & ~x643 & ~x652 & ~x670 & ~x672 & ~x674 & ~x694 & ~x695 & ~x713 & ~x741 & ~x747 & ~x759 & ~x760 & ~x763 & ~x769 & ~x780;
assign c049 =  x435 &  x461 &  x464 & ~x14 & ~x22 & ~x34 & ~x43 & ~x108 & ~x136 & ~x311 & ~x323 & ~x351 & ~x614 & ~x640 & ~x773;
assign c051 =  x349 & ~x9 & ~x10 & ~x18 & ~x26 & ~x28 & ~x52 & ~x56 & ~x79 & ~x94 & ~x172 & ~x192 & ~x252 & ~x254 & ~x358 & ~x417 & ~x445 & ~x485 & ~x486 & ~x487 & ~x505 & ~x558 & ~x617 & ~x645 & ~x697 & ~x717 & ~x755;
assign c053 = ~x1 & ~x2 & ~x10 & ~x13 & ~x14 & ~x20 & ~x21 & ~x32 & ~x36 & ~x44 & ~x48 & ~x66 & ~x77 & ~x86 & ~x100 & ~x101 & ~x140 & ~x166 & ~x167 & ~x172 & ~x195 & ~x196 & ~x234 & ~x254 & ~x281 & ~x283 & ~x307 & ~x308 & ~x311 & ~x329 & ~x330 & ~x335 & ~x336 & ~x340 & ~x349 & ~x357 & ~x359 & ~x364 & ~x370 & ~x386 & ~x415 & ~x418 & ~x441 & ~x471 & ~x473 & ~x506 & ~x558 & ~x561 & ~x587 & ~x591 & ~x614 & ~x616 & ~x618 & ~x619 & ~x620 & ~x646 & ~x667 & ~x670 & ~x682 & ~x683 & ~x699 & ~x722 & ~x725 & ~x754 & ~x760 & ~x762 & ~x763 & ~x767 & ~x768 & ~x776 & ~x777 & ~x779 & ~x781 & ~x782;
assign c055 =  x439 &  x495 & ~x319 & ~x401 & ~x629 & ~x656 & ~x765;
assign c057 = ~x0 & ~x1 & ~x4 & ~x10 & ~x14 & ~x20 & ~x23 & ~x24 & ~x30 & ~x31 & ~x36 & ~x39 & ~x40 & ~x49 & ~x50 & ~x62 & ~x63 & ~x66 & ~x71 & ~x73 & ~x76 & ~x79 & ~x82 & ~x83 & ~x85 & ~x88 & ~x97 & ~x109 & ~x113 & ~x116 & ~x117 & ~x119 & ~x120 & ~x121 & ~x141 & ~x143 & ~x145 & ~x146 & ~x195 & ~x198 & ~x199 & ~x200 & ~x202 & ~x204 & ~x221 & ~x226 & ~x253 & ~x255 & ~x258 & ~x272 & ~x273 & ~x275 & ~x283 & ~x284 & ~x285 & ~x298 & ~x299 & ~x300 & ~x301 & ~x303 & ~x310 & ~x327 & ~x328 & ~x329 & ~x335 & ~x336 & ~x359 & ~x362 & ~x368 & ~x385 & ~x386 & ~x387 & ~x390 & ~x395 & ~x396 & ~x397 & ~x416 & ~x417 & ~x425 & ~x447 & ~x478 & ~x480 & ~x508 & ~x529 & ~x532 & ~x565 & ~x589 & ~x591 & ~x612 & ~x614 & ~x617 & ~x618 & ~x643 & ~x644 & ~x648 & ~x650 & ~x669 & ~x679 & ~x681 & ~x687 & ~x690 & ~x692 & ~x694 & ~x695 & ~x697 & ~x698 & ~x700 & ~x701 & ~x704 & ~x705 & ~x707 & ~x721 & ~x723 & ~x726 & ~x731 & ~x733 & ~x735 & ~x739 & ~x747 & ~x752 & ~x753 & ~x759 & ~x771 & ~x772 & ~x775 & ~x776;
assign c059 =  x350 &  x351 &  x352 & ~x4 & ~x21 & ~x23 & ~x28 & ~x31 & ~x35 & ~x36 & ~x38 & ~x47 & ~x55 & ~x56 & ~x61 & ~x79 & ~x80 & ~x106 & ~x109 & ~x111 & ~x140 & ~x195 & ~x197 & ~x225 & ~x226 & ~x249 & ~x253 & ~x263 & ~x305 & ~x331 & ~x336 & ~x339 & ~x358 & ~x362 & ~x363 & ~x387 & ~x392 & ~x423 & ~x461 & ~x463 & ~x530 & ~x561 & ~x587 & ~x588 & ~x614 & ~x644 & ~x645 & ~x647 & ~x648 & ~x667 & ~x669 & ~x671 & ~x673 & ~x675 & ~x677 & ~x679 & ~x691 & ~x696 & ~x698 & ~x710 & ~x723 & ~x725 & ~x726 & ~x732 & ~x743 & ~x754 & ~x755 & ~x757 & ~x765 & ~x768 & ~x773 & ~x774 & ~x780 & ~x781;
assign c061 =  x234 &  x463 &  x464 &  x465 & ~x26 & ~x35 & ~x39 & ~x40 & ~x45 & ~x51 & ~x53 & ~x57 & ~x58 & ~x59 & ~x61 & ~x63 & ~x66 & ~x91 & ~x95 & ~x116 & ~x117 & ~x118 & ~x141 & ~x143 & ~x145 & ~x147 & ~x165 & ~x167 & ~x169 & ~x172 & ~x173 & ~x196 & ~x198 & ~x221 & ~x222 & ~x252 & ~x277 & ~x278 & ~x306 & ~x311 & ~x337 & ~x338 & ~x362 & ~x365 & ~x391 & ~x421 & ~x422 & ~x450 & ~x474 & ~x476 & ~x506 & ~x530 & ~x564 & ~x589 & ~x619 & ~x647 & ~x667 & ~x695 & ~x698 & ~x700 & ~x704 & ~x733 & ~x743 & ~x752 & ~x763 & ~x770 & ~x772 & ~x775 & ~x777 & ~x779 & ~x783;
assign c063 =  x432 &  x461 &  x462 & ~x71 & ~x103 & ~x365 & ~x589 & ~x612 & ~x739 & ~x740 & ~x780;
assign c065 =  x328 & ~x10 & ~x18 & ~x25 & ~x43 & ~x47 & ~x82 & ~x101 & ~x102 & ~x108 & ~x110 & ~x114 & ~x145 & ~x163 & ~x223 & ~x225 & ~x337 & ~x390 & ~x419 & ~x445 & ~x454 & ~x507 & ~x513 & ~x539 & ~x556 & ~x721 & ~x749 & ~x765;
assign c067 = ~x2 & ~x5 & ~x8 & ~x9 & ~x21 & ~x22 & ~x27 & ~x31 & ~x33 & ~x37 & ~x42 & ~x43 & ~x46 & ~x48 & ~x50 & ~x55 & ~x62 & ~x64 & ~x65 & ~x69 & ~x70 & ~x74 & ~x75 & ~x78 & ~x79 & ~x81 & ~x84 & ~x85 & ~x89 & ~x90 & ~x92 & ~x97 & ~x98 & ~x101 & ~x103 & ~x106 & ~x111 & ~x119 & ~x135 & ~x140 & ~x142 & ~x145 & ~x147 & ~x162 & ~x166 & ~x197 & ~x198 & ~x199 & ~x227 & ~x252 & ~x253 & ~x279 & ~x284 & ~x308 & ~x338 & ~x339 & ~x360 & ~x361 & ~x363 & ~x364 & ~x393 & ~x395 & ~x417 & ~x419 & ~x421 & ~x422 & ~x423 & ~x424 & ~x425 & ~x452 & ~x453 & ~x454 & ~x455 & ~x475 & ~x476 & ~x478 & ~x480 & ~x484 & ~x485 & ~x486 & ~x500 & ~x502 & ~x503 & ~x515 & ~x516 & ~x533 & ~x559 & ~x615 & ~x639 & ~x640 & ~x642 & ~x645 & ~x646 & ~x668 & ~x675 & ~x678 & ~x701 & ~x704 & ~x705 & ~x706 & ~x722 & ~x726 & ~x729 & ~x730 & ~x732 & ~x733 & ~x736 & ~x741 & ~x744 & ~x752 & ~x754 & ~x757 & ~x760 & ~x765 & ~x766 & ~x767 & ~x768;
assign c069 =  x717;
assign c071 =  x263 & ~x8 & ~x11 & ~x75 & ~x127 & ~x153 & ~x154 & ~x196 & ~x352 & ~x353 & ~x377 & ~x387 & ~x475 & ~x508 & ~x526 & ~x528 & ~x537 & ~x539 & ~x554 & ~x699;
assign c073 = ~x1 & ~x5 & ~x7 & ~x12 & ~x13 & ~x15 & ~x21 & ~x23 & ~x27 & ~x28 & ~x31 & ~x39 & ~x40 & ~x41 & ~x44 & ~x49 & ~x52 & ~x53 & ~x60 & ~x63 & ~x65 & ~x67 & ~x68 & ~x69 & ~x70 & ~x71 & ~x73 & ~x77 & ~x78 & ~x88 & ~x97 & ~x102 & ~x103 & ~x105 & ~x108 & ~x116 & ~x117 & ~x119 & ~x134 & ~x136 & ~x138 & ~x139 & ~x141 & ~x144 & ~x193 & ~x194 & ~x198 & ~x199 & ~x220 & ~x222 & ~x225 & ~x254 & ~x280 & ~x281 & ~x307 & ~x309 & ~x337 & ~x361 & ~x363 & ~x365 & ~x388 & ~x391 & ~x393 & ~x395 & ~x416 & ~x421 & ~x422 & ~x425 & ~x426 & ~x427 & ~x429 & ~x430 & ~x431 & ~x433 & ~x445 & ~x448 & ~x450 & ~x453 & ~x456 & ~x458 & ~x460 & ~x476 & ~x478 & ~x480 & ~x481 & ~x482 & ~x483 & ~x484 & ~x500 & ~x501 & ~x502 & ~x508 & ~x532 & ~x559 & ~x561 & ~x584 & ~x587 & ~x589 & ~x590 & ~x614 & ~x642 & ~x643 & ~x644 & ~x665 & ~x667 & ~x671 & ~x672 & ~x673 & ~x674 & ~x676 & ~x692 & ~x696 & ~x697 & ~x701 & ~x702 & ~x703 & ~x704 & ~x715 & ~x720 & ~x727 & ~x735 & ~x738 & ~x743 & ~x745 & ~x748 & ~x750 & ~x755 & ~x756 & ~x759 & ~x762 & ~x764 & ~x768 & ~x775 & ~x776 & ~x779 & ~x783;
assign c075 =  x693;
assign c077 =  x434 & ~x8 & ~x168 & ~x480 & ~x593 & ~x657 & ~x706;
assign c079 =  x437 &  x466 & ~x2 & ~x4 & ~x27 & ~x40 & ~x50 & ~x84 & ~x142 & ~x194 & ~x267 & ~x334 & ~x363 & ~x421 & ~x448 & ~x503 & ~x506 & ~x534 & ~x559 & ~x587 & ~x595 & ~x613 & ~x638 & ~x648 & ~x720 & ~x725;
assign c081 =  x521 & ~x10 & ~x17 & ~x18 & ~x22 & ~x26 & ~x36 & ~x43 & ~x47 & ~x61 & ~x69 & ~x83 & ~x84 & ~x100 & ~x104 & ~x131 & ~x137 & ~x140 & ~x143 & ~x196 & ~x225 & ~x249 & ~x253 & ~x254 & ~x283 & ~x305 & ~x306 & ~x335 & ~x359 & ~x414 & ~x446 & ~x448 & ~x476 & ~x503 & ~x528 & ~x557 & ~x591 & ~x600 & ~x614 & ~x628 & ~x641 & ~x650 & ~x651 & ~x669 & ~x676 & ~x683 & ~x707 & ~x721 & ~x725 & ~x726 & ~x751 & ~x761 & ~x774 & ~x778;
assign c083 =  x363;
assign c085 =  x662 & ~x39 & ~x275 & ~x331 & ~x332 & ~x358 & ~x385 & ~x472 & ~x506 & ~x680 & ~x738;
assign c087 = ~x1 & ~x7 & ~x8 & ~x35 & ~x43 & ~x76 & ~x96 & ~x101 & ~x107 & ~x122 & ~x137 & ~x144 & ~x166 & ~x338 & ~x388 & ~x390 & ~x404 & ~x416 & ~x446 & ~x474 & ~x499 & ~x503 & ~x512 & ~x513 & ~x530 & ~x536 & ~x537 & ~x539 & ~x542 & ~x564 & ~x567 & ~x568 & ~x587 & ~x593 & ~x596 & ~x623 & ~x694 & ~x696 & ~x701 & ~x705 & ~x753 & ~x754 & ~x757 & ~x773;
assign c089 =  x463 & ~x4 & ~x92 & ~x272 & ~x306 & ~x308 & ~x312 & ~x322 & ~x450 & ~x536 & ~x615 & ~x616 & ~x651 & ~x730;
assign c091 =  x380 &  x404 &  x405 &  x406 &  x407 &  x431 & ~x31 & ~x123 & ~x224 & ~x278 & ~x337 & ~x393 & ~x448 & ~x591 & ~x761;
assign c093 = ~x28 & ~x45 & ~x85 & ~x228 & ~x272 & ~x273 & ~x298 & ~x299 & ~x300 & ~x302 & ~x305 & ~x332 & ~x360 & ~x369 & ~x373 & ~x395 & ~x503 & ~x587 & ~x612 & ~x684 & ~x723 & ~x733 & ~x768 & ~x772;
assign c095 =  x379 & ~x519;
assign c097 = ~x1 & ~x8 & ~x9 & ~x17 & ~x18 & ~x19 & ~x23 & ~x25 & ~x41 & ~x42 & ~x44 & ~x45 & ~x46 & ~x47 & ~x48 & ~x52 & ~x55 & ~x57 & ~x59 & ~x61 & ~x69 & ~x79 & ~x84 & ~x85 & ~x86 & ~x87 & ~x88 & ~x94 & ~x96 & ~x97 & ~x98 & ~x106 & ~x110 & ~x123 & ~x124 & ~x139 & ~x141 & ~x142 & ~x143 & ~x145 & ~x146 & ~x147 & ~x152 & ~x169 & ~x172 & ~x175 & ~x196 & ~x200 & ~x223 & ~x226 & ~x228 & ~x229 & ~x231 & ~x253 & ~x256 & ~x257 & ~x278 & ~x282 & ~x283 & ~x285 & ~x307 & ~x315 & ~x334 & ~x335 & ~x336 & ~x353 & ~x354 & ~x355 & ~x356 & ~x357 & ~x358 & ~x359 & ~x362 & ~x366 & ~x370 & ~x386 & ~x387 & ~x390 & ~x398 & ~x412 & ~x413 & ~x416 & ~x420 & ~x422 & ~x423 & ~x424 & ~x442 & ~x447 & ~x448 & ~x450 & ~x472 & ~x474 & ~x502 & ~x528 & ~x529 & ~x530 & ~x531 & ~x532 & ~x557 & ~x558 & ~x560 & ~x585 & ~x593 & ~x615 & ~x616 & ~x618 & ~x619 & ~x637 & ~x639 & ~x644 & ~x645 & ~x668 & ~x669 & ~x670 & ~x676 & ~x677 & ~x678 & ~x697 & ~x698 & ~x702 & ~x705 & ~x708 & ~x720 & ~x722 & ~x728 & ~x731 & ~x732 & ~x733 & ~x738 & ~x739 & ~x743 & ~x748 & ~x756 & ~x758 & ~x763 & ~x771 & ~x772 & ~x781 & ~x783;
assign c099 =  x518 & ~x23 & ~x51 & ~x86 & ~x136 & ~x164 & ~x266 & ~x268 & ~x321 & ~x338 & ~x370 & ~x371 & ~x389 & ~x446 & ~x477 & ~x557 & ~x560 & ~x591 & ~x618 & ~x672 & ~x727 & ~x747 & ~x757;
assign c0101 = ~x4 & ~x30 & ~x33 & ~x35 & ~x39 & ~x40 & ~x67 & ~x68 & ~x88 & ~x108 & ~x199 & ~x242 & ~x245 & ~x248 & ~x249 & ~x268 & ~x269 & ~x272 & ~x273 & ~x299 & ~x300 & ~x301 & ~x303 & ~x305 & ~x339 & ~x360 & ~x363 & ~x418 & ~x424 & ~x451 & ~x503 & ~x506 & ~x561 & ~x586 & ~x650 & ~x671 & ~x691 & ~x692 & ~x710 & ~x723 & ~x730 & ~x757 & ~x760 & ~x772 & ~x774;
assign c0103 = ~x2 & ~x6 & ~x26 & ~x53 & ~x57 & ~x81 & ~x82 & ~x106 & ~x112 & ~x114 & ~x133 & ~x144 & ~x186 & ~x196 & ~x229 & ~x279 & ~x285 & ~x309 & ~x335 & ~x341 & ~x368 & ~x369 & ~x417 & ~x453 & ~x467 & ~x472 & ~x474 & ~x478 & ~x505 & ~x526 & ~x530 & ~x531 & ~x532 & ~x554 & ~x559 & ~x561 & ~x614 & ~x675 & ~x695 & ~x700 & ~x713 & ~x727 & ~x731 & ~x733 & ~x739 & ~x744 & ~x746 & ~x765 & ~x772 & ~x779;
assign c0105 =  x407 & ~x39 & ~x44 & ~x338 & ~x632 & ~x633 & ~x648 & ~x651 & ~x653 & ~x655 & ~x674 & ~x758;
assign c0107 =  x348 &  x349 &  x351 & ~x32 & ~x57 & ~x75 & ~x88 & ~x93 & ~x304 & ~x305 & ~x335 & ~x338 & ~x359 & ~x361 & ~x388 & ~x394 & ~x459 & ~x504 & ~x512 & ~x589 & ~x615 & ~x616 & ~x670 & ~x694 & ~x706 & ~x725 & ~x728 & ~x755 & ~x759 & ~x770;
assign c0109 =  x711;
assign c0111 = ~x4 & ~x209 & ~x216 & ~x239 & ~x285 & ~x367 & ~x397 & ~x686;
assign c0113 =  x460 &  x461 & ~x45 & ~x61 & ~x75 & ~x221 & ~x295 & ~x339 & ~x343 & ~x645 & ~x669 & ~x698 & ~x748;
assign c0115 = ~x35 & ~x36 & ~x46 & ~x87 & ~x106 & ~x109 & ~x145 & ~x170 & ~x224 & ~x250 & ~x255 & ~x268 & ~x337 & ~x341 & ~x344 & ~x345 & ~x347 & ~x361 & ~x369 & ~x389 & ~x393 & ~x414 & ~x441 & ~x447 & ~x588 & ~x646 & ~x649 & ~x665 & ~x692 & ~x699 & ~x707 & ~x718 & ~x730 & ~x745 & ~x749 & ~x750 & ~x759;
assign c0117 =  x102 & ~x301;
assign c0119 =  x379 & ~x1 & ~x8 & ~x57 & ~x70 & ~x110 & ~x123 & ~x229 & ~x267 & ~x361 & ~x446 & ~x453 & ~x506 & ~x698 & ~x700 & ~x741;
assign c0121 =  x535;
assign c0123 = ~x1 & ~x52 & ~x92 & ~x165 & ~x167 & ~x251 & ~x254 & ~x366 & ~x392 & ~x419 & ~x422 & ~x425 & ~x426 & ~x427 & ~x484 & ~x493 & ~x508 & ~x509 & ~x523 & ~x525 & ~x526 & ~x551 & ~x554 & ~x560 & ~x638 & ~x701 & ~x724 & ~x776;
assign c0125 = ~x22 & ~x26 & ~x91 & ~x118 & ~x168 & ~x170 & ~x187 & ~x192 & ~x215 & ~x222 & ~x240 & ~x313 & ~x425 & ~x451 & ~x452 & ~x530 & ~x533 & ~x559 & ~x561 & ~x611 & ~x613 & ~x619 & ~x667 & ~x673 & ~x678 & ~x711 & ~x722 & ~x725 & ~x727 & ~x751 & ~x777;
assign c0127 =  x406 & ~x324 & ~x770;
assign c0129 = ~x0 & ~x9 & ~x10 & ~x38 & ~x69 & ~x70 & ~x95 & ~x178 & ~x196 & ~x197 & ~x225 & ~x229 & ~x279 & ~x331 & ~x336 & ~x359 & ~x389 & ~x500 & ~x525 & ~x526 & ~x552 & ~x554 & ~x564 & ~x571 & ~x585 & ~x590 & ~x593 & ~x597 & ~x622 & ~x651 & ~x672 & ~x677 & ~x734 & ~x754 & ~x769;
assign c0131 = ~x2 & ~x3 & ~x4 & ~x5 & ~x6 & ~x7 & ~x9 & ~x11 & ~x12 & ~x14 & ~x17 & ~x19 & ~x20 & ~x21 & ~x24 & ~x25 & ~x35 & ~x44 & ~x45 & ~x46 & ~x50 & ~x60 & ~x61 & ~x65 & ~x70 & ~x73 & ~x79 & ~x80 & ~x85 & ~x90 & ~x91 & ~x97 & ~x99 & ~x104 & ~x112 & ~x118 & ~x120 & ~x138 & ~x139 & ~x140 & ~x144 & ~x145 & ~x149 & ~x150 & ~x164 & ~x168 & ~x169 & ~x173 & ~x197 & ~x198 & ~x228 & ~x250 & ~x252 & ~x253 & ~x254 & ~x281 & ~x283 & ~x305 & ~x309 & ~x332 & ~x362 & ~x366 & ~x367 & ~x388 & ~x390 & ~x417 & ~x444 & ~x445 & ~x448 & ~x472 & ~x477 & ~x479 & ~x500 & ~x502 & ~x506 & ~x509 & ~x528 & ~x530 & ~x531 & ~x537 & ~x539 & ~x540 & ~x541 & ~x542 & ~x556 & ~x586 & ~x609 & ~x613 & ~x614 & ~x615 & ~x636 & ~x640 & ~x668 & ~x672 & ~x673 & ~x675 & ~x676 & ~x689 & ~x701 & ~x716 & ~x717 & ~x725 & ~x726 & ~x730 & ~x738 & ~x748 & ~x754 & ~x770 & ~x772 & ~x781 & ~x782;
assign c0133 = ~x0 & ~x2 & ~x3 & ~x12 & ~x13 & ~x14 & ~x15 & ~x16 & ~x20 & ~x21 & ~x22 & ~x25 & ~x26 & ~x28 & ~x29 & ~x32 & ~x33 & ~x34 & ~x35 & ~x38 & ~x39 & ~x41 & ~x42 & ~x43 & ~x44 & ~x45 & ~x46 & ~x47 & ~x49 & ~x51 & ~x53 & ~x57 & ~x58 & ~x61 & ~x64 & ~x66 & ~x67 & ~x70 & ~x71 & ~x73 & ~x75 & ~x77 & ~x80 & ~x83 & ~x84 & ~x86 & ~x87 & ~x88 & ~x89 & ~x101 & ~x107 & ~x110 & ~x111 & ~x113 & ~x114 & ~x115 & ~x118 & ~x119 & ~x120 & ~x133 & ~x134 & ~x135 & ~x136 & ~x137 & ~x138 & ~x139 & ~x141 & ~x143 & ~x145 & ~x168 & ~x169 & ~x170 & ~x171 & ~x172 & ~x174 & ~x193 & ~x195 & ~x196 & ~x197 & ~x198 & ~x200 & ~x202 & ~x220 & ~x223 & ~x224 & ~x226 & ~x227 & ~x248 & ~x249 & ~x251 & ~x253 & ~x254 & ~x277 & ~x280 & ~x282 & ~x305 & ~x307 & ~x332 & ~x333 & ~x334 & ~x336 & ~x338 & ~x339 & ~x360 & ~x361 & ~x363 & ~x367 & ~x388 & ~x392 & ~x393 & ~x395 & ~x396 & ~x415 & ~x416 & ~x417 & ~x418 & ~x419 & ~x420 & ~x421 & ~x424 & ~x425 & ~x430 & ~x432 & ~x443 & ~x446 & ~x448 & ~x450 & ~x455 & ~x456 & ~x457 & ~x458 & ~x459 & ~x474 & ~x476 & ~x479 & ~x501 & ~x502 & ~x504 & ~x529 & ~x530 & ~x531 & ~x532 & ~x533 & ~x535 & ~x557 & ~x559 & ~x560 & ~x562 & ~x585 & ~x591 & ~x611 & ~x613 & ~x615 & ~x617 & ~x619 & ~x639 & ~x640 & ~x642 & ~x644 & ~x645 & ~x647 & ~x665 & ~x668 & ~x670 & ~x671 & ~x672 & ~x673 & ~x674 & ~x675 & ~x693 & ~x694 & ~x695 & ~x696 & ~x698 & ~x699 & ~x700 & ~x703 & ~x708 & ~x709 & ~x713 & ~x714 & ~x715 & ~x717 & ~x718 & ~x719 & ~x720 & ~x721 & ~x725 & ~x726 & ~x727 & ~x728 & ~x729 & ~x731 & ~x733 & ~x736 & ~x737 & ~x741 & ~x743 & ~x745 & ~x746 & ~x747 & ~x749 & ~x750 & ~x751 & ~x755 & ~x758 & ~x759 & ~x761 & ~x763 & ~x764 & ~x765 & ~x767 & ~x768 & ~x771 & ~x772 & ~x773 & ~x774 & ~x775 & ~x778 & ~x780;
assign c0135 = ~x6 & ~x14 & ~x24 & ~x25 & ~x29 & ~x34 & ~x36 & ~x38 & ~x44 & ~x57 & ~x58 & ~x65 & ~x68 & ~x73 & ~x75 & ~x83 & ~x87 & ~x97 & ~x103 & ~x112 & ~x137 & ~x141 & ~x143 & ~x166 & ~x172 & ~x195 & ~x197 & ~x222 & ~x223 & ~x229 & ~x280 & ~x282 & ~x284 & ~x305 & ~x358 & ~x362 & ~x365 & ~x366 & ~x387 & ~x388 & ~x390 & ~x414 & ~x418 & ~x419 & ~x420 & ~x443 & ~x450 & ~x455 & ~x471 & ~x478 & ~x479 & ~x485 & ~x486 & ~x488 & ~x500 & ~x501 & ~x503 & ~x513 & ~x514 & ~x515 & ~x516 & ~x527 & ~x529 & ~x531 & ~x558 & ~x560 & ~x585 & ~x587 & ~x590 & ~x642 & ~x665 & ~x675 & ~x692 & ~x703 & ~x704 & ~x722 & ~x726 & ~x744 & ~x750 & ~x754 & ~x770 & ~x782 & ~x783;
assign c0137 =  x549 & ~x227 & ~x328 & ~x330 & ~x369 & ~x382 & ~x422 & ~x565;
assign c0139 = ~x109 & ~x185 & ~x357 & ~x453 & ~x481 & ~x514;
assign c0141 = ~x2 & ~x7 & ~x10 & ~x12 & ~x13 & ~x16 & ~x18 & ~x20 & ~x39 & ~x41 & ~x44 & ~x46 & ~x47 & ~x50 & ~x53 & ~x59 & ~x64 & ~x67 & ~x71 & ~x85 & ~x86 & ~x87 & ~x92 & ~x107 & ~x116 & ~x139 & ~x166 & ~x169 & ~x172 & ~x198 & ~x199 & ~x243 & ~x244 & ~x245 & ~x250 & ~x270 & ~x271 & ~x278 & ~x283 & ~x285 & ~x297 & ~x302 & ~x306 & ~x312 & ~x330 & ~x332 & ~x334 & ~x336 & ~x361 & ~x365 & ~x367 & ~x368 & ~x369 & ~x388 & ~x392 & ~x394 & ~x398 & ~x421 & ~x449 & ~x474 & ~x475 & ~x478 & ~x534 & ~x557 & ~x586 & ~x590 & ~x593 & ~x611 & ~x614 & ~x621 & ~x639 & ~x646 & ~x647 & ~x667 & ~x668 & ~x673 & ~x675 & ~x678 & ~x679 & ~x681 & ~x689 & ~x693 & ~x698 & ~x699 & ~x700 & ~x709 & ~x711 & ~x714 & ~x721 & ~x723 & ~x736 & ~x741 & ~x743 & ~x745 & ~x749 & ~x751 & ~x756 & ~x769 & ~x770 & ~x778 & ~x781;
assign c0143 =  x249;
assign c0145 =  x350 &  x352 &  x603 & ~x0 & ~x2 & ~x16 & ~x23 & ~x30 & ~x40 & ~x41 & ~x43 & ~x49 & ~x66 & ~x73 & ~x75 & ~x78 & ~x90 & ~x104 & ~x169 & ~x170 & ~x172 & ~x174 & ~x197 & ~x201 & ~x225 & ~x226 & ~x229 & ~x255 & ~x275 & ~x278 & ~x311 & ~x363 & ~x364 & ~x365 & ~x367 & ~x394 & ~x396 & ~x418 & ~x419 & ~x445 & ~x488 & ~x502 & ~x516 & ~x558 & ~x586 & ~x591 & ~x610 & ~x642 & ~x643 & ~x646 & ~x670 & ~x673 & ~x697 & ~x709 & ~x710 & ~x718 & ~x720 & ~x723 & ~x725 & ~x737 & ~x739 & ~x747 & ~x755 & ~x763 & ~x768 & ~x776 & ~x777;
assign c0147 =  x511 &  x522 &  x550 & ~x6 & ~x79 & ~x196 & ~x341 & ~x356 & ~x389 & ~x413 & ~x414 & ~x502 & ~x531 & ~x618 & ~x681 & ~x777 & ~x780 & ~x782;
assign c0149 =  x379 &  x406 & ~x2 & ~x3 & ~x4 & ~x6 & ~x12 & ~x29 & ~x30 & ~x35 & ~x37 & ~x40 & ~x41 & ~x43 & ~x45 & ~x51 & ~x53 & ~x73 & ~x87 & ~x91 & ~x108 & ~x140 & ~x143 & ~x148 & ~x172 & ~x195 & ~x227 & ~x311 & ~x356 & ~x357 & ~x358 & ~x362 & ~x387 & ~x388 & ~x390 & ~x393 & ~x419 & ~x449 & ~x451 & ~x473 & ~x505 & ~x530 & ~x533 & ~x562 & ~x617 & ~x640 & ~x641 & ~x642 & ~x644 & ~x666 & ~x669 & ~x672 & ~x673 & ~x676 & ~x690 & ~x693 & ~x696 & ~x700 & ~x703 & ~x721 & ~x722 & ~x726 & ~x731 & ~x733 & ~x734 & ~x735 & ~x742 & ~x745 & ~x751 & ~x752 & ~x763 & ~x764 & ~x771 & ~x779 & ~x782;
assign c0151 = ~x43 & ~x54 & ~x61 & ~x62 & ~x86 & ~x107 & ~x110 & ~x116 & ~x146 & ~x165 & ~x172 & ~x187 & ~x215 & ~x220 & ~x241 & ~x242 & ~x249 & ~x268 & ~x282 & ~x359 & ~x448 & ~x478 & ~x564 & ~x584 & ~x587 & ~x592 & ~x621 & ~x622 & ~x639 & ~x683 & ~x684 & ~x687 & ~x713 & ~x717 & ~x725 & ~x735 & ~x739 & ~x741 & ~x761 & ~x773 & ~x780;
assign c0153 =  x406 &  x433 & ~x686 & ~x776 & ~x783;
assign c0155 =  x492 & ~x114 & ~x194 & ~x291 & ~x318 & ~x319 & ~x321 & ~x475 & ~x476 & ~x630 & ~x675 & ~x731;
assign c0157 =  x492 &  x520 & ~x359 & ~x387 & ~x571 & ~x572 & ~x573;
assign c0159 =  x324 & ~x453 & ~x454 & ~x455 & ~x458 & ~x483;
assign c0161 =  x464 & ~x2 & ~x9 & ~x16 & ~x19 & ~x22 & ~x32 & ~x36 & ~x37 & ~x38 & ~x43 & ~x44 & ~x51 & ~x52 & ~x59 & ~x64 & ~x75 & ~x80 & ~x90 & ~x167 & ~x198 & ~x224 & ~x253 & ~x292 & ~x294 & ~x337 & ~x389 & ~x393 & ~x423 & ~x424 & ~x447 & ~x452 & ~x475 & ~x532 & ~x562 & ~x585 & ~x676 & ~x680 & ~x691 & ~x702 & ~x721 & ~x722 & ~x723 & ~x734 & ~x749 & ~x750 & ~x751 & ~x778 & ~x783;
assign c0163 =  x520 & ~x13 & ~x35 & ~x60 & ~x67 & ~x80 & ~x82 & ~x83 & ~x114 & ~x138 & ~x198 & ~x228 & ~x248 & ~x254 & ~x277 & ~x284 & ~x308 & ~x314 & ~x319 & ~x321 & ~x333 & ~x369 & ~x529 & ~x533 & ~x535 & ~x558 & ~x620 & ~x657 & ~x668 & ~x685 & ~x688 & ~x731 & ~x736 & ~x759 & ~x760 & ~x763 & ~x764 & ~x769 & ~x777;
assign c0165 =  x404 &  x405 &  x406 & ~x29 & ~x32 & ~x56 & ~x86 & ~x98 & ~x138 & ~x141 & ~x197 & ~x279 & ~x307 & ~x357 & ~x358 & ~x368 & ~x393 & ~x395 & ~x444 & ~x480 & ~x563 & ~x610 & ~x619 & ~x642 & ~x666 & ~x668 & ~x675 & ~x701 & ~x712 & ~x715 & ~x738 & ~x753 & ~x772 & ~x775;
assign c0167 = ~x26 & ~x265 & ~x282 & ~x356 & ~x384 & ~x386 & ~x413 & ~x415 & ~x618 & ~x654 & ~x655 & ~x762;
assign c0169 = ~x5 & ~x182 & ~x190 & ~x514 & ~x526 & ~x529 & ~x542 & ~x567 & ~x593;
assign c0171 =  x436 & ~x242 & ~x269 & ~x475 & ~x618;
assign c0173 =  x327 & ~x240 & ~x242;
assign c0175 =  x406 & ~x10 & ~x12 & ~x20 & ~x31 & ~x52 & ~x86 & ~x113 & ~x170 & ~x171 & ~x199 & ~x422 & ~x423 & ~x449 & ~x468 & ~x480 & ~x494 & ~x495 & ~x537 & ~x589 & ~x618 & ~x761 & ~x777 & ~x783;
assign c0177 =  x465 & ~x154 & ~x155 & ~x156 & ~x415 & ~x498 & ~x569 & ~x593 & ~x594 & ~x595 & ~x596 & ~x622 & ~x624 & ~x633;
assign c0179 =  x409 & ~x213 & ~x268 & ~x297 & ~x322;
assign c0181 = ~x0 & ~x1 & ~x6 & ~x7 & ~x8 & ~x9 & ~x10 & ~x14 & ~x15 & ~x16 & ~x17 & ~x18 & ~x19 & ~x21 & ~x23 & ~x24 & ~x25 & ~x29 & ~x30 & ~x32 & ~x34 & ~x37 & ~x38 & ~x39 & ~x40 & ~x41 & ~x42 & ~x43 & ~x45 & ~x46 & ~x47 & ~x49 & ~x50 & ~x51 & ~x52 & ~x53 & ~x54 & ~x55 & ~x57 & ~x58 & ~x59 & ~x62 & ~x66 & ~x67 & ~x69 & ~x70 & ~x71 & ~x72 & ~x73 & ~x76 & ~x77 & ~x79 & ~x80 & ~x81 & ~x83 & ~x85 & ~x86 & ~x90 & ~x91 & ~x92 & ~x93 & ~x94 & ~x95 & ~x97 & ~x98 & ~x102 & ~x103 & ~x105 & ~x106 & ~x107 & ~x108 & ~x109 & ~x110 & ~x112 & ~x113 & ~x115 & ~x117 & ~x119 & ~x120 & ~x135 & ~x136 & ~x137 & ~x138 & ~x141 & ~x142 & ~x143 & ~x145 & ~x167 & ~x170 & ~x194 & ~x197 & ~x198 & ~x199 & ~x223 & ~x228 & ~x250 & ~x251 & ~x252 & ~x253 & ~x255 & ~x256 & ~x276 & ~x278 & ~x280 & ~x281 & ~x283 & ~x285 & ~x304 & ~x306 & ~x307 & ~x308 & ~x309 & ~x310 & ~x312 & ~x331 & ~x332 & ~x334 & ~x336 & ~x337 & ~x361 & ~x363 & ~x365 & ~x367 & ~x368 & ~x370 & ~x388 & ~x389 & ~x391 & ~x394 & ~x397 & ~x398 & ~x416 & ~x417 & ~x423 & ~x424 & ~x425 & ~x426 & ~x427 & ~x428 & ~x430 & ~x431 & ~x432 & ~x445 & ~x446 & ~x447 & ~x448 & ~x449 & ~x450 & ~x452 & ~x453 & ~x454 & ~x455 & ~x456 & ~x473 & ~x474 & ~x475 & ~x476 & ~x483 & ~x501 & ~x502 & ~x504 & ~x505 & ~x507 & ~x528 & ~x529 & ~x531 & ~x532 & ~x557 & ~x562 & ~x563 & ~x583 & ~x584 & ~x586 & ~x587 & ~x589 & ~x610 & ~x611 & ~x613 & ~x615 & ~x637 & ~x638 & ~x640 & ~x642 & ~x644 & ~x646 & ~x665 & ~x666 & ~x668 & ~x669 & ~x671 & ~x672 & ~x676 & ~x692 & ~x694 & ~x696 & ~x697 & ~x700 & ~x703 & ~x704 & ~x707 & ~x708 & ~x710 & ~x712 & ~x714 & ~x717 & ~x718 & ~x719 & ~x724 & ~x725 & ~x727 & ~x728 & ~x732 & ~x733 & ~x739 & ~x743 & ~x744 & ~x746 & ~x747 & ~x749 & ~x750 & ~x753 & ~x754 & ~x755 & ~x756 & ~x757 & ~x759 & ~x760 & ~x761 & ~x764 & ~x766 & ~x768 & ~x769 & ~x771 & ~x772 & ~x773 & ~x776 & ~x777 & ~x778 & ~x779 & ~x780 & ~x781 & ~x782;
assign c0183 =  x317 & ~x22 & ~x125 & ~x128 & ~x132 & ~x139 & ~x148 & ~x154 & ~x156 & ~x251 & ~x255 & ~x351 & ~x361 & ~x393 & ~x395 & ~x442 & ~x470 & ~x480 & ~x498 & ~x537 & ~x539 & ~x552 & ~x564 & ~x593 & ~x615 & ~x621 & ~x760 & ~x761;
assign c0185 =  x716;
assign c0187 =  x434 &  x435 &  x436 & ~x446;
assign c0189 = ~x12 & ~x13 & ~x30 & ~x34 & ~x61 & ~x66 & ~x86 & ~x108 & ~x111 & ~x141 & ~x171 & ~x204 & ~x242 & ~x244 & ~x269 & ~x286 & ~x341 & ~x359 & ~x360 & ~x369 & ~x386 & ~x387 & ~x445 & ~x557 & ~x561 & ~x562 & ~x565 & ~x585 & ~x594 & ~x624 & ~x707 & ~x710 & ~x717 & ~x742 & ~x773;
assign c0191 = ~x49 & ~x154 & ~x444 & ~x514 & ~x541 & ~x544 & ~x564 & ~x571 & ~x595 & ~x622 & ~x626;
assign c0193 =  x433;
assign c0195 =  x565 & ~x5 & ~x37 & ~x45 & ~x51 & ~x53 & ~x70 & ~x79 & ~x92 & ~x108 & ~x225 & ~x338 & ~x344 & ~x363 & ~x365 & ~x369 & ~x370 & ~x373 & ~x374 & ~x395 & ~x396 & ~x398 & ~x445 & ~x501 & ~x556 & ~x559 & ~x562 & ~x611 & ~x640 & ~x646 & ~x676 & ~x736 & ~x746 & ~x774 & ~x776 & ~x777 & ~x780 & ~x782;
assign c0197 =  x408 &  x513 & ~x8 & ~x18 & ~x27 & ~x37 & ~x44 & ~x63 & ~x86 & ~x89 & ~x91 & ~x109 & ~x113 & ~x125 & ~x128 & ~x130 & ~x131 & ~x140 & ~x145 & ~x199 & ~x221 & ~x226 & ~x249 & ~x252 & ~x306 & ~x336 & ~x362 & ~x363 & ~x390 & ~x420 & ~x446 & ~x531 & ~x585 & ~x590 & ~x614 & ~x643 & ~x697 & ~x721 & ~x723 & ~x729 & ~x753 & ~x763 & ~x777 & ~x783;
assign c0199 =  x462 & ~x35 & ~x87 & ~x137 & ~x229 & ~x287 & ~x343 & ~x351 & ~x400 & ~x425 & ~x453 & ~x473 & ~x640 & ~x701 & ~x721 & ~x726 & ~x751 & ~x757;
assign c0201 = ~x97 & ~x168 & ~x271 & ~x301 & ~x337 & ~x339 & ~x425 & ~x453 & ~x454 & ~x460 & ~x490 & ~x517 & ~x561 & ~x735 & ~x746 & ~x748 & ~x757 & ~x782;
assign c0203 =  x461 & ~x629 & ~x655;
assign c0205 =  x324 & ~x301 & ~x425 & ~x426 & ~x427 & ~x464 & ~x516 & ~x745;
assign c0207 = ~x24 & ~x41 & ~x54 & ~x81 & ~x130 & ~x150 & ~x176 & ~x200 & ~x311 & ~x354 & ~x365 & ~x411 & ~x413 & ~x443 & ~x474 & ~x478 & ~x498 & ~x523 & ~x560 & ~x620 & ~x639 & ~x644 & ~x666 & ~x694 & ~x695 & ~x701 & ~x717 & ~x725 & ~x730 & ~x767 & ~x771;
assign c0209 = ~x1 & ~x4 & ~x5 & ~x10 & ~x11 & ~x12 & ~x15 & ~x17 & ~x22 & ~x30 & ~x33 & ~x36 & ~x37 & ~x45 & ~x47 & ~x49 & ~x50 & ~x51 & ~x52 & ~x53 & ~x54 & ~x59 & ~x68 & ~x69 & ~x72 & ~x75 & ~x78 & ~x83 & ~x85 & ~x90 & ~x106 & ~x110 & ~x135 & ~x136 & ~x143 & ~x164 & ~x167 & ~x168 & ~x193 & ~x199 & ~x226 & ~x336 & ~x339 & ~x342 & ~x360 & ~x361 & ~x362 & ~x368 & ~x369 & ~x390 & ~x392 & ~x394 & ~x396 & ~x397 & ~x398 & ~x399 & ~x401 & ~x402 & ~x403 & ~x416 & ~x423 & ~x424 & ~x425 & ~x426 & ~x427 & ~x428 & ~x429 & ~x444 & ~x445 & ~x449 & ~x454 & ~x455 & ~x456 & ~x472 & ~x474 & ~x479 & ~x480 & ~x501 & ~x502 & ~x506 & ~x527 & ~x531 & ~x532 & ~x534 & ~x559 & ~x586 & ~x613 & ~x615 & ~x616 & ~x640 & ~x646 & ~x648 & ~x667 & ~x668 & ~x671 & ~x672 & ~x676 & ~x691 & ~x696 & ~x705 & ~x706 & ~x714 & ~x718 & ~x721 & ~x727 & ~x731 & ~x733 & ~x735 & ~x736 & ~x739 & ~x740 & ~x742 & ~x747 & ~x755 & ~x757 & ~x760 & ~x770 & ~x779 & ~x780 & ~x781;
assign c0211 = ~x37 & ~x83 & ~x215 & ~x239 & ~x240 & ~x242 & ~x266 & ~x336 & ~x446 & ~x621 & ~x655 & ~x656 & ~x657 & ~x659 & ~x662 & ~x683 & ~x734;
assign c0213 = ~x32 & ~x33 & ~x90 & ~x168 & ~x197 & ~x199 & ~x230 & ~x233 & ~x258 & ~x269 & ~x270 & ~x272 & ~x274 & ~x275 & ~x297 & ~x298 & ~x303 & ~x363 & ~x447 & ~x536 & ~x562 & ~x565 & ~x584 & ~x594 & ~x614 & ~x624 & ~x644 & ~x674 & ~x728 & ~x730 & ~x765 & ~x767;
assign c0215 =  x350 &  x378 &  x380 & ~x30 & ~x33 & ~x48 & ~x59 & ~x66 & ~x81 & ~x85 & ~x221 & ~x255 & ~x331 & ~x332 & ~x391 & ~x451 & ~x478 & ~x491 & ~x501 & ~x517 & ~x518 & ~x615 & ~x648 & ~x704 & ~x729 & ~x748 & ~x755;
assign c0217 =  x487 &  x489 & ~x6 & ~x9 & ~x14 & ~x23 & ~x37 & ~x49 & ~x51 & ~x59 & ~x61 & ~x69 & ~x76 & ~x78 & ~x107 & ~x111 & ~x113 & ~x115 & ~x137 & ~x145 & ~x169 & ~x170 & ~x222 & ~x281 & ~x359 & ~x362 & ~x377 & ~x386 & ~x387 & ~x393 & ~x403 & ~x422 & ~x423 & ~x424 & ~x445 & ~x446 & ~x451 & ~x473 & ~x561 & ~x642 & ~x696 & ~x716 & ~x717 & ~x737 & ~x738 & ~x740 & ~x742 & ~x753 & ~x760 & ~x761 & ~x766 & ~x772 & ~x777;
assign c0219 = ~x4 & ~x8 & ~x19 & ~x24 & ~x41 & ~x42 & ~x44 & ~x52 & ~x66 & ~x67 & ~x70 & ~x87 & ~x97 & ~x114 & ~x134 & ~x140 & ~x142 & ~x143 & ~x169 & ~x195 & ~x222 & ~x251 & ~x276 & ~x304 & ~x310 & ~x393 & ~x417 & ~x422 & ~x473 & ~x481 & ~x482 & ~x484 & ~x485 & ~x507 & ~x508 & ~x510 & ~x511 & ~x514 & ~x515 & ~x558 & ~x562 & ~x564 & ~x588 & ~x644 & ~x669 & ~x699 & ~x714 & ~x717 & ~x720 & ~x723 & ~x725 & ~x728 & ~x729 & ~x740 & ~x756 & ~x762 & ~x781;
assign c0221 = ~x6 & ~x10 & ~x28 & ~x33 & ~x35 & ~x38 & ~x51 & ~x53 & ~x77 & ~x79 & ~x110 & ~x117 & ~x120 & ~x134 & ~x138 & ~x142 & ~x169 & ~x193 & ~x194 & ~x219 & ~x336 & ~x359 & ~x419 & ~x499 & ~x507 & ~x561 & ~x563 & ~x570 & ~x572 & ~x592 & ~x595 & ~x596 & ~x597 & ~x599 & ~x621 & ~x626 & ~x677 & ~x679 & ~x697 & ~x699 & ~x703 & ~x705 & ~x708 & ~x723 & ~x726 & ~x759 & ~x760 & ~x767 & ~x777;
assign c0223 = ~x3 & ~x6 & ~x8 & ~x10 & ~x15 & ~x23 & ~x26 & ~x29 & ~x34 & ~x42 & ~x52 & ~x55 & ~x56 & ~x57 & ~x65 & ~x69 & ~x77 & ~x82 & ~x84 & ~x85 & ~x86 & ~x111 & ~x112 & ~x141 & ~x197 & ~x224 & ~x250 & ~x251 & ~x257 & ~x279 & ~x280 & ~x283 & ~x290 & ~x307 & ~x332 & ~x333 & ~x357 & ~x358 & ~x361 & ~x362 & ~x368 & ~x386 & ~x387 & ~x392 & ~x445 & ~x447 & ~x465 & ~x532 & ~x533 & ~x562 & ~x588 & ~x589 & ~x618 & ~x641 & ~x646 & ~x664 & ~x671 & ~x684 & ~x687 & ~x697 & ~x701 & ~x702 & ~x709 & ~x713 & ~x718 & ~x726 & ~x729 & ~x734 & ~x737 & ~x739 & ~x740 & ~x748 & ~x752 & ~x760 & ~x763 & ~x764 & ~x766 & ~x768 & ~x774 & ~x777 & ~x779 & ~x782;
assign c0225 =  x235 &  x376 &  x380 & ~x130 & ~x505;
assign c0227 =  x490 &  x491 & ~x4 & ~x11 & ~x37 & ~x46 & ~x65 & ~x73 & ~x80 & ~x86 & ~x88 & ~x102 & ~x106 & ~x110 & ~x111 & ~x135 & ~x141 & ~x169 & ~x171 & ~x172 & ~x173 & ~x191 & ~x192 & ~x196 & ~x221 & ~x227 & ~x228 & ~x251 & ~x253 & ~x254 & ~x278 & ~x281 & ~x307 & ~x321 & ~x338 & ~x387 & ~x422 & ~x474 & ~x475 & ~x534 & ~x559 & ~x586 & ~x587 & ~x592 & ~x614 & ~x619 & ~x621 & ~x622 & ~x645 & ~x646 & ~x649 & ~x674 & ~x696 & ~x698 & ~x699 & ~x701 & ~x703 & ~x718 & ~x725 & ~x731 & ~x739 & ~x743 & ~x752 & ~x769 & ~x772 & ~x774;
assign c0229 =  x351 & ~x14 & ~x21 & ~x23 & ~x24 & ~x25 & ~x49 & ~x58 & ~x61 & ~x70 & ~x79 & ~x113 & ~x118 & ~x220 & ~x221 & ~x222 & ~x267 & ~x280 & ~x283 & ~x294 & ~x335 & ~x360 & ~x391 & ~x393 & ~x420 & ~x506 & ~x613 & ~x616 & ~x641 & ~x644 & ~x648 & ~x674 & ~x675 & ~x676 & ~x678 & ~x690 & ~x729 & ~x753;
assign c0231 =  x352 &  x377 & ~x11 & ~x15 & ~x22 & ~x49 & ~x56 & ~x57 & ~x66 & ~x74 & ~x77 & ~x82 & ~x89 & ~x116 & ~x140 & ~x169 & ~x222 & ~x281 & ~x304 & ~x329 & ~x476 & ~x477 & ~x488 & ~x491 & ~x556 & ~x557 & ~x588 & ~x614 & ~x748 & ~x761;
assign c0233 =  x461 &  x518 &  x567;
assign c0235 =  x466 &  x545 & ~x370 & ~x402 & ~x426 & ~x443;
assign c0237 =  x542 &  x573 & ~x53 & ~x170 & ~x173 & ~x242 & ~x255 & ~x268 & ~x365 & ~x529 & ~x592 & ~x652 & ~x674 & ~x695 & ~x718 & ~x753;
assign c0239 =  x408 & ~x2 & ~x3 & ~x11 & ~x12 & ~x17 & ~x20 & ~x35 & ~x37 & ~x44 & ~x51 & ~x60 & ~x81 & ~x110 & ~x141 & ~x164 & ~x170 & ~x192 & ~x195 & ~x197 & ~x198 & ~x200 & ~x223 & ~x224 & ~x227 & ~x252 & ~x280 & ~x337 & ~x473 & ~x478 & ~x533 & ~x535 & ~x585 & ~x587 & ~x595 & ~x611 & ~x613 & ~x644 & ~x652 & ~x654 & ~x655 & ~x657 & ~x677 & ~x679 & ~x700 & ~x703 & ~x713 & ~x761 & ~x767 & ~x774 & ~x776 & ~x782;
assign c0241 =  x157 & ~x25 & ~x33 & ~x34 & ~x50 & ~x51 & ~x68 & ~x86 & ~x87 & ~x93 & ~x95 & ~x98 & ~x109 & ~x138 & ~x145 & ~x170 & ~x173 & ~x197 & ~x221 & ~x249 & ~x253 & ~x254 & ~x255 & ~x285 & ~x286 & ~x299 & ~x300 & ~x303 & ~x308 & ~x330 & ~x331 & ~x357 & ~x368 & ~x389 & ~x390 & ~x391 & ~x421 & ~x436 & ~x451 & ~x558 & ~x559 & ~x615 & ~x616 & ~x647 & ~x661 & ~x672 & ~x689 & ~x695 & ~x696 & ~x700 & ~x709 & ~x713 & ~x718 & ~x728 & ~x734 & ~x736 & ~x745 & ~x758 & ~x776 & ~x779 & ~x783;
assign c0243 =  x107;
assign c0245 =  x352 &  x378 & ~x21 & ~x46 & ~x385;
assign c0247 = ~x0 & ~x9 & ~x27 & ~x63 & ~x91 & ~x129 & ~x182 & ~x183 & ~x184 & ~x227 & ~x305 & ~x399 & ~x425 & ~x426 & ~x453 & ~x456 & ~x512 & ~x605 & ~x659 & ~x670;
assign c0249 =  x352 &  x353 &  x377 &  x378 &  x379 &  x404 & ~x97;
assign c0251 = ~x14 & ~x20 & ~x27 & ~x31 & ~x38 & ~x48 & ~x74 & ~x76 & ~x78 & ~x99 & ~x102 & ~x108 & ~x116 & ~x194 & ~x195 & ~x203 & ~x285 & ~x311 & ~x312 & ~x334 & ~x338 & ~x339 & ~x340 & ~x366 & ~x386 & ~x411 & ~x412 & ~x413 & ~x414 & ~x415 & ~x438 & ~x449 & ~x469 & ~x473 & ~x497 & ~x554 & ~x670 & ~x673 & ~x705 & ~x742 & ~x761;
assign c0253 =  x376 &  x378 &  x379 &  x380 & ~x5 & ~x10 & ~x44 & ~x54 & ~x61 & ~x73 & ~x78 & ~x94 & ~x121 & ~x366 & ~x388 & ~x423 & ~x506 & ~x515 & ~x535 & ~x557 & ~x644 & ~x650 & ~x698 & ~x722 & ~x728 & ~x769;
assign c0255 =  x434 &  x436 & ~x324 & ~x443 & ~x674;
assign c0257 =  x539 &  x596 &  x597 &  x598 & ~x1 & ~x2 & ~x5 & ~x9 & ~x13 & ~x14 & ~x15 & ~x16 & ~x19 & ~x32 & ~x34 & ~x36 & ~x39 & ~x50 & ~x60 & ~x61 & ~x65 & ~x71 & ~x74 & ~x77 & ~x78 & ~x79 & ~x83 & ~x84 & ~x87 & ~x90 & ~x106 & ~x109 & ~x112 & ~x113 & ~x114 & ~x134 & ~x140 & ~x142 & ~x143 & ~x161 & ~x170 & ~x171 & ~x193 & ~x194 & ~x196 & ~x197 & ~x198 & ~x221 & ~x222 & ~x223 & ~x224 & ~x225 & ~x227 & ~x228 & ~x252 & ~x253 & ~x276 & ~x278 & ~x280 & ~x281 & ~x282 & ~x285 & ~x303 & ~x308 & ~x309 & ~x316 & ~x333 & ~x334 & ~x337 & ~x338 & ~x339 & ~x341 & ~x343 & ~x362 & ~x367 & ~x368 & ~x369 & ~x370 & ~x371 & ~x387 & ~x392 & ~x397 & ~x399 & ~x400 & ~x419 & ~x424 & ~x450 & ~x473 & ~x474 & ~x478 & ~x533 & ~x560 & ~x588 & ~x590 & ~x613 & ~x614 & ~x619 & ~x638 & ~x639 & ~x640 & ~x644 & ~x645 & ~x669 & ~x671 & ~x679 & ~x680 & ~x683 & ~x685 & ~x686 & ~x687 & ~x689 & ~x690 & ~x692 & ~x693 & ~x695 & ~x702 & ~x707 & ~x712 & ~x713 & ~x714 & ~x718 & ~x721 & ~x724 & ~x726 & ~x730 & ~x737 & ~x742 & ~x749 & ~x751 & ~x753 & ~x755 & ~x759 & ~x763 & ~x767 & ~x769 & ~x770 & ~x774 & ~x775 & ~x776 & ~x777;
assign c0259 =  x492 & ~x20 & ~x28 & ~x39 & ~x63 & ~x89 & ~x136 & ~x141 & ~x171 & ~x337 & ~x339 & ~x352 & ~x353 & ~x354 & ~x378 & ~x389 & ~x415 & ~x425 & ~x443 & ~x503 & ~x586 & ~x640 & ~x694 & ~x713 & ~x732 & ~x749 & ~x775;
assign c0261 =  x713;
assign c0263 =  x158 &  x577 & ~x48 & ~x386 & ~x394 & ~x396 & ~x401 & ~x682 & ~x740;
assign c0265 =  x507;
assign c0267 =  x100;
assign c0269 =  x462 &  x463 &  x492 &  x548 &  x576 & ~x24 & ~x61 & ~x114 & ~x280 & ~x305 & ~x332 & ~x365 & ~x395 & ~x530 & ~x612 & ~x617 & ~x628 & ~x695 & ~x754 & ~x768 & ~x778;
assign c0271 =  x406 &  x407 & ~x178 & ~x297;
assign c0273 =  x488 & ~x5 & ~x18 & ~x32 & ~x37 & ~x77 & ~x139 & ~x140 & ~x141 & ~x230 & ~x254 & ~x286 & ~x311 & ~x314 & ~x325 & ~x326 & ~x369 & ~x378 & ~x387 & ~x414 & ~x442 & ~x470 & ~x500 & ~x502 & ~x506 & ~x590 & ~x613 & ~x752 & ~x759;
assign c0275 =  x494 &  x523 & ~x1 & ~x2 & ~x8 & ~x18 & ~x19 & ~x28 & ~x33 & ~x35 & ~x42 & ~x56 & ~x74 & ~x82 & ~x88 & ~x110 & ~x117 & ~x143 & ~x225 & ~x277 & ~x283 & ~x309 & ~x368 & ~x416 & ~x476 & ~x501 & ~x503 & ~x505 & ~x506 & ~x533 & ~x560 & ~x562 & ~x588 & ~x630 & ~x651 & ~x658 & ~x677 & ~x680 & ~x699 & ~x705 & ~x724 & ~x733 & ~x747 & ~x762 & ~x778;
assign c0277 =  x607 & ~x301 & ~x359 & ~x425 & ~x426;
assign c0279 =  x708;
assign c0281 =  x434 &  x461 & ~x11 & ~x15 & ~x21 & ~x23 & ~x35 & ~x39 & ~x43 & ~x44 & ~x54 & ~x58 & ~x63 & ~x80 & ~x82 & ~x83 & ~x90 & ~x108 & ~x115 & ~x140 & ~x141 & ~x220 & ~x254 & ~x280 & ~x365 & ~x385 & ~x391 & ~x395 & ~x419 & ~x421 & ~x423 & ~x475 & ~x498 & ~x507 & ~x532 & ~x534 & ~x557 & ~x560 & ~x563 & ~x614 & ~x643 & ~x671 & ~x675 & ~x678 & ~x730 & ~x734 & ~x736 & ~x740 & ~x744 & ~x752 & ~x753 & ~x782;
assign c0283 = ~x1 & ~x6 & ~x11 & ~x17 & ~x23 & ~x25 & ~x27 & ~x47 & ~x50 & ~x51 & ~x62 & ~x65 & ~x69 & ~x76 & ~x77 & ~x79 & ~x81 & ~x85 & ~x87 & ~x93 & ~x97 & ~x108 & ~x115 & ~x144 & ~x165 & ~x167 & ~x195 & ~x196 & ~x199 & ~x220 & ~x221 & ~x247 & ~x253 & ~x274 & ~x280 & ~x282 & ~x299 & ~x301 & ~x302 & ~x332 & ~x336 & ~x361 & ~x367 & ~x390 & ~x396 & ~x417 & ~x449 & ~x460 & ~x461 & ~x487 & ~x489 & ~x506 & ~x514 & ~x515 & ~x517 & ~x530 & ~x532 & ~x535 & ~x560 & ~x562 & ~x586 & ~x587 & ~x613 & ~x643 & ~x644 & ~x645 & ~x648 & ~x671 & ~x673 & ~x674 & ~x675 & ~x679 & ~x697 & ~x708 & ~x722 & ~x726 & ~x727 & ~x729 & ~x730 & ~x754 & ~x758 & ~x763 & ~x769 & ~x774 & ~x776 & ~x778 & ~x779 & ~x780 & ~x782 & ~x783;
assign c0285 = ~x11 & ~x17 & ~x19 & ~x21 & ~x53 & ~x60 & ~x68 & ~x79 & ~x80 & ~x87 & ~x91 & ~x128 & ~x129 & ~x145 & ~x153 & ~x154 & ~x155 & ~x157 & ~x167 & ~x179 & ~x224 & ~x360 & ~x388 & ~x390 & ~x415 & ~x417 & ~x420 & ~x475 & ~x500 & ~x510 & ~x526 & ~x527 & ~x531 & ~x537 & ~x542 & ~x554 & ~x565 & ~x568 & ~x592 & ~x642 & ~x671 & ~x700 & ~x732 & ~x733 & ~x753 & ~x759;
assign c0287 =  x448;
assign c0289 =  x407 &  x408 & ~x0 & ~x13 & ~x54 & ~x68 & ~x114 & ~x137 & ~x166 & ~x167 & ~x172 & ~x174 & ~x200 & ~x201 & ~x254 & ~x280 & ~x324 & ~x351 & ~x422 & ~x447 & ~x448 & ~x474 & ~x530 & ~x589 & ~x590 & ~x614 & ~x619 & ~x669 & ~x675 & ~x692 & ~x694 & ~x699 & ~x700 & ~x709 & ~x727 & ~x736 & ~x739 & ~x752 & ~x769;
assign c0291 =  x602 & ~x4 & ~x10 & ~x12 & ~x22 & ~x37 & ~x38 & ~x43 & ~x62 & ~x109 & ~x111 & ~x163 & ~x187 & ~x225 & ~x240 & ~x242 & ~x283 & ~x306 & ~x447 & ~x474 & ~x504 & ~x508 & ~x584 & ~x617 & ~x637 & ~x638 & ~x641 & ~x646 & ~x668 & ~x675 & ~x686 & ~x736 & ~x743 & ~x757 & ~x762 & ~x772 & ~x775;
assign c0293 =  x572 & ~x25 & ~x217 & ~x240 & ~x253 & ~x315 & ~x342 & ~x368 & ~x504 & ~x616;
assign c0295 =  x380 & ~x0 & ~x2 & ~x3 & ~x6 & ~x9 & ~x17 & ~x18 & ~x22 & ~x24 & ~x27 & ~x32 & ~x36 & ~x46 & ~x48 & ~x49 & ~x57 & ~x68 & ~x76 & ~x80 & ~x83 & ~x85 & ~x90 & ~x113 & ~x115 & ~x137 & ~x169 & ~x192 & ~x194 & ~x197 & ~x200 & ~x220 & ~x254 & ~x266 & ~x281 & ~x282 & ~x307 & ~x363 & ~x419 & ~x423 & ~x478 & ~x488 & ~x502 & ~x505 & ~x614 & ~x616 & ~x643 & ~x670 & ~x676 & ~x690 & ~x691 & ~x693 & ~x696 & ~x698 & ~x704 & ~x707 & ~x708 & ~x716 & ~x717 & ~x721 & ~x736 & ~x740 & ~x745 & ~x752 & ~x760 & ~x761 & ~x762 & ~x764 & ~x767 & ~x776 & ~x777 & ~x780;
assign c0297 =  x461;
assign c0299 =  x179 &  x491 & ~x7 & ~x41 & ~x658 & ~x751;
assign c10 = ~x0 & ~x6 & ~x9 & ~x10 & ~x11 & ~x12 & ~x15 & ~x16 & ~x18 & ~x19 & ~x22 & ~x23 & ~x26 & ~x27 & ~x28 & ~x29 & ~x30 & ~x33 & ~x34 & ~x36 & ~x37 & ~x39 & ~x40 & ~x41 & ~x42 & ~x43 & ~x45 & ~x46 & ~x47 & ~x49 & ~x51 & ~x54 & ~x55 & ~x57 & ~x58 & ~x60 & ~x64 & ~x65 & ~x67 & ~x69 & ~x73 & ~x74 & ~x76 & ~x78 & ~x81 & ~x82 & ~x84 & ~x86 & ~x87 & ~x88 & ~x89 & ~x90 & ~x93 & ~x94 & ~x96 & ~x98 & ~x99 & ~x101 & ~x103 & ~x105 & ~x107 & ~x108 & ~x109 & ~x111 & ~x112 & ~x114 & ~x116 & ~x117 & ~x118 & ~x121 & ~x124 & ~x128 & ~x135 & ~x136 & ~x138 & ~x139 & ~x140 & ~x143 & ~x144 & ~x145 & ~x148 & ~x149 & ~x153 & ~x154 & ~x156 & ~x166 & ~x167 & ~x168 & ~x169 & ~x170 & ~x174 & ~x193 & ~x194 & ~x195 & ~x197 & ~x199 & ~x203 & ~x204 & ~x205 & ~x207 & ~x208 & ~x209 & ~x210 & ~x221 & ~x223 & ~x225 & ~x229 & ~x230 & ~x235 & ~x236 & ~x237 & ~x238 & ~x248 & ~x249 & ~x251 & ~x254 & ~x256 & ~x259 & ~x260 & ~x261 & ~x262 & ~x263 & ~x264 & ~x265 & ~x266 & ~x277 & ~x278 & ~x280 & ~x281 & ~x282 & ~x284 & ~x287 & ~x288 & ~x289 & ~x290 & ~x291 & ~x292 & ~x293 & ~x303 & ~x304 & ~x306 & ~x307 & ~x308 & ~x309 & ~x314 & ~x318 & ~x319 & ~x320 & ~x329 & ~x330 & ~x331 & ~x336 & ~x338 & ~x339 & ~x341 & ~x343 & ~x344 & ~x345 & ~x346 & ~x347 & ~x355 & ~x356 & ~x358 & ~x359 & ~x360 & ~x362 & ~x363 & ~x364 & ~x365 & ~x369 & ~x371 & ~x372 & ~x373 & ~x383 & ~x384 & ~x386 & ~x387 & ~x394 & ~x397 & ~x398 & ~x399 & ~x400 & ~x409 & ~x410 & ~x412 & ~x419 & ~x423 & ~x424 & ~x425 & ~x437 & ~x438 & ~x439 & ~x440 & ~x441 & ~x442 & ~x443 & ~x452 & ~x465 & ~x466 & ~x467 & ~x470 & ~x471 & ~x473 & ~x475 & ~x492 & ~x493 & ~x496 & ~x498 & ~x501 & ~x502 & ~x503 & ~x504 & ~x506 & ~x508 & ~x520 & ~x521 & ~x527 & ~x529 & ~x537 & ~x547 & ~x548 & ~x549 & ~x551 & ~x552 & ~x554 & ~x560 & ~x562 & ~x563 & ~x575 & ~x576 & ~x578 & ~x579 & ~x581 & ~x583 & ~x584 & ~x585 & ~x586 & ~x587 & ~x590 & ~x591 & ~x603 & ~x604 & ~x605 & ~x606 & ~x607 & ~x608 & ~x609 & ~x610 & ~x611 & ~x616 & ~x617 & ~x631 & ~x633 & ~x636 & ~x637 & ~x638 & ~x639 & ~x640 & ~x641 & ~x642 & ~x644 & ~x647 & ~x660 & ~x664 & ~x666 & ~x670 & ~x671 & ~x673 & ~x674 & ~x676 & ~x677 & ~x682 & ~x688 & ~x691 & ~x692 & ~x695 & ~x697 & ~x699 & ~x700 & ~x702 & ~x703 & ~x707 & ~x709 & ~x711 & ~x714 & ~x716 & ~x718 & ~x719 & ~x721 & ~x722 & ~x723 & ~x724 & ~x727 & ~x729 & ~x730 & ~x731 & ~x735 & ~x738 & ~x740 & ~x743 & ~x744 & ~x745 & ~x747 & ~x748 & ~x749 & ~x750 & ~x751 & ~x752 & ~x753 & ~x758 & ~x760 & ~x761 & ~x765 & ~x766 & ~x767 & ~x768 & ~x769 & ~x771 & ~x772 & ~x774 & ~x775 & ~x777 & ~x780 & ~x781 & ~x783;
assign c12 =  x265 &  x293 &  x321 & ~x9 & ~x14 & ~x29 & ~x68 & ~x77 & ~x88 & ~x160 & ~x174 & ~x175 & ~x190 & ~x227 & ~x232 & ~x274 & ~x329 & ~x374 & ~x398 & ~x430 & ~x512 & ~x538 & ~x586 & ~x597 & ~x624 & ~x676 & ~x690 & ~x707 & ~x718 & ~x726 & ~x748 & ~x762 & ~x779;
assign c14 =  x294 &  x322 &  x378 & ~x8 & ~x18 & ~x38 & ~x51 & ~x89 & ~x93 & ~x103 & ~x105 & ~x122 & ~x133 & ~x145 & ~x158 & ~x171 & ~x188 & ~x221 & ~x223 & ~x224 & ~x226 & ~x228 & ~x241 & ~x242 & ~x243 & ~x253 & ~x269 & ~x270 & ~x274 & ~x278 & ~x280 & ~x284 & ~x285 & ~x326 & ~x354 & ~x365 & ~x388 & ~x389 & ~x426 & ~x438 & ~x443 & ~x444 & ~x458 & ~x506 & ~x508 & ~x534 & ~x565 & ~x582 & ~x584 & ~x585 & ~x586 & ~x608 & ~x617 & ~x618 & ~x665 & ~x672 & ~x674 & ~x675 & ~x676 & ~x700 & ~x711 & ~x714 & ~x716 & ~x724 & ~x737 & ~x738 & ~x742 & ~x749 & ~x752 & ~x756 & ~x757 & ~x761 & ~x773 & ~x777 & ~x778 & ~x781;
assign c16 =  x724;
assign c18 =  x407 & ~x5 & ~x12 & ~x13 & ~x27 & ~x31 & ~x42 & ~x53 & ~x57 & ~x61 & ~x130 & ~x137 & ~x149 & ~x165 & ~x166 & ~x171 & ~x177 & ~x196 & ~x202 & ~x204 & ~x228 & ~x250 & ~x258 & ~x263 & ~x277 & ~x278 & ~x283 & ~x304 & ~x314 & ~x316 & ~x328 & ~x330 & ~x337 & ~x343 & ~x359 & ~x364 & ~x367 & ~x383 & ~x384 & ~x385 & ~x396 & ~x403 & ~x419 & ~x420 & ~x440 & ~x441 & ~x449 & ~x456 & ~x458 & ~x472 & ~x476 & ~x486 & ~x504 & ~x510 & ~x537 & ~x557 & ~x564 & ~x566 & ~x568 & ~x581 & ~x582 & ~x588 & ~x614 & ~x616 & ~x643 & ~x646 & ~x648 & ~x649 & ~x650 & ~x667 & ~x669 & ~x689 & ~x702 & ~x710 & ~x716 & ~x720 & ~x725 & ~x744 & ~x755 & ~x768 & ~x778 & ~x779;
assign c110 =  x562;
assign c112 =  x19;
assign c114 =  x503;
assign c116 =  x239 &  x240 &  x295 &  x323 &  x324 &  x350 &  x406 &  x407 &  x461 &  x489 &  x517 &  x545 & ~x0 & ~x4 & ~x10 & ~x25 & ~x27 & ~x28 & ~x31 & ~x33 & ~x45 & ~x53 & ~x59 & ~x61 & ~x64 & ~x66 & ~x75 & ~x78 & ~x81 & ~x83 & ~x88 & ~x90 & ~x97 & ~x101 & ~x106 & ~x107 & ~x113 & ~x119 & ~x121 & ~x123 & ~x131 & ~x135 & ~x136 & ~x139 & ~x140 & ~x142 & ~x144 & ~x146 & ~x148 & ~x149 & ~x151 & ~x161 & ~x164 & ~x165 & ~x166 & ~x167 & ~x171 & ~x173 & ~x192 & ~x195 & ~x202 & ~x204 & ~x206 & ~x216 & ~x219 & ~x223 & ~x229 & ~x234 & ~x244 & ~x250 & ~x254 & ~x255 & ~x260 & ~x272 & ~x279 & ~x281 & ~x282 & ~x286 & ~x288 & ~x289 & ~x304 & ~x305 & ~x311 & ~x316 & ~x341 & ~x342 & ~x358 & ~x363 & ~x364 & ~x365 & ~x366 & ~x367 & ~x371 & ~x372 & ~x384 & ~x385 & ~x387 & ~x391 & ~x393 & ~x394 & ~x399 & ~x415 & ~x417 & ~x418 & ~x419 & ~x420 & ~x423 & ~x426 & ~x427 & ~x442 & ~x445 & ~x447 & ~x448 & ~x456 & ~x470 & ~x471 & ~x476 & ~x481 & ~x482 & ~x508 & ~x525 & ~x528 & ~x531 & ~x532 & ~x536 & ~x540 & ~x551 & ~x559 & ~x560 & ~x561 & ~x563 & ~x564 & ~x565 & ~x581 & ~x583 & ~x585 & ~x588 & ~x590 & ~x591 & ~x592 & ~x594 & ~x595 & ~x607 & ~x610 & ~x615 & ~x621 & ~x641 & ~x643 & ~x650 & ~x651 & ~x667 & ~x676 & ~x689 & ~x693 & ~x696 & ~x699 & ~x709 & ~x722 & ~x723 & ~x725 & ~x726 & ~x728 & ~x730 & ~x735 & ~x737 & ~x738 & ~x739 & ~x740 & ~x744 & ~x747 & ~x748 & ~x749 & ~x755 & ~x759 & ~x761 & ~x762 & ~x766 & ~x770 & ~x771 & ~x772 & ~x776 & ~x778 & ~x781 & ~x782 & ~x783;
assign c118 =  x379 & ~x5 & ~x12 & ~x21 & ~x27 & ~x34 & ~x39 & ~x40 & ~x53 & ~x57 & ~x71 & ~x73 & ~x76 & ~x84 & ~x117 & ~x119 & ~x136 & ~x141 & ~x145 & ~x162 & ~x167 & ~x218 & ~x219 & ~x220 & ~x242 & ~x262 & ~x301 & ~x308 & ~x311 & ~x341 & ~x361 & ~x394 & ~x402 & ~x420 & ~x427 & ~x437 & ~x449 & ~x469 & ~x471 & ~x478 & ~x498 & ~x500 & ~x512 & ~x515 & ~x531 & ~x533 & ~x561 & ~x585 & ~x588 & ~x642 & ~x645 & ~x653 & ~x668 & ~x676 & ~x700 & ~x701 & ~x716 & ~x721 & ~x725 & ~x730 & ~x742 & ~x746 & ~x751 & ~x754 & ~x755 & ~x758 & ~x764;
assign c120 =  x448;
assign c122 =  x42;
assign c124 =  x325 &  x352 & ~x0 & ~x1 & ~x2 & ~x4 & ~x5 & ~x6 & ~x7 & ~x8 & ~x10 & ~x13 & ~x14 & ~x16 & ~x19 & ~x20 & ~x25 & ~x26 & ~x28 & ~x30 & ~x32 & ~x37 & ~x39 & ~x41 & ~x42 & ~x44 & ~x47 & ~x51 & ~x54 & ~x56 & ~x60 & ~x62 & ~x63 & ~x66 & ~x67 & ~x70 & ~x72 & ~x73 & ~x76 & ~x80 & ~x82 & ~x83 & ~x86 & ~x87 & ~x88 & ~x90 & ~x92 & ~x96 & ~x97 & ~x98 & ~x99 & ~x100 & ~x101 & ~x108 & ~x110 & ~x111 & ~x114 & ~x116 & ~x117 & ~x123 & ~x125 & ~x126 & ~x128 & ~x137 & ~x138 & ~x139 & ~x141 & ~x143 & ~x144 & ~x147 & ~x149 & ~x150 & ~x151 & ~x152 & ~x154 & ~x155 & ~x156 & ~x167 & ~x169 & ~x170 & ~x171 & ~x173 & ~x174 & ~x175 & ~x178 & ~x181 & ~x182 & ~x183 & ~x195 & ~x199 & ~x200 & ~x202 & ~x203 & ~x208 & ~x210 & ~x221 & ~x222 & ~x223 & ~x224 & ~x225 & ~x226 & ~x227 & ~x228 & ~x229 & ~x231 & ~x234 & ~x235 & ~x236 & ~x237 & ~x238 & ~x239 & ~x248 & ~x251 & ~x252 & ~x254 & ~x258 & ~x262 & ~x264 & ~x265 & ~x266 & ~x275 & ~x277 & ~x279 & ~x281 & ~x283 & ~x285 & ~x287 & ~x288 & ~x292 & ~x293 & ~x303 & ~x304 & ~x305 & ~x306 & ~x308 & ~x313 & ~x317 & ~x318 & ~x319 & ~x320 & ~x321 & ~x332 & ~x335 & ~x336 & ~x337 & ~x338 & ~x340 & ~x342 & ~x343 & ~x345 & ~x346 & ~x347 & ~x348 & ~x357 & ~x358 & ~x365 & ~x366 & ~x368 & ~x370 & ~x371 & ~x374 & ~x385 & ~x386 & ~x387 & ~x389 & ~x391 & ~x395 & ~x397 & ~x398 & ~x399 & ~x400 & ~x401 & ~x415 & ~x419 & ~x420 & ~x421 & ~x425 & ~x426 & ~x427 & ~x429 & ~x438 & ~x440 & ~x444 & ~x445 & ~x446 & ~x447 & ~x448 & ~x450 & ~x451 & ~x452 & ~x454 & ~x455 & ~x469 & ~x471 & ~x475 & ~x476 & ~x480 & ~x481 & ~x482 & ~x496 & ~x498 & ~x499 & ~x502 & ~x504 & ~x506 & ~x507 & ~x508 & ~x510 & ~x520 & ~x521 & ~x522 & ~x523 & ~x524 & ~x526 & ~x528 & ~x529 & ~x530 & ~x531 & ~x533 & ~x534 & ~x536 & ~x537 & ~x550 & ~x551 & ~x554 & ~x555 & ~x556 & ~x557 & ~x558 & ~x559 & ~x563 & ~x575 & ~x576 & ~x577 & ~x578 & ~x581 & ~x582 & ~x584 & ~x585 & ~x586 & ~x589 & ~x591 & ~x604 & ~x605 & ~x606 & ~x608 & ~x614 & ~x615 & ~x619 & ~x620 & ~x631 & ~x634 & ~x635 & ~x636 & ~x638 & ~x640 & ~x641 & ~x644 & ~x658 & ~x659 & ~x665 & ~x670 & ~x672 & ~x673 & ~x674 & ~x675 & ~x676 & ~x686 & ~x688 & ~x689 & ~x694 & ~x700 & ~x701 & ~x703 & ~x704 & ~x705 & ~x707 & ~x709 & ~x710 & ~x711 & ~x714 & ~x715 & ~x716 & ~x717 & ~x718 & ~x720 & ~x721 & ~x722 & ~x724 & ~x726 & ~x727 & ~x728 & ~x729 & ~x732 & ~x733 & ~x734 & ~x735 & ~x738 & ~x739 & ~x740 & ~x741 & ~x742 & ~x744 & ~x746 & ~x747 & ~x753 & ~x757 & ~x758 & ~x759 & ~x760 & ~x763 & ~x764 & ~x766 & ~x768 & ~x770 & ~x771 & ~x773 & ~x776 & ~x777 & ~x779 & ~x781 & ~x782 & ~x783;
assign c126 =  x17;
assign c128 =  x293 &  x516 &  x545 & ~x15 & ~x16 & ~x18 & ~x22 & ~x25 & ~x32 & ~x48 & ~x50 & ~x60 & ~x61 & ~x70 & ~x81 & ~x90 & ~x93 & ~x111 & ~x147 & ~x172 & ~x175 & ~x190 & ~x197 & ~x201 & ~x204 & ~x215 & ~x217 & ~x218 & ~x233 & ~x243 & ~x244 & ~x250 & ~x253 & ~x254 & ~x271 & ~x280 & ~x313 & ~x326 & ~x331 & ~x333 & ~x334 & ~x336 & ~x341 & ~x359 & ~x374 & ~x414 & ~x452 & ~x473 & ~x482 & ~x484 & ~x485 & ~x486 & ~x503 & ~x528 & ~x582 & ~x613 & ~x635 & ~x636 & ~x664 & ~x674 & ~x677 & ~x693 & ~x705 & ~x711 & ~x712 & ~x735 & ~x764 & ~x766;
assign c130 =  x462 & ~x9 & ~x14 & ~x16 & ~x19 & ~x37 & ~x50 & ~x51 & ~x57 & ~x80 & ~x85 & ~x87 & ~x108 & ~x130 & ~x133 & ~x134 & ~x136 & ~x164 & ~x173 & ~x231 & ~x233 & ~x251 & ~x256 & ~x273 & ~x297 & ~x306 & ~x309 & ~x331 & ~x381 & ~x383 & ~x393 & ~x398 & ~x429 & ~x430 & ~x442 & ~x447 & ~x456 & ~x466 & ~x469 & ~x472 & ~x486 & ~x487 & ~x511 & ~x583 & ~x585 & ~x591 & ~x640 & ~x643 & ~x651 & ~x654 & ~x688 & ~x696 & ~x711 & ~x718 & ~x722 & ~x730 & ~x745 & ~x758 & ~x766 & ~x774 & ~x781;
assign c132 = ~x13 & ~x29 & ~x30 & ~x61 & ~x93 & ~x102 & ~x110 & ~x135 & ~x146 & ~x167 & ~x171 & ~x177 & ~x179 & ~x218 & ~x231 & ~x235 & ~x246 & ~x248 & ~x251 & ~x256 & ~x260 & ~x302 & ~x314 & ~x354 & ~x363 & ~x425 & ~x429 & ~x487 & ~x589 & ~x595 & ~x650 & ~x652 & ~x666 & ~x674 & ~x693 & ~x702 & ~x726 & ~x756;
assign c134 =  x324 &  x325 &  x351 &  x352 &  x434 & ~x1 & ~x4 & ~x5 & ~x8 & ~x9 & ~x10 & ~x12 & ~x14 & ~x17 & ~x18 & ~x19 & ~x20 & ~x21 & ~x23 & ~x24 & ~x25 & ~x26 & ~x27 & ~x28 & ~x30 & ~x35 & ~x37 & ~x39 & ~x41 & ~x42 & ~x48 & ~x49 & ~x53 & ~x55 & ~x56 & ~x60 & ~x61 & ~x63 & ~x64 & ~x66 & ~x68 & ~x70 & ~x71 & ~x72 & ~x73 & ~x75 & ~x77 & ~x79 & ~x81 & ~x83 & ~x84 & ~x85 & ~x86 & ~x89 & ~x92 & ~x93 & ~x94 & ~x95 & ~x96 & ~x97 & ~x98 & ~x99 & ~x100 & ~x103 & ~x104 & ~x107 & ~x108 & ~x109 & ~x110 & ~x111 & ~x113 & ~x115 & ~x116 & ~x117 & ~x118 & ~x120 & ~x121 & ~x122 & ~x123 & ~x124 & ~x127 & ~x128 & ~x136 & ~x138 & ~x139 & ~x140 & ~x144 & ~x146 & ~x147 & ~x148 & ~x149 & ~x150 & ~x151 & ~x152 & ~x153 & ~x154 & ~x155 & ~x164 & ~x168 & ~x169 & ~x170 & ~x171 & ~x175 & ~x177 & ~x182 & ~x183 & ~x195 & ~x196 & ~x199 & ~x202 & ~x203 & ~x204 & ~x205 & ~x206 & ~x207 & ~x208 & ~x209 & ~x210 & ~x211 & ~x220 & ~x221 & ~x223 & ~x224 & ~x226 & ~x227 & ~x230 & ~x231 & ~x232 & ~x233 & ~x235 & ~x236 & ~x237 & ~x247 & ~x248 & ~x249 & ~x251 & ~x252 & ~x253 & ~x256 & ~x257 & ~x260 & ~x262 & ~x263 & ~x264 & ~x265 & ~x275 & ~x276 & ~x277 & ~x278 & ~x280 & ~x282 & ~x283 & ~x285 & ~x288 & ~x289 & ~x291 & ~x293 & ~x301 & ~x302 & ~x303 & ~x304 & ~x305 & ~x306 & ~x307 & ~x309 & ~x312 & ~x313 & ~x314 & ~x318 & ~x319 & ~x320 & ~x332 & ~x334 & ~x335 & ~x336 & ~x338 & ~x339 & ~x340 & ~x342 & ~x343 & ~x344 & ~x345 & ~x356 & ~x357 & ~x359 & ~x360 & ~x361 & ~x362 & ~x364 & ~x365 & ~x369 & ~x370 & ~x371 & ~x372 & ~x384 & ~x385 & ~x386 & ~x389 & ~x390 & ~x391 & ~x397 & ~x398 & ~x399 & ~x412 & ~x414 & ~x415 & ~x416 & ~x418 & ~x419 & ~x420 & ~x422 & ~x423 & ~x426 & ~x439 & ~x440 & ~x442 & ~x443 & ~x444 & ~x446 & ~x448 & ~x452 & ~x453 & ~x454 & ~x466 & ~x469 & ~x471 & ~x472 & ~x473 & ~x476 & ~x478 & ~x480 & ~x482 & ~x493 & ~x495 & ~x496 & ~x497 & ~x499 & ~x502 & ~x503 & ~x504 & ~x505 & ~x506 & ~x508 & ~x510 & ~x522 & ~x523 & ~x525 & ~x526 & ~x527 & ~x528 & ~x529 & ~x530 & ~x531 & ~x535 & ~x537 & ~x538 & ~x549 & ~x550 & ~x551 & ~x552 & ~x557 & ~x559 & ~x560 & ~x562 & ~x563 & ~x565 & ~x577 & ~x579 & ~x580 & ~x581 & ~x589 & ~x590 & ~x591 & ~x592 & ~x603 & ~x606 & ~x610 & ~x613 & ~x615 & ~x616 & ~x617 & ~x619 & ~x635 & ~x638 & ~x639 & ~x640 & ~x643 & ~x644 & ~x645 & ~x647 & ~x648 & ~x658 & ~x661 & ~x662 & ~x663 & ~x664 & ~x667 & ~x669 & ~x671 & ~x673 & ~x674 & ~x677 & ~x678 & ~x688 & ~x689 & ~x692 & ~x694 & ~x695 & ~x699 & ~x700 & ~x702 & ~x703 & ~x705 & ~x708 & ~x710 & ~x714 & ~x715 & ~x718 & ~x719 & ~x721 & ~x723 & ~x724 & ~x726 & ~x728 & ~x730 & ~x731 & ~x734 & ~x736 & ~x737 & ~x738 & ~x739 & ~x741 & ~x742 & ~x743 & ~x745 & ~x747 & ~x748 & ~x751 & ~x754 & ~x755 & ~x756 & ~x761 & ~x763 & ~x764 & ~x771 & ~x772 & ~x773 & ~x774 & ~x775 & ~x776 & ~x777 & ~x778 & ~x779 & ~x780 & ~x782;
assign c136 =  x756;
assign c138 =  x337;
assign c140 =  x85;
assign c142 =  x241 &  x267 &  x296 &  x323 &  x351 &  x378 &  x460 &  x488 &  x516 &  x517 &  x545 &  x572 & ~x0 & ~x3 & ~x6 & ~x7 & ~x13 & ~x17 & ~x19 & ~x23 & ~x25 & ~x27 & ~x33 & ~x34 & ~x36 & ~x42 & ~x45 & ~x50 & ~x52 & ~x53 & ~x54 & ~x56 & ~x58 & ~x62 & ~x63 & ~x69 & ~x71 & ~x72 & ~x76 & ~x77 & ~x84 & ~x86 & ~x92 & ~x93 & ~x96 & ~x99 & ~x100 & ~x101 & ~x104 & ~x112 & ~x114 & ~x115 & ~x117 & ~x120 & ~x123 & ~x124 & ~x136 & ~x146 & ~x147 & ~x148 & ~x151 & ~x162 & ~x171 & ~x172 & ~x176 & ~x177 & ~x179 & ~x192 & ~x193 & ~x194 & ~x196 & ~x205 & ~x206 & ~x207 & ~x219 & ~x222 & ~x226 & ~x230 & ~x234 & ~x235 & ~x247 & ~x248 & ~x249 & ~x250 & ~x251 & ~x253 & ~x258 & ~x259 & ~x263 & ~x273 & ~x275 & ~x288 & ~x301 & ~x305 & ~x308 & ~x309 & ~x310 & ~x315 & ~x332 & ~x336 & ~x343 & ~x345 & ~x346 & ~x358 & ~x359 & ~x369 & ~x370 & ~x374 & ~x383 & ~x389 & ~x392 & ~x396 & ~x398 & ~x401 & ~x417 & ~x421 & ~x426 & ~x428 & ~x439 & ~x442 & ~x449 & ~x450 & ~x470 & ~x472 & ~x473 & ~x475 & ~x476 & ~x478 & ~x479 & ~x480 & ~x482 & ~x484 & ~x503 & ~x504 & ~x507 & ~x508 & ~x512 & ~x521 & ~x529 & ~x530 & ~x533 & ~x534 & ~x536 & ~x539 & ~x551 & ~x552 & ~x559 & ~x563 & ~x567 & ~x577 & ~x580 & ~x581 & ~x583 & ~x586 & ~x588 & ~x589 & ~x605 & ~x608 & ~x609 & ~x610 & ~x618 & ~x620 & ~x622 & ~x633 & ~x636 & ~x643 & ~x644 & ~x649 & ~x663 & ~x666 & ~x667 & ~x668 & ~x671 & ~x672 & ~x677 & ~x688 & ~x689 & ~x690 & ~x691 & ~x696 & ~x700 & ~x702 & ~x703 & ~x705 & ~x718 & ~x722 & ~x724 & ~x725 & ~x726 & ~x727 & ~x730 & ~x733 & ~x736 & ~x740 & ~x741 & ~x746 & ~x751 & ~x761 & ~x764 & ~x771 & ~x773 & ~x777 & ~x779;
assign c144 =  x671;
assign c146 =  x293 & ~x5 & ~x18 & ~x21 & ~x51 & ~x58 & ~x60 & ~x88 & ~x118 & ~x166 & ~x176 & ~x177 & ~x198 & ~x229 & ~x284 & ~x310 & ~x336 & ~x356 & ~x360 & ~x387 & ~x391 & ~x399 & ~x420 & ~x421 & ~x483 & ~x487 & ~x507 & ~x515 & ~x523 & ~x525 & ~x534 & ~x538 & ~x557 & ~x579 & ~x586 & ~x593 & ~x612 & ~x615 & ~x619 & ~x621 & ~x646 & ~x670 & ~x676 & ~x693 & ~x708 & ~x719 & ~x772 & ~x775 & ~x780;
assign c148 =  x81;
assign c150 = ~x2 & ~x5 & ~x7 & ~x17 & ~x24 & ~x25 & ~x26 & ~x31 & ~x35 & ~x37 & ~x39 & ~x40 & ~x44 & ~x47 & ~x48 & ~x49 & ~x50 & ~x51 & ~x54 & ~x58 & ~x60 & ~x61 & ~x65 & ~x68 & ~x69 & ~x71 & ~x74 & ~x76 & ~x83 & ~x84 & ~x86 & ~x87 & ~x95 & ~x98 & ~x101 & ~x106 & ~x107 & ~x109 & ~x110 & ~x113 & ~x114 & ~x115 & ~x119 & ~x122 & ~x125 & ~x126 & ~x127 & ~x131 & ~x137 & ~x140 & ~x141 & ~x144 & ~x149 & ~x152 & ~x166 & ~x168 & ~x169 & ~x171 & ~x173 & ~x178 & ~x180 & ~x196 & ~x198 & ~x199 & ~x200 & ~x201 & ~x203 & ~x205 & ~x208 & ~x209 & ~x210 & ~x221 & ~x223 & ~x228 & ~x234 & ~x235 & ~x236 & ~x237 & ~x250 & ~x251 & ~x257 & ~x258 & ~x260 & ~x261 & ~x263 & ~x277 & ~x283 & ~x302 & ~x306 & ~x308 & ~x309 & ~x310 & ~x312 & ~x315 & ~x316 & ~x317 & ~x318 & ~x319 & ~x331 & ~x337 & ~x338 & ~x344 & ~x346 & ~x361 & ~x366 & ~x371 & ~x385 & ~x387 & ~x388 & ~x390 & ~x393 & ~x400 & ~x402 & ~x410 & ~x412 & ~x421 & ~x425 & ~x428 & ~x440 & ~x443 & ~x455 & ~x456 & ~x465 & ~x466 & ~x467 & ~x470 & ~x471 & ~x472 & ~x473 & ~x478 & ~x481 & ~x482 & ~x491 & ~x494 & ~x495 & ~x496 & ~x497 & ~x502 & ~x504 & ~x505 & ~x507 & ~x508 & ~x509 & ~x510 & ~x511 & ~x519 & ~x520 & ~x522 & ~x525 & ~x530 & ~x531 & ~x533 & ~x546 & ~x549 & ~x552 & ~x554 & ~x559 & ~x562 & ~x573 & ~x574 & ~x575 & ~x576 & ~x580 & ~x581 & ~x585 & ~x586 & ~x588 & ~x589 & ~x602 & ~x603 & ~x610 & ~x618 & ~x632 & ~x640 & ~x645 & ~x648 & ~x656 & ~x657 & ~x660 & ~x665 & ~x668 & ~x671 & ~x676 & ~x677 & ~x686 & ~x692 & ~x694 & ~x695 & ~x701 & ~x702 & ~x710 & ~x711 & ~x714 & ~x715 & ~x716 & ~x717 & ~x719 & ~x721 & ~x722 & ~x723 & ~x726 & ~x728 & ~x730 & ~x734 & ~x745 & ~x746 & ~x747 & ~x750 & ~x751 & ~x752 & ~x759 & ~x760 & ~x761 & ~x771 & ~x773 & ~x775 & ~x776 & ~x779 & ~x782 & ~x783;
assign c152 =  x326 &  x567 &  x568 &  x622 & ~x156 & ~x184 & ~x211 & ~x265 & ~x266;
assign c154 = ~x10 & ~x37 & ~x42 & ~x48 & ~x50 & ~x56 & ~x81 & ~x84 & ~x106 & ~x132 & ~x147 & ~x170 & ~x172 & ~x190 & ~x202 & ~x204 & ~x251 & ~x252 & ~x269 & ~x278 & ~x280 & ~x346 & ~x361 & ~x408 & ~x437 & ~x458 & ~x485 & ~x493 & ~x512 & ~x513 & ~x526 & ~x541 & ~x553 & ~x556 & ~x560 & ~x567 & ~x584 & ~x611 & ~x649 & ~x650 & ~x668 & ~x669 & ~x686 & ~x709 & ~x710 & ~x719 & ~x730 & ~x732 & ~x737 & ~x746 & ~x763 & ~x764 & ~x778;
assign c156 =  x36;
assign c158 =  x42;
assign c160 =  x434 &  x546 &  x574 & ~x10 & ~x16 & ~x17 & ~x20 & ~x29 & ~x37 & ~x42 & ~x49 & ~x53 & ~x57 & ~x60 & ~x62 & ~x93 & ~x96 & ~x98 & ~x105 & ~x110 & ~x114 & ~x117 & ~x122 & ~x146 & ~x147 & ~x159 & ~x160 & ~x166 & ~x177 & ~x190 & ~x200 & ~x203 & ~x218 & ~x244 & ~x245 & ~x246 & ~x251 & ~x257 & ~x271 & ~x272 & ~x280 & ~x281 & ~x289 & ~x328 & ~x362 & ~x382 & ~x392 & ~x427 & ~x438 & ~x447 & ~x448 & ~x452 & ~x467 & ~x475 & ~x479 & ~x482 & ~x494 & ~x508 & ~x511 & ~x527 & ~x534 & ~x535 & ~x537 & ~x583 & ~x612 & ~x619 & ~x620 & ~x635 & ~x636 & ~x665 & ~x699 & ~x724 & ~x725 & ~x747 & ~x750 & ~x760 & ~x775;
assign c162 = ~x3 & ~x12 & ~x14 & ~x16 & ~x24 & ~x29 & ~x47 & ~x50 & ~x51 & ~x56 & ~x64 & ~x68 & ~x71 & ~x102 & ~x113 & ~x129 & ~x158 & ~x170 & ~x219 & ~x232 & ~x250 & ~x269 & ~x273 & ~x277 & ~x278 & ~x285 & ~x299 & ~x314 & ~x327 & ~x336 & ~x337 & ~x338 & ~x359 & ~x360 & ~x420 & ~x422 & ~x446 & ~x474 & ~x480 & ~x481 & ~x506 & ~x509 & ~x531 & ~x537 & ~x539 & ~x542 & ~x559 & ~x584 & ~x613 & ~x616 & ~x641 & ~x647 & ~x685 & ~x688 & ~x692 & ~x696 & ~x697 & ~x702 & ~x709 & ~x714 & ~x715 & ~x719 & ~x740 & ~x744 & ~x755 & ~x760 & ~x766 & ~x767 & ~x773 & ~x779;
assign c164 = ~x4 & ~x7 & ~x25 & ~x28 & ~x34 & ~x51 & ~x53 & ~x57 & ~x60 & ~x66 & ~x80 & ~x89 & ~x109 & ~x122 & ~x137 & ~x159 & ~x179 & ~x189 & ~x195 & ~x197 & ~x232 & ~x269 & ~x298 & ~x341 & ~x353 & ~x354 & ~x400 & ~x443 & ~x451 & ~x464 & ~x557 & ~x617 & ~x652 & ~x674 & ~x680 & ~x739 & ~x743 & ~x747 & ~x764;
assign c166 =  x762;
assign c168 =  x518 &  x603 & ~x3 & ~x6 & ~x17 & ~x33 & ~x36 & ~x37 & ~x40 & ~x49 & ~x68 & ~x72 & ~x81 & ~x88 & ~x91 & ~x94 & ~x101 & ~x103 & ~x104 & ~x105 & ~x110 & ~x118 & ~x122 & ~x130 & ~x132 & ~x138 & ~x140 & ~x141 & ~x142 & ~x146 & ~x149 & ~x160 & ~x188 & ~x189 & ~x194 & ~x195 & ~x215 & ~x218 & ~x220 & ~x224 & ~x249 & ~x257 & ~x277 & ~x304 & ~x318 & ~x328 & ~x338 & ~x339 & ~x343 & ~x367 & ~x368 & ~x371 & ~x382 & ~x395 & ~x424 & ~x430 & ~x441 & ~x444 & ~x457 & ~x458 & ~x481 & ~x485 & ~x497 & ~x509 & ~x533 & ~x539 & ~x562 & ~x592 & ~x593 & ~x594 & ~x620 & ~x646 & ~x647 & ~x670 & ~x678 & ~x679 & ~x683 & ~x691 & ~x692 & ~x698 & ~x701 & ~x703 & ~x706 & ~x711 & ~x715 & ~x719 & ~x723 & ~x725 & ~x729 & ~x733 & ~x734 & ~x742 & ~x759 & ~x765 & ~x771 & ~x775 & ~x780 & ~x781;
assign c170 =  x325 &  x326 &  x352 &  x353 &  x379 &  x380 &  x406 &  x433 &  x461 &  x487 &  x488 &  x515 &  x542 &  x569 & ~x0 & ~x3 & ~x6 & ~x8 & ~x20 & ~x21 & ~x26 & ~x28 & ~x29 & ~x30 & ~x31 & ~x36 & ~x38 & ~x43 & ~x45 & ~x46 & ~x52 & ~x56 & ~x57 & ~x58 & ~x63 & ~x64 & ~x70 & ~x72 & ~x74 & ~x79 & ~x81 & ~x83 & ~x85 & ~x88 & ~x90 & ~x95 & ~x98 & ~x99 & ~x100 & ~x101 & ~x102 & ~x106 & ~x109 & ~x110 & ~x118 & ~x119 & ~x121 & ~x122 & ~x126 & ~x127 & ~x128 & ~x136 & ~x139 & ~x140 & ~x141 & ~x142 & ~x143 & ~x144 & ~x147 & ~x148 & ~x150 & ~x151 & ~x154 & ~x156 & ~x165 & ~x166 & ~x167 & ~x168 & ~x173 & ~x174 & ~x175 & ~x176 & ~x178 & ~x179 & ~x181 & ~x182 & ~x183 & ~x195 & ~x196 & ~x199 & ~x200 & ~x201 & ~x203 & ~x205 & ~x208 & ~x209 & ~x210 & ~x230 & ~x231 & ~x232 & ~x234 & ~x235 & ~x236 & ~x237 & ~x249 & ~x250 & ~x251 & ~x254 & ~x257 & ~x258 & ~x259 & ~x260 & ~x262 & ~x264 & ~x265 & ~x278 & ~x279 & ~x280 & ~x281 & ~x283 & ~x286 & ~x287 & ~x289 & ~x290 & ~x291 & ~x292 & ~x305 & ~x308 & ~x309 & ~x310 & ~x311 & ~x312 & ~x315 & ~x316 & ~x319 & ~x330 & ~x332 & ~x333 & ~x335 & ~x336 & ~x338 & ~x341 & ~x344 & ~x358 & ~x359 & ~x361 & ~x363 & ~x364 & ~x365 & ~x369 & ~x371 & ~x373 & ~x374 & ~x384 & ~x390 & ~x396 & ~x397 & ~x398 & ~x399 & ~x400 & ~x411 & ~x412 & ~x413 & ~x416 & ~x417 & ~x418 & ~x420 & ~x426 & ~x427 & ~x428 & ~x429 & ~x438 & ~x439 & ~x442 & ~x443 & ~x445 & ~x448 & ~x449 & ~x452 & ~x454 & ~x455 & ~x466 & ~x470 & ~x471 & ~x474 & ~x477 & ~x480 & ~x483 & ~x495 & ~x496 & ~x499 & ~x501 & ~x509 & ~x520 & ~x521 & ~x522 & ~x523 & ~x524 & ~x526 & ~x527 & ~x528 & ~x529 & ~x532 & ~x534 & ~x535 & ~x536 & ~x537 & ~x548 & ~x549 & ~x550 & ~x551 & ~x554 & ~x558 & ~x563 & ~x575 & ~x578 & ~x580 & ~x583 & ~x592 & ~x602 & ~x603 & ~x604 & ~x606 & ~x607 & ~x608 & ~x609 & ~x610 & ~x614 & ~x616 & ~x618 & ~x630 & ~x634 & ~x635 & ~x638 & ~x640 & ~x643 & ~x646 & ~x658 & ~x660 & ~x662 & ~x665 & ~x666 & ~x672 & ~x673 & ~x674 & ~x675 & ~x676 & ~x687 & ~x690 & ~x691 & ~x695 & ~x698 & ~x701 & ~x702 & ~x703 & ~x704 & ~x705 & ~x706 & ~x709 & ~x712 & ~x714 & ~x718 & ~x723 & ~x724 & ~x726 & ~x728 & ~x732 & ~x733 & ~x735 & ~x737 & ~x739 & ~x742 & ~x743 & ~x747 & ~x749 & ~x750 & ~x751 & ~x754 & ~x755 & ~x756 & ~x757 & ~x759 & ~x760 & ~x762 & ~x763 & ~x764 & ~x765 & ~x767 & ~x769 & ~x773 & ~x774 & ~x775 & ~x776 & ~x781 & ~x783;
assign c172 = ~x3 & ~x6 & ~x7 & ~x8 & ~x9 & ~x12 & ~x20 & ~x24 & ~x28 & ~x30 & ~x33 & ~x39 & ~x41 & ~x43 & ~x47 & ~x54 & ~x57 & ~x58 & ~x60 & ~x64 & ~x68 & ~x69 & ~x70 & ~x74 & ~x77 & ~x79 & ~x80 & ~x83 & ~x86 & ~x87 & ~x96 & ~x99 & ~x100 & ~x103 & ~x104 & ~x109 & ~x111 & ~x113 & ~x115 & ~x117 & ~x124 & ~x138 & ~x139 & ~x140 & ~x144 & ~x147 & ~x148 & ~x151 & ~x152 & ~x167 & ~x170 & ~x174 & ~x176 & ~x177 & ~x178 & ~x179 & ~x181 & ~x195 & ~x197 & ~x203 & ~x204 & ~x205 & ~x206 & ~x207 & ~x208 & ~x222 & ~x224 & ~x225 & ~x229 & ~x231 & ~x232 & ~x233 & ~x236 & ~x237 & ~x238 & ~x251 & ~x254 & ~x256 & ~x259 & ~x263 & ~x264 & ~x265 & ~x276 & ~x279 & ~x287 & ~x288 & ~x290 & ~x291 & ~x292 & ~x293 & ~x304 & ~x307 & ~x309 & ~x310 & ~x314 & ~x317 & ~x318 & ~x321 & ~x330 & ~x335 & ~x337 & ~x340 & ~x342 & ~x343 & ~x345 & ~x347 & ~x348 & ~x356 & ~x357 & ~x358 & ~x361 & ~x368 & ~x371 & ~x373 & ~x385 & ~x388 & ~x390 & ~x393 & ~x396 & ~x397 & ~x400 & ~x403 & ~x411 & ~x415 & ~x417 & ~x419 & ~x421 & ~x422 & ~x423 & ~x426 & ~x427 & ~x428 & ~x439 & ~x440 & ~x441 & ~x443 & ~x444 & ~x446 & ~x448 & ~x449 & ~x451 & ~x467 & ~x470 & ~x472 & ~x475 & ~x477 & ~x478 & ~x482 & ~x483 & ~x484 & ~x492 & ~x493 & ~x494 & ~x496 & ~x507 & ~x509 & ~x510 & ~x520 & ~x523 & ~x525 & ~x531 & ~x537 & ~x548 & ~x551 & ~x561 & ~x562 & ~x563 & ~x575 & ~x577 & ~x578 & ~x579 & ~x583 & ~x587 & ~x592 & ~x605 & ~x606 & ~x607 & ~x611 & ~x614 & ~x617 & ~x619 & ~x631 & ~x632 & ~x634 & ~x639 & ~x641 & ~x642 & ~x647 & ~x648 & ~x660 & ~x663 & ~x668 & ~x670 & ~x672 & ~x674 & ~x676 & ~x677 & ~x689 & ~x693 & ~x695 & ~x696 & ~x697 & ~x698 & ~x705 & ~x707 & ~x709 & ~x711 & ~x712 & ~x715 & ~x716 & ~x718 & ~x720 & ~x721 & ~x722 & ~x723 & ~x726 & ~x727 & ~x728 & ~x730 & ~x733 & ~x738 & ~x739 & ~x740 & ~x745 & ~x746 & ~x747 & ~x748 & ~x750 & ~x751 & ~x752 & ~x760 & ~x765 & ~x766 & ~x767 & ~x768 & ~x769 & ~x774 & ~x778 & ~x782;
assign c174 =  x269 &  x296 &  x324 &  x325 &  x350 &  x351 &  x405 &  x406 &  x460 &  x515 &  x516 &  x542 &  x543 &  x570 &  x597 & ~x2 & ~x6 & ~x10 & ~x13 & ~x14 & ~x17 & ~x23 & ~x25 & ~x26 & ~x27 & ~x28 & ~x29 & ~x32 & ~x33 & ~x34 & ~x35 & ~x36 & ~x38 & ~x44 & ~x45 & ~x46 & ~x47 & ~x55 & ~x56 & ~x59 & ~x61 & ~x62 & ~x63 & ~x65 & ~x67 & ~x68 & ~x69 & ~x70 & ~x72 & ~x73 & ~x75 & ~x77 & ~x79 & ~x80 & ~x84 & ~x88 & ~x89 & ~x91 & ~x93 & ~x98 & ~x99 & ~x100 & ~x101 & ~x108 & ~x110 & ~x117 & ~x118 & ~x123 & ~x124 & ~x125 & ~x127 & ~x128 & ~x135 & ~x139 & ~x142 & ~x143 & ~x146 & ~x148 & ~x152 & ~x153 & ~x154 & ~x155 & ~x165 & ~x167 & ~x170 & ~x171 & ~x172 & ~x175 & ~x177 & ~x178 & ~x180 & ~x194 & ~x197 & ~x198 & ~x202 & ~x207 & ~x210 & ~x222 & ~x225 & ~x226 & ~x231 & ~x233 & ~x235 & ~x236 & ~x237 & ~x248 & ~x249 & ~x250 & ~x256 & ~x258 & ~x260 & ~x261 & ~x263 & ~x264 & ~x265 & ~x277 & ~x281 & ~x284 & ~x287 & ~x288 & ~x291 & ~x305 & ~x306 & ~x309 & ~x311 & ~x316 & ~x318 & ~x335 & ~x336 & ~x337 & ~x341 & ~x342 & ~x344 & ~x357 & ~x359 & ~x360 & ~x361 & ~x366 & ~x368 & ~x369 & ~x370 & ~x373 & ~x384 & ~x385 & ~x388 & ~x389 & ~x392 & ~x393 & ~x395 & ~x411 & ~x412 & ~x414 & ~x416 & ~x417 & ~x418 & ~x419 & ~x420 & ~x424 & ~x425 & ~x426 & ~x427 & ~x438 & ~x439 & ~x440 & ~x444 & ~x448 & ~x451 & ~x452 & ~x455 & ~x468 & ~x473 & ~x475 & ~x478 & ~x482 & ~x493 & ~x494 & ~x498 & ~x502 & ~x503 & ~x506 & ~x507 & ~x508 & ~x525 & ~x526 & ~x530 & ~x531 & ~x532 & ~x536 & ~x537 & ~x550 & ~x552 & ~x558 & ~x559 & ~x560 & ~x561 & ~x562 & ~x575 & ~x578 & ~x579 & ~x580 & ~x582 & ~x585 & ~x591 & ~x602 & ~x604 & ~x605 & ~x609 & ~x610 & ~x615 & ~x620 & ~x633 & ~x634 & ~x635 & ~x636 & ~x642 & ~x643 & ~x646 & ~x647 & ~x648 & ~x658 & ~x659 & ~x671 & ~x676 & ~x685 & ~x686 & ~x688 & ~x691 & ~x692 & ~x694 & ~x698 & ~x700 & ~x702 & ~x705 & ~x706 & ~x707 & ~x711 & ~x714 & ~x724 & ~x725 & ~x726 & ~x727 & ~x728 & ~x731 & ~x734 & ~x735 & ~x737 & ~x738 & ~x739 & ~x740 & ~x744 & ~x745 & ~x746 & ~x749 & ~x750 & ~x753 & ~x754 & ~x760 & ~x761 & ~x762 & ~x770 & ~x781;
assign c176 =  x156 &  x267 &  x406 &  x490 &  x545 & ~x1 & ~x2 & ~x3 & ~x9 & ~x19 & ~x21 & ~x28 & ~x33 & ~x40 & ~x66 & ~x78 & ~x91 & ~x95 & ~x111 & ~x162 & ~x168 & ~x177 & ~x192 & ~x203 & ~x220 & ~x224 & ~x244 & ~x246 & ~x253 & ~x255 & ~x256 & ~x272 & ~x276 & ~x336 & ~x339 & ~x355 & ~x368 & ~x382 & ~x383 & ~x386 & ~x392 & ~x398 & ~x399 & ~x411 & ~x412 & ~x419 & ~x439 & ~x441 & ~x443 & ~x467 & ~x474 & ~x504 & ~x510 & ~x528 & ~x554 & ~x557 & ~x588 & ~x608 & ~x635 & ~x638 & ~x648 & ~x662 & ~x666 & ~x674 & ~x690 & ~x696 & ~x713 & ~x751 & ~x769;
assign c178 =  x322 & ~x3 & ~x89 & ~x129 & ~x132 & ~x134 & ~x188 & ~x212 & ~x220 & ~x231 & ~x250 & ~x325 & ~x382 & ~x411 & ~x442 & ~x455 & ~x478 & ~x505 & ~x513 & ~x531 & ~x539 & ~x561 & ~x616 & ~x669 & ~x708 & ~x720;
assign c180 =  x490 & ~x26 & ~x51 & ~x56 & ~x84 & ~x94 & ~x119 & ~x120 & ~x157 & ~x173 & ~x192 & ~x205 & ~x214 & ~x362 & ~x369 & ~x375 & ~x383 & ~x391 & ~x393 & ~x402 & ~x403 & ~x509 & ~x535 & ~x536 & ~x586 & ~x588 & ~x593 & ~x596 & ~x614 & ~x617 & ~x621 & ~x706 & ~x709 & ~x716 & ~x717 & ~x730 & ~x754 & ~x757 & ~x783;
assign c182 =  x216 &  x271 &  x325 &  x352 &  x380 &  x460 &  x487 &  x488 &  x515 &  x568 &  x595 & ~x182 & ~x235 & ~x236 & ~x262 & ~x292 & ~x400 & ~x438 & ~x573 & ~x574 & ~x578 & ~x629 & ~x633 & ~x635;
assign c184 =  x1;
assign c186 =  x295 &  x322 &  x407 &  x462 &  x517 & ~x2 & ~x3 & ~x4 & ~x6 & ~x7 & ~x12 & ~x15 & ~x16 & ~x20 & ~x23 & ~x26 & ~x29 & ~x37 & ~x38 & ~x40 & ~x45 & ~x51 & ~x55 & ~x58 & ~x59 & ~x79 & ~x80 & ~x82 & ~x85 & ~x90 & ~x91 & ~x98 & ~x99 & ~x102 & ~x107 & ~x118 & ~x120 & ~x123 & ~x132 & ~x135 & ~x144 & ~x145 & ~x160 & ~x165 & ~x175 & ~x178 & ~x189 & ~x191 & ~x195 & ~x196 & ~x197 & ~x202 & ~x203 & ~x205 & ~x226 & ~x229 & ~x230 & ~x245 & ~x246 & ~x251 & ~x252 & ~x255 & ~x259 & ~x261 & ~x272 & ~x273 & ~x288 & ~x289 & ~x304 & ~x306 & ~x313 & ~x315 & ~x329 & ~x331 & ~x334 & ~x337 & ~x342 & ~x361 & ~x367 & ~x382 & ~x390 & ~x395 & ~x410 & ~x411 & ~x413 & ~x415 & ~x416 & ~x421 & ~x422 & ~x440 & ~x445 & ~x447 & ~x450 & ~x451 & ~x452 & ~x455 & ~x456 & ~x467 & ~x469 & ~x470 & ~x473 & ~x482 & ~x483 & ~x484 & ~x494 & ~x495 & ~x523 & ~x524 & ~x527 & ~x530 & ~x532 & ~x540 & ~x551 & ~x553 & ~x564 & ~x582 & ~x587 & ~x589 & ~x591 & ~x592 & ~x593 & ~x609 & ~x611 & ~x613 & ~x619 & ~x620 & ~x621 & ~x622 & ~x640 & ~x644 & ~x646 & ~x651 & ~x669 & ~x670 & ~x672 & ~x674 & ~x677 & ~x678 & ~x679 & ~x689 & ~x692 & ~x693 & ~x694 & ~x695 & ~x696 & ~x697 & ~x699 & ~x704 & ~x706 & ~x707 & ~x708 & ~x720 & ~x728 & ~x731 & ~x732 & ~x738 & ~x743 & ~x748 & ~x750 & ~x753 & ~x763 & ~x764 & ~x765 & ~x766 & ~x770 & ~x772 & ~x773 & ~x775 & ~x778 & ~x781;
assign c188 =  x238 &  x323 &  x350 &  x378 &  x379 &  x407 &  x518 & ~x0 & ~x5 & ~x9 & ~x11 & ~x29 & ~x31 & ~x34 & ~x49 & ~x55 & ~x57 & ~x66 & ~x88 & ~x93 & ~x95 & ~x106 & ~x118 & ~x121 & ~x131 & ~x132 & ~x135 & ~x136 & ~x143 & ~x147 & ~x163 & ~x167 & ~x170 & ~x173 & ~x174 & ~x189 & ~x191 & ~x193 & ~x195 & ~x201 & ~x222 & ~x249 & ~x251 & ~x259 & ~x276 & ~x277 & ~x301 & ~x302 & ~x304 & ~x336 & ~x338 & ~x355 & ~x361 & ~x362 & ~x368 & ~x370 & ~x394 & ~x398 & ~x411 & ~x416 & ~x418 & ~x419 & ~x423 & ~x439 & ~x447 & ~x454 & ~x468 & ~x469 & ~x473 & ~x481 & ~x483 & ~x499 & ~x503 & ~x504 & ~x506 & ~x507 & ~x509 & ~x529 & ~x530 & ~x557 & ~x561 & ~x566 & ~x583 & ~x586 & ~x593 & ~x616 & ~x617 & ~x620 & ~x642 & ~x649 & ~x650 & ~x653 & ~x668 & ~x670 & ~x683 & ~x691 & ~x693 & ~x701 & ~x702 & ~x709 & ~x714 & ~x721 & ~x729 & ~x756 & ~x758 & ~x759 & ~x768 & ~x773 & ~x779;
assign c190 =  x590;
assign c192 =  x170;
assign c194 =  x141;
assign c196 =  x269 &  x489 & ~x40 & ~x48 & ~x52 & ~x68 & ~x75 & ~x76 & ~x80 & ~x94 & ~x98 & ~x106 & ~x123 & ~x124 & ~x136 & ~x147 & ~x149 & ~x150 & ~x151 & ~x162 & ~x172 & ~x179 & ~x181 & ~x191 & ~x195 & ~x203 & ~x232 & ~x234 & ~x235 & ~x236 & ~x237 & ~x246 & ~x247 & ~x259 & ~x263 & ~x264 & ~x265 & ~x278 & ~x288 & ~x291 & ~x293 & ~x302 & ~x311 & ~x314 & ~x317 & ~x318 & ~x319 & ~x328 & ~x339 & ~x341 & ~x345 & ~x346 & ~x348 & ~x355 & ~x357 & ~x372 & ~x373 & ~x390 & ~x400 & ~x402 & ~x403 & ~x440 & ~x445 & ~x466 & ~x475 & ~x479 & ~x482 & ~x484 & ~x492 & ~x493 & ~x495 & ~x496 & ~x519 & ~x520 & ~x521 & ~x523 & ~x530 & ~x538 & ~x540 & ~x547 & ~x548 & ~x550 & ~x566 & ~x577 & ~x579 & ~x594 & ~x595 & ~x607 & ~x613 & ~x614 & ~x632 & ~x644 & ~x658 & ~x659 & ~x665 & ~x676 & ~x685 & ~x692 & ~x704 & ~x736 & ~x759 & ~x769;
assign c198 =  x15;
assign c1102 =  x14;
assign c1104 =  x0;
assign c1106 =  x14 &  x113 &  x306;
assign c1108 =  x19;
assign c1110 =  x724;
assign c1112 =  x269 &  x296 &  x297 &  x324 &  x325 &  x326 &  x353 &  x378 &  x380 &  x406 &  x407 &  x461 &  x488 &  x515 &  x516 & ~x3 & ~x44 & ~x53 & ~x59 & ~x61 & ~x76 & ~x97 & ~x115 & ~x117 & ~x118 & ~x122 & ~x124 & ~x125 & ~x149 & ~x153 & ~x167 & ~x177 & ~x179 & ~x180 & ~x181 & ~x207 & ~x209 & ~x210 & ~x232 & ~x234 & ~x236 & ~x237 & ~x262 & ~x278 & ~x283 & ~x287 & ~x289 & ~x290 & ~x292 & ~x315 & ~x317 & ~x320 & ~x330 & ~x342 & ~x346 & ~x347 & ~x360 & ~x384 & ~x386 & ~x389 & ~x399 & ~x401 & ~x411 & ~x424 & ~x438 & ~x439 & ~x442 & ~x453 & ~x455 & ~x456 & ~x481 & ~x493 & ~x494 & ~x502 & ~x523 & ~x527 & ~x528 & ~x550 & ~x604 & ~x605 & ~x610 & ~x617 & ~x638 & ~x639 & ~x673 & ~x683 & ~x685 & ~x692 & ~x698 & ~x705 & ~x713 & ~x733 & ~x747 & ~x753 & ~x773 & ~x777;
assign c1114 =  x72 &  x127 & ~x487;
assign c1116 =  x6;
assign c1118 =  x156 &  x267 &  x296 &  x407 &  x463 &  x547 & ~x1 & ~x2 & ~x28 & ~x29 & ~x39 & ~x41 & ~x45 & ~x46 & ~x51 & ~x64 & ~x74 & ~x78 & ~x82 & ~x83 & ~x97 & ~x99 & ~x100 & ~x105 & ~x117 & ~x122 & ~x135 & ~x138 & ~x146 & ~x161 & ~x163 & ~x166 & ~x175 & ~x223 & ~x228 & ~x231 & ~x261 & ~x277 & ~x278 & ~x289 & ~x303 & ~x307 & ~x334 & ~x338 & ~x365 & ~x387 & ~x392 & ~x397 & ~x416 & ~x419 & ~x421 & ~x423 & ~x439 & ~x451 & ~x452 & ~x468 & ~x498 & ~x499 & ~x502 & ~x509 & ~x524 & ~x525 & ~x535 & ~x537 & ~x558 & ~x567 & ~x579 & ~x622 & ~x623 & ~x636 & ~x638 & ~x641 & ~x649 & ~x651 & ~x652 & ~x669 & ~x676 & ~x691 & ~x696 & ~x702 & ~x706 & ~x712 & ~x716 & ~x739 & ~x751 & ~x753 & ~x779 & ~x780;
assign c1120 =  x487 & ~x14 & ~x16 & ~x24 & ~x29 & ~x43 & ~x45 & ~x47 & ~x48 & ~x61 & ~x74 & ~x77 & ~x95 & ~x116 & ~x125 & ~x129 & ~x130 & ~x147 & ~x152 & ~x155 & ~x156 & ~x157 & ~x175 & ~x184 & ~x198 & ~x203 & ~x204 & ~x211 & ~x221 & ~x226 & ~x235 & ~x248 & ~x249 & ~x251 & ~x257 & ~x259 & ~x261 & ~x262 & ~x263 & ~x277 & ~x280 & ~x286 & ~x288 & ~x289 & ~x290 & ~x309 & ~x315 & ~x316 & ~x317 & ~x318 & ~x330 & ~x333 & ~x336 & ~x343 & ~x344 & ~x368 & ~x372 & ~x374 & ~x395 & ~x398 & ~x400 & ~x401 & ~x402 & ~x415 & ~x426 & ~x427 & ~x429 & ~x438 & ~x440 & ~x444 & ~x450 & ~x453 & ~x454 & ~x456 & ~x466 & ~x467 & ~x470 & ~x475 & ~x483 & ~x496 & ~x497 & ~x518 & ~x530 & ~x537 & ~x546 & ~x552 & ~x554 & ~x556 & ~x559 & ~x573 & ~x574 & ~x575 & ~x586 & ~x589 & ~x601 & ~x602 & ~x604 & ~x609 & ~x618 & ~x630 & ~x631 & ~x638 & ~x647 & ~x656 & ~x657 & ~x658 & ~x660 & ~x661 & ~x665 & ~x688 & ~x713 & ~x714 & ~x719 & ~x736 & ~x757 & ~x761 & ~x762 & ~x765 & ~x776 & ~x778;
assign c1122 =  x420;
assign c1124 =  x166;
assign c1126 =  x490 & ~x13 & ~x65 & ~x82 & ~x91 & ~x112 & ~x130 & ~x131 & ~x143 & ~x144 & ~x186 & ~x189 & ~x233 & ~x328 & ~x337 & ~x341 & ~x354 & ~x360 & ~x361 & ~x384 & ~x387 & ~x400 & ~x423 & ~x431 & ~x459 & ~x479 & ~x481 & ~x484 & ~x528 & ~x533 & ~x556 & ~x588 & ~x610 & ~x614 & ~x653 & ~x670 & ~x676 & ~x679 & ~x685 & ~x686 & ~x696 & ~x704 & ~x710 & ~x720 & ~x763 & ~x778 & ~x780;
assign c1128 =  x33;
assign c1130 =  x266 &  x294 &  x406 &  x490 & ~x14 & ~x29 & ~x43 & ~x49 & ~x72 & ~x88 & ~x91 & ~x116 & ~x120 & ~x144 & ~x167 & ~x185 & ~x200 & ~x204 & ~x231 & ~x241 & ~x245 & ~x251 & ~x273 & ~x314 & ~x335 & ~x411 & ~x428 & ~x451 & ~x454 & ~x485 & ~x486 & ~x509 & ~x530 & ~x587 & ~x589 & ~x622 & ~x647 & ~x650 & ~x652 & ~x674 & ~x690 & ~x695 & ~x729 & ~x754 & ~x755 & ~x758 & ~x778;
assign c1132 = ~x0 & ~x1 & ~x3 & ~x4 & ~x5 & ~x7 & ~x8 & ~x10 & ~x11 & ~x13 & ~x14 & ~x15 & ~x17 & ~x18 & ~x19 & ~x20 & ~x22 & ~x24 & ~x25 & ~x26 & ~x27 & ~x28 & ~x30 & ~x32 & ~x35 & ~x37 & ~x38 & ~x39 & ~x41 & ~x42 & ~x46 & ~x48 & ~x50 & ~x51 & ~x52 & ~x53 & ~x54 & ~x55 & ~x59 & ~x60 & ~x61 & ~x62 & ~x64 & ~x65 & ~x67 & ~x70 & ~x72 & ~x73 & ~x74 & ~x76 & ~x77 & ~x78 & ~x80 & ~x82 & ~x84 & ~x86 & ~x89 & ~x91 & ~x92 & ~x93 & ~x94 & ~x95 & ~x96 & ~x97 & ~x98 & ~x99 & ~x100 & ~x102 & ~x104 & ~x105 & ~x107 & ~x109 & ~x111 & ~x116 & ~x117 & ~x118 & ~x120 & ~x121 & ~x122 & ~x125 & ~x134 & ~x136 & ~x137 & ~x138 & ~x140 & ~x142 & ~x145 & ~x146 & ~x147 & ~x148 & ~x149 & ~x150 & ~x151 & ~x152 & ~x162 & ~x163 & ~x166 & ~x167 & ~x168 & ~x169 & ~x171 & ~x172 & ~x173 & ~x174 & ~x175 & ~x178 & ~x180 & ~x191 & ~x194 & ~x196 & ~x199 & ~x201 & ~x202 & ~x203 & ~x205 & ~x207 & ~x208 & ~x209 & ~x218 & ~x219 & ~x220 & ~x221 & ~x222 & ~x226 & ~x228 & ~x229 & ~x230 & ~x231 & ~x232 & ~x233 & ~x234 & ~x235 & ~x236 & ~x245 & ~x246 & ~x247 & ~x248 & ~x249 & ~x250 & ~x252 & ~x253 & ~x254 & ~x258 & ~x260 & ~x262 & ~x264 & ~x272 & ~x273 & ~x274 & ~x277 & ~x278 & ~x279 & ~x280 & ~x281 & ~x282 & ~x284 & ~x285 & ~x286 & ~x287 & ~x288 & ~x290 & ~x300 & ~x301 & ~x302 & ~x304 & ~x305 & ~x306 & ~x307 & ~x308 & ~x309 & ~x313 & ~x314 & ~x315 & ~x317 & ~x319 & ~x328 & ~x330 & ~x331 & ~x332 & ~x333 & ~x334 & ~x336 & ~x338 & ~x339 & ~x340 & ~x341 & ~x342 & ~x345 & ~x346 & ~x355 & ~x356 & ~x357 & ~x359 & ~x360 & ~x361 & ~x362 & ~x363 & ~x365 & ~x366 & ~x367 & ~x370 & ~x371 & ~x372 & ~x374 & ~x382 & ~x384 & ~x386 & ~x387 & ~x388 & ~x389 & ~x390 & ~x391 & ~x393 & ~x394 & ~x395 & ~x396 & ~x397 & ~x401 & ~x410 & ~x412 & ~x416 & ~x420 & ~x421 & ~x422 & ~x423 & ~x425 & ~x426 & ~x427 & ~x438 & ~x439 & ~x443 & ~x447 & ~x448 & ~x449 & ~x450 & ~x453 & ~x454 & ~x465 & ~x466 & ~x467 & ~x468 & ~x470 & ~x472 & ~x476 & ~x477 & ~x480 & ~x482 & ~x494 & ~x495 & ~x501 & ~x503 & ~x504 & ~x506 & ~x508 & ~x509 & ~x511 & ~x520 & ~x521 & ~x523 & ~x524 & ~x526 & ~x529 & ~x530 & ~x531 & ~x533 & ~x534 & ~x536 & ~x538 & ~x539 & ~x540 & ~x549 & ~x550 & ~x551 & ~x552 & ~x553 & ~x555 & ~x557 & ~x559 & ~x561 & ~x562 & ~x563 & ~x564 & ~x566 & ~x577 & ~x579 & ~x580 & ~x581 & ~x582 & ~x586 & ~x587 & ~x590 & ~x591 & ~x592 & ~x593 & ~x595 & ~x605 & ~x607 & ~x609 & ~x610 & ~x611 & ~x615 & ~x618 & ~x620 & ~x621 & ~x622 & ~x623 & ~x640 & ~x641 & ~x644 & ~x646 & ~x647 & ~x662 & ~x663 & ~x664 & ~x666 & ~x667 & ~x668 & ~x670 & ~x673 & ~x675 & ~x676 & ~x678 & ~x679 & ~x692 & ~x693 & ~x696 & ~x697 & ~x698 & ~x702 & ~x703 & ~x704 & ~x705 & ~x711 & ~x712 & ~x715 & ~x716 & ~x717 & ~x721 & ~x722 & ~x723 & ~x726 & ~x729 & ~x730 & ~x731 & ~x734 & ~x735 & ~x736 & ~x737 & ~x738 & ~x739 & ~x740 & ~x742 & ~x743 & ~x744 & ~x745 & ~x747 & ~x748 & ~x750 & ~x751 & ~x752 & ~x753 & ~x755 & ~x759 & ~x762 & ~x764 & ~x766 & ~x767 & ~x770 & ~x773 & ~x774 & ~x775 & ~x776 & ~x779 & ~x780 & ~x782;
assign c1134 =  x240 &  x267 &  x295 &  x296 &  x297 &  x380 &  x406 &  x407 &  x434 &  x435 &  x436 &  x462 &  x517 &  x518 &  x573 &  x600 &  x601 & ~x3 & ~x4 & ~x6 & ~x9 & ~x11 & ~x16 & ~x19 & ~x22 & ~x24 & ~x28 & ~x29 & ~x36 & ~x38 & ~x39 & ~x40 & ~x41 & ~x43 & ~x55 & ~x58 & ~x59 & ~x67 & ~x71 & ~x72 & ~x73 & ~x74 & ~x75 & ~x76 & ~x78 & ~x82 & ~x85 & ~x89 & ~x91 & ~x92 & ~x96 & ~x97 & ~x100 & ~x101 & ~x106 & ~x107 & ~x112 & ~x114 & ~x115 & ~x118 & ~x119 & ~x122 & ~x138 & ~x139 & ~x142 & ~x147 & ~x166 & ~x170 & ~x171 & ~x174 & ~x175 & ~x176 & ~x178 & ~x191 & ~x192 & ~x193 & ~x198 & ~x201 & ~x204 & ~x219 & ~x224 & ~x227 & ~x230 & ~x233 & ~x247 & ~x250 & ~x253 & ~x258 & ~x262 & ~x273 & ~x285 & ~x287 & ~x289 & ~x290 & ~x301 & ~x313 & ~x317 & ~x328 & ~x329 & ~x333 & ~x337 & ~x338 & ~x339 & ~x340 & ~x341 & ~x342 & ~x343 & ~x357 & ~x362 & ~x368 & ~x384 & ~x386 & ~x397 & ~x400 & ~x417 & ~x418 & ~x440 & ~x442 & ~x443 & ~x446 & ~x450 & ~x451 & ~x467 & ~x469 & ~x470 & ~x471 & ~x476 & ~x479 & ~x481 & ~x497 & ~x498 & ~x500 & ~x508 & ~x509 & ~x510 & ~x511 & ~x529 & ~x539 & ~x550 & ~x552 & ~x553 & ~x557 & ~x559 & ~x564 & ~x565 & ~x579 & ~x582 & ~x586 & ~x590 & ~x608 & ~x610 & ~x613 & ~x618 & ~x619 & ~x637 & ~x638 & ~x642 & ~x648 & ~x649 & ~x662 & ~x671 & ~x674 & ~x675 & ~x677 & ~x689 & ~x694 & ~x695 & ~x699 & ~x707 & ~x708 & ~x709 & ~x710 & ~x711 & ~x716 & ~x718 & ~x721 & ~x722 & ~x723 & ~x727 & ~x729 & ~x730 & ~x734 & ~x740 & ~x745 & ~x748 & ~x759 & ~x763 & ~x764 & ~x765 & ~x767 & ~x768 & ~x773 & ~x774 & ~x779;
assign c1136 =  x24;
assign c1138 =  x379 &  x406 & ~x1 & ~x3 & ~x6 & ~x7 & ~x8 & ~x15 & ~x16 & ~x17 & ~x18 & ~x19 & ~x20 & ~x21 & ~x22 & ~x24 & ~x25 & ~x28 & ~x29 & ~x30 & ~x31 & ~x32 & ~x34 & ~x36 & ~x38 & ~x39 & ~x40 & ~x41 & ~x45 & ~x46 & ~x47 & ~x49 & ~x50 & ~x51 & ~x52 & ~x55 & ~x56 & ~x57 & ~x60 & ~x61 & ~x62 & ~x66 & ~x68 & ~x69 & ~x70 & ~x71 & ~x72 & ~x73 & ~x74 & ~x75 & ~x76 & ~x77 & ~x79 & ~x81 & ~x82 & ~x83 & ~x85 & ~x86 & ~x87 & ~x88 & ~x89 & ~x91 & ~x92 & ~x93 & ~x96 & ~x99 & ~x100 & ~x101 & ~x104 & ~x106 & ~x107 & ~x108 & ~x111 & ~x114 & ~x115 & ~x116 & ~x117 & ~x118 & ~x119 & ~x120 & ~x125 & ~x126 & ~x127 & ~x128 & ~x136 & ~x137 & ~x138 & ~x139 & ~x140 & ~x141 & ~x142 & ~x143 & ~x145 & ~x147 & ~x148 & ~x150 & ~x153 & ~x154 & ~x155 & ~x166 & ~x168 & ~x170 & ~x171 & ~x172 & ~x173 & ~x174 & ~x176 & ~x181 & ~x182 & ~x183 & ~x192 & ~x193 & ~x196 & ~x197 & ~x198 & ~x199 & ~x200 & ~x204 & ~x205 & ~x206 & ~x209 & ~x211 & ~x219 & ~x220 & ~x222 & ~x224 & ~x225 & ~x228 & ~x229 & ~x231 & ~x232 & ~x233 & ~x234 & ~x248 & ~x249 & ~x250 & ~x254 & ~x255 & ~x256 & ~x258 & ~x259 & ~x261 & ~x274 & ~x275 & ~x276 & ~x278 & ~x279 & ~x283 & ~x284 & ~x286 & ~x287 & ~x288 & ~x289 & ~x290 & ~x301 & ~x304 & ~x305 & ~x306 & ~x307 & ~x313 & ~x314 & ~x315 & ~x316 & ~x317 & ~x318 & ~x330 & ~x333 & ~x336 & ~x337 & ~x338 & ~x339 & ~x341 & ~x342 & ~x343 & ~x344 & ~x345 & ~x346 & ~x347 & ~x357 & ~x358 & ~x364 & ~x365 & ~x366 & ~x367 & ~x369 & ~x371 & ~x372 & ~x373 & ~x375 & ~x385 & ~x386 & ~x387 & ~x388 & ~x389 & ~x391 & ~x393 & ~x399 & ~x400 & ~x401 & ~x413 & ~x416 & ~x417 & ~x420 & ~x421 & ~x423 & ~x424 & ~x425 & ~x428 & ~x429 & ~x438 & ~x440 & ~x441 & ~x443 & ~x444 & ~x447 & ~x448 & ~x454 & ~x455 & ~x466 & ~x470 & ~x471 & ~x473 & ~x475 & ~x476 & ~x477 & ~x478 & ~x480 & ~x495 & ~x496 & ~x497 & ~x499 & ~x500 & ~x501 & ~x502 & ~x503 & ~x505 & ~x506 & ~x507 & ~x508 & ~x509 & ~x510 & ~x520 & ~x522 & ~x525 & ~x526 & ~x527 & ~x528 & ~x529 & ~x530 & ~x533 & ~x534 & ~x535 & ~x536 & ~x537 & ~x552 & ~x553 & ~x555 & ~x557 & ~x558 & ~x559 & ~x560 & ~x561 & ~x562 & ~x563 & ~x579 & ~x580 & ~x581 & ~x583 & ~x584 & ~x585 & ~x586 & ~x587 & ~x588 & ~x589 & ~x592 & ~x608 & ~x610 & ~x611 & ~x612 & ~x613 & ~x614 & ~x615 & ~x616 & ~x618 & ~x619 & ~x620 & ~x629 & ~x635 & ~x636 & ~x637 & ~x639 & ~x640 & ~x641 & ~x642 & ~x643 & ~x644 & ~x646 & ~x647 & ~x657 & ~x658 & ~x665 & ~x666 & ~x667 & ~x668 & ~x669 & ~x670 & ~x672 & ~x676 & ~x684 & ~x686 & ~x688 & ~x690 & ~x694 & ~x695 & ~x696 & ~x698 & ~x699 & ~x701 & ~x702 & ~x705 & ~x706 & ~x707 & ~x710 & ~x711 & ~x712 & ~x714 & ~x715 & ~x716 & ~x717 & ~x718 & ~x724 & ~x725 & ~x727 & ~x730 & ~x734 & ~x735 & ~x736 & ~x737 & ~x738 & ~x739 & ~x740 & ~x741 & ~x742 & ~x743 & ~x744 & ~x745 & ~x748 & ~x749 & ~x750 & ~x751 & ~x752 & ~x754 & ~x755 & ~x758 & ~x759 & ~x761 & ~x764 & ~x767 & ~x768 & ~x769 & ~x770 & ~x771 & ~x773 & ~x775 & ~x776 & ~x777 & ~x778 & ~x780 & ~x781 & ~x782;
assign c1140 =  x154 &  x210 & ~x4 & ~x39 & ~x52 & ~x57 & ~x61 & ~x68 & ~x73 & ~x143 & ~x159 & ~x202 & ~x270 & ~x298 & ~x299 & ~x327 & ~x328 & ~x376 & ~x427 & ~x430 & ~x431 & ~x432 & ~x459 & ~x482 & ~x504 & ~x560 & ~x658 & ~x694 & ~x712 & ~x745;
assign c1142 =  x90;
assign c1146 =  x162 &  x622 & ~x157 & ~x265;
assign c1148 =  x294 &  x350 &  x406 &  x462 &  x518 & ~x7 & ~x8 & ~x17 & ~x30 & ~x35 & ~x36 & ~x72 & ~x76 & ~x80 & ~x89 & ~x116 & ~x117 & ~x118 & ~x129 & ~x130 & ~x141 & ~x146 & ~x167 & ~x195 & ~x216 & ~x220 & ~x227 & ~x242 & ~x246 & ~x249 & ~x257 & ~x270 & ~x302 & ~x304 & ~x309 & ~x311 & ~x331 & ~x358 & ~x363 & ~x364 & ~x365 & ~x366 & ~x388 & ~x392 & ~x394 & ~x398 & ~x420 & ~x421 & ~x439 & ~x447 & ~x478 & ~x510 & ~x529 & ~x552 & ~x558 & ~x560 & ~x565 & ~x566 & ~x569 & ~x625 & ~x641 & ~x645 & ~x651 & ~x680 & ~x694 & ~x708 & ~x709 & ~x729 & ~x755 & ~x769 & ~x777;
assign c1150 =  x22;
assign c1152 =  x505;
assign c1154 =  x767;
assign c1156 =  x238 & ~x28 & ~x42 & ~x47 & ~x49 & ~x57 & ~x71 & ~x75 & ~x104 & ~x120 & ~x132 & ~x134 & ~x146 & ~x158 & ~x160 & ~x170 & ~x176 & ~x189 & ~x245 & ~x277 & ~x279 & ~x280 & ~x282 & ~x298 & ~x299 & ~x307 & ~x314 & ~x328 & ~x344 & ~x356 & ~x362 & ~x367 & ~x368 & ~x387 & ~x388 & ~x389 & ~x397 & ~x410 & ~x414 & ~x416 & ~x417 & ~x420 & ~x438 & ~x447 & ~x451 & ~x452 & ~x466 & ~x479 & ~x487 & ~x497 & ~x504 & ~x507 & ~x511 & ~x533 & ~x540 & ~x554 & ~x555 & ~x557 & ~x587 & ~x591 & ~x639 & ~x646 & ~x663 & ~x674 & ~x698 & ~x699 & ~x713 & ~x716 & ~x721 & ~x725 & ~x741 & ~x752 & ~x756 & ~x758;
assign c1158 =  x212 &  x239 &  x240 &  x267 &  x268 &  x295 &  x323 &  x378 & ~x0 & ~x2 & ~x4 & ~x6 & ~x7 & ~x8 & ~x13 & ~x14 & ~x17 & ~x20 & ~x21 & ~x24 & ~x26 & ~x29 & ~x31 & ~x32 & ~x33 & ~x34 & ~x35 & ~x41 & ~x43 & ~x44 & ~x45 & ~x46 & ~x50 & ~x51 & ~x54 & ~x57 & ~x58 & ~x59 & ~x60 & ~x61 & ~x62 & ~x63 & ~x66 & ~x70 & ~x71 & ~x73 & ~x80 & ~x83 & ~x86 & ~x92 & ~x95 & ~x98 & ~x103 & ~x105 & ~x106 & ~x109 & ~x110 & ~x113 & ~x116 & ~x117 & ~x118 & ~x120 & ~x122 & ~x123 & ~x125 & ~x132 & ~x134 & ~x135 & ~x138 & ~x140 & ~x141 & ~x150 & ~x152 & ~x153 & ~x162 & ~x163 & ~x164 & ~x165 & ~x167 & ~x168 & ~x171 & ~x172 & ~x174 & ~x176 & ~x178 & ~x193 & ~x194 & ~x195 & ~x196 & ~x198 & ~x202 & ~x203 & ~x206 & ~x207 & ~x217 & ~x218 & ~x220 & ~x221 & ~x222 & ~x223 & ~x224 & ~x225 & ~x227 & ~x228 & ~x233 & ~x234 & ~x236 & ~x246 & ~x247 & ~x249 & ~x250 & ~x252 & ~x254 & ~x259 & ~x260 & ~x261 & ~x262 & ~x273 & ~x274 & ~x275 & ~x276 & ~x277 & ~x278 & ~x279 & ~x280 & ~x284 & ~x285 & ~x286 & ~x290 & ~x305 & ~x308 & ~x309 & ~x312 & ~x313 & ~x314 & ~x316 & ~x327 & ~x331 & ~x334 & ~x336 & ~x337 & ~x338 & ~x339 & ~x341 & ~x342 & ~x344 & ~x346 & ~x356 & ~x359 & ~x360 & ~x361 & ~x362 & ~x364 & ~x365 & ~x366 & ~x368 & ~x369 & ~x371 & ~x372 & ~x383 & ~x386 & ~x387 & ~x388 & ~x390 & ~x393 & ~x394 & ~x398 & ~x399 & ~x415 & ~x416 & ~x419 & ~x421 & ~x423 & ~x426 & ~x427 & ~x428 & ~x438 & ~x439 & ~x444 & ~x445 & ~x446 & ~x447 & ~x448 & ~x449 & ~x450 & ~x451 & ~x453 & ~x454 & ~x455 & ~x466 & ~x469 & ~x471 & ~x472 & ~x473 & ~x474 & ~x476 & ~x477 & ~x478 & ~x483 & ~x484 & ~x493 & ~x494 & ~x499 & ~x500 & ~x501 & ~x502 & ~x503 & ~x506 & ~x509 & ~x510 & ~x521 & ~x522 & ~x526 & ~x527 & ~x529 & ~x531 & ~x532 & ~x533 & ~x534 & ~x539 & ~x549 & ~x553 & ~x554 & ~x555 & ~x556 & ~x559 & ~x560 & ~x562 & ~x567 & ~x587 & ~x589 & ~x591 & ~x592 & ~x594 & ~x611 & ~x612 & ~x614 & ~x615 & ~x617 & ~x618 & ~x619 & ~x641 & ~x642 & ~x643 & ~x647 & ~x663 & ~x664 & ~x665 & ~x669 & ~x672 & ~x673 & ~x675 & ~x676 & ~x677 & ~x690 & ~x691 & ~x693 & ~x694 & ~x699 & ~x700 & ~x702 & ~x703 & ~x705 & ~x710 & ~x715 & ~x716 & ~x718 & ~x719 & ~x720 & ~x724 & ~x725 & ~x727 & ~x728 & ~x729 & ~x730 & ~x731 & ~x733 & ~x739 & ~x741 & ~x743 & ~x744 & ~x746 & ~x748 & ~x749 & ~x751 & ~x754 & ~x756 & ~x757 & ~x759 & ~x766 & ~x774 & ~x775 & ~x776 & ~x780;
assign c1160 = ~x4 & ~x8 & ~x9 & ~x10 & ~x15 & ~x19 & ~x20 & ~x24 & ~x36 & ~x40 & ~x43 & ~x46 & ~x52 & ~x57 & ~x59 & ~x60 & ~x62 & ~x69 & ~x74 & ~x81 & ~x82 & ~x84 & ~x85 & ~x90 & ~x93 & ~x94 & ~x97 & ~x105 & ~x107 & ~x110 & ~x112 & ~x116 & ~x118 & ~x119 & ~x120 & ~x123 & ~x127 & ~x139 & ~x146 & ~x150 & ~x168 & ~x169 & ~x171 & ~x176 & ~x178 & ~x190 & ~x192 & ~x194 & ~x195 & ~x205 & ~x219 & ~x221 & ~x225 & ~x226 & ~x227 & ~x229 & ~x232 & ~x233 & ~x234 & ~x247 & ~x249 & ~x251 & ~x252 & ~x254 & ~x256 & ~x258 & ~x262 & ~x276 & ~x277 & ~x281 & ~x288 & ~x290 & ~x292 & ~x309 & ~x312 & ~x319 & ~x328 & ~x330 & ~x331 & ~x332 & ~x334 & ~x335 & ~x385 & ~x386 & ~x388 & ~x393 & ~x395 & ~x398 & ~x410 & ~x416 & ~x442 & ~x445 & ~x449 & ~x452 & ~x465 & ~x466 & ~x469 & ~x470 & ~x471 & ~x472 & ~x479 & ~x480 & ~x494 & ~x500 & ~x501 & ~x503 & ~x506 & ~x509 & ~x540 & ~x549 & ~x550 & ~x553 & ~x554 & ~x559 & ~x563 & ~x577 & ~x584 & ~x585 & ~x588 & ~x589 & ~x592 & ~x594 & ~x597 & ~x608 & ~x612 & ~x615 & ~x616 & ~x621 & ~x623 & ~x624 & ~x625 & ~x636 & ~x638 & ~x641 & ~x643 & ~x644 & ~x646 & ~x647 & ~x648 & ~x654 & ~x663 & ~x669 & ~x679 & ~x690 & ~x691 & ~x704 & ~x708 & ~x710 & ~x717 & ~x720 & ~x721 & ~x722 & ~x726 & ~x732 & ~x734 & ~x737 & ~x742 & ~x747 & ~x754 & ~x755 & ~x759 & ~x768 & ~x769 & ~x775 & ~x783;
assign c1162 =  x46;
assign c1164 = ~x3 & ~x14 & ~x22 & ~x50 & ~x70 & ~x82 & ~x85 & ~x89 & ~x107 & ~x110 & ~x115 & ~x137 & ~x162 & ~x164 & ~x173 & ~x190 & ~x194 & ~x202 & ~x215 & ~x224 & ~x226 & ~x230 & ~x253 & ~x256 & ~x260 & ~x272 & ~x279 & ~x302 & ~x306 & ~x307 & ~x331 & ~x332 & ~x337 & ~x341 & ~x344 & ~x355 & ~x385 & ~x386 & ~x438 & ~x439 & ~x455 & ~x468 & ~x475 & ~x481 & ~x495 & ~x544 & ~x559 & ~x565 & ~x566 & ~x572 & ~x591 & ~x594 & ~x600 & ~x616 & ~x647 & ~x649 & ~x652 & ~x657 & ~x666 & ~x677 & ~x703 & ~x707 & ~x708 & ~x714 & ~x716 & ~x730 & ~x733 & ~x734 & ~x745 & ~x753 & ~x761 & ~x766 & ~x768 & ~x774;
assign c1166 = ~x6 & ~x12 & ~x15 & ~x19 & ~x21 & ~x28 & ~x33 & ~x37 & ~x38 & ~x50 & ~x54 & ~x55 & ~x56 & ~x67 & ~x70 & ~x80 & ~x83 & ~x85 & ~x92 & ~x93 & ~x98 & ~x99 & ~x104 & ~x107 & ~x111 & ~x112 & ~x130 & ~x132 & ~x137 & ~x140 & ~x144 & ~x151 & ~x160 & ~x167 & ~x169 & ~x173 & ~x189 & ~x191 & ~x192 & ~x218 & ~x219 & ~x227 & ~x228 & ~x230 & ~x231 & ~x233 & ~x234 & ~x235 & ~x254 & ~x256 & ~x260 & ~x274 & ~x280 & ~x282 & ~x288 & ~x301 & ~x302 & ~x305 & ~x307 & ~x309 & ~x344 & ~x353 & ~x354 & ~x362 & ~x364 & ~x368 & ~x371 & ~x383 & ~x392 & ~x399 & ~x421 & ~x423 & ~x443 & ~x444 & ~x445 & ~x451 & ~x452 & ~x453 & ~x465 & ~x474 & ~x498 & ~x502 & ~x508 & ~x510 & ~x521 & ~x522 & ~x527 & ~x530 & ~x535 & ~x539 & ~x540 & ~x557 & ~x559 & ~x562 & ~x565 & ~x566 & ~x592 & ~x614 & ~x617 & ~x646 & ~x647 & ~x665 & ~x670 & ~x674 & ~x681 & ~x695 & ~x698 & ~x701 & ~x703 & ~x718 & ~x720 & ~x729 & ~x735 & ~x737 & ~x739 & ~x745 & ~x748 & ~x749 & ~x757 & ~x762 & ~x766 & ~x767 & ~x770 & ~x776 & ~x783;
assign c1168 =  x297 &  x324 &  x406 &  x460 & ~x1 & ~x3 & ~x6 & ~x7 & ~x11 & ~x12 & ~x14 & ~x16 & ~x19 & ~x22 & ~x26 & ~x29 & ~x31 & ~x32 & ~x35 & ~x38 & ~x41 & ~x44 & ~x45 & ~x48 & ~x53 & ~x54 & ~x55 & ~x56 & ~x58 & ~x61 & ~x62 & ~x64 & ~x65 & ~x67 & ~x70 & ~x72 & ~x74 & ~x76 & ~x77 & ~x81 & ~x84 & ~x85 & ~x86 & ~x87 & ~x88 & ~x89 & ~x90 & ~x93 & ~x94 & ~x96 & ~x97 & ~x98 & ~x102 & ~x106 & ~x107 & ~x108 & ~x110 & ~x111 & ~x112 & ~x116 & ~x121 & ~x122 & ~x124 & ~x126 & ~x137 & ~x144 & ~x150 & ~x151 & ~x152 & ~x153 & ~x165 & ~x166 & ~x167 & ~x169 & ~x170 & ~x173 & ~x174 & ~x175 & ~x176 & ~x179 & ~x180 & ~x181 & ~x183 & ~x198 & ~x200 & ~x202 & ~x205 & ~x206 & ~x207 & ~x209 & ~x221 & ~x222 & ~x223 & ~x225 & ~x226 & ~x228 & ~x229 & ~x233 & ~x234 & ~x235 & ~x236 & ~x237 & ~x248 & ~x249 & ~x252 & ~x253 & ~x256 & ~x257 & ~x258 & ~x259 & ~x260 & ~x262 & ~x264 & ~x275 & ~x278 & ~x284 & ~x285 & ~x287 & ~x289 & ~x290 & ~x291 & ~x303 & ~x305 & ~x306 & ~x307 & ~x309 & ~x310 & ~x314 & ~x315 & ~x316 & ~x318 & ~x329 & ~x338 & ~x342 & ~x346 & ~x360 & ~x361 & ~x367 & ~x368 & ~x370 & ~x383 & ~x384 & ~x385 & ~x388 & ~x392 & ~x395 & ~x396 & ~x399 & ~x412 & ~x420 & ~x421 & ~x424 & ~x425 & ~x427 & ~x437 & ~x441 & ~x444 & ~x447 & ~x449 & ~x452 & ~x454 & ~x464 & ~x465 & ~x468 & ~x469 & ~x472 & ~x474 & ~x477 & ~x479 & ~x480 & ~x482 & ~x492 & ~x496 & ~x497 & ~x498 & ~x499 & ~x501 & ~x502 & ~x503 & ~x508 & ~x510 & ~x518 & ~x521 & ~x522 & ~x523 & ~x524 & ~x526 & ~x527 & ~x528 & ~x529 & ~x530 & ~x531 & ~x536 & ~x546 & ~x547 & ~x548 & ~x549 & ~x550 & ~x551 & ~x554 & ~x555 & ~x559 & ~x560 & ~x561 & ~x562 & ~x564 & ~x565 & ~x575 & ~x576 & ~x579 & ~x584 & ~x586 & ~x589 & ~x605 & ~x609 & ~x611 & ~x614 & ~x615 & ~x617 & ~x618 & ~x619 & ~x635 & ~x638 & ~x639 & ~x642 & ~x644 & ~x645 & ~x646 & ~x647 & ~x661 & ~x662 & ~x665 & ~x667 & ~x668 & ~x670 & ~x672 & ~x675 & ~x684 & ~x685 & ~x687 & ~x688 & ~x689 & ~x690 & ~x691 & ~x695 & ~x696 & ~x701 & ~x702 & ~x704 & ~x706 & ~x710 & ~x711 & ~x714 & ~x715 & ~x717 & ~x719 & ~x721 & ~x722 & ~x724 & ~x726 & ~x728 & ~x730 & ~x731 & ~x732 & ~x733 & ~x735 & ~x736 & ~x738 & ~x741 & ~x745 & ~x746 & ~x747 & ~x749 & ~x750 & ~x752 & ~x753 & ~x755 & ~x759 & ~x760 & ~x762 & ~x766 & ~x768 & ~x777 & ~x778 & ~x779;
assign c1170 =  x350 &  x520 &  x548 &  x576 &  x633 & ~x43 & ~x213 & ~x246 & ~x269 & ~x515;
assign c1172 =  x223;
assign c1174 =  x324 &  x351 &  x406 & ~x0 & ~x11 & ~x14 & ~x15 & ~x16 & ~x17 & ~x20 & ~x22 & ~x28 & ~x29 & ~x31 & ~x33 & ~x35 & ~x36 & ~x39 & ~x40 & ~x42 & ~x46 & ~x47 & ~x48 & ~x49 & ~x50 & ~x53 & ~x56 & ~x58 & ~x59 & ~x61 & ~x62 & ~x64 & ~x67 & ~x68 & ~x69 & ~x72 & ~x74 & ~x79 & ~x82 & ~x84 & ~x85 & ~x86 & ~x89 & ~x91 & ~x94 & ~x95 & ~x97 & ~x98 & ~x109 & ~x112 & ~x115 & ~x118 & ~x120 & ~x121 & ~x125 & ~x126 & ~x128 & ~x135 & ~x136 & ~x139 & ~x140 & ~x142 & ~x143 & ~x148 & ~x150 & ~x152 & ~x153 & ~x154 & ~x155 & ~x164 & ~x166 & ~x170 & ~x172 & ~x173 & ~x174 & ~x175 & ~x179 & ~x180 & ~x181 & ~x191 & ~x193 & ~x196 & ~x197 & ~x198 & ~x199 & ~x203 & ~x204 & ~x205 & ~x209 & ~x210 & ~x218 & ~x219 & ~x220 & ~x221 & ~x222 & ~x223 & ~x225 & ~x228 & ~x229 & ~x230 & ~x231 & ~x232 & ~x233 & ~x235 & ~x236 & ~x237 & ~x238 & ~x246 & ~x247 & ~x248 & ~x249 & ~x251 & ~x252 & ~x253 & ~x257 & ~x258 & ~x260 & ~x261 & ~x264 & ~x265 & ~x273 & ~x274 & ~x275 & ~x276 & ~x278 & ~x280 & ~x284 & ~x285 & ~x286 & ~x287 & ~x288 & ~x289 & ~x290 & ~x291 & ~x301 & ~x302 & ~x303 & ~x304 & ~x306 & ~x307 & ~x308 & ~x309 & ~x310 & ~x311 & ~x313 & ~x315 & ~x316 & ~x318 & ~x328 & ~x329 & ~x330 & ~x334 & ~x335 & ~x336 & ~x337 & ~x338 & ~x339 & ~x342 & ~x343 & ~x344 & ~x345 & ~x347 & ~x356 & ~x357 & ~x358 & ~x359 & ~x363 & ~x369 & ~x371 & ~x372 & ~x373 & ~x383 & ~x384 & ~x385 & ~x391 & ~x393 & ~x394 & ~x398 & ~x409 & ~x410 & ~x412 & ~x415 & ~x417 & ~x426 & ~x437 & ~x438 & ~x439 & ~x440 & ~x441 & ~x443 & ~x444 & ~x445 & ~x447 & ~x449 & ~x450 & ~x454 & ~x465 & ~x466 & ~x469 & ~x470 & ~x475 & ~x477 & ~x492 & ~x497 & ~x505 & ~x506 & ~x509 & ~x519 & ~x521 & ~x522 & ~x524 & ~x526 & ~x528 & ~x530 & ~x532 & ~x534 & ~x535 & ~x536 & ~x537 & ~x538 & ~x547 & ~x548 & ~x549 & ~x552 & ~x553 & ~x554 & ~x555 & ~x557 & ~x559 & ~x561 & ~x563 & ~x565 & ~x566 & ~x577 & ~x578 & ~x579 & ~x580 & ~x581 & ~x588 & ~x590 & ~x591 & ~x592 & ~x593 & ~x594 & ~x609 & ~x610 & ~x614 & ~x617 & ~x619 & ~x621 & ~x632 & ~x635 & ~x637 & ~x638 & ~x639 & ~x641 & ~x642 & ~x645 & ~x646 & ~x647 & ~x659 & ~x665 & ~x666 & ~x669 & ~x671 & ~x679 & ~x688 & ~x690 & ~x691 & ~x692 & ~x698 & ~x699 & ~x701 & ~x702 & ~x703 & ~x704 & ~x707 & ~x711 & ~x712 & ~x714 & ~x715 & ~x720 & ~x721 & ~x722 & ~x723 & ~x724 & ~x726 & ~x727 & ~x728 & ~x729 & ~x731 & ~x733 & ~x734 & ~x735 & ~x739 & ~x740 & ~x741 & ~x742 & ~x746 & ~x747 & ~x748 & ~x751 & ~x752 & ~x756 & ~x758 & ~x759 & ~x760 & ~x762 & ~x763 & ~x765 & ~x768 & ~x770 & ~x777 & ~x781 & ~x782;
assign c1176 =  x46;
assign c1178 = ~x3 & ~x8 & ~x9 & ~x12 & ~x13 & ~x14 & ~x28 & ~x30 & ~x37 & ~x39 & ~x40 & ~x42 & ~x43 & ~x53 & ~x55 & ~x59 & ~x60 & ~x65 & ~x74 & ~x77 & ~x94 & ~x115 & ~x122 & ~x123 & ~x137 & ~x145 & ~x162 & ~x163 & ~x169 & ~x171 & ~x173 & ~x175 & ~x191 & ~x192 & ~x194 & ~x199 & ~x201 & ~x203 & ~x206 & ~x219 & ~x231 & ~x232 & ~x233 & ~x234 & ~x245 & ~x246 & ~x249 & ~x250 & ~x253 & ~x271 & ~x273 & ~x284 & ~x300 & ~x304 & ~x314 & ~x318 & ~x320 & ~x326 & ~x327 & ~x334 & ~x338 & ~x341 & ~x343 & ~x345 & ~x348 & ~x354 & ~x358 & ~x365 & ~x381 & ~x394 & ~x400 & ~x409 & ~x414 & ~x416 & ~x417 & ~x419 & ~x421 & ~x423 & ~x425 & ~x429 & ~x430 & ~x436 & ~x438 & ~x439 & ~x454 & ~x456 & ~x458 & ~x464 & ~x465 & ~x466 & ~x467 & ~x468 & ~x471 & ~x473 & ~x474 & ~x485 & ~x492 & ~x495 & ~x505 & ~x506 & ~x507 & ~x508 & ~x536 & ~x565 & ~x585 & ~x588 & ~x590 & ~x610 & ~x639 & ~x641 & ~x663 & ~x668 & ~x675 & ~x685 & ~x687 & ~x688 & ~x689 & ~x692 & ~x694 & ~x695 & ~x698 & ~x709 & ~x716 & ~x721 & ~x723 & ~x727 & ~x742 & ~x749 & ~x751 & ~x752 & ~x756 & ~x759 & ~x764 & ~x773 & ~x778;
assign c1180 =  x376 &  x377 &  x404 &  x405 &  x432 &  x460 &  x487 &  x515 &  x543 & ~x0 & ~x17 & ~x35 & ~x49 & ~x52 & ~x58 & ~x68 & ~x94 & ~x97 & ~x109 & ~x123 & ~x125 & ~x141 & ~x143 & ~x146 & ~x147 & ~x148 & ~x152 & ~x177 & ~x179 & ~x180 & ~x205 & ~x206 & ~x234 & ~x236 & ~x247 & ~x261 & ~x263 & ~x275 & ~x276 & ~x285 & ~x291 & ~x317 & ~x318 & ~x336 & ~x343 & ~x345 & ~x363 & ~x371 & ~x373 & ~x374 & ~x396 & ~x400 & ~x425 & ~x455 & ~x465 & ~x468 & ~x491 & ~x493 & ~x500 & ~x504 & ~x519 & ~x529 & ~x532 & ~x546 & ~x547 & ~x554 & ~x561 & ~x565 & ~x574 & ~x575 & ~x576 & ~x585 & ~x602 & ~x603 & ~x615 & ~x632 & ~x640 & ~x658 & ~x685 & ~x726 & ~x729 & ~x739 & ~x744 & ~x754;
assign c1182 =  x678;
assign c1184 =  x29;
assign c1186 =  x728;
assign c1188 =  x80;
assign c1190 =  x267 & ~x1 & ~x2 & ~x12 & ~x30 & ~x35 & ~x49 & ~x51 & ~x52 & ~x56 & ~x57 & ~x65 & ~x68 & ~x74 & ~x88 & ~x89 & ~x92 & ~x106 & ~x108 & ~x112 & ~x117 & ~x118 & ~x122 & ~x141 & ~x144 & ~x148 & ~x152 & ~x160 & ~x163 & ~x166 & ~x178 & ~x191 & ~x192 & ~x206 & ~x217 & ~x220 & ~x221 & ~x224 & ~x233 & ~x259 & ~x263 & ~x271 & ~x286 & ~x305 & ~x311 & ~x315 & ~x317 & ~x336 & ~x347 & ~x367 & ~x370 & ~x390 & ~x393 & ~x399 & ~x410 & ~x411 & ~x412 & ~x419 & ~x427 & ~x438 & ~x442 & ~x445 & ~x449 & ~x471 & ~x472 & ~x478 & ~x508 & ~x528 & ~x529 & ~x531 & ~x553 & ~x566 & ~x569 & ~x584 & ~x592 & ~x595 & ~x614 & ~x615 & ~x617 & ~x648 & ~x650 & ~x670 & ~x675 & ~x677 & ~x680 & ~x698 & ~x707 & ~x717 & ~x722 & ~x724 & ~x725 & ~x741 & ~x744 & ~x751 & ~x758 & ~x767;
assign c1192 =  x15;
assign c1194 =  x293 &  x321 &  x349 &  x406 & ~x14 & ~x19 & ~x22 & ~x69 & ~x77 & ~x80 & ~x86 & ~x91 & ~x95 & ~x103 & ~x190 & ~x201 & ~x221 & ~x249 & ~x284 & ~x327 & ~x329 & ~x333 & ~x361 & ~x370 & ~x371 & ~x412 & ~x421 & ~x425 & ~x438 & ~x441 & ~x481 & ~x487 & ~x515 & ~x561 & ~x585 & ~x615 & ~x622 & ~x652 & ~x653 & ~x655 & ~x657 & ~x673 & ~x678 & ~x702 & ~x707 & ~x714 & ~x733 & ~x747 & ~x749 & ~x754 & ~x764;
assign c1196 =  x40;
assign c1198 =  x491 &  x547 & ~x3 & ~x8 & ~x28 & ~x29 & ~x32 & ~x37 & ~x42 & ~x47 & ~x50 & ~x54 & ~x55 & ~x65 & ~x81 & ~x94 & ~x111 & ~x112 & ~x114 & ~x118 & ~x140 & ~x166 & ~x171 & ~x187 & ~x190 & ~x191 & ~x193 & ~x202 & ~x226 & ~x242 & ~x244 & ~x246 & ~x247 & ~x254 & ~x258 & ~x269 & ~x276 & ~x300 & ~x311 & ~x326 & ~x338 & ~x339 & ~x341 & ~x361 & ~x363 & ~x383 & ~x386 & ~x392 & ~x395 & ~x411 & ~x414 & ~x428 & ~x437 & ~x449 & ~x485 & ~x500 & ~x515 & ~x530 & ~x565 & ~x583 & ~x591 & ~x620 & ~x646 & ~x649 & ~x651 & ~x652 & ~x672 & ~x685 & ~x694 & ~x709 & ~x717 & ~x723 & ~x732 & ~x733 & ~x734 & ~x741 & ~x746 & ~x748 & ~x752 & ~x767 & ~x769 & ~x772 & ~x779;
assign c1200 =  x154 &  x295 & ~x4 & ~x13 & ~x47 & ~x86 & ~x89 & ~x117 & ~x120 & ~x121 & ~x137 & ~x146 & ~x214 & ~x225 & ~x242 & ~x247 & ~x273 & ~x300 & ~x329 & ~x338 & ~x360 & ~x397 & ~x425 & ~x429 & ~x430 & ~x451 & ~x453 & ~x460 & ~x473 & ~x478 & ~x486 & ~x500 & ~x507 & ~x533 & ~x534 & ~x685 & ~x687 & ~x688 & ~x706 & ~x742 & ~x771 & ~x772 & ~x782;
assign c1202 =  x433 &  x460 & ~x3 & ~x8 & ~x15 & ~x18 & ~x19 & ~x35 & ~x38 & ~x39 & ~x40 & ~x47 & ~x52 & ~x55 & ~x57 & ~x58 & ~x59 & ~x71 & ~x72 & ~x76 & ~x78 & ~x82 & ~x91 & ~x93 & ~x94 & ~x95 & ~x98 & ~x102 & ~x114 & ~x122 & ~x124 & ~x139 & ~x141 & ~x143 & ~x148 & ~x152 & ~x165 & ~x168 & ~x173 & ~x176 & ~x177 & ~x179 & ~x181 & ~x194 & ~x200 & ~x208 & ~x223 & ~x227 & ~x230 & ~x231 & ~x232 & ~x235 & ~x247 & ~x259 & ~x261 & ~x262 & ~x274 & ~x275 & ~x277 & ~x284 & ~x287 & ~x288 & ~x291 & ~x292 & ~x303 & ~x313 & ~x314 & ~x317 & ~x332 & ~x333 & ~x338 & ~x345 & ~x359 & ~x367 & ~x372 & ~x374 & ~x375 & ~x398 & ~x402 & ~x409 & ~x410 & ~x414 & ~x415 & ~x416 & ~x421 & ~x423 & ~x424 & ~x426 & ~x428 & ~x437 & ~x442 & ~x443 & ~x454 & ~x456 & ~x463 & ~x464 & ~x467 & ~x479 & ~x481 & ~x483 & ~x493 & ~x504 & ~x510 & ~x521 & ~x529 & ~x535 & ~x547 & ~x552 & ~x554 & ~x559 & ~x562 & ~x563 & ~x574 & ~x575 & ~x580 & ~x585 & ~x586 & ~x587 & ~x588 & ~x603 & ~x609 & ~x613 & ~x614 & ~x617 & ~x618 & ~x633 & ~x638 & ~x639 & ~x645 & ~x648 & ~x658 & ~x659 & ~x661 & ~x662 & ~x663 & ~x666 & ~x669 & ~x671 & ~x672 & ~x673 & ~x676 & ~x678 & ~x679 & ~x689 & ~x691 & ~x717 & ~x719 & ~x720 & ~x724 & ~x725 & ~x726 & ~x729 & ~x730 & ~x732 & ~x735 & ~x740 & ~x751 & ~x754 & ~x756 & ~x759 & ~x760 & ~x769 & ~x771 & ~x773 & ~x777 & ~x779;
assign c1204 =  x614;
assign c1206 =  x769;
assign c1208 =  x294 &  x322 & ~x8 & ~x28 & ~x32 & ~x33 & ~x39 & ~x48 & ~x52 & ~x53 & ~x62 & ~x66 & ~x69 & ~x76 & ~x83 & ~x85 & ~x86 & ~x88 & ~x95 & ~x104 & ~x105 & ~x108 & ~x117 & ~x120 & ~x141 & ~x160 & ~x164 & ~x194 & ~x202 & ~x204 & ~x214 & ~x217 & ~x219 & ~x241 & ~x243 & ~x246 & ~x258 & ~x271 & ~x332 & ~x333 & ~x353 & ~x357 & ~x364 & ~x371 & ~x381 & ~x386 & ~x390 & ~x398 & ~x403 & ~x413 & ~x428 & ~x454 & ~x456 & ~x458 & ~x471 & ~x474 & ~x486 & ~x507 & ~x512 & ~x535 & ~x557 & ~x588 & ~x594 & ~x610 & ~x621 & ~x623 & ~x638 & ~x649 & ~x650 & ~x669 & ~x674 & ~x677 & ~x680 & ~x689 & ~x690 & ~x696 & ~x698 & ~x706 & ~x712 & ~x719 & ~x725 & ~x730 & ~x733 & ~x734 & ~x739 & ~x761 & ~x764 & ~x769 & ~x776 & ~x780 & ~x782;
assign c1210 =  x351 &  x433 &  x460 &  x487 &  x542 &  x568 &  x569 & ~x125 & ~x151 & ~x154 & ~x178 & ~x180 & ~x230 & ~x231 & ~x234 & ~x237 & ~x263 & ~x265 & ~x287 & ~x318 & ~x319 & ~x330 & ~x346 & ~x363 & ~x372 & ~x373 & ~x374 & ~x384 & ~x399 & ~x438 & ~x482 & ~x491 & ~x492 & ~x509 & ~x519 & ~x531 & ~x546 & ~x547 & ~x552 & ~x574 & ~x575 & ~x576 & ~x585 & ~x601 & ~x602 & ~x628 & ~x629 & ~x630 & ~x656;
assign c1212 =  x518 &  x519 &  x547 &  x604 & ~x30 & ~x44 & ~x56 & ~x65 & ~x67 & ~x72 & ~x86 & ~x88 & ~x94 & ~x100 & ~x116 & ~x137 & ~x140 & ~x162 & ~x191 & ~x222 & ~x223 & ~x230 & ~x231 & ~x245 & ~x299 & ~x300 & ~x305 & ~x315 & ~x316 & ~x326 & ~x328 & ~x343 & ~x354 & ~x355 & ~x356 & ~x362 & ~x366 & ~x392 & ~x413 & ~x416 & ~x425 & ~x452 & ~x467 & ~x472 & ~x473 & ~x474 & ~x497 & ~x499 & ~x529 & ~x557 & ~x584 & ~x591 & ~x592 & ~x595 & ~x599 & ~x610 & ~x615 & ~x667 & ~x671 & ~x678 & ~x679 & ~x685 & ~x692 & ~x695 & ~x710 & ~x716 & ~x717 & ~x718 & ~x723 & ~x736 & ~x737 & ~x738 & ~x741 & ~x744 & ~x745 & ~x754 & ~x755 & ~x758 & ~x761 & ~x775 & ~x781 & ~x782 & ~x783;
assign c1214 =  x186 &  x212 &  x241 &  x242 &  x268 &  x269 &  x296 &  x297 &  x324 &  x325 &  x379 &  x408 &  x434 &  x435 &  x462 &  x517 & ~x2 & ~x3 & ~x5 & ~x18 & ~x20 & ~x24 & ~x25 & ~x27 & ~x29 & ~x30 & ~x37 & ~x39 & ~x54 & ~x58 & ~x59 & ~x75 & ~x76 & ~x77 & ~x79 & ~x83 & ~x87 & ~x89 & ~x91 & ~x93 & ~x94 & ~x97 & ~x98 & ~x99 & ~x100 & ~x102 & ~x103 & ~x106 & ~x114 & ~x119 & ~x122 & ~x123 & ~x135 & ~x136 & ~x143 & ~x148 & ~x149 & ~x152 & ~x165 & ~x167 & ~x168 & ~x169 & ~x171 & ~x172 & ~x175 & ~x177 & ~x178 & ~x193 & ~x194 & ~x197 & ~x198 & ~x199 & ~x200 & ~x201 & ~x202 & ~x207 & ~x223 & ~x226 & ~x231 & ~x232 & ~x233 & ~x235 & ~x246 & ~x249 & ~x250 & ~x253 & ~x254 & ~x260 & ~x261 & ~x275 & ~x280 & ~x284 & ~x290 & ~x301 & ~x311 & ~x312 & ~x328 & ~x329 & ~x330 & ~x332 & ~x338 & ~x341 & ~x342 & ~x356 & ~x358 & ~x363 & ~x365 & ~x368 & ~x373 & ~x384 & ~x388 & ~x390 & ~x393 & ~x399 & ~x412 & ~x419 & ~x421 & ~x426 & ~x439 & ~x442 & ~x443 & ~x444 & ~x445 & ~x450 & ~x451 & ~x453 & ~x455 & ~x466 & ~x467 & ~x468 & ~x469 & ~x472 & ~x476 & ~x479 & ~x481 & ~x494 & ~x498 & ~x500 & ~x505 & ~x508 & ~x525 & ~x526 & ~x530 & ~x537 & ~x550 & ~x555 & ~x556 & ~x558 & ~x562 & ~x563 & ~x565 & ~x582 & ~x584 & ~x585 & ~x586 & ~x588 & ~x589 & ~x591 & ~x592 & ~x608 & ~x611 & ~x612 & ~x613 & ~x615 & ~x618 & ~x620 & ~x621 & ~x633 & ~x634 & ~x636 & ~x637 & ~x661 & ~x662 & ~x663 & ~x664 & ~x665 & ~x668 & ~x671 & ~x672 & ~x673 & ~x674 & ~x675 & ~x689 & ~x690 & ~x692 & ~x696 & ~x697 & ~x698 & ~x699 & ~x703 & ~x704 & ~x710 & ~x711 & ~x715 & ~x717 & ~x720 & ~x725 & ~x729 & ~x731 & ~x734 & ~x735 & ~x737 & ~x739 & ~x741 & ~x749 & ~x753 & ~x756 & ~x758 & ~x759 & ~x763 & ~x766 & ~x767 & ~x768 & ~x778 & ~x781 & ~x782 & ~x783;
assign c1218 =  x253 &  x703;
assign c1220 = ~x1 & ~x8 & ~x18 & ~x21 & ~x23 & ~x24 & ~x26 & ~x27 & ~x29 & ~x31 & ~x40 & ~x46 & ~x48 & ~x64 & ~x66 & ~x76 & ~x80 & ~x82 & ~x86 & ~x88 & ~x89 & ~x105 & ~x107 & ~x109 & ~x111 & ~x112 & ~x121 & ~x135 & ~x161 & ~x168 & ~x170 & ~x171 & ~x172 & ~x178 & ~x190 & ~x191 & ~x192 & ~x196 & ~x199 & ~x200 & ~x201 & ~x202 & ~x204 & ~x206 & ~x218 & ~x221 & ~x231 & ~x245 & ~x248 & ~x254 & ~x255 & ~x256 & ~x258 & ~x260 & ~x263 & ~x272 & ~x278 & ~x280 & ~x281 & ~x284 & ~x288 & ~x290 & ~x305 & ~x307 & ~x313 & ~x314 & ~x317 & ~x327 & ~x334 & ~x335 & ~x337 & ~x339 & ~x340 & ~x343 & ~x345 & ~x354 & ~x358 & ~x359 & ~x369 & ~x372 & ~x383 & ~x394 & ~x398 & ~x411 & ~x413 & ~x415 & ~x423 & ~x425 & ~x439 & ~x440 & ~x443 & ~x450 & ~x453 & ~x465 & ~x467 & ~x468 & ~x470 & ~x473 & ~x475 & ~x482 & ~x483 & ~x492 & ~x493 & ~x506 & ~x512 & ~x527 & ~x530 & ~x531 & ~x534 & ~x537 & ~x540 & ~x562 & ~x569 & ~x589 & ~x592 & ~x593 & ~x606 & ~x613 & ~x614 & ~x616 & ~x622 & ~x634 & ~x635 & ~x640 & ~x643 & ~x652 & ~x662 & ~x667 & ~x668 & ~x672 & ~x673 & ~x677 & ~x680 & ~x691 & ~x694 & ~x696 & ~x703 & ~x705 & ~x718 & ~x721 & ~x724 & ~x726 & ~x727 & ~x728 & ~x731 & ~x732 & ~x736 & ~x743 & ~x745 & ~x749 & ~x757 & ~x762 & ~x764 & ~x768 & ~x769 & ~x776 & ~x779 & ~x783;
assign c1222 =  x489 &  x543 &  x544 &  x571 &  x600 & ~x18 & ~x19 & ~x23 & ~x40 & ~x41 & ~x52 & ~x61 & ~x64 & ~x75 & ~x81 & ~x83 & ~x90 & ~x105 & ~x117 & ~x120 & ~x126 & ~x134 & ~x146 & ~x148 & ~x151 & ~x152 & ~x164 & ~x175 & ~x189 & ~x195 & ~x198 & ~x203 & ~x206 & ~x219 & ~x220 & ~x221 & ~x225 & ~x227 & ~x233 & ~x235 & ~x246 & ~x251 & ~x273 & ~x276 & ~x280 & ~x282 & ~x285 & ~x304 & ~x313 & ~x316 & ~x333 & ~x338 & ~x342 & ~x346 & ~x347 & ~x355 & ~x372 & ~x384 & ~x390 & ~x399 & ~x401 & ~x427 & ~x439 & ~x442 & ~x443 & ~x444 & ~x448 & ~x457 & ~x469 & ~x474 & ~x475 & ~x482 & ~x483 & ~x509 & ~x512 & ~x525 & ~x538 & ~x539 & ~x548 & ~x550 & ~x554 & ~x565 & ~x567 & ~x580 & ~x581 & ~x583 & ~x584 & ~x595 & ~x622 & ~x640 & ~x643 & ~x659 & ~x662 & ~x687 & ~x693 & ~x700 & ~x707 & ~x711 & ~x712 & ~x714 & ~x718 & ~x725 & ~x731 & ~x734 & ~x738 & ~x742 & ~x754 & ~x755 & ~x761 & ~x765 & ~x766 & ~x767 & ~x775 & ~x776;
assign c1224 =  x729;
assign c1226 =  x186 &  x241 &  x268 &  x269 &  x296 &  x297 &  x324 &  x352 &  x380 &  x406 &  x407 &  x408 & ~x1 & ~x2 & ~x3 & ~x4 & ~x8 & ~x12 & ~x16 & ~x20 & ~x21 & ~x24 & ~x26 & ~x28 & ~x29 & ~x30 & ~x33 & ~x34 & ~x35 & ~x37 & ~x40 & ~x42 & ~x45 & ~x47 & ~x48 & ~x49 & ~x50 & ~x51 & ~x53 & ~x54 & ~x56 & ~x59 & ~x60 & ~x64 & ~x66 & ~x67 & ~x69 & ~x71 & ~x72 & ~x73 & ~x75 & ~x76 & ~x77 & ~x78 & ~x80 & ~x81 & ~x83 & ~x86 & ~x88 & ~x90 & ~x91 & ~x92 & ~x93 & ~x94 & ~x95 & ~x97 & ~x99 & ~x104 & ~x108 & ~x109 & ~x111 & ~x115 & ~x118 & ~x120 & ~x121 & ~x122 & ~x135 & ~x137 & ~x138 & ~x139 & ~x141 & ~x142 & ~x145 & ~x151 & ~x152 & ~x153 & ~x154 & ~x155 & ~x163 & ~x167 & ~x168 & ~x170 & ~x172 & ~x175 & ~x177 & ~x178 & ~x179 & ~x181 & ~x190 & ~x192 & ~x194 & ~x195 & ~x201 & ~x202 & ~x204 & ~x205 & ~x207 & ~x209 & ~x210 & ~x219 & ~x221 & ~x222 & ~x224 & ~x228 & ~x230 & ~x231 & ~x232 & ~x235 & ~x236 & ~x251 & ~x252 & ~x255 & ~x257 & ~x258 & ~x260 & ~x261 & ~x262 & ~x263 & ~x265 & ~x274 & ~x278 & ~x281 & ~x283 & ~x286 & ~x289 & ~x290 & ~x302 & ~x303 & ~x307 & ~x310 & ~x311 & ~x312 & ~x318 & ~x328 & ~x330 & ~x331 & ~x332 & ~x334 & ~x336 & ~x338 & ~x341 & ~x343 & ~x356 & ~x357 & ~x359 & ~x360 & ~x361 & ~x363 & ~x364 & ~x369 & ~x372 & ~x384 & ~x385 & ~x386 & ~x387 & ~x388 & ~x390 & ~x391 & ~x395 & ~x398 & ~x400 & ~x411 & ~x413 & ~x414 & ~x417 & ~x418 & ~x421 & ~x422 & ~x426 & ~x438 & ~x439 & ~x440 & ~x444 & ~x445 & ~x446 & ~x447 & ~x448 & ~x450 & ~x451 & ~x452 & ~x453 & ~x465 & ~x466 & ~x467 & ~x470 & ~x477 & ~x478 & ~x482 & ~x483 & ~x493 & ~x494 & ~x497 & ~x499 & ~x500 & ~x502 & ~x503 & ~x509 & ~x510 & ~x522 & ~x523 & ~x524 & ~x526 & ~x527 & ~x528 & ~x531 & ~x536 & ~x550 & ~x552 & ~x554 & ~x555 & ~x556 & ~x557 & ~x558 & ~x560 & ~x562 & ~x563 & ~x579 & ~x580 & ~x581 & ~x582 & ~x584 & ~x585 & ~x586 & ~x592 & ~x605 & ~x606 & ~x607 & ~x609 & ~x612 & ~x615 & ~x617 & ~x618 & ~x619 & ~x620 & ~x621 & ~x635 & ~x636 & ~x637 & ~x639 & ~x643 & ~x644 & ~x645 & ~x648 & ~x661 & ~x662 & ~x663 & ~x668 & ~x670 & ~x671 & ~x675 & ~x689 & ~x691 & ~x693 & ~x696 & ~x697 & ~x698 & ~x699 & ~x703 & ~x705 & ~x708 & ~x711 & ~x715 & ~x722 & ~x723 & ~x724 & ~x725 & ~x729 & ~x730 & ~x731 & ~x732 & ~x733 & ~x735 & ~x736 & ~x738 & ~x739 & ~x740 & ~x741 & ~x742 & ~x745 & ~x746 & ~x747 & ~x750 & ~x751 & ~x753 & ~x756 & ~x758 & ~x759 & ~x760 & ~x761 & ~x764 & ~x765 & ~x771 & ~x772 & ~x773 & ~x775 & ~x781 & ~x783;
assign c1228 =  x266 &  x350 &  x378 &  x517 & ~x1 & ~x4 & ~x5 & ~x11 & ~x15 & ~x18 & ~x26 & ~x40 & ~x41 & ~x63 & ~x70 & ~x77 & ~x81 & ~x91 & ~x96 & ~x98 & ~x99 & ~x105 & ~x107 & ~x113 & ~x118 & ~x120 & ~x122 & ~x131 & ~x134 & ~x138 & ~x144 & ~x148 & ~x160 & ~x169 & ~x173 & ~x198 & ~x201 & ~x203 & ~x216 & ~x219 & ~x227 & ~x229 & ~x230 & ~x246 & ~x251 & ~x252 & ~x276 & ~x287 & ~x316 & ~x330 & ~x337 & ~x342 & ~x354 & ~x392 & ~x394 & ~x401 & ~x416 & ~x418 & ~x420 & ~x428 & ~x443 & ~x447 & ~x470 & ~x472 & ~x504 & ~x506 & ~x507 & ~x509 & ~x511 & ~x526 & ~x533 & ~x537 & ~x540 & ~x554 & ~x563 & ~x583 & ~x587 & ~x589 & ~x619 & ~x637 & ~x663 & ~x664 & ~x669 & ~x670 & ~x672 & ~x693 & ~x696 & ~x698 & ~x708 & ~x711 & ~x716 & ~x723 & ~x739 & ~x741 & ~x750 & ~x751 & ~x754 & ~x769 & ~x778 & ~x783;
assign c1230 =  x53;
assign c1232 =  x61;
assign c1234 =  x112;
assign c1236 =  x675;
assign c1238 =  x336;
assign c1240 =  x196;
assign c1242 = ~x0 & ~x2 & ~x3 & ~x4 & ~x5 & ~x6 & ~x7 & ~x9 & ~x11 & ~x13 & ~x14 & ~x15 & ~x17 & ~x18 & ~x19 & ~x20 & ~x21 & ~x23 & ~x27 & ~x28 & ~x31 & ~x32 & ~x34 & ~x37 & ~x38 & ~x39 & ~x41 & ~x42 & ~x44 & ~x47 & ~x48 & ~x50 & ~x51 & ~x56 & ~x58 & ~x62 & ~x64 & ~x65 & ~x67 & ~x68 & ~x69 & ~x72 & ~x73 & ~x76 & ~x77 & ~x79 & ~x80 & ~x81 & ~x83 & ~x84 & ~x86 & ~x92 & ~x94 & ~x95 & ~x96 & ~x98 & ~x99 & ~x100 & ~x106 & ~x109 & ~x110 & ~x111 & ~x112 & ~x113 & ~x114 & ~x115 & ~x118 & ~x120 & ~x121 & ~x122 & ~x123 & ~x124 & ~x136 & ~x140 & ~x143 & ~x144 & ~x149 & ~x150 & ~x151 & ~x152 & ~x153 & ~x165 & ~x167 & ~x173 & ~x174 & ~x175 & ~x176 & ~x177 & ~x178 & ~x179 & ~x180 & ~x181 & ~x192 & ~x193 & ~x194 & ~x195 & ~x196 & ~x198 & ~x199 & ~x200 & ~x204 & ~x206 & ~x207 & ~x210 & ~x221 & ~x222 & ~x225 & ~x227 & ~x228 & ~x229 & ~x230 & ~x231 & ~x232 & ~x236 & ~x238 & ~x248 & ~x249 & ~x250 & ~x251 & ~x252 & ~x253 & ~x254 & ~x257 & ~x259 & ~x260 & ~x263 & ~x264 & ~x265 & ~x266 & ~x276 & ~x278 & ~x279 & ~x280 & ~x281 & ~x282 & ~x283 & ~x284 & ~x285 & ~x286 & ~x287 & ~x289 & ~x290 & ~x291 & ~x303 & ~x304 & ~x305 & ~x307 & ~x311 & ~x316 & ~x318 & ~x320 & ~x330 & ~x331 & ~x332 & ~x333 & ~x336 & ~x337 & ~x338 & ~x339 & ~x341 & ~x342 & ~x343 & ~x344 & ~x346 & ~x348 & ~x358 & ~x361 & ~x363 & ~x364 & ~x365 & ~x367 & ~x370 & ~x371 & ~x372 & ~x373 & ~x374 & ~x384 & ~x385 & ~x387 & ~x389 & ~x390 & ~x391 & ~x393 & ~x396 & ~x397 & ~x399 & ~x400 & ~x401 & ~x402 & ~x411 & ~x415 & ~x417 & ~x425 & ~x428 & ~x429 & ~x438 & ~x440 & ~x443 & ~x444 & ~x446 & ~x449 & ~x450 & ~x452 & ~x453 & ~x454 & ~x455 & ~x456 & ~x466 & ~x467 & ~x468 & ~x470 & ~x471 & ~x474 & ~x476 & ~x477 & ~x478 & ~x480 & ~x481 & ~x482 & ~x494 & ~x499 & ~x501 & ~x502 & ~x503 & ~x506 & ~x509 & ~x521 & ~x522 & ~x524 & ~x527 & ~x528 & ~x531 & ~x532 & ~x534 & ~x536 & ~x537 & ~x548 & ~x549 & ~x550 & ~x551 & ~x552 & ~x553 & ~x561 & ~x562 & ~x563 & ~x574 & ~x575 & ~x576 & ~x577 & ~x578 & ~x579 & ~x581 & ~x582 & ~x583 & ~x585 & ~x589 & ~x590 & ~x601 & ~x602 & ~x605 & ~x606 & ~x608 & ~x610 & ~x611 & ~x613 & ~x616 & ~x617 & ~x618 & ~x619 & ~x628 & ~x629 & ~x631 & ~x632 & ~x634 & ~x636 & ~x637 & ~x638 & ~x639 & ~x640 & ~x643 & ~x644 & ~x645 & ~x646 & ~x647 & ~x656 & ~x658 & ~x660 & ~x662 & ~x667 & ~x670 & ~x673 & ~x674 & ~x675 & ~x682 & ~x685 & ~x686 & ~x688 & ~x692 & ~x698 & ~x699 & ~x701 & ~x702 & ~x703 & ~x706 & ~x707 & ~x708 & ~x710 & ~x713 & ~x715 & ~x718 & ~x719 & ~x725 & ~x726 & ~x728 & ~x729 & ~x730 & ~x731 & ~x733 & ~x734 & ~x739 & ~x742 & ~x746 & ~x748 & ~x750 & ~x751 & ~x752 & ~x753 & ~x756 & ~x757 & ~x758 & ~x760 & ~x761 & ~x764 & ~x767 & ~x769 & ~x770 & ~x771 & ~x772 & ~x773 & ~x778 & ~x779;
assign c1244 =  x195;
assign c1246 =  x60;
assign c1248 =  x532;
assign c1250 =  x295 &  x322 &  x350 &  x351 &  x404 &  x405 &  x406 &  x461 &  x488 &  x517 &  x543 &  x545 &  x599 &  x600 & ~x2 & ~x4 & ~x14 & ~x15 & ~x35 & ~x49 & ~x51 & ~x65 & ~x68 & ~x74 & ~x76 & ~x77 & ~x90 & ~x101 & ~x109 & ~x116 & ~x121 & ~x132 & ~x143 & ~x144 & ~x146 & ~x163 & ~x172 & ~x195 & ~x198 & ~x203 & ~x204 & ~x253 & ~x257 & ~x258 & ~x280 & ~x286 & ~x302 & ~x308 & ~x310 & ~x313 & ~x316 & ~x317 & ~x318 & ~x331 & ~x341 & ~x345 & ~x358 & ~x360 & ~x361 & ~x369 & ~x370 & ~x374 & ~x400 & ~x412 & ~x417 & ~x423 & ~x427 & ~x441 & ~x444 & ~x449 & ~x453 & ~x468 & ~x476 & ~x479 & ~x497 & ~x498 & ~x525 & ~x539 & ~x553 & ~x556 & ~x565 & ~x580 & ~x583 & ~x585 & ~x622 & ~x643 & ~x650 & ~x670 & ~x677 & ~x699 & ~x715 & ~x716 & ~x718 & ~x732 & ~x740 & ~x747 & ~x749 & ~x754 & ~x757 & ~x774;
assign c1252 =  x239 &  x322 &  x489 &  x517 &  x545 & ~x7 & ~x19 & ~x33 & ~x37 & ~x57 & ~x58 & ~x64 & ~x85 & ~x86 & ~x94 & ~x118 & ~x119 & ~x130 & ~x133 & ~x141 & ~x168 & ~x206 & ~x223 & ~x226 & ~x227 & ~x233 & ~x275 & ~x278 & ~x286 & ~x342 & ~x359 & ~x373 & ~x386 & ~x411 & ~x427 & ~x428 & ~x445 & ~x446 & ~x452 & ~x456 & ~x471 & ~x472 & ~x502 & ~x508 & ~x525 & ~x530 & ~x532 & ~x533 & ~x534 & ~x566 & ~x596 & ~x624 & ~x637 & ~x642 & ~x668 & ~x670 & ~x677 & ~x707 & ~x720 & ~x721 & ~x722 & ~x724 & ~x726 & ~x727 & ~x736 & ~x775 & ~x777 & ~x783;
assign c1254 =  x732;
assign c1256 =  x295 &  x322 &  x350 &  x546 &  x574 & ~x0 & ~x5 & ~x28 & ~x39 & ~x52 & ~x57 & ~x59 & ~x66 & ~x67 & ~x70 & ~x76 & ~x78 & ~x79 & ~x81 & ~x82 & ~x83 & ~x95 & ~x98 & ~x100 & ~x110 & ~x112 & ~x118 & ~x121 & ~x123 & ~x142 & ~x147 & ~x164 & ~x165 & ~x169 & ~x171 & ~x173 & ~x174 & ~x188 & ~x190 & ~x191 & ~x192 & ~x195 & ~x198 & ~x201 & ~x202 & ~x203 & ~x227 & ~x251 & ~x257 & ~x258 & ~x261 & ~x262 & ~x277 & ~x279 & ~x282 & ~x290 & ~x307 & ~x314 & ~x336 & ~x338 & ~x340 & ~x341 & ~x365 & ~x366 & ~x368 & ~x369 & ~x371 & ~x389 & ~x394 & ~x396 & ~x411 & ~x426 & ~x427 & ~x440 & ~x443 & ~x446 & ~x447 & ~x448 & ~x451 & ~x467 & ~x468 & ~x474 & ~x476 & ~x478 & ~x483 & ~x502 & ~x508 & ~x509 & ~x524 & ~x526 & ~x527 & ~x534 & ~x535 & ~x557 & ~x560 & ~x565 & ~x568 & ~x584 & ~x590 & ~x593 & ~x596 & ~x617 & ~x638 & ~x642 & ~x648 & ~x666 & ~x675 & ~x676 & ~x679 & ~x692 & ~x700 & ~x701 & ~x702 & ~x722 & ~x727 & ~x728 & ~x730 & ~x732 & ~x733 & ~x737 & ~x738 & ~x746 & ~x747 & ~x751 & ~x764 & ~x768 & ~x770 & ~x771 & ~x773 & ~x774 & ~x775 & ~x782 & ~x783;
assign c1258 =  x489 & ~x5 & ~x13 & ~x19 & ~x43 & ~x44 & ~x60 & ~x65 & ~x72 & ~x88 & ~x97 & ~x100 & ~x117 & ~x134 & ~x137 & ~x147 & ~x151 & ~x153 & ~x174 & ~x178 & ~x190 & ~x192 & ~x197 & ~x201 & ~x206 & ~x207 & ~x208 & ~x209 & ~x220 & ~x228 & ~x231 & ~x232 & ~x248 & ~x264 & ~x274 & ~x275 & ~x280 & ~x289 & ~x310 & ~x317 & ~x318 & ~x319 & ~x328 & ~x335 & ~x343 & ~x348 & ~x356 & ~x362 & ~x370 & ~x375 & ~x382 & ~x402 & ~x409 & ~x418 & ~x421 & ~x423 & ~x437 & ~x446 & ~x457 & ~x464 & ~x466 & ~x468 & ~x519 & ~x521 & ~x526 & ~x527 & ~x529 & ~x537 & ~x538 & ~x540 & ~x547 & ~x553 & ~x558 & ~x566 & ~x588 & ~x591 & ~x594 & ~x595 & ~x603 & ~x612 & ~x634 & ~x646 & ~x662 & ~x666 & ~x677 & ~x678 & ~x690 & ~x691 & ~x700 & ~x706 & ~x710 & ~x712 & ~x714 & ~x723 & ~x747 & ~x750 & ~x758 & ~x759 & ~x778;
assign c1260 =  x782;
assign c1262 =  x335;
assign c1264 =  x55;
assign c1266 =  x87;
assign c1268 = ~x0 & ~x20 & ~x24 & ~x29 & ~x33 & ~x50 & ~x63 & ~x81 & ~x92 & ~x117 & ~x120 & ~x176 & ~x187 & ~x199 & ~x203 & ~x231 & ~x233 & ~x258 & ~x272 & ~x279 & ~x290 & ~x312 & ~x319 & ~x336 & ~x386 & ~x418 & ~x419 & ~x425 & ~x437 & ~x442 & ~x447 & ~x449 & ~x457 & ~x494 & ~x500 & ~x515 & ~x523 & ~x563 & ~x582 & ~x584 & ~x588 & ~x619 & ~x620 & ~x640 & ~x671 & ~x693 & ~x713 & ~x745 & ~x758;
assign c1270 =  x14;
assign c1272 =  x351 &  x378 &  x406 &  x433 & ~x0 & ~x2 & ~x3 & ~x4 & ~x7 & ~x10 & ~x11 & ~x13 & ~x14 & ~x15 & ~x18 & ~x19 & ~x23 & ~x25 & ~x27 & ~x28 & ~x29 & ~x32 & ~x34 & ~x35 & ~x37 & ~x40 & ~x41 & ~x43 & ~x44 & ~x48 & ~x49 & ~x51 & ~x53 & ~x58 & ~x60 & ~x61 & ~x62 & ~x64 & ~x66 & ~x68 & ~x70 & ~x72 & ~x76 & ~x78 & ~x79 & ~x82 & ~x86 & ~x87 & ~x88 & ~x89 & ~x90 & ~x91 & ~x92 & ~x97 & ~x100 & ~x105 & ~x109 & ~x110 & ~x111 & ~x112 & ~x113 & ~x114 & ~x117 & ~x119 & ~x120 & ~x122 & ~x125 & ~x126 & ~x135 & ~x136 & ~x141 & ~x142 & ~x143 & ~x144 & ~x145 & ~x146 & ~x149 & ~x150 & ~x151 & ~x152 & ~x153 & ~x163 & ~x165 & ~x166 & ~x169 & ~x170 & ~x173 & ~x176 & ~x177 & ~x179 & ~x192 & ~x195 & ~x199 & ~x204 & ~x220 & ~x221 & ~x222 & ~x227 & ~x233 & ~x234 & ~x237 & ~x245 & ~x246 & ~x247 & ~x248 & ~x251 & ~x253 & ~x254 & ~x258 & ~x261 & ~x262 & ~x264 & ~x273 & ~x274 & ~x276 & ~x282 & ~x283 & ~x286 & ~x287 & ~x289 & ~x292 & ~x302 & ~x303 & ~x304 & ~x305 & ~x309 & ~x310 & ~x312 & ~x313 & ~x314 & ~x315 & ~x316 & ~x318 & ~x320 & ~x328 & ~x330 & ~x334 & ~x335 & ~x336 & ~x337 & ~x338 & ~x339 & ~x340 & ~x342 & ~x344 & ~x345 & ~x346 & ~x347 & ~x348 & ~x356 & ~x358 & ~x359 & ~x360 & ~x362 & ~x364 & ~x365 & ~x366 & ~x368 & ~x372 & ~x373 & ~x374 & ~x375 & ~x383 & ~x388 & ~x393 & ~x395 & ~x396 & ~x398 & ~x399 & ~x400 & ~x401 & ~x415 & ~x416 & ~x422 & ~x427 & ~x428 & ~x429 & ~x438 & ~x439 & ~x442 & ~x443 & ~x444 & ~x446 & ~x447 & ~x449 & ~x450 & ~x452 & ~x454 & ~x455 & ~x466 & ~x468 & ~x470 & ~x472 & ~x474 & ~x476 & ~x480 & ~x481 & ~x482 & ~x493 & ~x494 & ~x495 & ~x499 & ~x500 & ~x502 & ~x504 & ~x506 & ~x510 & ~x511 & ~x521 & ~x522 & ~x527 & ~x528 & ~x533 & ~x536 & ~x537 & ~x538 & ~x547 & ~x548 & ~x549 & ~x550 & ~x554 & ~x555 & ~x560 & ~x564 & ~x565 & ~x566 & ~x575 & ~x582 & ~x584 & ~x587 & ~x588 & ~x589 & ~x591 & ~x603 & ~x608 & ~x612 & ~x615 & ~x619 & ~x620 & ~x621 & ~x634 & ~x635 & ~x638 & ~x640 & ~x641 & ~x644 & ~x648 & ~x662 & ~x666 & ~x671 & ~x672 & ~x674 & ~x677 & ~x678 & ~x686 & ~x690 & ~x692 & ~x695 & ~x703 & ~x704 & ~x705 & ~x707 & ~x708 & ~x709 & ~x711 & ~x713 & ~x714 & ~x717 & ~x718 & ~x720 & ~x722 & ~x723 & ~x730 & ~x733 & ~x735 & ~x742 & ~x743 & ~x745 & ~x748 & ~x749 & ~x751 & ~x755 & ~x757 & ~x759 & ~x760 & ~x762 & ~x765 & ~x773 & ~x774 & ~x775 & ~x778 & ~x783;
assign c1274 =  x268 &  x269 &  x296 &  x324 &  x351 &  x352 &  x406 &  x462 &  x544 &  x572 & ~x3 & ~x7 & ~x8 & ~x9 & ~x11 & ~x13 & ~x15 & ~x17 & ~x23 & ~x26 & ~x33 & ~x36 & ~x38 & ~x42 & ~x44 & ~x47 & ~x48 & ~x51 & ~x54 & ~x55 & ~x61 & ~x63 & ~x64 & ~x68 & ~x71 & ~x75 & ~x76 & ~x81 & ~x82 & ~x89 & ~x91 & ~x92 & ~x94 & ~x97 & ~x98 & ~x99 & ~x104 & ~x110 & ~x111 & ~x114 & ~x120 & ~x122 & ~x124 & ~x125 & ~x134 & ~x135 & ~x143 & ~x144 & ~x146 & ~x153 & ~x164 & ~x165 & ~x166 & ~x171 & ~x173 & ~x174 & ~x175 & ~x176 & ~x178 & ~x179 & ~x180 & ~x181 & ~x191 & ~x192 & ~x194 & ~x196 & ~x198 & ~x199 & ~x201 & ~x202 & ~x204 & ~x206 & ~x208 & ~x209 & ~x220 & ~x221 & ~x224 & ~x228 & ~x232 & ~x234 & ~x235 & ~x236 & ~x245 & ~x246 & ~x247 & ~x248 & ~x250 & ~x251 & ~x256 & ~x257 & ~x258 & ~x259 & ~x260 & ~x261 & ~x273 & ~x276 & ~x277 & ~x280 & ~x285 & ~x289 & ~x301 & ~x302 & ~x303 & ~x311 & ~x312 & ~x313 & ~x315 & ~x316 & ~x330 & ~x335 & ~x336 & ~x339 & ~x341 & ~x355 & ~x359 & ~x361 & ~x364 & ~x369 & ~x370 & ~x384 & ~x387 & ~x394 & ~x397 & ~x399 & ~x401 & ~x422 & ~x438 & ~x439 & ~x440 & ~x443 & ~x445 & ~x446 & ~x447 & ~x449 & ~x450 & ~x451 & ~x452 & ~x456 & ~x466 & ~x471 & ~x475 & ~x476 & ~x478 & ~x480 & ~x481 & ~x483 & ~x494 & ~x497 & ~x498 & ~x499 & ~x501 & ~x503 & ~x504 & ~x508 & ~x511 & ~x512 & ~x522 & ~x526 & ~x527 & ~x537 & ~x539 & ~x555 & ~x556 & ~x560 & ~x564 & ~x565 & ~x566 & ~x578 & ~x580 & ~x581 & ~x582 & ~x585 & ~x589 & ~x590 & ~x591 & ~x607 & ~x608 & ~x610 & ~x613 & ~x614 & ~x618 & ~x619 & ~x621 & ~x635 & ~x650 & ~x661 & ~x662 & ~x663 & ~x665 & ~x668 & ~x670 & ~x672 & ~x675 & ~x677 & ~x679 & ~x692 & ~x694 & ~x695 & ~x696 & ~x697 & ~x701 & ~x706 & ~x707 & ~x716 & ~x720 & ~x725 & ~x726 & ~x737 & ~x742 & ~x743 & ~x744 & ~x745 & ~x746 & ~x747 & ~x752 & ~x754 & ~x755 & ~x765 & ~x772 & ~x774 & ~x779 & ~x781;
assign c1276 = ~x4 & ~x5 & ~x8 & ~x10 & ~x16 & ~x17 & ~x25 & ~x26 & ~x31 & ~x32 & ~x34 & ~x36 & ~x37 & ~x40 & ~x44 & ~x45 & ~x46 & ~x47 & ~x50 & ~x51 & ~x53 & ~x55 & ~x56 & ~x59 & ~x63 & ~x68 & ~x73 & ~x75 & ~x77 & ~x80 & ~x84 & ~x89 & ~x93 & ~x94 & ~x98 & ~x112 & ~x113 & ~x120 & ~x124 & ~x133 & ~x136 & ~x138 & ~x141 & ~x145 & ~x146 & ~x147 & ~x148 & ~x149 & ~x151 & ~x172 & ~x174 & ~x190 & ~x191 & ~x192 & ~x196 & ~x204 & ~x207 & ~x220 & ~x221 & ~x222 & ~x223 & ~x232 & ~x245 & ~x248 & ~x249 & ~x251 & ~x252 & ~x255 & ~x256 & ~x261 & ~x263 & ~x276 & ~x280 & ~x282 & ~x283 & ~x284 & ~x288 & ~x291 & ~x303 & ~x308 & ~x311 & ~x312 & ~x315 & ~x331 & ~x332 & ~x339 & ~x340 & ~x344 & ~x353 & ~x360 & ~x369 & ~x370 & ~x371 & ~x372 & ~x381 & ~x386 & ~x388 & ~x391 & ~x394 & ~x400 & ~x401 & ~x402 & ~x408 & ~x419 & ~x420 & ~x422 & ~x429 & ~x444 & ~x448 & ~x452 & ~x454 & ~x455 & ~x465 & ~x468 & ~x470 & ~x471 & ~x474 & ~x477 & ~x482 & ~x483 & ~x484 & ~x491 & ~x493 & ~x504 & ~x505 & ~x519 & ~x520 & ~x521 & ~x523 & ~x527 & ~x533 & ~x539 & ~x540 & ~x553 & ~x557 & ~x560 & ~x561 & ~x565 & ~x567 & ~x588 & ~x613 & ~x614 & ~x619 & ~x641 & ~x643 & ~x647 & ~x649 & ~x659 & ~x660 & ~x661 & ~x662 & ~x666 & ~x669 & ~x679 & ~x690 & ~x691 & ~x693 & ~x694 & ~x696 & ~x698 & ~x705 & ~x707 & ~x708 & ~x711 & ~x712 & ~x715 & ~x717 & ~x718 & ~x719 & ~x720 & ~x722 & ~x723 & ~x730 & ~x736 & ~x738 & ~x740 & ~x758 & ~x759 & ~x761 & ~x769 & ~x771 & ~x773 & ~x775 & ~x780 & ~x781;
assign c1278 =  x239 &  x267 &  x295 &  x323 &  x350 &  x378 &  x405 &  x434 &  x461 &  x489 &  x490 &  x544 &  x572 &  x600 & ~x1 & ~x4 & ~x7 & ~x17 & ~x20 & ~x21 & ~x23 & ~x24 & ~x26 & ~x29 & ~x33 & ~x34 & ~x35 & ~x37 & ~x40 & ~x41 & ~x46 & ~x48 & ~x49 & ~x50 & ~x54 & ~x55 & ~x57 & ~x58 & ~x62 & ~x63 & ~x67 & ~x68 & ~x75 & ~x77 & ~x78 & ~x83 & ~x87 & ~x89 & ~x95 & ~x100 & ~x101 & ~x104 & ~x110 & ~x120 & ~x123 & ~x124 & ~x136 & ~x143 & ~x144 & ~x147 & ~x150 & ~x163 & ~x164 & ~x168 & ~x170 & ~x172 & ~x177 & ~x190 & ~x200 & ~x202 & ~x203 & ~x220 & ~x225 & ~x227 & ~x245 & ~x248 & ~x254 & ~x257 & ~x277 & ~x306 & ~x307 & ~x312 & ~x328 & ~x329 & ~x332 & ~x334 & ~x337 & ~x344 & ~x359 & ~x362 & ~x368 & ~x372 & ~x374 & ~x383 & ~x384 & ~x386 & ~x394 & ~x397 & ~x399 & ~x400 & ~x415 & ~x417 & ~x420 & ~x423 & ~x429 & ~x439 & ~x444 & ~x447 & ~x449 & ~x451 & ~x452 & ~x456 & ~x469 & ~x474 & ~x476 & ~x477 & ~x493 & ~x497 & ~x499 & ~x502 & ~x506 & ~x507 & ~x510 & ~x525 & ~x530 & ~x532 & ~x534 & ~x538 & ~x556 & ~x558 & ~x561 & ~x564 & ~x582 & ~x591 & ~x609 & ~x612 & ~x617 & ~x640 & ~x669 & ~x674 & ~x688 & ~x689 & ~x693 & ~x701 & ~x702 & ~x704 & ~x706 & ~x707 & ~x711 & ~x715 & ~x716 & ~x717 & ~x718 & ~x724 & ~x725 & ~x726 & ~x728 & ~x731 & ~x732 & ~x740 & ~x741 & ~x743 & ~x745 & ~x746 & ~x747 & ~x748 & ~x753 & ~x755 & ~x756 & ~x757 & ~x761 & ~x765 & ~x767 & ~x768 & ~x771 & ~x773;
assign c1280 =  x325 &  x352 &  x379 &  x406 &  x460 &  x461 &  x487 &  x488 &  x515 &  x542 & ~x6 & ~x10 & ~x12 & ~x14 & ~x20 & ~x27 & ~x36 & ~x38 & ~x45 & ~x52 & ~x56 & ~x62 & ~x64 & ~x70 & ~x77 & ~x91 & ~x94 & ~x95 & ~x96 & ~x100 & ~x101 & ~x113 & ~x124 & ~x125 & ~x127 & ~x129 & ~x136 & ~x144 & ~x150 & ~x152 & ~x154 & ~x155 & ~x167 & ~x169 & ~x174 & ~x178 & ~x179 & ~x180 & ~x182 & ~x183 & ~x196 & ~x203 & ~x204 & ~x206 & ~x207 & ~x228 & ~x231 & ~x236 & ~x237 & ~x257 & ~x261 & ~x262 & ~x265 & ~x292 & ~x307 & ~x308 & ~x318 & ~x320 & ~x334 & ~x344 & ~x345 & ~x347 & ~x348 & ~x357 & ~x365 & ~x367 & ~x372 & ~x373 & ~x384 & ~x394 & ~x397 & ~x398 & ~x411 & ~x412 & ~x438 & ~x444 & ~x455 & ~x466 & ~x467 & ~x478 & ~x503 & ~x506 & ~x508 & ~x520 & ~x521 & ~x522 & ~x524 & ~x525 & ~x526 & ~x533 & ~x537 & ~x548 & ~x549 & ~x553 & ~x556 & ~x558 & ~x575 & ~x581 & ~x601 & ~x602 & ~x604 & ~x610 & ~x617 & ~x629 & ~x630 & ~x631 & ~x644 & ~x646 & ~x647 & ~x660 & ~x668 & ~x671 & ~x675 & ~x676 & ~x683 & ~x684 & ~x706 & ~x715 & ~x716 & ~x718 & ~x722 & ~x729 & ~x739 & ~x741 & ~x747 & ~x754;
assign c1282 =  x292 & ~x20 & ~x49 & ~x56 & ~x68 & ~x89 & ~x108 & ~x185 & ~x250 & ~x259 & ~x307 & ~x311 & ~x364 & ~x416 & ~x423 & ~x430 & ~x442 & ~x443 & ~x487 & ~x503 & ~x592 & ~x596 & ~x613 & ~x616 & ~x645 & ~x665 & ~x685 & ~x760 & ~x782;
assign c1284 =  x154 &  x211 &  x295 &  x322 &  x350 &  x378 & ~x2 & ~x12 & ~x14 & ~x23 & ~x26 & ~x29 & ~x36 & ~x57 & ~x63 & ~x75 & ~x85 & ~x93 & ~x111 & ~x115 & ~x116 & ~x121 & ~x139 & ~x143 & ~x148 & ~x166 & ~x187 & ~x188 & ~x199 & ~x202 & ~x205 & ~x216 & ~x227 & ~x229 & ~x242 & ~x253 & ~x270 & ~x271 & ~x274 & ~x280 & ~x298 & ~x302 & ~x305 & ~x309 & ~x327 & ~x369 & ~x396 & ~x401 & ~x411 & ~x453 & ~x454 & ~x468 & ~x483 & ~x497 & ~x532 & ~x539 & ~x583 & ~x618 & ~x621 & ~x636 & ~x639 & ~x650 & ~x663 & ~x665 & ~x668 & ~x672 & ~x683 & ~x692 & ~x702 & ~x715 & ~x718 & ~x727 & ~x735 & ~x752 & ~x759 & ~x764 & ~x770 & ~x777 & ~x781 & ~x782;
assign c1286 =  x645;
assign c1288 =  x674;
assign c1290 =  x37;
assign c1292 =  x323 &  x407 & ~x3 & ~x9 & ~x17 & ~x20 & ~x28 & ~x41 & ~x72 & ~x87 & ~x93 & ~x94 & ~x105 & ~x112 & ~x119 & ~x142 & ~x160 & ~x172 & ~x199 & ~x219 & ~x220 & ~x223 & ~x227 & ~x231 & ~x250 & ~x253 & ~x262 & ~x270 & ~x273 & ~x289 & ~x298 & ~x332 & ~x376 & ~x383 & ~x390 & ~x391 & ~x393 & ~x398 & ~x403 & ~x422 & ~x428 & ~x429 & ~x432 & ~x442 & ~x447 & ~x450 & ~x475 & ~x478 & ~x487 & ~x500 & ~x512 & ~x533 & ~x534 & ~x584 & ~x590 & ~x615 & ~x619 & ~x642 & ~x645 & ~x647 & ~x665 & ~x687 & ~x697 & ~x701 & ~x719 & ~x732 & ~x736 & ~x772 & ~x773;
assign c1294 =  x308 &  x698;
assign c1296 =  x297 &  x298 &  x324 &  x325 &  x351 &  x379 &  x435 &  x570 &  x624 & ~x97 & ~x123 & ~x124 & ~x154 & ~x183 & ~x208 & ~x210 & ~x228 & ~x265 & ~x292 & ~x293 & ~x318 & ~x320 & ~x374 & ~x400 & ~x453 & ~x465 & ~x493 & ~x629;
assign c1298 =  x268 &  x351 &  x378 &  x406 &  x434 &  x488 &  x489 &  x515 &  x516 &  x544 &  x572 &  x600 &  x627 & ~x3 & ~x6 & ~x7 & ~x9 & ~x10 & ~x11 & ~x12 & ~x14 & ~x18 & ~x30 & ~x31 & ~x33 & ~x34 & ~x37 & ~x42 & ~x46 & ~x50 & ~x51 & ~x52 & ~x56 & ~x57 & ~x59 & ~x62 & ~x63 & ~x69 & ~x70 & ~x73 & ~x75 & ~x77 & ~x78 & ~x80 & ~x81 & ~x84 & ~x85 & ~x86 & ~x89 & ~x90 & ~x94 & ~x95 & ~x98 & ~x99 & ~x101 & ~x103 & ~x106 & ~x107 & ~x111 & ~x113 & ~x119 & ~x120 & ~x121 & ~x123 & ~x124 & ~x125 & ~x134 & ~x136 & ~x137 & ~x140 & ~x142 & ~x143 & ~x146 & ~x148 & ~x149 & ~x151 & ~x164 & ~x165 & ~x167 & ~x172 & ~x174 & ~x175 & ~x177 & ~x178 & ~x181 & ~x192 & ~x195 & ~x200 & ~x201 & ~x205 & ~x207 & ~x218 & ~x219 & ~x220 & ~x221 & ~x222 & ~x224 & ~x229 & ~x230 & ~x233 & ~x235 & ~x246 & ~x247 & ~x249 & ~x250 & ~x252 & ~x257 & ~x258 & ~x259 & ~x260 & ~x264 & ~x276 & ~x279 & ~x280 & ~x282 & ~x284 & ~x287 & ~x289 & ~x290 & ~x291 & ~x302 & ~x304 & ~x305 & ~x306 & ~x307 & ~x309 & ~x310 & ~x311 & ~x312 & ~x313 & ~x317 & ~x318 & ~x330 & ~x337 & ~x339 & ~x340 & ~x343 & ~x345 & ~x346 & ~x361 & ~x366 & ~x367 & ~x370 & ~x371 & ~x372 & ~x374 & ~x387 & ~x392 & ~x393 & ~x396 & ~x397 & ~x398 & ~x400 & ~x401 & ~x414 & ~x416 & ~x417 & ~x418 & ~x419 & ~x423 & ~x425 & ~x427 & ~x428 & ~x444 & ~x445 & ~x448 & ~x451 & ~x454 & ~x455 & ~x456 & ~x467 & ~x468 & ~x469 & ~x471 & ~x474 & ~x476 & ~x477 & ~x479 & ~x480 & ~x481 & ~x482 & ~x483 & ~x497 & ~x501 & ~x503 & ~x504 & ~x509 & ~x521 & ~x524 & ~x527 & ~x530 & ~x532 & ~x535 & ~x538 & ~x552 & ~x553 & ~x557 & ~x558 & ~x562 & ~x563 & ~x564 & ~x565 & ~x566 & ~x581 & ~x582 & ~x585 & ~x591 & ~x605 & ~x606 & ~x608 & ~x610 & ~x612 & ~x614 & ~x618 & ~x632 & ~x637 & ~x641 & ~x642 & ~x643 & ~x646 & ~x647 & ~x666 & ~x672 & ~x674 & ~x675 & ~x679 & ~x680 & ~x694 & ~x695 & ~x696 & ~x700 & ~x703 & ~x707 & ~x708 & ~x710 & ~x719 & ~x721 & ~x722 & ~x724 & ~x726 & ~x727 & ~x728 & ~x730 & ~x732 & ~x733 & ~x735 & ~x737 & ~x738 & ~x741 & ~x742 & ~x743 & ~x745 & ~x746 & ~x751 & ~x752 & ~x753 & ~x754 & ~x756 & ~x757 & ~x760 & ~x761 & ~x762 & ~x764 & ~x766 & ~x768 & ~x769 & ~x772 & ~x774 & ~x777;
assign c11 =  x542 & ~x30 & ~x34 & ~x42 & ~x61 & ~x72 & ~x109 & ~x115 & ~x161 & ~x195 & ~x199 & ~x215 & ~x218 & ~x224 & ~x243 & ~x250 & ~x293 & ~x308 & ~x310 & ~x312 & ~x332 & ~x335 & ~x394 & ~x474 & ~x529 & ~x564 & ~x566 & ~x615 & ~x647 & ~x666 & ~x729 & ~x761 & ~x766 & ~x772 & ~x778;
assign c13 =  x316 & ~x1 & ~x4 & ~x22 & ~x23 & ~x26 & ~x28 & ~x41 & ~x43 & ~x50 & ~x51 & ~x53 & ~x55 & ~x59 & ~x69 & ~x73 & ~x76 & ~x81 & ~x84 & ~x90 & ~x99 & ~x100 & ~x106 & ~x107 & ~x111 & ~x113 & ~x118 & ~x125 & ~x127 & ~x131 & ~x133 & ~x136 & ~x139 & ~x140 & ~x142 & ~x143 & ~x172 & ~x198 & ~x222 & ~x225 & ~x226 & ~x279 & ~x280 & ~x308 & ~x334 & ~x335 & ~x337 & ~x362 & ~x365 & ~x418 & ~x419 & ~x445 & ~x448 & ~x451 & ~x474 & ~x506 & ~x529 & ~x534 & ~x555 & ~x561 & ~x587 & ~x588 & ~x615 & ~x619 & ~x620 & ~x622 & ~x623 & ~x644 & ~x669 & ~x679 & ~x699 & ~x701 & ~x702 & ~x704 & ~x725 & ~x730 & ~x752 & ~x753 & ~x765 & ~x766 & ~x770 & ~x779 & ~x783;
assign c15 =  x352 &  x406 & ~x11 & ~x17 & ~x27 & ~x45 & ~x82 & ~x85 & ~x105 & ~x115 & ~x159 & ~x161 & ~x163 & ~x170 & ~x174 & ~x188 & ~x195 & ~x201 & ~x217 & ~x225 & ~x230 & ~x257 & ~x309 & ~x322 & ~x369 & ~x388 & ~x447 & ~x454 & ~x473 & ~x479 & ~x498 & ~x553 & ~x559 & ~x563 & ~x590 & ~x594 & ~x614 & ~x615 & ~x616 & ~x621 & ~x675 & ~x691 & ~x696 & ~x700 & ~x702 & ~x726 & ~x729 & ~x748 & ~x753 & ~x759 & ~x762;
assign c17 =  x217 &  x238 & ~x27 & ~x174 & ~x201 & ~x254 & ~x398 & ~x504 & ~x751;
assign c19 =  x573 & ~x1 & ~x25 & ~x39 & ~x40 & ~x56 & ~x61 & ~x62 & ~x78 & ~x82 & ~x83 & ~x111 & ~x114 & ~x140 & ~x177 & ~x203 & ~x224 & ~x232 & ~x260 & ~x288 & ~x307 & ~x314 & ~x323 & ~x339 & ~x361 & ~x370 & ~x396 & ~x398 & ~x411 & ~x415 & ~x418 & ~x445 & ~x450 & ~x452 & ~x470 & ~x500 & ~x530 & ~x531 & ~x532 & ~x584 & ~x592 & ~x612 & ~x613 & ~x616 & ~x618 & ~x634 & ~x640 & ~x643 & ~x660 & ~x666 & ~x667 & ~x669 & ~x670 & ~x687 & ~x689 & ~x697 & ~x704 & ~x714 & ~x716 & ~x727 & ~x732 & ~x745 & ~x748 & ~x749 & ~x752 & ~x753 & ~x758 & ~x762 & ~x774 & ~x777;
assign c111 =  x383 & ~x0 & ~x24 & ~x28 & ~x43 & ~x53 & ~x55 & ~x62 & ~x67 & ~x86 & ~x90 & ~x143 & ~x163 & ~x251 & ~x278 & ~x335 & ~x376 & ~x449 & ~x476 & ~x502 & ~x506 & ~x531 & ~x558 & ~x589 & ~x640 & ~x643 & ~x645 & ~x669 & ~x673 & ~x694 & ~x700 & ~x727 & ~x744 & ~x752 & ~x754 & ~x765 & ~x768 & ~x769;
assign c113 =  x510 & ~x15 & ~x35 & ~x55 & ~x61 & ~x83 & ~x84 & ~x87 & ~x173 & ~x198 & ~x199 & ~x280 & ~x336 & ~x418 & ~x424 & ~x474 & ~x503 & ~x585 & ~x674 & ~x678 & ~x701 & ~x743 & ~x766 & ~x783;
assign c115 =  x521 & ~x30 & ~x46 & ~x75 & ~x83 & ~x262 & ~x335 & ~x443 & ~x490 & ~x532 & ~x581 & ~x583 & ~x586 & ~x648 & ~x737 & ~x782;
assign c117 =  x401 &  x431 & ~x31 & ~x44 & ~x49 & ~x55 & ~x59 & ~x70 & ~x88 & ~x118 & ~x123 & ~x128 & ~x224 & ~x225 & ~x311 & ~x334 & ~x336 & ~x392 & ~x416 & ~x421 & ~x476 & ~x479 & ~x502 & ~x507 & ~x529 & ~x531 & ~x591 & ~x612 & ~x619 & ~x641 & ~x643 & ~x645 & ~x695 & ~x706 & ~x734 & ~x755 & ~x775;
assign c119 = ~x0 & ~x3 & ~x5 & ~x9 & ~x16 & ~x20 & ~x22 & ~x37 & ~x45 & ~x46 & ~x65 & ~x76 & ~x78 & ~x91 & ~x94 & ~x100 & ~x101 & ~x105 & ~x106 & ~x110 & ~x117 & ~x139 & ~x141 & ~x144 & ~x145 & ~x172 & ~x198 & ~x223 & ~x280 & ~x308 & ~x309 & ~x361 & ~x362 & ~x363 & ~x423 & ~x433 & ~x434 & ~x447 & ~x449 & ~x463 & ~x529 & ~x531 & ~x532 & ~x534 & ~x557 & ~x641 & ~x642 & ~x644 & ~x669 & ~x674 & ~x697 & ~x702 & ~x703 & ~x707 & ~x722 & ~x724 & ~x730 & ~x732 & ~x735 & ~x736 & ~x743 & ~x748 & ~x754 & ~x762 & ~x765 & ~x770;
assign c121 = ~x5 & ~x9 & ~x11 & ~x14 & ~x25 & ~x27 & ~x29 & ~x30 & ~x37 & ~x47 & ~x48 & ~x51 & ~x64 & ~x67 & ~x71 & ~x75 & ~x82 & ~x83 & ~x85 & ~x86 & ~x87 & ~x90 & ~x95 & ~x100 & ~x106 & ~x111 & ~x112 & ~x117 & ~x122 & ~x123 & ~x130 & ~x131 & ~x132 & ~x133 & ~x136 & ~x148 & ~x149 & ~x156 & ~x158 & ~x159 & ~x163 & ~x164 & ~x166 & ~x169 & ~x170 & ~x171 & ~x178 & ~x181 & ~x182 & ~x188 & ~x189 & ~x197 & ~x223 & ~x224 & ~x251 & ~x252 & ~x281 & ~x282 & ~x285 & ~x309 & ~x313 & ~x335 & ~x336 & ~x341 & ~x361 & ~x363 & ~x364 & ~x365 & ~x368 & ~x387 & ~x388 & ~x389 & ~x395 & ~x417 & ~x418 & ~x420 & ~x422 & ~x424 & ~x440 & ~x469 & ~x475 & ~x477 & ~x478 & ~x480 & ~x497 & ~x506 & ~x507 & ~x529 & ~x533 & ~x555 & ~x557 & ~x566 & ~x579 & ~x584 & ~x585 & ~x586 & ~x589 & ~x592 & ~x608 & ~x615 & ~x616 & ~x617 & ~x618 & ~x621 & ~x622 & ~x636 & ~x637 & ~x645 & ~x646 & ~x648 & ~x691 & ~x694 & ~x696 & ~x703 & ~x723 & ~x729 & ~x730 & ~x737 & ~x738 & ~x751 & ~x755 & ~x757 & ~x761 & ~x764 & ~x771 & ~x776 & ~x778 & ~x779;
assign c123 = ~x4 & ~x7 & ~x10 & ~x17 & ~x18 & ~x26 & ~x39 & ~x40 & ~x41 & ~x42 & ~x46 & ~x52 & ~x53 & ~x56 & ~x60 & ~x61 & ~x62 & ~x65 & ~x73 & ~x80 & ~x83 & ~x84 & ~x85 & ~x87 & ~x90 & ~x109 & ~x117 & ~x136 & ~x139 & ~x140 & ~x144 & ~x165 & ~x166 & ~x167 & ~x169 & ~x170 & ~x173 & ~x196 & ~x198 & ~x203 & ~x224 & ~x249 & ~x251 & ~x253 & ~x256 & ~x281 & ~x308 & ~x312 & ~x339 & ~x340 & ~x366 & ~x377 & ~x378 & ~x379 & ~x391 & ~x446 & ~x475 & ~x500 & ~x506 & ~x528 & ~x560 & ~x561 & ~x586 & ~x587 & ~x589 & ~x590 & ~x613 & ~x617 & ~x640 & ~x645 & ~x646 & ~x647 & ~x692 & ~x700 & ~x703 & ~x723 & ~x724 & ~x728 & ~x729 & ~x731 & ~x734 & ~x746 & ~x755 & ~x758 & ~x760 & ~x773 & ~x776 & ~x778;
assign c125 =  x298 & ~x3 & ~x4 & ~x8 & ~x15 & ~x19 & ~x20 & ~x21 & ~x25 & ~x27 & ~x28 & ~x29 & ~x39 & ~x41 & ~x44 & ~x45 & ~x48 & ~x50 & ~x54 & ~x55 & ~x57 & ~x60 & ~x70 & ~x77 & ~x84 & ~x87 & ~x99 & ~x103 & ~x107 & ~x109 & ~x113 & ~x117 & ~x136 & ~x141 & ~x158 & ~x168 & ~x187 & ~x196 & ~x197 & ~x215 & ~x216 & ~x224 & ~x249 & ~x251 & ~x252 & ~x304 & ~x306 & ~x307 & ~x309 & ~x310 & ~x332 & ~x335 & ~x336 & ~x389 & ~x391 & ~x395 & ~x447 & ~x474 & ~x476 & ~x481 & ~x502 & ~x505 & ~x507 & ~x533 & ~x558 & ~x559 & ~x564 & ~x567 & ~x585 & ~x590 & ~x595 & ~x614 & ~x621 & ~x644 & ~x650 & ~x670 & ~x674 & ~x677 & ~x678 & ~x694 & ~x696 & ~x697 & ~x698 & ~x699 & ~x700 & ~x727 & ~x749 & ~x750 & ~x770 & ~x780 & ~x783;
assign c127 =  x437 & ~x7 & ~x9 & ~x10 & ~x14 & ~x25 & ~x28 & ~x54 & ~x56 & ~x59 & ~x61 & ~x66 & ~x84 & ~x88 & ~x90 & ~x92 & ~x93 & ~x113 & ~x137 & ~x144 & ~x152 & ~x174 & ~x192 & ~x197 & ~x215 & ~x222 & ~x225 & ~x280 & ~x284 & ~x337 & ~x391 & ~x392 & ~x394 & ~x395 & ~x419 & ~x420 & ~x444 & ~x473 & ~x476 & ~x502 & ~x505 & ~x532 & ~x554 & ~x556 & ~x560 & ~x562 & ~x579 & ~x580 & ~x589 & ~x634 & ~x636 & ~x645 & ~x647 & ~x663 & ~x666 & ~x691 & ~x698 & ~x699 & ~x701 & ~x703 & ~x716 & ~x718 & ~x723 & ~x733 & ~x745 & ~x754 & ~x759 & ~x780;
assign c129 =  x326 & ~x0 & ~x1 & ~x4 & ~x12 & ~x16 & ~x21 & ~x32 & ~x41 & ~x68 & ~x89 & ~x102 & ~x135 & ~x140 & ~x143 & ~x161 & ~x168 & ~x196 & ~x296 & ~x307 & ~x310 & ~x312 & ~x368 & ~x393 & ~x453 & ~x506 & ~x508 & ~x613 & ~x665 & ~x668 & ~x671 & ~x675 & ~x702 & ~x723 & ~x761 & ~x768 & ~x773 & ~x778 & ~x781 & ~x783;
assign c131 =  x374 &  x403 &  x405 & ~x16 & ~x20 & ~x37 & ~x42 & ~x64 & ~x84 & ~x104 & ~x113 & ~x136 & ~x172 & ~x252 & ~x279 & ~x281 & ~x311 & ~x332 & ~x415 & ~x449 & ~x453 & ~x532 & ~x536 & ~x556 & ~x644 & ~x671 & ~x675 & ~x702 & ~x703 & ~x715 & ~x729 & ~x733 & ~x735 & ~x750 & ~x756 & ~x758 & ~x768 & ~x777 & ~x778;
assign c133 =  x271 & ~x1 & ~x3 & ~x6 & ~x10 & ~x16 & ~x17 & ~x20 & ~x30 & ~x32 & ~x33 & ~x34 & ~x40 & ~x41 & ~x42 & ~x44 & ~x50 & ~x61 & ~x64 & ~x70 & ~x71 & ~x74 & ~x84 & ~x88 & ~x91 & ~x98 & ~x99 & ~x103 & ~x104 & ~x105 & ~x111 & ~x113 & ~x114 & ~x132 & ~x135 & ~x136 & ~x141 & ~x149 & ~x154 & ~x157 & ~x164 & ~x168 & ~x188 & ~x222 & ~x252 & ~x253 & ~x281 & ~x282 & ~x307 & ~x309 & ~x335 & ~x361 & ~x362 & ~x364 & ~x390 & ~x418 & ~x419 & ~x422 & ~x451 & ~x474 & ~x477 & ~x504 & ~x505 & ~x526 & ~x527 & ~x529 & ~x531 & ~x533 & ~x555 & ~x557 & ~x558 & ~x559 & ~x564 & ~x584 & ~x585 & ~x586 & ~x587 & ~x589 & ~x609 & ~x611 & ~x613 & ~x615 & ~x640 & ~x642 & ~x643 & ~x647 & ~x649 & ~x650 & ~x665 & ~x673 & ~x678 & ~x698 & ~x702 & ~x703 & ~x704 & ~x726 & ~x727 & ~x728 & ~x731 & ~x754 & ~x755 & ~x756 & ~x759 & ~x764 & ~x771 & ~x777 & ~x778;
assign c135 =  x457 & ~x14 & ~x37 & ~x54 & ~x64 & ~x75 & ~x77 & ~x84 & ~x106 & ~x110 & ~x115 & ~x194 & ~x197 & ~x225 & ~x253 & ~x278 & ~x310 & ~x336 & ~x364 & ~x366 & ~x391 & ~x393 & ~x394 & ~x481 & ~x504 & ~x560 & ~x687 & ~x701 & ~x703 & ~x727 & ~x747 & ~x758 & ~x771;
assign c137 = ~x10 & ~x22 & ~x32 & ~x33 & ~x40 & ~x44 & ~x49 & ~x50 & ~x59 & ~x61 & ~x67 & ~x69 & ~x70 & ~x71 & ~x78 & ~x79 & ~x85 & ~x90 & ~x92 & ~x95 & ~x96 & ~x100 & ~x104 & ~x106 & ~x107 & ~x109 & ~x111 & ~x121 & ~x133 & ~x134 & ~x138 & ~x144 & ~x146 & ~x161 & ~x164 & ~x187 & ~x188 & ~x190 & ~x200 & ~x223 & ~x228 & ~x229 & ~x279 & ~x307 & ~x310 & ~x334 & ~x336 & ~x338 & ~x360 & ~x361 & ~x366 & ~x367 & ~x368 & ~x391 & ~x394 & ~x395 & ~x414 & ~x415 & ~x416 & ~x417 & ~x421 & ~x422 & ~x445 & ~x447 & ~x449 & ~x450 & ~x468 & ~x469 & ~x470 & ~x473 & ~x474 & ~x478 & ~x486 & ~x487 & ~x502 & ~x507 & ~x523 & ~x529 & ~x532 & ~x557 & ~x561 & ~x579 & ~x580 & ~x591 & ~x605 & ~x615 & ~x617 & ~x619 & ~x644 & ~x647 & ~x665 & ~x666 & ~x669 & ~x675 & ~x690 & ~x693 & ~x698 & ~x701 & ~x718 & ~x719 & ~x721 & ~x725 & ~x727 & ~x729 & ~x745 & ~x748 & ~x749 & ~x754 & ~x755 & ~x757 & ~x760 & ~x761 & ~x763 & ~x772 & ~x775 & ~x776 & ~x777 & ~x778 & ~x781 & ~x783;
assign c139 =  x356 &  x381 &  x382 & ~x1 & ~x3 & ~x8 & ~x11 & ~x26 & ~x33 & ~x38 & ~x53 & ~x81 & ~x88 & ~x106 & ~x110 & ~x142 & ~x143 & ~x225 & ~x448 & ~x535 & ~x590 & ~x615 & ~x671 & ~x740 & ~x779;
assign c141 = ~x2 & ~x5 & ~x7 & ~x15 & ~x16 & ~x17 & ~x18 & ~x19 & ~x20 & ~x21 & ~x24 & ~x25 & ~x27 & ~x32 & ~x33 & ~x34 & ~x38 & ~x41 & ~x42 & ~x46 & ~x47 & ~x48 & ~x50 & ~x52 & ~x58 & ~x67 & ~x72 & ~x79 & ~x85 & ~x100 & ~x111 & ~x115 & ~x117 & ~x134 & ~x136 & ~x141 & ~x169 & ~x198 & ~x247 & ~x248 & ~x250 & ~x251 & ~x279 & ~x307 & ~x364 & ~x394 & ~x420 & ~x450 & ~x452 & ~x460 & ~x461 & ~x473 & ~x475 & ~x477 & ~x478 & ~x490 & ~x491 & ~x504 & ~x506 & ~x529 & ~x530 & ~x531 & ~x532 & ~x537 & ~x560 & ~x561 & ~x562 & ~x566 & ~x584 & ~x615 & ~x616 & ~x640 & ~x641 & ~x646 & ~x670 & ~x671 & ~x680 & ~x682 & ~x695 & ~x701 & ~x704 & ~x707 & ~x708 & ~x713 & ~x732 & ~x737 & ~x741 & ~x757 & ~x758 & ~x763 & ~x770 & ~x777 & ~x778 & ~x780 & ~x783;
assign c143 =  x408 & ~x5 & ~x24 & ~x36 & ~x46 & ~x61 & ~x63 & ~x69 & ~x70 & ~x71 & ~x80 & ~x84 & ~x110 & ~x137 & ~x140 & ~x195 & ~x200 & ~x201 & ~x233 & ~x251 & ~x311 & ~x314 & ~x324 & ~x340 & ~x358 & ~x371 & ~x391 & ~x417 & ~x418 & ~x424 & ~x445 & ~x447 & ~x449 & ~x450 & ~x454 & ~x471 & ~x474 & ~x499 & ~x500 & ~x502 & ~x506 & ~x535 & ~x582 & ~x588 & ~x617 & ~x646 & ~x648 & ~x661 & ~x667 & ~x669 & ~x671 & ~x724 & ~x729 & ~x731 & ~x734 & ~x740 & ~x741 & ~x750 & ~x752 & ~x757 & ~x765 & ~x766 & ~x781;
assign c145 =  x409 & ~x22 & ~x41 & ~x58 & ~x73 & ~x74 & ~x83 & ~x114 & ~x129 & ~x265 & ~x271 & ~x307 & ~x364 & ~x388 & ~x499 & ~x506 & ~x560 & ~x621 & ~x714 & ~x753;
assign c147 =  x521 & ~x0 & ~x1 & ~x9 & ~x14 & ~x16 & ~x17 & ~x22 & ~x24 & ~x34 & ~x43 & ~x45 & ~x50 & ~x60 & ~x64 & ~x67 & ~x68 & ~x73 & ~x78 & ~x79 & ~x82 & ~x85 & ~x95 & ~x97 & ~x99 & ~x105 & ~x109 & ~x113 & ~x136 & ~x142 & ~x148 & ~x165 & ~x168 & ~x169 & ~x197 & ~x224 & ~x250 & ~x251 & ~x278 & ~x282 & ~x307 & ~x361 & ~x362 & ~x390 & ~x393 & ~x416 & ~x417 & ~x420 & ~x445 & ~x490 & ~x506 & ~x528 & ~x530 & ~x531 & ~x553 & ~x557 & ~x584 & ~x608 & ~x610 & ~x636 & ~x638 & ~x645 & ~x664 & ~x665 & ~x674 & ~x675 & ~x694 & ~x698 & ~x703 & ~x724 & ~x727 & ~x729 & ~x730 & ~x737 & ~x740 & ~x742 & ~x750 & ~x753 & ~x754 & ~x761 & ~x766 & ~x767 & ~x771;
assign c149 =  x184 & ~x18 & ~x21 & ~x29 & ~x31 & ~x33 & ~x56 & ~x77 & ~x89 & ~x99 & ~x105 & ~x106 & ~x229 & ~x295 & ~x309 & ~x310 & ~x315 & ~x368 & ~x417 & ~x451 & ~x453 & ~x482 & ~x504 & ~x505 & ~x527 & ~x590 & ~x607 & ~x615 & ~x616 & ~x634 & ~x670 & ~x694 & ~x698 & ~x727 & ~x740 & ~x743;
assign c151 =  x151 &  x153 &  x178 & ~x0 & ~x15 & ~x24 & ~x28 & ~x39 & ~x43 & ~x51 & ~x56 & ~x69 & ~x85 & ~x87 & ~x88 & ~x90 & ~x94 & ~x100 & ~x102 & ~x105 & ~x115 & ~x116 & ~x133 & ~x143 & ~x193 & ~x197 & ~x252 & ~x279 & ~x305 & ~x306 & ~x337 & ~x365 & ~x474 & ~x478 & ~x503 & ~x504 & ~x533 & ~x558 & ~x587 & ~x589 & ~x593 & ~x621 & ~x672 & ~x692 & ~x746 & ~x764 & ~x780 & ~x783;
assign c153 =  x604 & ~x5 & ~x17 & ~x27 & ~x31 & ~x47 & ~x58 & ~x65 & ~x82 & ~x84 & ~x87 & ~x113 & ~x136 & ~x165 & ~x193 & ~x220 & ~x225 & ~x277 & ~x279 & ~x305 & ~x306 & ~x336 & ~x365 & ~x366 & ~x476 & ~x492 & ~x502 & ~x518 & ~x519 & ~x560 & ~x562 & ~x616 & ~x641 & ~x644 & ~x671 & ~x675 & ~x678 & ~x689 & ~x696 & ~x745 & ~x754 & ~x755 & ~x758 & ~x781;
assign c155 =  x442 & ~x13;
assign c157 =  x488 &  x550 & ~x25 & ~x26 & ~x41 & ~x42 & ~x56 & ~x60 & ~x61 & ~x72 & ~x73 & ~x74 & ~x77 & ~x107 & ~x112 & ~x114 & ~x115 & ~x141 & ~x171 & ~x194 & ~x197 & ~x309 & ~x311 & ~x422 & ~x559 & ~x562 & ~x586 & ~x587 & ~x642 & ~x643 & ~x666 & ~x672 & ~x673 & ~x681 & ~x696 & ~x706 & ~x707 & ~x728 & ~x762 & ~x767 & ~x778 & ~x779 & ~x780;
assign c159 =  x210 & ~x9 & ~x45 & ~x74 & ~x99 & ~x118 & ~x126 & ~x127 & ~x128 & ~x139 & ~x140 & ~x171 & ~x220 & ~x292 & ~x364 & ~x384 & ~x398 & ~x400 & ~x416 & ~x424 & ~x429 & ~x441 & ~x445 & ~x458 & ~x472 & ~x474 & ~x532 & ~x593 & ~x669 & ~x677 & ~x721 & ~x725 & ~x727 & ~x730 & ~x782;
assign c161 =  x154 &  x298 & ~x9 & ~x26 & ~x49 & ~x67 & ~x87 & ~x103 & ~x105 & ~x106 & ~x108 & ~x109 & ~x113 & ~x114 & ~x169 & ~x171 & ~x172 & ~x196 & ~x226 & ~x250 & ~x280 & ~x308 & ~x331 & ~x332 & ~x334 & ~x336 & ~x364 & ~x391 & ~x425 & ~x447 & ~x616 & ~x672 & ~x698 & ~x709 & ~x713 & ~x716 & ~x742 & ~x743 & ~x756 & ~x763 & ~x781;
assign c163 =  x155 & ~x7 & ~x12 & ~x15 & ~x16 & ~x17 & ~x37 & ~x44 & ~x48 & ~x51 & ~x55 & ~x64 & ~x72 & ~x75 & ~x78 & ~x87 & ~x91 & ~x102 & ~x106 & ~x107 & ~x112 & ~x117 & ~x118 & ~x119 & ~x133 & ~x135 & ~x139 & ~x141 & ~x164 & ~x169 & ~x171 & ~x173 & ~x191 & ~x193 & ~x194 & ~x195 & ~x197 & ~x219 & ~x220 & ~x221 & ~x223 & ~x225 & ~x228 & ~x238 & ~x249 & ~x303 & ~x310 & ~x313 & ~x329 & ~x330 & ~x365 & ~x369 & ~x385 & ~x395 & ~x398 & ~x399 & ~x421 & ~x427 & ~x443 & ~x480 & ~x501 & ~x528 & ~x534 & ~x537 & ~x560 & ~x561 & ~x588 & ~x645 & ~x649 & ~x674 & ~x675 & ~x677 & ~x681 & ~x696 & ~x699 & ~x700 & ~x706 & ~x707 & ~x713 & ~x714 & ~x717 & ~x720 & ~x721 & ~x723 & ~x726 & ~x728 & ~x737 & ~x749 & ~x756 & ~x762 & ~x772 & ~x774;
assign c165 =  x374 &  x403 & ~x14 & ~x29 & ~x53 & ~x66 & ~x114 & ~x198 & ~x253 & ~x311 & ~x312 & ~x334 & ~x419 & ~x445 & ~x456 & ~x512 & ~x532 & ~x556 & ~x583 & ~x665 & ~x689 & ~x737;
assign c167 =  x182 & ~x6 & ~x7 & ~x9 & ~x13 & ~x19 & ~x27 & ~x35 & ~x37 & ~x56 & ~x60 & ~x61 & ~x82 & ~x127 & ~x170 & ~x171 & ~x194 & ~x198 & ~x251 & ~x276 & ~x278 & ~x311 & ~x312 & ~x334 & ~x336 & ~x368 & ~x419 & ~x475 & ~x477 & ~x518 & ~x616 & ~x646 & ~x698 & ~x724 & ~x730 & ~x731 & ~x742 & ~x745 & ~x750 & ~x762 & ~x766 & ~x769 & ~x772;
assign c169 =  x511 & ~x2 & ~x3 & ~x5 & ~x10 & ~x14 & ~x15 & ~x16 & ~x20 & ~x22 & ~x25 & ~x26 & ~x35 & ~x43 & ~x46 & ~x51 & ~x55 & ~x58 & ~x61 & ~x62 & ~x63 & ~x66 & ~x67 & ~x68 & ~x82 & ~x83 & ~x86 & ~x88 & ~x89 & ~x90 & ~x91 & ~x113 & ~x115 & ~x145 & ~x147 & ~x168 & ~x171 & ~x173 & ~x200 & ~x224 & ~x227 & ~x256 & ~x258 & ~x280 & ~x281 & ~x368 & ~x392 & ~x395 & ~x421 & ~x423 & ~x450 & ~x474 & ~x476 & ~x479 & ~x504 & ~x507 & ~x508 & ~x529 & ~x533 & ~x535 & ~x559 & ~x615 & ~x619 & ~x641 & ~x644 & ~x645 & ~x646 & ~x650 & ~x670 & ~x672 & ~x673 & ~x680 & ~x684 & ~x685 & ~x686 & ~x697 & ~x702 & ~x703 & ~x710 & ~x713 & ~x719 & ~x728 & ~x735 & ~x741 & ~x746 & ~x748 & ~x753 & ~x759 & ~x760 & ~x761 & ~x767 & ~x768 & ~x770 & ~x780 & ~x783;
assign c171 = ~x1 & ~x21 & ~x45 & ~x49 & ~x51 & ~x88 & ~x93 & ~x116 & ~x138 & ~x140 & ~x167 & ~x168 & ~x194 & ~x306 & ~x340 & ~x419 & ~x421 & ~x435 & ~x475 & ~x505 & ~x515 & ~x529 & ~x589 & ~x618 & ~x715 & ~x729 & ~x731 & ~x732 & ~x776 & ~x780;
assign c173 =  x454 & ~x3 & ~x4 & ~x26 & ~x83 & ~x282 & ~x333 & ~x446 & ~x505 & ~x644 & ~x649;
assign c175 = ~x4 & ~x6 & ~x10 & ~x16 & ~x31 & ~x35 & ~x36 & ~x38 & ~x58 & ~x68 & ~x74 & ~x83 & ~x97 & ~x110 & ~x141 & ~x155 & ~x198 & ~x223 & ~x248 & ~x254 & ~x279 & ~x338 & ~x363 & ~x368 & ~x393 & ~x396 & ~x405 & ~x406 & ~x421 & ~x448 & ~x481 & ~x502 & ~x509 & ~x561 & ~x585 & ~x587 & ~x598 & ~x615 & ~x626 & ~x671 & ~x697 & ~x700 & ~x733 & ~x735 & ~x736 & ~x756 & ~x762 & ~x767 & ~x776 & ~x777;
assign c177 =  x486 &  x542 &  x570 & ~x13 & ~x15 & ~x19 & ~x23 & ~x61 & ~x77 & ~x83 & ~x110 & ~x112 & ~x165 & ~x167 & ~x168 & ~x194 & ~x199 & ~x221 & ~x224 & ~x247 & ~x252 & ~x276 & ~x278 & ~x286 & ~x329 & ~x332 & ~x336 & ~x337 & ~x355 & ~x362 & ~x382 & ~x388 & ~x396 & ~x411 & ~x413 & ~x420 & ~x425 & ~x475 & ~x615 & ~x619 & ~x640 & ~x647 & ~x652 & ~x653 & ~x654 & ~x670 & ~x674 & ~x700 & ~x710 & ~x750 & ~x756 & ~x763 & ~x782;
assign c179 =  x258 & ~x14 & ~x17 & ~x26 & ~x49 & ~x73 & ~x78 & ~x88 & ~x99 & ~x112 & ~x127 & ~x129 & ~x139 & ~x140 & ~x158 & ~x278 & ~x307 & ~x309 & ~x422 & ~x475 & ~x480 & ~x503 & ~x529 & ~x560 & ~x561 & ~x563 & ~x585 & ~x594 & ~x617 & ~x641 & ~x668 & ~x733 & ~x752 & ~x757 & ~x767 & ~x770 & ~x778 & ~x780;
assign c181 =  x263 & ~x15 & ~x16 & ~x22 & ~x25 & ~x26 & ~x54 & ~x57 & ~x75 & ~x81 & ~x86 & ~x89 & ~x107 & ~x119 & ~x125 & ~x127 & ~x129 & ~x137 & ~x141 & ~x146 & ~x150 & ~x151 & ~x154 & ~x157 & ~x168 & ~x224 & ~x278 & ~x283 & ~x360 & ~x394 & ~x417 & ~x424 & ~x444 & ~x450 & ~x455 & ~x471 & ~x474 & ~x477 & ~x482 & ~x483 & ~x528 & ~x533 & ~x538 & ~x554 & ~x564 & ~x568 & ~x589 & ~x616 & ~x619 & ~x637 & ~x670 & ~x673 & ~x691 & ~x701 & ~x721 & ~x723 & ~x737 & ~x765 & ~x775;
assign c183 =  x520 & ~x0 & ~x2 & ~x6 & ~x8 & ~x11 & ~x23 & ~x41 & ~x54 & ~x56 & ~x58 & ~x61 & ~x76 & ~x169 & ~x191 & ~x193 & ~x200 & ~x227 & ~x281 & ~x293 & ~x301 & ~x309 & ~x313 & ~x332 & ~x362 & ~x363 & ~x563 & ~x588 & ~x591 & ~x594 & ~x607 & ~x615 & ~x616 & ~x620 & ~x634 & ~x648 & ~x670 & ~x673 & ~x677 & ~x702 & ~x704 & ~x706 & ~x709 & ~x728 & ~x730 & ~x735 & ~x739 & ~x755 & ~x762 & ~x765 & ~x770 & ~x776;
assign c185 = ~x36 & ~x99 & ~x128 & ~x291 & ~x391 & ~x450 & ~x771 & ~x772;
assign c187 =  x402 & ~x0 & ~x4 & ~x7 & ~x9 & ~x19 & ~x22 & ~x28 & ~x39 & ~x40 & ~x41 & ~x45 & ~x46 & ~x47 & ~x49 & ~x51 & ~x52 & ~x58 & ~x62 & ~x64 & ~x66 & ~x77 & ~x80 & ~x83 & ~x88 & ~x114 & ~x115 & ~x117 & ~x139 & ~x197 & ~x199 & ~x201 & ~x226 & ~x250 & ~x251 & ~x253 & ~x279 & ~x321 & ~x363 & ~x368 & ~x419 & ~x421 & ~x446 & ~x449 & ~x473 & ~x503 & ~x529 & ~x530 & ~x533 & ~x557 & ~x562 & ~x585 & ~x591 & ~x614 & ~x615 & ~x617 & ~x619 & ~x642 & ~x647 & ~x648 & ~x672 & ~x673 & ~x702 & ~x725 & ~x732 & ~x742 & ~x748 & ~x755 & ~x757 & ~x768;
assign c189 =  x316 & ~x0 & ~x1 & ~x5 & ~x8 & ~x11 & ~x18 & ~x21 & ~x29 & ~x33 & ~x36 & ~x40 & ~x41 & ~x47 & ~x51 & ~x57 & ~x58 & ~x59 & ~x60 & ~x63 & ~x67 & ~x69 & ~x71 & ~x77 & ~x82 & ~x84 & ~x92 & ~x101 & ~x105 & ~x110 & ~x111 & ~x112 & ~x121 & ~x124 & ~x125 & ~x126 & ~x127 & ~x134 & ~x141 & ~x145 & ~x152 & ~x164 & ~x169 & ~x198 & ~x199 & ~x279 & ~x332 & ~x336 & ~x361 & ~x391 & ~x394 & ~x419 & ~x420 & ~x450 & ~x475 & ~x476 & ~x478 & ~x500 & ~x501 & ~x504 & ~x507 & ~x531 & ~x536 & ~x557 & ~x564 & ~x565 & ~x584 & ~x585 & ~x587 & ~x593 & ~x594 & ~x618 & ~x640 & ~x642 & ~x644 & ~x645 & ~x647 & ~x669 & ~x671 & ~x674 & ~x675 & ~x677 & ~x697 & ~x701 & ~x702 & ~x707 & ~x708 & ~x723 & ~x727 & ~x751 & ~x752 & ~x754 & ~x756 & ~x759 & ~x764 & ~x766 & ~x768 & ~x776 & ~x777 & ~x779 & ~x782;
assign c191 =  x438 & ~x5 & ~x12 & ~x14 & ~x18 & ~x19 & ~x21 & ~x22 & ~x23 & ~x26 & ~x42 & ~x48 & ~x49 & ~x50 & ~x64 & ~x65 & ~x69 & ~x87 & ~x89 & ~x140 & ~x144 & ~x196 & ~x198 & ~x220 & ~x225 & ~x282 & ~x307 & ~x309 & ~x361 & ~x362 & ~x363 & ~x366 & ~x394 & ~x395 & ~x448 & ~x473 & ~x477 & ~x500 & ~x533 & ~x555 & ~x559 & ~x561 & ~x615 & ~x641 & ~x646 & ~x655 & ~x658 & ~x684 & ~x700 & ~x710 & ~x712 & ~x714 & ~x726 & ~x727 & ~x730 & ~x734 & ~x735 & ~x739 & ~x741 & ~x744 & ~x763 & ~x767 & ~x773 & ~x780;
assign c193 =  x459 &  x492 & ~x26 & ~x29 & ~x33 & ~x37 & ~x52 & ~x73 & ~x92 & ~x174 & ~x175 & ~x222 & ~x307 & ~x311 & ~x332 & ~x337 & ~x367 & ~x382 & ~x411 & ~x420 & ~x423 & ~x502 & ~x531 & ~x559 & ~x592 & ~x593 & ~x616 & ~x648 & ~x669 & ~x698 & ~x700 & ~x743 & ~x769 & ~x773 & ~x781;
assign c195 =  x208 &  x326 & ~x3 & ~x7 & ~x10 & ~x19 & ~x27 & ~x30 & ~x43 & ~x65 & ~x85 & ~x115 & ~x135 & ~x139 & ~x142 & ~x282 & ~x308 & ~x334 & ~x337 & ~x339 & ~x396 & ~x449 & ~x475 & ~x504 & ~x531 & ~x532 & ~x556 & ~x617 & ~x673 & ~x693 & ~x703 & ~x758 & ~x764 & ~x765;
assign c197 =  x487 & ~x1 & ~x7 & ~x16 & ~x20 & ~x28 & ~x34 & ~x38 & ~x50 & ~x54 & ~x59 & ~x69 & ~x77 & ~x81 & ~x83 & ~x88 & ~x106 & ~x111 & ~x165 & ~x191 & ~x222 & ~x252 & ~x254 & ~x256 & ~x279 & ~x281 & ~x282 & ~x307 & ~x310 & ~x334 & ~x337 & ~x338 & ~x361 & ~x393 & ~x450 & ~x479 & ~x481 & ~x502 & ~x505 & ~x506 & ~x507 & ~x531 & ~x535 & ~x617 & ~x642 & ~x644 & ~x667 & ~x669 & ~x670 & ~x675 & ~x681 & ~x696 & ~x697 & ~x709 & ~x719 & ~x721 & ~x726 & ~x731 & ~x736 & ~x738 & ~x740 & ~x741 & ~x743 & ~x745 & ~x746 & ~x747 & ~x750 & ~x754 & ~x762 & ~x777 & ~x778;
assign c199 =  x525 & ~x4 & ~x5 & ~x22 & ~x23 & ~x26 & ~x34 & ~x38 & ~x42 & ~x44 & ~x54 & ~x57 & ~x58 & ~x59 & ~x62 & ~x64 & ~x72 & ~x79 & ~x83 & ~x86 & ~x87 & ~x88 & ~x91 & ~x113 & ~x117 & ~x135 & ~x139 & ~x142 & ~x172 & ~x191 & ~x221 & ~x223 & ~x226 & ~x249 & ~x251 & ~x305 & ~x310 & ~x338 & ~x366 & ~x391 & ~x421 & ~x447 & ~x475 & ~x478 & ~x532 & ~x561 & ~x562 & ~x563 & ~x586 & ~x589 & ~x615 & ~x616 & ~x617 & ~x619 & ~x643 & ~x647 & ~x669 & ~x672 & ~x673 & ~x675 & ~x700 & ~x703 & ~x706 & ~x718 & ~x722 & ~x728 & ~x730 & ~x733 & ~x735 & ~x739 & ~x745 & ~x749 & ~x751 & ~x752 & ~x753 & ~x754 & ~x755 & ~x758 & ~x759 & ~x764 & ~x768 & ~x769 & ~x770 & ~x772 & ~x773 & ~x778 & ~x779 & ~x783;
assign c1101 =  x493 & ~x1 & ~x15 & ~x25 & ~x44 & ~x46 & ~x82 & ~x144 & ~x196 & ~x305 & ~x306 & ~x320 & ~x334 & ~x340 & ~x366 & ~x418 & ~x421 & ~x447 & ~x478 & ~x503 & ~x557 & ~x602 & ~x646 & ~x669 & ~x674 & ~x679 & ~x694 & ~x728 & ~x764;
assign c1103 =  x440 & ~x0 & ~x15 & ~x18 & ~x22 & ~x32 & ~x37 & ~x43 & ~x49 & ~x53 & ~x82 & ~x87 & ~x88 & ~x90 & ~x91 & ~x92 & ~x112 & ~x114 & ~x118 & ~x136 & ~x144 & ~x166 & ~x167 & ~x193 & ~x222 & ~x223 & ~x279 & ~x305 & ~x306 & ~x333 & ~x336 & ~x361 & ~x418 & ~x420 & ~x473 & ~x501 & ~x502 & ~x530 & ~x533 & ~x584 & ~x587 & ~x612 & ~x614 & ~x615 & ~x643 & ~x645 & ~x647 & ~x667 & ~x673 & ~x675 & ~x676 & ~x680 & ~x696 & ~x698 & ~x699 & ~x705 & ~x706 & ~x723 & ~x725 & ~x727 & ~x735 & ~x755 & ~x757 & ~x759 & ~x760 & ~x762 & ~x767 & ~x775 & ~x780 & ~x781;
assign c1105 = ~x11 & ~x12 & ~x13 & ~x14 & ~x17 & ~x18 & ~x20 & ~x23 & ~x25 & ~x26 & ~x28 & ~x40 & ~x42 & ~x45 & ~x46 & ~x48 & ~x49 & ~x51 & ~x53 & ~x57 & ~x59 & ~x65 & ~x73 & ~x76 & ~x79 & ~x80 & ~x81 & ~x82 & ~x83 & ~x84 & ~x86 & ~x90 & ~x91 & ~x92 & ~x94 & ~x96 & ~x97 & ~x98 & ~x99 & ~x100 & ~x106 & ~x110 & ~x114 & ~x115 & ~x136 & ~x138 & ~x139 & ~x140 & ~x141 & ~x165 & ~x167 & ~x169 & ~x170 & ~x194 & ~x195 & ~x201 & ~x224 & ~x230 & ~x248 & ~x249 & ~x252 & ~x272 & ~x280 & ~x306 & ~x307 & ~x311 & ~x328 & ~x330 & ~x337 & ~x363 & ~x386 & ~x389 & ~x390 & ~x391 & ~x392 & ~x417 & ~x420 & ~x422 & ~x471 & ~x474 & ~x475 & ~x479 & ~x489 & ~x490 & ~x499 & ~x505 & ~x506 & ~x513 & ~x514 & ~x516 & ~x529 & ~x535 & ~x537 & ~x553 & ~x558 & ~x589 & ~x611 & ~x612 & ~x613 & ~x615 & ~x617 & ~x620 & ~x640 & ~x641 & ~x643 & ~x647 & ~x665 & ~x670 & ~x671 & ~x673 & ~x676 & ~x694 & ~x701 & ~x705 & ~x707 & ~x708 & ~x722 & ~x723 & ~x727 & ~x728 & ~x732 & ~x736 & ~x743 & ~x750 & ~x751 & ~x754 & ~x757 & ~x758 & ~x768 & ~x770 & ~x775 & ~x781 & ~x783;
assign c1107 =  x407 & ~x23 & ~x32 & ~x37 & ~x45 & ~x47 & ~x56 & ~x61 & ~x65 & ~x67 & ~x71 & ~x76 & ~x104 & ~x111 & ~x113 & ~x132 & ~x159 & ~x165 & ~x218 & ~x223 & ~x225 & ~x275 & ~x278 & ~x280 & ~x303 & ~x321 & ~x322 & ~x330 & ~x335 & ~x340 & ~x422 & ~x507 & ~x530 & ~x532 & ~x559 & ~x595 & ~x598 & ~x650 & ~x729 & ~x732 & ~x735 & ~x753 & ~x754 & ~x765;
assign c1109 =  x156 &  x188 & ~x9 & ~x15 & ~x29 & ~x41 & ~x61 & ~x71 & ~x78 & ~x106 & ~x335 & ~x366 & ~x588 & ~x644 & ~x763;
assign c1111 =  x686 & ~x12 & ~x23 & ~x37 & ~x38 & ~x42 & ~x46 & ~x48 & ~x69 & ~x76 & ~x77 & ~x86 & ~x103 & ~x104 & ~x108 & ~x109 & ~x110 & ~x121 & ~x122 & ~x123 & ~x126 & ~x128 & ~x132 & ~x135 & ~x143 & ~x165 & ~x197 & ~x250 & ~x332 & ~x334 & ~x364 & ~x365 & ~x389 & ~x392 & ~x393 & ~x394 & ~x418 & ~x421 & ~x445 & ~x451 & ~x454 & ~x456 & ~x504 & ~x509 & ~x514 & ~x535 & ~x545 & ~x573 & ~x586 & ~x618 & ~x675 & ~x676 & ~x693 & ~x700 & ~x705 & ~x727 & ~x739 & ~x747 & ~x765 & ~x768 & ~x774 & ~x777;
assign c1113 =  x511 &  x540 & ~x0 & ~x7 & ~x8 & ~x14 & ~x19 & ~x25 & ~x45 & ~x46 & ~x53 & ~x55 & ~x56 & ~x74 & ~x75 & ~x80 & ~x82 & ~x83 & ~x84 & ~x90 & ~x110 & ~x116 & ~x136 & ~x139 & ~x142 & ~x173 & ~x251 & ~x254 & ~x278 & ~x281 & ~x282 & ~x310 & ~x336 & ~x338 & ~x339 & ~x368 & ~x392 & ~x394 & ~x395 & ~x419 & ~x422 & ~x423 & ~x504 & ~x531 & ~x532 & ~x560 & ~x587 & ~x615 & ~x616 & ~x639 & ~x641 & ~x643 & ~x644 & ~x649 & ~x666 & ~x671 & ~x674 & ~x695 & ~x702 & ~x704 & ~x707 & ~x708 & ~x710 & ~x713 & ~x717 & ~x726 & ~x731 & ~x738 & ~x739 & ~x753 & ~x755 & ~x769 & ~x777 & ~x781 & ~x783;
assign c1115 = ~x13 & ~x16 & ~x42 & ~x47 & ~x58 & ~x61 & ~x72 & ~x93 & ~x94 & ~x97 & ~x111 & ~x112 & ~x113 & ~x119 & ~x121 & ~x125 & ~x129 & ~x139 & ~x142 & ~x143 & ~x170 & ~x171 & ~x226 & ~x255 & ~x307 & ~x308 & ~x364 & ~x390 & ~x407 & ~x423 & ~x424 & ~x447 & ~x479 & ~x499 & ~x504 & ~x506 & ~x528 & ~x529 & ~x531 & ~x584 & ~x592 & ~x613 & ~x614 & ~x638 & ~x642 & ~x670 & ~x671 & ~x672 & ~x678 & ~x693 & ~x695 & ~x697 & ~x698 & ~x701 & ~x706 & ~x723 & ~x725 & ~x730 & ~x736 & ~x737 & ~x739 & ~x754 & ~x755 & ~x756 & ~x763 & ~x764 & ~x768 & ~x775 & ~x777 & ~x779 & ~x783;
assign c1117 =  x463 & ~x18 & ~x42 & ~x44 & ~x74 & ~x77 & ~x83 & ~x92 & ~x102 & ~x108 & ~x131 & ~x141 & ~x144 & ~x151 & ~x176 & ~x281 & ~x351 & ~x396 & ~x417 & ~x444 & ~x449 & ~x473 & ~x504 & ~x505 & ~x533 & ~x635 & ~x641 & ~x698 & ~x712 & ~x757 & ~x779;
assign c1119 =  x208 & ~x13 & ~x30 & ~x59 & ~x75 & ~x80 & ~x83 & ~x91 & ~x127 & ~x134 & ~x160 & ~x224 & ~x293 & ~x336 & ~x413 & ~x420 & ~x526 & ~x562 & ~x570 & ~x587 & ~x596 & ~x616 & ~x625 & ~x645 & ~x723;
assign c1121 = ~x11 & ~x14 & ~x18 & ~x22 & ~x23 & ~x24 & ~x29 & ~x40 & ~x51 & ~x53 & ~x61 & ~x75 & ~x80 & ~x81 & ~x83 & ~x86 & ~x95 & ~x109 & ~x110 & ~x113 & ~x120 & ~x122 & ~x139 & ~x140 & ~x146 & ~x147 & ~x163 & ~x166 & ~x167 & ~x177 & ~x199 & ~x226 & ~x279 & ~x285 & ~x302 & ~x309 & ~x311 & ~x313 & ~x322 & ~x330 & ~x333 & ~x337 & ~x356 & ~x384 & ~x397 & ~x420 & ~x421 & ~x422 & ~x423 & ~x446 & ~x449 & ~x476 & ~x478 & ~x499 & ~x507 & ~x534 & ~x538 & ~x558 & ~x560 & ~x564 & ~x584 & ~x588 & ~x591 & ~x609 & ~x618 & ~x624 & ~x632 & ~x640 & ~x650 & ~x662 & ~x663 & ~x666 & ~x703 & ~x728 & ~x732 & ~x735 & ~x754 & ~x765 & ~x766 & ~x772 & ~x773 & ~x776 & ~x779;
assign c1123 =  x543 &  x578 & ~x59 & ~x74 & ~x163 & ~x293 & ~x338 & ~x502 & ~x558 & ~x642 & ~x647 & ~x683 & ~x716 & ~x768;
assign c1125 =  x523 & ~x1 & ~x2 & ~x13 & ~x36 & ~x58 & ~x72 & ~x78 & ~x113 & ~x195 & ~x221 & ~x252 & ~x280 & ~x282 & ~x292 & ~x293 & ~x334 & ~x395 & ~x475 & ~x479 & ~x560 & ~x615 & ~x643 & ~x668 & ~x669 & ~x674 & ~x677 & ~x712 & ~x739 & ~x746 & ~x757 & ~x768 & ~x771 & ~x773;
assign c1127 =  x494 & ~x8 & ~x14 & ~x18 & ~x26 & ~x34 & ~x40 & ~x43 & ~x50 & ~x57 & ~x62 & ~x70 & ~x71 & ~x72 & ~x74 & ~x110 & ~x141 & ~x222 & ~x236 & ~x252 & ~x279 & ~x337 & ~x341 & ~x387 & ~x392 & ~x422 & ~x450 & ~x451 & ~x478 & ~x479 & ~x502 & ~x643 & ~x645 & ~x665 & ~x666 & ~x717 & ~x724 & ~x726 & ~x752 & ~x783;
assign c1129 =  x291 & ~x14 & ~x27 & ~x28 & ~x36 & ~x49 & ~x54 & ~x56 & ~x77 & ~x84 & ~x85 & ~x117 & ~x122 & ~x135 & ~x145 & ~x167 & ~x171 & ~x174 & ~x179 & ~x201 & ~x310 & ~x335 & ~x393 & ~x394 & ~x418 & ~x420 & ~x444 & ~x477 & ~x503 & ~x533 & ~x576 & ~x603 & ~x631 & ~x661 & ~x728 & ~x746 & ~x766 & ~x767;
assign c1131 =  x657 &  x658 & ~x26 & ~x43 & ~x166 & ~x223 & ~x277 & ~x303 & ~x359 & ~x392 & ~x420 & ~x428 & ~x453 & ~x546 & ~x562 & ~x612 & ~x617 & ~x696;
assign c1133 =  x654 &  x656 & ~x5 & ~x7 & ~x20 & ~x38 & ~x78 & ~x102 & ~x197 & ~x253 & ~x306 & ~x307 & ~x308 & ~x367 & ~x392 & ~x422 & ~x476 & ~x477 & ~x502 & ~x571 & ~x619 & ~x621 & ~x668 & ~x674 & ~x703 & ~x704 & ~x714 & ~x734 & ~x752 & ~x760 & ~x762 & ~x763 & ~x765 & ~x767 & ~x768;
assign c1135 =  x577 & ~x0 & ~x4 & ~x8 & ~x43 & ~x46 & ~x58 & ~x73 & ~x80 & ~x86 & ~x88 & ~x107 & ~x115 & ~x140 & ~x141 & ~x142 & ~x143 & ~x166 & ~x219 & ~x223 & ~x253 & ~x277 & ~x332 & ~x333 & ~x361 & ~x395 & ~x407 & ~x423 & ~x434 & ~x475 & ~x478 & ~x506 & ~x507 & ~x533 & ~x534 & ~x590 & ~x592 & ~x593 & ~x615 & ~x620 & ~x644 & ~x648 & ~x649 & ~x669 & ~x674 & ~x679 & ~x700 & ~x702 & ~x703 & ~x704 & ~x711 & ~x727 & ~x729 & ~x759;
assign c1137 =  x156 & ~x1 & ~x2 & ~x28 & ~x42 & ~x44 & ~x50 & ~x58 & ~x63 & ~x72 & ~x76 & ~x97 & ~x104 & ~x112 & ~x115 & ~x146 & ~x166 & ~x169 & ~x229 & ~x240 & ~x276 & ~x313 & ~x331 & ~x337 & ~x358 & ~x364 & ~x388 & ~x390 & ~x394 & ~x395 & ~x397 & ~x449 & ~x526 & ~x639 & ~x643 & ~x674 & ~x713 & ~x720 & ~x721 & ~x729 & ~x730 & ~x732 & ~x744 & ~x755 & ~x759 & ~x776 & ~x779;
assign c1139 =  x407 &  x460 & ~x18 & ~x26 & ~x36 & ~x54 & ~x82 & ~x83 & ~x93 & ~x112 & ~x116 & ~x138 & ~x140 & ~x256 & ~x258 & ~x309 & ~x323 & ~x335 & ~x359 & ~x364 & ~x367 & ~x395 & ~x397 & ~x413 & ~x415 & ~x419 & ~x423 & ~x425 & ~x441 & ~x453 & ~x471 & ~x479 & ~x500 & ~x504 & ~x531 & ~x535 & ~x564 & ~x588 & ~x616 & ~x665 & ~x674 & ~x698 & ~x703 & ~x705 & ~x723 & ~x731 & ~x747 & ~x773 & ~x776;
assign c1141 =  x239 & ~x6 & ~x30 & ~x35 & ~x44 & ~x48 & ~x52 & ~x61 & ~x62 & ~x76 & ~x85 & ~x87 & ~x106 & ~x110 & ~x113 & ~x136 & ~x140 & ~x143 & ~x164 & ~x170 & ~x173 & ~x174 & ~x224 & ~x280 & ~x281 & ~x295 & ~x302 & ~x312 & ~x339 & ~x363 & ~x364 & ~x392 & ~x448 & ~x451 & ~x563 & ~x591 & ~x594 & ~x610 & ~x618 & ~x623 & ~x650 & ~x663 & ~x664 & ~x667 & ~x697 & ~x699 & ~x756 & ~x759 & ~x760 & ~x763 & ~x766 & ~x769 & ~x776;
assign c1143 =  x300 & ~x4 & ~x5 & ~x11 & ~x15 & ~x22 & ~x23 & ~x26 & ~x28 & ~x31 & ~x41 & ~x53 & ~x54 & ~x55 & ~x68 & ~x72 & ~x76 & ~x83 & ~x89 & ~x105 & ~x108 & ~x109 & ~x110 & ~x115 & ~x116 & ~x138 & ~x143 & ~x144 & ~x162 & ~x163 & ~x164 & ~x165 & ~x170 & ~x192 & ~x194 & ~x254 & ~x279 & ~x307 & ~x309 & ~x312 & ~x337 & ~x339 & ~x366 & ~x367 & ~x392 & ~x413 & ~x418 & ~x420 & ~x440 & ~x447 & ~x449 & ~x504 & ~x506 & ~x507 & ~x559 & ~x588 & ~x615 & ~x641 & ~x669 & ~x670 & ~x696 & ~x720 & ~x723 & ~x731 & ~x732 & ~x740 & ~x743 & ~x752 & ~x753 & ~x755 & ~x756 & ~x758 & ~x760 & ~x761 & ~x762 & ~x763 & ~x772 & ~x773 & ~x774 & ~x775;
assign c1145 =  x521 &  x549 & ~x60 & ~x62 & ~x140 & ~x179 & ~x205 & ~x207 & ~x208 & ~x234 & ~x343 & ~x362 & ~x418 & ~x445 & ~x446 & ~x530 & ~x560 & ~x663 & ~x674 & ~x683 & ~x684 & ~x702 & ~x704 & ~x726;
assign c1147 =  x154 &  x543 & ~x24 & ~x28 & ~x34 & ~x43 & ~x55 & ~x73 & ~x79 & ~x105 & ~x170 & ~x173 & ~x197 & ~x219 & ~x250 & ~x252 & ~x266 & ~x281 & ~x300 & ~x305 & ~x336 & ~x423 & ~x424 & ~x448 & ~x451 & ~x503 & ~x535 & ~x591 & ~x620 & ~x675 & ~x677 & ~x707 & ~x708 & ~x739 & ~x752 & ~x756 & ~x757 & ~x769 & ~x772 & ~x775;
assign c1149 =  x467 & ~x8 & ~x10 & ~x12 & ~x15 & ~x20 & ~x21 & ~x26 & ~x29 & ~x31 & ~x37 & ~x39 & ~x41 & ~x46 & ~x48 & ~x53 & ~x57 & ~x59 & ~x60 & ~x61 & ~x66 & ~x67 & ~x74 & ~x78 & ~x79 & ~x82 & ~x85 & ~x86 & ~x89 & ~x112 & ~x114 & ~x139 & ~x140 & ~x143 & ~x144 & ~x165 & ~x280 & ~x282 & ~x308 & ~x334 & ~x363 & ~x393 & ~x394 & ~x395 & ~x416 & ~x418 & ~x419 & ~x475 & ~x476 & ~x477 & ~x503 & ~x508 & ~x527 & ~x530 & ~x532 & ~x534 & ~x557 & ~x586 & ~x613 & ~x615 & ~x644 & ~x645 & ~x670 & ~x671 & ~x672 & ~x674 & ~x675 & ~x680 & ~x681 & ~x697 & ~x699 & ~x704 & ~x706 & ~x708 & ~x724 & ~x725 & ~x730 & ~x737 & ~x750 & ~x753 & ~x778 & ~x779 & ~x781 & ~x782;
assign c1151 =  x181 &  x214 & ~x17 & ~x45 & ~x58 & ~x72 & ~x80 & ~x96 & ~x104 & ~x107 & ~x112 & ~x121 & ~x227 & ~x419 & ~x530 & ~x670 & ~x723 & ~x741 & ~x743;
assign c1153 =  x543 & ~x24 & ~x37 & ~x74 & ~x75 & ~x79 & ~x90 & ~x117 & ~x143 & ~x144 & ~x169 & ~x171 & ~x276 & ~x277 & ~x305 & ~x311 & ~x322 & ~x323 & ~x333 & ~x390 & ~x420 & ~x421 & ~x445 & ~x503 & ~x505 & ~x534 & ~x591 & ~x613 & ~x615 & ~x645 & ~x672 & ~x716 & ~x754 & ~x762 & ~x763 & ~x767 & ~x773;
assign c1155 =  x317 & ~x41 & ~x52 & ~x56 & ~x75 & ~x78 & ~x96 & ~x99 & ~x120 & ~x123 & ~x125 & ~x127 & ~x134 & ~x147 & ~x228 & ~x307 & ~x308 & ~x367 & ~x369 & ~x397 & ~x418 & ~x424 & ~x449 & ~x477 & ~x479 & ~x535 & ~x555 & ~x596 & ~x620 & ~x622 & ~x623 & ~x639 & ~x674 & ~x721 & ~x771;
assign c1157 = ~x10 & ~x13 & ~x16 & ~x27 & ~x41 & ~x46 & ~x53 & ~x58 & ~x60 & ~x63 & ~x74 & ~x76 & ~x85 & ~x101 & ~x102 & ~x116 & ~x163 & ~x168 & ~x186 & ~x188 & ~x198 & ~x220 & ~x228 & ~x243 & ~x264 & ~x273 & ~x276 & ~x277 & ~x281 & ~x312 & ~x320 & ~x337 & ~x395 & ~x531 & ~x648 & ~x652 & ~x654 & ~x684 & ~x699 & ~x701 & ~x702 & ~x734 & ~x742 & ~x750 & ~x775 & ~x777;
assign c1159 =  x627 & ~x14 & ~x17 & ~x18 & ~x19 & ~x38 & ~x47 & ~x48 & ~x53 & ~x70 & ~x87 & ~x93 & ~x138 & ~x139 & ~x203 & ~x233 & ~x252 & ~x259 & ~x283 & ~x305 & ~x306 & ~x324 & ~x412 & ~x419 & ~x423 & ~x424 & ~x505 & ~x580 & ~x592 & ~x610 & ~x646 & ~x672 & ~x696 & ~x733 & ~x734 & ~x735 & ~x750 & ~x760 & ~x775;
assign c1161 = ~x1 & ~x5 & ~x11 & ~x14 & ~x20 & ~x48 & ~x60 & ~x76 & ~x78 & ~x88 & ~x93 & ~x114 & ~x140 & ~x142 & ~x163 & ~x167 & ~x172 & ~x199 & ~x218 & ~x257 & ~x282 & ~x295 & ~x308 & ~x338 & ~x389 & ~x473 & ~x503 & ~x558 & ~x565 & ~x566 & ~x587 & ~x590 & ~x596 & ~x611 & ~x614 & ~x622 & ~x623 & ~x625 & ~x634 & ~x636 & ~x637 & ~x638 & ~x648 & ~x653 & ~x665 & ~x668 & ~x718 & ~x750 & ~x754 & ~x757 & ~x764 & ~x779;
assign c1163 =  x272 & ~x3 & ~x54 & ~x88 & ~x99 & ~x103 & ~x128 & ~x129 & ~x131 & ~x132 & ~x141 & ~x142 & ~x143 & ~x475 & ~x487 & ~x616 & ~x645 & ~x668 & ~x726 & ~x770;
assign c1165 =  x290 & ~x35 & ~x39 & ~x40 & ~x48 & ~x50 & ~x53 & ~x59 & ~x61 & ~x62 & ~x73 & ~x86 & ~x91 & ~x94 & ~x95 & ~x97 & ~x105 & ~x110 & ~x119 & ~x120 & ~x123 & ~x124 & ~x127 & ~x128 & ~x142 & ~x158 & ~x167 & ~x169 & ~x198 & ~x201 & ~x223 & ~x251 & ~x252 & ~x279 & ~x308 & ~x333 & ~x334 & ~x349 & ~x350 & ~x361 & ~x390 & ~x449 & ~x451 & ~x592 & ~x615 & ~x619 & ~x621 & ~x622 & ~x623 & ~x646 & ~x704 & ~x705 & ~x706 & ~x724 & ~x728 & ~x747 & ~x748 & ~x753 & ~x754 & ~x756 & ~x761 & ~x775;
assign c1167 =  x205 & ~x52 & ~x117 & ~x606 & ~x766;
assign c1169 =  x346 & ~x5 & ~x8 & ~x11 & ~x14 & ~x19 & ~x23 & ~x32 & ~x33 & ~x44 & ~x59 & ~x65 & ~x68 & ~x76 & ~x102 & ~x112 & ~x118 & ~x120 & ~x123 & ~x138 & ~x143 & ~x148 & ~x172 & ~x173 & ~x175 & ~x176 & ~x177 & ~x230 & ~x254 & ~x282 & ~x284 & ~x308 & ~x365 & ~x392 & ~x525 & ~x528 & ~x554 & ~x556 & ~x560 & ~x562 & ~x565 & ~x582 & ~x606 & ~x607 & ~x609 & ~x613 & ~x615 & ~x618 & ~x620 & ~x634 & ~x636 & ~x640 & ~x643 & ~x664 & ~x670 & ~x675 & ~x703 & ~x709 & ~x736 & ~x743 & ~x744 & ~x765 & ~x766 & ~x782;
assign c1171 =  x235 &  x270 & ~x4 & ~x8 & ~x9 & ~x11 & ~x14 & ~x22 & ~x31 & ~x37 & ~x41 & ~x42 & ~x44 & ~x49 & ~x66 & ~x87 & ~x91 & ~x92 & ~x100 & ~x115 & ~x116 & ~x122 & ~x123 & ~x131 & ~x147 & ~x149 & ~x167 & ~x195 & ~x222 & ~x250 & ~x389 & ~x390 & ~x418 & ~x480 & ~x509 & ~x534 & ~x538 & ~x557 & ~x559 & ~x585 & ~x607 & ~x675 & ~x676 & ~x696 & ~x736 & ~x755 & ~x777;
assign c1173 =  x566 &  x625 & ~x16 & ~x34 & ~x67 & ~x75 & ~x87 & ~x89 & ~x118 & ~x167 & ~x171 & ~x196 & ~x306 & ~x307 & ~x365 & ~x390 & ~x417 & ~x419 & ~x561 & ~x587 & ~x588 & ~x616 & ~x647 & ~x677 & ~x700 & ~x711 & ~x721 & ~x734 & ~x753 & ~x756 & ~x758 & ~x760 & ~x762 & ~x768 & ~x770 & ~x775;
assign c1175 = ~x5 & ~x8 & ~x10 & ~x12 & ~x15 & ~x30 & ~x43 & ~x53 & ~x58 & ~x61 & ~x67 & ~x68 & ~x77 & ~x79 & ~x90 & ~x94 & ~x112 & ~x122 & ~x123 & ~x125 & ~x194 & ~x195 & ~x197 & ~x224 & ~x226 & ~x253 & ~x280 & ~x296 & ~x307 & ~x310 & ~x317 & ~x332 & ~x345 & ~x417 & ~x427 & ~x440 & ~x444 & ~x448 & ~x449 & ~x450 & ~x475 & ~x496 & ~x497 & ~x530 & ~x557 & ~x559 & ~x587 & ~x589 & ~x608 & ~x620 & ~x641 & ~x647 & ~x669 & ~x674 & ~x691 & ~x696 & ~x701 & ~x716 & ~x731 & ~x732 & ~x737 & ~x763 & ~x769 & ~x773 & ~x775;
assign c1177 =  x205 & ~x5 & ~x11 & ~x29 & ~x72 & ~x79 & ~x100 & ~x107 & ~x116 & ~x132 & ~x170 & ~x291 & ~x364 & ~x453 & ~x480 & ~x617 & ~x678 & ~x681 & ~x704 & ~x724 & ~x730 & ~x743 & ~x758 & ~x762 & ~x766 & ~x772;
assign c1179 =  x437 & ~x6 & ~x8 & ~x10 & ~x13 & ~x17 & ~x18 & ~x23 & ~x25 & ~x28 & ~x36 & ~x37 & ~x42 & ~x43 & ~x44 & ~x46 & ~x53 & ~x54 & ~x56 & ~x62 & ~x64 & ~x67 & ~x68 & ~x69 & ~x70 & ~x79 & ~x81 & ~x98 & ~x108 & ~x114 & ~x117 & ~x118 & ~x120 & ~x139 & ~x145 & ~x167 & ~x169 & ~x171 & ~x197 & ~x222 & ~x223 & ~x250 & ~x253 & ~x254 & ~x277 & ~x332 & ~x334 & ~x335 & ~x336 & ~x364 & ~x365 & ~x393 & ~x416 & ~x419 & ~x421 & ~x425 & ~x449 & ~x501 & ~x503 & ~x505 & ~x528 & ~x531 & ~x555 & ~x556 & ~x557 & ~x584 & ~x612 & ~x614 & ~x641 & ~x644 & ~x668 & ~x673 & ~x676 & ~x697 & ~x701 & ~x722 & ~x725 & ~x727 & ~x733 & ~x738 & ~x739 & ~x746 & ~x763 & ~x767 & ~x776;
assign c1181 =  x204 & ~x6 & ~x9 & ~x18 & ~x30 & ~x116 & ~x117 & ~x132 & ~x138 & ~x161 & ~x171 & ~x279 & ~x291 & ~x362 & ~x366 & ~x385 & ~x388 & ~x426 & ~x448 & ~x720 & ~x740 & ~x747 & ~x755 & ~x776;
assign c1183 =  x494 & ~x11 & ~x23 & ~x26 & ~x30 & ~x31 & ~x34 & ~x40 & ~x44 & ~x52 & ~x77 & ~x80 & ~x92 & ~x115 & ~x120 & ~x122 & ~x139 & ~x145 & ~x149 & ~x150 & ~x152 & ~x171 & ~x193 & ~x198 & ~x199 & ~x220 & ~x227 & ~x279 & ~x305 & ~x310 & ~x331 & ~x366 & ~x387 & ~x392 & ~x393 & ~x450 & ~x476 & ~x615 & ~x616 & ~x642 & ~x665 & ~x667 & ~x725 & ~x731 & ~x755 & ~x757 & ~x765;
assign c1185 =  x485 &  x492 &  x513 & ~x2 & ~x7 & ~x28 & ~x30 & ~x74 & ~x76 & ~x81 & ~x139 & ~x142 & ~x199 & ~x200 & ~x201 & ~x229 & ~x257 & ~x280 & ~x306 & ~x336 & ~x339 & ~x340 & ~x363 & ~x368 & ~x388 & ~x448 & ~x449 & ~x498 & ~x504 & ~x532 & ~x533 & ~x558 & ~x584 & ~x585 & ~x587 & ~x588 & ~x590 & ~x591 & ~x619 & ~x640 & ~x645 & ~x646 & ~x648 & ~x660 & ~x672 & ~x688 & ~x692 & ~x726 & ~x737 & ~x743 & ~x751 & ~x752 & ~x766 & ~x771 & ~x776 & ~x780;
assign c1187 =  x382 &  x383 & ~x10 & ~x24 & ~x26 & ~x31 & ~x47 & ~x57 & ~x88 & ~x109 & ~x114 & ~x115 & ~x136 & ~x137 & ~x142 & ~x144 & ~x193 & ~x225 & ~x252 & ~x277 & ~x278 & ~x307 & ~x340 & ~x366 & ~x393 & ~x476 & ~x478 & ~x502 & ~x534 & ~x587 & ~x642 & ~x690 & ~x691 & ~x693 & ~x694 & ~x697 & ~x701 & ~x741 & ~x754 & ~x755 & ~x764;
assign c1189 =  x209 &  x298 & ~x4 & ~x21 & ~x30 & ~x42 & ~x44 & ~x55 & ~x73 & ~x104 & ~x109 & ~x113 & ~x140 & ~x225 & ~x254 & ~x281 & ~x365 & ~x393 & ~x445 & ~x453 & ~x454 & ~x477 & ~x479 & ~x534 & ~x675 & ~x701 & ~x717 & ~x762 & ~x765 & ~x771;
assign c1191 =  x432 & ~x45 & ~x54 & ~x108 & ~x140 & ~x223 & ~x256 & ~x378 & ~x526 & ~x561 & ~x637 & ~x662 & ~x772;
assign c1193 =  x289 & ~x7 & ~x10 & ~x35 & ~x59 & ~x63 & ~x68 & ~x79 & ~x84 & ~x98 & ~x110 & ~x114 & ~x145 & ~x169 & ~x170 & ~x223 & ~x225 & ~x280 & ~x335 & ~x361 & ~x366 & ~x446 & ~x450 & ~x503 & ~x509 & ~x532 & ~x561 & ~x578 & ~x593 & ~x607 & ~x616 & ~x619 & ~x624 & ~x640 & ~x643 & ~x672 & ~x694 & ~x729 & ~x731 & ~x749 & ~x752 & ~x756 & ~x772 & ~x780 & ~x782 & ~x783;
assign c1195 =  x456 & ~x3 & ~x6 & ~x9 & ~x13 & ~x15 & ~x23 & ~x25 & ~x32 & ~x42 & ~x50 & ~x51 & ~x58 & ~x59 & ~x61 & ~x87 & ~x117 & ~x118 & ~x137 & ~x169 & ~x170 & ~x195 & ~x198 & ~x252 & ~x253 & ~x254 & ~x255 & ~x256 & ~x278 & ~x279 & ~x283 & ~x362 & ~x393 & ~x423 & ~x449 & ~x452 & ~x503 & ~x585 & ~x586 & ~x592 & ~x614 & ~x644 & ~x645 & ~x649 & ~x668 & ~x672 & ~x674 & ~x675 & ~x676 & ~x677 & ~x680 & ~x691 & ~x698 & ~x702 & ~x722 & ~x725 & ~x727 & ~x730 & ~x735 & ~x740 & ~x754 & ~x755 & ~x758 & ~x769 & ~x771 & ~x782;
assign c1197 =  x629 & ~x86 & ~x109 & ~x113 & ~x192 & ~x340 & ~x390 & ~x499 & ~x517 & ~x537 & ~x593 & ~x701 & ~x711 & ~x726 & ~x762 & ~x777;
assign c1199 =  x181 &  x243 & ~x2 & ~x3 & ~x6 & ~x8 & ~x17 & ~x19 & ~x31 & ~x32 & ~x36 & ~x38 & ~x40 & ~x42 & ~x45 & ~x56 & ~x59 & ~x62 & ~x69 & ~x70 & ~x73 & ~x77 & ~x82 & ~x85 & ~x89 & ~x94 & ~x95 & ~x105 & ~x109 & ~x112 & ~x116 & ~x117 & ~x118 & ~x122 & ~x123 & ~x136 & ~x192 & ~x199 & ~x200 & ~x221 & ~x224 & ~x228 & ~x252 & ~x253 & ~x255 & ~x277 & ~x282 & ~x283 & ~x305 & ~x333 & ~x334 & ~x336 & ~x337 & ~x338 & ~x360 & ~x361 & ~x366 & ~x391 & ~x393 & ~x416 & ~x417 & ~x421 & ~x423 & ~x445 & ~x448 & ~x449 & ~x473 & ~x477 & ~x501 & ~x529 & ~x532 & ~x584 & ~x585 & ~x615 & ~x641 & ~x642 & ~x646 & ~x670 & ~x672 & ~x674 & ~x696 & ~x700 & ~x731 & ~x733 & ~x738 & ~x743 & ~x744 & ~x745 & ~x746 & ~x747 & ~x751 & ~x753 & ~x763 & ~x764 & ~x767 & ~x779 & ~x782;
assign c1201 =  x430 & ~x3 & ~x16 & ~x283 & ~x337 & ~x351 & ~x587 & ~x643 & ~x646 & ~x695 & ~x703 & ~x717 & ~x753 & ~x767 & ~x774;
assign c1203 =  x151 & ~x11 & ~x14 & ~x16 & ~x30 & ~x35 & ~x41 & ~x45 & ~x60 & ~x61 & ~x76 & ~x78 & ~x101 & ~x109 & ~x111 & ~x130 & ~x137 & ~x164 & ~x216 & ~x218 & ~x245 & ~x249 & ~x250 & ~x262 & ~x282 & ~x292 & ~x309 & ~x332 & ~x395 & ~x396 & ~x419 & ~x449 & ~x477 & ~x479 & ~x509 & ~x534 & ~x640 & ~x642 & ~x645 & ~x698 & ~x712 & ~x716 & ~x731 & ~x736 & ~x756 & ~x759 & ~x766;
assign c1205 =  x493 & ~x16 & ~x19 & ~x28 & ~x29 & ~x33 & ~x34 & ~x35 & ~x42 & ~x48 & ~x59 & ~x60 & ~x78 & ~x80 & ~x86 & ~x110 & ~x112 & ~x141 & ~x142 & ~x143 & ~x147 & ~x150 & ~x151 & ~x163 & ~x164 & ~x177 & ~x204 & ~x222 & ~x224 & ~x229 & ~x252 & ~x280 & ~x281 & ~x283 & ~x286 & ~x305 & ~x307 & ~x317 & ~x339 & ~x370 & ~x390 & ~x415 & ~x442 & ~x443 & ~x447 & ~x452 & ~x478 & ~x498 & ~x499 & ~x502 & ~x523 & ~x527 & ~x561 & ~x587 & ~x607 & ~x617 & ~x634 & ~x636 & ~x639 & ~x690 & ~x697 & ~x703 & ~x706 & ~x720 & ~x727 & ~x728 & ~x737 & ~x738 & ~x740 & ~x741 & ~x759 & ~x761 & ~x762 & ~x767 & ~x778 & ~x780 & ~x781 & ~x782;
assign c1207 =  x236 &  x353 & ~x11 & ~x28 & ~x53 & ~x76 & ~x125 & ~x166 & ~x196 & ~x197 & ~x250 & ~x308 & ~x361 & ~x531 & ~x539 & ~x596 & ~x644 & ~x699 & ~x701 & ~x704 & ~x738 & ~x781;
assign c1209 =  x181 &  x269 & ~x1 & ~x22 & ~x23 & ~x25 & ~x28 & ~x30 & ~x67 & ~x70 & ~x74 & ~x76 & ~x88 & ~x100 & ~x115 & ~x133 & ~x138 & ~x249 & ~x250 & ~x265 & ~x281 & ~x308 & ~x331 & ~x341 & ~x366 & ~x416 & ~x419 & ~x455 & ~x479 & ~x480 & ~x501 & ~x585 & ~x588 & ~x589 & ~x644 & ~x673 & ~x695 & ~x701 & ~x702 & ~x703 & ~x746 & ~x747 & ~x756 & ~x770 & ~x776 & ~x781;
assign c1211 =  x631 & ~x9 & ~x45 & ~x46 & ~x54 & ~x55 & ~x66 & ~x67 & ~x71 & ~x81 & ~x88 & ~x97 & ~x112 & ~x116 & ~x196 & ~x199 & ~x227 & ~x229 & ~x246 & ~x250 & ~x259 & ~x284 & ~x307 & ~x309 & ~x312 & ~x317 & ~x332 & ~x387 & ~x392 & ~x393 & ~x394 & ~x398 & ~x413 & ~x415 & ~x419 & ~x420 & ~x427 & ~x446 & ~x448 & ~x472 & ~x506 & ~x546 & ~x557 & ~x560 & ~x585 & ~x590 & ~x593 & ~x615 & ~x617 & ~x649 & ~x681 & ~x709 & ~x710 & ~x728 & ~x748 & ~x750 & ~x758;
assign c1213 =  x185 &  x405 &  x434 & ~x13 & ~x15 & ~x23 & ~x24 & ~x25 & ~x52 & ~x79 & ~x113 & ~x167 & ~x201 & ~x204 & ~x280 & ~x323 & ~x392 & ~x395 & ~x613 & ~x690 & ~x698 & ~x720 & ~x783;
assign c1215 =  x437 &  x438 & ~x0 & ~x34 & ~x35 & ~x37 & ~x39 & ~x41 & ~x42 & ~x43 & ~x45 & ~x48 & ~x49 & ~x54 & ~x57 & ~x64 & ~x65 & ~x67 & ~x78 & ~x80 & ~x91 & ~x111 & ~x112 & ~x114 & ~x116 & ~x118 & ~x142 & ~x168 & ~x196 & ~x198 & ~x223 & ~x249 & ~x251 & ~x333 & ~x334 & ~x338 & ~x393 & ~x395 & ~x531 & ~x554 & ~x556 & ~x558 & ~x561 & ~x583 & ~x643 & ~x669 & ~x671 & ~x673 & ~x686 & ~x704 & ~x707 & ~x709 & ~x714 & ~x724 & ~x726 & ~x732 & ~x735 & ~x749 & ~x765 & ~x774;
assign c1217 =  x269 &  x491 & ~x10 & ~x24 & ~x25 & ~x60 & ~x62 & ~x65 & ~x88 & ~x90 & ~x105 & ~x112 & ~x116 & ~x129 & ~x130 & ~x146 & ~x156 & ~x158 & ~x159 & ~x186 & ~x197 & ~x251 & ~x283 & ~x306 & ~x313 & ~x354 & ~x361 & ~x362 & ~x393 & ~x417 & ~x421 & ~x448 & ~x449 & ~x473 & ~x503 & ~x530 & ~x534 & ~x535 & ~x557 & ~x562 & ~x588 & ~x621 & ~x623 & ~x642 & ~x671 & ~x678 & ~x693 & ~x702 & ~x738 & ~x747 & ~x749 & ~x763 & ~x774 & ~x775 & ~x780;
assign c1219 =  x537 & ~x9 & ~x24 & ~x53 & ~x78 & ~x86 & ~x307 & ~x340 & ~x726 & ~x756;
assign c1221 =  x324 & ~x24 & ~x34 & ~x62 & ~x65 & ~x83 & ~x89 & ~x91 & ~x102 & ~x108 & ~x136 & ~x146 & ~x159 & ~x162 & ~x187 & ~x190 & ~x195 & ~x198 & ~x267 & ~x306 & ~x310 & ~x313 & ~x315 & ~x337 & ~x340 & ~x342 & ~x363 & ~x369 & ~x396 & ~x411 & ~x413 & ~x425 & ~x505 & ~x560 & ~x619 & ~x620 & ~x633 & ~x642 & ~x664 & ~x689 & ~x706 & ~x707 & ~x723 & ~x726 & ~x728 & ~x732 & ~x744 & ~x747 & ~x760 & ~x763 & ~x775;
assign c1223 =  x272 &  x273 & ~x52 & ~x106 & ~x161 & ~x163 & ~x179 & ~x195 & ~x200 & ~x256 & ~x502 & ~x613 & ~x617;
assign c1225 =  x605 & ~x4 & ~x14 & ~x17 & ~x19 & ~x21 & ~x22 & ~x23 & ~x31 & ~x33 & ~x36 & ~x38 & ~x40 & ~x42 & ~x44 & ~x45 & ~x49 & ~x53 & ~x57 & ~x62 & ~x64 & ~x67 & ~x71 & ~x73 & ~x79 & ~x82 & ~x87 & ~x88 & ~x90 & ~x101 & ~x108 & ~x112 & ~x118 & ~x139 & ~x140 & ~x141 & ~x163 & ~x164 & ~x168 & ~x195 & ~x197 & ~x221 & ~x222 & ~x224 & ~x227 & ~x247 & ~x280 & ~x307 & ~x333 & ~x337 & ~x362 & ~x366 & ~x417 & ~x418 & ~x422 & ~x444 & ~x448 & ~x449 & ~x477 & ~x478 & ~x519 & ~x556 & ~x557 & ~x558 & ~x560 & ~x562 & ~x588 & ~x612 & ~x643 & ~x664 & ~x675 & ~x676 & ~x694 & ~x695 & ~x698 & ~x700 & ~x702 & ~x703 & ~x705 & ~x708 & ~x713 & ~x720 & ~x721 & ~x727 & ~x729 & ~x730 & ~x731 & ~x736 & ~x754 & ~x757 & ~x759 & ~x763 & ~x768 & ~x773 & ~x775 & ~x782;
assign c1227 =  x657 & ~x7 & ~x33 & ~x50 & ~x51 & ~x67 & ~x98 & ~x99 & ~x144 & ~x172 & ~x194 & ~x197 & ~x223 & ~x367 & ~x369 & ~x478 & ~x502 & ~x531 & ~x532 & ~x545 & ~x560 & ~x574 & ~x589 & ~x615 & ~x639 & ~x641 & ~x642 & ~x670 & ~x676 & ~x720 & ~x723 & ~x724 & ~x729 & ~x747 & ~x756 & ~x759 & ~x776 & ~x782;
assign c1229 =  x237 &  x244 & ~x10 & ~x12 & ~x19 & ~x44 & ~x103 & ~x142 & ~x150 & ~x283 & ~x391 & ~x397 & ~x693 & ~x753 & ~x762 & ~x777;
assign c1231 =  x235 & ~x26 & ~x35 & ~x39 & ~x43 & ~x54 & ~x62 & ~x106 & ~x107 & ~x110 & ~x114 & ~x116 & ~x128 & ~x137 & ~x139 & ~x148 & ~x151 & ~x154 & ~x155 & ~x191 & ~x218 & ~x283 & ~x339 & ~x420 & ~x473 & ~x505 & ~x536 & ~x559 & ~x561 & ~x582 & ~x619 & ~x634 & ~x646 & ~x699 & ~x720 & ~x728 & ~x749 & ~x756 & ~x759;
assign c1233 =  x410 &  x411 & ~x8 & ~x11 & ~x13 & ~x25 & ~x26 & ~x37 & ~x39 & ~x40 & ~x46 & ~x57 & ~x59 & ~x66 & ~x80 & ~x87 & ~x88 & ~x93 & ~x107 & ~x110 & ~x123 & ~x138 & ~x140 & ~x143 & ~x146 & ~x165 & ~x197 & ~x223 & ~x224 & ~x225 & ~x226 & ~x250 & ~x252 & ~x307 & ~x335 & ~x366 & ~x391 & ~x393 & ~x395 & ~x422 & ~x448 & ~x475 & ~x501 & ~x506 & ~x531 & ~x533 & ~x556 & ~x560 & ~x562 & ~x583 & ~x585 & ~x616 & ~x618 & ~x640 & ~x644 & ~x645 & ~x647 & ~x670 & ~x672 & ~x674 & ~x696 & ~x699 & ~x701 & ~x703 & ~x724 & ~x728 & ~x744 & ~x749 & ~x752 & ~x755 & ~x757 & ~x760 & ~x767 & ~x773 & ~x774 & ~x783;
assign c1235 =  x407 & ~x10 & ~x13 & ~x21 & ~x38 & ~x42 & ~x59 & ~x71 & ~x80 & ~x88 & ~x136 & ~x153 & ~x195 & ~x198 & ~x279 & ~x296 & ~x365 & ~x366 & ~x416 & ~x505 & ~x508 & ~x556 & ~x557 & ~x577 & ~x606 & ~x633 & ~x642 & ~x646 & ~x664 & ~x672 & ~x699 & ~x726 & ~x746 & ~x751 & ~x757 & ~x769;
assign c1237 =  x406 &  x407 &  x630 & ~x11 & ~x12 & ~x46 & ~x73 & ~x96 & ~x107 & ~x194 & ~x195 & ~x256 & ~x282 & ~x358 & ~x421 & ~x480 & ~x546 & ~x561 & ~x668 & ~x727 & ~x769 & ~x774 & ~x775 & ~x778 & ~x780 & ~x783;
assign c1239 =  x498 & ~x31 & ~x33 & ~x58 & ~x72 & ~x141 & ~x395 & ~x563 & ~x673 & ~x735 & ~x749 & ~x773;
assign c1241 =  x510 & ~x19 & ~x38 & ~x66 & ~x74 & ~x140 & ~x144 & ~x668 & ~x713 & ~x735 & ~x737 & ~x752 & ~x768;
assign c1243 =  x433 &  x577 & ~x20 & ~x32 & ~x35 & ~x172 & ~x196 & ~x219 & ~x228 & ~x282 & ~x423 & ~x507 & ~x557 & ~x618 & ~x681 & ~x683 & ~x726 & ~x732 & ~x739 & ~x743;
assign c1245 =  x684 & ~x1 & ~x2 & ~x19 & ~x23 & ~x28 & ~x30 & ~x31 & ~x34 & ~x37 & ~x38 & ~x39 & ~x40 & ~x41 & ~x44 & ~x45 & ~x50 & ~x55 & ~x58 & ~x61 & ~x70 & ~x85 & ~x86 & ~x88 & ~x90 & ~x92 & ~x102 & ~x103 & ~x104 & ~x109 & ~x110 & ~x115 & ~x118 & ~x122 & ~x123 & ~x125 & ~x132 & ~x135 & ~x139 & ~x145 & ~x176 & ~x196 & ~x197 & ~x200 & ~x201 & ~x223 & ~x227 & ~x229 & ~x251 & ~x256 & ~x280 & ~x282 & ~x309 & ~x361 & ~x365 & ~x366 & ~x367 & ~x368 & ~x391 & ~x422 & ~x426 & ~x445 & ~x447 & ~x450 & ~x470 & ~x471 & ~x473 & ~x476 & ~x479 & ~x480 & ~x481 & ~x510 & ~x526 & ~x535 & ~x553 & ~x564 & ~x587 & ~x588 & ~x590 & ~x592 & ~x614 & ~x634 & ~x637 & ~x644 & ~x645 & ~x648 & ~x661 & ~x669 & ~x670 & ~x671 & ~x674 & ~x687 & ~x693 & ~x694 & ~x698 & ~x699 & ~x700 & ~x702 & ~x714 & ~x718 & ~x720 & ~x730 & ~x736 & ~x743 & ~x746 & ~x747 & ~x748 & ~x749 & ~x750 & ~x752 & ~x755 & ~x757 & ~x759 & ~x760 & ~x761 & ~x763 & ~x770 & ~x779 & ~x780;
assign c1247 =  x438 & ~x9 & ~x23 & ~x42 & ~x54 & ~x139 & ~x145 & ~x166 & ~x223 & ~x224 & ~x333 & ~x369 & ~x388 & ~x418 & ~x448 & ~x533 & ~x545 & ~x584 & ~x613 & ~x665 & ~x673 & ~x721 & ~x732 & ~x763;
assign c1249 =  x460 &  x549 & ~x4 & ~x20 & ~x26 & ~x33 & ~x34 & ~x39 & ~x45 & ~x51 & ~x52 & ~x53 & ~x55 & ~x65 & ~x68 & ~x70 & ~x84 & ~x114 & ~x136 & ~x140 & ~x144 & ~x170 & ~x172 & ~x193 & ~x194 & ~x195 & ~x197 & ~x198 & ~x251 & ~x256 & ~x282 & ~x283 & ~x301 & ~x302 & ~x307 & ~x310 & ~x329 & ~x338 & ~x386 & ~x410 & ~x417 & ~x473 & ~x476 & ~x478 & ~x503 & ~x504 & ~x505 & ~x506 & ~x558 & ~x560 & ~x585 & ~x588 & ~x590 & ~x619 & ~x640 & ~x648 & ~x652 & ~x666 & ~x670 & ~x673 & ~x675 & ~x695 & ~x697 & ~x703 & ~x708 & ~x725 & ~x731 & ~x744 & ~x751 & ~x752 & ~x753 & ~x755 & ~x765 & ~x767 & ~x771 & ~x772 & ~x773 & ~x775;
assign c1251 =  x403 & ~x59 & ~x108 & ~x109 & ~x225 & ~x454 & ~x457 & ~x472 & ~x529 & ~x533 & ~x543 & ~x583 & ~x605 & ~x616 & ~x663 & ~x718 & ~x731 & ~x736 & ~x762 & ~x771;
assign c1253 =  x520 & ~x28 & ~x35 & ~x37 & ~x48 & ~x49 & ~x51 & ~x56 & ~x65 & ~x84 & ~x89 & ~x97 & ~x121 & ~x125 & ~x144 & ~x151 & ~x179 & ~x221 & ~x222 & ~x223 & ~x225 & ~x308 & ~x324 & ~x363 & ~x366 & ~x368 & ~x391 & ~x421 & ~x450 & ~x474 & ~x523 & ~x555 & ~x563 & ~x580 & ~x621 & ~x638 & ~x650 & ~x668 & ~x673 & ~x674 & ~x676 & ~x679 & ~x700 & ~x761 & ~x769 & ~x773 & ~x775;
assign c1255 =  x457 & ~x3 & ~x15 & ~x27 & ~x46 & ~x51 & ~x52 & ~x56 & ~x57 & ~x58 & ~x87 & ~x138 & ~x162 & ~x165 & ~x166 & ~x167 & ~x171 & ~x228 & ~x284 & ~x311 & ~x312 & ~x417 & ~x453 & ~x506 & ~x534 & ~x613 & ~x616 & ~x637 & ~x640 & ~x642 & ~x643 & ~x645 & ~x650 & ~x651 & ~x666 & ~x679 & ~x684 & ~x688 & ~x696 & ~x698 & ~x704 & ~x712 & ~x714 & ~x725 & ~x729 & ~x738 & ~x739 & ~x742 & ~x745 & ~x748 & ~x751 & ~x758;
assign c1257 =  x301 & ~x17 & ~x19 & ~x29 & ~x34 & ~x49 & ~x68 & ~x74 & ~x76 & ~x83 & ~x86 & ~x88 & ~x90 & ~x107 & ~x109 & ~x115 & ~x135 & ~x139 & ~x140 & ~x142 & ~x163 & ~x164 & ~x168 & ~x172 & ~x198 & ~x307 & ~x310 & ~x335 & ~x336 & ~x364 & ~x367 & ~x420 & ~x447 & ~x450 & ~x473 & ~x501 & ~x588 & ~x591 & ~x618 & ~x644 & ~x646 & ~x647 & ~x648 & ~x668 & ~x674 & ~x676 & ~x695 & ~x725 & ~x727 & ~x741 & ~x754 & ~x757 & ~x758 & ~x772 & ~x776 & ~x777;
assign c1259 =  x432 & ~x3 & ~x12 & ~x40 & ~x58 & ~x76 & ~x94 & ~x107 & ~x116 & ~x137 & ~x139 & ~x162 & ~x166 & ~x200 & ~x216 & ~x274 & ~x275 & ~x281 & ~x286 & ~x343 & ~x349 & ~x390 & ~x445 & ~x452 & ~x480 & ~x559 & ~x566 & ~x593 & ~x594 & ~x674 & ~x676 & ~x702 & ~x703 & ~x704 & ~x724 & ~x742 & ~x748 & ~x769 & ~x777 & ~x780 & ~x783;
assign c1261 = ~x1 & ~x13 & ~x14 & ~x15 & ~x17 & ~x24 & ~x30 & ~x31 & ~x32 & ~x35 & ~x37 & ~x39 & ~x42 & ~x46 & ~x47 & ~x52 & ~x55 & ~x63 & ~x64 & ~x87 & ~x90 & ~x107 & ~x110 & ~x114 & ~x115 & ~x118 & ~x132 & ~x141 & ~x160 & ~x167 & ~x171 & ~x172 & ~x174 & ~x227 & ~x280 & ~x307 & ~x350 & ~x351 & ~x361 & ~x362 & ~x364 & ~x389 & ~x395 & ~x396 & ~x421 & ~x423 & ~x449 & ~x477 & ~x503 & ~x504 & ~x507 & ~x532 & ~x534 & ~x560 & ~x564 & ~x594 & ~x613 & ~x616 & ~x633 & ~x635 & ~x643 & ~x663 & ~x674 & ~x675 & ~x692 & ~x719 & ~x721 & ~x723 & ~x725 & ~x731 & ~x751 & ~x755 & ~x766 & ~x771 & ~x775;
assign c1263 =  x469 & ~x0 & ~x10 & ~x28 & ~x42 & ~x54 & ~x60 & ~x79 & ~x80 & ~x108 & ~x115 & ~x194 & ~x282 & ~x335 & ~x338 & ~x476 & ~x479 & ~x504 & ~x614 & ~x615 & ~x617 & ~x645 & ~x673 & ~x712 & ~x726 & ~x728 & ~x761 & ~x762 & ~x766 & ~x773 & ~x778;
assign c1265 = ~x2 & ~x42 & ~x46 & ~x48 & ~x53 & ~x63 & ~x69 & ~x71 & ~x72 & ~x76 & ~x78 & ~x80 & ~x82 & ~x110 & ~x112 & ~x142 & ~x154 & ~x170 & ~x171 & ~x195 & ~x201 & ~x229 & ~x250 & ~x362 & ~x363 & ~x364 & ~x366 & ~x379 & ~x394 & ~x420 & ~x451 & ~x503 & ~x506 & ~x557 & ~x559 & ~x607 & ~x614 & ~x619 & ~x640 & ~x641 & ~x642 & ~x644 & ~x658 & ~x664 & ~x675 & ~x676 & ~x685 & ~x700 & ~x712 & ~x719 & ~x722 & ~x728 & ~x731 & ~x734 & ~x750 & ~x754 & ~x758 & ~x759 & ~x763 & ~x764 & ~x766 & ~x772 & ~x773 & ~x775 & ~x776 & ~x777 & ~x780 & ~x782 & ~x783;
assign c1267 =  x513 &  x540 &  x541 &  x601 & ~x47 & ~x62 & ~x71 & ~x73 & ~x86 & ~x136 & ~x142 & ~x168 & ~x172 & ~x286 & ~x306 & ~x314 & ~x329 & ~x341 & ~x382 & ~x503 & ~x504 & ~x589 & ~x614 & ~x710 & ~x733 & ~x750 & ~x774 & ~x781;
assign c1269 =  x468 & ~x0 & ~x1 & ~x5 & ~x7 & ~x12 & ~x13 & ~x14 & ~x16 & ~x19 & ~x20 & ~x21 & ~x23 & ~x29 & ~x32 & ~x37 & ~x38 & ~x40 & ~x42 & ~x44 & ~x46 & ~x48 & ~x51 & ~x55 & ~x56 & ~x65 & ~x73 & ~x74 & ~x78 & ~x82 & ~x84 & ~x87 & ~x106 & ~x111 & ~x112 & ~x114 & ~x115 & ~x137 & ~x138 & ~x140 & ~x143 & ~x163 & ~x165 & ~x168 & ~x169 & ~x171 & ~x192 & ~x221 & ~x222 & ~x249 & ~x277 & ~x305 & ~x308 & ~x333 & ~x335 & ~x360 & ~x361 & ~x363 & ~x364 & ~x366 & ~x393 & ~x447 & ~x476 & ~x503 & ~x504 & ~x556 & ~x558 & ~x560 & ~x585 & ~x586 & ~x587 & ~x588 & ~x617 & ~x618 & ~x619 & ~x641 & ~x644 & ~x645 & ~x673 & ~x676 & ~x696 & ~x701 & ~x702 & ~x703 & ~x720 & ~x725 & ~x726 & ~x728 & ~x733 & ~x734 & ~x736 & ~x737 & ~x741 & ~x748 & ~x749 & ~x750 & ~x753 & ~x754 & ~x755 & ~x758 & ~x767 & ~x777 & ~x778 & ~x779 & ~x780 & ~x782;
assign c1271 =  x604 & ~x6 & ~x7 & ~x11 & ~x14 & ~x20 & ~x25 & ~x26 & ~x29 & ~x30 & ~x34 & ~x46 & ~x53 & ~x55 & ~x57 & ~x60 & ~x69 & ~x73 & ~x101 & ~x108 & ~x113 & ~x130 & ~x167 & ~x170 & ~x197 & ~x252 & ~x308 & ~x309 & ~x334 & ~x339 & ~x364 & ~x391 & ~x392 & ~x396 & ~x418 & ~x419 & ~x420 & ~x423 & ~x447 & ~x463 & ~x476 & ~x477 & ~x479 & ~x504 & ~x532 & ~x559 & ~x560 & ~x615 & ~x617 & ~x618 & ~x642 & ~x646 & ~x666 & ~x675 & ~x689 & ~x692 & ~x694 & ~x695 & ~x696 & ~x698 & ~x702 & ~x709 & ~x722 & ~x726 & ~x729 & ~x731 & ~x735 & ~x757 & ~x765 & ~x770 & ~x778 & ~x783;
assign c1273 =  x216 & ~x13 & ~x23 & ~x25 & ~x27 & ~x28 & ~x33 & ~x36 & ~x41 & ~x42 & ~x43 & ~x45 & ~x57 & ~x58 & ~x61 & ~x64 & ~x70 & ~x72 & ~x73 & ~x78 & ~x89 & ~x106 & ~x112 & ~x120 & ~x134 & ~x228 & ~x250 & ~x258 & ~x279 & ~x284 & ~x306 & ~x340 & ~x381 & ~x394 & ~x419 & ~x424 & ~x449 & ~x452 & ~x475 & ~x500 & ~x560 & ~x562 & ~x586 & ~x587 & ~x612 & ~x614 & ~x642 & ~x645 & ~x669 & ~x672 & ~x697 & ~x701 & ~x716 & ~x733 & ~x745 & ~x748 & ~x752 & ~x755 & ~x756 & ~x758 & ~x760 & ~x766 & ~x773 & ~x782 & ~x783;
assign c1275 =  x210 & ~x25 & ~x53 & ~x64 & ~x77 & ~x97 & ~x109 & ~x129 & ~x154 & ~x155 & ~x157 & ~x158 & ~x164 & ~x171 & ~x191 & ~x220 & ~x293 & ~x312 & ~x357 & ~x364 & ~x371 & ~x441 & ~x540 & ~x589 & ~x595 & ~x650 & ~x733 & ~x754 & ~x774 & ~x776;
assign c1277 =  x232 & ~x7 & ~x8 & ~x13 & ~x26 & ~x36 & ~x48 & ~x49 & ~x56 & ~x62 & ~x87 & ~x97 & ~x99 & ~x104 & ~x106 & ~x108 & ~x109 & ~x111 & ~x116 & ~x119 & ~x128 & ~x166 & ~x169 & ~x173 & ~x199 & ~x275 & ~x283 & ~x304 & ~x337 & ~x339 & ~x395 & ~x422 & ~x475 & ~x476 & ~x534 & ~x562 & ~x589 & ~x614 & ~x756 & ~x758 & ~x760 & ~x780 & ~x782;
assign c1279 =  x440 & ~x0 & ~x1 & ~x7 & ~x8 & ~x15 & ~x16 & ~x24 & ~x25 & ~x29 & ~x32 & ~x37 & ~x40 & ~x43 & ~x46 & ~x49 & ~x50 & ~x51 & ~x53 & ~x60 & ~x89 & ~x91 & ~x103 & ~x111 & ~x113 & ~x137 & ~x141 & ~x164 & ~x165 & ~x167 & ~x191 & ~x194 & ~x222 & ~x223 & ~x251 & ~x252 & ~x253 & ~x277 & ~x278 & ~x279 & ~x308 & ~x366 & ~x393 & ~x419 & ~x420 & ~x503 & ~x507 & ~x531 & ~x534 & ~x558 & ~x561 & ~x586 & ~x587 & ~x642 & ~x646 & ~x703 & ~x708 & ~x724 & ~x736 & ~x759 & ~x763 & ~x764 & ~x769 & ~x781 & ~x782 & ~x783;
assign c1281 =  x271 &  x272 & ~x9 & ~x10 & ~x44 & ~x45 & ~x59 & ~x74 & ~x81 & ~x160 & ~x171 & ~x190 & ~x226 & ~x307 & ~x368 & ~x392 & ~x395 & ~x396 & ~x419 & ~x421 & ~x448 & ~x503 & ~x584 & ~x667 & ~x699 & ~x733 & ~x740 & ~x757 & ~x760;
assign c1283 =  x259 & ~x0 & ~x17 & ~x18 & ~x24 & ~x31 & ~x36 & ~x37 & ~x43 & ~x44 & ~x47 & ~x64 & ~x72 & ~x74 & ~x77 & ~x79 & ~x84 & ~x88 & ~x106 & ~x109 & ~x128 & ~x131 & ~x132 & ~x138 & ~x159 & ~x160 & ~x161 & ~x164 & ~x188 & ~x223 & ~x251 & ~x366 & ~x391 & ~x421 & ~x447 & ~x476 & ~x479 & ~x505 & ~x507 & ~x508 & ~x532 & ~x562 & ~x586 & ~x587 & ~x589 & ~x615 & ~x621 & ~x642 & ~x644 & ~x645 & ~x669 & ~x673 & ~x677 & ~x679 & ~x700 & ~x725 & ~x726 & ~x727 & ~x729 & ~x740 & ~x756 & ~x759 & ~x763 & ~x773 & ~x782 & ~x783;
assign c1285 =  x151 & ~x15 & ~x18 & ~x20 & ~x28 & ~x30 & ~x31 & ~x48 & ~x57 & ~x66 & ~x72 & ~x74 & ~x75 & ~x83 & ~x89 & ~x133 & ~x264 & ~x275 & ~x276 & ~x278 & ~x304 & ~x309 & ~x330 & ~x339 & ~x365 & ~x368 & ~x390 & ~x393 & ~x425 & ~x446 & ~x453 & ~x529 & ~x587 & ~x591 & ~x617 & ~x642 & ~x672 & ~x697 & ~x715 & ~x720 & ~x732 & ~x741 & ~x743 & ~x773 & ~x775;
assign c1287 =  x180 &  x433 & ~x11 & ~x17 & ~x40 & ~x57 & ~x62 & ~x64 & ~x67 & ~x68 & ~x71 & ~x75 & ~x85 & ~x88 & ~x107 & ~x117 & ~x145 & ~x229 & ~x250 & ~x252 & ~x278 & ~x280 & ~x305 & ~x306 & ~x308 & ~x321 & ~x331 & ~x337 & ~x363 & ~x392 & ~x476 & ~x477 & ~x532 & ~x533 & ~x588 & ~x672 & ~x689 & ~x691 & ~x700 & ~x709 & ~x720 & ~x730 & ~x741 & ~x769 & ~x774;
assign c1289 =  x515 & ~x2 & ~x20 & ~x48 & ~x54 & ~x78 & ~x88 & ~x90 & ~x103 & ~x113 & ~x158 & ~x164 & ~x188 & ~x191 & ~x200 & ~x215 & ~x217 & ~x225 & ~x251 & ~x253 & ~x284 & ~x303 & ~x308 & ~x335 & ~x358 & ~x361 & ~x368 & ~x395 & ~x418 & ~x419 & ~x451 & ~x504 & ~x536 & ~x537 & ~x560 & ~x563 & ~x566 & ~x617 & ~x653 & ~x669 & ~x671 & ~x684 & ~x698 & ~x709 & ~x711 & ~x718 & ~x724 & ~x743 & ~x744 & ~x752 & ~x758 & ~x760 & ~x765 & ~x769 & ~x775;
assign c1291 =  x461 &  x489 &  x490 & ~x115 & ~x227 & ~x315 & ~x378 & ~x394 & ~x640 & ~x675 & ~x679 & ~x759 & ~x769;
assign c1293 =  x374 & ~x4 & ~x7 & ~x16 & ~x25 & ~x29 & ~x36 & ~x37 & ~x39 & ~x42 & ~x43 & ~x45 & ~x61 & ~x70 & ~x88 & ~x95 & ~x102 & ~x106 & ~x144 & ~x166 & ~x171 & ~x194 & ~x225 & ~x227 & ~x255 & ~x285 & ~x306 & ~x308 & ~x336 & ~x422 & ~x424 & ~x451 & ~x475 & ~x476 & ~x479 & ~x501 & ~x504 & ~x520 & ~x529 & ~x592 & ~x614 & ~x616 & ~x639 & ~x643 & ~x646 & ~x648 & ~x671 & ~x695 & ~x696 & ~x697 & ~x698 & ~x699 & ~x716 & ~x718 & ~x730 & ~x731 & ~x741 & ~x751 & ~x756 & ~x772 & ~x775 & ~x779 & ~x780;
assign c1295 =  x263 &  x264 & ~x3 & ~x7 & ~x8 & ~x12 & ~x17 & ~x24 & ~x32 & ~x36 & ~x43 & ~x44 & ~x45 & ~x47 & ~x51 & ~x65 & ~x73 & ~x77 & ~x78 & ~x79 & ~x88 & ~x97 & ~x99 & ~x125 & ~x126 & ~x130 & ~x151 & ~x155 & ~x169 & ~x172 & ~x173 & ~x174 & ~x193 & ~x199 & ~x220 & ~x225 & ~x253 & ~x254 & ~x301 & ~x308 & ~x336 & ~x368 & ~x369 & ~x384 & ~x391 & ~x393 & ~x425 & ~x450 & ~x453 & ~x455 & ~x456 & ~x472 & ~x473 & ~x499 & ~x527 & ~x557 & ~x578 & ~x618 & ~x620 & ~x623 & ~x645 & ~x662 & ~x666 & ~x678 & ~x699 & ~x729 & ~x761 & ~x764 & ~x766 & ~x778;
assign c1297 =  x236 &  x240 & ~x16 & ~x30 & ~x36 & ~x43 & ~x72 & ~x87 & ~x93 & ~x110 & ~x115 & ~x119 & ~x124 & ~x128 & ~x132 & ~x133 & ~x222 & ~x253 & ~x256 & ~x311 & ~x362 & ~x363 & ~x393 & ~x505 & ~x606 & ~x614 & ~x619 & ~x697 & ~x713 & ~x757 & ~x780;
assign c1299 =  x382 & ~x1 & ~x5 & ~x10 & ~x12 & ~x14 & ~x19 & ~x27 & ~x28 & ~x32 & ~x33 & ~x37 & ~x55 & ~x59 & ~x61 & ~x63 & ~x80 & ~x84 & ~x86 & ~x88 & ~x109 & ~x110 & ~x132 & ~x133 & ~x135 & ~x140 & ~x160 & ~x162 & ~x164 & ~x165 & ~x169 & ~x189 & ~x192 & ~x196 & ~x220 & ~x222 & ~x247 & ~x276 & ~x304 & ~x333 & ~x335 & ~x337 & ~x368 & ~x392 & ~x417 & ~x422 & ~x426 & ~x432 & ~x444 & ~x445 & ~x531 & ~x559 & ~x585 & ~x586 & ~x619 & ~x643 & ~x645 & ~x699 & ~x702 & ~x704 & ~x724 & ~x729 & ~x731 & ~x733 & ~x748 & ~x752 & ~x755 & ~x756 & ~x758 & ~x761 & ~x765 & ~x769 & ~x778 & ~x780;
assign c20 =  x516 & ~x14 & ~x23 & ~x27 & ~x28 & ~x39 & ~x42 & ~x48 & ~x59 & ~x78 & ~x82 & ~x99 & ~x142 & ~x188 & ~x191 & ~x245 & ~x273 & ~x280 & ~x300 & ~x302 & ~x310 & ~x336 & ~x391 & ~x394 & ~x396 & ~x397 & ~x399 & ~x425 & ~x450 & ~x533 & ~x564 & ~x643 & ~x673 & ~x688 & ~x689 & ~x690 & ~x702 & ~x704 & ~x708 & ~x710 & ~x712 & ~x713 & ~x719 & ~x757 & ~x761 & ~x766 & ~x770;
assign c22 =  x474;
assign c24 =  x582 & ~x497;
assign c26 =  x477;
assign c28 =  x569 & ~x2 & ~x4 & ~x7 & ~x9 & ~x10 & ~x11 & ~x12 & ~x13 & ~x15 & ~x16 & ~x18 & ~x19 & ~x21 & ~x25 & ~x31 & ~x42 & ~x43 & ~x50 & ~x51 & ~x59 & ~x61 & ~x68 & ~x69 & ~x71 & ~x73 & ~x79 & ~x83 & ~x84 & ~x85 & ~x95 & ~x96 & ~x98 & ~x99 & ~x101 & ~x105 & ~x107 & ~x108 & ~x111 & ~x112 & ~x117 & ~x122 & ~x123 & ~x135 & ~x137 & ~x139 & ~x140 & ~x141 & ~x143 & ~x146 & ~x149 & ~x167 & ~x174 & ~x193 & ~x201 & ~x219 & ~x221 & ~x222 & ~x230 & ~x248 & ~x252 & ~x256 & ~x257 & ~x277 & ~x281 & ~x283 & ~x309 & ~x334 & ~x335 & ~x337 & ~x338 & ~x339 & ~x340 & ~x341 & ~x361 & ~x362 & ~x366 & ~x368 & ~x370 & ~x371 & ~x372 & ~x376 & ~x377 & ~x393 & ~x394 & ~x414 & ~x416 & ~x417 & ~x420 & ~x448 & ~x475 & ~x496 & ~x504 & ~x505 & ~x528 & ~x529 & ~x531 & ~x554 & ~x560 & ~x585 & ~x587 & ~x589 & ~x614 & ~x615 & ~x640 & ~x641 & ~x668 & ~x669 & ~x671 & ~x672 & ~x690 & ~x692 & ~x693 & ~x695 & ~x699 & ~x700 & ~x702 & ~x704 & ~x705 & ~x706 & ~x709 & ~x710 & ~x723 & ~x726 & ~x731 & ~x732 & ~x735 & ~x739 & ~x742 & ~x743 & ~x747 & ~x764 & ~x766 & ~x768 & ~x769 & ~x774 & ~x775 & ~x776 & ~x781 & ~x783;
assign c210 =  x485 & ~x11 & ~x25 & ~x27 & ~x28 & ~x34 & ~x47 & ~x61 & ~x64 & ~x68 & ~x82 & ~x87 & ~x93 & ~x95 & ~x104 & ~x114 & ~x136 & ~x140 & ~x141 & ~x145 & ~x147 & ~x164 & ~x191 & ~x199 & ~x201 & ~x202 & ~x203 & ~x221 & ~x222 & ~x223 & ~x225 & ~x226 & ~x227 & ~x229 & ~x230 & ~x231 & ~x249 & ~x252 & ~x255 & ~x279 & ~x285 & ~x293 & ~x311 & ~x314 & ~x318 & ~x333 & ~x335 & ~x343 & ~x361 & ~x392 & ~x473 & ~x479 & ~x528 & ~x529 & ~x588 & ~x615 & ~x649 & ~x650 & ~x668 & ~x669 & ~x674 & ~x685 & ~x690 & ~x691 & ~x693 & ~x699 & ~x707 & ~x715 & ~x716 & ~x723 & ~x731 & ~x735 & ~x746 & ~x747 & ~x750 & ~x752 & ~x763 & ~x764 & ~x772 & ~x783;
assign c212 =  x543 &  x577 & ~x291 & ~x315 & ~x321 & ~x506 & ~x586;
assign c214 =  x667;
assign c216 =  x641;
assign c218 = ~x0 & ~x2 & ~x3 & ~x6 & ~x7 & ~x8 & ~x9 & ~x10 & ~x15 & ~x16 & ~x19 & ~x21 & ~x25 & ~x28 & ~x29 & ~x36 & ~x39 & ~x41 & ~x45 & ~x46 & ~x47 & ~x50 & ~x56 & ~x59 & ~x61 & ~x62 & ~x64 & ~x70 & ~x80 & ~x81 & ~x83 & ~x85 & ~x87 & ~x88 & ~x89 & ~x90 & ~x92 & ~x94 & ~x95 & ~x97 & ~x98 & ~x103 & ~x105 & ~x106 & ~x108 & ~x110 & ~x112 & ~x115 & ~x122 & ~x123 & ~x133 & ~x135 & ~x136 & ~x140 & ~x142 & ~x145 & ~x150 & ~x155 & ~x158 & ~x162 & ~x163 & ~x165 & ~x166 & ~x169 & ~x172 & ~x176 & ~x188 & ~x189 & ~x191 & ~x195 & ~x198 & ~x200 & ~x216 & ~x217 & ~x218 & ~x219 & ~x224 & ~x251 & ~x254 & ~x277 & ~x278 & ~x305 & ~x307 & ~x308 & ~x334 & ~x336 & ~x337 & ~x338 & ~x366 & ~x369 & ~x392 & ~x395 & ~x396 & ~x448 & ~x449 & ~x450 & ~x451 & ~x476 & ~x477 & ~x503 & ~x505 & ~x533 & ~x535 & ~x574 & ~x575 & ~x576 & ~x580 & ~x581 & ~x582 & ~x583 & ~x587 & ~x591 & ~x593 & ~x600 & ~x601 & ~x602 & ~x603 & ~x604 & ~x605 & ~x606 & ~x607 & ~x608 & ~x609 & ~x610 & ~x611 & ~x612 & ~x613 & ~x616 & ~x624 & ~x625 & ~x626 & ~x627 & ~x628 & ~x632 & ~x634 & ~x635 & ~x636 & ~x639 & ~x644 & ~x646 & ~x648 & ~x651 & ~x652 & ~x653 & ~x654 & ~x655 & ~x656 & ~x659 & ~x661 & ~x662 & ~x663 & ~x665 & ~x666 & ~x667 & ~x668 & ~x670 & ~x671 & ~x677 & ~x678 & ~x681 & ~x682 & ~x683 & ~x685 & ~x687 & ~x688 & ~x690 & ~x691 & ~x693 & ~x694 & ~x695 & ~x700 & ~x701 & ~x702 & ~x712 & ~x715 & ~x716 & ~x720 & ~x724 & ~x725 & ~x727 & ~x728 & ~x729 & ~x730 & ~x732 & ~x733 & ~x735 & ~x740 & ~x741 & ~x742 & ~x745 & ~x747 & ~x750 & ~x754 & ~x757 & ~x759 & ~x763 & ~x766 & ~x772 & ~x773 & ~x775 & ~x780 & ~x781 & ~x782;
assign c220 =  x151 &  x210 & ~x23 & ~x98 & ~x100 & ~x113 & ~x138 & ~x244 & ~x250 & ~x275 & ~x281 & ~x318 & ~x362 & ~x366 & ~x369 & ~x422 & ~x558 & ~x621 & ~x643 & ~x677 & ~x709 & ~x717 & ~x769;
assign c222 =  x418;
assign c224 = ~x0 & ~x6 & ~x7 & ~x10 & ~x16 & ~x23 & ~x29 & ~x30 & ~x33 & ~x39 & ~x42 & ~x43 & ~x46 & ~x49 & ~x58 & ~x61 & ~x63 & ~x68 & ~x74 & ~x75 & ~x76 & ~x79 & ~x84 & ~x85 & ~x115 & ~x116 & ~x117 & ~x119 & ~x137 & ~x138 & ~x140 & ~x144 & ~x165 & ~x171 & ~x192 & ~x199 & ~x248 & ~x254 & ~x276 & ~x280 & ~x284 & ~x288 & ~x309 & ~x311 & ~x312 & ~x315 & ~x333 & ~x334 & ~x336 & ~x340 & ~x353 & ~x363 & ~x366 & ~x369 & ~x370 & ~x374 & ~x380 & ~x397 & ~x407 & ~x420 & ~x421 & ~x447 & ~x477 & ~x500 & ~x501 & ~x530 & ~x561 & ~x562 & ~x588 & ~x613 & ~x617 & ~x618 & ~x641 & ~x643 & ~x645 & ~x666 & ~x667 & ~x669 & ~x670 & ~x671 & ~x685 & ~x689 & ~x692 & ~x700 & ~x704 & ~x707 & ~x709 & ~x713 & ~x715 & ~x717 & ~x718 & ~x720 & ~x725 & ~x727 & ~x728 & ~x729 & ~x731 & ~x734 & ~x736 & ~x737 & ~x743 & ~x746 & ~x749 & ~x751 & ~x754 & ~x756 & ~x757 & ~x758 & ~x760 & ~x761 & ~x763 & ~x765 & ~x769 & ~x773 & ~x777 & ~x783;
assign c226 =  x473;
assign c228 =  x731;
assign c230 =  x403 & ~x5 & ~x8 & ~x11 & ~x12 & ~x26 & ~x29 & ~x35 & ~x41 & ~x44 & ~x45 & ~x46 & ~x47 & ~x51 & ~x53 & ~x54 & ~x56 & ~x58 & ~x75 & ~x76 & ~x90 & ~x107 & ~x108 & ~x118 & ~x136 & ~x139 & ~x142 & ~x146 & ~x147 & ~x168 & ~x170 & ~x191 & ~x193 & ~x197 & ~x200 & ~x224 & ~x249 & ~x251 & ~x276 & ~x277 & ~x278 & ~x287 & ~x304 & ~x313 & ~x317 & ~x319 & ~x320 & ~x336 & ~x363 & ~x393 & ~x418 & ~x422 & ~x503 & ~x504 & ~x588 & ~x643 & ~x644 & ~x645 & ~x646 & ~x650 & ~x658 & ~x668 & ~x669 & ~x673 & ~x674 & ~x677 & ~x678 & ~x679 & ~x680 & ~x681 & ~x682 & ~x684 & ~x686 & ~x692 & ~x698 & ~x703 & ~x715 & ~x717 & ~x720 & ~x740 & ~x744 & ~x749 & ~x762 & ~x767 & ~x776;
assign c232 = ~x1 & ~x7 & ~x22 & ~x24 & ~x25 & ~x35 & ~x36 & ~x37 & ~x53 & ~x55 & ~x56 & ~x58 & ~x62 & ~x72 & ~x86 & ~x103 & ~x105 & ~x109 & ~x161 & ~x168 & ~x187 & ~x190 & ~x196 & ~x223 & ~x227 & ~x255 & ~x273 & ~x291 & ~x300 & ~x302 & ~x307 & ~x313 & ~x317 & ~x320 & ~x329 & ~x337 & ~x340 & ~x342 & ~x344 & ~x364 & ~x477 & ~x479 & ~x504 & ~x506 & ~x508 & ~x509 & ~x529 & ~x531 & ~x532 & ~x536 & ~x558 & ~x586 & ~x593 & ~x618 & ~x639 & ~x650 & ~x653 & ~x654 & ~x656 & ~x667 & ~x673 & ~x675 & ~x678 & ~x687 & ~x689 & ~x700 & ~x702 & ~x706 & ~x707 & ~x708 & ~x713 & ~x716 & ~x720 & ~x741 & ~x742 & ~x745 & ~x761 & ~x774 & ~x780 & ~x781 & ~x783;
assign c234 =  x281;
assign c236 =  x306 &  x420;
assign c238 = ~x7 & ~x13 & ~x16 & ~x18 & ~x20 & ~x22 & ~x23 & ~x24 & ~x28 & ~x31 & ~x35 & ~x38 & ~x39 & ~x40 & ~x44 & ~x46 & ~x48 & ~x50 & ~x54 & ~x57 & ~x59 & ~x63 & ~x66 & ~x78 & ~x82 & ~x92 & ~x93 & ~x109 & ~x110 & ~x112 & ~x113 & ~x116 & ~x138 & ~x139 & ~x140 & ~x141 & ~x144 & ~x145 & ~x146 & ~x165 & ~x194 & ~x195 & ~x196 & ~x199 & ~x221 & ~x224 & ~x227 & ~x252 & ~x253 & ~x277 & ~x278 & ~x282 & ~x286 & ~x307 & ~x314 & ~x316 & ~x317 & ~x318 & ~x319 & ~x321 & ~x323 & ~x324 & ~x335 & ~x337 & ~x338 & ~x340 & ~x341 & ~x343 & ~x351 & ~x361 & ~x362 & ~x363 & ~x364 & ~x365 & ~x366 & ~x392 & ~x394 & ~x396 & ~x417 & ~x418 & ~x421 & ~x450 & ~x472 & ~x475 & ~x503 & ~x505 & ~x507 & ~x531 & ~x535 & ~x557 & ~x559 & ~x561 & ~x583 & ~x585 & ~x589 & ~x612 & ~x640 & ~x666 & ~x670 & ~x680 & ~x690 & ~x695 & ~x697 & ~x700 & ~x701 & ~x702 & ~x704 & ~x706 & ~x707 & ~x710 & ~x711 & ~x712 & ~x720 & ~x723 & ~x726 & ~x727 & ~x730 & ~x731 & ~x732 & ~x734 & ~x735 & ~x736 & ~x740 & ~x745 & ~x748 & ~x752 & ~x756 & ~x763 & ~x768 & ~x769 & ~x771 & ~x773 & ~x774 & ~x777 & ~x779 & ~x781 & ~x783;
assign c240 =  x464 & ~x1 & ~x2 & ~x9 & ~x10 & ~x16 & ~x17 & ~x22 & ~x23 & ~x25 & ~x28 & ~x29 & ~x30 & ~x34 & ~x38 & ~x41 & ~x42 & ~x45 & ~x48 & ~x51 & ~x53 & ~x54 & ~x57 & ~x58 & ~x59 & ~x61 & ~x62 & ~x63 & ~x69 & ~x70 & ~x73 & ~x74 & ~x75 & ~x76 & ~x79 & ~x80 & ~x83 & ~x86 & ~x87 & ~x88 & ~x90 & ~x91 & ~x106 & ~x109 & ~x110 & ~x111 & ~x113 & ~x114 & ~x117 & ~x118 & ~x131 & ~x132 & ~x135 & ~x139 & ~x146 & ~x148 & ~x161 & ~x165 & ~x166 & ~x169 & ~x170 & ~x171 & ~x174 & ~x175 & ~x189 & ~x192 & ~x197 & ~x198 & ~x216 & ~x217 & ~x219 & ~x220 & ~x221 & ~x222 & ~x223 & ~x228 & ~x254 & ~x255 & ~x280 & ~x281 & ~x305 & ~x307 & ~x311 & ~x335 & ~x339 & ~x365 & ~x368 & ~x393 & ~x394 & ~x419 & ~x421 & ~x451 & ~x474 & ~x503 & ~x505 & ~x506 & ~x507 & ~x508 & ~x531 & ~x532 & ~x534 & ~x535 & ~x558 & ~x561 & ~x577 & ~x578 & ~x593 & ~x604 & ~x606 & ~x616 & ~x618 & ~x619 & ~x621 & ~x622 & ~x623 & ~x634 & ~x635 & ~x639 & ~x642 & ~x645 & ~x646 & ~x649 & ~x650 & ~x654 & ~x656 & ~x657 & ~x659 & ~x660 & ~x661 & ~x662 & ~x664 & ~x666 & ~x669 & ~x670 & ~x672 & ~x673 & ~x680 & ~x684 & ~x688 & ~x689 & ~x690 & ~x696 & ~x699 & ~x701 & ~x702 & ~x705 & ~x706 & ~x711 & ~x712 & ~x713 & ~x714 & ~x717 & ~x722 & ~x724 & ~x728 & ~x732 & ~x742 & ~x743 & ~x750 & ~x755 & ~x758 & ~x760 & ~x763 & ~x765 & ~x768 & ~x769 & ~x772 & ~x773 & ~x774 & ~x775 & ~x777 & ~x778 & ~x779 & ~x780 & ~x781;
assign c242 =  x152 &  x636 & ~x29 & ~x60 & ~x115 & ~x142 & ~x196 & ~x256 & ~x304 & ~x363 & ~x368 & ~x396 & ~x468 & ~x470 & ~x731 & ~x747;
assign c244 =  x770;
assign c246 =  x583 & ~x499;
assign c248 =  x363;
assign c250 = ~x1 & ~x8 & ~x9 & ~x34 & ~x39 & ~x45 & ~x46 & ~x47 & ~x52 & ~x66 & ~x68 & ~x72 & ~x76 & ~x78 & ~x84 & ~x87 & ~x92 & ~x96 & ~x100 & ~x103 & ~x104 & ~x114 & ~x116 & ~x136 & ~x140 & ~x141 & ~x142 & ~x144 & ~x145 & ~x147 & ~x159 & ~x169 & ~x170 & ~x188 & ~x189 & ~x191 & ~x193 & ~x195 & ~x196 & ~x220 & ~x244 & ~x246 & ~x255 & ~x274 & ~x275 & ~x301 & ~x311 & ~x329 & ~x331 & ~x332 & ~x339 & ~x356 & ~x358 & ~x363 & ~x365 & ~x377 & ~x390 & ~x404 & ~x413 & ~x417 & ~x442 & ~x445 & ~x455 & ~x457 & ~x458 & ~x467 & ~x468 & ~x505 & ~x508 & ~x512 & ~x513 & ~x530 & ~x534 & ~x536 & ~x558 & ~x562 & ~x587 & ~x588 & ~x589 & ~x590 & ~x622 & ~x650 & ~x667 & ~x672 & ~x679 & ~x705 & ~x711 & ~x713 & ~x720 & ~x728 & ~x745 & ~x749 & ~x759 & ~x765 & ~x767 & ~x776 & ~x781;
assign c252 = ~x0 & ~x6 & ~x7 & ~x8 & ~x20 & ~x22 & ~x23 & ~x25 & ~x35 & ~x39 & ~x40 & ~x42 & ~x46 & ~x56 & ~x60 & ~x63 & ~x64 & ~x79 & ~x80 & ~x83 & ~x86 & ~x89 & ~x112 & ~x113 & ~x114 & ~x115 & ~x166 & ~x168 & ~x199 & ~x223 & ~x224 & ~x225 & ~x231 & ~x254 & ~x258 & ~x260 & ~x284 & ~x285 & ~x286 & ~x287 & ~x289 & ~x305 & ~x312 & ~x314 & ~x317 & ~x319 & ~x320 & ~x321 & ~x324 & ~x339 & ~x366 & ~x367 & ~x389 & ~x391 & ~x417 & ~x423 & ~x443 & ~x446 & ~x471 & ~x477 & ~x502 & ~x503 & ~x506 & ~x531 & ~x534 & ~x556 & ~x588 & ~x590 & ~x618 & ~x619 & ~x643 & ~x644 & ~x645 & ~x646 & ~x664 & ~x665 & ~x668 & ~x677 & ~x683 & ~x690 & ~x702 & ~x705 & ~x706 & ~x710 & ~x715 & ~x716 & ~x719 & ~x721 & ~x724 & ~x727 & ~x739 & ~x759 & ~x765 & ~x778 & ~x782 & ~x783;
assign c254 =  x779;
assign c256 =  x558;
assign c258 =  x561;
assign c260 =  x429 & ~x3 & ~x11 & ~x15 & ~x17 & ~x19 & ~x20 & ~x29 & ~x36 & ~x44 & ~x45 & ~x59 & ~x60 & ~x62 & ~x63 & ~x66 & ~x67 & ~x68 & ~x72 & ~x75 & ~x77 & ~x80 & ~x81 & ~x86 & ~x88 & ~x91 & ~x107 & ~x111 & ~x113 & ~x114 & ~x115 & ~x137 & ~x139 & ~x141 & ~x142 & ~x145 & ~x164 & ~x172 & ~x173 & ~x174 & ~x193 & ~x199 & ~x220 & ~x221 & ~x223 & ~x227 & ~x250 & ~x252 & ~x276 & ~x277 & ~x285 & ~x306 & ~x309 & ~x310 & ~x311 & ~x312 & ~x313 & ~x314 & ~x315 & ~x332 & ~x336 & ~x337 & ~x338 & ~x342 & ~x344 & ~x346 & ~x363 & ~x369 & ~x370 & ~x391 & ~x396 & ~x420 & ~x421 & ~x422 & ~x423 & ~x444 & ~x449 & ~x477 & ~x478 & ~x506 & ~x533 & ~x534 & ~x556 & ~x559 & ~x560 & ~x562 & ~x587 & ~x588 & ~x590 & ~x613 & ~x619 & ~x640 & ~x642 & ~x647 & ~x660 & ~x667 & ~x668 & ~x671 & ~x672 & ~x675 & ~x677 & ~x680 & ~x682 & ~x683 & ~x684 & ~x687 & ~x688 & ~x689 & ~x691 & ~x692 & ~x695 & ~x699 & ~x700 & ~x701 & ~x702 & ~x704 & ~x705 & ~x706 & ~x709 & ~x710 & ~x711 & ~x713 & ~x716 & ~x719 & ~x725 & ~x727 & ~x728 & ~x730 & ~x731 & ~x737 & ~x739 & ~x740 & ~x747 & ~x749 & ~x751 & ~x753 & ~x755 & ~x762 & ~x763 & ~x769 & ~x770 & ~x771 & ~x775 & ~x781 & ~x782 & ~x783;
assign c262 =  x486 & ~x1 & ~x2 & ~x3 & ~x10 & ~x11 & ~x22 & ~x23 & ~x34 & ~x42 & ~x44 & ~x47 & ~x51 & ~x54 & ~x57 & ~x59 & ~x60 & ~x84 & ~x87 & ~x221 & ~x222 & ~x230 & ~x252 & ~x256 & ~x277 & ~x321 & ~x347 & ~x348 & ~x365 & ~x373 & ~x374 & ~x389 & ~x400 & ~x401 & ~x423 & ~x426 & ~x427 & ~x448 & ~x656 & ~x682 & ~x685 & ~x688 & ~x699 & ~x707 & ~x711 & ~x717 & ~x721 & ~x733 & ~x744 & ~x745 & ~x769 & ~x770 & ~x781;
assign c264 =  x514 & ~x1 & ~x10 & ~x12 & ~x16 & ~x22 & ~x32 & ~x36 & ~x44 & ~x56 & ~x60 & ~x64 & ~x67 & ~x77 & ~x83 & ~x84 & ~x88 & ~x102 & ~x104 & ~x115 & ~x136 & ~x137 & ~x139 & ~x161 & ~x164 & ~x167 & ~x172 & ~x173 & ~x189 & ~x194 & ~x220 & ~x226 & ~x227 & ~x256 & ~x274 & ~x275 & ~x278 & ~x279 & ~x280 & ~x281 & ~x285 & ~x292 & ~x302 & ~x305 & ~x307 & ~x312 & ~x319 & ~x328 & ~x341 & ~x343 & ~x345 & ~x346 & ~x397 & ~x420 & ~x448 & ~x450 & ~x451 & ~x476 & ~x479 & ~x480 & ~x502 & ~x503 & ~x558 & ~x588 & ~x613 & ~x620 & ~x641 & ~x650 & ~x667 & ~x670 & ~x671 & ~x672 & ~x676 & ~x678 & ~x685 & ~x686 & ~x688 & ~x691 & ~x696 & ~x697 & ~x703 & ~x705 & ~x708 & ~x710 & ~x711 & ~x712 & ~x713 & ~x715 & ~x716 & ~x720 & ~x721 & ~x726 & ~x727 & ~x728 & ~x729 & ~x733 & ~x741 & ~x746 & ~x760 & ~x764 & ~x765 & ~x767 & ~x768 & ~x771 & ~x774 & ~x778;
assign c266 =  x180 & ~x29 & ~x31 & ~x32 & ~x56 & ~x72 & ~x83 & ~x92 & ~x112 & ~x118 & ~x128 & ~x138 & ~x193 & ~x199 & ~x245 & ~x308 & ~x321 & ~x335 & ~x349 & ~x358 & ~x375 & ~x376 & ~x377 & ~x399 & ~x404 & ~x426 & ~x429 & ~x430 & ~x432 & ~x455 & ~x456 & ~x459 & ~x481 & ~x510 & ~x511 & ~x512 & ~x530 & ~x537 & ~x567 & ~x650 & ~x651 & ~x679 & ~x680 & ~x699 & ~x727 & ~x753 & ~x759 & ~x766 & ~x772;
assign c268 =  x404 & ~x1 & ~x2 & ~x4 & ~x8 & ~x17 & ~x26 & ~x28 & ~x29 & ~x42 & ~x44 & ~x57 & ~x63 & ~x64 & ~x76 & ~x107 & ~x136 & ~x139 & ~x166 & ~x173 & ~x199 & ~x221 & ~x229 & ~x253 & ~x254 & ~x257 & ~x258 & ~x281 & ~x288 & ~x289 & ~x292 & ~x293 & ~x307 & ~x318 & ~x338 & ~x416 & ~x417 & ~x445 & ~x504 & ~x561 & ~x639 & ~x649 & ~x653 & ~x656 & ~x663 & ~x679 & ~x680 & ~x686 & ~x691 & ~x713 & ~x723 & ~x726 & ~x728 & ~x730 & ~x731 & ~x735 & ~x753 & ~x767 & ~x770 & ~x778;
assign c270 =  x82;
assign c272 = ~x3 & ~x4 & ~x8 & ~x9 & ~x10 & ~x13 & ~x14 & ~x16 & ~x23 & ~x31 & ~x32 & ~x34 & ~x37 & ~x45 & ~x51 & ~x52 & ~x59 & ~x63 & ~x65 & ~x75 & ~x79 & ~x80 & ~x81 & ~x86 & ~x90 & ~x104 & ~x114 & ~x116 & ~x135 & ~x136 & ~x139 & ~x141 & ~x168 & ~x169 & ~x192 & ~x199 & ~x224 & ~x225 & ~x227 & ~x248 & ~x255 & ~x261 & ~x265 & ~x277 & ~x279 & ~x293 & ~x295 & ~x306 & ~x316 & ~x319 & ~x332 & ~x335 & ~x338 & ~x340 & ~x342 & ~x343 & ~x350 & ~x361 & ~x362 & ~x364 & ~x365 & ~x368 & ~x390 & ~x391 & ~x395 & ~x418 & ~x419 & ~x446 & ~x447 & ~x449 & ~x476 & ~x506 & ~x530 & ~x531 & ~x533 & ~x589 & ~x611 & ~x646 & ~x648 & ~x668 & ~x678 & ~x680 & ~x681 & ~x683 & ~x687 & ~x688 & ~x692 & ~x703 & ~x704 & ~x711 & ~x713 & ~x717 & ~x718 & ~x724 & ~x727 & ~x728 & ~x730 & ~x731 & ~x738 & ~x739 & ~x740 & ~x745 & ~x753 & ~x757 & ~x761 & ~x763 & ~x768 & ~x778 & ~x779 & ~x782;
assign c276 =  x493 & ~x2 & ~x8 & ~x14 & ~x15 & ~x18 & ~x20 & ~x25 & ~x28 & ~x32 & ~x37 & ~x38 & ~x39 & ~x46 & ~x47 & ~x50 & ~x59 & ~x71 & ~x74 & ~x79 & ~x93 & ~x117 & ~x133 & ~x134 & ~x142 & ~x167 & ~x168 & ~x171 & ~x190 & ~x194 & ~x228 & ~x253 & ~x274 & ~x280 & ~x281 & ~x310 & ~x311 & ~x313 & ~x331 & ~x332 & ~x335 & ~x357 & ~x358 & ~x360 & ~x385 & ~x387 & ~x392 & ~x396 & ~x422 & ~x424 & ~x449 & ~x452 & ~x480 & ~x504 & ~x506 & ~x576 & ~x577 & ~x587 & ~x603 & ~x604 & ~x606 & ~x612 & ~x614 & ~x632 & ~x634 & ~x636 & ~x640 & ~x646 & ~x658 & ~x659 & ~x661 & ~x662 & ~x664 & ~x665 & ~x669 & ~x670 & ~x676 & ~x682 & ~x683 & ~x684 & ~x685 & ~x687 & ~x688 & ~x689 & ~x692 & ~x694 & ~x703 & ~x709 & ~x712 & ~x713 & ~x716 & ~x717 & ~x723 & ~x730 & ~x732 & ~x735 & ~x745 & ~x749 & ~x755 & ~x756 & ~x757 & ~x758 & ~x763 & ~x764 & ~x771 & ~x779;
assign c278 = ~x31 & ~x84 & ~x263 & ~x281 & ~x289 & ~x294 & ~x319 & ~x323 & ~x340 & ~x343 & ~x349 & ~x350 & ~x390 & ~x432 & ~x442 & ~x444 & ~x474 & ~x501 & ~x527 & ~x595 & ~x621 & ~x679 & ~x708 & ~x730;
assign c280 =  x154 &  x180 &  x625 &  x626 &  x654 & ~x49 & ~x87 & ~x140 & ~x221 & ~x248 & ~x249 & ~x350 & ~x361 & ~x395 & ~x402 & ~x403 & ~x404 & ~x424 & ~x444 & ~x452 & ~x456 & ~x482 & ~x563 & ~x722 & ~x737;
assign c282 =  x389;
assign c284 =  x756;
assign c286 =  x512 & ~x0 & ~x9 & ~x11 & ~x17 & ~x26 & ~x27 & ~x34 & ~x41 & ~x48 & ~x51 & ~x62 & ~x63 & ~x79 & ~x84 & ~x93 & ~x107 & ~x109 & ~x144 & ~x145 & ~x166 & ~x190 & ~x194 & ~x196 & ~x200 & ~x202 & ~x220 & ~x249 & ~x252 & ~x253 & ~x255 & ~x289 & ~x293 & ~x306 & ~x307 & ~x308 & ~x313 & ~x317 & ~x335 & ~x340 & ~x342 & ~x343 & ~x363 & ~x395 & ~x420 & ~x476 & ~x503 & ~x584 & ~x589 & ~x592 & ~x641 & ~x646 & ~x673 & ~x682 & ~x684 & ~x687 & ~x688 & ~x690 & ~x700 & ~x701 & ~x702 & ~x711 & ~x713 & ~x724 & ~x731 & ~x734 & ~x738 & ~x741 & ~x745 & ~x746 & ~x747 & ~x750 & ~x752 & ~x755 & ~x760 & ~x762 & ~x769 & ~x779;
assign c288 =  x487 &  x545 & ~x4 & ~x6 & ~x28 & ~x29 & ~x38 & ~x54 & ~x78 & ~x84 & ~x91 & ~x94 & ~x111 & ~x113 & ~x117 & ~x135 & ~x197 & ~x202 & ~x225 & ~x248 & ~x331 & ~x335 & ~x347 & ~x373 & ~x392 & ~x393 & ~x395 & ~x398 & ~x429 & ~x559 & ~x588 & ~x655 & ~x682 & ~x705 & ~x706 & ~x712 & ~x728 & ~x731 & ~x736 & ~x746 & ~x750;
assign c290 =  x434 &  x490 &  x491 & ~x0 & ~x2 & ~x5 & ~x7 & ~x8 & ~x9 & ~x12 & ~x14 & ~x16 & ~x18 & ~x19 & ~x20 & ~x23 & ~x27 & ~x30 & ~x36 & ~x38 & ~x39 & ~x40 & ~x41 & ~x42 & ~x43 & ~x53 & ~x54 & ~x55 & ~x59 & ~x61 & ~x62 & ~x65 & ~x66 & ~x68 & ~x70 & ~x71 & ~x74 & ~x77 & ~x79 & ~x80 & ~x81 & ~x83 & ~x85 & ~x86 & ~x108 & ~x109 & ~x110 & ~x112 & ~x115 & ~x116 & ~x118 & ~x119 & ~x120 & ~x135 & ~x136 & ~x137 & ~x138 & ~x143 & ~x145 & ~x146 & ~x148 & ~x164 & ~x165 & ~x171 & ~x173 & ~x192 & ~x193 & ~x202 & ~x220 & ~x225 & ~x228 & ~x229 & ~x248 & ~x250 & ~x251 & ~x253 & ~x256 & ~x259 & ~x277 & ~x278 & ~x283 & ~x285 & ~x312 & ~x332 & ~x336 & ~x337 & ~x340 & ~x364 & ~x365 & ~x391 & ~x392 & ~x393 & ~x414 & ~x416 & ~x419 & ~x444 & ~x448 & ~x449 & ~x471 & ~x474 & ~x476 & ~x478 & ~x501 & ~x504 & ~x534 & ~x558 & ~x562 & ~x586 & ~x587 & ~x588 & ~x589 & ~x616 & ~x619 & ~x628 & ~x630 & ~x639 & ~x642 & ~x644 & ~x645 & ~x652 & ~x657 & ~x658 & ~x669 & ~x670 & ~x671 & ~x673 & ~x674 & ~x677 & ~x679 & ~x681 & ~x682 & ~x683 & ~x686 & ~x695 & ~x696 & ~x697 & ~x699 & ~x705 & ~x706 & ~x707 & ~x708 & ~x716 & ~x718 & ~x723 & ~x726 & ~x727 & ~x728 & ~x729 & ~x731 & ~x735 & ~x741 & ~x742 & ~x744 & ~x747 & ~x749 & ~x750 & ~x751 & ~x752 & ~x754 & ~x755 & ~x756 & ~x758 & ~x760 & ~x761 & ~x763 & ~x768 & ~x769 & ~x775 & ~x776 & ~x778 & ~x781 & ~x783;
assign c292 =  x525 & ~x13 & ~x107 & ~x134 & ~x190 & ~x228 & ~x256 & ~x277 & ~x308 & ~x333 & ~x336 & ~x339 & ~x357 & ~x358 & ~x416 & ~x439 & ~x536 & ~x613 & ~x667 & ~x674 & ~x686 & ~x689 & ~x692 & ~x733;
assign c294 = ~x2 & ~x3 & ~x10 & ~x12 & ~x13 & ~x15 & ~x17 & ~x20 & ~x21 & ~x22 & ~x23 & ~x25 & ~x26 & ~x27 & ~x28 & ~x31 & ~x41 & ~x42 & ~x44 & ~x53 & ~x62 & ~x66 & ~x71 & ~x72 & ~x73 & ~x74 & ~x76 & ~x78 & ~x82 & ~x84 & ~x88 & ~x89 & ~x92 & ~x97 & ~x99 & ~x101 & ~x102 & ~x103 & ~x107 & ~x110 & ~x113 & ~x115 & ~x120 & ~x136 & ~x138 & ~x139 & ~x140 & ~x145 & ~x163 & ~x164 & ~x193 & ~x194 & ~x196 & ~x198 & ~x220 & ~x221 & ~x223 & ~x227 & ~x253 & ~x276 & ~x277 & ~x282 & ~x305 & ~x309 & ~x333 & ~x346 & ~x347 & ~x348 & ~x349 & ~x351 & ~x364 & ~x366 & ~x367 & ~x368 & ~x371 & ~x372 & ~x373 & ~x374 & ~x391 & ~x397 & ~x398 & ~x420 & ~x423 & ~x445 & ~x447 & ~x452 & ~x477 & ~x502 & ~x503 & ~x505 & ~x507 & ~x529 & ~x531 & ~x534 & ~x557 & ~x562 & ~x585 & ~x587 & ~x589 & ~x612 & ~x616 & ~x617 & ~x618 & ~x645 & ~x648 & ~x666 & ~x667 & ~x673 & ~x674 & ~x675 & ~x677 & ~x678 & ~x681 & ~x682 & ~x684 & ~x685 & ~x689 & ~x694 & ~x696 & ~x698 & ~x699 & ~x702 & ~x705 & ~x707 & ~x709 & ~x713 & ~x714 & ~x715 & ~x716 & ~x718 & ~x722 & ~x723 & ~x724 & ~x731 & ~x732 & ~x733 & ~x734 & ~x735 & ~x736 & ~x737 & ~x738 & ~x739 & ~x740 & ~x742 & ~x746 & ~x749 & ~x750 & ~x751 & ~x755 & ~x756 & ~x757 & ~x762 & ~x766 & ~x767 & ~x769 & ~x770 & ~x771 & ~x772 & ~x773 & ~x774 & ~x775 & ~x779 & ~x782 & ~x783;
assign c296 =  x155 &  x465 &  x492 & ~x53 & ~x168 & ~x294 & ~x352 & ~x395;
assign c298 =  x182 &  x516 & ~x80 & ~x101 & ~x102 & ~x171 & ~x173 & ~x221 & ~x274 & ~x320 & ~x374 & ~x426 & ~x456 & ~x644 & ~x680;
assign c2100 =  x460 & ~x34 & ~x62 & ~x91 & ~x145 & ~x165 & ~x265 & ~x292 & ~x306 & ~x321 & ~x375 & ~x391 & ~x401 & ~x454 & ~x722;
assign c2102 =  x459 &  x485 & ~x6 & ~x14 & ~x23 & ~x25 & ~x33 & ~x34 & ~x51 & ~x53 & ~x60 & ~x65 & ~x80 & ~x85 & ~x87 & ~x104 & ~x114 & ~x115 & ~x135 & ~x136 & ~x143 & ~x144 & ~x168 & ~x171 & ~x193 & ~x199 & ~x200 & ~x219 & ~x249 & ~x285 & ~x302 & ~x303 & ~x304 & ~x309 & ~x311 & ~x312 & ~x313 & ~x341 & ~x342 & ~x358 & ~x369 & ~x387 & ~x388 & ~x391 & ~x414 & ~x421 & ~x439 & ~x450 & ~x531 & ~x533 & ~x559 & ~x619 & ~x642 & ~x643 & ~x657 & ~x672 & ~x677 & ~x680 & ~x682 & ~x709 & ~x713 & ~x715 & ~x717 & ~x718 & ~x719 & ~x721 & ~x737 & ~x738 & ~x744 & ~x746 & ~x765 & ~x773 & ~x775 & ~x777 & ~x780 & ~x781 & ~x782;
assign c2104 =  x545 &  x571 &  x572 &  x598 &  x599 & ~x2 & ~x5 & ~x7 & ~x8 & ~x18 & ~x25 & ~x26 & ~x27 & ~x38 & ~x39 & ~x45 & ~x46 & ~x47 & ~x54 & ~x59 & ~x60 & ~x63 & ~x65 & ~x67 & ~x70 & ~x71 & ~x76 & ~x77 & ~x78 & ~x80 & ~x81 & ~x88 & ~x90 & ~x92 & ~x104 & ~x110 & ~x112 & ~x117 & ~x120 & ~x134 & ~x135 & ~x140 & ~x144 & ~x162 & ~x164 & ~x169 & ~x171 & ~x172 & ~x191 & ~x197 & ~x219 & ~x222 & ~x223 & ~x225 & ~x248 & ~x276 & ~x304 & ~x306 & ~x311 & ~x312 & ~x323 & ~x324 & ~x331 & ~x332 & ~x337 & ~x351 & ~x359 & ~x360 & ~x387 & ~x392 & ~x397 & ~x415 & ~x422 & ~x442 & ~x443 & ~x470 & ~x472 & ~x475 & ~x477 & ~x502 & ~x503 & ~x557 & ~x588 & ~x617 & ~x619 & ~x644 & ~x669 & ~x671 & ~x673 & ~x687 & ~x691 & ~x697 & ~x698 & ~x702 & ~x708 & ~x709 & ~x717 & ~x725 & ~x726 & ~x728 & ~x730 & ~x731 & ~x735 & ~x737 & ~x738 & ~x741 & ~x745 & ~x748 & ~x749 & ~x750 & ~x756 & ~x758 & ~x759 & ~x761 & ~x763 & ~x765 & ~x771 & ~x778;
assign c2106 =  x458 & ~x5 & ~x8 & ~x10 & ~x12 & ~x14 & ~x16 & ~x19 & ~x20 & ~x23 & ~x37 & ~x38 & ~x42 & ~x47 & ~x51 & ~x53 & ~x67 & ~x73 & ~x83 & ~x108 & ~x115 & ~x117 & ~x122 & ~x123 & ~x134 & ~x135 & ~x137 & ~x140 & ~x141 & ~x143 & ~x165 & ~x171 & ~x173 & ~x195 & ~x203 & ~x225 & ~x229 & ~x249 & ~x256 & ~x277 & ~x280 & ~x338 & ~x362 & ~x363 & ~x364 & ~x365 & ~x371 & ~x373 & ~x374 & ~x394 & ~x396 & ~x397 & ~x400 & ~x401 & ~x419 & ~x424 & ~x425 & ~x475 & ~x477 & ~x534 & ~x562 & ~x585 & ~x587 & ~x609 & ~x611 & ~x629 & ~x630 & ~x638 & ~x639 & ~x641 & ~x642 & ~x644 & ~x646 & ~x655 & ~x658 & ~x666 & ~x667 & ~x669 & ~x670 & ~x673 & ~x674 & ~x678 & ~x680 & ~x682 & ~x684 & ~x685 & ~x687 & ~x690 & ~x693 & ~x694 & ~x695 & ~x697 & ~x698 & ~x703 & ~x706 & ~x710 & ~x711 & ~x714 & ~x718 & ~x719 & ~x723 & ~x725 & ~x726 & ~x727 & ~x735 & ~x744 & ~x753 & ~x754 & ~x757 & ~x759 & ~x765 & ~x768 & ~x773 & ~x779 & ~x780 & ~x782;
assign c2108 = ~x0 & ~x3 & ~x6 & ~x11 & ~x21 & ~x26 & ~x28 & ~x32 & ~x33 & ~x34 & ~x35 & ~x37 & ~x45 & ~x46 & ~x58 & ~x61 & ~x64 & ~x68 & ~x73 & ~x77 & ~x81 & ~x82 & ~x85 & ~x87 & ~x89 & ~x93 & ~x96 & ~x98 & ~x104 & ~x107 & ~x109 & ~x113 & ~x115 & ~x116 & ~x134 & ~x137 & ~x140 & ~x141 & ~x144 & ~x169 & ~x171 & ~x192 & ~x195 & ~x196 & ~x222 & ~x252 & ~x255 & ~x278 & ~x280 & ~x283 & ~x284 & ~x303 & ~x308 & ~x310 & ~x331 & ~x332 & ~x333 & ~x334 & ~x335 & ~x336 & ~x337 & ~x346 & ~x348 & ~x359 & ~x361 & ~x362 & ~x367 & ~x371 & ~x372 & ~x374 & ~x378 & ~x379 & ~x387 & ~x390 & ~x392 & ~x397 & ~x399 & ~x417 & ~x424 & ~x446 & ~x478 & ~x504 & ~x507 & ~x533 & ~x558 & ~x560 & ~x561 & ~x562 & ~x589 & ~x590 & ~x615 & ~x639 & ~x647 & ~x668 & ~x671 & ~x674 & ~x678 & ~x680 & ~x682 & ~x683 & ~x696 & ~x697 & ~x699 & ~x700 & ~x704 & ~x705 & ~x711 & ~x712 & ~x714 & ~x715 & ~x719 & ~x722 & ~x723 & ~x733 & ~x735 & ~x736 & ~x737 & ~x741 & ~x742 & ~x745 & ~x749 & ~x762 & ~x763 & ~x768 & ~x770 & ~x773 & ~x781;
assign c2110 = ~x0 & ~x1 & ~x5 & ~x6 & ~x8 & ~x13 & ~x15 & ~x28 & ~x31 & ~x39 & ~x45 & ~x46 & ~x47 & ~x49 & ~x52 & ~x54 & ~x60 & ~x62 & ~x63 & ~x65 & ~x68 & ~x69 & ~x71 & ~x75 & ~x77 & ~x78 & ~x79 & ~x81 & ~x94 & ~x107 & ~x108 & ~x110 & ~x135 & ~x137 & ~x138 & ~x143 & ~x144 & ~x163 & ~x164 & ~x167 & ~x192 & ~x196 & ~x198 & ~x219 & ~x221 & ~x223 & ~x224 & ~x277 & ~x281 & ~x305 & ~x307 & ~x308 & ~x311 & ~x322 & ~x336 & ~x337 & ~x338 & ~x347 & ~x348 & ~x349 & ~x367 & ~x369 & ~x370 & ~x373 & ~x378 & ~x394 & ~x395 & ~x396 & ~x399 & ~x418 & ~x419 & ~x422 & ~x448 & ~x449 & ~x476 & ~x477 & ~x478 & ~x506 & ~x532 & ~x533 & ~x534 & ~x558 & ~x586 & ~x587 & ~x589 & ~x591 & ~x592 & ~x619 & ~x638 & ~x640 & ~x644 & ~x645 & ~x648 & ~x665 & ~x667 & ~x670 & ~x673 & ~x678 & ~x679 & ~x683 & ~x684 & ~x686 & ~x687 & ~x688 & ~x691 & ~x695 & ~x696 & ~x697 & ~x698 & ~x707 & ~x709 & ~x710 & ~x711 & ~x712 & ~x715 & ~x716 & ~x720 & ~x725 & ~x726 & ~x741 & ~x745 & ~x746 & ~x748 & ~x754 & ~x757 & ~x758 & ~x762 & ~x764 & ~x765 & ~x769 & ~x772 & ~x780 & ~x782;
assign c2112 =  x157 &  x214 &  x271 &  x517 & ~x0 & ~x5 & ~x11 & ~x23 & ~x30 & ~x39 & ~x48 & ~x53 & ~x56 & ~x60 & ~x63 & ~x64 & ~x65 & ~x71 & ~x73 & ~x75 & ~x78 & ~x80 & ~x117 & ~x120 & ~x135 & ~x140 & ~x147 & ~x167 & ~x219 & ~x224 & ~x227 & ~x229 & ~x252 & ~x254 & ~x279 & ~x282 & ~x284 & ~x302 & ~x313 & ~x334 & ~x335 & ~x336 & ~x339 & ~x360 & ~x361 & ~x364 & ~x386 & ~x387 & ~x396 & ~x415 & ~x419 & ~x448 & ~x505 & ~x506 & ~x532 & ~x588 & ~x589 & ~x640 & ~x645 & ~x659 & ~x660 & ~x669 & ~x671 & ~x672 & ~x674 & ~x688 & ~x724 & ~x725 & ~x726 & ~x744 & ~x745 & ~x768 & ~x776 & ~x783;
assign c2114 =  x301 &  x464 &  x509 & ~x287 & ~x289 & ~x315 & ~x342;
assign c2116 =  x210 &  x211 &  x543 &  x599 & ~x2 & ~x37 & ~x38 & ~x48 & ~x52 & ~x65 & ~x70 & ~x74 & ~x81 & ~x98 & ~x99 & ~x102 & ~x171 & ~x225 & ~x255 & ~x276 & ~x333 & ~x335 & ~x336 & ~x349 & ~x364 & ~x402 & ~x417 & ~x421 & ~x455 & ~x476 & ~x481 & ~x499 & ~x503 & ~x505 & ~x508 & ~x564 & ~x590 & ~x614 & ~x615 & ~x643 & ~x645 & ~x646 & ~x667 & ~x668 & ~x669 & ~x673 & ~x677 & ~x679 & ~x680 & ~x708 & ~x724 & ~x729 & ~x733 & ~x735 & ~x750 & ~x756 & ~x757 & ~x758 & ~x763 & ~x771 & ~x777 & ~x779;
assign c2118 =  x391;
assign c2120 =  x405 &  x515 &  x539 & ~x315 & ~x316 & ~x630 & ~x632 & ~x633;
assign c2122 =  x700;
assign c2124 =  x526 & ~x4 & ~x13 & ~x22 & ~x41 & ~x52 & ~x59 & ~x64 & ~x73 & ~x75 & ~x78 & ~x80 & ~x89 & ~x106 & ~x113 & ~x142 & ~x144 & ~x169 & ~x170 & ~x190 & ~x191 & ~x197 & ~x200 & ~x220 & ~x223 & ~x224 & ~x225 & ~x227 & ~x228 & ~x248 & ~x252 & ~x275 & ~x278 & ~x281 & ~x284 & ~x303 & ~x330 & ~x331 & ~x359 & ~x361 & ~x366 & ~x385 & ~x386 & ~x387 & ~x389 & ~x394 & ~x413 & ~x414 & ~x417 & ~x425 & ~x449 & ~x480 & ~x532 & ~x534 & ~x559 & ~x609 & ~x611 & ~x635 & ~x636 & ~x637 & ~x641 & ~x644 & ~x645 & ~x660 & ~x665 & ~x667 & ~x682 & ~x685 & ~x688 & ~x690 & ~x692 & ~x693 & ~x711 & ~x713 & ~x714 & ~x716 & ~x717 & ~x719 & ~x720 & ~x732 & ~x734 & ~x738 & ~x742 & ~x753 & ~x757 & ~x781;
assign c2126 =  x429 &  x430 & ~x18 & ~x29 & ~x38 & ~x39 & ~x42 & ~x45 & ~x50 & ~x51 & ~x91 & ~x106 & ~x111 & ~x117 & ~x138 & ~x139 & ~x141 & ~x144 & ~x145 & ~x167 & ~x174 & ~x191 & ~x198 & ~x200 & ~x202 & ~x229 & ~x232 & ~x277 & ~x285 & ~x286 & ~x287 & ~x303 & ~x304 & ~x305 & ~x307 & ~x309 & ~x319 & ~x340 & ~x341 & ~x343 & ~x345 & ~x363 & ~x392 & ~x393 & ~x394 & ~x419 & ~x420 & ~x447 & ~x505 & ~x530 & ~x532 & ~x640 & ~x643 & ~x652 & ~x680 & ~x681 & ~x683 & ~x689 & ~x698 & ~x699 & ~x712 & ~x715 & ~x722 & ~x741 & ~x754 & ~x759 & ~x760 & ~x770 & ~x781;
assign c2128 =  x532;
assign c2130 =  x522 &  x546 & ~x0 & ~x3 & ~x6 & ~x8 & ~x9 & ~x11 & ~x16 & ~x21 & ~x23 & ~x26 & ~x30 & ~x31 & ~x32 & ~x33 & ~x34 & ~x37 & ~x38 & ~x46 & ~x48 & ~x49 & ~x56 & ~x61 & ~x62 & ~x64 & ~x68 & ~x77 & ~x81 & ~x83 & ~x84 & ~x86 & ~x87 & ~x88 & ~x89 & ~x90 & ~x92 & ~x99 & ~x101 & ~x106 & ~x107 & ~x110 & ~x111 & ~x113 & ~x114 & ~x117 & ~x119 & ~x136 & ~x137 & ~x140 & ~x142 & ~x145 & ~x146 & ~x162 & ~x164 & ~x166 & ~x168 & ~x191 & ~x192 & ~x194 & ~x196 & ~x197 & ~x198 & ~x199 & ~x218 & ~x223 & ~x247 & ~x248 & ~x252 & ~x254 & ~x255 & ~x277 & ~x278 & ~x279 & ~x302 & ~x308 & ~x311 & ~x330 & ~x331 & ~x333 & ~x336 & ~x361 & ~x362 & ~x367 & ~x386 & ~x387 & ~x413 & ~x420 & ~x421 & ~x424 & ~x448 & ~x477 & ~x478 & ~x479 & ~x503 & ~x505 & ~x506 & ~x533 & ~x534 & ~x557 & ~x559 & ~x563 & ~x587 & ~x589 & ~x618 & ~x619 & ~x631 & ~x634 & ~x645 & ~x647 & ~x659 & ~x662 & ~x663 & ~x669 & ~x672 & ~x683 & ~x684 & ~x686 & ~x687 & ~x688 & ~x689 & ~x690 & ~x691 & ~x694 & ~x695 & ~x697 & ~x700 & ~x703 & ~x706 & ~x708 & ~x709 & ~x710 & ~x712 & ~x713 & ~x715 & ~x717 & ~x719 & ~x720 & ~x721 & ~x725 & ~x726 & ~x730 & ~x736 & ~x743 & ~x744 & ~x755 & ~x760 & ~x763 & ~x764 & ~x766 & ~x770 & ~x772 & ~x776 & ~x778 & ~x781;
assign c2132 =  x327 &  x355 &  x463 &  x542 & ~x11 & ~x34 & ~x36 & ~x37 & ~x41 & ~x48 & ~x54 & ~x56 & ~x60 & ~x68 & ~x78 & ~x88 & ~x111 & ~x135 & ~x142 & ~x143 & ~x144 & ~x163 & ~x175 & ~x201 & ~x220 & ~x251 & ~x256 & ~x314 & ~x331 & ~x335 & ~x360 & ~x420 & ~x447 & ~x557 & ~x558 & ~x559 & ~x586 & ~x588 & ~x647 & ~x650 & ~x658 & ~x679 & ~x687 & ~x694 & ~x699 & ~x704 & ~x707 & ~x719 & ~x721 & ~x737 & ~x746 & ~x750 & ~x753 & ~x757 & ~x762 & ~x780;
assign c2134 = ~x5 & ~x6 & ~x7 & ~x9 & ~x11 & ~x14 & ~x24 & ~x25 & ~x37 & ~x42 & ~x58 & ~x76 & ~x83 & ~x89 & ~x112 & ~x114 & ~x136 & ~x140 & ~x169 & ~x199 & ~x221 & ~x223 & ~x248 & ~x254 & ~x280 & ~x285 & ~x287 & ~x294 & ~x306 & ~x310 & ~x312 & ~x315 & ~x317 & ~x319 & ~x321 & ~x332 & ~x338 & ~x341 & ~x359 & ~x362 & ~x367 & ~x380 & ~x394 & ~x417 & ~x421 & ~x447 & ~x475 & ~x476 & ~x500 & ~x533 & ~x534 & ~x563 & ~x587 & ~x619 & ~x620 & ~x640 & ~x641 & ~x673 & ~x680 & ~x699 & ~x706 & ~x711 & ~x712 & ~x714 & ~x720 & ~x726 & ~x727 & ~x731 & ~x749 & ~x752 & ~x754 & ~x756 & ~x758 & ~x763 & ~x771 & ~x774;
assign c2136 =  x224;
assign c2138 = ~x0 & ~x5 & ~x12 & ~x36 & ~x44 & ~x50 & ~x57 & ~x69 & ~x75 & ~x77 & ~x80 & ~x81 & ~x90 & ~x100 & ~x101 & ~x102 & ~x103 & ~x106 & ~x107 & ~x108 & ~x116 & ~x136 & ~x157 & ~x158 & ~x162 & ~x163 & ~x190 & ~x191 & ~x194 & ~x196 & ~x199 & ~x200 & ~x214 & ~x215 & ~x224 & ~x244 & ~x248 & ~x251 & ~x272 & ~x273 & ~x276 & ~x281 & ~x299 & ~x306 & ~x310 & ~x329 & ~x330 & ~x331 & ~x337 & ~x358 & ~x363 & ~x365 & ~x383 & ~x394 & ~x412 & ~x413 & ~x420 & ~x424 & ~x452 & ~x503 & ~x560 & ~x561 & ~x564 & ~x565 & ~x603 & ~x612 & ~x615 & ~x631 & ~x632 & ~x633 & ~x646 & ~x648 & ~x656 & ~x657 & ~x658 & ~x659 & ~x660 & ~x661 & ~x669 & ~x671 & ~x674 & ~x677 & ~x678 & ~x681 & ~x683 & ~x686 & ~x688 & ~x689 & ~x691 & ~x704 & ~x705 & ~x706 & ~x717 & ~x721 & ~x722 & ~x725 & ~x726 & ~x729 & ~x735 & ~x736 & ~x737 & ~x741 & ~x748 & ~x755 & ~x759 & ~x761 & ~x763 & ~x765 & ~x775 & ~x776;
assign c2140 =  x590;
assign c2142 =  x501;
assign c2144 =  x639;
assign c2146 =  x461 &  x488 & ~x0 & ~x1 & ~x3 & ~x5 & ~x8 & ~x9 & ~x13 & ~x14 & ~x16 & ~x17 & ~x20 & ~x24 & ~x30 & ~x33 & ~x35 & ~x39 & ~x42 & ~x49 & ~x50 & ~x57 & ~x58 & ~x62 & ~x65 & ~x66 & ~x74 & ~x75 & ~x78 & ~x84 & ~x85 & ~x87 & ~x89 & ~x91 & ~x93 & ~x97 & ~x105 & ~x113 & ~x133 & ~x135 & ~x136 & ~x144 & ~x145 & ~x148 & ~x149 & ~x150 & ~x151 & ~x164 & ~x170 & ~x171 & ~x173 & ~x174 & ~x177 & ~x191 & ~x201 & ~x203 & ~x205 & ~x219 & ~x229 & ~x230 & ~x233 & ~x253 & ~x256 & ~x279 & ~x309 & ~x338 & ~x362 & ~x363 & ~x365 & ~x366 & ~x367 & ~x392 & ~x393 & ~x395 & ~x419 & ~x421 & ~x424 & ~x530 & ~x560 & ~x599 & ~x600 & ~x604 & ~x605 & ~x613 & ~x618 & ~x626 & ~x627 & ~x629 & ~x632 & ~x633 & ~x635 & ~x636 & ~x642 & ~x645 & ~x647 & ~x648 & ~x652 & ~x653 & ~x655 & ~x657 & ~x659 & ~x660 & ~x662 & ~x667 & ~x681 & ~x682 & ~x683 & ~x688 & ~x690 & ~x691 & ~x697 & ~x704 & ~x706 & ~x708 & ~x713 & ~x714 & ~x715 & ~x717 & ~x719 & ~x727 & ~x730 & ~x734 & ~x740 & ~x743 & ~x750 & ~x754 & ~x756 & ~x757 & ~x761 & ~x762 & ~x763 & ~x764 & ~x766 & ~x774 & ~x776 & ~x777 & ~x779 & ~x782;
assign c2148 =  x171;
assign c2150 =  x181 &  x543 & ~x8 & ~x195 & ~x285 & ~x313 & ~x315 & ~x319 & ~x321 & ~x343 & ~x349 & ~x440 & ~x441 & ~x502 & ~x585 & ~x645 & ~x711;
assign c2152 = ~x0 & ~x2 & ~x7 & ~x12 & ~x15 & ~x19 & ~x24 & ~x27 & ~x28 & ~x34 & ~x38 & ~x40 & ~x42 & ~x43 & ~x44 & ~x46 & ~x49 & ~x63 & ~x66 & ~x79 & ~x80 & ~x94 & ~x96 & ~x107 & ~x108 & ~x114 & ~x115 & ~x118 & ~x137 & ~x139 & ~x168 & ~x194 & ~x195 & ~x222 & ~x248 & ~x266 & ~x277 & ~x278 & ~x279 & ~x281 & ~x292 & ~x294 & ~x306 & ~x318 & ~x319 & ~x321 & ~x322 & ~x324 & ~x336 & ~x337 & ~x343 & ~x344 & ~x352 & ~x359 & ~x363 & ~x365 & ~x366 & ~x369 & ~x370 & ~x387 & ~x392 & ~x395 & ~x415 & ~x417 & ~x420 & ~x445 & ~x448 & ~x449 & ~x474 & ~x502 & ~x507 & ~x530 & ~x533 & ~x534 & ~x535 & ~x558 & ~x562 & ~x585 & ~x587 & ~x615 & ~x616 & ~x642 & ~x643 & ~x669 & ~x671 & ~x672 & ~x678 & ~x698 & ~x702 & ~x704 & ~x708 & ~x729 & ~x737 & ~x747 & ~x748 & ~x753 & ~x769 & ~x772 & ~x773 & ~x775 & ~x776 & ~x777 & ~x779;
assign c2154 =  x418;
assign c2156 =  x581 &  x582 & ~x1 & ~x10 & ~x22 & ~x65 & ~x79 & ~x88 & ~x133 & ~x199 & ~x253 & ~x255 & ~x282 & ~x311 & ~x337 & ~x360 & ~x386 & ~x415 & ~x448 & ~x530 & ~x643 & ~x663 & ~x672 & ~x690 & ~x708 & ~x726 & ~x738 & ~x748 & ~x757 & ~x779 & ~x781;
assign c2158 =  x756;
assign c2160 =  x239 &  x488 &  x489 &  x542 & ~x19 & ~x129 & ~x146 & ~x164 & ~x194 & ~x200 & ~x230 & ~x260 & ~x286 & ~x413 & ~x414 & ~x441 & ~x468 & ~x717 & ~x763 & ~x772;
assign c2162 =  x519 &  x548 &  x549 &  x583;
assign c2164 = ~x7 & ~x10 & ~x15 & ~x38 & ~x42 & ~x56 & ~x75 & ~x76 & ~x85 & ~x101 & ~x103 & ~x117 & ~x127 & ~x129 & ~x136 & ~x141 & ~x162 & ~x185 & ~x186 & ~x187 & ~x188 & ~x220 & ~x246 & ~x247 & ~x249 & ~x270 & ~x298 & ~x327 & ~x339 & ~x354 & ~x382 & ~x396 & ~x452 & ~x503 & ~x537 & ~x560 & ~x603 & ~x615 & ~x620 & ~x630 & ~x632 & ~x633 & ~x635 & ~x637 & ~x646 & ~x658 & ~x659 & ~x660 & ~x663 & ~x670 & ~x673 & ~x684 & ~x685 & ~x687 & ~x688 & ~x699 & ~x700 & ~x705 & ~x714 & ~x751 & ~x766 & ~x776;
assign c2166 =  x696;
assign c2168 =  x21;
assign c2170 =  x212 &  x571 &  x606 & ~x0 & ~x2 & ~x14 & ~x17 & ~x27 & ~x28 & ~x32 & ~x34 & ~x36 & ~x49 & ~x103 & ~x141 & ~x171 & ~x221 & ~x279 & ~x304 & ~x311 & ~x360 & ~x386 & ~x387 & ~x388 & ~x426 & ~x441 & ~x442 & ~x443 & ~x449 & ~x468 & ~x469 & ~x470 & ~x471 & ~x474 & ~x494 & ~x495 & ~x496 & ~x507 & ~x535 & ~x558 & ~x559 & ~x616 & ~x669 & ~x688 & ~x703 & ~x710 & ~x727 & ~x737 & ~x739 & ~x755 & ~x756 & ~x764;
assign c2174 =  x156 &  x297 &  x486 & ~x466;
assign c2176 = ~x6 & ~x10 & ~x16 & ~x17 & ~x22 & ~x25 & ~x26 & ~x28 & ~x35 & ~x36 & ~x37 & ~x42 & ~x43 & ~x46 & ~x47 & ~x48 & ~x49 & ~x52 & ~x53 & ~x55 & ~x56 & ~x58 & ~x60 & ~x61 & ~x62 & ~x64 & ~x65 & ~x70 & ~x73 & ~x74 & ~x77 & ~x81 & ~x82 & ~x84 & ~x86 & ~x88 & ~x92 & ~x93 & ~x95 & ~x99 & ~x100 & ~x102 & ~x105 & ~x107 & ~x109 & ~x110 & ~x111 & ~x113 & ~x114 & ~x115 & ~x117 & ~x120 & ~x121 & ~x123 & ~x134 & ~x135 & ~x136 & ~x141 & ~x144 & ~x145 & ~x164 & ~x169 & ~x171 & ~x172 & ~x192 & ~x193 & ~x196 & ~x197 & ~x199 & ~x200 & ~x220 & ~x227 & ~x248 & ~x250 & ~x252 & ~x253 & ~x255 & ~x256 & ~x276 & ~x279 & ~x280 & ~x283 & ~x284 & ~x305 & ~x307 & ~x308 & ~x310 & ~x311 & ~x332 & ~x334 & ~x335 & ~x336 & ~x338 & ~x339 & ~x351 & ~x359 & ~x361 & ~x362 & ~x363 & ~x364 & ~x366 & ~x367 & ~x368 & ~x373 & ~x374 & ~x376 & ~x377 & ~x378 & ~x379 & ~x391 & ~x393 & ~x394 & ~x396 & ~x398 & ~x399 & ~x414 & ~x415 & ~x419 & ~x420 & ~x421 & ~x423 & ~x424 & ~x425 & ~x426 & ~x442 & ~x443 & ~x447 & ~x449 & ~x451 & ~x452 & ~x473 & ~x477 & ~x480 & ~x506 & ~x508 & ~x534 & ~x536 & ~x559 & ~x561 & ~x585 & ~x586 & ~x590 & ~x591 & ~x612 & ~x619 & ~x643 & ~x644 & ~x645 & ~x669 & ~x673 & ~x675 & ~x676 & ~x677 & ~x692 & ~x696 & ~x698 & ~x700 & ~x701 & ~x704 & ~x706 & ~x708 & ~x709 & ~x710 & ~x711 & ~x712 & ~x718 & ~x721 & ~x725 & ~x728 & ~x729 & ~x730 & ~x731 & ~x732 & ~x734 & ~x736 & ~x737 & ~x738 & ~x740 & ~x742 & ~x743 & ~x744 & ~x746 & ~x747 & ~x749 & ~x750 & ~x751 & ~x753 & ~x757 & ~x759 & ~x763 & ~x765 & ~x766 & ~x769 & ~x771 & ~x773 & ~x777 & ~x778 & ~x783;
assign c2178 =  x778;
assign c2180 =  x460 &  x569 & ~x313 & ~x342 & ~x400 & ~x480 & ~x701 & ~x769;
assign c2182 =  x608 & ~x7 & ~x9 & ~x10 & ~x13 & ~x19 & ~x29 & ~x30 & ~x33 & ~x68 & ~x77 & ~x87 & ~x91 & ~x116 & ~x141 & ~x142 & ~x166 & ~x221 & ~x254 & ~x280 & ~x281 & ~x285 & ~x305 & ~x306 & ~x310 & ~x335 & ~x339 & ~x362 & ~x363 & ~x390 & ~x392 & ~x393 & ~x397 & ~x417 & ~x446 & ~x496 & ~x498 & ~x499 & ~x529 & ~x587 & ~x589 & ~x617 & ~x644 & ~x647 & ~x662 & ~x669 & ~x673 & ~x674 & ~x679 & ~x690 & ~x694 & ~x697 & ~x712 & ~x718 & ~x731 & ~x739 & ~x744 & ~x748 & ~x754 & ~x759 & ~x765 & ~x768 & ~x770 & ~x779;
assign c2184 =  x153 & ~x2 & ~x3 & ~x4 & ~x5 & ~x8 & ~x10 & ~x12 & ~x14 & ~x23 & ~x27 & ~x31 & ~x33 & ~x36 & ~x37 & ~x41 & ~x46 & ~x47 & ~x48 & ~x50 & ~x51 & ~x55 & ~x63 & ~x70 & ~x72 & ~x74 & ~x75 & ~x76 & ~x79 & ~x87 & ~x89 & ~x91 & ~x92 & ~x105 & ~x106 & ~x111 & ~x115 & ~x118 & ~x132 & ~x135 & ~x136 & ~x138 & ~x139 & ~x141 & ~x142 & ~x144 & ~x145 & ~x168 & ~x169 & ~x192 & ~x195 & ~x196 & ~x197 & ~x219 & ~x221 & ~x227 & ~x253 & ~x279 & ~x283 & ~x294 & ~x304 & ~x305 & ~x307 & ~x309 & ~x311 & ~x322 & ~x331 & ~x334 & ~x348 & ~x359 & ~x366 & ~x367 & ~x369 & ~x375 & ~x376 & ~x387 & ~x388 & ~x394 & ~x397 & ~x398 & ~x399 & ~x402 & ~x415 & ~x416 & ~x419 & ~x420 & ~x424 & ~x425 & ~x428 & ~x443 & ~x445 & ~x446 & ~x450 & ~x455 & ~x456 & ~x472 & ~x478 & ~x480 & ~x500 & ~x503 & ~x504 & ~x508 & ~x533 & ~x534 & ~x556 & ~x558 & ~x563 & ~x565 & ~x566 & ~x585 & ~x590 & ~x591 & ~x593 & ~x616 & ~x620 & ~x621 & ~x645 & ~x647 & ~x671 & ~x676 & ~x677 & ~x679 & ~x700 & ~x702 & ~x704 & ~x708 & ~x710 & ~x712 & ~x713 & ~x714 & ~x718 & ~x724 & ~x728 & ~x733 & ~x735 & ~x737 & ~x740 & ~x743 & ~x744 & ~x746 & ~x749 & ~x751 & ~x754 & ~x760 & ~x763 & ~x766 & ~x769 & ~x771 & ~x777 & ~x780 & ~x782 & ~x783;
assign c2186 =  x156 &  x184 &  x463 & ~x2 & ~x8 & ~x10 & ~x35 & ~x36 & ~x38 & ~x52 & ~x72 & ~x77 & ~x100 & ~x102 & ~x109 & ~x112 & ~x113 & ~x117 & ~x166 & ~x192 & ~x196 & ~x199 & ~x221 & ~x228 & ~x250 & ~x257 & ~x259 & ~x332 & ~x350 & ~x394 & ~x451 & ~x475 & ~x532 & ~x585 & ~x637 & ~x643 & ~x647 & ~x669 & ~x674 & ~x686 & ~x689 & ~x690 & ~x694 & ~x701 & ~x704 & ~x706 & ~x707 & ~x712 & ~x719 & ~x735 & ~x738 & ~x746 & ~x753 & ~x765 & ~x767 & ~x772;
assign c2188 =  x182 &  x628 & ~x8 & ~x14 & ~x15 & ~x17 & ~x18 & ~x23 & ~x25 & ~x30 & ~x31 & ~x34 & ~x44 & ~x52 & ~x53 & ~x57 & ~x59 & ~x66 & ~x68 & ~x69 & ~x80 & ~x82 & ~x87 & ~x95 & ~x100 & ~x102 & ~x109 & ~x113 & ~x121 & ~x123 & ~x132 & ~x133 & ~x135 & ~x137 & ~x143 & ~x167 & ~x198 & ~x220 & ~x254 & ~x282 & ~x306 & ~x307 & ~x334 & ~x336 & ~x351 & ~x362 & ~x378 & ~x379 & ~x389 & ~x391 & ~x396 & ~x402 & ~x403 & ~x404 & ~x406 & ~x415 & ~x424 & ~x428 & ~x430 & ~x442 & ~x443 & ~x447 & ~x454 & ~x479 & ~x480 & ~x503 & ~x504 & ~x506 & ~x507 & ~x508 & ~x510 & ~x533 & ~x613 & ~x615 & ~x646 & ~x698 & ~x707 & ~x708 & ~x710 & ~x711 & ~x712 & ~x724 & ~x726 & ~x736 & ~x742 & ~x753 & ~x758 & ~x768 & ~x769 & ~x771 & ~x780;
assign c2190 =  x570 &  x605 & ~x39 & ~x42 & ~x74 & ~x86 & ~x103 & ~x106 & ~x277 & ~x308 & ~x395 & ~x439 & ~x441 & ~x442 & ~x449 & ~x467 & ~x468 & ~x472 & ~x494 & ~x496 & ~x508 & ~x556 & ~x557 & ~x562 & ~x563 & ~x613 & ~x641 & ~x645 & ~x686 & ~x731 & ~x779;
assign c2192 =  x153 & ~x2 & ~x10 & ~x20 & ~x25 & ~x103 & ~x104 & ~x134 & ~x144 & ~x196 & ~x217 & ~x273 & ~x274 & ~x281 & ~x301 & ~x321 & ~x334 & ~x341 & ~x366 & ~x391 & ~x420 & ~x450 & ~x471 & ~x496 & ~x551 & ~x586 & ~x589 & ~x590 & ~x593 & ~x623 & ~x669 & ~x711 & ~x712 & ~x737 & ~x782;
assign c2194 =  x754;
assign c2196 =  x703;
assign c2198 =  x184 & ~x64 & ~x68 & ~x70 & ~x73 & ~x74 & ~x92 & ~x97 & ~x101 & ~x176 & ~x222 & ~x247 & ~x274 & ~x307 & ~x330 & ~x348 & ~x350 & ~x385 & ~x418 & ~x422 & ~x468 & ~x494 & ~x528 & ~x535 & ~x536 & ~x620 & ~x642 & ~x695 & ~x696 & ~x701 & ~x714 & ~x721 & ~x729 & ~x766 & ~x773;
assign c2200 =  x182 & ~x16 & ~x25 & ~x34 & ~x41 & ~x46 & ~x71 & ~x78 & ~x90 & ~x103 & ~x113 & ~x114 & ~x173 & ~x192 & ~x221 & ~x294 & ~x305 & ~x311 & ~x322 & ~x331 & ~x346 & ~x349 & ~x363 & ~x366 & ~x368 & ~x387 & ~x393 & ~x399 & ~x444 & ~x452 & ~x483 & ~x501 & ~x551 & ~x616 & ~x621 & ~x648 & ~x673 & ~x701 & ~x712 & ~x713 & ~x747 & ~x749 & ~x757 & ~x759 & ~x783;
assign c2202 =  x458 &  x512 & ~x2 & ~x3 & ~x4 & ~x9 & ~x14 & ~x15 & ~x16 & ~x17 & ~x19 & ~x20 & ~x21 & ~x22 & ~x29 & ~x30 & ~x34 & ~x36 & ~x39 & ~x40 & ~x49 & ~x54 & ~x55 & ~x63 & ~x77 & ~x78 & ~x80 & ~x82 & ~x88 & ~x90 & ~x91 & ~x107 & ~x108 & ~x109 & ~x112 & ~x114 & ~x117 & ~x118 & ~x119 & ~x139 & ~x144 & ~x168 & ~x170 & ~x171 & ~x193 & ~x197 & ~x199 & ~x223 & ~x226 & ~x227 & ~x249 & ~x305 & ~x320 & ~x336 & ~x338 & ~x344 & ~x347 & ~x362 & ~x367 & ~x369 & ~x371 & ~x396 & ~x421 & ~x445 & ~x450 & ~x475 & ~x476 & ~x477 & ~x506 & ~x558 & ~x561 & ~x588 & ~x589 & ~x619 & ~x637 & ~x643 & ~x662 & ~x663 & ~x665 & ~x670 & ~x676 & ~x677 & ~x683 & ~x684 & ~x685 & ~x698 & ~x704 & ~x705 & ~x707 & ~x708 & ~x710 & ~x713 & ~x716 & ~x719 & ~x722 & ~x723 & ~x726 & ~x728 & ~x729 & ~x730 & ~x731 & ~x733 & ~x735 & ~x740 & ~x742 & ~x749 & ~x750 & ~x752 & ~x756 & ~x758 & ~x759 & ~x760 & ~x763 & ~x776 & ~x779;
assign c2204 =  x250;
assign c2206 =  x465 &  x547 &  x599 & ~x3 & ~x4 & ~x5 & ~x10 & ~x11 & ~x14 & ~x19 & ~x24 & ~x30 & ~x31 & ~x34 & ~x38 & ~x39 & ~x40 & ~x44 & ~x47 & ~x49 & ~x51 & ~x56 & ~x59 & ~x70 & ~x73 & ~x75 & ~x77 & ~x79 & ~x82 & ~x85 & ~x89 & ~x90 & ~x107 & ~x110 & ~x112 & ~x114 & ~x115 & ~x119 & ~x134 & ~x139 & ~x140 & ~x142 & ~x143 & ~x163 & ~x170 & ~x173 & ~x192 & ~x193 & ~x196 & ~x198 & ~x199 & ~x201 & ~x220 & ~x221 & ~x225 & ~x227 & ~x248 & ~x251 & ~x252 & ~x255 & ~x257 & ~x258 & ~x276 & ~x280 & ~x282 & ~x283 & ~x284 & ~x295 & ~x304 & ~x308 & ~x311 & ~x312 & ~x323 & ~x336 & ~x337 & ~x338 & ~x340 & ~x341 & ~x361 & ~x363 & ~x365 & ~x366 & ~x369 & ~x389 & ~x392 & ~x395 & ~x396 & ~x417 & ~x419 & ~x421 & ~x446 & ~x451 & ~x472 & ~x473 & ~x474 & ~x476 & ~x477 & ~x502 & ~x507 & ~x531 & ~x533 & ~x535 & ~x560 & ~x584 & ~x588 & ~x590 & ~x591 & ~x618 & ~x640 & ~x641 & ~x644 & ~x645 & ~x657 & ~x658 & ~x667 & ~x668 & ~x671 & ~x674 & ~x685 & ~x686 & ~x687 & ~x698 & ~x703 & ~x704 & ~x706 & ~x708 & ~x709 & ~x712 & ~x714 & ~x716 & ~x722 & ~x723 & ~x734 & ~x736 & ~x739 & ~x740 & ~x742 & ~x743 & ~x746 & ~x748 & ~x750 & ~x756 & ~x761 & ~x763 & ~x765 & ~x770 & ~x771 & ~x775 & ~x777 & ~x779;
assign c2208 =  x375 & ~x192 & ~x202 & ~x232 & ~x234 & ~x259 & ~x262 & ~x263 & ~x265 & ~x287 & ~x288 & ~x290 & ~x292 & ~x293 & ~x294 & ~x295 & ~x658 & ~x686;
assign c2210 =  x527 & ~x331 & ~x398 & ~x632 & ~x660;
assign c2212 =  x432 &  x461 & ~x8 & ~x9 & ~x10 & ~x11 & ~x12 & ~x15 & ~x16 & ~x20 & ~x21 & ~x23 & ~x24 & ~x26 & ~x27 & ~x29 & ~x30 & ~x33 & ~x41 & ~x45 & ~x46 & ~x49 & ~x50 & ~x52 & ~x53 & ~x55 & ~x60 & ~x64 & ~x80 & ~x81 & ~x85 & ~x88 & ~x91 & ~x92 & ~x94 & ~x95 & ~x103 & ~x104 & ~x105 & ~x107 & ~x109 & ~x110 & ~x111 & ~x113 & ~x114 & ~x117 & ~x123 & ~x139 & ~x141 & ~x143 & ~x144 & ~x145 & ~x147 & ~x149 & ~x164 & ~x166 & ~x169 & ~x170 & ~x171 & ~x172 & ~x191 & ~x192 & ~x195 & ~x197 & ~x198 & ~x200 & ~x203 & ~x221 & ~x223 & ~x224 & ~x248 & ~x250 & ~x254 & ~x276 & ~x277 & ~x278 & ~x281 & ~x283 & ~x284 & ~x304 & ~x308 & ~x309 & ~x332 & ~x333 & ~x335 & ~x336 & ~x341 & ~x362 & ~x364 & ~x365 & ~x367 & ~x391 & ~x418 & ~x419 & ~x421 & ~x448 & ~x449 & ~x476 & ~x477 & ~x504 & ~x530 & ~x532 & ~x534 & ~x560 & ~x562 & ~x589 & ~x590 & ~x601 & ~x613 & ~x615 & ~x617 & ~x628 & ~x629 & ~x631 & ~x643 & ~x647 & ~x652 & ~x653 & ~x654 & ~x658 & ~x659 & ~x666 & ~x668 & ~x670 & ~x673 & ~x675 & ~x676 & ~x677 & ~x678 & ~x679 & ~x680 & ~x681 & ~x682 & ~x683 & ~x685 & ~x686 & ~x690 & ~x692 & ~x694 & ~x695 & ~x697 & ~x700 & ~x702 & ~x707 & ~x709 & ~x710 & ~x715 & ~x716 & ~x717 & ~x719 & ~x723 & ~x724 & ~x726 & ~x727 & ~x728 & ~x733 & ~x742 & ~x744 & ~x747 & ~x749 & ~x756 & ~x758 & ~x761 & ~x762 & ~x763 & ~x770 & ~x774 & ~x782 & ~x783;
assign c2214 =  x488 & ~x1 & ~x53 & ~x57 & ~x64 & ~x66 & ~x87 & ~x102 & ~x136 & ~x138 & ~x162 & ~x191 & ~x218 & ~x219 & ~x251 & ~x278 & ~x311 & ~x319 & ~x320 & ~x338 & ~x346 & ~x348 & ~x373 & ~x397 & ~x399 & ~x424 & ~x473 & ~x522 & ~x589 & ~x591 & ~x619 & ~x642 & ~x646 & ~x653 & ~x675 & ~x679 & ~x681 & ~x682 & ~x703 & ~x709 & ~x712 & ~x733 & ~x737 & ~x745 & ~x758 & ~x777;
assign c2216 =  x431 &  x497 &  x500;
assign c2218 = ~x3 & ~x11 & ~x16 & ~x17 & ~x19 & ~x20 & ~x27 & ~x28 & ~x40 & ~x45 & ~x47 & ~x49 & ~x51 & ~x56 & ~x61 & ~x62 & ~x64 & ~x71 & ~x75 & ~x80 & ~x84 & ~x85 & ~x86 & ~x106 & ~x111 & ~x117 & ~x118 & ~x131 & ~x137 & ~x140 & ~x141 & ~x162 & ~x167 & ~x175 & ~x176 & ~x187 & ~x196 & ~x198 & ~x215 & ~x217 & ~x222 & ~x246 & ~x254 & ~x255 & ~x276 & ~x279 & ~x281 & ~x283 & ~x309 & ~x335 & ~x338 & ~x356 & ~x364 & ~x373 & ~x392 & ~x395 & ~x396 & ~x398 & ~x419 & ~x422 & ~x423 & ~x476 & ~x477 & ~x478 & ~x503 & ~x531 & ~x536 & ~x560 & ~x576 & ~x587 & ~x589 & ~x593 & ~x603 & ~x633 & ~x642 & ~x647 & ~x648 & ~x654 & ~x658 & ~x660 & ~x662 & ~x664 & ~x665 & ~x672 & ~x673 & ~x676 & ~x679 & ~x683 & ~x686 & ~x687 & ~x690 & ~x708 & ~x714 & ~x716 & ~x720 & ~x728 & ~x731 & ~x732 & ~x745 & ~x747 & ~x749 & ~x752 & ~x753 & ~x764 & ~x767 & ~x768 & ~x770 & ~x772 & ~x774 & ~x777;
assign c2220 =  x186 &  x517 & ~x0 & ~x3 & ~x4 & ~x5 & ~x8 & ~x9 & ~x12 & ~x14 & ~x17 & ~x33 & ~x34 & ~x35 & ~x38 & ~x45 & ~x46 & ~x47 & ~x49 & ~x50 & ~x51 & ~x53 & ~x59 & ~x60 & ~x64 & ~x65 & ~x66 & ~x75 & ~x77 & ~x78 & ~x80 & ~x81 & ~x82 & ~x84 & ~x87 & ~x88 & ~x92 & ~x95 & ~x108 & ~x109 & ~x110 & ~x112 & ~x115 & ~x117 & ~x118 & ~x119 & ~x120 & ~x121 & ~x122 & ~x135 & ~x136 & ~x138 & ~x139 & ~x140 & ~x141 & ~x142 & ~x143 & ~x146 & ~x147 & ~x148 & ~x149 & ~x150 & ~x164 & ~x166 & ~x170 & ~x171 & ~x173 & ~x175 & ~x192 & ~x195 & ~x196 & ~x200 & ~x220 & ~x221 & ~x223 & ~x224 & ~x225 & ~x228 & ~x229 & ~x230 & ~x250 & ~x255 & ~x258 & ~x276 & ~x277 & ~x278 & ~x279 & ~x281 & ~x283 & ~x284 & ~x285 & ~x286 & ~x287 & ~x296 & ~x304 & ~x305 & ~x308 & ~x312 & ~x334 & ~x335 & ~x339 & ~x364 & ~x366 & ~x368 & ~x387 & ~x391 & ~x394 & ~x416 & ~x417 & ~x418 & ~x420 & ~x422 & ~x446 & ~x448 & ~x449 & ~x450 & ~x473 & ~x477 & ~x500 & ~x502 & ~x504 & ~x505 & ~x506 & ~x529 & ~x530 & ~x534 & ~x557 & ~x558 & ~x559 & ~x562 & ~x586 & ~x588 & ~x589 & ~x612 & ~x614 & ~x618 & ~x642 & ~x643 & ~x646 & ~x655 & ~x656 & ~x658 & ~x668 & ~x669 & ~x670 & ~x674 & ~x675 & ~x681 & ~x683 & ~x684 & ~x687 & ~x693 & ~x695 & ~x698 & ~x700 & ~x703 & ~x705 & ~x711 & ~x718 & ~x719 & ~x720 & ~x721 & ~x724 & ~x726 & ~x728 & ~x729 & ~x730 & ~x735 & ~x737 & ~x738 & ~x739 & ~x740 & ~x741 & ~x745 & ~x746 & ~x752 & ~x755 & ~x756 & ~x760 & ~x761 & ~x768 & ~x769 & ~x774 & ~x776 & ~x777 & ~x781;
assign c2222 =  x602 & ~x10 & ~x25 & ~x48 & ~x62 & ~x75 & ~x77 & ~x80 & ~x81 & ~x91 & ~x107 & ~x138 & ~x142 & ~x228 & ~x255 & ~x285 & ~x308 & ~x310 & ~x327 & ~x330 & ~x333 & ~x338 & ~x340 & ~x383 & ~x400 & ~x421 & ~x423 & ~x426 & ~x438 & ~x449 & ~x452 & ~x492 & ~x531 & ~x560 & ~x563 & ~x645 & ~x646 & ~x667 & ~x676 & ~x695 & ~x704 & ~x709 & ~x721 & ~x729 & ~x730 & ~x743 & ~x753;
assign c2224 =  x150 & ~x4 & ~x9 & ~x30 & ~x33 & ~x38 & ~x61 & ~x63 & ~x73 & ~x134 & ~x138 & ~x189 & ~x192 & ~x198 & ~x220 & ~x256 & ~x263 & ~x291 & ~x310 & ~x312 & ~x319 & ~x335 & ~x345 & ~x346 & ~x370 & ~x372 & ~x388 & ~x397 & ~x398 & ~x427 & ~x449 & ~x475 & ~x510 & ~x565 & ~x591 & ~x650 & ~x651 & ~x677 & ~x680 & ~x699 & ~x712 & ~x723 & ~x730 & ~x732 & ~x753 & ~x754 & ~x757 & ~x759 & ~x773 & ~x783;
assign c2226 =  x701;
assign c2228 =  x540 & ~x2 & ~x3 & ~x8 & ~x13 & ~x16 & ~x41 & ~x45 & ~x50 & ~x54 & ~x59 & ~x60 & ~x71 & ~x72 & ~x74 & ~x77 & ~x83 & ~x111 & ~x133 & ~x137 & ~x142 & ~x144 & ~x165 & ~x197 & ~x218 & ~x219 & ~x247 & ~x252 & ~x254 & ~x275 & ~x294 & ~x304 & ~x305 & ~x311 & ~x322 & ~x334 & ~x335 & ~x342 & ~x343 & ~x389 & ~x397 & ~x398 & ~x419 & ~x423 & ~x425 & ~x446 & ~x447 & ~x450 & ~x452 & ~x476 & ~x478 & ~x504 & ~x505 & ~x506 & ~x535 & ~x562 & ~x588 & ~x614 & ~x641 & ~x645 & ~x647 & ~x648 & ~x649 & ~x660 & ~x668 & ~x675 & ~x680 & ~x681 & ~x684 & ~x695 & ~x696 & ~x702 & ~x704 & ~x710 & ~x714 & ~x724 & ~x728 & ~x737 & ~x738 & ~x741 & ~x751 & ~x753 & ~x755 & ~x767;
assign c2230 = ~x0 & ~x1 & ~x2 & ~x4 & ~x5 & ~x10 & ~x12 & ~x13 & ~x15 & ~x16 & ~x17 & ~x19 & ~x20 & ~x24 & ~x25 & ~x30 & ~x31 & ~x35 & ~x38 & ~x40 & ~x41 & ~x42 & ~x43 & ~x45 & ~x46 & ~x49 & ~x52 & ~x54 & ~x61 & ~x65 & ~x69 & ~x73 & ~x74 & ~x75 & ~x76 & ~x77 & ~x78 & ~x83 & ~x85 & ~x87 & ~x89 & ~x94 & ~x95 & ~x96 & ~x98 & ~x109 & ~x114 & ~x117 & ~x120 & ~x123 & ~x130 & ~x131 & ~x133 & ~x142 & ~x146 & ~x147 & ~x160 & ~x161 & ~x163 & ~x165 & ~x166 & ~x167 & ~x168 & ~x170 & ~x171 & ~x173 & ~x176 & ~x192 & ~x194 & ~x196 & ~x225 & ~x227 & ~x252 & ~x253 & ~x276 & ~x279 & ~x280 & ~x281 & ~x282 & ~x304 & ~x306 & ~x309 & ~x310 & ~x311 & ~x334 & ~x336 & ~x362 & ~x365 & ~x367 & ~x368 & ~x369 & ~x371 & ~x372 & ~x393 & ~x395 & ~x417 & ~x419 & ~x477 & ~x479 & ~x502 & ~x503 & ~x507 & ~x533 & ~x534 & ~x557 & ~x558 & ~x561 & ~x585 & ~x587 & ~x589 & ~x591 & ~x605 & ~x608 & ~x609 & ~x613 & ~x614 & ~x616 & ~x617 & ~x629 & ~x630 & ~x631 & ~x633 & ~x642 & ~x645 & ~x648 & ~x650 & ~x651 & ~x652 & ~x653 & ~x654 & ~x655 & ~x656 & ~x665 & ~x666 & ~x668 & ~x669 & ~x671 & ~x673 & ~x674 & ~x675 & ~x676 & ~x677 & ~x680 & ~x681 & ~x682 & ~x683 & ~x684 & ~x685 & ~x688 & ~x689 & ~x692 & ~x696 & ~x699 & ~x701 & ~x702 & ~x703 & ~x706 & ~x707 & ~x708 & ~x712 & ~x713 & ~x714 & ~x718 & ~x720 & ~x722 & ~x727 & ~x734 & ~x735 & ~x737 & ~x739 & ~x742 & ~x743 & ~x744 & ~x745 & ~x747 & ~x748 & ~x749 & ~x751 & ~x755 & ~x756 & ~x761 & ~x768 & ~x769 & ~x770 & ~x773 & ~x776 & ~x778 & ~x779 & ~x780;
assign c2232 =  x438 &  x518 &  x544 &  x570 & ~x6 & ~x25 & ~x39 & ~x42 & ~x47 & ~x56 & ~x58 & ~x59 & ~x62 & ~x85 & ~x106 & ~x110 & ~x137 & ~x142 & ~x170 & ~x195 & ~x226 & ~x249 & ~x254 & ~x280 & ~x283 & ~x310 & ~x320 & ~x335 & ~x347 & ~x369 & ~x395 & ~x397 & ~x446 & ~x451 & ~x477 & ~x505 & ~x534 & ~x559 & ~x562 & ~x585 & ~x589 & ~x616 & ~x671 & ~x679 & ~x706 & ~x708 & ~x710 & ~x711 & ~x724 & ~x725 & ~x732 & ~x739 & ~x753 & ~x760 & ~x762 & ~x763 & ~x767 & ~x772 & ~x774;
assign c2234 =  x600 & ~x26 & ~x35 & ~x37 & ~x42 & ~x57 & ~x63 & ~x64 & ~x67 & ~x91 & ~x109 & ~x136 & ~x143 & ~x196 & ~x197 & ~x279 & ~x302 & ~x306 & ~x357 & ~x372 & ~x414 & ~x417 & ~x439 & ~x441 & ~x447 & ~x465 & ~x467 & ~x519 & ~x559 & ~x561 & ~x586 & ~x613 & ~x615 & ~x643 & ~x746 & ~x749 & ~x759 & ~x760 & ~x778 & ~x780;
assign c2236 =  x463 &  x490 &  x517 & ~x4 & ~x19 & ~x22 & ~x23 & ~x30 & ~x36 & ~x50 & ~x52 & ~x53 & ~x54 & ~x55 & ~x57 & ~x61 & ~x66 & ~x67 & ~x71 & ~x73 & ~x76 & ~x78 & ~x86 & ~x87 & ~x93 & ~x94 & ~x100 & ~x102 & ~x104 & ~x110 & ~x113 & ~x116 & ~x123 & ~x135 & ~x141 & ~x163 & ~x165 & ~x166 & ~x170 & ~x172 & ~x192 & ~x194 & ~x200 & ~x201 & ~x220 & ~x221 & ~x226 & ~x228 & ~x247 & ~x249 & ~x256 & ~x281 & ~x312 & ~x329 & ~x331 & ~x332 & ~x339 & ~x359 & ~x367 & ~x391 & ~x396 & ~x404 & ~x415 & ~x416 & ~x422 & ~x429 & ~x430 & ~x439 & ~x440 & ~x441 & ~x451 & ~x473 & ~x478 & ~x481 & ~x505 & ~x506 & ~x591 & ~x641 & ~x672 & ~x705 & ~x708 & ~x709 & ~x710 & ~x715 & ~x717 & ~x719 & ~x722 & ~x732 & ~x734 & ~x735 & ~x736 & ~x742 & ~x743 & ~x746 & ~x747 & ~x750 & ~x758 & ~x768 & ~x770 & ~x771 & ~x779 & ~x780 & ~x782;
assign c2238 =  x458 &  x541 & ~x2 & ~x33 & ~x35 & ~x43 & ~x71 & ~x76 & ~x78 & ~x107 & ~x132 & ~x135 & ~x163 & ~x219 & ~x228 & ~x276 & ~x279 & ~x280 & ~x281 & ~x285 & ~x289 & ~x293 & ~x363 & ~x365 & ~x504 & ~x648 & ~x684 & ~x700 & ~x708 & ~x712 & ~x763 & ~x771 & ~x782;
assign c2240 =  x647;
assign c2242 =  x600 & ~x0 & ~x4 & ~x9 & ~x11 & ~x13 & ~x16 & ~x29 & ~x31 & ~x38 & ~x39 & ~x40 & ~x44 & ~x45 & ~x46 & ~x47 & ~x48 & ~x51 & ~x53 & ~x56 & ~x58 & ~x60 & ~x61 & ~x76 & ~x78 & ~x80 & ~x82 & ~x83 & ~x89 & ~x105 & ~x109 & ~x112 & ~x113 & ~x114 & ~x139 & ~x162 & ~x164 & ~x170 & ~x190 & ~x191 & ~x192 & ~x198 & ~x219 & ~x220 & ~x221 & ~x225 & ~x249 & ~x279 & ~x282 & ~x283 & ~x292 & ~x294 & ~x306 & ~x307 & ~x308 & ~x315 & ~x318 & ~x319 & ~x322 & ~x332 & ~x338 & ~x363 & ~x368 & ~x389 & ~x395 & ~x420 & ~x442 & ~x444 & ~x446 & ~x450 & ~x451 & ~x501 & ~x503 & ~x505 & ~x507 & ~x527 & ~x528 & ~x530 & ~x563 & ~x586 & ~x588 & ~x592 & ~x615 & ~x619 & ~x641 & ~x643 & ~x667 & ~x669 & ~x675 & ~x683 & ~x695 & ~x699 & ~x701 & ~x702 & ~x704 & ~x708 & ~x709 & ~x711 & ~x712 & ~x726 & ~x727 & ~x729 & ~x742 & ~x743 & ~x749 & ~x751 & ~x752 & ~x754 & ~x763 & ~x764 & ~x772 & ~x774 & ~x776 & ~x777 & ~x778 & ~x782;
assign c2244 =  x516 &  x570 &  x665 & ~x524;
assign c2246 = ~x295 & ~x297 & ~x316 & ~x318 & ~x322 & ~x325 & ~x344 & ~x345 & ~x347 & ~x348 & ~x349 & ~x350 & ~x352 & ~x353 & ~x380 & ~x397 & ~x398 & ~x425 & ~x697 & ~x705 & ~x763;
assign c2248 =  x182 & ~x3 & ~x24 & ~x25 & ~x29 & ~x32 & ~x37 & ~x44 & ~x54 & ~x78 & ~x84 & ~x96 & ~x100 & ~x103 & ~x104 & ~x139 & ~x141 & ~x144 & ~x167 & ~x220 & ~x224 & ~x225 & ~x226 & ~x228 & ~x294 & ~x307 & ~x334 & ~x348 & ~x359 & ~x360 & ~x369 & ~x374 & ~x376 & ~x392 & ~x393 & ~x421 & ~x424 & ~x429 & ~x465 & ~x478 & ~x479 & ~x501 & ~x506 & ~x533 & ~x536 & ~x557 & ~x585 & ~x586 & ~x641 & ~x643 & ~x647 & ~x666 & ~x671 & ~x674 & ~x678 & ~x679 & ~x695 & ~x710 & ~x733 & ~x737 & ~x751 & ~x760;
assign c2250 =  x592;
assign c2254 =  x583 & ~x74 & ~x372 & ~x500 & ~x662;
assign c2256 =  x456 & ~x28 & ~x41 & ~x48 & ~x54 & ~x59 & ~x62 & ~x68 & ~x70 & ~x78 & ~x86 & ~x87 & ~x109 & ~x111 & ~x135 & ~x143 & ~x165 & ~x167 & ~x168 & ~x199 & ~x222 & ~x248 & ~x265 & ~x276 & ~x286 & ~x311 & ~x313 & ~x317 & ~x320 & ~x322 & ~x342 & ~x362 & ~x367 & ~x368 & ~x392 & ~x418 & ~x451 & ~x532 & ~x589 & ~x617 & ~x620 & ~x646 & ~x659 & ~x668 & ~x669 & ~x684 & ~x687 & ~x692 & ~x699 & ~x706 & ~x708 & ~x714 & ~x745 & ~x746 & ~x749 & ~x764 & ~x776;
assign c2258 =  x475;
assign c2260 =  x432 &  x454 &  x509 & ~x287 & ~x316 & ~x340 & ~x664 & ~x691;
assign c2262 =  x175 & ~x290 & ~x346 & ~x348 & ~x362 & ~x371 & ~x373 & ~x417 & ~x592 & ~x678 & ~x764;
assign c2264 =  x702;
assign c2266 =  x295 &  x515 & ~x4 & ~x23 & ~x46 & ~x65 & ~x72 & ~x73 & ~x86 & ~x105 & ~x130 & ~x133 & ~x134 & ~x158 & ~x162 & ~x163 & ~x195 & ~x216 & ~x218 & ~x245 & ~x248 & ~x256 & ~x309 & ~x339 & ~x505 & ~x531 & ~x534 & ~x558 & ~x563 & ~x642 & ~x645 & ~x652 & ~x658 & ~x659 & ~x660 & ~x663 & ~x671 & ~x686 & ~x688 & ~x689 & ~x693 & ~x712 & ~x717 & ~x748 & ~x752 & ~x754 & ~x761 & ~x763 & ~x765 & ~x767 & ~x773 & ~x777;
assign c2268 = ~x2 & ~x5 & ~x6 & ~x10 & ~x14 & ~x17 & ~x18 & ~x21 & ~x23 & ~x25 & ~x26 & ~x28 & ~x33 & ~x34 & ~x37 & ~x38 & ~x42 & ~x44 & ~x45 & ~x46 & ~x47 & ~x49 & ~x50 & ~x51 & ~x55 & ~x56 & ~x58 & ~x60 & ~x63 & ~x64 & ~x67 & ~x69 & ~x72 & ~x73 & ~x75 & ~x77 & ~x78 & ~x79 & ~x80 & ~x82 & ~x84 & ~x85 & ~x86 & ~x87 & ~x89 & ~x90 & ~x92 & ~x93 & ~x95 & ~x106 & ~x107 & ~x110 & ~x115 & ~x119 & ~x122 & ~x124 & ~x135 & ~x136 & ~x138 & ~x142 & ~x143 & ~x144 & ~x146 & ~x147 & ~x149 & ~x161 & ~x163 & ~x165 & ~x167 & ~x168 & ~x175 & ~x190 & ~x191 & ~x192 & ~x194 & ~x201 & ~x202 & ~x219 & ~x220 & ~x221 & ~x222 & ~x224 & ~x225 & ~x226 & ~x227 & ~x229 & ~x230 & ~x250 & ~x251 & ~x252 & ~x254 & ~x275 & ~x276 & ~x277 & ~x279 & ~x282 & ~x304 & ~x306 & ~x308 & ~x310 & ~x311 & ~x312 & ~x336 & ~x337 & ~x338 & ~x339 & ~x340 & ~x342 & ~x393 & ~x394 & ~x395 & ~x420 & ~x421 & ~x448 & ~x449 & ~x477 & ~x478 & ~x505 & ~x506 & ~x531 & ~x534 & ~x557 & ~x558 & ~x560 & ~x561 & ~x575 & ~x590 & ~x591 & ~x602 & ~x603 & ~x605 & ~x611 & ~x613 & ~x614 & ~x616 & ~x617 & ~x618 & ~x619 & ~x626 & ~x627 & ~x629 & ~x632 & ~x633 & ~x641 & ~x647 & ~x650 & ~x651 & ~x652 & ~x659 & ~x660 & ~x663 & ~x666 & ~x669 & ~x671 & ~x672 & ~x673 & ~x676 & ~x678 & ~x679 & ~x680 & ~x682 & ~x684 & ~x688 & ~x689 & ~x696 & ~x700 & ~x703 & ~x704 & ~x705 & ~x710 & ~x711 & ~x712 & ~x713 & ~x714 & ~x715 & ~x716 & ~x717 & ~x718 & ~x721 & ~x722 & ~x723 & ~x724 & ~x726 & ~x728 & ~x734 & ~x735 & ~x737 & ~x739 & ~x740 & ~x748 & ~x749 & ~x751 & ~x753 & ~x755 & ~x756 & ~x757 & ~x758 & ~x759 & ~x763 & ~x766 & ~x769 & ~x770 & ~x771 & ~x772 & ~x773 & ~x778 & ~x781 & ~x782;
assign c2270 =  x449;
assign c2272 =  x446;
assign c2274 =  x553 & ~x26 & ~x40 & ~x415 & ~x424 & ~x441 & ~x443 & ~x448 & ~x449 & ~x451 & ~x562 & ~x608 & ~x633 & ~x638 & ~x659 & ~x686;
assign c2276 =  x782;
assign c2278 = ~x1 & ~x10 & ~x14 & ~x24 & ~x36 & ~x46 & ~x78 & ~x104 & ~x107 & ~x115 & ~x134 & ~x136 & ~x137 & ~x142 & ~x144 & ~x166 & ~x208 & ~x221 & ~x226 & ~x260 & ~x261 & ~x276 & ~x281 & ~x289 & ~x293 & ~x297 & ~x304 & ~x306 & ~x307 & ~x314 & ~x325 & ~x363 & ~x367 & ~x391 & ~x534 & ~x561 & ~x585 & ~x613 & ~x614 & ~x615 & ~x642 & ~x645 & ~x658 & ~x659 & ~x663 & ~x667 & ~x682 & ~x686 & ~x691 & ~x698 & ~x699 & ~x700 & ~x708 & ~x712 & ~x717 & ~x719 & ~x720 & ~x722 & ~x735 & ~x743 & ~x752 & ~x754 & ~x758 & ~x762 & ~x768 & ~x773 & ~x776;
assign c2280 =  x158 &  x159 &  x272 & ~x25 & ~x35 & ~x47 & ~x64 & ~x140 & ~x173 & ~x174 & ~x241 & ~x256 & ~x257 & ~x258 & ~x281 & ~x323 & ~x331 & ~x333 & ~x359 & ~x364 & ~x395 & ~x476 & ~x500 & ~x657 & ~x658 & ~x662 & ~x694 & ~x696 & ~x704 & ~x710 & ~x715 & ~x722 & ~x728 & ~x730;
assign c2282 =  x667;
assign c2284 =  x724;
assign c2286 =  x647;
assign c2288 =  x773;
assign c2290 =  x157 &  x516 & ~x55 & ~x267 & ~x276 & ~x280 & ~x320 & ~x335 & ~x347 & ~x364 & ~x402 & ~x414 & ~x474 & ~x532 & ~x562 & ~x705 & ~x725 & ~x731 & ~x777 & ~x782;
assign c2292 =  x517 & ~x6 & ~x8 & ~x21 & ~x40 & ~x45 & ~x46 & ~x50 & ~x51 & ~x53 & ~x61 & ~x76 & ~x81 & ~x87 & ~x97 & ~x104 & ~x105 & ~x110 & ~x112 & ~x115 & ~x130 & ~x142 & ~x143 & ~x159 & ~x192 & ~x193 & ~x196 & ~x199 & ~x249 & ~x277 & ~x278 & ~x301 & ~x305 & ~x336 & ~x338 & ~x343 & ~x363 & ~x364 & ~x367 & ~x375 & ~x395 & ~x400 & ~x419 & ~x429 & ~x448 & ~x451 & ~x453 & ~x476 & ~x506 & ~x508 & ~x532 & ~x537 & ~x538 & ~x562 & ~x586 & ~x588 & ~x590 & ~x591 & ~x595 & ~x620 & ~x642 & ~x645 & ~x646 & ~x648 & ~x685 & ~x688 & ~x698 & ~x699 & ~x703 & ~x705 & ~x707 & ~x711 & ~x716 & ~x717 & ~x723 & ~x724 & ~x729 & ~x742 & ~x743 & ~x761 & ~x763 & ~x772 & ~x773 & ~x781 & ~x783;
assign c2294 =  x418;
assign c2296 =  x553 & ~x10 & ~x15 & ~x18 & ~x24 & ~x36 & ~x45 & ~x60 & ~x73 & ~x84 & ~x102 & ~x110 & ~x116 & ~x134 & ~x192 & ~x196 & ~x197 & ~x220 & ~x221 & ~x253 & ~x254 & ~x280 & ~x309 & ~x310 & ~x331 & ~x359 & ~x360 & ~x362 & ~x385 & ~x393 & ~x395 & ~x443 & ~x448 & ~x502 & ~x589 & ~x614 & ~x634 & ~x659 & ~x660 & ~x663 & ~x675 & ~x686 & ~x688 & ~x689 & ~x694 & ~x695 & ~x699 & ~x702 & ~x705 & ~x707 & ~x719 & ~x722 & ~x724 & ~x733 & ~x736 & ~x739 & ~x745 & ~x747 & ~x754 & ~x764 & ~x765;
assign c2298 =  x92;
assign c21 =  x269 & ~x5 & ~x32 & ~x101 & ~x118 & ~x133 & ~x143 & ~x150 & ~x155 & ~x159 & ~x308 & ~x332 & ~x388 & ~x393 & ~x447 & ~x499 & ~x507 & ~x525 & ~x536 & ~x633 & ~x641 & ~x646 & ~x661 & ~x667 & ~x669 & ~x716 & ~x728 & ~x744 & ~x751;
assign c23 = ~x1 & ~x5 & ~x6 & ~x13 & ~x14 & ~x19 & ~x21 & ~x32 & ~x37 & ~x38 & ~x40 & ~x44 & ~x46 & ~x48 & ~x49 & ~x52 & ~x53 & ~x59 & ~x64 & ~x65 & ~x78 & ~x85 & ~x87 & ~x103 & ~x104 & ~x106 & ~x109 & ~x111 & ~x115 & ~x122 & ~x138 & ~x140 & ~x144 & ~x170 & ~x194 & ~x197 & ~x198 & ~x199 & ~x200 & ~x227 & ~x246 & ~x247 & ~x254 & ~x283 & ~x285 & ~x307 & ~x308 & ~x309 & ~x313 & ~x314 & ~x315 & ~x331 & ~x332 & ~x334 & ~x338 & ~x339 & ~x363 & ~x364 & ~x369 & ~x386 & ~x387 & ~x394 & ~x396 & ~x399 & ~x415 & ~x417 & ~x422 & ~x423 & ~x424 & ~x425 & ~x447 & ~x449 & ~x450 & ~x471 & ~x501 & ~x502 & ~x503 & ~x510 & ~x528 & ~x536 & ~x540 & ~x541 & ~x554 & ~x555 & ~x556 & ~x559 & ~x562 & ~x570 & ~x583 & ~x585 & ~x588 & ~x610 & ~x613 & ~x614 & ~x617 & ~x638 & ~x643 & ~x645 & ~x665 & ~x668 & ~x673 & ~x675 & ~x686 & ~x695 & ~x697 & ~x700 & ~x704 & ~x707 & ~x720 & ~x727 & ~x730 & ~x741 & ~x749 & ~x753 & ~x756 & ~x757 & ~x759 & ~x769 & ~x777;
assign c25 =  x343 &  x427 & ~x642;
assign c27 =  x573 & ~x1 & ~x3 & ~x5 & ~x7 & ~x15 & ~x17 & ~x18 & ~x23 & ~x26 & ~x29 & ~x30 & ~x33 & ~x36 & ~x39 & ~x40 & ~x42 & ~x43 & ~x54 & ~x62 & ~x63 & ~x83 & ~x84 & ~x86 & ~x87 & ~x89 & ~x94 & ~x105 & ~x111 & ~x115 & ~x139 & ~x141 & ~x142 & ~x144 & ~x146 & ~x147 & ~x148 & ~x165 & ~x166 & ~x167 & ~x168 & ~x169 & ~x170 & ~x174 & ~x192 & ~x194 & ~x196 & ~x199 & ~x200 & ~x220 & ~x221 & ~x222 & ~x224 & ~x229 & ~x230 & ~x250 & ~x252 & ~x253 & ~x257 & ~x271 & ~x272 & ~x274 & ~x283 & ~x284 & ~x296 & ~x297 & ~x307 & ~x311 & ~x312 & ~x336 & ~x337 & ~x363 & ~x364 & ~x366 & ~x368 & ~x391 & ~x393 & ~x395 & ~x420 & ~x421 & ~x423 & ~x424 & ~x446 & ~x447 & ~x477 & ~x479 & ~x480 & ~x502 & ~x506 & ~x507 & ~x560 & ~x563 & ~x565 & ~x588 & ~x593 & ~x617 & ~x620 & ~x623 & ~x638 & ~x639 & ~x643 & ~x648 & ~x649 & ~x652 & ~x664 & ~x665 & ~x666 & ~x667 & ~x671 & ~x672 & ~x673 & ~x674 & ~x680 & ~x682 & ~x685 & ~x693 & ~x694 & ~x696 & ~x697 & ~x700 & ~x703 & ~x705 & ~x708 & ~x709 & ~x711 & ~x713 & ~x715 & ~x716 & ~x720 & ~x722 & ~x726 & ~x727 & ~x737 & ~x738 & ~x739 & ~x740 & ~x741 & ~x746 & ~x750 & ~x752 & ~x755 & ~x757 & ~x759 & ~x760 & ~x761 & ~x764 & ~x765 & ~x767 & ~x773 & ~x775 & ~x776 & ~x777 & ~x778 & ~x779 & ~x780 & ~x781 & ~x782 & ~x783;
assign c29 =  x383 &  x495 & ~x51 & ~x77 & ~x147 & ~x204 & ~x436 & ~x501 & ~x584 & ~x644;
assign c211 =  x374 & ~x3 & ~x35 & ~x115 & ~x116 & ~x122 & ~x123 & ~x124 & ~x126 & ~x392 & ~x425 & ~x426 & ~x451 & ~x453 & ~x473 & ~x479 & ~x516 & ~x529 & ~x589 & ~x670 & ~x697 & ~x738 & ~x777;
assign c213 =  x323 &  x351 & ~x4 & ~x5 & ~x6 & ~x9 & ~x10 & ~x18 & ~x22 & ~x23 & ~x28 & ~x39 & ~x45 & ~x48 & ~x53 & ~x57 & ~x68 & ~x74 & ~x77 & ~x82 & ~x108 & ~x110 & ~x112 & ~x113 & ~x114 & ~x116 & ~x139 & ~x142 & ~x167 & ~x171 & ~x196 & ~x199 & ~x222 & ~x254 & ~x278 & ~x308 & ~x310 & ~x333 & ~x336 & ~x339 & ~x363 & ~x368 & ~x390 & ~x395 & ~x422 & ~x474 & ~x484 & ~x486 & ~x487 & ~x488 & ~x489 & ~x503 & ~x512 & ~x515 & ~x532 & ~x557 & ~x585 & ~x589 & ~x614 & ~x642 & ~x665 & ~x667 & ~x669 & ~x673 & ~x675 & ~x694 & ~x695 & ~x701 & ~x702 & ~x710 & ~x722 & ~x724 & ~x727 & ~x731 & ~x733 & ~x738 & ~x742 & ~x743 & ~x744 & ~x752 & ~x754 & ~x760 & ~x763 & ~x765 & ~x768 & ~x770 & ~x774 & ~x779 & ~x781;
assign c215 =  x315 &  x371 & ~x79 & ~x171 & ~x336 & ~x590 & ~x623 & ~x643 & ~x644 & ~x652 & ~x682 & ~x769 & ~x783;
assign c217 = ~x18 & ~x23 & ~x58 & ~x60 & ~x95 & ~x97 & ~x107 & ~x109 & ~x135 & ~x137 & ~x196 & ~x221 & ~x229 & ~x252 & ~x310 & ~x338 & ~x366 & ~x432 & ~x436 & ~x450 & ~x461 & ~x516 & ~x530 & ~x563 & ~x588 & ~x591 & ~x616 & ~x618 & ~x620 & ~x638 & ~x668 & ~x676 & ~x679 & ~x725 & ~x741 & ~x752 & ~x776 & ~x783;
assign c219 =  x498 & ~x18 & ~x50 & ~x253 & ~x491 & ~x492 & ~x493 & ~x756 & ~x776;
assign c221 =  x212 & ~x32 & ~x38 & ~x55 & ~x105 & ~x141 & ~x143 & ~x173 & ~x232 & ~x255 & ~x312 & ~x315 & ~x337 & ~x365 & ~x366 & ~x388 & ~x415 & ~x471 & ~x498 & ~x504 & ~x515 & ~x526 & ~x529 & ~x531 & ~x552 & ~x562 & ~x590 & ~x607 & ~x609 & ~x610 & ~x635 & ~x643 & ~x672 & ~x688 & ~x689 & ~x691 & ~x693 & ~x706 & ~x731 & ~x742 & ~x767 & ~x776;
assign c223 = ~x0 & ~x1 & ~x4 & ~x10 & ~x11 & ~x18 & ~x20 & ~x21 & ~x24 & ~x28 & ~x29 & ~x30 & ~x31 & ~x36 & ~x40 & ~x41 & ~x45 & ~x46 & ~x47 & ~x50 & ~x53 & ~x55 & ~x59 & ~x65 & ~x67 & ~x69 & ~x73 & ~x74 & ~x76 & ~x78 & ~x80 & ~x82 & ~x87 & ~x89 & ~x92 & ~x93 & ~x94 & ~x95 & ~x97 & ~x98 & ~x99 & ~x100 & ~x103 & ~x104 & ~x105 & ~x109 & ~x110 & ~x111 & ~x115 & ~x116 & ~x119 & ~x129 & ~x133 & ~x134 & ~x135 & ~x136 & ~x138 & ~x141 & ~x145 & ~x162 & ~x164 & ~x190 & ~x191 & ~x197 & ~x219 & ~x220 & ~x221 & ~x248 & ~x250 & ~x252 & ~x276 & ~x280 & ~x281 & ~x304 & ~x306 & ~x307 & ~x309 & ~x336 & ~x337 & ~x338 & ~x360 & ~x363 & ~x364 & ~x365 & ~x395 & ~x416 & ~x418 & ~x422 & ~x423 & ~x443 & ~x444 & ~x445 & ~x448 & ~x449 & ~x450 & ~x474 & ~x479 & ~x498 & ~x501 & ~x502 & ~x503 & ~x504 & ~x506 & ~x507 & ~x527 & ~x528 & ~x529 & ~x533 & ~x535 & ~x537 & ~x538 & ~x544 & ~x556 & ~x557 & ~x558 & ~x560 & ~x572 & ~x573 & ~x582 & ~x584 & ~x586 & ~x587 & ~x592 & ~x609 & ~x615 & ~x638 & ~x641 & ~x643 & ~x645 & ~x646 & ~x648 & ~x665 & ~x666 & ~x670 & ~x672 & ~x673 & ~x676 & ~x693 & ~x697 & ~x703 & ~x704 & ~x707 & ~x710 & ~x723 & ~x726 & ~x728 & ~x730 & ~x731 & ~x734 & ~x735 & ~x736 & ~x737 & ~x740 & ~x750 & ~x753 & ~x754 & ~x758 & ~x760 & ~x761 & ~x764 & ~x766 & ~x773 & ~x776 & ~x778 & ~x782;
assign c225 = ~x3 & ~x14 & ~x18 & ~x24 & ~x36 & ~x44 & ~x45 & ~x51 & ~x52 & ~x54 & ~x62 & ~x73 & ~x78 & ~x108 & ~x110 & ~x116 & ~x171 & ~x174 & ~x198 & ~x199 & ~x202 & ~x222 & ~x226 & ~x228 & ~x231 & ~x249 & ~x251 & ~x256 & ~x280 & ~x313 & ~x331 & ~x361 & ~x362 & ~x369 & ~x371 & ~x372 & ~x388 & ~x400 & ~x423 & ~x428 & ~x446 & ~x472 & ~x485 & ~x499 & ~x515 & ~x516 & ~x531 & ~x560 & ~x584 & ~x585 & ~x587 & ~x618 & ~x634 & ~x664 & ~x666 & ~x667 & ~x672 & ~x680 & ~x686 & ~x693 & ~x695 & ~x702 & ~x715 & ~x720 & ~x724 & ~x731 & ~x736 & ~x739 & ~x740 & ~x748 & ~x752 & ~x762 & ~x767 & ~x771 & ~x778;
assign c227 =  x318 &  x346 & ~x8 & ~x28 & ~x137 & ~x140 & ~x144 & ~x254 & ~x268 & ~x285 & ~x314 & ~x424 & ~x534 & ~x609 & ~x670 & ~x716 & ~x742 & ~x756 & ~x761 & ~x762 & ~x778 & ~x783;
assign c229 =  x373 &  x402 & ~x0 & ~x10 & ~x12 & ~x14 & ~x25 & ~x31 & ~x34 & ~x36 & ~x37 & ~x45 & ~x46 & ~x47 & ~x53 & ~x61 & ~x64 & ~x65 & ~x66 & ~x77 & ~x83 & ~x85 & ~x110 & ~x114 & ~x116 & ~x135 & ~x136 & ~x139 & ~x140 & ~x142 & ~x145 & ~x169 & ~x219 & ~x220 & ~x247 & ~x333 & ~x363 & ~x366 & ~x390 & ~x395 & ~x417 & ~x418 & ~x425 & ~x447 & ~x453 & ~x454 & ~x473 & ~x474 & ~x475 & ~x478 & ~x481 & ~x501 & ~x509 & ~x530 & ~x532 & ~x537 & ~x557 & ~x565 & ~x584 & ~x585 & ~x587 & ~x593 & ~x594 & ~x621 & ~x623 & ~x639 & ~x668 & ~x674 & ~x702 & ~x705 & ~x721 & ~x722 & ~x724 & ~x725 & ~x734 & ~x737 & ~x741 & ~x754 & ~x757 & ~x760 & ~x772 & ~x783;
assign c231 =  x407 &  x434 & ~x3 & ~x13 & ~x17 & ~x38 & ~x40 & ~x52 & ~x53 & ~x55 & ~x60 & ~x71 & ~x82 & ~x86 & ~x93 & ~x99 & ~x105 & ~x107 & ~x117 & ~x122 & ~x124 & ~x136 & ~x141 & ~x143 & ~x147 & ~x164 & ~x169 & ~x175 & ~x193 & ~x196 & ~x200 & ~x202 & ~x225 & ~x257 & ~x275 & ~x276 & ~x279 & ~x306 & ~x315 & ~x335 & ~x345 & ~x363 & ~x366 & ~x371 & ~x372 & ~x386 & ~x387 & ~x393 & ~x395 & ~x399 & ~x415 & ~x416 & ~x420 & ~x421 & ~x424 & ~x426 & ~x447 & ~x455 & ~x479 & ~x480 & ~x481 & ~x497 & ~x502 & ~x526 & ~x533 & ~x535 & ~x579 & ~x583 & ~x589 & ~x616 & ~x634 & ~x636 & ~x640 & ~x648 & ~x661 & ~x663 & ~x671 & ~x674 & ~x689 & ~x692 & ~x717 & ~x718 & ~x719 & ~x732 & ~x750 & ~x753 & ~x764 & ~x773 & ~x778 & ~x780;
assign c233 =  x288 &  x371 & ~x50 & ~x319;
assign c235 =  x239 & ~x3 & ~x10 & ~x36 & ~x38 & ~x41 & ~x46 & ~x56 & ~x67 & ~x75 & ~x78 & ~x85 & ~x98 & ~x104 & ~x105 & ~x111 & ~x118 & ~x121 & ~x137 & ~x141 & ~x163 & ~x191 & ~x192 & ~x193 & ~x197 & ~x198 & ~x201 & ~x225 & ~x226 & ~x229 & ~x251 & ~x252 & ~x254 & ~x284 & ~x307 & ~x310 & ~x312 & ~x314 & ~x339 & ~x361 & ~x362 & ~x364 & ~x386 & ~x388 & ~x393 & ~x414 & ~x415 & ~x416 & ~x420 & ~x423 & ~x444 & ~x445 & ~x448 & ~x468 & ~x480 & ~x503 & ~x507 & ~x525 & ~x533 & ~x534 & ~x535 & ~x552 & ~x553 & ~x554 & ~x559 & ~x560 & ~x580 & ~x583 & ~x584 & ~x592 & ~x608 & ~x634 & ~x637 & ~x642 & ~x660 & ~x662 & ~x673 & ~x689 & ~x695 & ~x700 & ~x714 & ~x716 & ~x718 & ~x720 & ~x724 & ~x731 & ~x732 & ~x734 & ~x737 & ~x744 & ~x748 & ~x751 & ~x754 & ~x763 & ~x770 & ~x771 & ~x775 & ~x776 & ~x779;
assign c237 =  x579 &  x606 & ~x1 & ~x5 & ~x8 & ~x13 & ~x21 & ~x24 & ~x27 & ~x34 & ~x35 & ~x37 & ~x39 & ~x43 & ~x44 & ~x46 & ~x48 & ~x64 & ~x66 & ~x72 & ~x75 & ~x77 & ~x80 & ~x83 & ~x87 & ~x106 & ~x108 & ~x112 & ~x113 & ~x114 & ~x118 & ~x137 & ~x170 & ~x194 & ~x198 & ~x221 & ~x248 & ~x277 & ~x280 & ~x305 & ~x306 & ~x308 & ~x363 & ~x419 & ~x450 & ~x477 & ~x478 & ~x486 & ~x502 & ~x503 & ~x517 & ~x518 & ~x520 & ~x531 & ~x534 & ~x555 & ~x583 & ~x584 & ~x588 & ~x610 & ~x612 & ~x639 & ~x646 & ~x692 & ~x695 & ~x697 & ~x699 & ~x702 & ~x706 & ~x712 & ~x727 & ~x728 & ~x735 & ~x741 & ~x744 & ~x745 & ~x757 & ~x764 & ~x769 & ~x776 & ~x780 & ~x782;
assign c239 =  x350 &  x351 &  x380 & ~x39 & ~x44 & ~x89 & ~x105 & ~x132 & ~x134 & ~x135 & ~x306 & ~x360 & ~x454 & ~x515 & ~x517 & ~x528 & ~x532 & ~x587 & ~x612 & ~x617 & ~x639 & ~x677 & ~x721 & ~x726 & ~x728 & ~x731 & ~x738 & ~x739 & ~x749 & ~x764;
assign c241 =  x288 &  x343 &  x371 &  x399 & ~x87 & ~x367 & ~x395 & ~x476;
assign c243 = ~x4 & ~x6 & ~x8 & ~x9 & ~x11 & ~x14 & ~x17 & ~x23 & ~x25 & ~x29 & ~x36 & ~x38 & ~x40 & ~x41 & ~x47 & ~x55 & ~x57 & ~x62 & ~x63 & ~x67 & ~x69 & ~x70 & ~x73 & ~x75 & ~x80 & ~x82 & ~x85 & ~x94 & ~x97 & ~x98 & ~x105 & ~x106 & ~x115 & ~x117 & ~x142 & ~x165 & ~x197 & ~x224 & ~x277 & ~x305 & ~x307 & ~x333 & ~x336 & ~x339 & ~x360 & ~x364 & ~x391 & ~x392 & ~x393 & ~x416 & ~x421 & ~x423 & ~x444 & ~x445 & ~x449 & ~x456 & ~x457 & ~x478 & ~x489 & ~x505 & ~x506 & ~x514 & ~x529 & ~x532 & ~x533 & ~x542 & ~x583 & ~x588 & ~x613 & ~x639 & ~x668 & ~x670 & ~x671 & ~x695 & ~x702 & ~x704 & ~x707 & ~x724 & ~x725 & ~x726 & ~x727 & ~x731 & ~x735 & ~x739 & ~x740 & ~x743 & ~x751 & ~x753 & ~x754 & ~x756 & ~x759 & ~x766 & ~x779;
assign c245 = ~x12 & ~x13 & ~x14 & ~x15 & ~x21 & ~x33 & ~x42 & ~x44 & ~x57 & ~x59 & ~x70 & ~x71 & ~x73 & ~x84 & ~x94 & ~x95 & ~x119 & ~x123 & ~x124 & ~x125 & ~x126 & ~x137 & ~x140 & ~x196 & ~x197 & ~x220 & ~x248 & ~x276 & ~x278 & ~x335 & ~x417 & ~x443 & ~x491 & ~x505 & ~x534 & ~x546 & ~x556 & ~x559 & ~x564 & ~x602 & ~x603 & ~x616 & ~x618 & ~x645 & ~x682 & ~x701 & ~x704 & ~x711 & ~x713 & ~x726 & ~x728 & ~x734 & ~x741 & ~x752 & ~x753 & ~x777 & ~x779 & ~x783;
assign c247 = ~x1 & ~x22 & ~x53 & ~x55 & ~x58 & ~x80 & ~x104 & ~x106 & ~x172 & ~x184 & ~x185 & ~x220 & ~x226 & ~x238 & ~x240 & ~x267 & ~x293 & ~x389 & ~x417 & ~x449 & ~x451 & ~x537 & ~x558 & ~x560 & ~x562 & ~x586 & ~x594 & ~x639 & ~x644 & ~x696 & ~x715 & ~x716 & ~x777 & ~x782;
assign c249 =  x345 &  x373 &  x401 & ~x14 & ~x31 & ~x46 & ~x65 & ~x66 & ~x84 & ~x89 & ~x116 & ~x123 & ~x146 & ~x199 & ~x252 & ~x254 & ~x423 & ~x424 & ~x445 & ~x447 & ~x448 & ~x452 & ~x477 & ~x507 & ~x533 & ~x555 & ~x562 & ~x582 & ~x587 & ~x610 & ~x612 & ~x613 & ~x617 & ~x620 & ~x646 & ~x673 & ~x711 & ~x725 & ~x730 & ~x746 & ~x747 & ~x756 & ~x771 & ~x772 & ~x775 & ~x782;
assign c251 = ~x2 & ~x17 & ~x18 & ~x22 & ~x24 & ~x30 & ~x51 & ~x54 & ~x70 & ~x73 & ~x78 & ~x79 & ~x82 & ~x117 & ~x166 & ~x254 & ~x260 & ~x280 & ~x312 & ~x316 & ~x366 & ~x384 & ~x385 & ~x391 & ~x399 & ~x457 & ~x497 & ~x498 & ~x499 & ~x504 & ~x523 & ~x551 & ~x554 & ~x559 & ~x579 & ~x580 & ~x583 & ~x608 & ~x633 & ~x636 & ~x669 & ~x674 & ~x713 & ~x719 & ~x738 & ~x744 & ~x757 & ~x760 & ~x781;
assign c253 = ~x1 & ~x2 & ~x16 & ~x21 & ~x22 & ~x43 & ~x50 & ~x65 & ~x68 & ~x72 & ~x74 & ~x79 & ~x83 & ~x86 & ~x91 & ~x105 & ~x109 & ~x110 & ~x117 & ~x123 & ~x124 & ~x146 & ~x148 & ~x168 & ~x172 & ~x196 & ~x201 & ~x224 & ~x306 & ~x308 & ~x315 & ~x391 & ~x415 & ~x419 & ~x429 & ~x442 & ~x447 & ~x455 & ~x467 & ~x470 & ~x474 & ~x494 & ~x497 & ~x523 & ~x527 & ~x528 & ~x533 & ~x562 & ~x564 & ~x578 & ~x579 & ~x583 & ~x610 & ~x613 & ~x634 & ~x646 & ~x661 & ~x664 & ~x666 & ~x671 & ~x689 & ~x690 & ~x697 & ~x715 & ~x720 & ~x723 & ~x726 & ~x730 & ~x752 & ~x753 & ~x760 & ~x764 & ~x765 & ~x767 & ~x777;
assign c255 =  x406 & ~x7 & ~x11 & ~x27 & ~x32 & ~x33 & ~x37 & ~x38 & ~x43 & ~x47 & ~x50 & ~x62 & ~x82 & ~x85 & ~x104 & ~x107 & ~x171 & ~x194 & ~x196 & ~x224 & ~x248 & ~x253 & ~x257 & ~x303 & ~x305 & ~x311 & ~x331 & ~x341 & ~x345 & ~x357 & ~x369 & ~x386 & ~x393 & ~x395 & ~x423 & ~x441 & ~x443 & ~x446 & ~x451 & ~x454 & ~x469 & ~x473 & ~x481 & ~x483 & ~x502 & ~x510 & ~x511 & ~x529 & ~x532 & ~x543 & ~x544 & ~x583 & ~x637 & ~x664 & ~x665 & ~x691 & ~x705 & ~x720 & ~x733 & ~x740 & ~x742 & ~x751 & ~x757 & ~x763 & ~x775 & ~x777 & ~x779 & ~x783;
assign c257 =  x384 & ~x1 & ~x3 & ~x8 & ~x9 & ~x10 & ~x11 & ~x17 & ~x18 & ~x20 & ~x21 & ~x22 & ~x23 & ~x26 & ~x28 & ~x33 & ~x35 & ~x36 & ~x37 & ~x41 & ~x44 & ~x46 & ~x48 & ~x58 & ~x59 & ~x60 & ~x61 & ~x76 & ~x77 & ~x84 & ~x86 & ~x91 & ~x104 & ~x112 & ~x115 & ~x139 & ~x163 & ~x167 & ~x168 & ~x170 & ~x190 & ~x191 & ~x220 & ~x222 & ~x226 & ~x227 & ~x247 & ~x254 & ~x279 & ~x308 & ~x333 & ~x337 & ~x362 & ~x365 & ~x391 & ~x394 & ~x419 & ~x421 & ~x449 & ~x476 & ~x477 & ~x493 & ~x505 & ~x534 & ~x536 & ~x557 & ~x558 & ~x560 & ~x561 & ~x564 & ~x585 & ~x587 & ~x589 & ~x592 & ~x620 & ~x640 & ~x642 & ~x643 & ~x645 & ~x649 & ~x668 & ~x670 & ~x672 & ~x674 & ~x701 & ~x703 & ~x704 & ~x710 & ~x711 & ~x712 & ~x715 & ~x720 & ~x724 & ~x727 & ~x730 & ~x731 & ~x738 & ~x750 & ~x751 & ~x755 & ~x756 & ~x759 & ~x763 & ~x768 & ~x769 & ~x771 & ~x775 & ~x781;
assign c259 =  x220;
assign c261 = ~x56 & ~x62 & ~x153 & ~x335 & ~x348 & ~x441 & ~x499 & ~x523 & ~x539 & ~x577 & ~x605 & ~x641 & ~x689 & ~x717 & ~x728;
assign c263 =  x287 &  x370 &  x398 & ~x4 & ~x5 & ~x6 & ~x13 & ~x40 & ~x59 & ~x90 & ~x199 & ~x200 & ~x254 & ~x502 & ~x505 & ~x613 & ~x648 & ~x733;
assign c265 =  x351 & ~x5 & ~x11 & ~x16 & ~x23 & ~x24 & ~x26 & ~x27 & ~x34 & ~x36 & ~x50 & ~x91 & ~x95 & ~x100 & ~x101 & ~x118 & ~x120 & ~x121 & ~x122 & ~x141 & ~x143 & ~x148 & ~x169 & ~x172 & ~x290 & ~x308 & ~x316 & ~x360 & ~x366 & ~x414 & ~x423 & ~x426 & ~x442 & ~x446 & ~x455 & ~x498 & ~x499 & ~x527 & ~x554 & ~x613 & ~x635 & ~x642 & ~x661 & ~x662 & ~x672 & ~x714 & ~x738 & ~x747 & ~x749 & ~x769;
assign c267 =  x442 &  x470 & ~x167 & ~x465 & ~x532 & ~x757;
assign c269 =  x409 &  x574 & ~x244 & ~x297 & ~x623;
assign c271 =  x319 &  x347 & ~x4 & ~x6 & ~x18 & ~x58 & ~x63 & ~x82 & ~x92 & ~x108 & ~x109 & ~x146 & ~x169 & ~x202 & ~x223 & ~x341 & ~x389 & ~x391 & ~x396 & ~x422 & ~x463 & ~x476 & ~x477 & ~x503 & ~x504 & ~x529 & ~x557 & ~x559 & ~x582 & ~x618 & ~x638 & ~x644 & ~x666 & ~x669 & ~x699 & ~x704 & ~x706 & ~x720 & ~x723 & ~x732 & ~x742 & ~x747 & ~x753 & ~x756 & ~x763 & ~x764 & ~x777;
assign c273 =  x713 & ~x599;
assign c275 =  x525 &  x580 &  x607 & ~x12 & ~x141 & ~x250 & ~x279 & ~x492 & ~x518 & ~x519 & ~x520 & ~x584 & ~x614 & ~x616 & ~x678 & ~x727 & ~x760 & ~x766;
assign c277 =  x374 &  x601 & ~x15 & ~x20 & ~x28 & ~x35 & ~x121 & ~x125 & ~x138 & ~x154 & ~x337 & ~x452 & ~x473 & ~x588 & ~x698 & ~x727 & ~x780;
assign c279 =  x349 & ~x21 & ~x34 & ~x40 & ~x69 & ~x93 & ~x96 & ~x118 & ~x122 & ~x147 & ~x171 & ~x222 & ~x255 & ~x260 & ~x285 & ~x312 & ~x315 & ~x316 & ~x355 & ~x421 & ~x443 & ~x474 & ~x499 & ~x581 & ~x587 & ~x609 & ~x611 & ~x616 & ~x665 & ~x666 & ~x684 & ~x693 & ~x695 & ~x698 & ~x774;
assign c281 =  x548 & ~x4 & ~x9 & ~x11 & ~x18 & ~x19 & ~x20 & ~x21 & ~x22 & ~x32 & ~x34 & ~x42 & ~x44 & ~x51 & ~x53 & ~x56 & ~x58 & ~x60 & ~x61 & ~x82 & ~x83 & ~x85 & ~x86 & ~x90 & ~x109 & ~x113 & ~x115 & ~x116 & ~x121 & ~x136 & ~x137 & ~x141 & ~x146 & ~x147 & ~x148 & ~x168 & ~x169 & ~x171 & ~x176 & ~x193 & ~x198 & ~x203 & ~x204 & ~x222 & ~x225 & ~x226 & ~x230 & ~x257 & ~x277 & ~x280 & ~x282 & ~x287 & ~x307 & ~x308 & ~x311 & ~x312 & ~x327 & ~x328 & ~x334 & ~x337 & ~x339 & ~x358 & ~x360 & ~x362 & ~x392 & ~x393 & ~x417 & ~x419 & ~x421 & ~x422 & ~x423 & ~x425 & ~x446 & ~x449 & ~x451 & ~x471 & ~x472 & ~x474 & ~x476 & ~x478 & ~x479 & ~x500 & ~x505 & ~x506 & ~x526 & ~x529 & ~x532 & ~x534 & ~x555 & ~x557 & ~x561 & ~x580 & ~x581 & ~x582 & ~x589 & ~x590 & ~x607 & ~x615 & ~x636 & ~x642 & ~x645 & ~x664 & ~x666 & ~x668 & ~x675 & ~x691 & ~x692 & ~x693 & ~x700 & ~x701 & ~x702 & ~x703 & ~x709 & ~x711 & ~x716 & ~x719 & ~x727 & ~x728 & ~x729 & ~x732 & ~x740 & ~x745 & ~x748 & ~x749 & ~x750 & ~x753 & ~x756 & ~x758 & ~x759 & ~x760 & ~x765 & ~x767 & ~x770 & ~x772 & ~x773 & ~x777 & ~x778;
assign c283 =  x321 &  x322 &  x350 &  x379 & ~x0 & ~x7 & ~x51 & ~x59 & ~x96 & ~x115 & ~x118 & ~x120 & ~x137 & ~x171 & ~x223 & ~x279 & ~x283 & ~x305 & ~x306 & ~x308 & ~x361 & ~x362 & ~x367 & ~x368 & ~x388 & ~x389 & ~x398 & ~x400 & ~x419 & ~x422 & ~x423 & ~x444 & ~x445 & ~x452 & ~x454 & ~x471 & ~x473 & ~x498 & ~x502 & ~x525 & ~x526 & ~x527 & ~x530 & ~x559 & ~x581 & ~x584 & ~x586 & ~x590 & ~x610 & ~x612 & ~x616 & ~x619 & ~x642 & ~x643 & ~x664 & ~x665 & ~x666 & ~x669 & ~x676 & ~x699 & ~x702 & ~x706 & ~x728 & ~x730 & ~x733 & ~x740 & ~x752 & ~x769 & ~x771;
assign c285 =  x292 &  x347 &  x573 & ~x121 & ~x150 & ~x286 & ~x636 & ~x660 & ~x661;
assign c287 =  x578 & ~x2 & ~x3 & ~x8 & ~x9 & ~x20 & ~x22 & ~x25 & ~x37 & ~x39 & ~x51 & ~x53 & ~x57 & ~x58 & ~x60 & ~x61 & ~x62 & ~x72 & ~x78 & ~x81 & ~x86 & ~x89 & ~x90 & ~x91 & ~x99 & ~x107 & ~x110 & ~x111 & ~x115 & ~x117 & ~x119 & ~x127 & ~x138 & ~x140 & ~x141 & ~x143 & ~x144 & ~x145 & ~x147 & ~x165 & ~x168 & ~x191 & ~x192 & ~x193 & ~x226 & ~x247 & ~x254 & ~x255 & ~x277 & ~x281 & ~x309 & ~x335 & ~x336 & ~x343 & ~x360 & ~x364 & ~x367 & ~x370 & ~x371 & ~x392 & ~x393 & ~x394 & ~x396 & ~x398 & ~x417 & ~x420 & ~x444 & ~x447 & ~x448 & ~x450 & ~x454 & ~x472 & ~x477 & ~x478 & ~x500 & ~x508 & ~x528 & ~x530 & ~x533 & ~x536 & ~x554 & ~x555 & ~x556 & ~x557 & ~x562 & ~x563 & ~x585 & ~x589 & ~x593 & ~x594 & ~x609 & ~x610 & ~x637 & ~x639 & ~x643 & ~x645 & ~x665 & ~x667 & ~x669 & ~x670 & ~x676 & ~x680 & ~x695 & ~x702 & ~x703 & ~x720 & ~x723 & ~x725 & ~x730 & ~x736 & ~x739 & ~x753 & ~x756 & ~x757 & ~x758 & ~x759 & ~x761 & ~x766 & ~x770 & ~x771 & ~x773 & ~x779 & ~x783;
assign c289 = ~x1 & ~x10 & ~x12 & ~x16 & ~x51 & ~x70 & ~x82 & ~x89 & ~x106 & ~x108 & ~x118 & ~x123 & ~x149 & ~x166 & ~x193 & ~x197 & ~x252 & ~x256 & ~x308 & ~x338 & ~x342 & ~x360 & ~x364 & ~x373 & ~x390 & ~x392 & ~x399 & ~x414 & ~x440 & ~x451 & ~x471 & ~x475 & ~x477 & ~x479 & ~x483 & ~x498 & ~x522 & ~x523 & ~x528 & ~x534 & ~x551 & ~x561 & ~x578 & ~x589 & ~x605 & ~x607 & ~x643 & ~x660 & ~x669 & ~x695 & ~x726 & ~x730;
assign c291 =  x299 &  x302 & ~x158 & ~x187;
assign c293 =  x465 &  x685 & ~x63 & ~x71 & ~x80 & ~x82 & ~x125 & ~x252 & ~x447 & ~x564 & ~x694 & ~x734 & ~x759;
assign c295 =  x261 & ~x1 & ~x8 & ~x14 & ~x20 & ~x25 & ~x27 & ~x28 & ~x29 & ~x39 & ~x44 & ~x46 & ~x50 & ~x52 & ~x53 & ~x68 & ~x71 & ~x78 & ~x81 & ~x87 & ~x105 & ~x107 & ~x132 & ~x135 & ~x146 & ~x162 & ~x166 & ~x169 & ~x171 & ~x193 & ~x194 & ~x195 & ~x197 & ~x198 & ~x199 & ~x222 & ~x224 & ~x246 & ~x274 & ~x275 & ~x278 & ~x279 & ~x303 & ~x305 & ~x306 & ~x309 & ~x336 & ~x337 & ~x360 & ~x361 & ~x365 & ~x417 & ~x418 & ~x420 & ~x443 & ~x444 & ~x447 & ~x451 & ~x475 & ~x499 & ~x500 & ~x508 & ~x526 & ~x527 & ~x531 & ~x533 & ~x534 & ~x535 & ~x537 & ~x555 & ~x559 & ~x561 & ~x567 & ~x588 & ~x592 & ~x611 & ~x616 & ~x617 & ~x619 & ~x620 & ~x621 & ~x622 & ~x624 & ~x625 & ~x638 & ~x639 & ~x641 & ~x642 & ~x666 & ~x667 & ~x669 & ~x672 & ~x680 & ~x695 & ~x696 & ~x704 & ~x705 & ~x726 & ~x728 & ~x731 & ~x752 & ~x757 & ~x765 & ~x767 & ~x768 & ~x777 & ~x783;
assign c297 =  x682 & ~x156;
assign c299 = ~x3 & ~x5 & ~x12 & ~x14 & ~x16 & ~x19 & ~x21 & ~x24 & ~x25 & ~x27 & ~x33 & ~x41 & ~x42 & ~x45 & ~x48 & ~x50 & ~x54 & ~x56 & ~x57 & ~x68 & ~x72 & ~x73 & ~x79 & ~x84 & ~x85 & ~x91 & ~x107 & ~x110 & ~x112 & ~x115 & ~x137 & ~x194 & ~x197 & ~x220 & ~x227 & ~x249 & ~x277 & ~x328 & ~x333 & ~x390 & ~x391 & ~x394 & ~x417 & ~x418 & ~x457 & ~x458 & ~x474 & ~x478 & ~x485 & ~x486 & ~x488 & ~x489 & ~x490 & ~x514 & ~x516 & ~x517 & ~x519 & ~x529 & ~x587 & ~x615 & ~x643 & ~x694 & ~x695 & ~x704 & ~x706 & ~x714 & ~x728 & ~x730 & ~x733 & ~x735 & ~x744 & ~x749 & ~x751 & ~x774 & ~x776 & ~x778 & ~x779;
assign c2101 =  x380 &  x407 &  x492 &  x520 & ~x11 & ~x12 & ~x19 & ~x55 & ~x74 & ~x94 & ~x95 & ~x96 & ~x114 & ~x146 & ~x149 & ~x194 & ~x195 & ~x278 & ~x306 & ~x313 & ~x341 & ~x386 & ~x414 & ~x427 & ~x444 & ~x448 & ~x451 & ~x524 & ~x579 & ~x580 & ~x607 & ~x663 & ~x671 & ~x701 & ~x703 & ~x725 & ~x730 & ~x780;
assign c2103 =  x270 & ~x7 & ~x8 & ~x12 & ~x22 & ~x30 & ~x41 & ~x49 & ~x69 & ~x78 & ~x99 & ~x110 & ~x128 & ~x139 & ~x154 & ~x155 & ~x169 & ~x181 & ~x183 & ~x308 & ~x449 & ~x473 & ~x508 & ~x509 & ~x510 & ~x540 & ~x557 & ~x565 & ~x568 & ~x588 & ~x593 & ~x618 & ~x701 & ~x729 & ~x762;
assign c2105 =  x348 &  x381 &  x629 &  x630 & ~x8 & ~x9 & ~x12 & ~x15 & ~x18 & ~x19 & ~x28 & ~x35 & ~x38 & ~x46 & ~x48 & ~x58 & ~x59 & ~x60 & ~x62 & ~x71 & ~x79 & ~x88 & ~x105 & ~x107 & ~x110 & ~x113 & ~x116 & ~x142 & ~x167 & ~x168 & ~x251 & ~x252 & ~x279 & ~x282 & ~x311 & ~x361 & ~x365 & ~x366 & ~x369 & ~x390 & ~x399 & ~x419 & ~x421 & ~x422 & ~x423 & ~x443 & ~x472 & ~x476 & ~x503 & ~x506 & ~x557 & ~x586 & ~x588 & ~x639 & ~x649 & ~x669 & ~x671 & ~x675 & ~x678 & ~x695 & ~x696 & ~x698 & ~x704 & ~x708 & ~x717 & ~x718 & ~x719 & ~x723 & ~x734 & ~x739 & ~x740 & ~x744 & ~x748 & ~x751 & ~x765 & ~x767 & ~x778 & ~x781 & ~x782;
assign c2107 =  x496 &  x524 & ~x0 & ~x1 & ~x2 & ~x5 & ~x11 & ~x13 & ~x14 & ~x15 & ~x16 & ~x17 & ~x27 & ~x29 & ~x30 & ~x33 & ~x36 & ~x38 & ~x42 & ~x43 & ~x49 & ~x50 & ~x54 & ~x60 & ~x63 & ~x64 & ~x65 & ~x66 & ~x67 & ~x69 & ~x70 & ~x73 & ~x77 & ~x78 & ~x79 & ~x87 & ~x89 & ~x94 & ~x95 & ~x97 & ~x98 & ~x103 & ~x109 & ~x110 & ~x112 & ~x114 & ~x139 & ~x141 & ~x143 & ~x163 & ~x165 & ~x169 & ~x170 & ~x193 & ~x194 & ~x198 & ~x224 & ~x225 & ~x249 & ~x256 & ~x277 & ~x284 & ~x305 & ~x306 & ~x308 & ~x334 & ~x338 & ~x339 & ~x360 & ~x362 & ~x366 & ~x367 & ~x390 & ~x420 & ~x421 & ~x422 & ~x423 & ~x446 & ~x447 & ~x448 & ~x472 & ~x473 & ~x475 & ~x476 & ~x491 & ~x501 & ~x502 & ~x519 & ~x520 & ~x529 & ~x532 & ~x555 & ~x558 & ~x559 & ~x560 & ~x561 & ~x584 & ~x585 & ~x589 & ~x611 & ~x642 & ~x644 & ~x645 & ~x669 & ~x674 & ~x696 & ~x699 & ~x701 & ~x703 & ~x705 & ~x706 & ~x716 & ~x725 & ~x726 & ~x728 & ~x731 & ~x732 & ~x735 & ~x737 & ~x738 & ~x739 & ~x741 & ~x745 & ~x746 & ~x747 & ~x748 & ~x749 & ~x753 & ~x755 & ~x757 & ~x763 & ~x764 & ~x766 & ~x771 & ~x773 & ~x781;
assign c2109 =  x349 &  x377 & ~x2 & ~x35 & ~x36 & ~x37 & ~x39 & ~x45 & ~x56 & ~x60 & ~x62 & ~x63 & ~x64 & ~x65 & ~x68 & ~x75 & ~x76 & ~x90 & ~x93 & ~x95 & ~x98 & ~x99 & ~x101 & ~x106 & ~x110 & ~x113 & ~x135 & ~x138 & ~x141 & ~x147 & ~x169 & ~x176 & ~x199 & ~x250 & ~x256 & ~x278 & ~x306 & ~x307 & ~x310 & ~x314 & ~x332 & ~x368 & ~x369 & ~x370 & ~x391 & ~x396 & ~x414 & ~x469 & ~x470 & ~x471 & ~x472 & ~x476 & ~x499 & ~x507 & ~x524 & ~x525 & ~x526 & ~x528 & ~x529 & ~x533 & ~x552 & ~x553 & ~x557 & ~x581 & ~x582 & ~x584 & ~x609 & ~x610 & ~x614 & ~x636 & ~x637 & ~x639 & ~x665 & ~x669 & ~x690 & ~x691 & ~x700 & ~x711 & ~x720 & ~x723 & ~x727 & ~x729 & ~x752 & ~x753 & ~x764 & ~x770;
assign c2111 =  x350 &  x351 & ~x1 & ~x6 & ~x10 & ~x11 & ~x14 & ~x15 & ~x18 & ~x20 & ~x22 & ~x25 & ~x26 & ~x27 & ~x30 & ~x33 & ~x36 & ~x40 & ~x44 & ~x45 & ~x46 & ~x48 & ~x49 & ~x50 & ~x52 & ~x54 & ~x57 & ~x59 & ~x62 & ~x65 & ~x77 & ~x79 & ~x80 & ~x81 & ~x84 & ~x85 & ~x86 & ~x88 & ~x90 & ~x91 & ~x92 & ~x93 & ~x103 & ~x104 & ~x108 & ~x110 & ~x111 & ~x114 & ~x136 & ~x137 & ~x163 & ~x168 & ~x194 & ~x196 & ~x220 & ~x222 & ~x224 & ~x226 & ~x248 & ~x253 & ~x282 & ~x283 & ~x303 & ~x307 & ~x308 & ~x310 & ~x311 & ~x334 & ~x335 & ~x336 & ~x359 & ~x360 & ~x361 & ~x364 & ~x366 & ~x367 & ~x368 & ~x389 & ~x391 & ~x393 & ~x394 & ~x415 & ~x417 & ~x418 & ~x420 & ~x421 & ~x446 & ~x447 & ~x449 & ~x452 & ~x453 & ~x454 & ~x478 & ~x483 & ~x485 & ~x487 & ~x488 & ~x500 & ~x503 & ~x505 & ~x528 & ~x529 & ~x531 & ~x557 & ~x585 & ~x586 & ~x617 & ~x640 & ~x641 & ~x645 & ~x665 & ~x667 & ~x671 & ~x674 & ~x676 & ~x693 & ~x694 & ~x695 & ~x702 & ~x705 & ~x708 & ~x709 & ~x710 & ~x712 & ~x716 & ~x721 & ~x722 & ~x725 & ~x726 & ~x729 & ~x734 & ~x737 & ~x739 & ~x740 & ~x746 & ~x754 & ~x755 & ~x756 & ~x762 & ~x763 & ~x765 & ~x769 & ~x771 & ~x774 & ~x777 & ~x782 & ~x783;
assign c2113 =  x317 &  x372 & ~x111 & ~x424 & ~x449 & ~x667 & ~x738;
assign c2115 =  x318 & ~x62 & ~x226 & ~x251 & ~x270 & ~x293 & ~x451 & ~x481 & ~x501 & ~x561 & ~x564 & ~x615 & ~x668 & ~x714;
assign c2117 =  x287 &  x315 &  x343 & ~x389 & ~x546;
assign c2119 =  x346 &  x374 &  x544 & ~x26 & ~x27 & ~x148 & ~x198 & ~x307 & ~x340 & ~x418 & ~x425 & ~x476 & ~x554 & ~x558 & ~x611 & ~x619 & ~x620 & ~x636 & ~x640 & ~x643 & ~x741 & ~x744 & ~x783;
assign c2121 =  x348 & ~x10 & ~x13 & ~x14 & ~x17 & ~x18 & ~x23 & ~x27 & ~x34 & ~x37 & ~x57 & ~x60 & ~x61 & ~x62 & ~x66 & ~x69 & ~x74 & ~x77 & ~x82 & ~x83 & ~x88 & ~x89 & ~x90 & ~x93 & ~x104 & ~x105 & ~x108 & ~x111 & ~x112 & ~x136 & ~x137 & ~x139 & ~x141 & ~x143 & ~x166 & ~x195 & ~x197 & ~x221 & ~x222 & ~x225 & ~x226 & ~x251 & ~x252 & ~x253 & ~x283 & ~x284 & ~x311 & ~x330 & ~x336 & ~x338 & ~x339 & ~x341 & ~x363 & ~x364 & ~x367 & ~x370 & ~x371 & ~x387 & ~x394 & ~x395 & ~x399 & ~x416 & ~x419 & ~x421 & ~x426 & ~x445 & ~x454 & ~x457 & ~x473 & ~x475 & ~x485 & ~x528 & ~x585 & ~x586 & ~x616 & ~x640 & ~x642 & ~x643 & ~x644 & ~x653 & ~x654 & ~x665 & ~x675 & ~x678 & ~x693 & ~x694 & ~x696 & ~x700 & ~x704 & ~x706 & ~x708 & ~x709 & ~x710 & ~x711 & ~x720 & ~x721 & ~x731 & ~x737 & ~x740 & ~x755 & ~x756 & ~x759 & ~x764 & ~x765 & ~x766 & ~x768 & ~x772 & ~x773;
assign c2123 = ~x2 & ~x11 & ~x17 & ~x21 & ~x27 & ~x35 & ~x48 & ~x57 & ~x66 & ~x70 & ~x77 & ~x81 & ~x92 & ~x93 & ~x105 & ~x108 & ~x110 & ~x111 & ~x114 & ~x117 & ~x135 & ~x143 & ~x164 & ~x166 & ~x190 & ~x307 & ~x309 & ~x310 & ~x335 & ~x364 & ~x367 & ~x403 & ~x433 & ~x459 & ~x460 & ~x461 & ~x487 & ~x488 & ~x505 & ~x518 & ~x519 & ~x558 & ~x613 & ~x614 & ~x640 & ~x644 & ~x666 & ~x668 & ~x669 & ~x675 & ~x698 & ~x701 & ~x702 & ~x706 & ~x707 & ~x711 & ~x722 & ~x730 & ~x732 & ~x740 & ~x747 & ~x749 & ~x751 & ~x761 & ~x767 & ~x769 & ~x773 & ~x780;
assign c2125 = ~x3 & ~x4 & ~x12 & ~x15 & ~x25 & ~x26 & ~x27 & ~x29 & ~x30 & ~x32 & ~x35 & ~x44 & ~x50 & ~x52 & ~x56 & ~x57 & ~x59 & ~x60 & ~x63 & ~x64 & ~x68 & ~x76 & ~x77 & ~x79 & ~x81 & ~x85 & ~x87 & ~x89 & ~x90 & ~x92 & ~x115 & ~x116 & ~x119 & ~x120 & ~x121 & ~x123 & ~x135 & ~x141 & ~x142 & ~x147 & ~x149 & ~x163 & ~x166 & ~x167 & ~x168 & ~x171 & ~x172 & ~x193 & ~x194 & ~x195 & ~x196 & ~x198 & ~x199 & ~x200 & ~x224 & ~x226 & ~x227 & ~x248 & ~x249 & ~x253 & ~x282 & ~x307 & ~x309 & ~x310 & ~x313 & ~x334 & ~x336 & ~x337 & ~x339 & ~x342 & ~x359 & ~x360 & ~x362 & ~x363 & ~x364 & ~x365 & ~x388 & ~x389 & ~x390 & ~x396 & ~x417 & ~x418 & ~x424 & ~x442 & ~x443 & ~x444 & ~x448 & ~x449 & ~x451 & ~x452 & ~x471 & ~x498 & ~x499 & ~x501 & ~x502 & ~x503 & ~x505 & ~x508 & ~x510 & ~x526 & ~x529 & ~x532 & ~x533 & ~x534 & ~x535 & ~x553 & ~x554 & ~x555 & ~x557 & ~x558 & ~x566 & ~x567 & ~x579 & ~x580 & ~x581 & ~x583 & ~x584 & ~x587 & ~x592 & ~x593 & ~x594 & ~x607 & ~x611 & ~x618 & ~x622 & ~x624 & ~x635 & ~x636 & ~x637 & ~x638 & ~x639 & ~x645 & ~x646 & ~x648 & ~x649 & ~x651 & ~x652 & ~x664 & ~x670 & ~x671 & ~x674 & ~x675 & ~x679 & ~x680 & ~x688 & ~x689 & ~x693 & ~x694 & ~x697 & ~x698 & ~x702 & ~x703 & ~x706 & ~x713 & ~x716 & ~x719 & ~x720 & ~x725 & ~x726 & ~x728 & ~x729 & ~x734 & ~x735 & ~x738 & ~x748 & ~x749 & ~x752 & ~x755 & ~x756 & ~x757 & ~x759 & ~x765 & ~x766 & ~x768 & ~x772 & ~x780 & ~x781 & ~x782;
assign c2127 =  x319 &  x401 & ~x11 & ~x32 & ~x46 & ~x50 & ~x63 & ~x85 & ~x90 & ~x120 & ~x122 & ~x124 & ~x149 & ~x200 & ~x203 & ~x251 & ~x254 & ~x335 & ~x337 & ~x389 & ~x391 & ~x423 & ~x425 & ~x504 & ~x557 & ~x616 & ~x647 & ~x666 & ~x675 & ~x678 & ~x718 & ~x728 & ~x744 & ~x748 & ~x759 & ~x763 & ~x765 & ~x772 & ~x782;
assign c2129 =  x352 &  x377 & ~x10 & ~x58 & ~x60 & ~x87 & ~x98 & ~x103 & ~x111 & ~x112 & ~x134 & ~x139 & ~x168 & ~x171 & ~x252 & ~x277 & ~x334 & ~x385 & ~x394 & ~x415 & ~x417 & ~x454 & ~x478 & ~x484 & ~x486 & ~x502 & ~x504 & ~x614 & ~x644 & ~x645 & ~x667 & ~x695 & ~x700 & ~x701 & ~x740 & ~x744 & ~x753 & ~x760 & ~x774 & ~x780;
assign c2131 =  x687 & ~x16 & ~x23 & ~x339 & ~x473 & ~x566 & ~x573 & ~x588 & ~x596 & ~x696 & ~x700 & ~x768 & ~x770;
assign c2133 =  x399 &  x427 & ~x32 & ~x36 & ~x55 & ~x105 & ~x109 & ~x123 & ~x142 & ~x166 & ~x223 & ~x249 & ~x309 & ~x365 & ~x377 & ~x404 & ~x419 & ~x449 & ~x557 & ~x586 & ~x672 & ~x676 & ~x679 & ~x712 & ~x728 & ~x730 & ~x741 & ~x768 & ~x772 & ~x782;
assign c2135 =  x387 &  x398;
assign c2137 =  x707;
assign c2139 =  x216 &  x380 &  x381 & ~x3 & ~x50 & ~x100 & ~x102 & ~x103 & ~x361 & ~x477 & ~x661 & ~x697 & ~x730 & ~x761;
assign c2141 =  x353 &  x377 & ~x400 & ~x427 & ~x486;
assign c2143 = ~x0 & ~x22 & ~x34 & ~x55 & ~x66 & ~x89 & ~x99 & ~x102 & ~x103 & ~x107 & ~x111 & ~x116 & ~x128 & ~x133 & ~x139 & ~x151 & ~x153 & ~x164 & ~x170 & ~x196 & ~x224 & ~x225 & ~x249 & ~x348 & ~x389 & ~x394 & ~x416 & ~x473 & ~x477 & ~x482 & ~x499 & ~x500 & ~x527 & ~x536 & ~x539 & ~x554 & ~x555 & ~x568 & ~x570 & ~x581 & ~x612 & ~x616 & ~x636 & ~x637 & ~x645 & ~x664 & ~x692 & ~x693 & ~x696 & ~x698 & ~x720 & ~x724 & ~x749 & ~x750 & ~x752 & ~x758 & ~x775 & ~x776;
assign c2145 =  x522 &  x550 &  x577 & ~x0 & ~x1 & ~x2 & ~x3 & ~x6 & ~x7 & ~x8 & ~x9 & ~x10 & ~x11 & ~x13 & ~x15 & ~x16 & ~x17 & ~x18 & ~x19 & ~x23 & ~x24 & ~x26 & ~x27 & ~x29 & ~x32 & ~x33 & ~x35 & ~x36 & ~x37 & ~x38 & ~x39 & ~x40 & ~x41 & ~x42 & ~x43 & ~x44 & ~x45 & ~x46 & ~x47 & ~x48 & ~x49 & ~x50 & ~x51 & ~x52 & ~x53 & ~x54 & ~x57 & ~x58 & ~x59 & ~x60 & ~x61 & ~x64 & ~x65 & ~x67 & ~x71 & ~x73 & ~x79 & ~x80 & ~x81 & ~x83 & ~x84 & ~x86 & ~x87 & ~x89 & ~x90 & ~x92 & ~x93 & ~x106 & ~x107 & ~x109 & ~x110 & ~x111 & ~x112 & ~x115 & ~x116 & ~x117 & ~x118 & ~x119 & ~x120 & ~x135 & ~x136 & ~x137 & ~x139 & ~x140 & ~x143 & ~x144 & ~x145 & ~x146 & ~x147 & ~x148 & ~x167 & ~x171 & ~x172 & ~x174 & ~x192 & ~x195 & ~x197 & ~x198 & ~x199 & ~x200 & ~x202 & ~x219 & ~x220 & ~x221 & ~x224 & ~x225 & ~x227 & ~x228 & ~x230 & ~x246 & ~x247 & ~x248 & ~x249 & ~x252 & ~x253 & ~x255 & ~x256 & ~x257 & ~x258 & ~x259 & ~x275 & ~x276 & ~x278 & ~x279 & ~x280 & ~x283 & ~x284 & ~x285 & ~x286 & ~x302 & ~x303 & ~x304 & ~x305 & ~x306 & ~x307 & ~x308 & ~x309 & ~x331 & ~x333 & ~x334 & ~x337 & ~x340 & ~x341 & ~x363 & ~x365 & ~x366 & ~x367 & ~x389 & ~x391 & ~x392 & ~x393 & ~x394 & ~x418 & ~x419 & ~x420 & ~x421 & ~x423 & ~x444 & ~x445 & ~x446 & ~x447 & ~x448 & ~x449 & ~x452 & ~x472 & ~x474 & ~x475 & ~x478 & ~x500 & ~x502 & ~x503 & ~x504 & ~x506 & ~x526 & ~x527 & ~x528 & ~x532 & ~x554 & ~x555 & ~x557 & ~x559 & ~x580 & ~x581 & ~x583 & ~x589 & ~x590 & ~x608 & ~x609 & ~x611 & ~x612 & ~x617 & ~x618 & ~x619 & ~x621 & ~x636 & ~x638 & ~x639 & ~x640 & ~x641 & ~x642 & ~x645 & ~x647 & ~x648 & ~x649 & ~x665 & ~x666 & ~x667 & ~x668 & ~x670 & ~x673 & ~x674 & ~x675 & ~x676 & ~x677 & ~x678 & ~x681 & ~x682 & ~x691 & ~x692 & ~x696 & ~x697 & ~x698 & ~x699 & ~x700 & ~x702 & ~x705 & ~x707 & ~x708 & ~x709 & ~x711 & ~x712 & ~x714 & ~x723 & ~x724 & ~x725 & ~x726 & ~x727 & ~x730 & ~x731 & ~x733 & ~x734 & ~x735 & ~x736 & ~x737 & ~x738 & ~x740 & ~x741 & ~x742 & ~x743 & ~x744 & ~x745 & ~x749 & ~x750 & ~x752 & ~x758 & ~x759 & ~x761 & ~x762 & ~x763 & ~x766 & ~x768 & ~x769 & ~x770 & ~x772 & ~x774 & ~x775 & ~x777 & ~x778 & ~x779 & ~x780 & ~x781 & ~x783;
assign c2147 =  x348 & ~x2 & ~x26 & ~x30 & ~x39 & ~x40 & ~x45 & ~x47 & ~x65 & ~x85 & ~x116 & ~x122 & ~x125 & ~x127 & ~x167 & ~x194 & ~x198 & ~x305 & ~x310 & ~x333 & ~x341 & ~x388 & ~x419 & ~x443 & ~x470 & ~x475 & ~x476 & ~x497 & ~x499 & ~x500 & ~x526 & ~x528 & ~x560 & ~x581 & ~x582 & ~x608 & ~x611 & ~x614 & ~x616 & ~x639 & ~x643 & ~x691 & ~x697 & ~x698 & ~x701 & ~x705 & ~x711 & ~x758 & ~x765 & ~x777;
assign c2149 =  x242 & ~x6 & ~x23 & ~x25 & ~x34 & ~x51 & ~x61 & ~x65 & ~x71 & ~x86 & ~x88 & ~x92 & ~x98 & ~x111 & ~x112 & ~x127 & ~x145 & ~x153 & ~x155 & ~x169 & ~x393 & ~x445 & ~x474 & ~x479 & ~x484 & ~x505 & ~x529 & ~x532 & ~x534 & ~x540 & ~x614 & ~x616 & ~x639 & ~x641 & ~x667 & ~x690 & ~x691 & ~x698 & ~x700 & ~x719 & ~x721 & ~x731 & ~x749 & ~x757 & ~x762 & ~x763 & ~x778 & ~x782;
assign c2151 =  x376 &  x404 & ~x1 & ~x3 & ~x15 & ~x21 & ~x32 & ~x33 & ~x39 & ~x41 & ~x48 & ~x58 & ~x70 & ~x81 & ~x83 & ~x97 & ~x108 & ~x115 & ~x117 & ~x118 & ~x136 & ~x141 & ~x164 & ~x166 & ~x168 & ~x197 & ~x201 & ~x225 & ~x251 & ~x283 & ~x284 & ~x306 & ~x310 & ~x370 & ~x396 & ~x416 & ~x422 & ~x425 & ~x426 & ~x443 & ~x454 & ~x455 & ~x456 & ~x470 & ~x472 & ~x482 & ~x500 & ~x502 & ~x508 & ~x526 & ~x527 & ~x536 & ~x556 & ~x558 & ~x561 & ~x562 & ~x563 & ~x564 & ~x585 & ~x592 & ~x609 & ~x610 & ~x613 & ~x616 & ~x619 & ~x641 & ~x642 & ~x644 & ~x669 & ~x675 & ~x678 & ~x700 & ~x705 & ~x707 & ~x709 & ~x710 & ~x715 & ~x720 & ~x723 & ~x725 & ~x728 & ~x744 & ~x745 & ~x749 & ~x751 & ~x757 & ~x758 & ~x763 & ~x767 & ~x775;
assign c2153 =  x407 & ~x15 & ~x20 & ~x27 & ~x32 & ~x49 & ~x57 & ~x64 & ~x73 & ~x83 & ~x92 & ~x104 & ~x108 & ~x110 & ~x112 & ~x137 & ~x145 & ~x164 & ~x192 & ~x222 & ~x224 & ~x282 & ~x306 & ~x316 & ~x331 & ~x333 & ~x336 & ~x340 & ~x362 & ~x365 & ~x366 & ~x367 & ~x386 & ~x387 & ~x397 & ~x416 & ~x426 & ~x427 & ~x444 & ~x446 & ~x449 & ~x454 & ~x475 & ~x476 & ~x504 & ~x505 & ~x511 & ~x513 & ~x542 & ~x544 & ~x555 & ~x556 & ~x557 & ~x558 & ~x584 & ~x587 & ~x588 & ~x611 & ~x615 & ~x616 & ~x617 & ~x618 & ~x639 & ~x669 & ~x671 & ~x674 & ~x693 & ~x715 & ~x719 & ~x720 & ~x735 & ~x745 & ~x751 & ~x752 & ~x754 & ~x755 & ~x765 & ~x773 & ~x776 & ~x781 & ~x782;
assign c2155 = ~x37 & ~x58 & ~x124 & ~x200 & ~x284 & ~x397 & ~x417 & ~x418 & ~x442 & ~x472 & ~x524 & ~x580 & ~x585 & ~x591 & ~x607 & ~x635 & ~x643 & ~x693 & ~x699 & ~x718 & ~x750 & ~x764;
assign c2157 =  x288 &  x372 &  x400 & ~x99 & ~x249;
assign c2159 =  x550 &  x660 & ~x2 & ~x47 & ~x63 & ~x69 & ~x82 & ~x93 & ~x99 & ~x111 & ~x143 & ~x384 & ~x390 & ~x392 & ~x422 & ~x447 & ~x449 & ~x474 & ~x504 & ~x527 & ~x555 & ~x582 & ~x640 & ~x666 & ~x667 & ~x675 & ~x703 & ~x708 & ~x743 & ~x762 & ~x779;
assign c2161 =  x320 &  x375 & ~x1 & ~x9 & ~x27 & ~x34 & ~x35 & ~x38 & ~x42 & ~x43 & ~x57 & ~x58 & ~x59 & ~x62 & ~x64 & ~x66 & ~x68 & ~x81 & ~x84 & ~x109 & ~x113 & ~x117 & ~x124 & ~x140 & ~x146 & ~x149 & ~x168 & ~x169 & ~x170 & ~x171 & ~x222 & ~x251 & ~x255 & ~x280 & ~x313 & ~x314 & ~x333 & ~x338 & ~x344 & ~x389 & ~x418 & ~x444 & ~x449 & ~x477 & ~x498 & ~x506 & ~x525 & ~x527 & ~x528 & ~x533 & ~x552 & ~x554 & ~x558 & ~x582 & ~x614 & ~x637 & ~x642 & ~x647 & ~x664 & ~x696 & ~x699 & ~x701 & ~x724 & ~x731 & ~x732 & ~x735 & ~x742 & ~x748 & ~x762 & ~x763 & ~x767 & ~x773;
assign c2163 = ~x1 & ~x9 & ~x10 & ~x25 & ~x30 & ~x37 & ~x44 & ~x52 & ~x57 & ~x64 & ~x65 & ~x74 & ~x79 & ~x87 & ~x94 & ~x96 & ~x97 & ~x100 & ~x101 & ~x109 & ~x120 & ~x124 & ~x142 & ~x143 & ~x156 & ~x157 & ~x224 & ~x225 & ~x251 & ~x339 & ~x362 & ~x367 & ~x419 & ~x422 & ~x451 & ~x472 & ~x474 & ~x478 & ~x500 & ~x528 & ~x537 & ~x538 & ~x550 & ~x555 & ~x562 & ~x577 & ~x588 & ~x589 & ~x591 & ~x604 & ~x605 & ~x615 & ~x634 & ~x640 & ~x674 & ~x689 & ~x715 & ~x731 & ~x753 & ~x756 & ~x762 & ~x771 & ~x783;
assign c2165 = ~x2 & ~x5 & ~x8 & ~x11 & ~x19 & ~x20 & ~x21 & ~x22 & ~x26 & ~x36 & ~x41 & ~x42 & ~x52 & ~x53 & ~x54 & ~x59 & ~x60 & ~x62 & ~x64 & ~x65 & ~x68 & ~x69 & ~x77 & ~x78 & ~x80 & ~x81 & ~x86 & ~x91 & ~x93 & ~x95 & ~x96 & ~x100 & ~x111 & ~x113 & ~x123 & ~x132 & ~x135 & ~x140 & ~x142 & ~x144 & ~x145 & ~x159 & ~x162 & ~x164 & ~x167 & ~x189 & ~x191 & ~x193 & ~x194 & ~x195 & ~x198 & ~x220 & ~x225 & ~x250 & ~x279 & ~x309 & ~x335 & ~x337 & ~x338 & ~x363 & ~x364 & ~x365 & ~x366 & ~x370 & ~x387 & ~x388 & ~x390 & ~x391 & ~x396 & ~x418 & ~x420 & ~x424 & ~x444 & ~x445 & ~x446 & ~x471 & ~x478 & ~x497 & ~x499 & ~x500 & ~x501 & ~x506 & ~x525 & ~x526 & ~x528 & ~x535 & ~x537 & ~x539 & ~x540 & ~x553 & ~x557 & ~x559 & ~x560 & ~x562 & ~x563 & ~x568 & ~x569 & ~x580 & ~x581 & ~x586 & ~x587 & ~x589 & ~x592 & ~x595 & ~x609 & ~x610 & ~x611 & ~x618 & ~x623 & ~x636 & ~x637 & ~x640 & ~x642 & ~x647 & ~x649 & ~x651 & ~x667 & ~x668 & ~x670 & ~x671 & ~x672 & ~x691 & ~x693 & ~x694 & ~x696 & ~x698 & ~x701 & ~x702 & ~x719 & ~x720 & ~x727 & ~x731 & ~x745 & ~x747 & ~x749 & ~x752 & ~x753 & ~x755 & ~x757 & ~x758 & ~x765 & ~x766 & ~x777 & ~x782;
assign c2167 =  x371 &  x427 & ~x375 & ~x751;
assign c2169 =  x600 & ~x66 & ~x123 & ~x181 & ~x209 & ~x314 & ~x390 & ~x479 & ~x582 & ~x586 & ~x647 & ~x699 & ~x720 & ~x722 & ~x758 & ~x769;
assign c2171 =  x402 & ~x0 & ~x6 & ~x7 & ~x10 & ~x12 & ~x32 & ~x38 & ~x52 & ~x54 & ~x56 & ~x62 & ~x66 & ~x73 & ~x74 & ~x77 & ~x83 & ~x92 & ~x101 & ~x110 & ~x115 & ~x116 & ~x119 & ~x166 & ~x170 & ~x223 & ~x226 & ~x253 & ~x278 & ~x335 & ~x361 & ~x417 & ~x419 & ~x445 & ~x450 & ~x471 & ~x476 & ~x480 & ~x482 & ~x500 & ~x509 & ~x511 & ~x513 & ~x538 & ~x556 & ~x558 & ~x560 & ~x612 & ~x613 & ~x679 & ~x694 & ~x702 & ~x704 & ~x706 & ~x707 & ~x723 & ~x725 & ~x726 & ~x727 & ~x729 & ~x732 & ~x733 & ~x734 & ~x739 & ~x743 & ~x745 & ~x750 & ~x752 & ~x762 & ~x763 & ~x766 & ~x771 & ~x772 & ~x773 & ~x776;
assign c2173 =  x341;
assign c2175 =  x494 & ~x1 & ~x23 & ~x26 & ~x36 & ~x39 & ~x80 & ~x81 & ~x92 & ~x106 & ~x114 & ~x119 & ~x136 & ~x138 & ~x147 & ~x152 & ~x219 & ~x279 & ~x307 & ~x309 & ~x332 & ~x336 & ~x360 & ~x363 & ~x390 & ~x415 & ~x420 & ~x444 & ~x445 & ~x447 & ~x477 & ~x478 & ~x500 & ~x509 & ~x510 & ~x526 & ~x527 & ~x531 & ~x532 & ~x534 & ~x538 & ~x561 & ~x562 & ~x568 & ~x584 & ~x587 & ~x593 & ~x594 & ~x618 & ~x621 & ~x624 & ~x642 & ~x648 & ~x650 & ~x670 & ~x672 & ~x697 & ~x698 & ~x725 & ~x750 & ~x777 & ~x778 & ~x781;
assign c2177 =  x373 &  x400 &  x428 & ~x13 & ~x27 & ~x49 & ~x83 & ~x118 & ~x193 & ~x201 & ~x377 & ~x590 & ~x610 & ~x665 & ~x695 & ~x702 & ~x713 & ~x723 & ~x760;
assign c2179 = ~x1 & ~x3 & ~x5 & ~x9 & ~x12 & ~x14 & ~x17 & ~x18 & ~x23 & ~x24 & ~x25 & ~x27 & ~x29 & ~x30 & ~x33 & ~x38 & ~x39 & ~x41 & ~x42 & ~x43 & ~x45 & ~x49 & ~x50 & ~x51 & ~x52 & ~x54 & ~x55 & ~x60 & ~x61 & ~x63 & ~x65 & ~x66 & ~x68 & ~x69 & ~x82 & ~x83 & ~x84 & ~x87 & ~x92 & ~x93 & ~x107 & ~x108 & ~x109 & ~x111 & ~x113 & ~x116 & ~x137 & ~x138 & ~x139 & ~x165 & ~x167 & ~x170 & ~x171 & ~x192 & ~x194 & ~x198 & ~x221 & ~x222 & ~x225 & ~x252 & ~x254 & ~x277 & ~x279 & ~x280 & ~x281 & ~x305 & ~x306 & ~x307 & ~x309 & ~x310 & ~x334 & ~x337 & ~x338 & ~x362 & ~x365 & ~x371 & ~x389 & ~x391 & ~x399 & ~x419 & ~x421 & ~x423 & ~x428 & ~x445 & ~x456 & ~x458 & ~x472 & ~x477 & ~x478 & ~x486 & ~x501 & ~x502 & ~x503 & ~x506 & ~x515 & ~x516 & ~x517 & ~x530 & ~x531 & ~x533 & ~x534 & ~x545 & ~x556 & ~x559 & ~x560 & ~x561 & ~x562 & ~x587 & ~x588 & ~x611 & ~x613 & ~x615 & ~x616 & ~x617 & ~x618 & ~x639 & ~x642 & ~x644 & ~x647 & ~x666 & ~x668 & ~x671 & ~x673 & ~x674 & ~x680 & ~x701 & ~x703 & ~x705 & ~x708 & ~x711 & ~x712 & ~x715 & ~x720 & ~x722 & ~x724 & ~x727 & ~x728 & ~x731 & ~x732 & ~x733 & ~x734 & ~x736 & ~x738 & ~x740 & ~x748 & ~x751 & ~x752 & ~x753 & ~x756 & ~x760 & ~x761 & ~x762 & ~x763 & ~x767 & ~x768 & ~x776 & ~x779 & ~x781 & ~x783;
assign c2181 = ~x1 & ~x6 & ~x13 & ~x14 & ~x15 & ~x19 & ~x21 & ~x24 & ~x25 & ~x33 & ~x36 & ~x37 & ~x39 & ~x44 & ~x46 & ~x47 & ~x50 & ~x53 & ~x60 & ~x63 & ~x71 & ~x72 & ~x76 & ~x80 & ~x85 & ~x87 & ~x93 & ~x95 & ~x99 & ~x104 & ~x107 & ~x109 & ~x115 & ~x121 & ~x132 & ~x134 & ~x144 & ~x160 & ~x162 & ~x164 & ~x166 & ~x173 & ~x196 & ~x220 & ~x221 & ~x224 & ~x225 & ~x247 & ~x278 & ~x280 & ~x304 & ~x308 & ~x337 & ~x360 & ~x365 & ~x389 & ~x390 & ~x392 & ~x418 & ~x445 & ~x451 & ~x472 & ~x478 & ~x499 & ~x501 & ~x503 & ~x506 & ~x511 & ~x527 & ~x528 & ~x538 & ~x539 & ~x543 & ~x569 & ~x570 & ~x571 & ~x583 & ~x585 & ~x588 & ~x590 & ~x596 & ~x599 & ~x600 & ~x614 & ~x640 & ~x643 & ~x670 & ~x671 & ~x673 & ~x696 & ~x700 & ~x703 & ~x704 & ~x705 & ~x708 & ~x725 & ~x727 & ~x734 & ~x735 & ~x736 & ~x753 & ~x762 & ~x763 & ~x767 & ~x769 & ~x775 & ~x777;
assign c2183 = ~x5 & ~x22 & ~x23 & ~x45 & ~x46 & ~x54 & ~x84 & ~x89 & ~x111 & ~x121 & ~x144 & ~x156 & ~x359 & ~x387 & ~x389 & ~x390 & ~x444 & ~x448 & ~x449 & ~x455 & ~x472 & ~x499 & ~x508 & ~x509 & ~x528 & ~x529 & ~x554 & ~x555 & ~x561 & ~x565 & ~x566 & ~x570 & ~x583 & ~x590 & ~x596 & ~x608 & ~x610 & ~x614 & ~x619 & ~x663 & ~x666 & ~x690 & ~x691 & ~x718 & ~x734 & ~x747 & ~x751 & ~x768 & ~x781;
assign c2185 =  x382 & ~x4 & ~x12 & ~x64 & ~x82 & ~x105 & ~x144 & ~x182 & ~x195 & ~x223 & ~x331 & ~x420 & ~x565 & ~x567 & ~x570 & ~x587 & ~x588 & ~x650 & ~x766;
assign c2187 = ~x23 & ~x52 & ~x71 & ~x125 & ~x180 & ~x207 & ~x248 & ~x263 & ~x361 & ~x390 & ~x446 & ~x492 & ~x613 & ~x659;
assign c2189 =  x660 & ~x0 & ~x1 & ~x4 & ~x5 & ~x10 & ~x14 & ~x15 & ~x18 & ~x24 & ~x27 & ~x32 & ~x33 & ~x34 & ~x36 & ~x38 & ~x41 & ~x42 & ~x45 & ~x48 & ~x50 & ~x60 & ~x70 & ~x84 & ~x86 & ~x92 & ~x93 & ~x97 & ~x101 & ~x103 & ~x104 & ~x111 & ~x112 & ~x117 & ~x118 & ~x146 & ~x167 & ~x168 & ~x223 & ~x225 & ~x251 & ~x275 & ~x278 & ~x279 & ~x282 & ~x305 & ~x307 & ~x308 & ~x331 & ~x334 & ~x335 & ~x361 & ~x366 & ~x390 & ~x392 & ~x417 & ~x418 & ~x419 & ~x420 & ~x421 & ~x446 & ~x478 & ~x480 & ~x502 & ~x503 & ~x515 & ~x532 & ~x544 & ~x558 & ~x573 & ~x612 & ~x615 & ~x616 & ~x619 & ~x643 & ~x666 & ~x667 & ~x668 & ~x671 & ~x695 & ~x697 & ~x701 & ~x704 & ~x707 & ~x708 & ~x720 & ~x721 & ~x732 & ~x733 & ~x736 & ~x738 & ~x749 & ~x769 & ~x774 & ~x777 & ~x778 & ~x781 & ~x782 & ~x783;
assign c2191 =  x430 & ~x19 & ~x38 & ~x135 & ~x193 & ~x223 & ~x350 & ~x377 & ~x444 & ~x509 & ~x555 & ~x568 & ~x592 & ~x642 & ~x705 & ~x722;
assign c2193 =  x290 &  x345 &  x373 &  x401 & ~x13 & ~x198 & ~x333 & ~x502 & ~x529 & ~x645 & ~x751;
assign c2195 =  x319 &  x347 &  x374 &  x402 & ~x11 & ~x12 & ~x51 & ~x55 & ~x56 & ~x64 & ~x85 & ~x90 & ~x108 & ~x167 & ~x170 & ~x203 & ~x205 & ~x223 & ~x252 & ~x255 & ~x339 & ~x423 & ~x445 & ~x448 & ~x474 & ~x479 & ~x504 & ~x533 & ~x554 & ~x563 & ~x582 & ~x613 & ~x663 & ~x671 & ~x691 & ~x698 & ~x716 & ~x721 & ~x760 & ~x767 & ~x774 & ~x775 & ~x779 & ~x781;
assign c2197 = ~x1 & ~x2 & ~x7 & ~x33 & ~x34 & ~x51 & ~x57 & ~x64 & ~x71 & ~x73 & ~x81 & ~x84 & ~x85 & ~x88 & ~x108 & ~x109 & ~x110 & ~x138 & ~x167 & ~x195 & ~x196 & ~x197 & ~x203 & ~x226 & ~x232 & ~x279 & ~x280 & ~x282 & ~x335 & ~x366 & ~x367 & ~x394 & ~x396 & ~x444 & ~x460 & ~x463 & ~x486 & ~x487 & ~x490 & ~x491 & ~x531 & ~x556 & ~x610 & ~x612 & ~x613 & ~x615 & ~x666 & ~x690 & ~x693 & ~x699 & ~x709 & ~x711 & ~x719 & ~x721 & ~x722 & ~x735 & ~x736 & ~x751 & ~x758 & ~x763 & ~x764 & ~x766 & ~x774;
assign c2199 =  x404 &  x407 &  x433 & ~x1 & ~x3 & ~x7 & ~x11 & ~x12 & ~x22 & ~x26 & ~x32 & ~x38 & ~x42 & ~x50 & ~x61 & ~x66 & ~x67 & ~x77 & ~x81 & ~x83 & ~x87 & ~x94 & ~x107 & ~x108 & ~x110 & ~x136 & ~x138 & ~x139 & ~x140 & ~x142 & ~x143 & ~x170 & ~x172 & ~x221 & ~x225 & ~x226 & ~x251 & ~x268 & ~x283 & ~x390 & ~x391 & ~x416 & ~x423 & ~x425 & ~x444 & ~x472 & ~x473 & ~x481 & ~x482 & ~x499 & ~x503 & ~x504 & ~x510 & ~x511 & ~x556 & ~x586 & ~x611 & ~x613 & ~x617 & ~x639 & ~x698 & ~x699 & ~x705 & ~x721 & ~x723 & ~x729 & ~x735 & ~x742 & ~x749 & ~x756 & ~x764 & ~x770 & ~x780 & ~x781;
assign c2201 = ~x47 & ~x49 & ~x124 & ~x141 & ~x204 & ~x229 & ~x263 & ~x285 & ~x286 & ~x358 & ~x415 & ~x551 & ~x577 & ~x587 & ~x589 & ~x631 & ~x661 & ~x783;
assign c2203 =  x292 &  x347 &  x374 &  x402 & ~x49 & ~x50 & ~x63 & ~x68 & ~x108 & ~x111 & ~x113 & ~x121 & ~x149 & ~x175 & ~x195 & ~x204 & ~x226 & ~x228 & ~x308 & ~x333 & ~x337 & ~x366 & ~x368 & ~x392 & ~x395 & ~x396 & ~x447 & ~x527 & ~x529 & ~x590 & ~x610 & ~x611 & ~x612 & ~x619 & ~x638 & ~x667 & ~x668 & ~x677 & ~x678 & ~x679 & ~x696 & ~x749 & ~x758;
assign c2205 =  x406 & ~x149 & ~x440 & ~x577 & ~x605 & ~x632 & ~x714;
assign c2207 =  x604 & ~x2 & ~x8 & ~x12 & ~x29 & ~x51 & ~x56 & ~x66 & ~x68 & ~x82 & ~x84 & ~x94 & ~x134 & ~x138 & ~x200 & ~x251 & ~x385 & ~x413 & ~x425 & ~x427 & ~x440 & ~x452 & ~x455 & ~x509 & ~x544 & ~x555 & ~x564 & ~x581 & ~x587 & ~x609 & ~x636 & ~x663 & ~x670 & ~x694 & ~x719 & ~x746 & ~x757 & ~x771 & ~x779;
assign c2209 =  x405 & ~x7 & ~x51 & ~x101 & ~x105 & ~x115 & ~x139 & ~x196 & ~x312 & ~x360 & ~x373 & ~x387 & ~x401 & ~x413 & ~x440 & ~x445 & ~x455 & ~x468 & ~x469 & ~x470 & ~x471 & ~x474 & ~x495 & ~x498 & ~x505 & ~x523 & ~x524 & ~x529 & ~x551 & ~x560 & ~x581 & ~x606 & ~x613 & ~x634 & ~x638 & ~x662 & ~x690 & ~x752 & ~x778;
assign c2211 =  x317 &  x345 & ~x13 & ~x32 & ~x34 & ~x77 & ~x78 & ~x82 & ~x131 & ~x135 & ~x140 & ~x256 & ~x342 & ~x370 & ~x389 & ~x446 & ~x501 & ~x503 & ~x528 & ~x643 & ~x648 & ~x653 & ~x664 & ~x668 & ~x695 & ~x710 & ~x713 & ~x743 & ~x756 & ~x781;
assign c2213 =  x317 &  x345 &  x400 & ~x31 & ~x108 & ~x677;
assign c2215 =  x344 &  x372 & ~x2 & ~x25 & ~x69 & ~x299 & ~x361 & ~x615 & ~x619 & ~x772 & ~x778;
assign c2217 = ~x0 & ~x3 & ~x22 & ~x32 & ~x40 & ~x42 & ~x47 & ~x49 & ~x53 & ~x59 & ~x60 & ~x62 & ~x65 & ~x70 & ~x77 & ~x79 & ~x85 & ~x91 & ~x102 & ~x104 & ~x105 & ~x107 & ~x110 & ~x112 & ~x118 & ~x120 & ~x121 & ~x129 & ~x133 & ~x134 & ~x135 & ~x160 & ~x161 & ~x163 & ~x167 & ~x188 & ~x189 & ~x192 & ~x195 & ~x222 & ~x223 & ~x249 & ~x305 & ~x332 & ~x364 & ~x365 & ~x388 & ~x389 & ~x416 & ~x422 & ~x423 & ~x444 & ~x450 & ~x473 & ~x474 & ~x479 & ~x502 & ~x517 & ~x518 & ~x529 & ~x530 & ~x539 & ~x545 & ~x546 & ~x556 & ~x562 & ~x573 & ~x574 & ~x595 & ~x614 & ~x617 & ~x619 & ~x620 & ~x623 & ~x641 & ~x647 & ~x674 & ~x676 & ~x696 & ~x700 & ~x705 & ~x728 & ~x732 & ~x734 & ~x753 & ~x757 & ~x760 & ~x770 & ~x780;
assign c2219 =  x344 &  x428 & ~x281 & ~x449 & ~x474 & ~x610 & ~x762 & ~x776;
assign c2221 = ~x3 & ~x6 & ~x12 & ~x21 & ~x28 & ~x45 & ~x52 & ~x60 & ~x64 & ~x69 & ~x80 & ~x84 & ~x106 & ~x140 & ~x151 & ~x158 & ~x161 & ~x220 & ~x223 & ~x304 & ~x305 & ~x306 & ~x319 & ~x392 & ~x415 & ~x418 & ~x422 & ~x444 & ~x475 & ~x479 & ~x498 & ~x506 & ~x527 & ~x531 & ~x535 & ~x555 & ~x568 & ~x597 & ~x599 & ~x610 & ~x678 & ~x707 & ~x723 & ~x757 & ~x762 & ~x768;
assign c2223 =  x598 &  x599 & ~x0 & ~x3 & ~x5 & ~x8 & ~x15 & ~x22 & ~x23 & ~x26 & ~x27 & ~x33 & ~x36 & ~x44 & ~x52 & ~x55 & ~x60 & ~x62 & ~x64 & ~x80 & ~x83 & ~x84 & ~x85 & ~x86 & ~x89 & ~x90 & ~x91 & ~x92 & ~x93 & ~x97 & ~x99 & ~x100 & ~x109 & ~x120 & ~x167 & ~x196 & ~x201 & ~x202 & ~x203 & ~x225 & ~x227 & ~x230 & ~x251 & ~x255 & ~x258 & ~x259 & ~x279 & ~x283 & ~x286 & ~x287 & ~x308 & ~x312 & ~x333 & ~x334 & ~x342 & ~x357 & ~x359 & ~x367 & ~x369 & ~x370 & ~x371 & ~x386 & ~x390 & ~x394 & ~x398 & ~x414 & ~x415 & ~x416 & ~x417 & ~x419 & ~x427 & ~x428 & ~x441 & ~x442 & ~x448 & ~x449 & ~x450 & ~x456 & ~x469 & ~x470 & ~x475 & ~x476 & ~x497 & ~x498 & ~x500 & ~x502 & ~x504 & ~x527 & ~x529 & ~x532 & ~x552 & ~x553 & ~x554 & ~x555 & ~x556 & ~x560 & ~x582 & ~x587 & ~x607 & ~x608 & ~x611 & ~x617 & ~x635 & ~x640 & ~x642 & ~x643 & ~x645 & ~x646 & ~x663 & ~x664 & ~x666 & ~x671 & ~x672 & ~x676 & ~x689 & ~x692 & ~x697 & ~x700 & ~x704 & ~x712 & ~x714 & ~x715 & ~x717 & ~x718 & ~x719 & ~x720 & ~x724 & ~x729 & ~x738 & ~x740 & ~x743 & ~x744 & ~x749 & ~x751 & ~x755 & ~x758 & ~x762 & ~x766 & ~x769 & ~x770 & ~x772 & ~x779 & ~x783;
assign c2225 = ~x16 & ~x19 & ~x20 & ~x29 & ~x51 & ~x52 & ~x68 & ~x95 & ~x111 & ~x113 & ~x118 & ~x122 & ~x140 & ~x147 & ~x148 & ~x228 & ~x257 & ~x278 & ~x279 & ~x309 & ~x310 & ~x360 & ~x389 & ~x390 & ~x467 & ~x495 & ~x501 & ~x514 & ~x524 & ~x556 & ~x563 & ~x578 & ~x579 & ~x580 & ~x609 & ~x614 & ~x633 & ~x636 & ~x662 & ~x665 & ~x669 & ~x676 & ~x730 & ~x732 & ~x733 & ~x752 & ~x760 & ~x777 & ~x778;
assign c2227 =  x324 &  x551 &  x578 & ~x1 & ~x8 & ~x14 & ~x46 & ~x48 & ~x52 & ~x61 & ~x66 & ~x73 & ~x86 & ~x108 & ~x113 & ~x116 & ~x138 & ~x161 & ~x163 & ~x194 & ~x308 & ~x421 & ~x473 & ~x474 & ~x475 & ~x504 & ~x516 & ~x517 & ~x528 & ~x555 & ~x582 & ~x583 & ~x586 & ~x591 & ~x638 & ~x642 & ~x668 & ~x694 & ~x726 & ~x729 & ~x733 & ~x749 & ~x758 & ~x770 & ~x772 & ~x778;
assign c2229 =  x347 &  x375 &  x404 &  x407 & ~x5 & ~x52 & ~x59 & ~x67 & ~x117 & ~x165 & ~x399 & ~x419 & ~x427 & ~x471 & ~x480 & ~x528 & ~x589 & ~x612 & ~x674 & ~x744 & ~x745;
assign c2231 = ~x38 & ~x44 & ~x89 & ~x137 & ~x139 & ~x240 & ~x254 & ~x268 & ~x295 & ~x390 & ~x418 & ~x443 & ~x448 & ~x449 & ~x499 & ~x509 & ~x528 & ~x539 & ~x558 & ~x560 & ~x568 & ~x597 & ~x688;
assign c2233 =  x375 &  x404 &  x658 &  x659 & ~x3 & ~x9 & ~x10 & ~x18 & ~x25 & ~x49 & ~x57 & ~x61 & ~x142 & ~x224 & ~x362 & ~x450 & ~x475 & ~x506 & ~x508 & ~x533 & ~x561 & ~x592 & ~x644 & ~x675 & ~x699 & ~x720 & ~x728;
assign c2235 =  x232 &  x437 & ~x23 & ~x34 & ~x39 & ~x43 & ~x54 & ~x96 & ~x127 & ~x197 & ~x308 & ~x309 & ~x415 & ~x418 & ~x421 & ~x443 & ~x475 & ~x506 & ~x537 & ~x564 & ~x572 & ~x593 & ~x616 & ~x704 & ~x736 & ~x751 & ~x783;
assign c2237 = ~x10 & ~x12 & ~x17 & ~x19 & ~x23 & ~x34 & ~x38 & ~x39 & ~x43 & ~x50 & ~x53 & ~x60 & ~x62 & ~x66 & ~x83 & ~x84 & ~x85 & ~x86 & ~x92 & ~x93 & ~x94 & ~x97 & ~x123 & ~x124 & ~x143 & ~x145 & ~x171 & ~x176 & ~x197 & ~x220 & ~x226 & ~x227 & ~x253 & ~x255 & ~x270 & ~x277 & ~x279 & ~x283 & ~x297 & ~x303 & ~x309 & ~x312 & ~x335 & ~x336 & ~x338 & ~x362 & ~x366 & ~x387 & ~x395 & ~x415 & ~x416 & ~x419 & ~x422 & ~x426 & ~x454 & ~x471 & ~x498 & ~x502 & ~x505 & ~x507 & ~x510 & ~x525 & ~x527 & ~x531 & ~x536 & ~x537 & ~x538 & ~x558 & ~x562 & ~x581 & ~x584 & ~x586 & ~x587 & ~x588 & ~x589 & ~x591 & ~x593 & ~x608 & ~x610 & ~x615 & ~x636 & ~x638 & ~x644 & ~x650 & ~x663 & ~x665 & ~x667 & ~x671 & ~x674 & ~x675 & ~x678 & ~x691 & ~x696 & ~x712 & ~x722 & ~x726 & ~x729 & ~x731 & ~x732 & ~x733 & ~x737 & ~x738 & ~x739 & ~x749 & ~x754 & ~x769 & ~x770 & ~x773 & ~x775 & ~x776 & ~x777;
assign c2239 = ~x4 & ~x16 & ~x47 & ~x50 & ~x53 & ~x65 & ~x68 & ~x76 & ~x77 & ~x90 & ~x97 & ~x139 & ~x166 & ~x167 & ~x195 & ~x256 & ~x309 & ~x331 & ~x362 & ~x373 & ~x388 & ~x412 & ~x444 & ~x468 & ~x473 & ~x477 & ~x496 & ~x497 & ~x498 & ~x522 & ~x523 & ~x528 & ~x529 & ~x533 & ~x534 & ~x551 & ~x552 & ~x554 & ~x556 & ~x557 & ~x578 & ~x584 & ~x588 & ~x616 & ~x618 & ~x619 & ~x634 & ~x635 & ~x637 & ~x648 & ~x662 & ~x663 & ~x665 & ~x689 & ~x691 & ~x696 & ~x697 & ~x716 & ~x718 & ~x731 & ~x754 & ~x755 & ~x776 & ~x782;
assign c2241 =  x519 & ~x21 & ~x30 & ~x35 & ~x66 & ~x80 & ~x81 & ~x90 & ~x99 & ~x101 & ~x114 & ~x120 & ~x137 & ~x138 & ~x140 & ~x153 & ~x155 & ~x156 & ~x165 & ~x250 & ~x251 & ~x284 & ~x392 & ~x480 & ~x499 & ~x502 & ~x527 & ~x535 & ~x581 & ~x609 & ~x612 & ~x638 & ~x648 & ~x692 & ~x719 & ~x720 & ~x726 & ~x733 & ~x774 & ~x778 & ~x780 & ~x781;
assign c2243 =  x435 &  x658 &  x686 & ~x52 & ~x93 & ~x162;
assign c2245 =  x464 &  x493 & ~x2 & ~x3 & ~x9 & ~x12 & ~x14 & ~x17 & ~x20 & ~x22 & ~x24 & ~x26 & ~x28 & ~x29 & ~x31 & ~x32 & ~x35 & ~x39 & ~x42 & ~x43 & ~x47 & ~x55 & ~x59 & ~x60 & ~x62 & ~x64 & ~x65 & ~x68 & ~x69 & ~x72 & ~x74 & ~x75 & ~x76 & ~x78 & ~x84 & ~x87 & ~x94 & ~x95 & ~x99 & ~x100 & ~x107 & ~x108 & ~x110 & ~x113 & ~x115 & ~x116 & ~x119 & ~x122 & ~x130 & ~x133 & ~x138 & ~x140 & ~x163 & ~x166 & ~x168 & ~x169 & ~x223 & ~x249 & ~x252 & ~x275 & ~x308 & ~x333 & ~x360 & ~x365 & ~x387 & ~x388 & ~x392 & ~x413 & ~x417 & ~x442 & ~x445 & ~x479 & ~x499 & ~x500 & ~x506 & ~x509 & ~x536 & ~x537 & ~x556 & ~x562 & ~x584 & ~x589 & ~x593 & ~x599 & ~x617 & ~x620 & ~x622 & ~x643 & ~x671 & ~x698 & ~x699 & ~x700 & ~x701 & ~x724 & ~x728 & ~x730 & ~x731 & ~x732 & ~x738 & ~x754 & ~x761 & ~x762 & ~x774 & ~x780 & ~x781 & ~x782;
assign c2247 =  x454 & ~x9 & ~x17 & ~x22 & ~x44 & ~x109 & ~x138 & ~x145 & ~x221 & ~x278 & ~x366 & ~x405 & ~x406 & ~x430 & ~x475 & ~x477 & ~x501 & ~x646 & ~x667 & ~x728 & ~x773;
assign c2249 =  x710;
assign c2251 =  x375 &  x403 & ~x25 & ~x29 & ~x31 & ~x45 & ~x149 & ~x165 & ~x169 & ~x196 & ~x286 & ~x307 & ~x334 & ~x339 & ~x340 & ~x342 & ~x393 & ~x398 & ~x427 & ~x446 & ~x449 & ~x497 & ~x500 & ~x503 & ~x525 & ~x531 & ~x581 & ~x635 & ~x636 & ~x649 & ~x662 & ~x665 & ~x672 & ~x689 & ~x694 & ~x701 & ~x702 & ~x719 & ~x744 & ~x755 & ~x769 & ~x776 & ~x783;
assign c2253 =  x377 & ~x1 & ~x3 & ~x5 & ~x8 & ~x10 & ~x11 & ~x14 & ~x17 & ~x18 & ~x19 & ~x20 & ~x21 & ~x22 & ~x23 & ~x25 & ~x28 & ~x30 & ~x34 & ~x35 & ~x36 & ~x39 & ~x41 & ~x43 & ~x44 & ~x48 & ~x50 & ~x51 & ~x53 & ~x58 & ~x59 & ~x65 & ~x66 & ~x67 & ~x71 & ~x72 & ~x75 & ~x76 & ~x78 & ~x80 & ~x81 & ~x84 & ~x85 & ~x87 & ~x88 & ~x92 & ~x93 & ~x97 & ~x100 & ~x108 & ~x109 & ~x110 & ~x113 & ~x114 & ~x118 & ~x120 & ~x121 & ~x135 & ~x137 & ~x138 & ~x139 & ~x143 & ~x163 & ~x170 & ~x191 & ~x193 & ~x198 & ~x222 & ~x224 & ~x228 & ~x251 & ~x253 & ~x254 & ~x255 & ~x282 & ~x283 & ~x284 & ~x310 & ~x312 & ~x313 & ~x314 & ~x332 & ~x335 & ~x337 & ~x341 & ~x358 & ~x359 & ~x361 & ~x363 & ~x365 & ~x367 & ~x368 & ~x369 & ~x370 & ~x387 & ~x390 & ~x391 & ~x393 & ~x397 & ~x399 & ~x414 & ~x415 & ~x416 & ~x417 & ~x419 & ~x421 & ~x422 & ~x423 & ~x425 & ~x426 & ~x427 & ~x443 & ~x444 & ~x449 & ~x454 & ~x455 & ~x456 & ~x457 & ~x472 & ~x473 & ~x474 & ~x475 & ~x477 & ~x478 & ~x479 & ~x484 & ~x498 & ~x499 & ~x500 & ~x501 & ~x503 & ~x504 & ~x506 & ~x527 & ~x528 & ~x529 & ~x530 & ~x534 & ~x554 & ~x555 & ~x559 & ~x562 & ~x582 & ~x583 & ~x586 & ~x588 & ~x611 & ~x612 & ~x614 & ~x617 & ~x642 & ~x643 & ~x644 & ~x646 & ~x665 & ~x672 & ~x692 & ~x694 & ~x695 & ~x696 & ~x699 & ~x700 & ~x704 & ~x705 & ~x707 & ~x708 & ~x709 & ~x712 & ~x714 & ~x715 & ~x717 & ~x719 & ~x721 & ~x722 & ~x724 & ~x728 & ~x731 & ~x732 & ~x734 & ~x738 & ~x739 & ~x740 & ~x742 & ~x745 & ~x746 & ~x749 & ~x754 & ~x757 & ~x759 & ~x761 & ~x762 & ~x766 & ~x767 & ~x770 & ~x773 & ~x774 & ~x775 & ~x778 & ~x779 & ~x780;
assign c2255 = ~x1 & ~x3 & ~x17 & ~x19 & ~x29 & ~x53 & ~x83 & ~x86 & ~x111 & ~x140 & ~x146 & ~x147 & ~x166 & ~x221 & ~x299 & ~x325 & ~x328 & ~x332 & ~x352 & ~x359 & ~x369 & ~x390 & ~x413 & ~x414 & ~x442 & ~x448 & ~x480 & ~x508 & ~x526 & ~x531 & ~x536 & ~x583 & ~x589 & ~x616 & ~x621 & ~x638 & ~x639 & ~x675 & ~x693 & ~x712 & ~x737 & ~x740 & ~x747 & ~x756;
assign c2257 =  x321 &  x349 & ~x0 & ~x3 & ~x12 & ~x16 & ~x17 & ~x18 & ~x29 & ~x33 & ~x35 & ~x37 & ~x45 & ~x47 & ~x48 & ~x49 & ~x58 & ~x59 & ~x71 & ~x86 & ~x89 & ~x91 & ~x92 & ~x113 & ~x114 & ~x120 & ~x137 & ~x148 & ~x167 & ~x168 & ~x170 & ~x173 & ~x176 & ~x196 & ~x197 & ~x202 & ~x203 & ~x230 & ~x231 & ~x233 & ~x250 & ~x260 & ~x261 & ~x277 & ~x280 & ~x281 & ~x285 & ~x289 & ~x310 & ~x315 & ~x317 & ~x334 & ~x342 & ~x361 & ~x363 & ~x365 & ~x390 & ~x391 & ~x393 & ~x395 & ~x422 & ~x423 & ~x443 & ~x445 & ~x448 & ~x449 & ~x450 & ~x471 & ~x477 & ~x497 & ~x498 & ~x500 & ~x501 & ~x508 & ~x531 & ~x554 & ~x555 & ~x559 & ~x580 & ~x589 & ~x615 & ~x636 & ~x643 & ~x647 & ~x664 & ~x666 & ~x672 & ~x674 & ~x676 & ~x679 & ~x688 & ~x699 & ~x702 & ~x704 & ~x715 & ~x719 & ~x725 & ~x732 & ~x733 & ~x747 & ~x751 & ~x753 & ~x758 & ~x759 & ~x765 & ~x766 & ~x771 & ~x772;
assign c2259 =  x317 & ~x158 & ~x240 & ~x268 & ~x312 & ~x620 & ~x621 & ~x701;
assign c2261 =  x651 & ~x156 & ~x468 & ~x633;
assign c2263 = ~x0 & ~x1 & ~x2 & ~x6 & ~x10 & ~x16 & ~x17 & ~x19 & ~x20 & ~x33 & ~x38 & ~x41 & ~x42 & ~x44 & ~x45 & ~x46 & ~x49 & ~x59 & ~x68 & ~x87 & ~x96 & ~x101 & ~x111 & ~x117 & ~x120 & ~x123 & ~x127 & ~x154 & ~x155 & ~x158 & ~x159 & ~x174 & ~x194 & ~x195 & ~x200 & ~x223 & ~x225 & ~x255 & ~x309 & ~x312 & ~x338 & ~x360 & ~x387 & ~x415 & ~x417 & ~x422 & ~x444 & ~x445 & ~x473 & ~x478 & ~x498 & ~x499 & ~x501 & ~x506 & ~x528 & ~x529 & ~x531 & ~x536 & ~x554 & ~x557 & ~x560 & ~x563 & ~x584 & ~x586 & ~x588 & ~x590 & ~x591 & ~x618 & ~x619 & ~x634 & ~x638 & ~x639 & ~x640 & ~x646 & ~x667 & ~x701 & ~x704 & ~x715 & ~x718 & ~x719 & ~x720 & ~x724 & ~x731 & ~x732 & ~x746 & ~x747 & ~x753 & ~x755 & ~x758 & ~x772 & ~x776 & ~x783;
assign c2265 =  x348 &  x630 &  x631 &  x632 & ~x426 & ~x427 & ~x455 & ~x476 & ~x482;
assign c2267 =  x314 &  x426 & ~x11 & ~x31 & ~x109 & ~x474 & ~x535 & ~x699 & ~x712 & ~x750;
assign c2269 =  x682 & ~x543;
assign c2271 =  x357 & ~x34 & ~x336 & ~x537 & ~x626;
assign c2273 =  x292 &  x347 &  x573 & ~x10 & ~x22 & ~x50 & ~x59 & ~x63 & ~x70 & ~x85 & ~x86 & ~x114 & ~x145 & ~x149 & ~x173 & ~x228 & ~x259 & ~x287 & ~x363 & ~x418 & ~x422 & ~x582 & ~x589 & ~x607 & ~x609 & ~x610 & ~x641 & ~x659 & ~x663 & ~x674 & ~x684 & ~x710 & ~x712 & ~x749 & ~x768;
assign c2275 =  x269 &  x296 & ~x9 & ~x20 & ~x26 & ~x59 & ~x77 & ~x93 & ~x101 & ~x139 & ~x153 & ~x197 & ~x391 & ~x415 & ~x447 & ~x470 & ~x471 & ~x498 & ~x535 & ~x555 & ~x602 & ~x648 & ~x765 & ~x768;
assign c2277 =  x271 & ~x0 & ~x5 & ~x7 & ~x9 & ~x19 & ~x20 & ~x25 & ~x31 & ~x47 & ~x49 & ~x54 & ~x63 & ~x65 & ~x69 & ~x71 & ~x77 & ~x85 & ~x91 & ~x98 & ~x100 & ~x103 & ~x104 & ~x105 & ~x115 & ~x121 & ~x123 & ~x124 & ~x128 & ~x129 & ~x139 & ~x166 & ~x167 & ~x193 & ~x226 & ~x306 & ~x368 & ~x389 & ~x391 & ~x394 & ~x416 & ~x425 & ~x447 & ~x469 & ~x472 & ~x475 & ~x498 & ~x500 & ~x501 & ~x505 & ~x507 & ~x525 & ~x527 & ~x528 & ~x535 & ~x549 & ~x550 & ~x553 & ~x557 & ~x559 & ~x562 & ~x579 & ~x580 & ~x583 & ~x586 & ~x588 & ~x605 & ~x609 & ~x614 & ~x619 & ~x632 & ~x633 & ~x635 & ~x638 & ~x641 & ~x644 & ~x646 & ~x662 & ~x663 & ~x665 & ~x669 & ~x672 & ~x688 & ~x689 & ~x690 & ~x691 & ~x694 & ~x697 & ~x720 & ~x722 & ~x728 & ~x730 & ~x743 & ~x744 & ~x749 & ~x754 & ~x756 & ~x760 & ~x771 & ~x775 & ~x782;
assign c2279 =  x375 &  x659 & ~x25 & ~x97 & ~x133 & ~x224 & ~x574 & ~x726 & ~x731;
assign c2281 =  x400 & ~x130 & ~x185 & ~x240 & ~x706 & ~x751;
assign c2283 =  x426 & ~x11 & ~x14 & ~x18 & ~x34 & ~x36 & ~x48 & ~x61 & ~x86 & ~x91 & ~x99 & ~x119 & ~x137 & ~x166 & ~x196 & ~x197 & ~x250 & ~x254 & ~x309 & ~x338 & ~x376 & ~x403 & ~x421 & ~x532 & ~x562 & ~x563 & ~x586 & ~x591 & ~x613 & ~x676 & ~x679 & ~x724 & ~x736 & ~x756 & ~x765 & ~x772 & ~x774;
assign c2285 =  x318 &  x374 &  x402 & ~x111 & ~x528 & ~x537 & ~x666 & ~x698 & ~x748;
assign c2287 =  x601 & ~x31 & ~x82 & ~x90 & ~x114 & ~x115 & ~x151 & ~x173 & ~x241 & ~x242 & ~x270 & ~x271 & ~x364 & ~x366 & ~x368 & ~x369 & ~x398 & ~x416 & ~x418 & ~x561 & ~x587 & ~x591 & ~x636 & ~x643 & ~x661 & ~x667 & ~x715 & ~x721 & ~x746 & ~x762 & ~x763 & ~x783;
assign c2289 = ~x30 & ~x46 & ~x52 & ~x55 & ~x82 & ~x83 & ~x89 & ~x100 & ~x106 & ~x108 & ~x122 & ~x139 & ~x170 & ~x287 & ~x365 & ~x368 & ~x412 & ~x445 & ~x446 & ~x484 & ~x508 & ~x523 & ~x578 & ~x581 & ~x606 & ~x647 & ~x663 & ~x674 & ~x675 & ~x714 & ~x727 & ~x732 & ~x741 & ~x767;
assign c2291 = ~x16 & ~x18 & ~x21 & ~x26 & ~x27 & ~x32 & ~x67 & ~x72 & ~x79 & ~x82 & ~x87 & ~x89 & ~x93 & ~x116 & ~x195 & ~x199 & ~x227 & ~x334 & ~x384 & ~x393 & ~x421 & ~x423 & ~x429 & ~x448 & ~x462 & ~x487 & ~x491 & ~x502 & ~x504 & ~x506 & ~x531 & ~x532 & ~x586 & ~x611 & ~x613 & ~x639 & ~x641 & ~x668 & ~x672 & ~x694 & ~x714 & ~x715 & ~x720 & ~x726 & ~x734 & ~x736 & ~x744 & ~x764 & ~x767 & ~x777;
assign c2293 = ~x2 & ~x13 & ~x15 & ~x23 & ~x24 & ~x38 & ~x41 & ~x43 & ~x45 & ~x50 & ~x52 & ~x54 & ~x55 & ~x57 & ~x60 & ~x68 & ~x72 & ~x74 & ~x75 & ~x80 & ~x84 & ~x87 & ~x89 & ~x90 & ~x96 & ~x97 & ~x104 & ~x106 & ~x113 & ~x115 & ~x118 & ~x168 & ~x169 & ~x170 & ~x171 & ~x197 & ~x198 & ~x199 & ~x222 & ~x249 & ~x253 & ~x276 & ~x278 & ~x280 & ~x309 & ~x363 & ~x391 & ~x394 & ~x419 & ~x421 & ~x423 & ~x445 & ~x448 & ~x463 & ~x473 & ~x477 & ~x487 & ~x492 & ~x502 & ~x503 & ~x516 & ~x545 & ~x559 & ~x589 & ~x643 & ~x644 & ~x668 & ~x669 & ~x670 & ~x690 & ~x691 & ~x692 & ~x697 & ~x699 & ~x703 & ~x706 & ~x714 & ~x719 & ~x722 & ~x728 & ~x731 & ~x742 & ~x745 & ~x751 & ~x752 & ~x758 & ~x763 & ~x769 & ~x772;
assign c2295 = ~x12 & ~x13 & ~x19 & ~x34 & ~x43 & ~x49 & ~x50 & ~x53 & ~x70 & ~x71 & ~x73 & ~x85 & ~x92 & ~x93 & ~x95 & ~x97 & ~x119 & ~x123 & ~x127 & ~x128 & ~x144 & ~x149 & ~x165 & ~x167 & ~x170 & ~x171 & ~x173 & ~x198 & ~x201 & ~x222 & ~x228 & ~x249 & ~x253 & ~x280 & ~x336 & ~x343 & ~x360 & ~x366 & ~x371 & ~x387 & ~x388 & ~x421 & ~x425 & ~x442 & ~x443 & ~x445 & ~x446 & ~x468 & ~x469 & ~x470 & ~x471 & ~x477 & ~x501 & ~x506 & ~x524 & ~x551 & ~x559 & ~x561 & ~x562 & ~x579 & ~x592 & ~x606 & ~x608 & ~x616 & ~x633 & ~x640 & ~x663 & ~x667 & ~x688 & ~x698 & ~x715 & ~x717 & ~x739 & ~x753 & ~x759 & ~x762 & ~x772 & ~x778 & ~x781 & ~x782;
assign c2297 = ~x5 & ~x15 & ~x23 & ~x34 & ~x48 & ~x55 & ~x72 & ~x73 & ~x87 & ~x90 & ~x92 & ~x94 & ~x99 & ~x100 & ~x102 & ~x105 & ~x112 & ~x114 & ~x117 & ~x120 & ~x121 & ~x122 & ~x123 & ~x134 & ~x136 & ~x140 & ~x144 & ~x147 & ~x150 & ~x173 & ~x174 & ~x178 & ~x196 & ~x257 & ~x281 & ~x335 & ~x337 & ~x343 & ~x360 & ~x366 & ~x385 & ~x390 & ~x398 & ~x421 & ~x422 & ~x443 & ~x468 & ~x470 & ~x472 & ~x473 & ~x476 & ~x481 & ~x498 & ~x500 & ~x502 & ~x524 & ~x525 & ~x528 & ~x560 & ~x579 & ~x581 & ~x588 & ~x591 & ~x606 & ~x607 & ~x617 & ~x633 & ~x640 & ~x661 & ~x666 & ~x670 & ~x674 & ~x676 & ~x678 & ~x688 & ~x693 & ~x697 & ~x699 & ~x712 & ~x717 & ~x718 & ~x719 & ~x724 & ~x726 & ~x727 & ~x739 & ~x742 & ~x746 & ~x750 & ~x753 & ~x757 & ~x759 & ~x762 & ~x764 & ~x765 & ~x768 & ~x769 & ~x776 & ~x780;
assign c2299 = ~x51 & ~x58 & ~x109 & ~x125 & ~x203 & ~x314 & ~x399 & ~x481 & ~x484 & ~x506 & ~x522 & ~x523 & ~x589 & ~x607 & ~x616 & ~x621 & ~x634 & ~x689 & ~x752;
assign c30 =  x675;
assign c32 =  x32;
assign c34 =  x254;
assign c36 = ~x9 & ~x65 & ~x164 & ~x167 & ~x176 & ~x206 & ~x227 & ~x247 & ~x248 & ~x345 & ~x358 & ~x370 & ~x386 & ~x412 & ~x416 & ~x469 & ~x483 & ~x487 & ~x526 & ~x579 & ~x613 & ~x632 & ~x637 & ~x639 & ~x658 & ~x691 & ~x701 & ~x709 & ~x713 & ~x717 & ~x723 & ~x738 & ~x745 & ~x764 & ~x767;
assign c38 =  x178 &  x407 &  x658 &  x659 & ~x1 & ~x26 & ~x31 & ~x45 & ~x53 & ~x57 & ~x79 & ~x96 & ~x100 & ~x110 & ~x111 & ~x136 & ~x138 & ~x163 & ~x168 & ~x171 & ~x194 & ~x196 & ~x197 & ~x225 & ~x226 & ~x246 & ~x251 & ~x280 & ~x290 & ~x305 & ~x307 & ~x317 & ~x331 & ~x337 & ~x344 & ~x360 & ~x362 & ~x387 & ~x393 & ~x398 & ~x419 & ~x444 & ~x448 & ~x449 & ~x474 & ~x504 & ~x530 & ~x531 & ~x534 & ~x557 & ~x562 & ~x588 & ~x591 & ~x611 & ~x612 & ~x618 & ~x638 & ~x643 & ~x666 & ~x668 & ~x675 & ~x694 & ~x697 & ~x701 & ~x715 & ~x728 & ~x729 & ~x739 & ~x741 & ~x752 & ~x754 & ~x762 & ~x769 & ~x771;
assign c310 =  x324 &  x325 &  x350 & ~x1 & ~x5 & ~x10 & ~x14 & ~x15 & ~x22 & ~x24 & ~x34 & ~x36 & ~x42 & ~x43 & ~x44 & ~x46 & ~x54 & ~x55 & ~x61 & ~x65 & ~x75 & ~x76 & ~x80 & ~x81 & ~x82 & ~x84 & ~x88 & ~x89 & ~x92 & ~x94 & ~x96 & ~x109 & ~x112 & ~x114 & ~x138 & ~x141 & ~x142 & ~x163 & ~x165 & ~x193 & ~x224 & ~x225 & ~x226 & ~x250 & ~x252 & ~x260 & ~x277 & ~x281 & ~x282 & ~x284 & ~x287 & ~x288 & ~x289 & ~x291 & ~x304 & ~x308 & ~x313 & ~x314 & ~x330 & ~x336 & ~x364 & ~x367 & ~x393 & ~x445 & ~x446 & ~x448 & ~x459 & ~x460 & ~x473 & ~x475 & ~x504 & ~x505 & ~x529 & ~x533 & ~x557 & ~x559 & ~x560 & ~x561 & ~x587 & ~x588 & ~x589 & ~x613 & ~x615 & ~x617 & ~x639 & ~x666 & ~x671 & ~x684 & ~x685 & ~x690 & ~x692 & ~x694 & ~x697 & ~x701 & ~x702 & ~x705 & ~x707 & ~x711 & ~x712 & ~x714 & ~x715 & ~x720 & ~x726 & ~x727 & ~x733 & ~x737 & ~x740 & ~x745 & ~x748 & ~x753 & ~x766 & ~x767 & ~x774;
assign c312 =  x149 &  x265 &  x291;
assign c314 =  x626 &  x628 &  x629 & ~x0 & ~x6 & ~x8 & ~x15 & ~x27 & ~x28 & ~x29 & ~x30 & ~x33 & ~x34 & ~x35 & ~x42 & ~x56 & ~x64 & ~x69 & ~x80 & ~x86 & ~x90 & ~x104 & ~x108 & ~x110 & ~x131 & ~x140 & ~x161 & ~x163 & ~x165 & ~x167 & ~x168 & ~x174 & ~x189 & ~x197 & ~x201 & ~x218 & ~x219 & ~x223 & ~x225 & ~x247 & ~x254 & ~x275 & ~x277 & ~x284 & ~x304 & ~x306 & ~x333 & ~x337 & ~x359 & ~x361 & ~x387 & ~x420 & ~x421 & ~x422 & ~x447 & ~x454 & ~x455 & ~x474 & ~x477 & ~x503 & ~x506 & ~x513 & ~x514 & ~x526 & ~x532 & ~x533 & ~x534 & ~x555 & ~x557 & ~x560 & ~x562 & ~x585 & ~x609 & ~x613 & ~x619 & ~x639 & ~x641 & ~x646 & ~x665 & ~x669 & ~x670 & ~x680 & ~x683 & ~x692 & ~x693 & ~x697 & ~x702 & ~x706 & ~x711 & ~x713 & ~x714 & ~x717 & ~x728 & ~x737 & ~x751 & ~x754 & ~x755 & ~x756 & ~x759 & ~x762 & ~x764 & ~x769 & ~x778 & ~x779 & ~x782;
assign c316 =  x757;
assign c318 =  x535;
assign c320 =  x184 &  x269 &  x296 &  x322 & ~x1 & ~x25 & ~x48 & ~x71 & ~x76 & ~x117 & ~x138 & ~x164 & ~x191 & ~x247 & ~x300 & ~x301 & ~x309 & ~x339 & ~x370 & ~x452 & ~x485 & ~x505 & ~x507 & ~x515 & ~x516 & ~x535 & ~x542 & ~x561 & ~x670 & ~x694 & ~x718 & ~x725 & ~x730 & ~x732 & ~x759;
assign c322 =  x244 &  x300 & ~x18 & ~x58 & ~x141 & ~x259 & ~x279 & ~x289 & ~x361 & ~x417 & ~x455 & ~x485 & ~x486 & ~x584 & ~x702 & ~x748 & ~x764;
assign c324 =  x183 & ~x29 & ~x33 & ~x39 & ~x49 & ~x56 & ~x57 & ~x103 & ~x109 & ~x129 & ~x134 & ~x162 & ~x171 & ~x191 & ~x247 & ~x252 & ~x266 & ~x279 & ~x309 & ~x320 & ~x347 & ~x356 & ~x367 & ~x383 & ~x395 & ~x425 & ~x428 & ~x429 & ~x471 & ~x473 & ~x501 & ~x510 & ~x527 & ~x530 & ~x537 & ~x554 & ~x572 & ~x582 & ~x585 & ~x610 & ~x731 & ~x757 & ~x760 & ~x766 & ~x778;
assign c326 = ~x25 & ~x29 & ~x43 & ~x48 & ~x54 & ~x57 & ~x69 & ~x70 & ~x71 & ~x83 & ~x89 & ~x92 & ~x104 & ~x227 & ~x247 & ~x254 & ~x289 & ~x308 & ~x310 & ~x317 & ~x342 & ~x359 & ~x367 & ~x387 & ~x444 & ~x450 & ~x462 & ~x475 & ~x486 & ~x488 & ~x490 & ~x491 & ~x494 & ~x512 & ~x514 & ~x669 & ~x671 & ~x703 & ~x724 & ~x731 & ~x734 & ~x735 & ~x766 & ~x780;
assign c328 =  x298 &  x324 &  x325 &  x350 &  x351 & ~x0 & ~x1 & ~x6 & ~x9 & ~x11 & ~x13 & ~x14 & ~x21 & ~x25 & ~x30 & ~x31 & ~x37 & ~x38 & ~x49 & ~x54 & ~x55 & ~x69 & ~x71 & ~x72 & ~x79 & ~x81 & ~x85 & ~x90 & ~x93 & ~x111 & ~x115 & ~x118 & ~x119 & ~x120 & ~x135 & ~x145 & ~x165 & ~x166 & ~x169 & ~x224 & ~x225 & ~x228 & ~x251 & ~x255 & ~x276 & ~x282 & ~x307 & ~x308 & ~x309 & ~x331 & ~x335 & ~x340 & ~x342 & ~x359 & ~x361 & ~x363 & ~x365 & ~x387 & ~x447 & ~x449 & ~x450 & ~x458 & ~x461 & ~x463 & ~x475 & ~x489 & ~x503 & ~x531 & ~x532 & ~x534 & ~x558 & ~x560 & ~x585 & ~x586 & ~x612 & ~x613 & ~x615 & ~x618 & ~x619 & ~x642 & ~x645 & ~x646 & ~x666 & ~x671 & ~x672 & ~x676 & ~x692 & ~x698 & ~x703 & ~x704 & ~x705 & ~x706 & ~x716 & ~x717 & ~x722 & ~x723 & ~x725 & ~x726 & ~x728 & ~x730 & ~x734 & ~x735 & ~x739 & ~x742 & ~x744 & ~x745 & ~x747 & ~x748 & ~x751 & ~x755 & ~x758 & ~x759 & ~x766 & ~x770 & ~x771 & ~x775 & ~x777 & ~x778 & ~x781;
assign c330 =  x322 & ~x9 & ~x17 & ~x33 & ~x38 & ~x47 & ~x57 & ~x106 & ~x144 & ~x191 & ~x193 & ~x194 & ~x233 & ~x235 & ~x236 & ~x248 & ~x260 & ~x286 & ~x333 & ~x339 & ~x387 & ~x419 & ~x431 & ~x432 & ~x433 & ~x445 & ~x462 & ~x474 & ~x561 & ~x585 & ~x612 & ~x614 & ~x619 & ~x621 & ~x698 & ~x700 & ~x710 & ~x717 & ~x732 & ~x735 & ~x748 & ~x764 & ~x768 & ~x776 & ~x778 & ~x780;
assign c332 =  x406 &  x524 &  x607 & ~x5 & ~x13 & ~x30 & ~x32 & ~x43 & ~x45 & ~x70 & ~x90 & ~x114 & ~x126 & ~x127 & ~x132 & ~x133 & ~x161 & ~x166 & ~x191 & ~x195 & ~x248 & ~x280 & ~x334 & ~x338 & ~x387 & ~x396 & ~x423 & ~x452 & ~x484 & ~x485 & ~x504 & ~x515 & ~x534 & ~x557 & ~x560 & ~x561 & ~x615 & ~x619 & ~x641 & ~x645 & ~x666 & ~x677 & ~x678 & ~x692 & ~x695 & ~x697 & ~x721 & ~x736 & ~x746 & ~x747 & ~x752 & ~x761 & ~x767;
assign c334 =  x265 & ~x132 & ~x157 & ~x453 & ~x485 & ~x486 & ~x491 & ~x511 & ~x513;
assign c336 =  x49;
assign c338 =  x40;
assign c340 =  x432 &  x433 & ~x22 & ~x24 & ~x28 & ~x29 & ~x31 & ~x33 & ~x39 & ~x54 & ~x57 & ~x58 & ~x63 & ~x69 & ~x83 & ~x93 & ~x94 & ~x95 & ~x101 & ~x114 & ~x117 & ~x121 & ~x140 & ~x144 & ~x165 & ~x199 & ~x200 & ~x248 & ~x250 & ~x253 & ~x276 & ~x319 & ~x340 & ~x341 & ~x342 & ~x343 & ~x345 & ~x360 & ~x368 & ~x390 & ~x392 & ~x394 & ~x424 & ~x442 & ~x446 & ~x450 & ~x454 & ~x477 & ~x478 & ~x498 & ~x515 & ~x516 & ~x530 & ~x533 & ~x562 & ~x582 & ~x585 & ~x611 & ~x616 & ~x672 & ~x673 & ~x695 & ~x705 & ~x742 & ~x746 & ~x758 & ~x765 & ~x778;
assign c342 =  x705 &  x738;
assign c344 =  x476;
assign c346 =  x210 & ~x3 & ~x4 & ~x5 & ~x10 & ~x12 & ~x15 & ~x19 & ~x21 & ~x23 & ~x37 & ~x43 & ~x46 & ~x56 & ~x68 & ~x71 & ~x73 & ~x76 & ~x88 & ~x89 & ~x95 & ~x107 & ~x126 & ~x146 & ~x158 & ~x194 & ~x217 & ~x223 & ~x224 & ~x250 & ~x274 & ~x280 & ~x305 & ~x310 & ~x311 & ~x312 & ~x313 & ~x339 & ~x366 & ~x388 & ~x425 & ~x444 & ~x451 & ~x455 & ~x476 & ~x478 & ~x480 & ~x503 & ~x510 & ~x532 & ~x533 & ~x534 & ~x537 & ~x540 & ~x546 & ~x558 & ~x568 & ~x570 & ~x610 & ~x615 & ~x618 & ~x645 & ~x669 & ~x674 & ~x692 & ~x700 & ~x701 & ~x716 & ~x717 & ~x718 & ~x722 & ~x723 & ~x733 & ~x736 & ~x743 & ~x751 & ~x761 & ~x765 & ~x771 & ~x780;
assign c348 = ~x2 & ~x5 & ~x7 & ~x10 & ~x13 & ~x25 & ~x27 & ~x30 & ~x33 & ~x36 & ~x43 & ~x47 & ~x49 & ~x59 & ~x68 & ~x73 & ~x75 & ~x76 & ~x77 & ~x106 & ~x113 & ~x130 & ~x131 & ~x158 & ~x159 & ~x160 & ~x164 & ~x191 & ~x219 & ~x222 & ~x245 & ~x248 & ~x249 & ~x252 & ~x272 & ~x282 & ~x300 & ~x303 & ~x308 & ~x313 & ~x331 & ~x332 & ~x344 & ~x362 & ~x386 & ~x390 & ~x392 & ~x394 & ~x419 & ~x423 & ~x425 & ~x454 & ~x475 & ~x479 & ~x482 & ~x508 & ~x510 & ~x511 & ~x529 & ~x531 & ~x534 & ~x536 & ~x545 & ~x557 & ~x560 & ~x570 & ~x574 & ~x575 & ~x588 & ~x592 & ~x618 & ~x650 & ~x667 & ~x698 & ~x701 & ~x704 & ~x730 & ~x733 & ~x735 & ~x743 & ~x745 & ~x746 & ~x748 & ~x750 & ~x753 & ~x755 & ~x762 & ~x768;
assign c350 =  x172;
assign c352 =  x209 & ~x4 & ~x13 & ~x14 & ~x18 & ~x26 & ~x30 & ~x33 & ~x39 & ~x47 & ~x67 & ~x71 & ~x95 & ~x110 & ~x114 & ~x124 & ~x129 & ~x146 & ~x194 & ~x224 & ~x225 & ~x246 & ~x282 & ~x284 & ~x293 & ~x305 & ~x311 & ~x333 & ~x347 & ~x372 & ~x389 & ~x414 & ~x426 & ~x500 & ~x528 & ~x529 & ~x534 & ~x542 & ~x544 & ~x545 & ~x554 & ~x587 & ~x590 & ~x618 & ~x674 & ~x722 & ~x725 & ~x736 & ~x737 & ~x742 & ~x755 & ~x756 & ~x769 & ~x776 & ~x783;
assign c354 =  x269 &  x296 &  x322 & ~x9 & ~x13 & ~x14 & ~x15 & ~x17 & ~x21 & ~x25 & ~x28 & ~x30 & ~x34 & ~x37 & ~x41 & ~x49 & ~x57 & ~x62 & ~x66 & ~x68 & ~x70 & ~x78 & ~x89 & ~x91 & ~x102 & ~x111 & ~x113 & ~x118 & ~x133 & ~x134 & ~x135 & ~x136 & ~x144 & ~x146 & ~x164 & ~x166 & ~x172 & ~x190 & ~x191 & ~x192 & ~x195 & ~x196 & ~x220 & ~x225 & ~x247 & ~x248 & ~x249 & ~x252 & ~x253 & ~x273 & ~x279 & ~x281 & ~x300 & ~x302 & ~x305 & ~x308 & ~x313 & ~x330 & ~x331 & ~x333 & ~x335 & ~x340 & ~x360 & ~x364 & ~x387 & ~x389 & ~x417 & ~x418 & ~x419 & ~x423 & ~x424 & ~x445 & ~x447 & ~x449 & ~x450 & ~x451 & ~x472 & ~x473 & ~x475 & ~x478 & ~x488 & ~x489 & ~x504 & ~x505 & ~x506 & ~x530 & ~x535 & ~x556 & ~x560 & ~x561 & ~x564 & ~x586 & ~x591 & ~x592 & ~x612 & ~x617 & ~x618 & ~x641 & ~x646 & ~x664 & ~x669 & ~x671 & ~x687 & ~x694 & ~x698 & ~x702 & ~x704 & ~x709 & ~x714 & ~x716 & ~x720 & ~x721 & ~x722 & ~x727 & ~x730 & ~x733 & ~x736 & ~x741 & ~x746 & ~x752 & ~x757 & ~x758 & ~x760 & ~x762 & ~x766 & ~x779 & ~x780;
assign c356 =  x209 &  x434 &  x685 & ~x0 & ~x5 & ~x27 & ~x34 & ~x39 & ~x45 & ~x60 & ~x66 & ~x71 & ~x72 & ~x113 & ~x116 & ~x130 & ~x170 & ~x198 & ~x282 & ~x308 & ~x309 & ~x333 & ~x337 & ~x362 & ~x392 & ~x394 & ~x397 & ~x398 & ~x473 & ~x474 & ~x483 & ~x502 & ~x503 & ~x541 & ~x568 & ~x570 & ~x572 & ~x645 & ~x672 & ~x704 & ~x720 & ~x724 & ~x734 & ~x737 & ~x751 & ~x768 & ~x778 & ~x780;
assign c358 = ~x18 & ~x21 & ~x54 & ~x72 & ~x80 & ~x85 & ~x111 & ~x117 & ~x135 & ~x146 & ~x165 & ~x191 & ~x222 & ~x264 & ~x266 & ~x283 & ~x285 & ~x288 & ~x331 & ~x333 & ~x357 & ~x362 & ~x368 & ~x427 & ~x445 & ~x455 & ~x469 & ~x484 & ~x615 & ~x691 & ~x715 & ~x717 & ~x738 & ~x755 & ~x762;
assign c360 =  x449;
assign c362 =  x406 & ~x1 & ~x5 & ~x9 & ~x10 & ~x11 & ~x23 & ~x25 & ~x29 & ~x30 & ~x33 & ~x41 & ~x42 & ~x49 & ~x54 & ~x57 & ~x66 & ~x73 & ~x90 & ~x99 & ~x103 & ~x104 & ~x119 & ~x123 & ~x125 & ~x128 & ~x131 & ~x138 & ~x143 & ~x167 & ~x168 & ~x192 & ~x196 & ~x198 & ~x225 & ~x249 & ~x292 & ~x315 & ~x316 & ~x319 & ~x332 & ~x343 & ~x344 & ~x358 & ~x361 & ~x368 & ~x369 & ~x371 & ~x389 & ~x395 & ~x424 & ~x445 & ~x453 & ~x477 & ~x480 & ~x481 & ~x504 & ~x505 & ~x511 & ~x533 & ~x541 & ~x542 & ~x556 & ~x557 & ~x589 & ~x617 & ~x669 & ~x670 & ~x673 & ~x693 & ~x700 & ~x705 & ~x732 & ~x735 & ~x759 & ~x778 & ~x779;
assign c364 =  x353 &  x378 &  x469 &  x525 &  x580 & ~x109 & ~x371 & ~x399 & ~x640;
assign c366 =  x599 & ~x0 & ~x3 & ~x5 & ~x11 & ~x27 & ~x29 & ~x30 & ~x35 & ~x41 & ~x43 & ~x47 & ~x50 & ~x53 & ~x57 & ~x59 & ~x61 & ~x63 & ~x81 & ~x86 & ~x91 & ~x92 & ~x112 & ~x134 & ~x145 & ~x161 & ~x163 & ~x191 & ~x226 & ~x247 & ~x305 & ~x334 & ~x342 & ~x365 & ~x415 & ~x417 & ~x418 & ~x419 & ~x421 & ~x474 & ~x488 & ~x498 & ~x530 & ~x579 & ~x606 & ~x617 & ~x635 & ~x686 & ~x706 & ~x709 & ~x710 & ~x715 & ~x724 & ~x729 & ~x741 & ~x748 & ~x761 & ~x764 & ~x775;
assign c368 =  x564 & ~x482;
assign c370 =  x647;
assign c372 =  x267 &  x319 &  x321 & ~x6 & ~x10 & ~x26 & ~x28 & ~x61 & ~x63 & ~x65 & ~x75 & ~x104 & ~x109 & ~x113 & ~x187 & ~x248 & ~x272 & ~x273 & ~x288 & ~x303 & ~x393 & ~x427 & ~x473 & ~x533 & ~x563 & ~x610 & ~x695 & ~x697 & ~x707 & ~x720 & ~x734 & ~x742 & ~x780 & ~x781 & ~x783;
assign c374 =  x294 & ~x4 & ~x8 & ~x9 & ~x13 & ~x15 & ~x16 & ~x28 & ~x37 & ~x38 & ~x56 & ~x57 & ~x69 & ~x70 & ~x85 & ~x100 & ~x106 & ~x107 & ~x110 & ~x112 & ~x131 & ~x132 & ~x137 & ~x143 & ~x145 & ~x160 & ~x161 & ~x164 & ~x167 & ~x189 & ~x190 & ~x192 & ~x195 & ~x196 & ~x197 & ~x216 & ~x226 & ~x227 & ~x244 & ~x245 & ~x248 & ~x250 & ~x253 & ~x276 & ~x277 & ~x278 & ~x299 & ~x300 & ~x304 & ~x305 & ~x306 & ~x309 & ~x327 & ~x329 & ~x332 & ~x336 & ~x338 & ~x356 & ~x358 & ~x363 & ~x366 & ~x387 & ~x390 & ~x397 & ~x417 & ~x419 & ~x422 & ~x425 & ~x449 & ~x450 & ~x476 & ~x485 & ~x486 & ~x490 & ~x503 & ~x509 & ~x516 & ~x529 & ~x587 & ~x592 & ~x617 & ~x641 & ~x665 & ~x690 & ~x691 & ~x706 & ~x715 & ~x717 & ~x718 & ~x719 & ~x720 & ~x721 & ~x722 & ~x724 & ~x725 & ~x727 & ~x730 & ~x734 & ~x736 & ~x742 & ~x757 & ~x764 & ~x767 & ~x772 & ~x775 & ~x777;
assign c376 =  x168;
assign c378 =  x326 &  x536 & ~x429;
assign c380 =  x353 &  x378 & ~x5 & ~x14 & ~x15 & ~x17 & ~x24 & ~x27 & ~x30 & ~x37 & ~x42 & ~x44 & ~x53 & ~x57 & ~x59 & ~x60 & ~x62 & ~x63 & ~x77 & ~x81 & ~x85 & ~x91 & ~x94 & ~x95 & ~x106 & ~x107 & ~x114 & ~x136 & ~x142 & ~x143 & ~x165 & ~x172 & ~x196 & ~x199 & ~x227 & ~x283 & ~x305 & ~x308 & ~x318 & ~x336 & ~x344 & ~x362 & ~x363 & ~x366 & ~x371 & ~x388 & ~x399 & ~x418 & ~x456 & ~x485 & ~x486 & ~x487 & ~x488 & ~x529 & ~x530 & ~x531 & ~x556 & ~x560 & ~x585 & ~x638 & ~x640 & ~x642 & ~x669 & ~x670 & ~x673 & ~x676 & ~x704 & ~x706 & ~x709 & ~x711 & ~x715 & ~x724 & ~x737 & ~x742 & ~x748 & ~x750 & ~x751 & ~x753 & ~x755 & ~x761 & ~x762 & ~x775 & ~x779 & ~x781 & ~x783;
assign c382 =  x685 & ~x10 & ~x19 & ~x24 & ~x42 & ~x51 & ~x55 & ~x137 & ~x190 & ~x191 & ~x217 & ~x219 & ~x220 & ~x273 & ~x329 & ~x330 & ~x331 & ~x332 & ~x335 & ~x360 & ~x385 & ~x388 & ~x420 & ~x480 & ~x540 & ~x571 & ~x573 & ~x574 & ~x599 & ~x627 & ~x649 & ~x672 & ~x673 & ~x674 & ~x696 & ~x705 & ~x706 & ~x722 & ~x724 & ~x729 & ~x744 & ~x747 & ~x757 & ~x759 & ~x760 & ~x761 & ~x770;
assign c384 =  x127 &  x601 &  x626 & ~x0 & ~x1 & ~x12 & ~x13 & ~x14 & ~x17 & ~x18 & ~x26 & ~x29 & ~x30 & ~x37 & ~x56 & ~x61 & ~x64 & ~x67 & ~x86 & ~x87 & ~x88 & ~x90 & ~x91 & ~x92 & ~x94 & ~x106 & ~x110 & ~x114 & ~x118 & ~x135 & ~x145 & ~x165 & ~x172 & ~x173 & ~x174 & ~x195 & ~x197 & ~x202 & ~x206 & ~x221 & ~x232 & ~x234 & ~x247 & ~x257 & ~x259 & ~x260 & ~x302 & ~x310 & ~x311 & ~x329 & ~x341 & ~x357 & ~x358 & ~x359 & ~x363 & ~x364 & ~x391 & ~x416 & ~x420 & ~x443 & ~x445 & ~x500 & ~x531 & ~x533 & ~x555 & ~x557 & ~x581 & ~x586 & ~x611 & ~x612 & ~x615 & ~x636 & ~x641 & ~x643 & ~x660 & ~x672 & ~x680 & ~x682 & ~x684 & ~x690 & ~x694 & ~x702 & ~x710 & ~x711 & ~x723 & ~x731 & ~x732 & ~x737 & ~x739 & ~x749 & ~x750 & ~x751 & ~x761 & ~x763 & ~x765 & ~x766 & ~x767 & ~x776;
assign c386 =  x655 & ~x16 & ~x20 & ~x21 & ~x23 & ~x24 & ~x25 & ~x29 & ~x44 & ~x45 & ~x51 & ~x57 & ~x60 & ~x62 & ~x64 & ~x67 & ~x77 & ~x79 & ~x91 & ~x114 & ~x115 & ~x118 & ~x143 & ~x163 & ~x164 & ~x167 & ~x170 & ~x190 & ~x236 & ~x247 & ~x253 & ~x262 & ~x275 & ~x276 & ~x278 & ~x282 & ~x289 & ~x303 & ~x359 & ~x365 & ~x390 & ~x396 & ~x416 & ~x445 & ~x481 & ~x504 & ~x528 & ~x531 & ~x544 & ~x562 & ~x616 & ~x619 & ~x638 & ~x690 & ~x691 & ~x698 & ~x710 & ~x714 & ~x716 & ~x717 & ~x732 & ~x733 & ~x735 & ~x747 & ~x759 & ~x778 & ~x782;
assign c388 =  x21;
assign c390 =  x404 & ~x4 & ~x9 & ~x12 & ~x32 & ~x41 & ~x43 & ~x45 & ~x50 & ~x61 & ~x64 & ~x70 & ~x72 & ~x80 & ~x83 & ~x92 & ~x102 & ~x111 & ~x134 & ~x138 & ~x140 & ~x230 & ~x248 & ~x253 & ~x255 & ~x282 & ~x284 & ~x307 & ~x309 & ~x319 & ~x320 & ~x321 & ~x333 & ~x335 & ~x346 & ~x367 & ~x372 & ~x389 & ~x391 & ~x421 & ~x441 & ~x443 & ~x470 & ~x477 & ~x504 & ~x513 & ~x515 & ~x582 & ~x586 & ~x587 & ~x610 & ~x611 & ~x612 & ~x643 & ~x645 & ~x665 & ~x697 & ~x701 & ~x704 & ~x728 & ~x738 & ~x750 & ~x751 & ~x758 & ~x760 & ~x780;
assign c394 =  x185 &  x380 &  x381 &  x406 &  x407 &  x625 & ~x4 & ~x7 & ~x9 & ~x15 & ~x23 & ~x26 & ~x32 & ~x38 & ~x43 & ~x45 & ~x51 & ~x52 & ~x54 & ~x68 & ~x69 & ~x86 & ~x88 & ~x96 & ~x99 & ~x100 & ~x141 & ~x165 & ~x168 & ~x170 & ~x193 & ~x221 & ~x225 & ~x344 & ~x361 & ~x367 & ~x388 & ~x389 & ~x391 & ~x392 & ~x419 & ~x422 & ~x447 & ~x476 & ~x502 & ~x513 & ~x515 & ~x530 & ~x560 & ~x583 & ~x645 & ~x667 & ~x694 & ~x723 & ~x736 & ~x748 & ~x750 & ~x753 & ~x769 & ~x774 & ~x776 & ~x781;
assign c396 =  x224;
assign c398 = ~x44 & ~x73 & ~x79 & ~x87 & ~x129 & ~x139 & ~x158 & ~x160 & ~x190 & ~x219 & ~x243 & ~x244 & ~x273 & ~x274 & ~x304 & ~x449 & ~x458 & ~x460 & ~x490 & ~x502 & ~x519 & ~x559 & ~x594 & ~x614 & ~x641 & ~x686 & ~x695 & ~x701 & ~x741 & ~x743 & ~x759 & ~x774;
assign c3100 =  x266 & ~x1 & ~x3 & ~x5 & ~x11 & ~x13 & ~x14 & ~x15 & ~x17 & ~x18 & ~x19 & ~x22 & ~x24 & ~x25 & ~x26 & ~x27 & ~x30 & ~x32 & ~x33 & ~x34 & ~x36 & ~x38 & ~x40 & ~x42 & ~x47 & ~x49 & ~x50 & ~x51 & ~x52 & ~x53 & ~x55 & ~x57 & ~x58 & ~x60 & ~x69 & ~x71 & ~x73 & ~x74 & ~x76 & ~x77 & ~x78 & ~x79 & ~x84 & ~x87 & ~x90 & ~x103 & ~x104 & ~x105 & ~x106 & ~x108 & ~x111 & ~x112 & ~x115 & ~x116 & ~x132 & ~x135 & ~x141 & ~x142 & ~x143 & ~x144 & ~x166 & ~x169 & ~x171 & ~x172 & ~x188 & ~x189 & ~x190 & ~x191 & ~x192 & ~x196 & ~x197 & ~x199 & ~x216 & ~x218 & ~x220 & ~x221 & ~x222 & ~x223 & ~x224 & ~x227 & ~x246 & ~x247 & ~x248 & ~x250 & ~x251 & ~x253 & ~x254 & ~x272 & ~x275 & ~x277 & ~x278 & ~x279 & ~x280 & ~x282 & ~x302 & ~x305 & ~x306 & ~x307 & ~x309 & ~x311 & ~x312 & ~x329 & ~x330 & ~x331 & ~x332 & ~x333 & ~x337 & ~x339 & ~x358 & ~x360 & ~x361 & ~x363 & ~x364 & ~x368 & ~x388 & ~x389 & ~x392 & ~x393 & ~x394 & ~x395 & ~x416 & ~x419 & ~x420 & ~x421 & ~x422 & ~x423 & ~x444 & ~x446 & ~x448 & ~x456 & ~x474 & ~x479 & ~x480 & ~x483 & ~x485 & ~x486 & ~x488 & ~x489 & ~x490 & ~x502 & ~x505 & ~x507 & ~x514 & ~x515 & ~x529 & ~x530 & ~x534 & ~x535 & ~x556 & ~x558 & ~x560 & ~x562 & ~x563 & ~x585 & ~x587 & ~x589 & ~x590 & ~x614 & ~x616 & ~x618 & ~x620 & ~x641 & ~x642 & ~x643 & ~x644 & ~x645 & ~x646 & ~x649 & ~x667 & ~x669 & ~x670 & ~x671 & ~x672 & ~x675 & ~x677 & ~x689 & ~x691 & ~x692 & ~x694 & ~x699 & ~x700 & ~x701 & ~x704 & ~x706 & ~x709 & ~x711 & ~x718 & ~x719 & ~x720 & ~x721 & ~x723 & ~x725 & ~x727 & ~x728 & ~x731 & ~x732 & ~x733 & ~x734 & ~x740 & ~x741 & ~x742 & ~x743 & ~x745 & ~x746 & ~x747 & ~x749 & ~x750 & ~x751 & ~x753 & ~x756 & ~x757 & ~x758 & ~x759 & ~x761 & ~x765 & ~x767 & ~x769 & ~x770 & ~x772 & ~x773 & ~x774 & ~x775 & ~x776 & ~x778 & ~x780 & ~x781 & ~x782 & ~x783;
assign c3102 =  x154 & ~x2 & ~x9 & ~x27 & ~x46 & ~x55 & ~x72 & ~x77 & ~x87 & ~x132 & ~x166 & ~x209 & ~x219 & ~x235 & ~x248 & ~x261 & ~x274 & ~x283 & ~x302 & ~x303 & ~x330 & ~x394 & ~x395 & ~x463 & ~x490 & ~x503 & ~x531 & ~x555 & ~x583 & ~x611 & ~x638 & ~x643 & ~x696 & ~x710 & ~x718 & ~x731 & ~x741 & ~x749 & ~x761 & ~x776 & ~x780;
assign c3104 =  x34;
assign c3106 =  x336;
assign c3108 = ~x6 & ~x16 & ~x29 & ~x33 & ~x55 & ~x60 & ~x66 & ~x67 & ~x80 & ~x89 & ~x105 & ~x114 & ~x140 & ~x141 & ~x166 & ~x169 & ~x174 & ~x191 & ~x221 & ~x223 & ~x232 & ~x235 & ~x247 & ~x250 & ~x258 & ~x260 & ~x275 & ~x280 & ~x281 & ~x285 & ~x287 & ~x289 & ~x303 & ~x307 & ~x331 & ~x334 & ~x343 & ~x357 & ~x358 & ~x359 & ~x360 & ~x361 & ~x363 & ~x364 & ~x388 & ~x393 & ~x394 & ~x415 & ~x417 & ~x419 & ~x421 & ~x429 & ~x462 & ~x472 & ~x474 & ~x486 & ~x503 & ~x526 & ~x532 & ~x533 & ~x562 & ~x582 & ~x584 & ~x587 & ~x610 & ~x614 & ~x647 & ~x666 & ~x670 & ~x674 & ~x679 & ~x683 & ~x684 & ~x688 & ~x691 & ~x708 & ~x712 & ~x714 & ~x723 & ~x740 & ~x748 & ~x765 & ~x769 & ~x770 & ~x771 & ~x779;
assign c3110 =  x142;
assign c3112 =  x269 &  x297 &  x324 &  x377 & ~x10 & ~x11 & ~x31 & ~x35 & ~x56 & ~x62 & ~x64 & ~x65 & ~x66 & ~x78 & ~x85 & ~x87 & ~x105 & ~x114 & ~x115 & ~x134 & ~x166 & ~x192 & ~x194 & ~x195 & ~x222 & ~x225 & ~x226 & ~x247 & ~x250 & ~x275 & ~x283 & ~x290 & ~x291 & ~x306 & ~x358 & ~x359 & ~x362 & ~x363 & ~x387 & ~x419 & ~x421 & ~x474 & ~x475 & ~x487 & ~x488 & ~x531 & ~x559 & ~x584 & ~x587 & ~x590 & ~x642 & ~x665 & ~x666 & ~x674 & ~x715 & ~x721 & ~x723 & ~x730 & ~x734 & ~x736 & ~x738 & ~x743 & ~x755 & ~x768 & ~x774 & ~x782;
assign c3114 =  x216 &  x245 &  x326 &  x327 &  x352 &  x378 & ~x485 & ~x514;
assign c3116 = ~x3 & ~x7 & ~x14 & ~x23 & ~x26 & ~x32 & ~x33 & ~x34 & ~x36 & ~x39 & ~x47 & ~x48 & ~x57 & ~x91 & ~x95 & ~x147 & ~x162 & ~x163 & ~x164 & ~x172 & ~x174 & ~x191 & ~x196 & ~x197 & ~x198 & ~x205 & ~x219 & ~x221 & ~x248 & ~x262 & ~x266 & ~x287 & ~x291 & ~x305 & ~x308 & ~x389 & ~x414 & ~x415 & ~x417 & ~x441 & ~x472 & ~x474 & ~x482 & ~x500 & ~x516 & ~x526 & ~x532 & ~x533 & ~x535 & ~x558 & ~x583 & ~x586 & ~x588 & ~x611 & ~x636 & ~x637 & ~x638 & ~x667 & ~x668 & ~x673 & ~x703 & ~x711 & ~x731 & ~x735 & ~x736 & ~x745 & ~x759 & ~x767 & ~x770 & ~x780;
assign c3118 =  x390;
assign c3120 =  x405 &  x564 & ~x426 & ~x427 & ~x485;
assign c3122 =  x182 &  x184 &  x209 &  x210 &  x212 &  x213 &  x378 &  x404 &  x434 & ~x5 & ~x8 & ~x9 & ~x17 & ~x21 & ~x24 & ~x28 & ~x34 & ~x38 & ~x42 & ~x46 & ~x47 & ~x53 & ~x60 & ~x65 & ~x69 & ~x70 & ~x71 & ~x72 & ~x81 & ~x82 & ~x84 & ~x88 & ~x90 & ~x94 & ~x97 & ~x106 & ~x107 & ~x108 & ~x111 & ~x117 & ~x133 & ~x140 & ~x167 & ~x172 & ~x194 & ~x200 & ~x219 & ~x222 & ~x225 & ~x226 & ~x249 & ~x253 & ~x276 & ~x307 & ~x331 & ~x337 & ~x338 & ~x342 & ~x343 & ~x362 & ~x365 & ~x366 & ~x370 & ~x390 & ~x392 & ~x397 & ~x417 & ~x422 & ~x425 & ~x444 & ~x446 & ~x452 & ~x453 & ~x476 & ~x477 & ~x478 & ~x481 & ~x482 & ~x503 & ~x505 & ~x529 & ~x584 & ~x614 & ~x616 & ~x640 & ~x644 & ~x645 & ~x667 & ~x670 & ~x693 & ~x697 & ~x700 & ~x704 & ~x719 & ~x725 & ~x729 & ~x730 & ~x733 & ~x737 & ~x740 & ~x746 & ~x752 & ~x754 & ~x762 & ~x776 & ~x778 & ~x783;
assign c3124 =  x125 &  x321 & ~x33 & ~x141 & ~x163 & ~x191 & ~x208 & ~x234 & ~x246 & ~x391 & ~x476 & ~x555 & ~x745;
assign c3126 =  x124 &  x292 & ~x429;
assign c3128 =  x110;
assign c3130 = ~x2 & ~x15 & ~x16 & ~x19 & ~x21 & ~x24 & ~x26 & ~x35 & ~x38 & ~x43 & ~x44 & ~x49 & ~x53 & ~x56 & ~x59 & ~x61 & ~x63 & ~x65 & ~x69 & ~x71 & ~x74 & ~x86 & ~x91 & ~x108 & ~x109 & ~x113 & ~x115 & ~x117 & ~x129 & ~x130 & ~x132 & ~x158 & ~x161 & ~x162 & ~x167 & ~x168 & ~x170 & ~x172 & ~x174 & ~x195 & ~x197 & ~x201 & ~x202 & ~x219 & ~x227 & ~x247 & ~x254 & ~x256 & ~x258 & ~x277 & ~x279 & ~x284 & ~x304 & ~x305 & ~x307 & ~x308 & ~x309 & ~x318 & ~x334 & ~x338 & ~x343 & ~x360 & ~x365 & ~x366 & ~x370 & ~x388 & ~x395 & ~x412 & ~x419 & ~x445 & ~x450 & ~x451 & ~x452 & ~x453 & ~x473 & ~x475 & ~x478 & ~x512 & ~x514 & ~x531 & ~x533 & ~x535 & ~x543 & ~x544 & ~x545 & ~x557 & ~x561 & ~x562 & ~x563 & ~x590 & ~x591 & ~x609 & ~x611 & ~x616 & ~x617 & ~x621 & ~x622 & ~x637 & ~x639 & ~x640 & ~x645 & ~x646 & ~x666 & ~x669 & ~x674 & ~x691 & ~x693 & ~x694 & ~x702 & ~x703 & ~x717 & ~x724 & ~x727 & ~x728 & ~x729 & ~x730 & ~x732 & ~x733 & ~x747 & ~x748 & ~x749 & ~x750 & ~x752 & ~x754 & ~x756 & ~x758 & ~x764 & ~x766 & ~x767 & ~x769 & ~x771 & ~x774 & ~x781 & ~x783;
assign c3132 =  x200;
assign c3134 =  x272 &  x352 &  x575 & ~x15 & ~x26 & ~x46 & ~x65 & ~x92 & ~x111 & ~x229 & ~x257 & ~x287 & ~x291 & ~x292 & ~x309 & ~x479 & ~x502 & ~x526 & ~x530 & ~x552 & ~x557 & ~x607 & ~x608 & ~x714 & ~x723 & ~x762 & ~x766 & ~x773;
assign c3136 =  x187 &  x242 &  x550 &  x603 &  x604 & ~x3 & ~x4 & ~x12 & ~x16 & ~x73 & ~x88 & ~x90 & ~x92 & ~x94 & ~x109 & ~x115 & ~x163 & ~x192 & ~x201 & ~x249 & ~x275 & ~x332 & ~x336 & ~x338 & ~x345 & ~x346 & ~x362 & ~x369 & ~x371 & ~x445 & ~x446 & ~x472 & ~x502 & ~x527 & ~x533 & ~x555 & ~x556 & ~x562 & ~x610 & ~x614 & ~x638 & ~x643 & ~x665 & ~x674 & ~x675 & ~x716 & ~x717 & ~x732 & ~x735 & ~x754 & ~x770 & ~x772;
assign c3138 =  x155 &  x240 &  x266 &  x267 & ~x16 & ~x88 & ~x135 & ~x188 & ~x244 & ~x274 & ~x305 & ~x361 & ~x417 & ~x426 & ~x488 & ~x490 & ~x506 & ~x562 & ~x587 & ~x701 & ~x714 & ~x728;
assign c3140 = ~x5 & ~x11 & ~x19 & ~x23 & ~x50 & ~x52 & ~x78 & ~x81 & ~x96 & ~x97 & ~x102 & ~x137 & ~x147 & ~x162 & ~x164 & ~x189 & ~x193 & ~x194 & ~x226 & ~x227 & ~x229 & ~x253 & ~x282 & ~x292 & ~x293 & ~x310 & ~x317 & ~x318 & ~x319 & ~x342 & ~x345 & ~x362 & ~x388 & ~x399 & ~x412 & ~x422 & ~x447 & ~x480 & ~x497 & ~x527 & ~x542 & ~x572 & ~x592 & ~x636 & ~x676 & ~x690 & ~x693 & ~x696 & ~x697 & ~x699 & ~x705 & ~x718 & ~x720 & ~x721 & ~x744 & ~x746 & ~x747 & ~x760 & ~x761;
assign c3142 =  x209 &  x434 & ~x18 & ~x19 & ~x22 & ~x25 & ~x27 & ~x36 & ~x41 & ~x52 & ~x55 & ~x64 & ~x77 & ~x83 & ~x104 & ~x130 & ~x139 & ~x142 & ~x163 & ~x164 & ~x165 & ~x170 & ~x250 & ~x251 & ~x274 & ~x275 & ~x284 & ~x294 & ~x333 & ~x335 & ~x347 & ~x358 & ~x359 & ~x361 & ~x389 & ~x425 & ~x427 & ~x498 & ~x507 & ~x527 & ~x537 & ~x554 & ~x559 & ~x570 & ~x572 & ~x610 & ~x614 & ~x618 & ~x619 & ~x667 & ~x672 & ~x692 & ~x719 & ~x733 & ~x739 & ~x741 & ~x742 & ~x743 & ~x765 & ~x772 & ~x782;
assign c3144 =  x700;
assign c3146 =  x678;
assign c3148 =  x180 & ~x6 & ~x7 & ~x11 & ~x12 & ~x20 & ~x29 & ~x32 & ~x43 & ~x45 & ~x56 & ~x58 & ~x67 & ~x68 & ~x71 & ~x85 & ~x91 & ~x96 & ~x98 & ~x99 & ~x108 & ~x112 & ~x132 & ~x134 & ~x137 & ~x168 & ~x194 & ~x220 & ~x262 & ~x264 & ~x275 & ~x282 & ~x288 & ~x290 & ~x311 & ~x329 & ~x338 & ~x339 & ~x359 & ~x369 & ~x385 & ~x390 & ~x391 & ~x395 & ~x396 & ~x397 & ~x415 & ~x419 & ~x420 & ~x422 & ~x444 & ~x453 & ~x470 & ~x476 & ~x479 & ~x500 & ~x531 & ~x534 & ~x555 & ~x556 & ~x559 & ~x571 & ~x589 & ~x592 & ~x611 & ~x615 & ~x619 & ~x638 & ~x639 & ~x640 & ~x643 & ~x646 & ~x665 & ~x666 & ~x671 & ~x677 & ~x700 & ~x730 & ~x736 & ~x743 & ~x746 & ~x748 & ~x751 & ~x755 & ~x757 & ~x761 & ~x770 & ~x774 & ~x776;
assign c3150 =  x335 &  x615;
assign c3152 =  x376 & ~x1 & ~x2 & ~x3 & ~x6 & ~x8 & ~x9 & ~x10 & ~x12 & ~x13 & ~x15 & ~x16 & ~x19 & ~x22 & ~x26 & ~x28 & ~x29 & ~x32 & ~x35 & ~x42 & ~x46 & ~x51 & ~x52 & ~x55 & ~x63 & ~x68 & ~x71 & ~x72 & ~x73 & ~x81 & ~x83 & ~x85 & ~x86 & ~x91 & ~x93 & ~x95 & ~x97 & ~x102 & ~x104 & ~x105 & ~x107 & ~x109 & ~x112 & ~x129 & ~x131 & ~x133 & ~x135 & ~x136 & ~x139 & ~x143 & ~x158 & ~x159 & ~x160 & ~x161 & ~x164 & ~x170 & ~x188 & ~x190 & ~x191 & ~x192 & ~x196 & ~x198 & ~x199 & ~x217 & ~x218 & ~x221 & ~x223 & ~x224 & ~x244 & ~x245 & ~x246 & ~x249 & ~x250 & ~x271 & ~x272 & ~x274 & ~x276 & ~x277 & ~x281 & ~x282 & ~x299 & ~x301 & ~x302 & ~x307 & ~x327 & ~x332 & ~x335 & ~x338 & ~x339 & ~x360 & ~x361 & ~x362 & ~x365 & ~x390 & ~x391 & ~x393 & ~x394 & ~x395 & ~x415 & ~x416 & ~x417 & ~x423 & ~x424 & ~x425 & ~x446 & ~x449 & ~x450 & ~x454 & ~x455 & ~x456 & ~x475 & ~x476 & ~x478 & ~x479 & ~x484 & ~x485 & ~x486 & ~x487 & ~x489 & ~x504 & ~x506 & ~x509 & ~x510 & ~x512 & ~x531 & ~x533 & ~x534 & ~x540 & ~x556 & ~x557 & ~x560 & ~x585 & ~x586 & ~x588 & ~x592 & ~x612 & ~x615 & ~x617 & ~x618 & ~x621 & ~x645 & ~x646 & ~x648 & ~x651 & ~x671 & ~x675 & ~x692 & ~x693 & ~x696 & ~x697 & ~x699 & ~x700 & ~x705 & ~x722 & ~x727 & ~x728 & ~x729 & ~x736 & ~x739 & ~x740 & ~x741 & ~x742 & ~x744 & ~x745 & ~x747 & ~x750 & ~x754 & ~x755 & ~x756 & ~x757 & ~x758 & ~x760 & ~x765 & ~x766 & ~x768 & ~x769 & ~x772 & ~x774 & ~x775 & ~x777 & ~x781;
assign c3154 =  x323 &  x351 & ~x1 & ~x2 & ~x5 & ~x7 & ~x9 & ~x14 & ~x27 & ~x28 & ~x31 & ~x49 & ~x51 & ~x55 & ~x57 & ~x59 & ~x66 & ~x76 & ~x81 & ~x83 & ~x84 & ~x86 & ~x107 & ~x108 & ~x113 & ~x114 & ~x118 & ~x137 & ~x139 & ~x145 & ~x165 & ~x168 & ~x169 & ~x192 & ~x193 & ~x224 & ~x225 & ~x227 & ~x249 & ~x250 & ~x253 & ~x276 & ~x287 & ~x288 & ~x289 & ~x290 & ~x306 & ~x310 & ~x313 & ~x314 & ~x361 & ~x363 & ~x364 & ~x387 & ~x388 & ~x391 & ~x419 & ~x426 & ~x427 & ~x428 & ~x429 & ~x430 & ~x447 & ~x448 & ~x459 & ~x460 & ~x461 & ~x501 & ~x530 & ~x534 & ~x563 & ~x584 & ~x585 & ~x588 & ~x590 & ~x611 & ~x617 & ~x619 & ~x640 & ~x641 & ~x646 & ~x665 & ~x686 & ~x687 & ~x697 & ~x698 & ~x701 & ~x704 & ~x726 & ~x732 & ~x740 & ~x746 & ~x751 & ~x753 & ~x754 & ~x767 & ~x769 & ~x771 & ~x773 & ~x774 & ~x780;
assign c3156 =  x180 &  x404 & ~x0 & ~x4 & ~x8 & ~x9 & ~x13 & ~x24 & ~x31 & ~x36 & ~x49 & ~x51 & ~x57 & ~x65 & ~x72 & ~x78 & ~x82 & ~x91 & ~x94 & ~x99 & ~x101 & ~x117 & ~x136 & ~x173 & ~x192 & ~x194 & ~x196 & ~x220 & ~x225 & ~x248 & ~x256 & ~x276 & ~x278 & ~x280 & ~x286 & ~x291 & ~x303 & ~x305 & ~x313 & ~x342 & ~x394 & ~x419 & ~x420 & ~x444 & ~x446 & ~x476 & ~x483 & ~x503 & ~x512 & ~x563 & ~x582 & ~x583 & ~x585 & ~x589 & ~x590 & ~x610 & ~x611 & ~x612 & ~x615 & ~x640 & ~x669 & ~x671 & ~x692 & ~x702 & ~x720 & ~x742 & ~x749 & ~x756 & ~x767 & ~x782 & ~x783;
assign c3158 =  x183 & ~x56 & ~x222 & ~x292 & ~x302 & ~x317 & ~x332 & ~x468 & ~x543 & ~x544 & ~x545 & ~x664 & ~x772;
assign c3160 =  x174 &  x377 & ~x287;
assign c3162 =  x208 &  x234 &  x235 &  x236 &  x350 &  x377 &  x404 & ~x13 & ~x15 & ~x16 & ~x20 & ~x27 & ~x28 & ~x39 & ~x42 & ~x46 & ~x47 & ~x51 & ~x79 & ~x81 & ~x84 & ~x88 & ~x99 & ~x104 & ~x108 & ~x116 & ~x120 & ~x121 & ~x122 & ~x124 & ~x126 & ~x127 & ~x129 & ~x131 & ~x132 & ~x133 & ~x137 & ~x138 & ~x143 & ~x161 & ~x162 & ~x167 & ~x169 & ~x170 & ~x196 & ~x247 & ~x274 & ~x275 & ~x303 & ~x307 & ~x309 & ~x310 & ~x329 & ~x332 & ~x334 & ~x363 & ~x365 & ~x387 & ~x393 & ~x424 & ~x425 & ~x426 & ~x445 & ~x447 & ~x450 & ~x454 & ~x473 & ~x474 & ~x476 & ~x479 & ~x500 & ~x509 & ~x533 & ~x539 & ~x557 & ~x563 & ~x611 & ~x615 & ~x619 & ~x638 & ~x641 & ~x642 & ~x645 & ~x647 & ~x673 & ~x674 & ~x691 & ~x692 & ~x694 & ~x697 & ~x724 & ~x726 & ~x731 & ~x734 & ~x740 & ~x746 & ~x752 & ~x756 & ~x757 & ~x758 & ~x759 & ~x760 & ~x782;
assign c3164 = ~x7 & ~x34 & ~x43 & ~x45 & ~x54 & ~x80 & ~x96 & ~x105 & ~x111 & ~x114 & ~x134 & ~x191 & ~x278 & ~x292 & ~x344 & ~x397 & ~x398 & ~x445 & ~x542 & ~x545 & ~x546 & ~x560 & ~x571 & ~x573 & ~x575 & ~x599 & ~x746;
assign c3166 =  x326 &  x680 & ~x540 & ~x570;
assign c3168 =  x376 & ~x1 & ~x2 & ~x5 & ~x11 & ~x18 & ~x19 & ~x24 & ~x25 & ~x30 & ~x33 & ~x48 & ~x66 & ~x70 & ~x79 & ~x81 & ~x84 & ~x88 & ~x89 & ~x90 & ~x105 & ~x107 & ~x133 & ~x139 & ~x147 & ~x163 & ~x192 & ~x219 & ~x222 & ~x224 & ~x247 & ~x249 & ~x252 & ~x277 & ~x289 & ~x290 & ~x291 & ~x303 & ~x306 & ~x315 & ~x337 & ~x339 & ~x362 & ~x363 & ~x364 & ~x368 & ~x390 & ~x393 & ~x419 & ~x422 & ~x444 & ~x447 & ~x449 & ~x454 & ~x456 & ~x457 & ~x459 & ~x460 & ~x474 & ~x478 & ~x506 & ~x507 & ~x558 & ~x563 & ~x587 & ~x612 & ~x613 & ~x620 & ~x640 & ~x642 & ~x643 & ~x648 & ~x666 & ~x674 & ~x675 & ~x677 & ~x692 & ~x693 & ~x694 & ~x697 & ~x703 & ~x719 & ~x738 & ~x745 & ~x746 & ~x747 & ~x749 & ~x751 & ~x752 & ~x753 & ~x756 & ~x760 & ~x762 & ~x763 & ~x767 & ~x769 & ~x771 & ~x772 & ~x781;
assign c3170 =  x478;
assign c3172 =  x293 & ~x100 & ~x158 & ~x187 & ~x216 & ~x260 & ~x270 & ~x286 & ~x429 & ~x490;
assign c3174 =  x31;
assign c3176 =  x209 &  x235 &  x379 &  x406 &  x549 & ~x55 & ~x127 & ~x320 & ~x345 & ~x346;
assign c3178 =  x377 & ~x0 & ~x5 & ~x10 & ~x11 & ~x14 & ~x18 & ~x19 & ~x21 & ~x26 & ~x28 & ~x31 & ~x33 & ~x34 & ~x36 & ~x38 & ~x39 & ~x40 & ~x41 & ~x42 & ~x43 & ~x47 & ~x48 & ~x51 & ~x52 & ~x59 & ~x60 & ~x62 & ~x67 & ~x69 & ~x71 & ~x73 & ~x74 & ~x76 & ~x77 & ~x78 & ~x80 & ~x82 & ~x83 & ~x89 & ~x96 & ~x98 & ~x100 & ~x104 & ~x105 & ~x106 & ~x107 & ~x109 & ~x115 & ~x117 & ~x118 & ~x119 & ~x133 & ~x136 & ~x137 & ~x143 & ~x163 & ~x164 & ~x165 & ~x166 & ~x169 & ~x172 & ~x192 & ~x193 & ~x196 & ~x197 & ~x221 & ~x223 & ~x226 & ~x248 & ~x250 & ~x252 & ~x265 & ~x275 & ~x277 & ~x278 & ~x279 & ~x289 & ~x290 & ~x303 & ~x304 & ~x306 & ~x307 & ~x309 & ~x312 & ~x313 & ~x331 & ~x333 & ~x337 & ~x339 & ~x360 & ~x361 & ~x364 & ~x387 & ~x389 & ~x390 & ~x392 & ~x417 & ~x418 & ~x420 & ~x421 & ~x422 & ~x444 & ~x446 & ~x450 & ~x472 & ~x473 & ~x474 & ~x476 & ~x477 & ~x479 & ~x482 & ~x485 & ~x487 & ~x488 & ~x500 & ~x505 & ~x534 & ~x556 & ~x557 & ~x558 & ~x559 & ~x561 & ~x562 & ~x584 & ~x585 & ~x586 & ~x587 & ~x588 & ~x612 & ~x616 & ~x618 & ~x639 & ~x644 & ~x645 & ~x646 & ~x665 & ~x666 & ~x673 & ~x674 & ~x690 & ~x691 & ~x697 & ~x699 & ~x702 & ~x704 & ~x716 & ~x722 & ~x726 & ~x730 & ~x731 & ~x732 & ~x735 & ~x736 & ~x739 & ~x740 & ~x744 & ~x749 & ~x754 & ~x757 & ~x761 & ~x763 & ~x766 & ~x767 & ~x768 & ~x770 & ~x776 & ~x777 & ~x781 & ~x782 & ~x783;
assign c3180 =  x297 &  x325 &  x495 &  x570 & ~x6 & ~x11 & ~x64 & ~x76 & ~x85 & ~x109 & ~x119 & ~x170 & ~x197 & ~x201 & ~x334 & ~x338 & ~x359 & ~x463 & ~x500 & ~x530 & ~x532 & ~x558 & ~x588 & ~x665 & ~x679 & ~x704 & ~x715 & ~x730 & ~x738 & ~x760 & ~x769 & ~x770;
assign c3182 =  x213 &  x214 &  x380 &  x602 & ~x0 & ~x4 & ~x5 & ~x11 & ~x28 & ~x29 & ~x41 & ~x76 & ~x79 & ~x82 & ~x112 & ~x135 & ~x144 & ~x147 & ~x168 & ~x192 & ~x221 & ~x247 & ~x257 & ~x279 & ~x304 & ~x306 & ~x310 & ~x335 & ~x338 & ~x341 & ~x387 & ~x389 & ~x399 & ~x416 & ~x417 & ~x443 & ~x456 & ~x527 & ~x558 & ~x582 & ~x611 & ~x613 & ~x617 & ~x643 & ~x645 & ~x664 & ~x670 & ~x671 & ~x673 & ~x675 & ~x688 & ~x696 & ~x714 & ~x725 & ~x728 & ~x740 & ~x741 & ~x750 & ~x754 & ~x768;
assign c3184 =  x631 & ~x2 & ~x3 & ~x9 & ~x14 & ~x16 & ~x20 & ~x22 & ~x31 & ~x34 & ~x36 & ~x39 & ~x44 & ~x53 & ~x59 & ~x61 & ~x72 & ~x77 & ~x79 & ~x80 & ~x88 & ~x89 & ~x94 & ~x109 & ~x119 & ~x120 & ~x135 & ~x140 & ~x144 & ~x171 & ~x194 & ~x202 & ~x203 & ~x222 & ~x224 & ~x230 & ~x277 & ~x278 & ~x283 & ~x293 & ~x294 & ~x307 & ~x310 & ~x313 & ~x317 & ~x319 & ~x337 & ~x339 & ~x343 & ~x359 & ~x363 & ~x364 & ~x368 & ~x396 & ~x444 & ~x451 & ~x469 & ~x472 & ~x475 & ~x479 & ~x480 & ~x503 & ~x504 & ~x527 & ~x535 & ~x553 & ~x561 & ~x583 & ~x587 & ~x590 & ~x591 & ~x608 & ~x618 & ~x635 & ~x646 & ~x647 & ~x662 & ~x664 & ~x669 & ~x675 & ~x696 & ~x700 & ~x704 & ~x714 & ~x718 & ~x723 & ~x725 & ~x726 & ~x728 & ~x741 & ~x762 & ~x766 & ~x769 & ~x770 & ~x782 & ~x783;
assign c3186 =  x298 & ~x2 & ~x5 & ~x8 & ~x9 & ~x16 & ~x17 & ~x18 & ~x21 & ~x22 & ~x23 & ~x24 & ~x28 & ~x30 & ~x33 & ~x35 & ~x36 & ~x38 & ~x41 & ~x42 & ~x44 & ~x45 & ~x49 & ~x50 & ~x52 & ~x54 & ~x59 & ~x60 & ~x63 & ~x64 & ~x66 & ~x70 & ~x73 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x88 & ~x91 & ~x94 & ~x106 & ~x108 & ~x110 & ~x111 & ~x112 & ~x113 & ~x114 & ~x117 & ~x119 & ~x134 & ~x135 & ~x136 & ~x137 & ~x139 & ~x141 & ~x143 & ~x144 & ~x145 & ~x164 & ~x167 & ~x168 & ~x192 & ~x193 & ~x194 & ~x196 & ~x197 & ~x198 & ~x220 & ~x224 & ~x225 & ~x226 & ~x247 & ~x250 & ~x255 & ~x276 & ~x277 & ~x280 & ~x287 & ~x288 & ~x303 & ~x304 & ~x308 & ~x309 & ~x312 & ~x314 & ~x315 & ~x331 & ~x334 & ~x337 & ~x342 & ~x343 & ~x359 & ~x361 & ~x367 & ~x368 & ~x369 & ~x370 & ~x387 & ~x388 & ~x392 & ~x393 & ~x394 & ~x396 & ~x397 & ~x416 & ~x418 & ~x421 & ~x422 & ~x424 & ~x443 & ~x448 & ~x455 & ~x471 & ~x476 & ~x479 & ~x485 & ~x486 & ~x502 & ~x504 & ~x515 & ~x528 & ~x531 & ~x534 & ~x556 & ~x558 & ~x559 & ~x560 & ~x561 & ~x583 & ~x585 & ~x587 & ~x588 & ~x589 & ~x590 & ~x591 & ~x615 & ~x616 & ~x617 & ~x618 & ~x638 & ~x642 & ~x645 & ~x646 & ~x664 & ~x665 & ~x668 & ~x670 & ~x671 & ~x673 & ~x674 & ~x691 & ~x692 & ~x694 & ~x697 & ~x699 & ~x700 & ~x701 & ~x705 & ~x707 & ~x708 & ~x709 & ~x710 & ~x712 & ~x713 & ~x714 & ~x715 & ~x716 & ~x718 & ~x721 & ~x724 & ~x725 & ~x726 & ~x729 & ~x730 & ~x735 & ~x737 & ~x738 & ~x739 & ~x744 & ~x745 & ~x746 & ~x747 & ~x752 & ~x757 & ~x759 & ~x760 & ~x761 & ~x762 & ~x763 & ~x765 & ~x766 & ~x767 & ~x768 & ~x769 & ~x773 & ~x777 & ~x779;
assign c3188 =  x699;
assign c3190 =  x552 & ~x44 & ~x73 & ~x128 & ~x186 & ~x215 & ~x300 & ~x308 & ~x328 & ~x485 & ~x509 & ~x538 & ~x556 & ~x623 & ~x726 & ~x739 & ~x751;
assign c3192 =  x152 & ~x14 & ~x42 & ~x48 & ~x50 & ~x66 & ~x71 & ~x98 & ~x108 & ~x111 & ~x162 & ~x224 & ~x235 & ~x260 & ~x261 & ~x262 & ~x286 & ~x330 & ~x331 & ~x423 & ~x452 & ~x458 & ~x459 & ~x500 & ~x518 & ~x590 & ~x611 & ~x615 & ~x668 & ~x690 & ~x710 & ~x743 & ~x754 & ~x759 & ~x771 & ~x775;
assign c3194 =  x479;
assign c3196 =  x403 &  x404 & ~x4 & ~x11 & ~x13 & ~x14 & ~x20 & ~x21 & ~x22 & ~x28 & ~x29 & ~x30 & ~x32 & ~x37 & ~x39 & ~x56 & ~x60 & ~x66 & ~x75 & ~x79 & ~x80 & ~x85 & ~x87 & ~x94 & ~x97 & ~x100 & ~x102 & ~x105 & ~x110 & ~x112 & ~x114 & ~x116 & ~x131 & ~x134 & ~x141 & ~x145 & ~x167 & ~x171 & ~x172 & ~x196 & ~x197 & ~x221 & ~x249 & ~x250 & ~x276 & ~x279 & ~x292 & ~x304 & ~x309 & ~x314 & ~x317 & ~x319 & ~x332 & ~x333 & ~x337 & ~x338 & ~x339 & ~x340 & ~x344 & ~x366 & ~x369 & ~x391 & ~x415 & ~x418 & ~x419 & ~x421 & ~x424 & ~x445 & ~x453 & ~x472 & ~x474 & ~x475 & ~x478 & ~x500 & ~x501 & ~x511 & ~x528 & ~x533 & ~x557 & ~x560 & ~x589 & ~x617 & ~x638 & ~x639 & ~x640 & ~x642 & ~x645 & ~x667 & ~x668 & ~x691 & ~x693 & ~x694 & ~x695 & ~x703 & ~x714 & ~x715 & ~x716 & ~x722 & ~x723 & ~x724 & ~x727 & ~x740 & ~x741 & ~x743 & ~x746 & ~x748 & ~x752 & ~x756 & ~x757 & ~x763 & ~x764 & ~x765 & ~x766 & ~x767 & ~x774 & ~x776 & ~x782;
assign c3198 =  x146;
assign c3200 =  x731;
assign c3202 =  x208 & ~x7 & ~x29 & ~x38 & ~x42 & ~x46 & ~x47 & ~x74 & ~x78 & ~x83 & ~x93 & ~x106 & ~x130 & ~x157 & ~x159 & ~x166 & ~x167 & ~x252 & ~x273 & ~x276 & ~x301 & ~x331 & ~x336 & ~x343 & ~x371 & ~x384 & ~x423 & ~x444 & ~x510 & ~x539 & ~x540 & ~x546 & ~x547 & ~x560 & ~x561 & ~x584 & ~x586 & ~x590 & ~x600 & ~x614 & ~x653 & ~x702 & ~x709 & ~x723 & ~x725 & ~x750 & ~x756 & ~x764 & ~x773;
assign c3204 =  x21;
assign c3206 =  x772;
assign c3208 =  x267 &  x294 &  x348 &  x377 &  x469 & ~x133 & ~x302;
assign c3210 =  x754;
assign c3212 =  x646;
assign c3214 =  x39;
assign c3218 =  x56;
assign c3220 =  x27;
assign c3222 =  x207 &  x208 & ~x0 & ~x5 & ~x7 & ~x8 & ~x10 & ~x11 & ~x17 & ~x19 & ~x23 & ~x25 & ~x27 & ~x34 & ~x35 & ~x39 & ~x40 & ~x43 & ~x44 & ~x50 & ~x60 & ~x67 & ~x68 & ~x70 & ~x93 & ~x103 & ~x112 & ~x117 & ~x119 & ~x123 & ~x127 & ~x141 & ~x142 & ~x159 & ~x162 & ~x163 & ~x168 & ~x171 & ~x197 & ~x220 & ~x221 & ~x222 & ~x223 & ~x252 & ~x289 & ~x290 & ~x309 & ~x315 & ~x334 & ~x335 & ~x336 & ~x338 & ~x339 & ~x361 & ~x362 & ~x363 & ~x391 & ~x393 & ~x396 & ~x397 & ~x425 & ~x445 & ~x475 & ~x476 & ~x478 & ~x491 & ~x502 & ~x507 & ~x520 & ~x528 & ~x530 & ~x531 & ~x533 & ~x562 & ~x563 & ~x584 & ~x614 & ~x615 & ~x638 & ~x639 & ~x640 & ~x644 & ~x645 & ~x646 & ~x649 & ~x667 & ~x670 & ~x673 & ~x674 & ~x695 & ~x700 & ~x724 & ~x728 & ~x730 & ~x731 & ~x732 & ~x743 & ~x745 & ~x747 & ~x749 & ~x752 & ~x756 & ~x762 & ~x765 & ~x766 & ~x768 & ~x769 & ~x770 & ~x779;
assign c3224 =  x676;
assign c3226 =  x181 &  x182 &  x268 &  x295 &  x321 &  x348 & ~x1 & ~x2 & ~x8 & ~x15 & ~x26 & ~x32 & ~x53 & ~x58 & ~x63 & ~x66 & ~x68 & ~x73 & ~x75 & ~x77 & ~x78 & ~x81 & ~x82 & ~x86 & ~x92 & ~x96 & ~x104 & ~x106 & ~x108 & ~x112 & ~x114 & ~x136 & ~x138 & ~x140 & ~x141 & ~x164 & ~x168 & ~x171 & ~x191 & ~x193 & ~x194 & ~x199 & ~x226 & ~x247 & ~x249 & ~x250 & ~x251 & ~x282 & ~x284 & ~x304 & ~x311 & ~x329 & ~x332 & ~x334 & ~x338 & ~x360 & ~x387 & ~x388 & ~x391 & ~x393 & ~x394 & ~x416 & ~x420 & ~x446 & ~x476 & ~x477 & ~x478 & ~x479 & ~x488 & ~x506 & ~x530 & ~x531 & ~x533 & ~x558 & ~x559 & ~x586 & ~x588 & ~x613 & ~x615 & ~x646 & ~x667 & ~x670 & ~x672 & ~x676 & ~x696 & ~x701 & ~x717 & ~x718 & ~x720 & ~x721 & ~x722 & ~x734 & ~x741 & ~x755 & ~x756 & ~x758 & ~x762 & ~x764 & ~x771 & ~x776 & ~x778 & ~x779 & ~x780 & ~x781;
assign c3228 =  x421;
assign c3230 = ~x2 & ~x8 & ~x19 & ~x33 & ~x39 & ~x43 & ~x48 & ~x50 & ~x53 & ~x56 & ~x74 & ~x94 & ~x105 & ~x106 & ~x114 & ~x115 & ~x131 & ~x137 & ~x162 & ~x166 & ~x168 & ~x188 & ~x190 & ~x191 & ~x217 & ~x219 & ~x220 & ~x222 & ~x224 & ~x253 & ~x263 & ~x305 & ~x317 & ~x333 & ~x342 & ~x360 & ~x367 & ~x368 & ~x369 & ~x388 & ~x415 & ~x416 & ~x422 & ~x424 & ~x444 & ~x450 & ~x452 & ~x472 & ~x482 & ~x507 & ~x532 & ~x535 & ~x543 & ~x545 & ~x562 & ~x573 & ~x574 & ~x575 & ~x586 & ~x587 & ~x588 & ~x589 & ~x613 & ~x617 & ~x730 & ~x739 & ~x741 & ~x763 & ~x766 & ~x768 & ~x776;
assign c3232 =  x150 &  x319 & ~x232 & ~x233 & ~x273 & ~x454 & ~x704;
assign c3234 =  x143;
assign c3236 =  x209 &  x210 &  x211 &  x296 &  x350 &  x377 & ~x2 & ~x5 & ~x6 & ~x7 & ~x8 & ~x10 & ~x12 & ~x20 & ~x25 & ~x26 & ~x27 & ~x28 & ~x31 & ~x33 & ~x34 & ~x35 & ~x37 & ~x38 & ~x39 & ~x41 & ~x44 & ~x45 & ~x47 & ~x48 & ~x49 & ~x51 & ~x54 & ~x55 & ~x59 & ~x61 & ~x62 & ~x65 & ~x67 & ~x71 & ~x72 & ~x74 & ~x76 & ~x77 & ~x81 & ~x82 & ~x84 & ~x86 & ~x91 & ~x92 & ~x93 & ~x101 & ~x106 & ~x108 & ~x110 & ~x112 & ~x113 & ~x117 & ~x118 & ~x124 & ~x126 & ~x134 & ~x138 & ~x140 & ~x141 & ~x145 & ~x163 & ~x164 & ~x165 & ~x171 & ~x189 & ~x190 & ~x193 & ~x196 & ~x197 & ~x198 & ~x199 & ~x219 & ~x221 & ~x223 & ~x226 & ~x228 & ~x246 & ~x274 & ~x277 & ~x279 & ~x280 & ~x301 & ~x305 & ~x306 & ~x309 & ~x312 & ~x330 & ~x331 & ~x337 & ~x339 & ~x357 & ~x361 & ~x364 & ~x365 & ~x366 & ~x367 & ~x368 & ~x369 & ~x386 & ~x387 & ~x390 & ~x392 & ~x393 & ~x394 & ~x395 & ~x396 & ~x399 & ~x415 & ~x416 & ~x419 & ~x424 & ~x445 & ~x446 & ~x447 & ~x448 & ~x453 & ~x471 & ~x472 & ~x477 & ~x481 & ~x482 & ~x499 & ~x500 & ~x505 & ~x506 & ~x507 & ~x528 & ~x530 & ~x532 & ~x533 & ~x535 & ~x536 & ~x555 & ~x558 & ~x560 & ~x561 & ~x563 & ~x583 & ~x584 & ~x586 & ~x587 & ~x588 & ~x589 & ~x590 & ~x591 & ~x610 & ~x611 & ~x613 & ~x614 & ~x615 & ~x616 & ~x620 & ~x639 & ~x640 & ~x643 & ~x645 & ~x647 & ~x666 & ~x669 & ~x673 & ~x674 & ~x675 & ~x692 & ~x693 & ~x694 & ~x701 & ~x703 & ~x706 & ~x715 & ~x717 & ~x719 & ~x722 & ~x723 & ~x726 & ~x729 & ~x734 & ~x735 & ~x737 & ~x738 & ~x741 & ~x743 & ~x746 & ~x748 & ~x750 & ~x753 & ~x756 & ~x757 & ~x759 & ~x761 & ~x762 & ~x763 & ~x770 & ~x771 & ~x777 & ~x778 & ~x780;
assign c3238 =  x140;
assign c3240 = ~x3 & ~x9 & ~x10 & ~x12 & ~x24 & ~x63 & ~x79 & ~x83 & ~x88 & ~x95 & ~x96 & ~x101 & ~x115 & ~x140 & ~x143 & ~x222 & ~x318 & ~x319 & ~x338 & ~x344 & ~x358 & ~x366 & ~x370 & ~x387 & ~x415 & ~x445 & ~x447 & ~x449 & ~x452 & ~x475 & ~x502 & ~x504 & ~x505 & ~x506 & ~x510 & ~x541 & ~x543 & ~x557 & ~x563 & ~x574 & ~x584 & ~x587 & ~x601 & ~x614 & ~x665 & ~x694 & ~x700 & ~x706 & ~x723 & ~x735 & ~x744 & ~x746 & ~x757;
assign c3242 =  x181 &  x240 & ~x6 & ~x10 & ~x11 & ~x12 & ~x14 & ~x17 & ~x28 & ~x34 & ~x35 & ~x39 & ~x40 & ~x43 & ~x49 & ~x52 & ~x58 & ~x63 & ~x67 & ~x68 & ~x72 & ~x75 & ~x76 & ~x79 & ~x81 & ~x87 & ~x93 & ~x94 & ~x98 & ~x101 & ~x104 & ~x110 & ~x111 & ~x117 & ~x131 & ~x133 & ~x138 & ~x139 & ~x140 & ~x142 & ~x145 & ~x146 & ~x162 & ~x164 & ~x166 & ~x167 & ~x168 & ~x173 & ~x188 & ~x190 & ~x191 & ~x192 & ~x195 & ~x196 & ~x201 & ~x216 & ~x218 & ~x219 & ~x220 & ~x224 & ~x228 & ~x247 & ~x251 & ~x277 & ~x281 & ~x282 & ~x302 & ~x339 & ~x361 & ~x368 & ~x369 & ~x394 & ~x396 & ~x415 & ~x416 & ~x425 & ~x445 & ~x449 & ~x454 & ~x472 & ~x476 & ~x500 & ~x501 & ~x504 & ~x508 & ~x509 & ~x529 & ~x533 & ~x534 & ~x536 & ~x544 & ~x545 & ~x554 & ~x583 & ~x585 & ~x586 & ~x612 & ~x614 & ~x615 & ~x621 & ~x637 & ~x638 & ~x648 & ~x665 & ~x670 & ~x673 & ~x674 & ~x675 & ~x697 & ~x705 & ~x727 & ~x736 & ~x745 & ~x750 & ~x757 & ~x759 & ~x764 & ~x772 & ~x777 & ~x781;
assign c3244 = ~x11 & ~x19 & ~x28 & ~x32 & ~x35 & ~x39 & ~x43 & ~x47 & ~x49 & ~x57 & ~x59 & ~x61 & ~x67 & ~x71 & ~x78 & ~x81 & ~x82 & ~x83 & ~x84 & ~x91 & ~x92 & ~x93 & ~x97 & ~x99 & ~x106 & ~x107 & ~x110 & ~x120 & ~x127 & ~x129 & ~x131 & ~x132 & ~x135 & ~x138 & ~x144 & ~x164 & ~x166 & ~x170 & ~x174 & ~x192 & ~x194 & ~x196 & ~x198 & ~x200 & ~x221 & ~x223 & ~x225 & ~x251 & ~x276 & ~x277 & ~x281 & ~x308 & ~x320 & ~x339 & ~x340 & ~x346 & ~x359 & ~x363 & ~x369 & ~x370 & ~x371 & ~x373 & ~x386 & ~x387 & ~x390 & ~x395 & ~x398 & ~x400 & ~x444 & ~x448 & ~x450 & ~x452 & ~x475 & ~x501 & ~x505 & ~x506 & ~x507 & ~x513 & ~x514 & ~x515 & ~x529 & ~x535 & ~x541 & ~x544 & ~x546 & ~x559 & ~x562 & ~x563 & ~x571 & ~x572 & ~x584 & ~x611 & ~x614 & ~x638 & ~x643 & ~x644 & ~x645 & ~x673 & ~x675 & ~x694 & ~x696 & ~x700 & ~x701 & ~x717 & ~x724 & ~x729 & ~x731 & ~x732 & ~x742 & ~x752 & ~x757 & ~x764 & ~x772 & ~x773 & ~x779 & ~x782;
assign c3246 =  x199;
assign c3248 =  x563;
assign c3250 =  x351 &  x352 &  x379 &  x405 &  x494 &  x522 & ~x8 & ~x13 & ~x15 & ~x22 & ~x28 & ~x34 & ~x37 & ~x38 & ~x42 & ~x44 & ~x46 & ~x50 & ~x59 & ~x67 & ~x73 & ~x74 & ~x86 & ~x87 & ~x90 & ~x93 & ~x94 & ~x96 & ~x98 & ~x103 & ~x104 & ~x107 & ~x113 & ~x137 & ~x140 & ~x141 & ~x147 & ~x171 & ~x172 & ~x194 & ~x221 & ~x227 & ~x248 & ~x252 & ~x253 & ~x281 & ~x319 & ~x332 & ~x334 & ~x339 & ~x345 & ~x359 & ~x370 & ~x386 & ~x387 & ~x388 & ~x390 & ~x391 & ~x393 & ~x398 & ~x416 & ~x420 & ~x471 & ~x501 & ~x503 & ~x526 & ~x554 & ~x555 & ~x582 & ~x585 & ~x588 & ~x590 & ~x615 & ~x616 & ~x617 & ~x638 & ~x642 & ~x643 & ~x672 & ~x696 & ~x700 & ~x703 & ~x704 & ~x706 & ~x707 & ~x724 & ~x725 & ~x726 & ~x729 & ~x731 & ~x748 & ~x752 & ~x754 & ~x760 & ~x769 & ~x770 & ~x775 & ~x780 & ~x783;
assign c3252 =  x762;
assign c3254 =  x605 & ~x16 & ~x69 & ~x80 & ~x96 & ~x108 & ~x156 & ~x217 & ~x278 & ~x287 & ~x289 & ~x368 & ~x446 & ~x492 & ~x557 & ~x584 & ~x703 & ~x742 & ~x757;
assign c3256 =  x627 & ~x4 & ~x8 & ~x9 & ~x14 & ~x15 & ~x33 & ~x34 & ~x39 & ~x42 & ~x46 & ~x50 & ~x59 & ~x61 & ~x78 & ~x80 & ~x89 & ~x117 & ~x118 & ~x134 & ~x139 & ~x142 & ~x172 & ~x195 & ~x199 & ~x219 & ~x232 & ~x247 & ~x251 & ~x257 & ~x262 & ~x263 & ~x265 & ~x279 & ~x302 & ~x303 & ~x304 & ~x309 & ~x312 & ~x336 & ~x340 & ~x361 & ~x387 & ~x394 & ~x395 & ~x396 & ~x397 & ~x418 & ~x425 & ~x442 & ~x453 & ~x469 & ~x505 & ~x525 & ~x536 & ~x553 & ~x559 & ~x582 & ~x586 & ~x590 & ~x609 & ~x610 & ~x619 & ~x634 & ~x641 & ~x642 & ~x663 & ~x665 & ~x667 & ~x684 & ~x685 & ~x689 & ~x691 & ~x695 & ~x702 & ~x710 & ~x718 & ~x723 & ~x725 & ~x734 & ~x739 & ~x740 & ~x744 & ~x749 & ~x752 & ~x758 & ~x764 & ~x766 & ~x778 & ~x779 & ~x781;
assign c3258 =  x652 & ~x1 & ~x3 & ~x4 & ~x11 & ~x14 & ~x31 & ~x33 & ~x38 & ~x41 & ~x46 & ~x55 & ~x56 & ~x63 & ~x68 & ~x75 & ~x80 & ~x99 & ~x116 & ~x133 & ~x138 & ~x139 & ~x140 & ~x145 & ~x161 & ~x164 & ~x168 & ~x174 & ~x192 & ~x201 & ~x248 & ~x283 & ~x342 & ~x363 & ~x372 & ~x387 & ~x424 & ~x451 & ~x480 & ~x483 & ~x484 & ~x503 & ~x514 & ~x542 & ~x572 & ~x581 & ~x584 & ~x636 & ~x642 & ~x663 & ~x664 & ~x672 & ~x691 & ~x693 & ~x695 & ~x735 & ~x738 & ~x748 & ~x750 & ~x758 & ~x771;
assign c3260 =  x476;
assign c3262 =  x478;
assign c3264 =  x178 &  x321 &  x347 &  x375 &  x376 & ~x484 & ~x486;
assign c3266 =  x673;
assign c3268 =  x268 &  x295 &  x321 & ~x4 & ~x11 & ~x12 & ~x13 & ~x15 & ~x16 & ~x17 & ~x18 & ~x19 & ~x24 & ~x32 & ~x37 & ~x38 & ~x39 & ~x41 & ~x42 & ~x43 & ~x44 & ~x45 & ~x47 & ~x48 & ~x49 & ~x51 & ~x53 & ~x59 & ~x64 & ~x72 & ~x74 & ~x75 & ~x77 & ~x87 & ~x90 & ~x92 & ~x102 & ~x116 & ~x132 & ~x133 & ~x134 & ~x136 & ~x143 & ~x144 & ~x161 & ~x162 & ~x163 & ~x167 & ~x189 & ~x200 & ~x201 & ~x217 & ~x218 & ~x226 & ~x244 & ~x245 & ~x248 & ~x250 & ~x254 & ~x255 & ~x256 & ~x273 & ~x275 & ~x277 & ~x283 & ~x299 & ~x301 & ~x303 & ~x304 & ~x310 & ~x329 & ~x330 & ~x336 & ~x359 & ~x360 & ~x362 & ~x363 & ~x364 & ~x365 & ~x366 & ~x390 & ~x395 & ~x396 & ~x420 & ~x424 & ~x444 & ~x448 & ~x451 & ~x452 & ~x481 & ~x482 & ~x501 & ~x529 & ~x530 & ~x532 & ~x533 & ~x534 & ~x557 & ~x562 & ~x564 & ~x584 & ~x586 & ~x617 & ~x621 & ~x636 & ~x637 & ~x641 & ~x643 & ~x644 & ~x645 & ~x662 & ~x663 & ~x668 & ~x675 & ~x676 & ~x677 & ~x687 & ~x689 & ~x696 & ~x698 & ~x703 & ~x704 & ~x705 & ~x725 & ~x726 & ~x727 & ~x730 & ~x737 & ~x739 & ~x743 & ~x754 & ~x758 & ~x766 & ~x768 & ~x770 & ~x771 & ~x776 & ~x778 & ~x781;
assign c3270 =  x300 &  x380 & ~x36 & ~x91 & ~x196 & ~x331 & ~x333 & ~x484 & ~x485 & ~x486 & ~x487 & ~x527 & ~x553 & ~x607 & ~x614 & ~x617 & ~x635;
assign c3272 =  x185 &  x186 &  x298 &  x352 &  x378 &  x379 &  x575 &  x602 &  x627 & ~x3 & ~x24 & ~x25 & ~x43 & ~x52 & ~x57 & ~x71 & ~x81 & ~x85 & ~x106 & ~x109 & ~x114 & ~x122 & ~x136 & ~x137 & ~x138 & ~x142 & ~x165 & ~x191 & ~x194 & ~x200 & ~x201 & ~x222 & ~x226 & ~x252 & ~x276 & ~x285 & ~x303 & ~x304 & ~x310 & ~x313 & ~x333 & ~x334 & ~x358 & ~x359 & ~x362 & ~x365 & ~x369 & ~x390 & ~x391 & ~x393 & ~x416 & ~x417 & ~x443 & ~x446 & ~x449 & ~x450 & ~x473 & ~x478 & ~x500 & ~x504 & ~x526 & ~x535 & ~x555 & ~x558 & ~x559 & ~x560 & ~x582 & ~x583 & ~x586 & ~x588 & ~x613 & ~x617 & ~x637 & ~x640 & ~x643 & ~x644 & ~x645 & ~x663 & ~x668 & ~x694 & ~x695 & ~x702 & ~x712 & ~x714 & ~x724 & ~x730 & ~x741 & ~x748 & ~x752 & ~x755 & ~x756 & ~x761 & ~x772 & ~x773 & ~x778 & ~x780;
assign c3274 =  x244 &  x271 &  x299 &  x325 &  x351 &  x352 &  x599 & ~x0 & ~x8 & ~x16 & ~x19 & ~x26 & ~x27 & ~x35 & ~x37 & ~x39 & ~x41 & ~x46 & ~x49 & ~x69 & ~x74 & ~x86 & ~x106 & ~x110 & ~x113 & ~x118 & ~x138 & ~x143 & ~x194 & ~x222 & ~x248 & ~x280 & ~x304 & ~x334 & ~x364 & ~x366 & ~x388 & ~x392 & ~x394 & ~x415 & ~x445 & ~x449 & ~x475 & ~x478 & ~x502 & ~x506 & ~x531 & ~x557 & ~x608 & ~x612 & ~x616 & ~x645 & ~x668 & ~x674 & ~x676 & ~x701 & ~x711 & ~x714 & ~x715 & ~x723 & ~x727 & ~x729 & ~x740 & ~x759 & ~x766 & ~x770 & ~x775 & ~x779 & ~x783;
assign c3276 =  x629 & ~x2 & ~x4 & ~x6 & ~x10 & ~x14 & ~x17 & ~x19 & ~x22 & ~x28 & ~x31 & ~x43 & ~x46 & ~x50 & ~x52 & ~x59 & ~x67 & ~x72 & ~x75 & ~x80 & ~x82 & ~x83 & ~x91 & ~x101 & ~x103 & ~x105 & ~x136 & ~x143 & ~x157 & ~x161 & ~x167 & ~x188 & ~x198 & ~x218 & ~x219 & ~x220 & ~x249 & ~x252 & ~x283 & ~x305 & ~x306 & ~x331 & ~x334 & ~x336 & ~x358 & ~x362 & ~x364 & ~x366 & ~x387 & ~x389 & ~x398 & ~x399 & ~x402 & ~x418 & ~x422 & ~x423 & ~x444 & ~x445 & ~x459 & ~x472 & ~x474 & ~x475 & ~x476 & ~x477 & ~x489 & ~x500 & ~x503 & ~x504 & ~x516 & ~x517 & ~x518 & ~x531 & ~x532 & ~x562 & ~x585 & ~x588 & ~x612 & ~x638 & ~x641 & ~x643 & ~x644 & ~x646 & ~x648 & ~x665 & ~x666 & ~x668 & ~x671 & ~x703 & ~x724 & ~x730 & ~x732 & ~x734 & ~x742 & ~x749 & ~x754 & ~x758 & ~x761 & ~x764 & ~x769 & ~x774 & ~x777 & ~x778 & ~x780 & ~x782 & ~x783;
assign c3278 =  x185 & ~x0 & ~x1 & ~x2 & ~x3 & ~x6 & ~x7 & ~x16 & ~x22 & ~x24 & ~x31 & ~x38 & ~x40 & ~x41 & ~x43 & ~x47 & ~x50 & ~x51 & ~x53 & ~x55 & ~x56 & ~x58 & ~x61 & ~x62 & ~x64 & ~x70 & ~x71 & ~x72 & ~x73 & ~x74 & ~x75 & ~x77 & ~x78 & ~x79 & ~x82 & ~x85 & ~x89 & ~x90 & ~x91 & ~x92 & ~x94 & ~x97 & ~x98 & ~x99 & ~x101 & ~x102 & ~x103 & ~x104 & ~x107 & ~x109 & ~x114 & ~x117 & ~x120 & ~x130 & ~x131 & ~x132 & ~x134 & ~x135 & ~x136 & ~x141 & ~x144 & ~x145 & ~x163 & ~x164 & ~x167 & ~x172 & ~x174 & ~x191 & ~x192 & ~x193 & ~x194 & ~x197 & ~x201 & ~x223 & ~x225 & ~x226 & ~x227 & ~x229 & ~x253 & ~x277 & ~x279 & ~x281 & ~x282 & ~x283 & ~x304 & ~x309 & ~x312 & ~x332 & ~x333 & ~x335 & ~x339 & ~x362 & ~x363 & ~x364 & ~x366 & ~x368 & ~x369 & ~x370 & ~x372 & ~x392 & ~x393 & ~x395 & ~x414 & ~x417 & ~x420 & ~x422 & ~x424 & ~x444 & ~x451 & ~x470 & ~x472 & ~x474 & ~x476 & ~x478 & ~x479 & ~x499 & ~x501 & ~x502 & ~x503 & ~x505 & ~x510 & ~x511 & ~x513 & ~x529 & ~x542 & ~x544 & ~x559 & ~x560 & ~x583 & ~x586 & ~x610 & ~x611 & ~x613 & ~x615 & ~x641 & ~x643 & ~x645 & ~x664 & ~x668 & ~x670 & ~x671 & ~x672 & ~x673 & ~x689 & ~x690 & ~x691 & ~x693 & ~x695 & ~x696 & ~x698 & ~x700 & ~x702 & ~x713 & ~x715 & ~x721 & ~x726 & ~x728 & ~x732 & ~x734 & ~x736 & ~x737 & ~x738 & ~x742 & ~x745 & ~x747 & ~x750 & ~x754 & ~x755 & ~x756 & ~x757 & ~x758 & ~x759 & ~x760 & ~x762 & ~x763 & ~x768 & ~x769 & ~x776 & ~x777 & ~x780 & ~x782;
assign c3280 =  x270 &  x271 &  x297 &  x298 &  x325 &  x351 &  x574 &  x575 &  x600 & ~x10 & ~x12 & ~x13 & ~x16 & ~x18 & ~x21 & ~x22 & ~x23 & ~x26 & ~x29 & ~x33 & ~x41 & ~x43 & ~x60 & ~x67 & ~x86 & ~x91 & ~x118 & ~x141 & ~x144 & ~x149 & ~x166 & ~x167 & ~x169 & ~x170 & ~x192 & ~x228 & ~x248 & ~x253 & ~x259 & ~x284 & ~x287 & ~x288 & ~x303 & ~x305 & ~x307 & ~x313 & ~x314 & ~x331 & ~x335 & ~x365 & ~x367 & ~x368 & ~x370 & ~x387 & ~x393 & ~x417 & ~x418 & ~x445 & ~x449 & ~x474 & ~x503 & ~x504 & ~x531 & ~x535 & ~x557 & ~x558 & ~x560 & ~x582 & ~x590 & ~x611 & ~x613 & ~x617 & ~x641 & ~x643 & ~x644 & ~x645 & ~x646 & ~x665 & ~x670 & ~x671 & ~x674 & ~x688 & ~x692 & ~x697 & ~x698 & ~x704 & ~x712 & ~x713 & ~x716 & ~x720 & ~x730 & ~x744 & ~x746 & ~x751 & ~x753 & ~x756 & ~x765 & ~x767 & ~x771 & ~x781 & ~x782;
assign c3282 =  x266 &  x294 &  x627 & ~x13 & ~x15 & ~x18 & ~x22 & ~x56 & ~x58 & ~x84 & ~x91 & ~x104 & ~x111 & ~x132 & ~x161 & ~x162 & ~x168 & ~x169 & ~x192 & ~x194 & ~x195 & ~x219 & ~x245 & ~x246 & ~x254 & ~x272 & ~x273 & ~x311 & ~x312 & ~x333 & ~x339 & ~x358 & ~x415 & ~x447 & ~x448 & ~x472 & ~x485 & ~x507 & ~x512 & ~x590 & ~x610 & ~x613 & ~x614 & ~x617 & ~x641 & ~x644 & ~x647 & ~x725 & ~x731 & ~x735 & ~x749 & ~x757 & ~x778 & ~x783;
assign c3284 =  x779;
assign c3286 =  x306;
assign c3288 =  x210 &  x243 &  x326 &  x352 &  x378 &  x379 & ~x1 & ~x2 & ~x7 & ~x10 & ~x11 & ~x17 & ~x19 & ~x32 & ~x37 & ~x41 & ~x69 & ~x70 & ~x77 & ~x80 & ~x84 & ~x88 & ~x95 & ~x98 & ~x103 & ~x104 & ~x108 & ~x110 & ~x113 & ~x135 & ~x141 & ~x165 & ~x166 & ~x194 & ~x195 & ~x196 & ~x198 & ~x225 & ~x248 & ~x276 & ~x280 & ~x281 & ~x306 & ~x310 & ~x311 & ~x339 & ~x364 & ~x387 & ~x388 & ~x392 & ~x393 & ~x394 & ~x421 & ~x423 & ~x445 & ~x446 & ~x472 & ~x477 & ~x488 & ~x490 & ~x518 & ~x528 & ~x529 & ~x532 & ~x556 & ~x558 & ~x584 & ~x611 & ~x617 & ~x642 & ~x667 & ~x671 & ~x673 & ~x692 & ~x694 & ~x713 & ~x720 & ~x726 & ~x733 & ~x740 & ~x756 & ~x758 & ~x766 & ~x767 & ~x769 & ~x776;
assign c3292 =  x241 &  x296 &  x350 &  x466 &  x494 &  x577 &  x603 & ~x5 & ~x7 & ~x18 & ~x22 & ~x28 & ~x37 & ~x48 & ~x51 & ~x52 & ~x55 & ~x60 & ~x61 & ~x83 & ~x106 & ~x107 & ~x110 & ~x114 & ~x136 & ~x141 & ~x143 & ~x163 & ~x194 & ~x220 & ~x224 & ~x246 & ~x247 & ~x250 & ~x286 & ~x306 & ~x310 & ~x338 & ~x360 & ~x367 & ~x386 & ~x392 & ~x396 & ~x420 & ~x421 & ~x423 & ~x445 & ~x450 & ~x477 & ~x500 & ~x528 & ~x533 & ~x557 & ~x563 & ~x584 & ~x587 & ~x613 & ~x639 & ~x641 & ~x643 & ~x670 & ~x674 & ~x694 & ~x706 & ~x719 & ~x720 & ~x722 & ~x723 & ~x726 & ~x732 & ~x751 & ~x752 & ~x765 & ~x769 & ~x770 & ~x781;
assign c3294 =  x295 &  x349 & ~x1 & ~x6 & ~x11 & ~x12 & ~x20 & ~x21 & ~x22 & ~x23 & ~x24 & ~x27 & ~x29 & ~x32 & ~x35 & ~x39 & ~x40 & ~x45 & ~x46 & ~x58 & ~x67 & ~x71 & ~x73 & ~x74 & ~x79 & ~x80 & ~x83 & ~x86 & ~x92 & ~x100 & ~x102 & ~x106 & ~x110 & ~x116 & ~x132 & ~x133 & ~x138 & ~x141 & ~x143 & ~x164 & ~x167 & ~x169 & ~x170 & ~x189 & ~x191 & ~x192 & ~x195 & ~x217 & ~x221 & ~x226 & ~x227 & ~x246 & ~x271 & ~x272 & ~x273 & ~x274 & ~x280 & ~x281 & ~x303 & ~x304 & ~x308 & ~x333 & ~x336 & ~x339 & ~x359 & ~x363 & ~x393 & ~x395 & ~x421 & ~x422 & ~x425 & ~x426 & ~x444 & ~x447 & ~x472 & ~x473 & ~x474 & ~x476 & ~x478 & ~x479 & ~x480 & ~x487 & ~x489 & ~x516 & ~x534 & ~x556 & ~x559 & ~x560 & ~x564 & ~x584 & ~x585 & ~x588 & ~x589 & ~x591 & ~x617 & ~x618 & ~x640 & ~x648 & ~x667 & ~x668 & ~x675 & ~x677 & ~x693 & ~x694 & ~x698 & ~x701 & ~x703 & ~x705 & ~x706 & ~x719 & ~x720 & ~x723 & ~x738 & ~x740 & ~x742 & ~x747 & ~x748 & ~x759 & ~x760 & ~x766 & ~x771 & ~x772 & ~x773 & ~x776 & ~x778 & ~x779 & ~x781 & ~x782 & ~x783;
assign c3296 =  x114;
assign c3298 = ~x0 & ~x2 & ~x3 & ~x6 & ~x7 & ~x9 & ~x11 & ~x15 & ~x16 & ~x17 & ~x19 & ~x21 & ~x22 & ~x24 & ~x31 & ~x32 & ~x33 & ~x44 & ~x50 & ~x52 & ~x53 & ~x57 & ~x61 & ~x70 & ~x71 & ~x74 & ~x77 & ~x79 & ~x80 & ~x82 & ~x84 & ~x85 & ~x89 & ~x92 & ~x104 & ~x105 & ~x107 & ~x108 & ~x109 & ~x111 & ~x112 & ~x114 & ~x115 & ~x133 & ~x134 & ~x136 & ~x138 & ~x139 & ~x140 & ~x143 & ~x164 & ~x169 & ~x190 & ~x191 & ~x195 & ~x198 & ~x218 & ~x221 & ~x222 & ~x226 & ~x246 & ~x247 & ~x250 & ~x253 & ~x254 & ~x259 & ~x260 & ~x261 & ~x262 & ~x263 & ~x275 & ~x276 & ~x278 & ~x279 & ~x280 & ~x281 & ~x282 & ~x286 & ~x287 & ~x288 & ~x304 & ~x305 & ~x307 & ~x311 & ~x313 & ~x314 & ~x332 & ~x333 & ~x334 & ~x338 & ~x340 & ~x360 & ~x362 & ~x363 & ~x367 & ~x369 & ~x388 & ~x389 & ~x392 & ~x393 & ~x394 & ~x395 & ~x417 & ~x420 & ~x422 & ~x425 & ~x428 & ~x444 & ~x447 & ~x451 & ~x452 & ~x453 & ~x454 & ~x456 & ~x457 & ~x458 & ~x473 & ~x474 & ~x477 & ~x478 & ~x482 & ~x486 & ~x488 & ~x489 & ~x502 & ~x504 & ~x518 & ~x529 & ~x530 & ~x531 & ~x532 & ~x556 & ~x558 & ~x559 & ~x560 & ~x585 & ~x586 & ~x588 & ~x614 & ~x615 & ~x616 & ~x617 & ~x618 & ~x639 & ~x640 & ~x642 & ~x643 & ~x644 & ~x645 & ~x648 & ~x666 & ~x667 & ~x668 & ~x669 & ~x672 & ~x676 & ~x694 & ~x696 & ~x700 & ~x704 & ~x709 & ~x711 & ~x716 & ~x717 & ~x718 & ~x719 & ~x720 & ~x723 & ~x726 & ~x727 & ~x730 & ~x732 & ~x735 & ~x736 & ~x737 & ~x738 & ~x740 & ~x741 & ~x742 & ~x744 & ~x746 & ~x747 & ~x752 & ~x754 & ~x755 & ~x757 & ~x759 & ~x760 & ~x762 & ~x763 & ~x764 & ~x769 & ~x770 & ~x771 & ~x773 & ~x775 & ~x777 & ~x779 & ~x780 & ~x781;
assign c31 = ~x17 & ~x31 & ~x37 & ~x40 & ~x57 & ~x59 & ~x76 & ~x79 & ~x81 & ~x83 & ~x87 & ~x95 & ~x122 & ~x123 & ~x125 & ~x148 & ~x150 & ~x151 & ~x152 & ~x153 & ~x179 & ~x194 & ~x198 & ~x207 & ~x225 & ~x228 & ~x233 & ~x235 & ~x262 & ~x289 & ~x307 & ~x335 & ~x337 & ~x341 & ~x397 & ~x416 & ~x417 & ~x478 & ~x501 & ~x558 & ~x643 & ~x660 & ~x686 & ~x699 & ~x700 & ~x713 & ~x716 & ~x726 & ~x763;
assign c33 = ~x0 & ~x1 & ~x6 & ~x7 & ~x9 & ~x15 & ~x17 & ~x21 & ~x23 & ~x27 & ~x30 & ~x39 & ~x41 & ~x42 & ~x47 & ~x51 & ~x58 & ~x63 & ~x65 & ~x66 & ~x76 & ~x79 & ~x85 & ~x87 & ~x88 & ~x89 & ~x91 & ~x92 & ~x94 & ~x95 & ~x97 & ~x100 & ~x101 & ~x104 & ~x105 & ~x107 & ~x110 & ~x112 & ~x114 & ~x117 & ~x119 & ~x122 & ~x127 & ~x128 & ~x129 & ~x137 & ~x141 & ~x142 & ~x146 & ~x149 & ~x150 & ~x151 & ~x170 & ~x194 & ~x196 & ~x222 & ~x253 & ~x274 & ~x279 & ~x306 & ~x309 & ~x332 & ~x336 & ~x337 & ~x363 & ~x364 & ~x365 & ~x390 & ~x391 & ~x392 & ~x394 & ~x395 & ~x416 & ~x422 & ~x444 & ~x450 & ~x472 & ~x474 & ~x477 & ~x478 & ~x499 & ~x500 & ~x505 & ~x506 & ~x513 & ~x514 & ~x515 & ~x516 & ~x529 & ~x539 & ~x541 & ~x542 & ~x543 & ~x555 & ~x561 & ~x562 & ~x569 & ~x572 & ~x580 & ~x581 & ~x582 & ~x591 & ~x618 & ~x620 & ~x637 & ~x644 & ~x646 & ~x648 & ~x665 & ~x666 & ~x676 & ~x677 & ~x680 & ~x682 & ~x683 & ~x693 & ~x695 & ~x698 & ~x699 & ~x709 & ~x711 & ~x722 & ~x723 & ~x726 & ~x727 & ~x728 & ~x729 & ~x736 & ~x739 & ~x750 & ~x754 & ~x757 & ~x759 & ~x761 & ~x763 & ~x768 & ~x770 & ~x771 & ~x776 & ~x777 & ~x778 & ~x782 & ~x783;
assign c35 =  x357 & ~x16 & ~x248 & ~x381 & ~x640;
assign c37 =  x572 &  x600 & ~x3 & ~x7 & ~x9 & ~x17 & ~x18 & ~x23 & ~x31 & ~x34 & ~x39 & ~x47 & ~x49 & ~x61 & ~x62 & ~x76 & ~x77 & ~x81 & ~x82 & ~x89 & ~x90 & ~x93 & ~x95 & ~x104 & ~x115 & ~x120 & ~x121 & ~x122 & ~x135 & ~x138 & ~x140 & ~x141 & ~x142 & ~x146 & ~x160 & ~x164 & ~x165 & ~x170 & ~x173 & ~x174 & ~x222 & ~x225 & ~x254 & ~x277 & ~x279 & ~x282 & ~x284 & ~x285 & ~x305 & ~x311 & ~x313 & ~x314 & ~x334 & ~x339 & ~x360 & ~x368 & ~x370 & ~x387 & ~x391 & ~x394 & ~x397 & ~x398 & ~x399 & ~x416 & ~x418 & ~x420 & ~x421 & ~x422 & ~x446 & ~x447 & ~x451 & ~x452 & ~x470 & ~x476 & ~x477 & ~x479 & ~x480 & ~x481 & ~x498 & ~x506 & ~x513 & ~x530 & ~x531 & ~x534 & ~x536 & ~x540 & ~x556 & ~x563 & ~x567 & ~x569 & ~x583 & ~x587 & ~x593 & ~x615 & ~x616 & ~x618 & ~x620 & ~x621 & ~x639 & ~x640 & ~x642 & ~x646 & ~x647 & ~x649 & ~x668 & ~x673 & ~x675 & ~x676 & ~x677 & ~x700 & ~x702 & ~x704 & ~x705 & ~x717 & ~x721 & ~x727 & ~x730 & ~x744 & ~x745 & ~x747 & ~x749 & ~x753 & ~x756 & ~x765 & ~x766 & ~x768 & ~x769 & ~x779;
assign c39 =  x432 &  x459 &  x486 &  x540 & ~x24 & ~x27 & ~x39 & ~x51 & ~x85 & ~x116 & ~x143 & ~x166 & ~x257 & ~x278 & ~x284 & ~x362 & ~x365 & ~x425 & ~x427 & ~x477 & ~x560 & ~x588 & ~x616 & ~x687 & ~x696 & ~x712 & ~x713 & ~x726 & ~x731 & ~x745 & ~x754 & ~x755 & ~x756 & ~x759 & ~x766 & ~x770 & ~x783;
assign c311 =  x319 &  x347 &  x403 & ~x2 & ~x14 & ~x19 & ~x21 & ~x32 & ~x35 & ~x36 & ~x60 & ~x62 & ~x92 & ~x99 & ~x124 & ~x147 & ~x166 & ~x169 & ~x172 & ~x174 & ~x176 & ~x197 & ~x198 & ~x202 & ~x204 & ~x222 & ~x250 & ~x251 & ~x257 & ~x277 & ~x284 & ~x285 & ~x286 & ~x307 & ~x309 & ~x311 & ~x335 & ~x341 & ~x364 & ~x421 & ~x448 & ~x478 & ~x507 & ~x531 & ~x534 & ~x535 & ~x559 & ~x586 & ~x611 & ~x612 & ~x617 & ~x695 & ~x704 & ~x721 & ~x725 & ~x727 & ~x730 & ~x731 & ~x732 & ~x739 & ~x740 & ~x748 & ~x751 & ~x756 & ~x770 & ~x775 & ~x781 & ~x782;
assign c313 =  x315 &  x370 &  x398 & ~x58 & ~x83 & ~x141 & ~x251 & ~x448 & ~x767;
assign c315 =  x431 &  x485 &  x540 & ~x15 & ~x425 & ~x524 & ~x617;
assign c317 = ~x6 & ~x9 & ~x11 & ~x15 & ~x18 & ~x27 & ~x30 & ~x34 & ~x37 & ~x47 & ~x52 & ~x53 & ~x60 & ~x61 & ~x66 & ~x77 & ~x78 & ~x82 & ~x83 & ~x85 & ~x87 & ~x92 & ~x106 & ~x107 & ~x110 & ~x112 & ~x115 & ~x116 & ~x137 & ~x138 & ~x141 & ~x142 & ~x144 & ~x163 & ~x165 & ~x167 & ~x168 & ~x169 & ~x170 & ~x172 & ~x173 & ~x193 & ~x197 & ~x200 & ~x217 & ~x242 & ~x252 & ~x265 & ~x267 & ~x277 & ~x312 & ~x336 & ~x337 & ~x340 & ~x360 & ~x367 & ~x390 & ~x391 & ~x417 & ~x421 & ~x422 & ~x446 & ~x450 & ~x451 & ~x452 & ~x474 & ~x475 & ~x476 & ~x477 & ~x478 & ~x479 & ~x502 & ~x504 & ~x530 & ~x531 & ~x535 & ~x557 & ~x558 & ~x563 & ~x586 & ~x587 & ~x589 & ~x591 & ~x612 & ~x613 & ~x617 & ~x620 & ~x640 & ~x641 & ~x642 & ~x645 & ~x648 & ~x666 & ~x673 & ~x675 & ~x677 & ~x678 & ~x680 & ~x692 & ~x698 & ~x703 & ~x704 & ~x706 & ~x707 & ~x711 & ~x722 & ~x727 & ~x730 & ~x734 & ~x735 & ~x739 & ~x742 & ~x743 & ~x744 & ~x747 & ~x752 & ~x755 & ~x756 & ~x758 & ~x760 & ~x765 & ~x766 & ~x767 & ~x768 & ~x770 & ~x775 & ~x776 & ~x777 & ~x778 & ~x781 & ~x782;
assign c319 =  x263 &  x291 &  x319 & ~x20 & ~x22 & ~x31 & ~x34 & ~x40 & ~x43 & ~x45 & ~x49 & ~x50 & ~x53 & ~x58 & ~x64 & ~x80 & ~x90 & ~x97 & ~x142 & ~x143 & ~x145 & ~x147 & ~x166 & ~x175 & ~x195 & ~x198 & ~x221 & ~x225 & ~x231 & ~x255 & ~x256 & ~x258 & ~x282 & ~x284 & ~x286 & ~x288 & ~x307 & ~x309 & ~x315 & ~x338 & ~x361 & ~x363 & ~x388 & ~x417 & ~x419 & ~x421 & ~x422 & ~x423 & ~x472 & ~x476 & ~x479 & ~x503 & ~x561 & ~x563 & ~x583 & ~x584 & ~x613 & ~x641 & ~x642 & ~x645 & ~x646 & ~x668 & ~x696 & ~x710 & ~x711 & ~x714 & ~x716 & ~x726 & ~x730 & ~x731 & ~x739 & ~x751 & ~x770 & ~x776 & ~x783;
assign c321 = ~x2 & ~x5 & ~x10 & ~x16 & ~x18 & ~x22 & ~x27 & ~x29 & ~x31 & ~x40 & ~x41 & ~x74 & ~x79 & ~x82 & ~x87 & ~x108 & ~x112 & ~x113 & ~x115 & ~x116 & ~x165 & ~x168 & ~x196 & ~x198 & ~x225 & ~x227 & ~x228 & ~x252 & ~x253 & ~x295 & ~x322 & ~x324 & ~x333 & ~x334 & ~x349 & ~x364 & ~x366 & ~x378 & ~x390 & ~x394 & ~x417 & ~x418 & ~x419 & ~x422 & ~x450 & ~x476 & ~x502 & ~x504 & ~x532 & ~x560 & ~x587 & ~x613 & ~x642 & ~x671 & ~x672 & ~x674 & ~x676 & ~x678 & ~x687 & ~x698 & ~x703 & ~x710 & ~x719 & ~x725 & ~x729 & ~x745 & ~x747 & ~x752 & ~x765 & ~x766 & ~x770 & ~x776 & ~x781;
assign c323 =  x517 &  x572 & ~x4 & ~x6 & ~x10 & ~x12 & ~x13 & ~x20 & ~x21 & ~x22 & ~x23 & ~x26 & ~x28 & ~x32 & ~x34 & ~x36 & ~x37 & ~x41 & ~x46 & ~x52 & ~x59 & ~x61 & ~x62 & ~x66 & ~x73 & ~x76 & ~x83 & ~x84 & ~x99 & ~x100 & ~x104 & ~x108 & ~x109 & ~x110 & ~x111 & ~x115 & ~x118 & ~x133 & ~x142 & ~x163 & ~x193 & ~x197 & ~x198 & ~x220 & ~x221 & ~x223 & ~x224 & ~x247 & ~x251 & ~x254 & ~x276 & ~x282 & ~x283 & ~x306 & ~x308 & ~x312 & ~x313 & ~x335 & ~x338 & ~x341 & ~x360 & ~x361 & ~x363 & ~x364 & ~x387 & ~x388 & ~x391 & ~x395 & ~x400 & ~x417 & ~x423 & ~x426 & ~x428 & ~x452 & ~x453 & ~x456 & ~x469 & ~x470 & ~x476 & ~x480 & ~x503 & ~x508 & ~x531 & ~x533 & ~x538 & ~x539 & ~x541 & ~x565 & ~x567 & ~x587 & ~x588 & ~x589 & ~x590 & ~x591 & ~x594 & ~x595 & ~x614 & ~x616 & ~x622 & ~x623 & ~x640 & ~x643 & ~x645 & ~x650 & ~x667 & ~x672 & ~x674 & ~x676 & ~x696 & ~x699 & ~x700 & ~x703 & ~x705 & ~x706 & ~x721 & ~x724 & ~x726 & ~x729 & ~x730 & ~x731 & ~x741 & ~x744 & ~x749 & ~x753 & ~x754 & ~x761 & ~x764 & ~x767 & ~x771 & ~x773 & ~x782;
assign c325 =  x314 &  x342 & ~x2 & ~x3 & ~x19 & ~x76 & ~x82 & ~x90 & ~x123 & ~x306 & ~x307 & ~x336 & ~x587 & ~x652 & ~x674 & ~x682 & ~x706 & ~x709 & ~x738 & ~x751 & ~x759;
assign c327 =  x320 &  x348 &  x406 & ~x3 & ~x8 & ~x11 & ~x13 & ~x16 & ~x18 & ~x21 & ~x24 & ~x30 & ~x32 & ~x34 & ~x36 & ~x39 & ~x41 & ~x46 & ~x50 & ~x51 & ~x55 & ~x58 & ~x64 & ~x70 & ~x75 & ~x76 & ~x78 & ~x83 & ~x88 & ~x94 & ~x98 & ~x102 & ~x116 & ~x119 & ~x121 & ~x123 & ~x139 & ~x140 & ~x144 & ~x145 & ~x166 & ~x167 & ~x170 & ~x171 & ~x172 & ~x175 & ~x194 & ~x195 & ~x196 & ~x199 & ~x200 & ~x222 & ~x226 & ~x229 & ~x250 & ~x256 & ~x259 & ~x278 & ~x281 & ~x282 & ~x286 & ~x307 & ~x308 & ~x313 & ~x336 & ~x340 & ~x363 & ~x364 & ~x367 & ~x368 & ~x369 & ~x372 & ~x387 & ~x398 & ~x417 & ~x419 & ~x420 & ~x422 & ~x426 & ~x449 & ~x470 & ~x472 & ~x473 & ~x476 & ~x480 & ~x501 & ~x502 & ~x507 & ~x554 & ~x555 & ~x557 & ~x559 & ~x561 & ~x582 & ~x583 & ~x585 & ~x589 & ~x590 & ~x610 & ~x611 & ~x612 & ~x614 & ~x615 & ~x616 & ~x619 & ~x620 & ~x640 & ~x645 & ~x670 & ~x671 & ~x672 & ~x674 & ~x692 & ~x695 & ~x712 & ~x713 & ~x714 & ~x715 & ~x718 & ~x719 & ~x721 & ~x725 & ~x729 & ~x730 & ~x732 & ~x733 & ~x738 & ~x749 & ~x751 & ~x752 & ~x754 & ~x756 & ~x763 & ~x764 & ~x769 & ~x770 & ~x773;
assign c329 =  x325 &  x353 &  x464 &  x492 & ~x10 & ~x11 & ~x17 & ~x27 & ~x47 & ~x59 & ~x70 & ~x77 & ~x80 & ~x91 & ~x92 & ~x101 & ~x112 & ~x114 & ~x118 & ~x138 & ~x140 & ~x167 & ~x223 & ~x225 & ~x274 & ~x350 & ~x594 & ~x617 & ~x678 & ~x692 & ~x696 & ~x697 & ~x698 & ~x699 & ~x710 & ~x724 & ~x726 & ~x732 & ~x744 & ~x758 & ~x773;
assign c331 =  x338;
assign c333 =  x380 &  x408 &  x436 &  x464 & ~x1 & ~x4 & ~x8 & ~x12 & ~x16 & ~x20 & ~x21 & ~x33 & ~x35 & ~x41 & ~x45 & ~x52 & ~x55 & ~x59 & ~x61 & ~x62 & ~x64 & ~x66 & ~x69 & ~x72 & ~x75 & ~x76 & ~x82 & ~x88 & ~x89 & ~x94 & ~x98 & ~x104 & ~x106 & ~x110 & ~x128 & ~x140 & ~x159 & ~x163 & ~x194 & ~x195 & ~x222 & ~x227 & ~x248 & ~x280 & ~x337 & ~x359 & ~x362 & ~x368 & ~x389 & ~x397 & ~x416 & ~x417 & ~x421 & ~x423 & ~x424 & ~x451 & ~x453 & ~x474 & ~x475 & ~x476 & ~x478 & ~x480 & ~x496 & ~x499 & ~x501 & ~x506 & ~x509 & ~x512 & ~x513 & ~x527 & ~x531 & ~x533 & ~x551 & ~x561 & ~x564 & ~x585 & ~x591 & ~x611 & ~x615 & ~x616 & ~x617 & ~x619 & ~x620 & ~x621 & ~x622 & ~x623 & ~x640 & ~x644 & ~x646 & ~x650 & ~x668 & ~x670 & ~x678 & ~x698 & ~x704 & ~x707 & ~x708 & ~x722 & ~x723 & ~x726 & ~x756 & ~x758 & ~x762 & ~x765 & ~x774 & ~x777 & ~x778;
assign c335 =  x372 &  x427 & ~x1 & ~x9 & ~x35 & ~x709;
assign c337 = ~x0 & ~x50 & ~x51 & ~x54 & ~x55 & ~x66 & ~x79 & ~x90 & ~x96 & ~x98 & ~x137 & ~x141 & ~x196 & ~x278 & ~x350 & ~x352 & ~x379 & ~x406 & ~x420 & ~x435 & ~x500 & ~x528 & ~x587 & ~x588 & ~x590 & ~x704 & ~x706 & ~x723 & ~x728 & ~x756 & ~x757 & ~x759 & ~x761 & ~x763 & ~x779;
assign c339 =  x545 & ~x82 & ~x166 & ~x325 & ~x381 & ~x421 & ~x681 & ~x688;
assign c341 =  x432 &  x514 &  x542 &  x570 & ~x6 & ~x37 & ~x57 & ~x86 & ~x139 & ~x225 & ~x230 & ~x311 & ~x389 & ~x424 & ~x452 & ~x480 & ~x509 & ~x586 & ~x638 & ~x643 & ~x644 & ~x722 & ~x724 & ~x725 & ~x761;
assign c343 = ~x6 & ~x11 & ~x14 & ~x15 & ~x19 & ~x33 & ~x36 & ~x44 & ~x57 & ~x64 & ~x73 & ~x76 & ~x80 & ~x87 & ~x88 & ~x102 & ~x105 & ~x116 & ~x136 & ~x138 & ~x165 & ~x170 & ~x194 & ~x195 & ~x225 & ~x248 & ~x323 & ~x363 & ~x379 & ~x404 & ~x407 & ~x434 & ~x444 & ~x445 & ~x448 & ~x449 & ~x478 & ~x500 & ~x502 & ~x503 & ~x535 & ~x586 & ~x644 & ~x674 & ~x725 & ~x729 & ~x732 & ~x734 & ~x751 & ~x752 & ~x757 & ~x759 & ~x760;
assign c345 =  x329 & ~x14 & ~x16 & ~x17 & ~x28 & ~x70 & ~x91 & ~x92 & ~x114 & ~x169 & ~x171 & ~x198 & ~x338 & ~x380 & ~x391 & ~x418 & ~x503 & ~x616 & ~x668;
assign c347 =  x518 & ~x0 & ~x16 & ~x19 & ~x21 & ~x27 & ~x32 & ~x33 & ~x60 & ~x80 & ~x83 & ~x134 & ~x137 & ~x194 & ~x255 & ~x283 & ~x306 & ~x334 & ~x354 & ~x360 & ~x422 & ~x477 & ~x530 & ~x559 & ~x584 & ~x606 & ~x607 & ~x613 & ~x625 & ~x636 & ~x646 & ~x651 & ~x654 & ~x681 & ~x682 & ~x690 & ~x711 & ~x717 & ~x719 & ~x750 & ~x761 & ~x763;
assign c349 =  x409 &  x519 &  x546 & ~x44 & ~x86 & ~x89 & ~x107 & ~x164 & ~x165 & ~x169 & ~x194 & ~x199 & ~x275 & ~x323 & ~x450 & ~x533 & ~x560 & ~x591 & ~x612 & ~x617 & ~x662 & ~x679 & ~x734 & ~x754;
assign c351 =  x489 &  x544 & ~x18 & ~x39 & ~x49 & ~x54 & ~x73 & ~x78 & ~x82 & ~x87 & ~x162 & ~x193 & ~x221 & ~x222 & ~x251 & ~x254 & ~x279 & ~x293 & ~x303 & ~x305 & ~x338 & ~x348 & ~x361 & ~x365 & ~x420 & ~x506 & ~x679 & ~x681 & ~x686 & ~x701 & ~x714 & ~x718 & ~x719 & ~x724 & ~x743 & ~x746 & ~x773;
assign c353 =  x370 &  x398;
assign c355 =  x348 &  x376 &  x377 & ~x4 & ~x11 & ~x14 & ~x15 & ~x18 & ~x21 & ~x25 & ~x27 & ~x28 & ~x29 & ~x32 & ~x36 & ~x41 & ~x50 & ~x53 & ~x54 & ~x55 & ~x56 & ~x61 & ~x64 & ~x88 & ~x89 & ~x95 & ~x118 & ~x140 & ~x147 & ~x167 & ~x172 & ~x197 & ~x201 & ~x227 & ~x258 & ~x277 & ~x281 & ~x286 & ~x296 & ~x297 & ~x308 & ~x310 & ~x337 & ~x386 & ~x388 & ~x393 & ~x423 & ~x447 & ~x474 & ~x479 & ~x500 & ~x531 & ~x559 & ~x589 & ~x612 & ~x615 & ~x617 & ~x619 & ~x643 & ~x648 & ~x668 & ~x672 & ~x673 & ~x674 & ~x689 & ~x697 & ~x699 & ~x701 & ~x704 & ~x705 & ~x708 & ~x715 & ~x717 & ~x727 & ~x731 & ~x738 & ~x746 & ~x748 & ~x757 & ~x768 & ~x770 & ~x777 & ~x781;
assign c357 =  x771;
assign c359 =  x261 &  x289 &  x344 &  x632 & ~x517;
assign c361 =  x276;
assign c363 = ~x3 & ~x7 & ~x9 & ~x19 & ~x20 & ~x26 & ~x28 & ~x29 & ~x36 & ~x38 & ~x46 & ~x51 & ~x53 & ~x58 & ~x82 & ~x83 & ~x86 & ~x113 & ~x116 & ~x117 & ~x132 & ~x140 & ~x168 & ~x171 & ~x193 & ~x194 & ~x200 & ~x222 & ~x226 & ~x228 & ~x255 & ~x256 & ~x277 & ~x281 & ~x285 & ~x304 & ~x306 & ~x318 & ~x332 & ~x337 & ~x345 & ~x346 & ~x360 & ~x367 & ~x370 & ~x387 & ~x388 & ~x389 & ~x392 & ~x396 & ~x399 & ~x412 & ~x418 & ~x422 & ~x425 & ~x437 & ~x438 & ~x439 & ~x442 & ~x446 & ~x465 & ~x476 & ~x481 & ~x503 & ~x504 & ~x505 & ~x506 & ~x508 & ~x561 & ~x563 & ~x591 & ~x614 & ~x642 & ~x662 & ~x663 & ~x664 & ~x674 & ~x676 & ~x683 & ~x686 & ~x687 & ~x691 & ~x693 & ~x697 & ~x702 & ~x704 & ~x708 & ~x710 & ~x712 & ~x713 & ~x715 & ~x727 & ~x730 & ~x736 & ~x738 & ~x742 & ~x744 & ~x749 & ~x752 & ~x753 & ~x755 & ~x765 & ~x766 & ~x769 & ~x772 & ~x776 & ~x777 & ~x779 & ~x780 & ~x781;
assign c365 =  x386 & ~x252 & ~x279;
assign c367 =  x261 &  x317 & ~x4 & ~x38 & ~x62 & ~x72 & ~x89 & ~x109 & ~x114 & ~x144 & ~x171 & ~x308 & ~x391 & ~x419 & ~x434 & ~x474 & ~x475 & ~x516 & ~x528 & ~x529 & ~x530 & ~x557 & ~x558 & ~x586 & ~x619 & ~x648 & ~x649 & ~x651 & ~x665 & ~x675 & ~x729 & ~x751 & ~x755;
assign c369 =  x399 & ~x11 & ~x15 & ~x36 & ~x43 & ~x56 & ~x61 & ~x72 & ~x109 & ~x115 & ~x137 & ~x166 & ~x193 & ~x223 & ~x304 & ~x307 & ~x332 & ~x347 & ~x348 & ~x361 & ~x394 & ~x448 & ~x501 & ~x559 & ~x591 & ~x675 & ~x727 & ~x750 & ~x756 & ~x775 & ~x778;
assign c371 =  x462 &  x463 &  x490 & ~x0 & ~x1 & ~x3 & ~x5 & ~x6 & ~x9 & ~x11 & ~x12 & ~x13 & ~x16 & ~x20 & ~x25 & ~x27 & ~x28 & ~x29 & ~x30 & ~x34 & ~x35 & ~x36 & ~x37 & ~x38 & ~x40 & ~x41 & ~x43 & ~x46 & ~x48 & ~x49 & ~x51 & ~x54 & ~x55 & ~x56 & ~x58 & ~x59 & ~x60 & ~x62 & ~x63 & ~x67 & ~x68 & ~x74 & ~x79 & ~x82 & ~x85 & ~x86 & ~x88 & ~x90 & ~x107 & ~x112 & ~x113 & ~x114 & ~x117 & ~x137 & ~x138 & ~x140 & ~x141 & ~x142 & ~x144 & ~x163 & ~x166 & ~x167 & ~x191 & ~x196 & ~x197 & ~x199 & ~x219 & ~x221 & ~x223 & ~x224 & ~x225 & ~x248 & ~x249 & ~x250 & ~x252 & ~x253 & ~x254 & ~x255 & ~x256 & ~x275 & ~x280 & ~x281 & ~x283 & ~x306 & ~x311 & ~x332 & ~x333 & ~x334 & ~x335 & ~x362 & ~x366 & ~x367 & ~x389 & ~x390 & ~x391 & ~x392 & ~x393 & ~x395 & ~x417 & ~x418 & ~x420 & ~x422 & ~x447 & ~x450 & ~x475 & ~x476 & ~x478 & ~x503 & ~x506 & ~x529 & ~x530 & ~x531 & ~x533 & ~x558 & ~x562 & ~x587 & ~x588 & ~x590 & ~x614 & ~x616 & ~x618 & ~x629 & ~x642 & ~x643 & ~x645 & ~x646 & ~x647 & ~x649 & ~x657 & ~x658 & ~x666 & ~x667 & ~x669 & ~x672 & ~x673 & ~x683 & ~x684 & ~x685 & ~x686 & ~x690 & ~x691 & ~x692 & ~x695 & ~x697 & ~x698 & ~x700 & ~x703 & ~x704 & ~x712 & ~x713 & ~x714 & ~x715 & ~x716 & ~x717 & ~x718 & ~x719 & ~x720 & ~x721 & ~x722 & ~x723 & ~x724 & ~x725 & ~x726 & ~x727 & ~x733 & ~x738 & ~x739 & ~x741 & ~x744 & ~x746 & ~x747 & ~x748 & ~x749 & ~x750 & ~x752 & ~x754 & ~x755 & ~x758 & ~x759 & ~x763 & ~x765 & ~x766 & ~x768 & ~x769 & ~x773 & ~x774 & ~x776 & ~x781 & ~x782;
assign c373 =  x320 & ~x98 & ~x203 & ~x282 & ~x383 & ~x410 & ~x438 & ~x439 & ~x452 & ~x507 & ~x674 & ~x705 & ~x747;
assign c375 =  x245 & ~x5 & ~x77 & ~x310 & ~x325 & ~x354 & ~x355 & ~x762;
assign c377 =  x326 &  x354 &  x410 &  x438 & ~x0 & ~x20 & ~x29 & ~x30 & ~x33 & ~x42 & ~x44 & ~x91 & ~x95 & ~x109 & ~x139 & ~x151 & ~x154 & ~x169 & ~x189 & ~x196 & ~x252 & ~x361 & ~x364 & ~x507 & ~x508 & ~x515 & ~x533 & ~x542 & ~x570 & ~x595 & ~x596 & ~x616 & ~x621 & ~x623 & ~x650 & ~x672 & ~x736 & ~x753;
assign c379 = ~x8 & ~x69 & ~x87 & ~x168 & ~x224 & ~x311 & ~x319 & ~x344 & ~x376 & ~x453 & ~x460 & ~x501 & ~x543 & ~x565 & ~x568 & ~x569 & ~x592 & ~x620 & ~x677 & ~x704 & ~x723 & ~x731;
assign c381 =  x290 &  x346 &  x375 & ~x18 & ~x61 & ~x131 & ~x145 & ~x193 & ~x362 & ~x387 & ~x389 & ~x413 & ~x428 & ~x442 & ~x449 & ~x453 & ~x470 & ~x501 & ~x621 & ~x649 & ~x678 & ~x725 & ~x748 & ~x762;
assign c383 =  x541;
assign c385 =  x460 &  x515 & ~x4 & ~x9 & ~x18 & ~x27 & ~x28 & ~x31 & ~x39 & ~x45 & ~x56 & ~x57 & ~x64 & ~x73 & ~x77 & ~x84 & ~x85 & ~x100 & ~x104 & ~x108 & ~x113 & ~x117 & ~x132 & ~x139 & ~x140 & ~x143 & ~x145 & ~x194 & ~x195 & ~x199 & ~x221 & ~x256 & ~x281 & ~x305 & ~x343 & ~x369 & ~x389 & ~x393 & ~x394 & ~x401 & ~x413 & ~x430 & ~x451 & ~x453 & ~x455 & ~x457 & ~x478 & ~x508 & ~x535 & ~x536 & ~x586 & ~x591 & ~x615 & ~x644 & ~x646 & ~x668 & ~x670 & ~x694 & ~x695 & ~x696 & ~x697 & ~x703 & ~x713 & ~x715 & ~x719 & ~x720 & ~x724 & ~x730 & ~x739 & ~x744 & ~x751 & ~x752 & ~x763 & ~x775 & ~x780;
assign c387 =  x431 &  x486 & ~x4 & ~x5 & ~x6 & ~x10 & ~x11 & ~x13 & ~x16 & ~x46 & ~x47 & ~x50 & ~x51 & ~x53 & ~x78 & ~x87 & ~x106 & ~x108 & ~x110 & ~x141 & ~x144 & ~x145 & ~x165 & ~x168 & ~x173 & ~x192 & ~x194 & ~x201 & ~x223 & ~x225 & ~x227 & ~x253 & ~x255 & ~x281 & ~x282 & ~x286 & ~x307 & ~x311 & ~x336 & ~x338 & ~x343 & ~x363 & ~x369 & ~x370 & ~x390 & ~x397 & ~x418 & ~x422 & ~x425 & ~x446 & ~x448 & ~x449 & ~x451 & ~x477 & ~x480 & ~x507 & ~x533 & ~x589 & ~x617 & ~x645 & ~x651 & ~x667 & ~x669 & ~x680 & ~x688 & ~x689 & ~x693 & ~x694 & ~x698 & ~x700 & ~x705 & ~x708 & ~x709 & ~x711 & ~x713 & ~x714 & ~x716 & ~x717 & ~x726 & ~x728 & ~x729 & ~x730 & ~x731 & ~x735 & ~x736 & ~x749 & ~x756 & ~x761 & ~x765 & ~x768 & ~x770 & ~x779 & ~x782 & ~x783;
assign c389 =  x232 &  x288 & ~x4 & ~x10 & ~x13 & ~x28 & ~x30 & ~x39 & ~x41 & ~x51 & ~x58 & ~x61 & ~x72 & ~x73 & ~x84 & ~x87 & ~x88 & ~x89 & ~x96 & ~x141 & ~x142 & ~x144 & ~x169 & ~x194 & ~x195 & ~x278 & ~x306 & ~x366 & ~x391 & ~x395 & ~x423 & ~x447 & ~x475 & ~x478 & ~x480 & ~x506 & ~x530 & ~x533 & ~x534 & ~x535 & ~x551 & ~x585 & ~x592 & ~x639 & ~x644 & ~x673 & ~x674 & ~x695 & ~x700 & ~x701 & ~x703 & ~x723 & ~x732 & ~x750 & ~x754 & ~x755 & ~x757 & ~x760 & ~x762 & ~x763 & ~x783;
assign c391 =  x488 &  x543 & ~x15 & ~x56 & ~x101 & ~x106 & ~x112 & ~x164 & ~x224 & ~x251 & ~x277 & ~x283 & ~x369 & ~x389 & ~x392 & ~x401 & ~x412 & ~x456 & ~x505 & ~x512 & ~x538 & ~x539 & ~x557 & ~x613 & ~x641 & ~x643 & ~x703 & ~x752 & ~x760 & ~x776;
assign c393 =  x209 &  x263 &  x291 &  x319 &  x347 & ~x4 & ~x5 & ~x6 & ~x7 & ~x12 & ~x18 & ~x20 & ~x26 & ~x35 & ~x40 & ~x41 & ~x52 & ~x55 & ~x58 & ~x61 & ~x64 & ~x65 & ~x73 & ~x76 & ~x79 & ~x92 & ~x93 & ~x94 & ~x113 & ~x118 & ~x120 & ~x122 & ~x140 & ~x142 & ~x147 & ~x148 & ~x149 & ~x165 & ~x170 & ~x174 & ~x175 & ~x177 & ~x196 & ~x202 & ~x204 & ~x229 & ~x256 & ~x259 & ~x281 & ~x287 & ~x310 & ~x332 & ~x341 & ~x361 & ~x371 & ~x415 & ~x419 & ~x424 & ~x451 & ~x479 & ~x500 & ~x504 & ~x529 & ~x531 & ~x533 & ~x556 & ~x561 & ~x562 & ~x581 & ~x584 & ~x616 & ~x638 & ~x696 & ~x699 & ~x701 & ~x703 & ~x707 & ~x721 & ~x723 & ~x725 & ~x727 & ~x728 & ~x731 & ~x739 & ~x744 & ~x758 & ~x759 & ~x763 & ~x765 & ~x771 & ~x774 & ~x778 & ~x780;
assign c395 =  x460 &  x570 & ~x0 & ~x1 & ~x18 & ~x19 & ~x20 & ~x24 & ~x30 & ~x31 & ~x33 & ~x34 & ~x36 & ~x39 & ~x40 & ~x43 & ~x44 & ~x54 & ~x57 & ~x58 & ~x61 & ~x62 & ~x72 & ~x79 & ~x84 & ~x85 & ~x88 & ~x94 & ~x109 & ~x116 & ~x117 & ~x139 & ~x164 & ~x171 & ~x173 & ~x194 & ~x197 & ~x200 & ~x225 & ~x227 & ~x228 & ~x333 & ~x334 & ~x335 & ~x360 & ~x368 & ~x419 & ~x424 & ~x440 & ~x443 & ~x445 & ~x450 & ~x452 & ~x506 & ~x531 & ~x534 & ~x559 & ~x587 & ~x616 & ~x645 & ~x674 & ~x704 & ~x721 & ~x723 & ~x728 & ~x733 & ~x739 & ~x751 & ~x756 & ~x758 & ~x759 & ~x763 & ~x769 & ~x773 & ~x775;
assign c397 =  x316 &  x375 & ~x91 & ~x99 & ~x109 & ~x172 & ~x173 & ~x292 & ~x451 & ~x587 & ~x589 & ~x641 & ~x701 & ~x737 & ~x773;
assign c399 =  x320 & ~x1 & ~x2 & ~x7 & ~x9 & ~x10 & ~x14 & ~x20 & ~x22 & ~x23 & ~x25 & ~x28 & ~x30 & ~x35 & ~x42 & ~x43 & ~x45 & ~x46 & ~x50 & ~x53 & ~x55 & ~x56 & ~x57 & ~x58 & ~x63 & ~x64 & ~x69 & ~x74 & ~x77 & ~x80 & ~x84 & ~x86 & ~x91 & ~x95 & ~x99 & ~x108 & ~x110 & ~x111 & ~x115 & ~x118 & ~x119 & ~x121 & ~x139 & ~x143 & ~x145 & ~x164 & ~x165 & ~x168 & ~x169 & ~x171 & ~x172 & ~x173 & ~x174 & ~x194 & ~x195 & ~x196 & ~x197 & ~x220 & ~x223 & ~x227 & ~x228 & ~x230 & ~x248 & ~x249 & ~x250 & ~x251 & ~x252 & ~x259 & ~x267 & ~x284 & ~x305 & ~x306 & ~x308 & ~x309 & ~x330 & ~x336 & ~x337 & ~x338 & ~x341 & ~x357 & ~x360 & ~x366 & ~x367 & ~x372 & ~x388 & ~x391 & ~x393 & ~x394 & ~x396 & ~x397 & ~x399 & ~x419 & ~x421 & ~x423 & ~x427 & ~x446 & ~x447 & ~x451 & ~x452 & ~x454 & ~x455 & ~x473 & ~x475 & ~x477 & ~x479 & ~x502 & ~x503 & ~x504 & ~x507 & ~x528 & ~x532 & ~x533 & ~x559 & ~x564 & ~x565 & ~x586 & ~x587 & ~x588 & ~x612 & ~x616 & ~x617 & ~x620 & ~x637 & ~x640 & ~x641 & ~x644 & ~x646 & ~x649 & ~x665 & ~x670 & ~x672 & ~x677 & ~x678 & ~x679 & ~x692 & ~x693 & ~x694 & ~x695 & ~x697 & ~x700 & ~x701 & ~x702 & ~x704 & ~x709 & ~x714 & ~x715 & ~x717 & ~x724 & ~x726 & ~x728 & ~x732 & ~x733 & ~x735 & ~x736 & ~x740 & ~x744 & ~x745 & ~x746 & ~x753 & ~x754 & ~x756 & ~x759 & ~x760 & ~x761 & ~x769 & ~x770 & ~x774 & ~x775;
assign c3101 = ~x13 & ~x21 & ~x26 & ~x32 & ~x38 & ~x47 & ~x55 & ~x60 & ~x73 & ~x91 & ~x98 & ~x101 & ~x116 & ~x123 & ~x124 & ~x127 & ~x150 & ~x163 & ~x172 & ~x177 & ~x336 & ~x361 & ~x365 & ~x431 & ~x446 & ~x449 & ~x457 & ~x459 & ~x477 & ~x531 & ~x534 & ~x551 & ~x554 & ~x564 & ~x567 & ~x580 & ~x586 & ~x606 & ~x615 & ~x622 & ~x637 & ~x640 & ~x664 & ~x665 & ~x668 & ~x679 & ~x697 & ~x705;
assign c3103 = ~x1 & ~x2 & ~x5 & ~x12 & ~x14 & ~x23 & ~x34 & ~x39 & ~x46 & ~x47 & ~x52 & ~x57 & ~x62 & ~x64 & ~x68 & ~x75 & ~x81 & ~x82 & ~x86 & ~x89 & ~x90 & ~x92 & ~x94 & ~x95 & ~x97 & ~x113 & ~x114 & ~x121 & ~x122 & ~x123 & ~x138 & ~x142 & ~x143 & ~x147 & ~x148 & ~x149 & ~x176 & ~x177 & ~x198 & ~x204 & ~x205 & ~x251 & ~x260 & ~x269 & ~x278 & ~x284 & ~x286 & ~x287 & ~x300 & ~x308 & ~x314 & ~x315 & ~x332 & ~x337 & ~x338 & ~x343 & ~x363 & ~x365 & ~x366 & ~x394 & ~x397 & ~x398 & ~x419 & ~x424 & ~x445 & ~x447 & ~x449 & ~x452 & ~x471 & ~x479 & ~x498 & ~x505 & ~x507 & ~x529 & ~x530 & ~x534 & ~x557 & ~x559 & ~x561 & ~x582 & ~x584 & ~x587 & ~x589 & ~x592 & ~x616 & ~x617 & ~x636 & ~x637 & ~x638 & ~x645 & ~x670 & ~x672 & ~x688 & ~x695 & ~x701 & ~x707 & ~x710 & ~x717 & ~x719 & ~x720 & ~x724 & ~x725 & ~x727 & ~x728 & ~x730 & ~x732 & ~x733 & ~x734 & ~x741 & ~x747 & ~x748 & ~x749 & ~x752 & ~x754 & ~x757 & ~x760 & ~x766 & ~x767 & ~x769 & ~x772 & ~x778;
assign c3105 =  x514 &  x541 & ~x5 & ~x6 & ~x8 & ~x11 & ~x17 & ~x21 & ~x25 & ~x32 & ~x34 & ~x40 & ~x46 & ~x48 & ~x51 & ~x53 & ~x54 & ~x56 & ~x57 & ~x58 & ~x60 & ~x61 & ~x67 & ~x75 & ~x76 & ~x81 & ~x83 & ~x88 & ~x94 & ~x98 & ~x102 & ~x108 & ~x134 & ~x137 & ~x138 & ~x141 & ~x162 & ~x165 & ~x167 & ~x168 & ~x195 & ~x200 & ~x221 & ~x226 & ~x227 & ~x228 & ~x256 & ~x279 & ~x283 & ~x307 & ~x309 & ~x338 & ~x339 & ~x364 & ~x368 & ~x369 & ~x371 & ~x394 & ~x395 & ~x396 & ~x398 & ~x401 & ~x422 & ~x425 & ~x446 & ~x451 & ~x453 & ~x455 & ~x475 & ~x480 & ~x482 & ~x504 & ~x509 & ~x510 & ~x533 & ~x562 & ~x590 & ~x642 & ~x644 & ~x647 & ~x667 & ~x673 & ~x676 & ~x692 & ~x700 & ~x701 & ~x702 & ~x714 & ~x716 & ~x720 & ~x723 & ~x732 & ~x738 & ~x742 & ~x744 & ~x752 & ~x753 & ~x765 & ~x768 & ~x772 & ~x776 & ~x778 & ~x781;
assign c3107 =  x484 & ~x6 & ~x14 & ~x26 & ~x31 & ~x33 & ~x47 & ~x56 & ~x82 & ~x143 & ~x163 & ~x190 & ~x195 & ~x197 & ~x198 & ~x219 & ~x222 & ~x282 & ~x306 & ~x307 & ~x339 & ~x419 & ~x452 & ~x477 & ~x478 & ~x507 & ~x533 & ~x561 & ~x589 & ~x616 & ~x631 & ~x642 & ~x658 & ~x660 & ~x668 & ~x669 & ~x678 & ~x687 & ~x690 & ~x697 & ~x700 & ~x709 & ~x712 & ~x714 & ~x715 & ~x729 & ~x731 & ~x733 & ~x738 & ~x743 & ~x745 & ~x749 & ~x760 & ~x762 & ~x764 & ~x766;
assign c3109 = ~x7 & ~x9 & ~x11 & ~x12 & ~x13 & ~x15 & ~x17 & ~x22 & ~x31 & ~x36 & ~x43 & ~x44 & ~x47 & ~x48 & ~x55 & ~x59 & ~x78 & ~x83 & ~x104 & ~x105 & ~x110 & ~x114 & ~x133 & ~x136 & ~x138 & ~x141 & ~x143 & ~x144 & ~x161 & ~x166 & ~x171 & ~x173 & ~x174 & ~x189 & ~x190 & ~x191 & ~x193 & ~x194 & ~x195 & ~x197 & ~x200 & ~x201 & ~x202 & ~x217 & ~x218 & ~x221 & ~x224 & ~x229 & ~x230 & ~x255 & ~x257 & ~x273 & ~x278 & ~x280 & ~x281 & ~x285 & ~x308 & ~x312 & ~x313 & ~x333 & ~x342 & ~x359 & ~x364 & ~x365 & ~x368 & ~x391 & ~x395 & ~x396 & ~x420 & ~x421 & ~x423 & ~x424 & ~x453 & ~x474 & ~x477 & ~x480 & ~x504 & ~x508 & ~x533 & ~x536 & ~x559 & ~x561 & ~x592 & ~x593 & ~x616 & ~x628 & ~x643 & ~x645 & ~x647 & ~x649 & ~x657 & ~x671 & ~x674 & ~x676 & ~x680 & ~x684 & ~x685 & ~x686 & ~x692 & ~x699 & ~x703 & ~x711 & ~x712 & ~x714 & ~x715 & ~x720 & ~x722 & ~x723 & ~x728 & ~x732 & ~x733 & ~x735 & ~x738 & ~x739 & ~x742 & ~x744 & ~x755 & ~x759 & ~x762 & ~x763 & ~x764 & ~x765 & ~x766 & ~x767 & ~x768 & ~x770 & ~x772 & ~x776 & ~x778 & ~x780 & ~x781 & ~x783;
assign c3111 =  x263 &  x291 &  x348 & ~x0 & ~x6 & ~x7 & ~x8 & ~x21 & ~x24 & ~x30 & ~x35 & ~x39 & ~x44 & ~x51 & ~x60 & ~x64 & ~x75 & ~x80 & ~x97 & ~x112 & ~x113 & ~x117 & ~x142 & ~x145 & ~x147 & ~x148 & ~x167 & ~x170 & ~x175 & ~x176 & ~x199 & ~x203 & ~x221 & ~x222 & ~x223 & ~x225 & ~x252 & ~x256 & ~x260 & ~x280 & ~x313 & ~x314 & ~x343 & ~x419 & ~x420 & ~x449 & ~x471 & ~x502 & ~x503 & ~x507 & ~x557 & ~x558 & ~x560 & ~x561 & ~x565 & ~x582 & ~x587 & ~x592 & ~x637 & ~x638 & ~x644 & ~x646 & ~x667 & ~x669 & ~x670 & ~x674 & ~x676 & ~x691 & ~x694 & ~x695 & ~x697 & ~x701 & ~x702 & ~x706 & ~x719 & ~x721 & ~x726 & ~x728 & ~x732 & ~x733 & ~x742 & ~x749 & ~x752 & ~x753 & ~x759 & ~x778;
assign c3113 =  x154 & ~x0 & ~x4 & ~x11 & ~x12 & ~x20 & ~x26 & ~x38 & ~x39 & ~x46 & ~x49 & ~x51 & ~x52 & ~x53 & ~x54 & ~x56 & ~x59 & ~x60 & ~x73 & ~x74 & ~x75 & ~x76 & ~x78 & ~x80 & ~x87 & ~x90 & ~x109 & ~x111 & ~x115 & ~x135 & ~x136 & ~x137 & ~x139 & ~x141 & ~x163 & ~x164 & ~x170 & ~x199 & ~x223 & ~x225 & ~x226 & ~x227 & ~x251 & ~x252 & ~x257 & ~x282 & ~x292 & ~x306 & ~x307 & ~x311 & ~x321 & ~x322 & ~x332 & ~x335 & ~x350 & ~x363 & ~x421 & ~x447 & ~x448 & ~x477 & ~x479 & ~x504 & ~x530 & ~x532 & ~x585 & ~x615 & ~x617 & ~x618 & ~x647 & ~x668 & ~x676 & ~x679 & ~x682 & ~x685 & ~x690 & ~x697 & ~x702 & ~x703 & ~x708 & ~x711 & ~x723 & ~x733 & ~x738 & ~x741 & ~x746 & ~x761 & ~x762 & ~x763 & ~x769 & ~x774;
assign c3115 = ~x8 & ~x16 & ~x17 & ~x19 & ~x21 & ~x31 & ~x32 & ~x36 & ~x37 & ~x42 & ~x43 & ~x47 & ~x49 & ~x59 & ~x61 & ~x62 & ~x67 & ~x72 & ~x73 & ~x79 & ~x87 & ~x92 & ~x102 & ~x103 & ~x104 & ~x105 & ~x106 & ~x111 & ~x114 & ~x117 & ~x118 & ~x135 & ~x136 & ~x142 & ~x144 & ~x146 & ~x171 & ~x174 & ~x193 & ~x194 & ~x197 & ~x222 & ~x226 & ~x238 & ~x251 & ~x256 & ~x266 & ~x295 & ~x309 & ~x310 & ~x314 & ~x334 & ~x336 & ~x339 & ~x362 & ~x367 & ~x368 & ~x370 & ~x387 & ~x390 & ~x421 & ~x422 & ~x423 & ~x446 & ~x454 & ~x480 & ~x500 & ~x502 & ~x505 & ~x508 & ~x509 & ~x510 & ~x517 & ~x529 & ~x530 & ~x533 & ~x537 & ~x555 & ~x558 & ~x562 & ~x563 & ~x564 & ~x566 & ~x587 & ~x589 & ~x590 & ~x591 & ~x614 & ~x617 & ~x620 & ~x668 & ~x669 & ~x670 & ~x676 & ~x678 & ~x679 & ~x698 & ~x699 & ~x704 & ~x709 & ~x710 & ~x716 & ~x718 & ~x720 & ~x722 & ~x734 & ~x735 & ~x736 & ~x739 & ~x741 & ~x744 & ~x748 & ~x750 & ~x751 & ~x753 & ~x758 & ~x765 & ~x774 & ~x776 & ~x780 & ~x781 & ~x782;
assign c3117 =  x187 & ~x23 & ~x41 & ~x99 & ~x109 & ~x121 & ~x145 & ~x175 & ~x203 & ~x226 & ~x271 & ~x274 & ~x282 & ~x297 & ~x299 & ~x339 & ~x422 & ~x450 & ~x499 & ~x733;
assign c3119 =  x290 &  x345 &  x401 & ~x12 & ~x27 & ~x34 & ~x45 & ~x69 & ~x78 & ~x82 & ~x115 & ~x171 & ~x198 & ~x231 & ~x313 & ~x334 & ~x367 & ~x417 & ~x445 & ~x472 & ~x528 & ~x557 & ~x613 & ~x614 & ~x646 & ~x696 & ~x702 & ~x712 & ~x719;
assign c3121 =  x288 &  x344 &  x373 & ~x62 & ~x196 & ~x200 & ~x527 & ~x722;
assign c3123 =  x289 &  x317 &  x345 &  x375 & ~x1 & ~x23 & ~x30 & ~x43 & ~x52 & ~x56 & ~x78 & ~x87 & ~x90 & ~x92 & ~x99 & ~x102 & ~x106 & ~x224 & ~x253 & ~x310 & ~x365 & ~x422 & ~x448 & ~x450 & ~x451 & ~x452 & ~x474 & ~x503 & ~x530 & ~x586 & ~x589 & ~x743 & ~x746 & ~x748 & ~x767;
assign c3125 =  x438 &  x493 &  x521 & ~x17 & ~x27 & ~x31 & ~x59 & ~x69 & ~x84 & ~x126 & ~x165 & ~x378 & ~x420 & ~x567 & ~x697 & ~x709 & ~x730 & ~x737 & ~x752 & ~x760;
assign c3127 =  x459 &  x487 & ~x44 & ~x79 & ~x81 & ~x173 & ~x201 & ~x211 & ~x426 & ~x530 & ~x712 & ~x749;
assign c3129 =  x490 &  x518 &  x546 &  x602 & ~x14 & ~x30 & ~x39 & ~x71 & ~x98 & ~x130 & ~x142 & ~x223 & ~x282 & ~x418 & ~x531 & ~x625 & ~x644 & ~x665 & ~x672 & ~x678 & ~x682;
assign c3131 =  x316 &  x371 & ~x45 & ~x51 & ~x53 & ~x83 & ~x85 & ~x86 & ~x88 & ~x92 & ~x97 & ~x101 & ~x108 & ~x116 & ~x123 & ~x139 & ~x140 & ~x195 & ~x226 & ~x228 & ~x278 & ~x308 & ~x334 & ~x335 & ~x419 & ~x449 & ~x478 & ~x504 & ~x534 & ~x586 & ~x614 & ~x618 & ~x619 & ~x641 & ~x644 & ~x646 & ~x676 & ~x700 & ~x702 & ~x705 & ~x712 & ~x734 & ~x760 & ~x768 & ~x770 & ~x772;
assign c3133 =  x400 & ~x5 & ~x24 & ~x33 & ~x41 & ~x50 & ~x57 & ~x79 & ~x87 & ~x89 & ~x90 & ~x110 & ~x119 & ~x122 & ~x136 & ~x145 & ~x164 & ~x171 & ~x172 & ~x175 & ~x195 & ~x197 & ~x199 & ~x254 & ~x256 & ~x309 & ~x337 & ~x349 & ~x361 & ~x363 & ~x393 & ~x478 & ~x505 & ~x532 & ~x534 & ~x557 & ~x559 & ~x560 & ~x584 & ~x587 & ~x590 & ~x619 & ~x640 & ~x646 & ~x650 & ~x668 & ~x672 & ~x673 & ~x679 & ~x682 & ~x694 & ~x697 & ~x722 & ~x724 & ~x729 & ~x735 & ~x736 & ~x737 & ~x757 & ~x764 & ~x768 & ~x769 & ~x772 & ~x774 & ~x778 & ~x781;
assign c3135 = ~x2 & ~x7 & ~x8 & ~x10 & ~x14 & ~x16 & ~x18 & ~x19 & ~x23 & ~x25 & ~x27 & ~x30 & ~x33 & ~x34 & ~x38 & ~x39 & ~x41 & ~x42 & ~x43 & ~x44 & ~x46 & ~x51 & ~x52 & ~x58 & ~x59 & ~x64 & ~x70 & ~x72 & ~x78 & ~x81 & ~x86 & ~x90 & ~x92 & ~x105 & ~x107 & ~x110 & ~x111 & ~x112 & ~x116 & ~x118 & ~x122 & ~x135 & ~x143 & ~x162 & ~x167 & ~x168 & ~x171 & ~x193 & ~x194 & ~x197 & ~x198 & ~x219 & ~x222 & ~x224 & ~x225 & ~x246 & ~x249 & ~x251 & ~x253 & ~x255 & ~x256 & ~x279 & ~x281 & ~x283 & ~x304 & ~x306 & ~x330 & ~x336 & ~x338 & ~x358 & ~x364 & ~x366 & ~x390 & ~x393 & ~x418 & ~x420 & ~x421 & ~x450 & ~x451 & ~x478 & ~x505 & ~x506 & ~x507 & ~x533 & ~x534 & ~x558 & ~x559 & ~x560 & ~x565 & ~x584 & ~x587 & ~x589 & ~x592 & ~x596 & ~x603 & ~x604 & ~x612 & ~x613 & ~x632 & ~x640 & ~x643 & ~x644 & ~x646 & ~x647 & ~x648 & ~x651 & ~x661 & ~x669 & ~x670 & ~x673 & ~x674 & ~x676 & ~x677 & ~x678 & ~x696 & ~x699 & ~x705 & ~x706 & ~x717 & ~x718 & ~x728 & ~x731 & ~x732 & ~x745 & ~x746 & ~x752 & ~x755 & ~x760 & ~x762 & ~x766 & ~x767 & ~x768 & ~x769 & ~x770 & ~x772 & ~x774 & ~x776 & ~x782;
assign c3137 =  x291 &  x319 &  x347 &  x375 & ~x1 & ~x10 & ~x16 & ~x18 & ~x25 & ~x30 & ~x32 & ~x33 & ~x36 & ~x43 & ~x45 & ~x54 & ~x57 & ~x68 & ~x73 & ~x76 & ~x79 & ~x89 & ~x92 & ~x100 & ~x107 & ~x118 & ~x144 & ~x148 & ~x170 & ~x171 & ~x174 & ~x197 & ~x200 & ~x231 & ~x282 & ~x286 & ~x309 & ~x338 & ~x365 & ~x367 & ~x389 & ~x415 & ~x416 & ~x423 & ~x443 & ~x445 & ~x447 & ~x450 & ~x471 & ~x472 & ~x473 & ~x475 & ~x478 & ~x529 & ~x531 & ~x555 & ~x560 & ~x582 & ~x589 & ~x592 & ~x641 & ~x645 & ~x649 & ~x665 & ~x668 & ~x669 & ~x672 & ~x673 & ~x678 & ~x692 & ~x697 & ~x705 & ~x720 & ~x725 & ~x746 & ~x751 & ~x752 & ~x753 & ~x757 & ~x765 & ~x769 & ~x770 & ~x779 & ~x780 & ~x783;
assign c3139 =  x431 &  x486 & ~x11 & ~x18 & ~x27 & ~x29 & ~x30 & ~x34 & ~x35 & ~x46 & ~x47 & ~x50 & ~x52 & ~x54 & ~x55 & ~x56 & ~x57 & ~x58 & ~x61 & ~x63 & ~x66 & ~x68 & ~x75 & ~x79 & ~x88 & ~x89 & ~x112 & ~x116 & ~x142 & ~x144 & ~x146 & ~x168 & ~x169 & ~x170 & ~x171 & ~x172 & ~x201 & ~x223 & ~x227 & ~x230 & ~x250 & ~x255 & ~x257 & ~x281 & ~x282 & ~x283 & ~x284 & ~x311 & ~x335 & ~x337 & ~x340 & ~x341 & ~x369 & ~x388 & ~x391 & ~x395 & ~x420 & ~x421 & ~x422 & ~x423 & ~x424 & ~x452 & ~x475 & ~x480 & ~x505 & ~x530 & ~x531 & ~x532 & ~x535 & ~x536 & ~x557 & ~x559 & ~x561 & ~x589 & ~x590 & ~x591 & ~x592 & ~x613 & ~x616 & ~x617 & ~x619 & ~x643 & ~x645 & ~x646 & ~x667 & ~x668 & ~x675 & ~x678 & ~x682 & ~x694 & ~x695 & ~x698 & ~x701 & ~x703 & ~x705 & ~x711 & ~x715 & ~x720 & ~x721 & ~x722 & ~x726 & ~x729 & ~x731 & ~x737 & ~x746 & ~x749 & ~x750 & ~x751 & ~x755 & ~x757 & ~x758 & ~x761 & ~x763 & ~x769 & ~x770 & ~x771 & ~x772 & ~x773 & ~x778 & ~x779 & ~x780 & ~x782;
assign c3141 =  x159 & ~x90 & ~x227 & ~x268 & ~x298 & ~x302 & ~x332 & ~x336 & ~x395 & ~x585 & ~x646 & ~x678 & ~x694 & ~x710 & ~x718 & ~x725 & ~x775;
assign c3143 =  x519 &  x547 & ~x6 & ~x11 & ~x13 & ~x31 & ~x45 & ~x49 & ~x69 & ~x82 & ~x107 & ~x124 & ~x134 & ~x250 & ~x307 & ~x389 & ~x395 & ~x448 & ~x516 & ~x552 & ~x570 & ~x571 & ~x579 & ~x586 & ~x598 & ~x606 & ~x647 & ~x648 & ~x649 & ~x664 & ~x670 & ~x674 & ~x678 & ~x681 & ~x727 & ~x752 & ~x768 & ~x773 & ~x774 & ~x775 & ~x779;
assign c3145 = ~x0 & ~x10 & ~x12 & ~x18 & ~x30 & ~x35 & ~x43 & ~x48 & ~x52 & ~x88 & ~x89 & ~x91 & ~x114 & ~x123 & ~x139 & ~x149 & ~x151 & ~x179 & ~x206 & ~x207 & ~x261 & ~x262 & ~x279 & ~x282 & ~x283 & ~x284 & ~x315 & ~x316 & ~x325 & ~x425 & ~x502 & ~x561 & ~x608 & ~x618 & ~x634 & ~x635 & ~x662 & ~x664 & ~x693 & ~x704 & ~x722 & ~x725 & ~x735 & ~x748 & ~x757 & ~x760 & ~x767 & ~x769;
assign c3147 =  x434 &  x489 &  x516 &  x544 &  x572 & ~x3 & ~x6 & ~x8 & ~x10 & ~x11 & ~x14 & ~x19 & ~x20 & ~x25 & ~x26 & ~x30 & ~x31 & ~x33 & ~x36 & ~x38 & ~x39 & ~x40 & ~x45 & ~x49 & ~x53 & ~x54 & ~x58 & ~x59 & ~x69 & ~x70 & ~x74 & ~x75 & ~x77 & ~x78 & ~x79 & ~x80 & ~x81 & ~x83 & ~x84 & ~x88 & ~x93 & ~x97 & ~x99 & ~x100 & ~x101 & ~x111 & ~x112 & ~x113 & ~x114 & ~x117 & ~x119 & ~x134 & ~x136 & ~x138 & ~x161 & ~x168 & ~x169 & ~x172 & ~x192 & ~x195 & ~x198 & ~x221 & ~x222 & ~x226 & ~x249 & ~x252 & ~x276 & ~x279 & ~x305 & ~x311 & ~x332 & ~x333 & ~x334 & ~x335 & ~x337 & ~x359 & ~x361 & ~x363 & ~x365 & ~x366 & ~x367 & ~x388 & ~x389 & ~x391 & ~x395 & ~x417 & ~x421 & ~x422 & ~x423 & ~x446 & ~x451 & ~x476 & ~x479 & ~x507 & ~x532 & ~x534 & ~x535 & ~x558 & ~x559 & ~x564 & ~x586 & ~x587 & ~x588 & ~x591 & ~x592 & ~x615 & ~x640 & ~x642 & ~x669 & ~x670 & ~x671 & ~x674 & ~x675 & ~x677 & ~x703 & ~x728 & ~x731 & ~x733 & ~x737 & ~x739 & ~x743 & ~x744 & ~x745 & ~x747 & ~x748 & ~x750 & ~x751 & ~x753 & ~x755 & ~x759 & ~x761 & ~x765 & ~x770 & ~x774 & ~x778 & ~x781 & ~x782 & ~x783;
assign c3149 =  x490 &  x543 &  x571 & ~x11 & ~x30 & ~x33 & ~x48 & ~x56 & ~x57 & ~x62 & ~x64 & ~x78 & ~x86 & ~x89 & ~x110 & ~x112 & ~x140 & ~x251 & ~x254 & ~x305 & ~x309 & ~x350 & ~x363 & ~x389 & ~x451 & ~x501 & ~x532 & ~x558 & ~x562 & ~x617 & ~x671 & ~x695 & ~x697 & ~x698 & ~x713 & ~x722 & ~x724 & ~x743 & ~x754 & ~x756 & ~x758 & ~x771 & ~x775 & ~x783;
assign c3151 = ~x15 & ~x17 & ~x54 & ~x65 & ~x77 & ~x78 & ~x79 & ~x93 & ~x100 & ~x114 & ~x122 & ~x129 & ~x130 & ~x132 & ~x150 & ~x155 & ~x158 & ~x194 & ~x279 & ~x281 & ~x283 & ~x307 & ~x340 & ~x388 & ~x432 & ~x445 & ~x447 & ~x449 & ~x480 & ~x506 & ~x535 & ~x551 & ~x554 & ~x580 & ~x634 & ~x635 & ~x637 & ~x646 & ~x671 & ~x697 & ~x698 & ~x756 & ~x759 & ~x760 & ~x774 & ~x780 & ~x782;
assign c3153 =  x605 & ~x6 & ~x23 & ~x47 & ~x50 & ~x62 & ~x115 & ~x162 & ~x171 & ~x194 & ~x196 & ~x255 & ~x357 & ~x366 & ~x384 & ~x391 & ~x440 & ~x469 & ~x495 & ~x507 & ~x509 & ~x531 & ~x536 & ~x619 & ~x643 & ~x646 & ~x656 & ~x673 & ~x684 & ~x685 & ~x695 & ~x702 & ~x703 & ~x708 & ~x712 & ~x723 & ~x725;
assign c3155 = ~x9 & ~x20 & ~x32 & ~x35 & ~x37 & ~x39 & ~x43 & ~x50 & ~x66 & ~x80 & ~x86 & ~x91 & ~x95 & ~x108 & ~x116 & ~x138 & ~x139 & ~x141 & ~x148 & ~x150 & ~x175 & ~x177 & ~x178 & ~x189 & ~x195 & ~x217 & ~x225 & ~x253 & ~x275 & ~x281 & ~x307 & ~x312 & ~x335 & ~x338 & ~x340 & ~x370 & ~x395 & ~x425 & ~x449 & ~x473 & ~x479 & ~x502 & ~x504 & ~x505 & ~x506 & ~x533 & ~x535 & ~x558 & ~x560 & ~x597 & ~x626 & ~x645 & ~x647 & ~x651 & ~x662 & ~x679 & ~x689 & ~x691 & ~x697 & ~x710 & ~x721 & ~x727 & ~x748 & ~x751 & ~x763 & ~x769;
assign c3157 = ~x1 & ~x7 & ~x13 & ~x24 & ~x40 & ~x51 & ~x56 & ~x63 & ~x72 & ~x76 & ~x84 & ~x93 & ~x96 & ~x125 & ~x135 & ~x139 & ~x152 & ~x161 & ~x164 & ~x169 & ~x188 & ~x191 & ~x194 & ~x224 & ~x308 & ~x336 & ~x350 & ~x378 & ~x433 & ~x460 & ~x476 & ~x478 & ~x508 & ~x564 & ~x565 & ~x567 & ~x587 & ~x592 & ~x615 & ~x621 & ~x639 & ~x642 & ~x647 & ~x676 & ~x695 & ~x696 & ~x723 & ~x753 & ~x754 & ~x762 & ~x778;
assign c3159 =  x347 & ~x6 & ~x7 & ~x15 & ~x25 & ~x39 & ~x42 & ~x45 & ~x58 & ~x61 & ~x73 & ~x88 & ~x92 & ~x110 & ~x112 & ~x115 & ~x117 & ~x120 & ~x122 & ~x125 & ~x126 & ~x130 & ~x131 & ~x151 & ~x168 & ~x179 & ~x206 & ~x283 & ~x311 & ~x362 & ~x386 & ~x389 & ~x397 & ~x418 & ~x473 & ~x475 & ~x479 & ~x554 & ~x556 & ~x582 & ~x587 & ~x590 & ~x612 & ~x616 & ~x636 & ~x640 & ~x647 & ~x666 & ~x671 & ~x675 & ~x697 & ~x700 & ~x705 & ~x706 & ~x707 & ~x726 & ~x731 & ~x734 & ~x739 & ~x751 & ~x759 & ~x779;
assign c3161 =  x464 &  x491 & ~x6 & ~x27 & ~x34 & ~x40 & ~x88 & ~x106 & ~x138 & ~x159 & ~x161 & ~x167 & ~x193 & ~x223 & ~x251 & ~x337 & ~x339 & ~x341 & ~x368 & ~x369 & ~x394 & ~x396 & ~x448 & ~x452 & ~x498 & ~x525 & ~x526 & ~x555 & ~x560 & ~x588 & ~x591 & ~x593 & ~x598 & ~x622 & ~x644 & ~x646 & ~x651 & ~x675 & ~x680 & ~x699 & ~x705 & ~x722 & ~x732 & ~x755 & ~x760 & ~x772 & ~x774 & ~x778;
assign c3163 = ~x2 & ~x8 & ~x19 & ~x21 & ~x34 & ~x43 & ~x46 & ~x56 & ~x64 & ~x66 & ~x73 & ~x82 & ~x86 & ~x88 & ~x109 & ~x117 & ~x143 & ~x165 & ~x167 & ~x169 & ~x172 & ~x200 & ~x224 & ~x255 & ~x305 & ~x311 & ~x362 & ~x363 & ~x382 & ~x392 & ~x411 & ~x417 & ~x418 & ~x445 & ~x466 & ~x473 & ~x493 & ~x505 & ~x559 & ~x564 & ~x589 & ~x590 & ~x594 & ~x615 & ~x617 & ~x623 & ~x640 & ~x642 & ~x644 & ~x645 & ~x652 & ~x668 & ~x673 & ~x678 & ~x682 & ~x688 & ~x696 & ~x699 & ~x712 & ~x719 & ~x726 & ~x731 & ~x734 & ~x746 & ~x756 & ~x760 & ~x762 & ~x768 & ~x769 & ~x779;
assign c3165 =  x465 &  x492 & ~x68 & ~x73 & ~x96 & ~x99 & ~x139 & ~x142 & ~x157 & ~x308 & ~x335 & ~x377 & ~x405 & ~x423 & ~x448 & ~x507 & ~x557 & ~x562 & ~x584 & ~x612 & ~x620 & ~x640 & ~x647 & ~x674 & ~x710 & ~x729;
assign c3167 = ~x23 & ~x30 & ~x35 & ~x47 & ~x48 & ~x50 & ~x51 & ~x54 & ~x61 & ~x72 & ~x82 & ~x90 & ~x101 & ~x111 & ~x140 & ~x144 & ~x197 & ~x198 & ~x279 & ~x353 & ~x362 & ~x381 & ~x390 & ~x391 & ~x437 & ~x449 & ~x477 & ~x501 & ~x507 & ~x563 & ~x686 & ~x688 & ~x690 & ~x704 & ~x709 & ~x716 & ~x717 & ~x723 & ~x724 & ~x745 & ~x759 & ~x766 & ~x779;
assign c3169 = ~x8 & ~x14 & ~x57 & ~x96 & ~x99 & ~x126 & ~x146 & ~x147 & ~x148 & ~x176 & ~x198 & ~x202 & ~x204 & ~x222 & ~x226 & ~x227 & ~x231 & ~x259 & ~x269 & ~x270 & ~x271 & ~x273 & ~x275 & ~x277 & ~x287 & ~x310 & ~x344 & ~x395 & ~x396 & ~x421 & ~x422 & ~x424 & ~x451 & ~x453 & ~x470 & ~x498 & ~x501 & ~x536 & ~x553 & ~x673 & ~x702 & ~x706 & ~x709 & ~x712 & ~x741;
assign c3171 =  x287 & ~x5 & ~x10 & ~x11 & ~x12 & ~x13 & ~x18 & ~x23 & ~x38 & ~x47 & ~x50 & ~x66 & ~x67 & ~x68 & ~x69 & ~x73 & ~x78 & ~x79 & ~x80 & ~x85 & ~x88 & ~x93 & ~x94 & ~x96 & ~x100 & ~x107 & ~x109 & ~x113 & ~x116 & ~x119 & ~x140 & ~x145 & ~x169 & ~x251 & ~x252 & ~x277 & ~x281 & ~x390 & ~x422 & ~x434 & ~x448 & ~x461 & ~x475 & ~x504 & ~x505 & ~x559 & ~x613 & ~x614 & ~x616 & ~x617 & ~x618 & ~x643 & ~x644 & ~x670 & ~x679 & ~x697 & ~x698 & ~x705 & ~x706 & ~x734 & ~x752 & ~x753 & ~x755 & ~x757 & ~x760 & ~x762 & ~x770 & ~x774 & ~x775 & ~x783;
assign c3173 = ~x3 & ~x5 & ~x9 & ~x13 & ~x21 & ~x23 & ~x29 & ~x40 & ~x41 & ~x45 & ~x52 & ~x53 & ~x58 & ~x69 & ~x80 & ~x90 & ~x96 & ~x104 & ~x110 & ~x121 & ~x122 & ~x125 & ~x126 & ~x130 & ~x136 & ~x164 & ~x195 & ~x223 & ~x224 & ~x249 & ~x250 & ~x252 & ~x281 & ~x305 & ~x336 & ~x359 & ~x366 & ~x377 & ~x388 & ~x391 & ~x397 & ~x420 & ~x425 & ~x432 & ~x433 & ~x448 & ~x449 & ~x450 & ~x459 & ~x460 & ~x477 & ~x478 & ~x488 & ~x499 & ~x500 & ~x515 & ~x527 & ~x558 & ~x565 & ~x567 & ~x581 & ~x582 & ~x584 & ~x588 & ~x591 & ~x615 & ~x617 & ~x618 & ~x638 & ~x640 & ~x644 & ~x646 & ~x650 & ~x676 & ~x694 & ~x697 & ~x701 & ~x702 & ~x703 & ~x704 & ~x726 & ~x728 & ~x734 & ~x756 & ~x758 & ~x759 & ~x761 & ~x762 & ~x764 & ~x775 & ~x776 & ~x779 & ~x783;
assign c3175 = ~x3 & ~x7 & ~x15 & ~x21 & ~x33 & ~x36 & ~x37 & ~x43 & ~x46 & ~x48 & ~x49 & ~x51 & ~x56 & ~x66 & ~x87 & ~x90 & ~x95 & ~x96 & ~x97 & ~x105 & ~x106 & ~x110 & ~x113 & ~x114 & ~x117 & ~x122 & ~x128 & ~x137 & ~x151 & ~x152 & ~x161 & ~x162 & ~x163 & ~x164 & ~x175 & ~x226 & ~x335 & ~x337 & ~x362 & ~x363 & ~x365 & ~x418 & ~x444 & ~x447 & ~x448 & ~x470 & ~x471 & ~x472 & ~x487 & ~x488 & ~x506 & ~x514 & ~x516 & ~x525 & ~x528 & ~x533 & ~x542 & ~x560 & ~x561 & ~x563 & ~x564 & ~x565 & ~x569 & ~x580 & ~x581 & ~x586 & ~x587 & ~x589 & ~x593 & ~x595 & ~x598 & ~x608 & ~x609 & ~x617 & ~x622 & ~x625 & ~x626 & ~x648 & ~x649 & ~x654 & ~x674 & ~x677 & ~x681 & ~x694 & ~x703 & ~x705 & ~x707 & ~x723 & ~x724 & ~x727 & ~x735 & ~x749 & ~x761 & ~x775;
assign c3177 = ~x10 & ~x15 & ~x16 & ~x28 & ~x35 & ~x43 & ~x45 & ~x55 & ~x63 & ~x85 & ~x88 & ~x92 & ~x117 & ~x120 & ~x143 & ~x146 & ~x166 & ~x174 & ~x197 & ~x216 & ~x219 & ~x239 & ~x241 & ~x268 & ~x337 & ~x421 & ~x445 & ~x506 & ~x526 & ~x527 & ~x531 & ~x560 & ~x585 & ~x612 & ~x614 & ~x617 & ~x642 & ~x651 & ~x652 & ~x654 & ~x665 & ~x670 & ~x671 & ~x714 & ~x735 & ~x736 & ~x738 & ~x740 & ~x741 & ~x751 & ~x752 & ~x755 & ~x761 & ~x763 & ~x764 & ~x765 & ~x771 & ~x775;
assign c3179 =  x286 &  x314 &  x343 & ~x10;
assign c3181 =  x433 &  x460 &  x487 &  x514 &  x541 & ~x2 & ~x15 & ~x31 & ~x36 & ~x41 & ~x50 & ~x56 & ~x58 & ~x60 & ~x65 & ~x75 & ~x76 & ~x78 & ~x82 & ~x113 & ~x114 & ~x115 & ~x141 & ~x165 & ~x167 & ~x199 & ~x249 & ~x250 & ~x277 & ~x285 & ~x305 & ~x313 & ~x335 & ~x336 & ~x339 & ~x340 & ~x394 & ~x395 & ~x423 & ~x425 & ~x439 & ~x447 & ~x505 & ~x531 & ~x666 & ~x671 & ~x674 & ~x687 & ~x689 & ~x690 & ~x718 & ~x722 & ~x727 & ~x737 & ~x748 & ~x750 & ~x751 & ~x753 & ~x754 & ~x766 & ~x775 & ~x777 & ~x782;
assign c3183 =  x372 &  x401 & ~x0 & ~x3 & ~x18 & ~x35 & ~x41 & ~x49 & ~x59 & ~x65 & ~x72 & ~x104 & ~x112 & ~x113 & ~x126 & ~x165 & ~x169 & ~x192 & ~x255 & ~x279 & ~x280 & ~x283 & ~x365 & ~x392 & ~x449 & ~x473 & ~x479 & ~x507 & ~x560 & ~x562 & ~x563 & ~x621 & ~x643 & ~x644 & ~x648 & ~x671 & ~x677 & ~x702 & ~x727 & ~x733 & ~x741 & ~x782;
assign c3185 =  x318 & ~x0 & ~x1 & ~x3 & ~x31 & ~x32 & ~x40 & ~x41 & ~x42 & ~x50 & ~x75 & ~x82 & ~x88 & ~x93 & ~x100 & ~x105 & ~x106 & ~x114 & ~x120 & ~x130 & ~x133 & ~x148 & ~x165 & ~x168 & ~x195 & ~x201 & ~x224 & ~x227 & ~x228 & ~x293 & ~x334 & ~x336 & ~x365 & ~x392 & ~x414 & ~x421 & ~x446 & ~x449 & ~x474 & ~x477 & ~x478 & ~x505 & ~x506 & ~x526 & ~x531 & ~x535 & ~x538 & ~x553 & ~x559 & ~x564 & ~x615 & ~x619 & ~x644 & ~x646 & ~x694 & ~x726 & ~x770 & ~x773 & ~x779 & ~x782;
assign c3187 =  x293 &  x349 & ~x20 & ~x28 & ~x30 & ~x47 & ~x76 & ~x99 & ~x108 & ~x117 & ~x146 & ~x147 & ~x169 & ~x200 & ~x203 & ~x281 & ~x313 & ~x316 & ~x339 & ~x362 & ~x367 & ~x400 & ~x422 & ~x451 & ~x466 & ~x478 & ~x505 & ~x529 & ~x535 & ~x587 & ~x590 & ~x591 & ~x620 & ~x673 & ~x691 & ~x694 & ~x705 & ~x720 & ~x734 & ~x769;
assign c3189 =  x428 & ~x2 & ~x4 & ~x7 & ~x10 & ~x12 & ~x20 & ~x35 & ~x40 & ~x43 & ~x46 & ~x52 & ~x58 & ~x66 & ~x67 & ~x72 & ~x73 & ~x82 & ~x86 & ~x92 & ~x98 & ~x99 & ~x103 & ~x104 & ~x115 & ~x116 & ~x119 & ~x121 & ~x139 & ~x144 & ~x173 & ~x204 & ~x225 & ~x227 & ~x255 & ~x257 & ~x279 & ~x283 & ~x285 & ~x333 & ~x342 & ~x389 & ~x390 & ~x391 & ~x394 & ~x395 & ~x397 & ~x418 & ~x422 & ~x445 & ~x449 & ~x450 & ~x474 & ~x476 & ~x506 & ~x534 & ~x586 & ~x614 & ~x640 & ~x644 & ~x646 & ~x648 & ~x666 & ~x672 & ~x678 & ~x696 & ~x698 & ~x704 & ~x715 & ~x726 & ~x728 & ~x731 & ~x733 & ~x736 & ~x745 & ~x747 & ~x748 & ~x757 & ~x758 & ~x767 & ~x774 & ~x775 & ~x777;
assign c3191 =  x542 & ~x0 & ~x5 & ~x15 & ~x25 & ~x33 & ~x35 & ~x42 & ~x43 & ~x46 & ~x52 & ~x57 & ~x63 & ~x85 & ~x86 & ~x87 & ~x88 & ~x103 & ~x108 & ~x113 & ~x114 & ~x140 & ~x165 & ~x170 & ~x191 & ~x222 & ~x228 & ~x252 & ~x277 & ~x305 & ~x310 & ~x334 & ~x337 & ~x338 & ~x371 & ~x373 & ~x392 & ~x400 & ~x410 & ~x411 & ~x422 & ~x425 & ~x447 & ~x452 & ~x475 & ~x530 & ~x537 & ~x587 & ~x591 & ~x619 & ~x620 & ~x646 & ~x649 & ~x691 & ~x700 & ~x701 & ~x709 & ~x713 & ~x718 & ~x721 & ~x723 & ~x727 & ~x735 & ~x738 & ~x739 & ~x742 & ~x747 & ~x748 & ~x749 & ~x767 & ~x770 & ~x772;
assign c3193 =  x434 &  x461 &  x488 &  x515 &  x543 &  x570 & ~x3 & ~x5 & ~x12 & ~x16 & ~x21 & ~x27 & ~x31 & ~x41 & ~x48 & ~x50 & ~x58 & ~x61 & ~x62 & ~x65 & ~x70 & ~x74 & ~x80 & ~x88 & ~x100 & ~x107 & ~x111 & ~x137 & ~x138 & ~x170 & ~x172 & ~x195 & ~x199 & ~x226 & ~x228 & ~x251 & ~x252 & ~x256 & ~x280 & ~x283 & ~x284 & ~x307 & ~x309 & ~x310 & ~x332 & ~x334 & ~x364 & ~x367 & ~x369 & ~x389 & ~x390 & ~x393 & ~x395 & ~x396 & ~x397 & ~x422 & ~x423 & ~x449 & ~x475 & ~x476 & ~x477 & ~x478 & ~x479 & ~x480 & ~x585 & ~x586 & ~x614 & ~x616 & ~x641 & ~x642 & ~x643 & ~x645 & ~x695 & ~x698 & ~x703 & ~x717 & ~x718 & ~x720 & ~x721 & ~x722 & ~x723 & ~x724 & ~x725 & ~x726 & ~x732 & ~x735 & ~x742 & ~x746 & ~x747 & ~x748 & ~x749 & ~x750 & ~x756 & ~x758 & ~x767 & ~x774 & ~x777;
assign c3195 =  x190 & ~x300;
assign c3197 =  x374 &  x429 &  x457 & ~x137 & ~x201 & ~x203 & ~x257 & ~x258 & ~x418 & ~x506 & ~x669;
assign c3199 =  x374 & ~x4 & ~x9 & ~x10 & ~x12 & ~x14 & ~x15 & ~x17 & ~x18 & ~x19 & ~x21 & ~x22 & ~x23 & ~x26 & ~x30 & ~x39 & ~x41 & ~x44 & ~x49 & ~x59 & ~x60 & ~x61 & ~x63 & ~x65 & ~x66 & ~x69 & ~x72 & ~x80 & ~x83 & ~x87 & ~x88 & ~x92 & ~x94 & ~x97 & ~x105 & ~x108 & ~x110 & ~x114 & ~x123 & ~x141 & ~x142 & ~x167 & ~x173 & ~x176 & ~x197 & ~x200 & ~x225 & ~x227 & ~x229 & ~x250 & ~x252 & ~x253 & ~x254 & ~x257 & ~x276 & ~x278 & ~x279 & ~x280 & ~x282 & ~x284 & ~x303 & ~x306 & ~x310 & ~x311 & ~x322 & ~x332 & ~x334 & ~x339 & ~x360 & ~x361 & ~x393 & ~x422 & ~x423 & ~x445 & ~x447 & ~x448 & ~x450 & ~x454 & ~x472 & ~x477 & ~x479 & ~x498 & ~x500 & ~x506 & ~x529 & ~x530 & ~x532 & ~x534 & ~x536 & ~x555 & ~x561 & ~x563 & ~x564 & ~x586 & ~x589 & ~x592 & ~x612 & ~x613 & ~x615 & ~x617 & ~x637 & ~x638 & ~x640 & ~x665 & ~x668 & ~x669 & ~x695 & ~x697 & ~x698 & ~x724 & ~x725 & ~x730 & ~x731 & ~x732 & ~x733 & ~x735 & ~x748 & ~x750 & ~x751 & ~x754 & ~x763 & ~x764 & ~x769 & ~x773 & ~x774 & ~x781 & ~x783;
assign c3201 = ~x27 & ~x51 & ~x54 & ~x87 & ~x90 & ~x125 & ~x144 & ~x151 & ~x178 & ~x205 & ~x207 & ~x249 & ~x259 & ~x289 & ~x316 & ~x326 & ~x327 & ~x363 & ~x366 & ~x416 & ~x443 & ~x470 & ~x497 & ~x507 & ~x529 & ~x533 & ~x562 & ~x613 & ~x637 & ~x666 & ~x680 & ~x709 & ~x730 & ~x759 & ~x771 & ~x782;
assign c3203 =  x404 &  x431 &  x458 &  x485 & ~x1 & ~x3 & ~x8 & ~x12 & ~x17 & ~x20 & ~x21 & ~x33 & ~x35 & ~x37 & ~x38 & ~x41 & ~x45 & ~x50 & ~x59 & ~x61 & ~x64 & ~x66 & ~x75 & ~x87 & ~x92 & ~x107 & ~x108 & ~x116 & ~x119 & ~x137 & ~x141 & ~x166 & ~x168 & ~x174 & ~x196 & ~x200 & ~x225 & ~x226 & ~x228 & ~x278 & ~x284 & ~x307 & ~x309 & ~x334 & ~x338 & ~x342 & ~x364 & ~x368 & ~x419 & ~x420 & ~x422 & ~x423 & ~x424 & ~x426 & ~x479 & ~x503 & ~x504 & ~x533 & ~x534 & ~x536 & ~x558 & ~x559 & ~x561 & ~x586 & ~x589 & ~x613 & ~x616 & ~x640 & ~x641 & ~x644 & ~x646 & ~x669 & ~x672 & ~x674 & ~x676 & ~x690 & ~x692 & ~x697 & ~x698 & ~x704 & ~x706 & ~x711 & ~x716 & ~x723 & ~x739 & ~x749 & ~x750 & ~x756 & ~x762 & ~x773 & ~x775;
assign c3205 =  x358;
assign c3207 =  x459 &  x486 &  x541 & ~x5 & ~x6 & ~x13 & ~x19 & ~x21 & ~x25 & ~x27 & ~x30 & ~x31 & ~x34 & ~x37 & ~x38 & ~x41 & ~x53 & ~x55 & ~x57 & ~x61 & ~x72 & ~x79 & ~x81 & ~x87 & ~x89 & ~x91 & ~x135 & ~x136 & ~x139 & ~x142 & ~x166 & ~x170 & ~x195 & ~x196 & ~x199 & ~x225 & ~x226 & ~x256 & ~x257 & ~x279 & ~x283 & ~x308 & ~x311 & ~x315 & ~x334 & ~x337 & ~x339 & ~x340 & ~x343 & ~x344 & ~x362 & ~x363 & ~x366 & ~x369 & ~x393 & ~x400 & ~x418 & ~x425 & ~x427 & ~x450 & ~x452 & ~x474 & ~x508 & ~x530 & ~x535 & ~x562 & ~x586 & ~x614 & ~x615 & ~x616 & ~x640 & ~x644 & ~x646 & ~x667 & ~x668 & ~x672 & ~x674 & ~x691 & ~x695 & ~x697 & ~x705 & ~x708 & ~x710 & ~x711 & ~x716 & ~x717 & ~x726 & ~x733 & ~x735 & ~x738 & ~x744 & ~x746 & ~x751 & ~x754 & ~x757 & ~x765 & ~x771 & ~x774 & ~x775 & ~x776 & ~x779 & ~x781 & ~x783;
assign c3209 =  x315 &  x343 & ~x1 & ~x2 & ~x3 & ~x5 & ~x7 & ~x8 & ~x9 & ~x10 & ~x11 & ~x17 & ~x18 & ~x20 & ~x22 & ~x23 & ~x24 & ~x25 & ~x26 & ~x30 & ~x31 & ~x33 & ~x34 & ~x36 & ~x39 & ~x41 & ~x44 & ~x45 & ~x47 & ~x49 & ~x51 & ~x53 & ~x55 & ~x56 & ~x57 & ~x59 & ~x64 & ~x65 & ~x66 & ~x67 & ~x68 & ~x69 & ~x70 & ~x71 & ~x72 & ~x73 & ~x74 & ~x76 & ~x77 & ~x79 & ~x80 & ~x81 & ~x82 & ~x83 & ~x84 & ~x87 & ~x89 & ~x91 & ~x93 & ~x97 & ~x99 & ~x102 & ~x105 & ~x107 & ~x108 & ~x109 & ~x113 & ~x114 & ~x115 & ~x116 & ~x117 & ~x119 & ~x121 & ~x133 & ~x135 & ~x138 & ~x141 & ~x142 & ~x143 & ~x144 & ~x167 & ~x168 & ~x171 & ~x194 & ~x198 & ~x199 & ~x224 & ~x225 & ~x250 & ~x251 & ~x253 & ~x277 & ~x278 & ~x279 & ~x280 & ~x282 & ~x306 & ~x307 & ~x308 & ~x309 & ~x310 & ~x333 & ~x334 & ~x335 & ~x336 & ~x338 & ~x362 & ~x365 & ~x366 & ~x390 & ~x392 & ~x417 & ~x421 & ~x446 & ~x447 & ~x449 & ~x450 & ~x451 & ~x474 & ~x475 & ~x476 & ~x477 & ~x478 & ~x479 & ~x501 & ~x503 & ~x506 & ~x507 & ~x529 & ~x530 & ~x532 & ~x533 & ~x558 & ~x560 & ~x586 & ~x588 & ~x591 & ~x612 & ~x613 & ~x614 & ~x616 & ~x617 & ~x618 & ~x619 & ~x621 & ~x643 & ~x646 & ~x647 & ~x648 & ~x649 & ~x650 & ~x667 & ~x668 & ~x669 & ~x671 & ~x672 & ~x673 & ~x674 & ~x675 & ~x677 & ~x680 & ~x695 & ~x696 & ~x697 & ~x698 & ~x699 & ~x701 & ~x702 & ~x703 & ~x705 & ~x706 & ~x707 & ~x709 & ~x710 & ~x711 & ~x726 & ~x727 & ~x728 & ~x730 & ~x732 & ~x734 & ~x735 & ~x736 & ~x742 & ~x743 & ~x749 & ~x752 & ~x753 & ~x755 & ~x756 & ~x757 & ~x760 & ~x761 & ~x762 & ~x763 & ~x765 & ~x767 & ~x769 & ~x770 & ~x771 & ~x773 & ~x775 & ~x778 & ~x782;
assign c3211 =  x430 &  x456 & ~x1 & ~x6 & ~x10 & ~x13 & ~x14 & ~x23 & ~x29 & ~x30 & ~x31 & ~x35 & ~x40 & ~x46 & ~x48 & ~x57 & ~x58 & ~x59 & ~x61 & ~x65 & ~x73 & ~x81 & ~x87 & ~x92 & ~x111 & ~x116 & ~x118 & ~x139 & ~x140 & ~x141 & ~x143 & ~x144 & ~x145 & ~x163 & ~x169 & ~x170 & ~x172 & ~x192 & ~x193 & ~x195 & ~x197 & ~x198 & ~x200 & ~x223 & ~x252 & ~x253 & ~x256 & ~x281 & ~x305 & ~x310 & ~x312 & ~x335 & ~x336 & ~x339 & ~x364 & ~x388 & ~x393 & ~x394 & ~x422 & ~x423 & ~x446 & ~x449 & ~x450 & ~x451 & ~x472 & ~x474 & ~x501 & ~x503 & ~x504 & ~x532 & ~x533 & ~x617 & ~x642 & ~x646 & ~x647 & ~x649 & ~x677 & ~x678 & ~x679 & ~x683 & ~x684 & ~x686 & ~x688 & ~x690 & ~x694 & ~x701 & ~x702 & ~x703 & ~x705 & ~x707 & ~x708 & ~x710 & ~x711 & ~x712 & ~x715 & ~x722 & ~x725 & ~x726 & ~x732 & ~x744 & ~x745 & ~x752 & ~x753 & ~x757 & ~x763 & ~x765 & ~x769 & ~x771 & ~x773 & ~x775 & ~x776 & ~x779;
assign c3213 =  x429 &  x456 & ~x5 & ~x10 & ~x15 & ~x16 & ~x21 & ~x23 & ~x27 & ~x34 & ~x58 & ~x75 & ~x77 & ~x80 & ~x90 & ~x91 & ~x106 & ~x116 & ~x143 & ~x173 & ~x229 & ~x307 & ~x311 & ~x503 & ~x531 & ~x585 & ~x657 & ~x675 & ~x677 & ~x707 & ~x723 & ~x743 & ~x750 & ~x760 & ~x767;
assign c3215 =  x407 &  x434 &  x461 &  x488 &  x515 &  x570 & ~x5 & ~x6 & ~x13 & ~x23 & ~x25 & ~x32 & ~x50 & ~x52 & ~x68 & ~x70 & ~x73 & ~x86 & ~x88 & ~x105 & ~x115 & ~x143 & ~x169 & ~x195 & ~x276 & ~x283 & ~x312 & ~x331 & ~x332 & ~x336 & ~x340 & ~x369 & ~x370 & ~x400 & ~x421 & ~x425 & ~x440 & ~x443 & ~x448 & ~x501 & ~x614 & ~x641 & ~x645 & ~x671 & ~x673 & ~x675 & ~x696 & ~x700 & ~x741 & ~x754 & ~x755 & ~x757 & ~x761 & ~x771 & ~x774;
assign c3217 =  x461 &  x517 &  x544 &  x572 & ~x2 & ~x37 & ~x102 & ~x107 & ~x112 & ~x163 & ~x167 & ~x192 & ~x196 & ~x273 & ~x283 & ~x301 & ~x335 & ~x340 & ~x384 & ~x394 & ~x419 & ~x475 & ~x478 & ~x481 & ~x535 & ~x618 & ~x675 & ~x699 & ~x701 & ~x717 & ~x718 & ~x728 & ~x729 & ~x748 & ~x762 & ~x768 & ~x770 & ~x773 & ~x777 & ~x780;
assign c3219 =  x374 & ~x7 & ~x10 & ~x21 & ~x27 & ~x41 & ~x46 & ~x49 & ~x51 & ~x59 & ~x81 & ~x84 & ~x86 & ~x88 & ~x90 & ~x92 & ~x95 & ~x112 & ~x113 & ~x118 & ~x121 & ~x148 & ~x194 & ~x204 & ~x228 & ~x323 & ~x337 & ~x339 & ~x340 & ~x366 & ~x367 & ~x394 & ~x416 & ~x421 & ~x422 & ~x424 & ~x451 & ~x474 & ~x478 & ~x499 & ~x505 & ~x534 & ~x559 & ~x562 & ~x620 & ~x648 & ~x696 & ~x697 & ~x723 & ~x726 & ~x736 & ~x753 & ~x763 & ~x764 & ~x766 & ~x769 & ~x775 & ~x782 & ~x783;
assign c3221 = ~x4 & ~x6 & ~x18 & ~x21 & ~x28 & ~x33 & ~x34 & ~x47 & ~x51 & ~x58 & ~x68 & ~x79 & ~x87 & ~x93 & ~x94 & ~x101 & ~x109 & ~x117 & ~x120 & ~x169 & ~x170 & ~x200 & ~x219 & ~x246 & ~x277 & ~x333 & ~x334 & ~x389 & ~x392 & ~x418 & ~x435 & ~x463 & ~x474 & ~x477 & ~x491 & ~x498 & ~x502 & ~x506 & ~x508 & ~x532 & ~x534 & ~x553 & ~x584 & ~x602 & ~x611 & ~x615 & ~x618 & ~x643 & ~x648 & ~x651 & ~x669 & ~x671 & ~x679 & ~x681 & ~x701 & ~x724 & ~x731 & ~x733 & ~x764 & ~x765 & ~x769;
assign c3223 =  x465 & ~x5 & ~x26 & ~x62 & ~x66 & ~x76 & ~x127 & ~x191 & ~x422 & ~x452 & ~x477 & ~x537 & ~x540 & ~x553 & ~x579 & ~x580 & ~x585 & ~x593 & ~x597 & ~x614 & ~x626 & ~x638 & ~x647 & ~x665 & ~x678 & ~x706 & ~x710 & ~x711 & ~x739 & ~x772;
assign c3225 =  x317 &  x345 &  x401 & ~x11 & ~x20 & ~x100 & ~x102 & ~x113 & ~x143 & ~x202 & ~x229 & ~x286 & ~x313 & ~x335 & ~x339 & ~x392 & ~x446 & ~x527 & ~x586 & ~x589 & ~x676 & ~x702 & ~x725 & ~x747 & ~x778 & ~x781;
assign c3227 = ~x11 & ~x13 & ~x21 & ~x24 & ~x29 & ~x36 & ~x44 & ~x75 & ~x77 & ~x95 & ~x100 & ~x124 & ~x127 & ~x140 & ~x148 & ~x150 & ~x173 & ~x183 & ~x277 & ~x336 & ~x361 & ~x415 & ~x452 & ~x453 & ~x498 & ~x501 & ~x504 & ~x505 & ~x507 & ~x509 & ~x578 & ~x587 & ~x592 & ~x608 & ~x670 & ~x691 & ~x714 & ~x748 & ~x766;
assign c3229 = ~x3 & ~x5 & ~x7 & ~x12 & ~x24 & ~x30 & ~x37 & ~x38 & ~x42 & ~x63 & ~x75 & ~x76 & ~x77 & ~x95 & ~x110 & ~x111 & ~x112 & ~x123 & ~x130 & ~x141 & ~x145 & ~x168 & ~x178 & ~x195 & ~x249 & ~x274 & ~x332 & ~x334 & ~x335 & ~x361 & ~x394 & ~x414 & ~x417 & ~x450 & ~x479 & ~x498 & ~x508 & ~x510 & ~x511 & ~x512 & ~x528 & ~x530 & ~x533 & ~x552 & ~x553 & ~x561 & ~x566 & ~x583 & ~x586 & ~x587 & ~x648 & ~x654 & ~x668 & ~x673 & ~x677 & ~x678 & ~x682 & ~x683 & ~x685 & ~x726 & ~x729 & ~x732 & ~x733 & ~x740 & ~x752 & ~x754 & ~x755 & ~x760 & ~x761 & ~x766 & ~x782;
assign c3231 =  x374 & ~x2 & ~x12 & ~x15 & ~x16 & ~x19 & ~x40 & ~x47 & ~x49 & ~x51 & ~x52 & ~x53 & ~x54 & ~x55 & ~x58 & ~x63 & ~x66 & ~x68 & ~x69 & ~x71 & ~x73 & ~x76 & ~x82 & ~x84 & ~x87 & ~x91 & ~x92 & ~x94 & ~x101 & ~x109 & ~x114 & ~x115 & ~x119 & ~x120 & ~x123 & ~x124 & ~x125 & ~x143 & ~x150 & ~x151 & ~x153 & ~x167 & ~x171 & ~x174 & ~x176 & ~x177 & ~x205 & ~x222 & ~x225 & ~x230 & ~x250 & ~x256 & ~x279 & ~x281 & ~x311 & ~x314 & ~x332 & ~x336 & ~x339 & ~x340 & ~x341 & ~x359 & ~x388 & ~x389 & ~x392 & ~x393 & ~x396 & ~x416 & ~x446 & ~x447 & ~x448 & ~x474 & ~x478 & ~x501 & ~x503 & ~x504 & ~x507 & ~x528 & ~x529 & ~x534 & ~x535 & ~x556 & ~x559 & ~x560 & ~x561 & ~x562 & ~x581 & ~x590 & ~x611 & ~x613 & ~x614 & ~x617 & ~x637 & ~x642 & ~x644 & ~x668 & ~x672 & ~x692 & ~x694 & ~x700 & ~x702 & ~x727 & ~x729 & ~x732 & ~x733 & ~x756 & ~x758 & ~x759 & ~x762 & ~x764 & ~x771 & ~x776 & ~x780;
assign c3233 =  x706;
assign c3235 =  x431 &  x458 &  x485 &  x512 & ~x27 & ~x281 & ~x367 & ~x412 & ~x420 & ~x504 & ~x677 & ~x688 & ~x690 & ~x691 & ~x747 & ~x751 & ~x772 & ~x777;
assign c3237 =  x491 &  x519 & ~x13 & ~x36 & ~x38 & ~x70 & ~x76 & ~x170 & ~x171 & ~x250 & ~x253 & ~x280 & ~x284 & ~x308 & ~x342 & ~x364 & ~x365 & ~x366 & ~x392 & ~x395 & ~x446 & ~x476 & ~x508 & ~x533 & ~x559 & ~x564 & ~x590 & ~x615 & ~x628 & ~x642 & ~x655 & ~x675 & ~x683 & ~x698 & ~x712 & ~x721 & ~x746 & ~x749 & ~x762 & ~x769 & ~x775 & ~x778;
assign c3239 = ~x4 & ~x6 & ~x29 & ~x35 & ~x40 & ~x45 & ~x49 & ~x56 & ~x57 & ~x77 & ~x82 & ~x84 & ~x86 & ~x88 & ~x109 & ~x116 & ~x136 & ~x137 & ~x140 & ~x168 & ~x194 & ~x199 & ~x251 & ~x265 & ~x276 & ~x293 & ~x295 & ~x305 & ~x321 & ~x322 & ~x323 & ~x334 & ~x335 & ~x348 & ~x349 & ~x350 & ~x351 & ~x449 & ~x450 & ~x478 & ~x502 & ~x531 & ~x533 & ~x558 & ~x587 & ~x643 & ~x657 & ~x658 & ~x675 & ~x681 & ~x686 & ~x688 & ~x699 & ~x700 & ~x713 & ~x715 & ~x728 & ~x730 & ~x740 & ~x741 & ~x743 & ~x754 & ~x755 & ~x779;
assign c3241 = ~x14 & ~x27 & ~x30 & ~x36 & ~x62 & ~x65 & ~x87 & ~x99 & ~x101 & ~x107 & ~x109 & ~x114 & ~x125 & ~x126 & ~x152 & ~x159 & ~x172 & ~x179 & ~x180 & ~x181 & ~x189 & ~x191 & ~x194 & ~x223 & ~x251 & ~x254 & ~x281 & ~x307 & ~x312 & ~x329 & ~x330 & ~x362 & ~x391 & ~x393 & ~x394 & ~x418 & ~x449 & ~x476 & ~x479 & ~x480 & ~x536 & ~x551 & ~x552 & ~x562 & ~x579 & ~x583 & ~x590 & ~x592 & ~x593 & ~x605 & ~x607 & ~x608 & ~x620 & ~x634 & ~x635 & ~x641 & ~x644 & ~x645 & ~x650 & ~x661 & ~x664 & ~x668 & ~x707 & ~x718 & ~x720 & ~x726 & ~x744 & ~x745 & ~x753 & ~x759 & ~x766 & ~x774;
assign c3243 =  x464 & ~x8 & ~x13 & ~x23 & ~x49 & ~x50 & ~x59 & ~x61 & ~x62 & ~x72 & ~x77 & ~x78 & ~x79 & ~x80 & ~x109 & ~x115 & ~x117 & ~x138 & ~x139 & ~x141 & ~x166 & ~x167 & ~x197 & ~x199 & ~x222 & ~x223 & ~x230 & ~x251 & ~x255 & ~x277 & ~x283 & ~x286 & ~x294 & ~x295 & ~x302 & ~x309 & ~x312 & ~x335 & ~x341 & ~x351 & ~x367 & ~x393 & ~x416 & ~x420 & ~x422 & ~x445 & ~x475 & ~x504 & ~x585 & ~x611 & ~x613 & ~x618 & ~x641 & ~x675 & ~x695 & ~x699 & ~x701 & ~x703 & ~x707 & ~x716 & ~x717 & ~x718 & ~x723 & ~x743 & ~x748 & ~x754 & ~x760 & ~x763 & ~x768 & ~x769 & ~x779;
assign c3245 =  x219 & ~x326;
assign c3247 = ~x3 & ~x7 & ~x14 & ~x18 & ~x23 & ~x31 & ~x34 & ~x37 & ~x50 & ~x53 & ~x56 & ~x62 & ~x67 & ~x69 & ~x73 & ~x76 & ~x82 & ~x100 & ~x118 & ~x127 & ~x131 & ~x133 & ~x142 & ~x144 & ~x147 & ~x153 & ~x154 & ~x158 & ~x169 & ~x176 & ~x178 & ~x183 & ~x194 & ~x223 & ~x278 & ~x279 & ~x303 & ~x304 & ~x336 & ~x417 & ~x476 & ~x506 & ~x509 & ~x515 & ~x526 & ~x540 & ~x542 & ~x560 & ~x589 & ~x590 & ~x591 & ~x594 & ~x608 & ~x610 & ~x617 & ~x648 & ~x649 & ~x650 & ~x667 & ~x670 & ~x674 & ~x675 & ~x678 & ~x694 & ~x701 & ~x706 & ~x723 & ~x729 & ~x731 & ~x732 & ~x735;
assign c3249 =  x543 & ~x60 & ~x281 & ~x283 & ~x361 & ~x391 & ~x439 & ~x480 & ~x536 & ~x564 & ~x630 & ~x657 & ~x659 & ~x660 & ~x670 & ~x671 & ~x689 & ~x690 & ~x719 & ~x745 & ~x756 & ~x771;
assign c3251 = ~x14 & ~x16 & ~x35 & ~x50 & ~x53 & ~x57 & ~x60 & ~x64 & ~x68 & ~x85 & ~x90 & ~x113 & ~x167 & ~x175 & ~x230 & ~x258 & ~x282 & ~x298 & ~x303 & ~x309 & ~x337 & ~x396 & ~x397 & ~x465 & ~x466 & ~x498 & ~x508 & ~x521 & ~x531 & ~x564 & ~x586 & ~x592 & ~x621 & ~x641 & ~x675 & ~x677 & ~x704 & ~x712 & ~x730 & ~x739 & ~x740 & ~x744 & ~x747 & ~x749 & ~x770;
assign c3253 =  x346 & ~x6 & ~x7 & ~x16 & ~x25 & ~x28 & ~x32 & ~x39 & ~x40 & ~x41 & ~x43 & ~x47 & ~x49 & ~x55 & ~x57 & ~x58 & ~x65 & ~x67 & ~x76 & ~x77 & ~x80 & ~x85 & ~x87 & ~x88 & ~x90 & ~x93 & ~x104 & ~x117 & ~x118 & ~x119 & ~x121 & ~x137 & ~x139 & ~x144 & ~x173 & ~x174 & ~x193 & ~x195 & ~x226 & ~x254 & ~x255 & ~x266 & ~x269 & ~x278 & ~x280 & ~x307 & ~x310 & ~x333 & ~x335 & ~x366 & ~x388 & ~x419 & ~x447 & ~x473 & ~x477 & ~x502 & ~x505 & ~x508 & ~x509 & ~x529 & ~x531 & ~x534 & ~x560 & ~x561 & ~x564 & ~x583 & ~x584 & ~x585 & ~x587 & ~x589 & ~x591 & ~x611 & ~x612 & ~x615 & ~x617 & ~x618 & ~x619 & ~x620 & ~x638 & ~x639 & ~x640 & ~x645 & ~x664 & ~x665 & ~x697 & ~x703 & ~x716 & ~x718 & ~x719 & ~x720 & ~x725 & ~x741 & ~x742 & ~x746 & ~x755 & ~x761 & ~x763 & ~x766 & ~x769 & ~x771 & ~x774;
assign c3255 =  x289 &  x345 & ~x7 & ~x21 & ~x26 & ~x35 & ~x39 & ~x46 & ~x53 & ~x62 & ~x70 & ~x74 & ~x76 & ~x80 & ~x82 & ~x100 & ~x106 & ~x140 & ~x144 & ~x146 & ~x169 & ~x174 & ~x221 & ~x310 & ~x312 & ~x361 & ~x446 & ~x517 & ~x612 & ~x672 & ~x734 & ~x761 & ~x778;
assign c3257 =  x416;
assign c3259 = ~x0 & ~x5 & ~x6 & ~x10 & ~x12 & ~x15 & ~x17 & ~x19 & ~x20 & ~x26 & ~x29 & ~x32 & ~x37 & ~x40 & ~x45 & ~x47 & ~x51 & ~x52 & ~x53 & ~x61 & ~x68 & ~x70 & ~x79 & ~x83 & ~x88 & ~x90 & ~x104 & ~x105 & ~x108 & ~x109 & ~x110 & ~x111 & ~x113 & ~x135 & ~x136 & ~x138 & ~x141 & ~x143 & ~x163 & ~x165 & ~x166 & ~x167 & ~x196 & ~x197 & ~x224 & ~x255 & ~x278 & ~x283 & ~x322 & ~x333 & ~x350 & ~x365 & ~x378 & ~x379 & ~x392 & ~x394 & ~x417 & ~x447 & ~x449 & ~x475 & ~x476 & ~x504 & ~x505 & ~x530 & ~x531 & ~x533 & ~x534 & ~x561 & ~x587 & ~x615 & ~x616 & ~x617 & ~x632 & ~x641 & ~x643 & ~x645 & ~x670 & ~x673 & ~x675 & ~x686 & ~x695 & ~x698 & ~x699 & ~x702 & ~x704 & ~x705 & ~x713 & ~x727 & ~x728 & ~x730 & ~x731 & ~x733 & ~x737 & ~x740 & ~x752 & ~x753 & ~x755 & ~x764 & ~x765 & ~x766 & ~x767 & ~x772 & ~x777 & ~x782 & ~x783;
assign c3261 =  x492 &  x519 & ~x2 & ~x9 & ~x14 & ~x16 & ~x60 & ~x79 & ~x90 & ~x130 & ~x138 & ~x142 & ~x143 & ~x145 & ~x159 & ~x479 & ~x532 & ~x533 & ~x541 & ~x552 & ~x565 & ~x578 & ~x592 & ~x609 & ~x613 & ~x638 & ~x640 & ~x647 & ~x650 & ~x664;
assign c3263 =  x434 &  x461 &  x487 &  x513 &  x541 & ~x1 & ~x3 & ~x86 & ~x107 & ~x115 & ~x250 & ~x257 & ~x281 & ~x308 & ~x335 & ~x531 & ~x686 & ~x688 & ~x707 & ~x753 & ~x775;
assign c3265 =  x235 & ~x27 & ~x55 & ~x61 & ~x74 & ~x80 & ~x111 & ~x121 & ~x161 & ~x175 & ~x176 & ~x196 & ~x197 & ~x204 & ~x221 & ~x232 & ~x239 & ~x258 & ~x309 & ~x336 & ~x341 & ~x369 & ~x390 & ~x473 & ~x474 & ~x507 & ~x528 & ~x649 & ~x650 & ~x669 & ~x678 & ~x680 & ~x707 & ~x715 & ~x726 & ~x755 & ~x766 & ~x769 & ~x771 & ~x777;
assign c3267 =  x302 & ~x382;
assign c3269 =  x517 &  x572 &  x600 & ~x47 & ~x57 & ~x62 & ~x73 & ~x76 & ~x81 & ~x97 & ~x100 & ~x136 & ~x138 & ~x140 & ~x173 & ~x192 & ~x224 & ~x255 & ~x337 & ~x359 & ~x424 & ~x449 & ~x480 & ~x498 & ~x503 & ~x508 & ~x533 & ~x538 & ~x561 & ~x568 & ~x569 & ~x593 & ~x594 & ~x620 & ~x645 & ~x650 & ~x676 & ~x728 & ~x750 & ~x756 & ~x761 & ~x780;
assign c3271 =  x490 &  x518 & ~x9 & ~x22 & ~x26 & ~x35 & ~x38 & ~x41 & ~x52 & ~x64 & ~x66 & ~x67 & ~x68 & ~x74 & ~x95 & ~x97 & ~x99 & ~x100 & ~x101 & ~x114 & ~x115 & ~x116 & ~x122 & ~x131 & ~x135 & ~x142 & ~x149 & ~x150 & ~x152 & ~x160 & ~x164 & ~x170 & ~x194 & ~x195 & ~x197 & ~x220 & ~x225 & ~x250 & ~x252 & ~x254 & ~x304 & ~x311 & ~x334 & ~x340 & ~x367 & ~x391 & ~x392 & ~x424 & ~x425 & ~x450 & ~x453 & ~x473 & ~x480 & ~x502 & ~x530 & ~x533 & ~x534 & ~x540 & ~x557 & ~x562 & ~x563 & ~x565 & ~x566 & ~x577 & ~x582 & ~x588 & ~x591 & ~x606 & ~x611 & ~x612 & ~x613 & ~x620 & ~x634 & ~x641 & ~x645 & ~x677 & ~x698 & ~x727 & ~x744 & ~x755 & ~x756 & ~x761 & ~x770 & ~x773 & ~x774 & ~x775 & ~x778 & ~x779;
assign c3273 =  x484 & ~x29 & ~x31 & ~x37 & ~x50 & ~x51 & ~x62 & ~x67 & ~x81 & ~x86 & ~x141 & ~x173 & ~x200 & ~x229 & ~x248 & ~x252 & ~x254 & ~x257 & ~x277 & ~x284 & ~x322 & ~x395 & ~x504 & ~x531 & ~x561 & ~x588 & ~x657 & ~x672 & ~x677 & ~x680 & ~x681 & ~x682 & ~x683 & ~x712 & ~x718 & ~x733 & ~x734 & ~x740 & ~x745 & ~x746 & ~x748 & ~x750 & ~x764 & ~x782;
assign c3275 =  x490 & ~x251 & ~x279 & ~x325 & ~x365 & ~x521 & ~x754;
assign c3277 =  x488 &  x515 & ~x25 & ~x39 & ~x41 & ~x42 & ~x47 & ~x89 & ~x195 & ~x367 & ~x398 & ~x439 & ~x457 & ~x546 & ~x613 & ~x713;
assign c3279 =  x289 & ~x7 & ~x17 & ~x27 & ~x28 & ~x29 & ~x36 & ~x43 & ~x50 & ~x55 & ~x73 & ~x77 & ~x79 & ~x117 & ~x139 & ~x171 & ~x193 & ~x251 & ~x264 & ~x267 & ~x274 & ~x286 & ~x312 & ~x332 & ~x336 & ~x417 & ~x422 & ~x449 & ~x450 & ~x505 & ~x532 & ~x535 & ~x562 & ~x585 & ~x591 & ~x618 & ~x670 & ~x671 & ~x695 & ~x697 & ~x741 & ~x773 & ~x774;
assign c3281 = ~x2 & ~x5 & ~x9 & ~x12 & ~x17 & ~x18 & ~x25 & ~x26 & ~x30 & ~x32 & ~x42 & ~x54 & ~x55 & ~x58 & ~x71 & ~x74 & ~x84 & ~x88 & ~x107 & ~x109 & ~x110 & ~x111 & ~x142 & ~x166 & ~x167 & ~x171 & ~x197 & ~x199 & ~x226 & ~x282 & ~x305 & ~x309 & ~x310 & ~x323 & ~x335 & ~x337 & ~x350 & ~x363 & ~x366 & ~x378 & ~x379 & ~x395 & ~x405 & ~x418 & ~x421 & ~x445 & ~x447 & ~x478 & ~x501 & ~x557 & ~x558 & ~x586 & ~x613 & ~x616 & ~x617 & ~x643 & ~x670 & ~x673 & ~x674 & ~x676 & ~x678 & ~x687 & ~x688 & ~x697 & ~x700 & ~x705 & ~x714 & ~x715 & ~x717 & ~x718 & ~x719 & ~x720 & ~x721 & ~x745 & ~x751 & ~x752 & ~x759 & ~x764 & ~x774 & ~x776 & ~x777 & ~x780;
assign c3283 = ~x1 & ~x7 & ~x9 & ~x10 & ~x11 & ~x15 & ~x16 & ~x25 & ~x26 & ~x28 & ~x30 & ~x33 & ~x36 & ~x37 & ~x39 & ~x40 & ~x45 & ~x47 & ~x51 & ~x55 & ~x60 & ~x62 & ~x64 & ~x66 & ~x73 & ~x78 & ~x79 & ~x83 & ~x87 & ~x88 & ~x89 & ~x93 & ~x112 & ~x115 & ~x116 & ~x117 & ~x118 & ~x139 & ~x140 & ~x142 & ~x144 & ~x146 & ~x165 & ~x166 & ~x168 & ~x171 & ~x173 & ~x194 & ~x195 & ~x199 & ~x201 & ~x203 & ~x222 & ~x249 & ~x251 & ~x252 & ~x253 & ~x255 & ~x257 & ~x258 & ~x267 & ~x277 & ~x281 & ~x282 & ~x287 & ~x309 & ~x310 & ~x311 & ~x312 & ~x335 & ~x336 & ~x339 & ~x350 & ~x351 & ~x362 & ~x367 & ~x368 & ~x391 & ~x393 & ~x422 & ~x474 & ~x477 & ~x478 & ~x504 & ~x529 & ~x533 & ~x534 & ~x560 & ~x561 & ~x562 & ~x586 & ~x589 & ~x613 & ~x614 & ~x641 & ~x646 & ~x647 & ~x649 & ~x650 & ~x651 & ~x670 & ~x672 & ~x676 & ~x677 & ~x679 & ~x680 & ~x682 & ~x693 & ~x695 & ~x704 & ~x706 & ~x707 & ~x708 & ~x709 & ~x710 & ~x716 & ~x717 & ~x721 & ~x724 & ~x725 & ~x738 & ~x741 & ~x747 & ~x748 & ~x754 & ~x759 & ~x762 & ~x766 & ~x768 & ~x772 & ~x773 & ~x781;
assign c3285 = ~x4 & ~x6 & ~x12 & ~x29 & ~x52 & ~x53 & ~x86 & ~x116 & ~x117 & ~x192 & ~x197 & ~x247 & ~x248 & ~x269 & ~x337 & ~x364 & ~x406 & ~x408 & ~x451 & ~x479 & ~x534 & ~x535 & ~x644 & ~x735 & ~x736 & ~x749 & ~x754 & ~x756 & ~x760;
assign c3287 = ~x6 & ~x11 & ~x20 & ~x24 & ~x28 & ~x29 & ~x34 & ~x46 & ~x49 & ~x51 & ~x61 & ~x84 & ~x86 & ~x89 & ~x94 & ~x95 & ~x102 & ~x111 & ~x112 & ~x123 & ~x126 & ~x138 & ~x142 & ~x150 & ~x152 & ~x194 & ~x195 & ~x196 & ~x197 & ~x200 & ~x206 & ~x233 & ~x256 & ~x260 & ~x262 & ~x279 & ~x304 & ~x330 & ~x334 & ~x340 & ~x359 & ~x361 & ~x365 & ~x389 & ~x391 & ~x393 & ~x416 & ~x419 & ~x423 & ~x425 & ~x443 & ~x449 & ~x473 & ~x474 & ~x481 & ~x503 & ~x524 & ~x525 & ~x527 & ~x534 & ~x554 & ~x561 & ~x563 & ~x583 & ~x590 & ~x609 & ~x614 & ~x616 & ~x618 & ~x620 & ~x645 & ~x648 & ~x675 & ~x698 & ~x702 & ~x703 & ~x704 & ~x722 & ~x724 & ~x728 & ~x738 & ~x739 & ~x752 & ~x755 & ~x762 & ~x765 & ~x767 & ~x769 & ~x773 & ~x777;
assign c3289 =  x289 &  x317 &  x345 &  x373 & ~x9 & ~x17 & ~x21 & ~x22 & ~x28 & ~x29 & ~x32 & ~x44 & ~x46 & ~x47 & ~x48 & ~x49 & ~x54 & ~x60 & ~x73 & ~x78 & ~x79 & ~x81 & ~x82 & ~x108 & ~x110 & ~x111 & ~x112 & ~x116 & ~x135 & ~x143 & ~x146 & ~x166 & ~x170 & ~x223 & ~x227 & ~x229 & ~x230 & ~x251 & ~x254 & ~x278 & ~x279 & ~x309 & ~x337 & ~x362 & ~x364 & ~x393 & ~x422 & ~x448 & ~x474 & ~x504 & ~x506 & ~x507 & ~x530 & ~x562 & ~x586 & ~x589 & ~x613 & ~x616 & ~x638 & ~x640 & ~x666 & ~x672 & ~x676 & ~x693 & ~x696 & ~x706 & ~x724 & ~x746 & ~x753 & ~x767 & ~x768 & ~x769;
assign c3291 =  x435 &  x489 &  x517 & ~x11 & ~x61 & ~x83 & ~x84 & ~x167 & ~x190 & ~x191 & ~x228 & ~x255 & ~x309 & ~x316 & ~x327 & ~x343 & ~x397 & ~x423 & ~x447 & ~x450 & ~x476 & ~x566 & ~x587 & ~x619 & ~x641 & ~x648 & ~x679 & ~x689 & ~x690 & ~x703 & ~x707 & ~x708 & ~x717 & ~x719 & ~x729 & ~x735 & ~x736 & ~x747 & ~x749 & ~x750 & ~x752 & ~x756 & ~x766;
assign c3293 =  x488 &  x570 & ~x3 & ~x44 & ~x45 & ~x60 & ~x61 & ~x64 & ~x85 & ~x88 & ~x102 & ~x113 & ~x281 & ~x359 & ~x364 & ~x370 & ~x416 & ~x439 & ~x477 & ~x506 & ~x529 & ~x530 & ~x644 & ~x691 & ~x698 & ~x704 & ~x726 & ~x748 & ~x756 & ~x762;
assign c3295 =  x462 &  x489 &  x517 &  x571 & ~x1 & ~x4 & ~x5 & ~x7 & ~x9 & ~x12 & ~x23 & ~x29 & ~x33 & ~x34 & ~x44 & ~x52 & ~x56 & ~x57 & ~x60 & ~x64 & ~x65 & ~x69 & ~x72 & ~x73 & ~x74 & ~x80 & ~x87 & ~x91 & ~x95 & ~x101 & ~x111 & ~x116 & ~x138 & ~x139 & ~x142 & ~x164 & ~x166 & ~x167 & ~x169 & ~x172 & ~x196 & ~x198 & ~x199 & ~x221 & ~x225 & ~x226 & ~x249 & ~x251 & ~x252 & ~x284 & ~x305 & ~x335 & ~x337 & ~x338 & ~x341 & ~x359 & ~x364 & ~x390 & ~x393 & ~x396 & ~x397 & ~x417 & ~x419 & ~x421 & ~x424 & ~x452 & ~x475 & ~x476 & ~x477 & ~x500 & ~x501 & ~x559 & ~x590 & ~x615 & ~x616 & ~x641 & ~x643 & ~x670 & ~x673 & ~x674 & ~x675 & ~x693 & ~x698 & ~x701 & ~x712 & ~x713 & ~x717 & ~x719 & ~x722 & ~x723 & ~x725 & ~x741 & ~x751 & ~x753 & ~x754 & ~x756 & ~x757 & ~x758 & ~x768 & ~x777 & ~x780 & ~x783;
assign c3297 = ~x1 & ~x4 & ~x17 & ~x27 & ~x31 & ~x35 & ~x42 & ~x44 & ~x46 & ~x63 & ~x86 & ~x96 & ~x97 & ~x98 & ~x103 & ~x143 & ~x169 & ~x193 & ~x222 & ~x223 & ~x251 & ~x282 & ~x306 & ~x334 & ~x337 & ~x352 & ~x380 & ~x408 & ~x461 & ~x613 & ~x639 & ~x647 & ~x665 & ~x666 & ~x724 & ~x734;
assign c3299 =  x315 &  x343 &  x372 &  x373 & ~x4 & ~x16 & ~x19 & ~x41 & ~x72 & ~x84 & ~x129 & ~x131 & ~x144 & ~x199 & ~x333 & ~x445 & ~x446 & ~x448 & ~x475 & ~x503 & ~x505 & ~x616 & ~x643 & ~x736 & ~x741 & ~x755 & ~x774 & ~x775 & ~x777 & ~x780;
assign c40 =  x225;
assign c42 =  x399 &  x425 & ~x295;
assign c44 =  x381 &  x408 &  x409 & ~x19 & ~x67 & ~x74 & ~x88 & ~x96 & ~x101 & ~x138 & ~x194 & ~x209 & ~x264 & ~x276 & ~x334 & ~x417 & ~x475 & ~x516 & ~x541 & ~x557 & ~x569 & ~x587 & ~x588 & ~x620 & ~x625 & ~x626 & ~x643 & ~x653 & ~x655 & ~x682 & ~x707 & ~x709 & ~x710 & ~x738 & ~x739 & ~x747 & ~x753;
assign c46 =  x31;
assign c410 = ~x1 & ~x3 & ~x6 & ~x9 & ~x10 & ~x14 & ~x15 & ~x16 & ~x21 & ~x23 & ~x24 & ~x27 & ~x28 & ~x29 & ~x30 & ~x36 & ~x37 & ~x38 & ~x41 & ~x42 & ~x43 & ~x44 & ~x45 & ~x47 & ~x48 & ~x50 & ~x52 & ~x53 & ~x55 & ~x56 & ~x57 & ~x58 & ~x60 & ~x61 & ~x62 & ~x63 & ~x64 & ~x66 & ~x67 & ~x69 & ~x71 & ~x72 & ~x74 & ~x75 & ~x77 & ~x78 & ~x79 & ~x80 & ~x82 & ~x85 & ~x88 & ~x89 & ~x91 & ~x92 & ~x95 & ~x97 & ~x98 & ~x99 & ~x103 & ~x104 & ~x105 & ~x111 & ~x112 & ~x113 & ~x121 & ~x127 & ~x128 & ~x131 & ~x132 & ~x136 & ~x137 & ~x139 & ~x140 & ~x141 & ~x142 & ~x154 & ~x155 & ~x164 & ~x165 & ~x166 & ~x168 & ~x169 & ~x170 & ~x171 & ~x172 & ~x182 & ~x191 & ~x196 & ~x197 & ~x199 & ~x200 & ~x210 & ~x221 & ~x222 & ~x223 & ~x225 & ~x227 & ~x250 & ~x251 & ~x252 & ~x255 & ~x266 & ~x274 & ~x275 & ~x278 & ~x280 & ~x281 & ~x293 & ~x294 & ~x304 & ~x307 & ~x311 & ~x330 & ~x332 & ~x333 & ~x336 & ~x337 & ~x338 & ~x339 & ~x362 & ~x363 & ~x364 & ~x366 & ~x367 & ~x390 & ~x392 & ~x394 & ~x421 & ~x422 & ~x449 & ~x451 & ~x474 & ~x475 & ~x476 & ~x477 & ~x478 & ~x479 & ~x500 & ~x505 & ~x506 & ~x528 & ~x529 & ~x530 & ~x532 & ~x534 & ~x536 & ~x543 & ~x556 & ~x557 & ~x558 & ~x559 & ~x562 & ~x564 & ~x570 & ~x571 & ~x584 & ~x585 & ~x587 & ~x589 & ~x592 & ~x596 & ~x597 & ~x598 & ~x614 & ~x616 & ~x618 & ~x624 & ~x626 & ~x641 & ~x642 & ~x644 & ~x648 & ~x649 & ~x653 & ~x669 & ~x672 & ~x673 & ~x677 & ~x678 & ~x680 & ~x681 & ~x697 & ~x699 & ~x701 & ~x706 & ~x708 & ~x717 & ~x719 & ~x720 & ~x721 & ~x725 & ~x726 & ~x729 & ~x732 & ~x733 & ~x734 & ~x735 & ~x737 & ~x738 & ~x741 & ~x742 & ~x744 & ~x745 & ~x748 & ~x749 & ~x756 & ~x757 & ~x760 & ~x762 & ~x763 & ~x765 & ~x766 & ~x768 & ~x769 & ~x770 & ~x773 & ~x774 & ~x777 & ~x778 & ~x780 & ~x782;
assign c412 =  x535;
assign c414 =  x762;
assign c416 = ~x4 & ~x9 & ~x14 & ~x15 & ~x17 & ~x21 & ~x23 & ~x24 & ~x25 & ~x26 & ~x32 & ~x33 & ~x35 & ~x37 & ~x38 & ~x39 & ~x41 & ~x44 & ~x47 & ~x49 & ~x50 & ~x52 & ~x55 & ~x61 & ~x64 & ~x65 & ~x68 & ~x70 & ~x72 & ~x74 & ~x76 & ~x78 & ~x81 & ~x82 & ~x84 & ~x86 & ~x87 & ~x91 & ~x94 & ~x95 & ~x97 & ~x100 & ~x101 & ~x103 & ~x104 & ~x106 & ~x115 & ~x116 & ~x118 & ~x120 & ~x125 & ~x133 & ~x135 & ~x137 & ~x141 & ~x143 & ~x146 & ~x153 & ~x168 & ~x169 & ~x171 & ~x181 & ~x191 & ~x192 & ~x194 & ~x195 & ~x197 & ~x198 & ~x200 & ~x201 & ~x209 & ~x221 & ~x224 & ~x228 & ~x229 & ~x236 & ~x246 & ~x251 & ~x252 & ~x274 & ~x278 & ~x279 & ~x282 & ~x284 & ~x301 & ~x304 & ~x305 & ~x308 & ~x310 & ~x312 & ~x332 & ~x336 & ~x337 & ~x338 & ~x358 & ~x366 & ~x386 & ~x390 & ~x392 & ~x393 & ~x416 & ~x418 & ~x419 & ~x422 & ~x444 & ~x449 & ~x452 & ~x474 & ~x475 & ~x477 & ~x479 & ~x500 & ~x502 & ~x506 & ~x527 & ~x528 & ~x532 & ~x536 & ~x538 & ~x539 & ~x555 & ~x557 & ~x559 & ~x561 & ~x564 & ~x565 & ~x568 & ~x583 & ~x585 & ~x586 & ~x589 & ~x590 & ~x593 & ~x594 & ~x598 & ~x610 & ~x614 & ~x615 & ~x618 & ~x621 & ~x622 & ~x627 & ~x652 & ~x653 & ~x666 & ~x667 & ~x668 & ~x669 & ~x677 & ~x681 & ~x682 & ~x685 & ~x694 & ~x697 & ~x698 & ~x702 & ~x711 & ~x721 & ~x723 & ~x725 & ~x728 & ~x733 & ~x734 & ~x735 & ~x736 & ~x739 & ~x740 & ~x742 & ~x749 & ~x750 & ~x753 & ~x755 & ~x761 & ~x762 & ~x765 & ~x766 & ~x768 & ~x770 & ~x772 & ~x773 & ~x776 & ~x777;
assign c418 = ~x1 & ~x8 & ~x9 & ~x10 & ~x11 & ~x13 & ~x21 & ~x22 & ~x23 & ~x25 & ~x26 & ~x30 & ~x31 & ~x34 & ~x42 & ~x44 & ~x45 & ~x46 & ~x50 & ~x53 & ~x57 & ~x61 & ~x62 & ~x63 & ~x66 & ~x68 & ~x69 & ~x70 & ~x71 & ~x72 & ~x76 & ~x77 & ~x82 & ~x85 & ~x87 & ~x89 & ~x92 & ~x93 & ~x96 & ~x97 & ~x103 & ~x104 & ~x106 & ~x109 & ~x110 & ~x112 & ~x115 & ~x128 & ~x129 & ~x131 & ~x136 & ~x137 & ~x139 & ~x140 & ~x143 & ~x144 & ~x148 & ~x150 & ~x157 & ~x167 & ~x169 & ~x170 & ~x171 & ~x173 & ~x185 & ~x196 & ~x200 & ~x222 & ~x225 & ~x226 & ~x229 & ~x250 & ~x253 & ~x254 & ~x268 & ~x278 & ~x283 & ~x295 & ~x306 & ~x310 & ~x322 & ~x323 & ~x350 & ~x351 & ~x388 & ~x389 & ~x394 & ~x415 & ~x419 & ~x444 & ~x448 & ~x450 & ~x471 & ~x474 & ~x476 & ~x477 & ~x500 & ~x501 & ~x502 & ~x506 & ~x530 & ~x531 & ~x534 & ~x536 & ~x537 & ~x553 & ~x559 & ~x563 & ~x580 & ~x584 & ~x585 & ~x589 & ~x590 & ~x592 & ~x593 & ~x594 & ~x612 & ~x614 & ~x615 & ~x621 & ~x639 & ~x641 & ~x648 & ~x664 & ~x665 & ~x668 & ~x670 & ~x676 & ~x677 & ~x695 & ~x707 & ~x719 & ~x720 & ~x721 & ~x723 & ~x724 & ~x731 & ~x733 & ~x735 & ~x736 & ~x742 & ~x747 & ~x750 & ~x757 & ~x759 & ~x767 & ~x770 & ~x774 & ~x777 & ~x781;
assign c420 =  x300 &  x464 &  x465 & ~x129 & ~x130 & ~x131 & ~x185 & ~x241 & ~x242 & ~x323 & ~x757;
assign c422 =  x461 &  x464 &  x465 & ~x0 & ~x1 & ~x4 & ~x6 & ~x17 & ~x34 & ~x35 & ~x39 & ~x40 & ~x43 & ~x45 & ~x48 & ~x52 & ~x57 & ~x63 & ~x66 & ~x69 & ~x71 & ~x73 & ~x78 & ~x80 & ~x81 & ~x82 & ~x85 & ~x87 & ~x91 & ~x93 & ~x94 & ~x96 & ~x101 & ~x102 & ~x108 & ~x109 & ~x113 & ~x115 & ~x119 & ~x121 & ~x122 & ~x131 & ~x134 & ~x140 & ~x146 & ~x149 & ~x163 & ~x165 & ~x168 & ~x169 & ~x170 & ~x171 & ~x173 & ~x174 & ~x175 & ~x190 & ~x196 & ~x197 & ~x199 & ~x223 & ~x245 & ~x246 & ~x250 & ~x256 & ~x272 & ~x273 & ~x274 & ~x275 & ~x279 & ~x300 & ~x308 & ~x312 & ~x313 & ~x329 & ~x331 & ~x336 & ~x340 & ~x341 & ~x355 & ~x357 & ~x360 & ~x362 & ~x363 & ~x364 & ~x391 & ~x392 & ~x417 & ~x418 & ~x419 & ~x420 & ~x421 & ~x422 & ~x446 & ~x448 & ~x449 & ~x473 & ~x501 & ~x502 & ~x507 & ~x529 & ~x553 & ~x554 & ~x555 & ~x556 & ~x560 & ~x564 & ~x565 & ~x567 & ~x568 & ~x570 & ~x571 & ~x581 & ~x583 & ~x588 & ~x593 & ~x598 & ~x617 & ~x621 & ~x648 & ~x650 & ~x653 & ~x670 & ~x677 & ~x683 & ~x697 & ~x698 & ~x699 & ~x700 & ~x707 & ~x709 & ~x720 & ~x722 & ~x726 & ~x730 & ~x731 & ~x739 & ~x746 & ~x749 & ~x752 & ~x755 & ~x760 & ~x761 & ~x766 & ~x771 & ~x774 & ~x775 & ~x780;
assign c424 =  x460 &  x465 & ~x4 & ~x6 & ~x11 & ~x12 & ~x17 & ~x19 & ~x22 & ~x24 & ~x27 & ~x31 & ~x36 & ~x40 & ~x42 & ~x47 & ~x51 & ~x52 & ~x62 & ~x66 & ~x67 & ~x74 & ~x85 & ~x88 & ~x90 & ~x92 & ~x105 & ~x111 & ~x113 & ~x119 & ~x122 & ~x138 & ~x139 & ~x148 & ~x170 & ~x171 & ~x173 & ~x197 & ~x201 & ~x214 & ~x221 & ~x223 & ~x224 & ~x225 & ~x230 & ~x242 & ~x245 & ~x251 & ~x255 & ~x257 & ~x285 & ~x287 & ~x307 & ~x309 & ~x310 & ~x340 & ~x361 & ~x364 & ~x369 & ~x389 & ~x417 & ~x418 & ~x419 & ~x449 & ~x475 & ~x476 & ~x500 & ~x527 & ~x534 & ~x539 & ~x544 & ~x553 & ~x558 & ~x560 & ~x563 & ~x566 & ~x568 & ~x570 & ~x580 & ~x583 & ~x584 & ~x585 & ~x586 & ~x588 & ~x589 & ~x591 & ~x593 & ~x596 & ~x598 & ~x611 & ~x618 & ~x622 & ~x624 & ~x626 & ~x639 & ~x640 & ~x641 & ~x650 & ~x666 & ~x669 & ~x692 & ~x694 & ~x696 & ~x702 & ~x704 & ~x719 & ~x723 & ~x732 & ~x735 & ~x740 & ~x743 & ~x746 & ~x752 & ~x757 & ~x764 & ~x771 & ~x772 & ~x774 & ~x776 & ~x780 & ~x781 & ~x782;
assign c426 = ~x8 & ~x9 & ~x10 & ~x11 & ~x12 & ~x13 & ~x14 & ~x16 & ~x18 & ~x22 & ~x23 & ~x26 & ~x29 & ~x35 & ~x41 & ~x46 & ~x53 & ~x57 & ~x60 & ~x62 & ~x65 & ~x67 & ~x68 & ~x70 & ~x76 & ~x77 & ~x83 & ~x87 & ~x91 & ~x93 & ~x95 & ~x97 & ~x102 & ~x103 & ~x104 & ~x105 & ~x106 & ~x110 & ~x111 & ~x112 & ~x113 & ~x114 & ~x115 & ~x117 & ~x120 & ~x132 & ~x138 & ~x139 & ~x140 & ~x145 & ~x149 & ~x162 & ~x163 & ~x164 & ~x166 & ~x167 & ~x168 & ~x184 & ~x191 & ~x192 & ~x193 & ~x194 & ~x197 & ~x198 & ~x199 & ~x211 & ~x223 & ~x224 & ~x225 & ~x249 & ~x257 & ~x259 & ~x266 & ~x278 & ~x281 & ~x286 & ~x294 & ~x306 & ~x308 & ~x310 & ~x321 & ~x322 & ~x331 & ~x332 & ~x340 & ~x360 & ~x364 & ~x368 & ~x388 & ~x390 & ~x393 & ~x418 & ~x420 & ~x444 & ~x446 & ~x448 & ~x449 & ~x474 & ~x476 & ~x500 & ~x501 & ~x503 & ~x504 & ~x507 & ~x509 & ~x526 & ~x527 & ~x530 & ~x531 & ~x534 & ~x535 & ~x537 & ~x555 & ~x560 & ~x561 & ~x562 & ~x563 & ~x564 & ~x570 & ~x571 & ~x585 & ~x593 & ~x598 & ~x599 & ~x610 & ~x611 & ~x612 & ~x616 & ~x619 & ~x620 & ~x622 & ~x623 & ~x624 & ~x626 & ~x627 & ~x645 & ~x646 & ~x649 & ~x652 & ~x654 & ~x655 & ~x672 & ~x674 & ~x677 & ~x678 & ~x679 & ~x681 & ~x682 & ~x692 & ~x697 & ~x699 & ~x701 & ~x703 & ~x706 & ~x708 & ~x723 & ~x726 & ~x730 & ~x732 & ~x735 & ~x736 & ~x737 & ~x741 & ~x743 & ~x744 & ~x746 & ~x748 & ~x753 & ~x762 & ~x763 & ~x766 & ~x767 & ~x768 & ~x769 & ~x772 & ~x775 & ~x778 & ~x781 & ~x783;
assign c428 =  x382 & ~x0 & ~x1 & ~x5 & ~x6 & ~x10 & ~x17 & ~x19 & ~x22 & ~x23 & ~x25 & ~x34 & ~x41 & ~x42 & ~x47 & ~x56 & ~x58 & ~x62 & ~x66 & ~x72 & ~x73 & ~x74 & ~x78 & ~x80 & ~x86 & ~x87 & ~x94 & ~x96 & ~x97 & ~x98 & ~x100 & ~x103 & ~x107 & ~x111 & ~x113 & ~x115 & ~x118 & ~x120 & ~x121 & ~x124 & ~x128 & ~x142 & ~x146 & ~x149 & ~x157 & ~x158 & ~x163 & ~x170 & ~x174 & ~x196 & ~x198 & ~x203 & ~x213 & ~x225 & ~x226 & ~x241 & ~x251 & ~x254 & ~x255 & ~x268 & ~x280 & ~x306 & ~x311 & ~x323 & ~x335 & ~x336 & ~x339 & ~x341 & ~x359 & ~x362 & ~x368 & ~x396 & ~x417 & ~x418 & ~x420 & ~x424 & ~x445 & ~x448 & ~x451 & ~x479 & ~x480 & ~x506 & ~x540 & ~x558 & ~x562 & ~x587 & ~x592 & ~x607 & ~x639 & ~x645 & ~x664 & ~x672 & ~x675 & ~x691 & ~x699 & ~x700 & ~x704 & ~x717 & ~x722 & ~x724 & ~x726 & ~x727 & ~x729 & ~x744 & ~x752 & ~x766 & ~x772 & ~x776 & ~x777 & ~x778;
assign c430 =  x345 &  x464 &  x467 &  x491 & ~x89 & ~x99 & ~x125 & ~x143 & ~x149 & ~x150 & ~x151 & ~x200 & ~x233 & ~x254 & ~x255 & ~x257 & ~x285 & ~x287 & ~x303 & ~x332 & ~x341 & ~x360 & ~x368 & ~x477 & ~x567 & ~x624 & ~x642 & ~x645 & ~x671 & ~x673 & ~x720 & ~x771;
assign c432 =  x241 &  x408 & ~x0 & ~x1 & ~x2 & ~x13 & ~x15 & ~x24 & ~x28 & ~x30 & ~x33 & ~x43 & ~x44 & ~x46 & ~x52 & ~x54 & ~x65 & ~x70 & ~x72 & ~x74 & ~x76 & ~x77 & ~x88 & ~x89 & ~x95 & ~x99 & ~x100 & ~x103 & ~x105 & ~x110 & ~x111 & ~x116 & ~x119 & ~x121 & ~x122 & ~x126 & ~x127 & ~x140 & ~x144 & ~x154 & ~x155 & ~x166 & ~x167 & ~x193 & ~x196 & ~x198 & ~x199 & ~x202 & ~x210 & ~x220 & ~x225 & ~x274 & ~x280 & ~x285 & ~x286 & ~x305 & ~x306 & ~x308 & ~x312 & ~x333 & ~x335 & ~x338 & ~x390 & ~x393 & ~x394 & ~x420 & ~x421 & ~x449 & ~x451 & ~x478 & ~x500 & ~x502 & ~x526 & ~x529 & ~x533 & ~x539 & ~x541 & ~x552 & ~x553 & ~x559 & ~x565 & ~x566 & ~x571 & ~x582 & ~x583 & ~x586 & ~x591 & ~x592 & ~x598 & ~x610 & ~x615 & ~x621 & ~x624 & ~x626 & ~x640 & ~x641 & ~x644 & ~x645 & ~x652 & ~x653 & ~x665 & ~x675 & ~x682 & ~x693 & ~x696 & ~x700 & ~x704 & ~x711 & ~x721 & ~x724 & ~x726 & ~x727 & ~x730 & ~x732 & ~x736 & ~x741 & ~x742 & ~x744 & ~x745 & ~x750 & ~x757 & ~x760 & ~x762 & ~x763 & ~x766 & ~x771 & ~x773;
assign c434 =  x352 &  x374 &  x380 &  x402 &  x431 &  x434 &  x462 &  x490 & ~x2 & ~x4 & ~x5 & ~x7 & ~x14 & ~x21 & ~x22 & ~x28 & ~x33 & ~x36 & ~x37 & ~x39 & ~x41 & ~x44 & ~x46 & ~x49 & ~x52 & ~x54 & ~x62 & ~x64 & ~x65 & ~x69 & ~x72 & ~x74 & ~x82 & ~x83 & ~x84 & ~x87 & ~x95 & ~x97 & ~x101 & ~x102 & ~x103 & ~x105 & ~x108 & ~x109 & ~x113 & ~x114 & ~x116 & ~x117 & ~x121 & ~x137 & ~x140 & ~x141 & ~x142 & ~x147 & ~x148 & ~x150 & ~x173 & ~x176 & ~x177 & ~x198 & ~x203 & ~x204 & ~x218 & ~x221 & ~x229 & ~x232 & ~x248 & ~x253 & ~x258 & ~x273 & ~x277 & ~x279 & ~x281 & ~x284 & ~x302 & ~x308 & ~x310 & ~x311 & ~x313 & ~x327 & ~x329 & ~x334 & ~x335 & ~x341 & ~x361 & ~x369 & ~x387 & ~x389 & ~x390 & ~x394 & ~x395 & ~x416 & ~x418 & ~x419 & ~x421 & ~x423 & ~x450 & ~x451 & ~x477 & ~x479 & ~x501 & ~x505 & ~x506 & ~x507 & ~x529 & ~x532 & ~x533 & ~x534 & ~x535 & ~x541 & ~x556 & ~x562 & ~x565 & ~x567 & ~x579 & ~x581 & ~x584 & ~x586 & ~x589 & ~x607 & ~x608 & ~x610 & ~x613 & ~x634 & ~x637 & ~x641 & ~x643 & ~x667 & ~x668 & ~x670 & ~x672 & ~x673 & ~x675 & ~x690 & ~x694 & ~x695 & ~x697 & ~x699 & ~x700 & ~x703 & ~x707 & ~x709 & ~x710 & ~x721 & ~x723 & ~x725 & ~x729 & ~x734 & ~x735 & ~x738 & ~x739 & ~x744 & ~x747 & ~x753 & ~x756 & ~x758 & ~x761 & ~x774 & ~x779 & ~x780;
assign c436 =  x724;
assign c438 =  x409 & ~x3 & ~x4 & ~x8 & ~x10 & ~x11 & ~x17 & ~x20 & ~x23 & ~x24 & ~x25 & ~x26 & ~x30 & ~x32 & ~x36 & ~x39 & ~x47 & ~x48 & ~x52 & ~x54 & ~x56 & ~x64 & ~x66 & ~x67 & ~x69 & ~x70 & ~x72 & ~x74 & ~x76 & ~x77 & ~x81 & ~x83 & ~x86 & ~x87 & ~x88 & ~x90 & ~x92 & ~x93 & ~x95 & ~x96 & ~x98 & ~x100 & ~x101 & ~x104 & ~x105 & ~x109 & ~x110 & ~x114 & ~x116 & ~x128 & ~x131 & ~x132 & ~x139 & ~x140 & ~x141 & ~x152 & ~x158 & ~x166 & ~x168 & ~x175 & ~x194 & ~x197 & ~x205 & ~x223 & ~x224 & ~x226 & ~x227 & ~x228 & ~x231 & ~x251 & ~x253 & ~x255 & ~x257 & ~x268 & ~x278 & ~x282 & ~x283 & ~x284 & ~x285 & ~x286 & ~x296 & ~x306 & ~x307 & ~x308 & ~x313 & ~x335 & ~x337 & ~x338 & ~x362 & ~x363 & ~x366 & ~x367 & ~x388 & ~x390 & ~x394 & ~x395 & ~x446 & ~x452 & ~x470 & ~x473 & ~x477 & ~x480 & ~x497 & ~x498 & ~x499 & ~x500 & ~x503 & ~x505 & ~x506 & ~x507 & ~x528 & ~x530 & ~x532 & ~x534 & ~x557 & ~x560 & ~x564 & ~x580 & ~x582 & ~x583 & ~x584 & ~x585 & ~x586 & ~x587 & ~x588 & ~x590 & ~x609 & ~x616 & ~x637 & ~x640 & ~x641 & ~x643 & ~x646 & ~x647 & ~x650 & ~x663 & ~x665 & ~x672 & ~x675 & ~x677 & ~x688 & ~x689 & ~x691 & ~x692 & ~x696 & ~x698 & ~x700 & ~x703 & ~x715 & ~x717 & ~x718 & ~x719 & ~x721 & ~x726 & ~x728 & ~x734 & ~x740 & ~x743 & ~x754 & ~x756 & ~x757 & ~x760 & ~x765 & ~x772 & ~x773 & ~x780 & ~x783;
assign c440 =  x347 &  x407 &  x435 &  x436 & ~x8 & ~x11 & ~x33 & ~x43 & ~x49 & ~x54 & ~x62 & ~x63 & ~x67 & ~x68 & ~x80 & ~x96 & ~x97 & ~x108 & ~x122 & ~x123 & ~x124 & ~x140 & ~x148 & ~x153 & ~x167 & ~x168 & ~x169 & ~x174 & ~x188 & ~x189 & ~x190 & ~x191 & ~x194 & ~x197 & ~x209 & ~x227 & ~x229 & ~x244 & ~x245 & ~x258 & ~x272 & ~x273 & ~x277 & ~x281 & ~x303 & ~x310 & ~x327 & ~x364 & ~x368 & ~x418 & ~x423 & ~x473 & ~x478 & ~x499 & ~x503 & ~x528 & ~x531 & ~x534 & ~x537 & ~x557 & ~x558 & ~x580 & ~x583 & ~x586 & ~x594 & ~x596 & ~x618 & ~x649 & ~x667 & ~x693 & ~x694 & ~x697 & ~x701 & ~x703 & ~x708 & ~x712 & ~x723 & ~x724 & ~x732 & ~x735 & ~x736 & ~x738 & ~x740 & ~x742 & ~x743 & ~x750 & ~x763 & ~x770 & ~x771 & ~x780;
assign c442 =  x638;
assign c444 =  x346 & ~x13 & ~x101 & ~x124 & ~x165 & ~x187 & ~x232 & ~x233 & ~x242 & ~x256 & ~x258 & ~x259 & ~x270 & ~x283 & ~x284 & ~x447 & ~x505 & ~x512 & ~x527 & ~x549 & ~x576 & ~x605 & ~x618 & ~x642 & ~x660 & ~x661 & ~x688 & ~x716 & ~x718 & ~x730 & ~x735 & ~x736 & ~x739 & ~x745 & ~x747 & ~x749 & ~x760 & ~x765 & ~x769 & ~x781;
assign c446 =  x296 &  x352 &  x463 &  x464 & ~x0 & ~x1 & ~x2 & ~x4 & ~x11 & ~x20 & ~x28 & ~x29 & ~x31 & ~x35 & ~x38 & ~x39 & ~x44 & ~x45 & ~x50 & ~x56 & ~x57 & ~x58 & ~x59 & ~x61 & ~x64 & ~x66 & ~x70 & ~x71 & ~x72 & ~x73 & ~x75 & ~x80 & ~x84 & ~x85 & ~x92 & ~x94 & ~x98 & ~x105 & ~x108 & ~x109 & ~x111 & ~x112 & ~x114 & ~x115 & ~x117 & ~x120 & ~x121 & ~x122 & ~x126 & ~x137 & ~x138 & ~x139 & ~x140 & ~x142 & ~x143 & ~x164 & ~x165 & ~x167 & ~x191 & ~x198 & ~x201 & ~x203 & ~x217 & ~x220 & ~x221 & ~x227 & ~x243 & ~x247 & ~x250 & ~x252 & ~x254 & ~x256 & ~x274 & ~x280 & ~x282 & ~x284 & ~x286 & ~x300 & ~x301 & ~x304 & ~x305 & ~x307 & ~x308 & ~x312 & ~x327 & ~x334 & ~x339 & ~x355 & ~x358 & ~x360 & ~x361 & ~x365 & ~x396 & ~x397 & ~x417 & ~x421 & ~x422 & ~x424 & ~x445 & ~x448 & ~x450 & ~x472 & ~x473 & ~x474 & ~x501 & ~x502 & ~x503 & ~x505 & ~x508 & ~x509 & ~x510 & ~x529 & ~x533 & ~x537 & ~x557 & ~x562 & ~x564 & ~x569 & ~x585 & ~x586 & ~x589 & ~x593 & ~x595 & ~x597 & ~x610 & ~x611 & ~x615 & ~x617 & ~x644 & ~x650 & ~x651 & ~x652 & ~x656 & ~x667 & ~x668 & ~x669 & ~x683 & ~x684 & ~x697 & ~x701 & ~x702 & ~x707 & ~x712 & ~x713 & ~x714 & ~x717 & ~x719 & ~x725 & ~x726 & ~x727 & ~x728 & ~x730 & ~x731 & ~x732 & ~x737 & ~x739 & ~x741 & ~x743 & ~x745 & ~x749 & ~x756 & ~x767 & ~x768 & ~x771 & ~x776 & ~x779;
assign c448 =  x456 &  x464 &  x488 &  x490 &  x516 &  x517 & ~x377 & ~x385 & ~x746;
assign c450 =  x401 &  x411 &  x435 & ~x5 & ~x9 & ~x30 & ~x49 & ~x66 & ~x69 & ~x72 & ~x76 & ~x92 & ~x99 & ~x110 & ~x115 & ~x147 & ~x153 & ~x252 & ~x255 & ~x281 & ~x286 & ~x309 & ~x336 & ~x390 & ~x450 & ~x514 & ~x525 & ~x526 & ~x529 & ~x540 & ~x554 & ~x555 & ~x560 & ~x568 & ~x641 & ~x642 & ~x655 & ~x670 & ~x713 & ~x719 & ~x746 & ~x764;
assign c452 =  x374 &  x429 & ~x2 & ~x3 & ~x7 & ~x8 & ~x11 & ~x12 & ~x13 & ~x15 & ~x16 & ~x19 & ~x20 & ~x26 & ~x29 & ~x30 & ~x31 & ~x32 & ~x33 & ~x38 & ~x41 & ~x42 & ~x43 & ~x44 & ~x49 & ~x52 & ~x53 & ~x63 & ~x65 & ~x70 & ~x71 & ~x72 & ~x73 & ~x75 & ~x76 & ~x79 & ~x80 & ~x82 & ~x83 & ~x85 & ~x86 & ~x90 & ~x91 & ~x92 & ~x93 & ~x96 & ~x97 & ~x108 & ~x114 & ~x117 & ~x121 & ~x122 & ~x126 & ~x136 & ~x138 & ~x141 & ~x142 & ~x143 & ~x144 & ~x146 & ~x160 & ~x166 & ~x168 & ~x170 & ~x172 & ~x175 & ~x188 & ~x193 & ~x194 & ~x195 & ~x198 & ~x200 & ~x202 & ~x203 & ~x221 & ~x226 & ~x228 & ~x230 & ~x231 & ~x232 & ~x243 & ~x258 & ~x276 & ~x277 & ~x282 & ~x286 & ~x305 & ~x307 & ~x310 & ~x312 & ~x313 & ~x314 & ~x332 & ~x333 & ~x334 & ~x337 & ~x338 & ~x340 & ~x342 & ~x358 & ~x360 & ~x361 & ~x362 & ~x366 & ~x367 & ~x369 & ~x388 & ~x393 & ~x394 & ~x397 & ~x417 & ~x419 & ~x422 & ~x424 & ~x447 & ~x448 & ~x449 & ~x450 & ~x473 & ~x476 & ~x479 & ~x500 & ~x501 & ~x502 & ~x528 & ~x530 & ~x533 & ~x534 & ~x536 & ~x554 & ~x556 & ~x557 & ~x560 & ~x561 & ~x563 & ~x578 & ~x581 & ~x589 & ~x590 & ~x591 & ~x594 & ~x595 & ~x597 & ~x607 & ~x609 & ~x610 & ~x615 & ~x616 & ~x617 & ~x618 & ~x619 & ~x625 & ~x635 & ~x636 & ~x637 & ~x639 & ~x640 & ~x644 & ~x647 & ~x648 & ~x649 & ~x650 & ~x651 & ~x665 & ~x666 & ~x670 & ~x673 & ~x674 & ~x675 & ~x676 & ~x678 & ~x679 & ~x690 & ~x692 & ~x693 & ~x694 & ~x696 & ~x701 & ~x702 & ~x707 & ~x710 & ~x711 & ~x715 & ~x719 & ~x726 & ~x727 & ~x728 & ~x733 & ~x736 & ~x739 & ~x741 & ~x742 & ~x743 & ~x745 & ~x746 & ~x750 & ~x755 & ~x758 & ~x760 & ~x763 & ~x765 & ~x767 & ~x769 & ~x771 & ~x773 & ~x775 & ~x776 & ~x781 & ~x782;
assign c454 = ~x3 & ~x4 & ~x14 & ~x17 & ~x19 & ~x40 & ~x62 & ~x72 & ~x91 & ~x94 & ~x97 & ~x98 & ~x101 & ~x117 & ~x124 & ~x125 & ~x126 & ~x153 & ~x168 & ~x181 & ~x194 & ~x195 & ~x236 & ~x253 & ~x264 & ~x265 & ~x292 & ~x304 & ~x319 & ~x332 & ~x336 & ~x365 & ~x475 & ~x480 & ~x573 & ~x590 & ~x593 & ~x599 & ~x624 & ~x653 & ~x654 & ~x681 & ~x708 & ~x733 & ~x740 & ~x744 & ~x769 & ~x770;
assign c456 =  x426 &  x428 &  x438 &  x455 &  x456 & ~x19 & ~x20 & ~x21 & ~x24 & ~x34 & ~x42 & ~x80 & ~x81 & ~x95 & ~x137 & ~x144 & ~x221 & ~x225 & ~x281 & ~x309 & ~x368 & ~x588 & ~x589 & ~x592 & ~x597 & ~x624 & ~x625 & ~x642 & ~x644 & ~x651 & ~x680 & ~x681 & ~x710 & ~x715 & ~x719 & ~x722 & ~x730 & ~x741 & ~x742 & ~x747 & ~x748 & ~x755 & ~x768 & ~x776;
assign c458 =  x325 &  x380 &  x402 &  x430 &  x462 &  x463 & ~x1 & ~x3 & ~x6 & ~x7 & ~x9 & ~x11 & ~x12 & ~x14 & ~x15 & ~x17 & ~x19 & ~x23 & ~x24 & ~x26 & ~x30 & ~x32 & ~x38 & ~x43 & ~x45 & ~x50 & ~x54 & ~x57 & ~x63 & ~x64 & ~x65 & ~x66 & ~x70 & ~x72 & ~x74 & ~x78 & ~x84 & ~x85 & ~x88 & ~x89 & ~x90 & ~x94 & ~x96 & ~x98 & ~x106 & ~x107 & ~x109 & ~x111 & ~x114 & ~x129 & ~x135 & ~x139 & ~x140 & ~x141 & ~x143 & ~x146 & ~x147 & ~x148 & ~x163 & ~x164 & ~x166 & ~x168 & ~x170 & ~x174 & ~x175 & ~x177 & ~x190 & ~x192 & ~x194 & ~x197 & ~x198 & ~x200 & ~x203 & ~x221 & ~x223 & ~x226 & ~x227 & ~x228 & ~x230 & ~x232 & ~x246 & ~x252 & ~x255 & ~x256 & ~x257 & ~x259 & ~x273 & ~x276 & ~x280 & ~x282 & ~x285 & ~x286 & ~x301 & ~x302 & ~x303 & ~x306 & ~x308 & ~x311 & ~x313 & ~x328 & ~x329 & ~x332 & ~x336 & ~x360 & ~x364 & ~x365 & ~x366 & ~x368 & ~x392 & ~x394 & ~x395 & ~x396 & ~x419 & ~x445 & ~x450 & ~x451 & ~x472 & ~x473 & ~x474 & ~x499 & ~x503 & ~x507 & ~x527 & ~x529 & ~x532 & ~x534 & ~x537 & ~x553 & ~x558 & ~x559 & ~x562 & ~x564 & ~x565 & ~x580 & ~x581 & ~x585 & ~x589 & ~x590 & ~x591 & ~x592 & ~x595 & ~x610 & ~x612 & ~x616 & ~x620 & ~x637 & ~x639 & ~x640 & ~x641 & ~x647 & ~x649 & ~x665 & ~x666 & ~x667 & ~x668 & ~x669 & ~x672 & ~x675 & ~x679 & ~x691 & ~x692 & ~x694 & ~x700 & ~x702 & ~x703 & ~x704 & ~x706 & ~x707 & ~x708 & ~x709 & ~x714 & ~x715 & ~x720 & ~x722 & ~x723 & ~x724 & ~x725 & ~x726 & ~x727 & ~x729 & ~x734 & ~x736 & ~x737 & ~x738 & ~x741 & ~x749 & ~x750 & ~x757 & ~x758 & ~x761 & ~x762 & ~x763 & ~x767 & ~x770 & ~x771 & ~x772 & ~x774 & ~x776 & ~x778 & ~x779 & ~x780 & ~x781 & ~x782 & ~x783;
assign c460 = ~x22 & ~x54 & ~x84 & ~x85 & ~x89 & ~x94 & ~x95 & ~x123 & ~x127 & ~x129 & ~x207 & ~x213 & ~x233 & ~x241 & ~x250 & ~x252 & ~x254 & ~x268 & ~x283 & ~x295 & ~x323 & ~x363 & ~x392 & ~x443 & ~x445 & ~x479 & ~x577 & ~x583 & ~x634 & ~x675 & ~x700 & ~x719 & ~x731 & ~x733;
assign c462 =  x295 &  x323 &  x379 &  x380 &  x462 & ~x3 & ~x14 & ~x36 & ~x39 & ~x40 & ~x53 & ~x55 & ~x58 & ~x63 & ~x70 & ~x89 & ~x95 & ~x119 & ~x121 & ~x124 & ~x127 & ~x145 & ~x146 & ~x170 & ~x195 & ~x198 & ~x223 & ~x248 & ~x256 & ~x265 & ~x279 & ~x285 & ~x312 & ~x335 & ~x339 & ~x340 & ~x364 & ~x448 & ~x501 & ~x504 & ~x524 & ~x528 & ~x535 & ~x542 & ~x550 & ~x553 & ~x580 & ~x584 & ~x594 & ~x609 & ~x671 & ~x677 & ~x696 & ~x701 & ~x718 & ~x719 & ~x725 & ~x728 & ~x740 & ~x762 & ~x768 & ~x774;
assign c464 =  x492 & ~x1 & ~x2 & ~x3 & ~x6 & ~x7 & ~x8 & ~x11 & ~x12 & ~x17 & ~x18 & ~x21 & ~x22 & ~x23 & ~x24 & ~x25 & ~x26 & ~x27 & ~x30 & ~x31 & ~x34 & ~x36 & ~x40 & ~x44 & ~x45 & ~x47 & ~x49 & ~x51 & ~x53 & ~x54 & ~x57 & ~x66 & ~x67 & ~x68 & ~x72 & ~x76 & ~x77 & ~x81 & ~x84 & ~x87 & ~x89 & ~x90 & ~x92 & ~x94 & ~x95 & ~x104 & ~x106 & ~x109 & ~x110 & ~x111 & ~x114 & ~x115 & ~x117 & ~x118 & ~x119 & ~x121 & ~x125 & ~x126 & ~x131 & ~x135 & ~x136 & ~x137 & ~x138 & ~x142 & ~x146 & ~x149 & ~x160 & ~x162 & ~x165 & ~x166 & ~x167 & ~x168 & ~x169 & ~x170 & ~x174 & ~x175 & ~x177 & ~x190 & ~x192 & ~x193 & ~x198 & ~x200 & ~x201 & ~x205 & ~x217 & ~x219 & ~x220 & ~x222 & ~x225 & ~x227 & ~x228 & ~x232 & ~x244 & ~x248 & ~x251 & ~x252 & ~x253 & ~x254 & ~x256 & ~x257 & ~x258 & ~x259 & ~x272 & ~x275 & ~x277 & ~x278 & ~x279 & ~x282 & ~x287 & ~x302 & ~x305 & ~x314 & ~x332 & ~x333 & ~x338 & ~x340 & ~x341 & ~x357 & ~x358 & ~x359 & ~x360 & ~x361 & ~x363 & ~x365 & ~x368 & ~x386 & ~x389 & ~x391 & ~x394 & ~x396 & ~x417 & ~x420 & ~x421 & ~x422 & ~x424 & ~x446 & ~x447 & ~x449 & ~x450 & ~x451 & ~x452 & ~x473 & ~x475 & ~x476 & ~x501 & ~x504 & ~x505 & ~x508 & ~x529 & ~x530 & ~x532 & ~x533 & ~x536 & ~x556 & ~x558 & ~x565 & ~x567 & ~x584 & ~x590 & ~x591 & ~x592 & ~x594 & ~x595 & ~x597 & ~x599 & ~x608 & ~x609 & ~x611 & ~x612 & ~x613 & ~x618 & ~x619 & ~x621 & ~x622 & ~x626 & ~x635 & ~x637 & ~x638 & ~x639 & ~x648 & ~x650 & ~x652 & ~x654 & ~x655 & ~x665 & ~x666 & ~x668 & ~x669 & ~x670 & ~x673 & ~x675 & ~x676 & ~x677 & ~x678 & ~x679 & ~x681 & ~x698 & ~x701 & ~x703 & ~x704 & ~x705 & ~x708 & ~x709 & ~x712 & ~x714 & ~x716 & ~x717 & ~x720 & ~x721 & ~x722 & ~x723 & ~x724 & ~x725 & ~x729 & ~x730 & ~x731 & ~x732 & ~x733 & ~x740 & ~x741 & ~x745 & ~x746 & ~x747 & ~x749 & ~x752 & ~x754 & ~x755 & ~x756 & ~x763 & ~x764 & ~x765 & ~x766 & ~x767 & ~x769 & ~x770 & ~x778 & ~x779 & ~x781 & ~x782 & ~x783;
assign c466 =  x765;
assign c468 = ~x7 & ~x39 & ~x47 & ~x51 & ~x64 & ~x65 & ~x74 & ~x82 & ~x101 & ~x108 & ~x126 & ~x127 & ~x130 & ~x143 & ~x157 & ~x185 & ~x186 & ~x201 & ~x223 & ~x240 & ~x242 & ~x251 & ~x268 & ~x270 & ~x284 & ~x296 & ~x297 & ~x323 & ~x324 & ~x325 & ~x353 & ~x364 & ~x416 & ~x422 & ~x479 & ~x505 & ~x506 & ~x534 & ~x563 & ~x641 & ~x697 & ~x699 & ~x719 & ~x755;
assign c470 =  x355 &  x410 & ~x1 & ~x5 & ~x7 & ~x17 & ~x19 & ~x25 & ~x31 & ~x35 & ~x37 & ~x40 & ~x47 & ~x54 & ~x70 & ~x72 & ~x76 & ~x78 & ~x85 & ~x94 & ~x102 & ~x103 & ~x120 & ~x124 & ~x126 & ~x133 & ~x142 & ~x143 & ~x144 & ~x146 & ~x156 & ~x158 & ~x159 & ~x167 & ~x170 & ~x175 & ~x187 & ~x196 & ~x198 & ~x199 & ~x214 & ~x226 & ~x227 & ~x241 & ~x253 & ~x268 & ~x296 & ~x306 & ~x308 & ~x336 & ~x338 & ~x360 & ~x361 & ~x362 & ~x363 & ~x417 & ~x421 & ~x445 & ~x447 & ~x451 & ~x474 & ~x503 & ~x506 & ~x528 & ~x532 & ~x533 & ~x559 & ~x565 & ~x585 & ~x606 & ~x608 & ~x613 & ~x620 & ~x641 & ~x644 & ~x649 & ~x689 & ~x692 & ~x699 & ~x703 & ~x718 & ~x727 & ~x730 & ~x736 & ~x741 & ~x746 & ~x748 & ~x749 & ~x752 & ~x758 & ~x759 & ~x773 & ~x780 & ~x782;
assign c472 =  x411 & ~x9 & ~x10 & ~x15 & ~x18 & ~x32 & ~x41 & ~x48 & ~x66 & ~x82 & ~x88 & ~x89 & ~x90 & ~x100 & ~x103 & ~x105 & ~x107 & ~x109 & ~x112 & ~x128 & ~x137 & ~x138 & ~x142 & ~x166 & ~x167 & ~x184 & ~x211 & ~x239 & ~x254 & ~x267 & ~x279 & ~x283 & ~x305 & ~x309 & ~x323 & ~x339 & ~x361 & ~x367 & ~x446 & ~x473 & ~x477 & ~x500 & ~x505 & ~x507 & ~x528 & ~x560 & ~x562 & ~x572 & ~x573 & ~x583 & ~x584 & ~x598 & ~x599 & ~x600 & ~x612 & ~x617 & ~x621 & ~x629 & ~x675 & ~x676 & ~x678 & ~x704 & ~x711 & ~x713 & ~x726 & ~x728 & ~x729 & ~x739 & ~x747 & ~x750 & ~x755 & ~x756 & ~x767 & ~x770 & ~x776 & ~x779;
assign c474 =  x456 &  x487 &  x489 &  x491 & ~x4 & ~x62 & ~x63 & ~x108 & ~x115 & ~x129 & ~x130 & ~x222 & ~x260 & ~x304 & ~x479 & ~x539 & ~x549 & ~x581 & ~x622 & ~x635 & ~x700 & ~x747 & ~x777;
assign c476 = ~x1 & ~x5 & ~x8 & ~x13 & ~x14 & ~x24 & ~x35 & ~x40 & ~x43 & ~x44 & ~x45 & ~x46 & ~x48 & ~x51 & ~x52 & ~x54 & ~x58 & ~x62 & ~x66 & ~x67 & ~x68 & ~x69 & ~x70 & ~x71 & ~x75 & ~x76 & ~x78 & ~x79 & ~x80 & ~x88 & ~x89 & ~x98 & ~x106 & ~x109 & ~x111 & ~x116 & ~x126 & ~x130 & ~x133 & ~x138 & ~x141 & ~x145 & ~x154 & ~x164 & ~x165 & ~x167 & ~x169 & ~x172 & ~x182 & ~x192 & ~x195 & ~x197 & ~x198 & ~x210 & ~x221 & ~x222 & ~x224 & ~x226 & ~x227 & ~x248 & ~x250 & ~x255 & ~x265 & ~x280 & ~x281 & ~x282 & ~x293 & ~x303 & ~x304 & ~x306 & ~x310 & ~x332 & ~x335 & ~x364 & ~x365 & ~x390 & ~x392 & ~x418 & ~x443 & ~x446 & ~x449 & ~x452 & ~x472 & ~x475 & ~x478 & ~x501 & ~x527 & ~x531 & ~x532 & ~x534 & ~x536 & ~x556 & ~x563 & ~x572 & ~x573 & ~x587 & ~x589 & ~x590 & ~x591 & ~x593 & ~x611 & ~x612 & ~x616 & ~x629 & ~x641 & ~x642 & ~x645 & ~x646 & ~x656 & ~x657 & ~x669 & ~x670 & ~x673 & ~x674 & ~x675 & ~x679 & ~x680 & ~x685 & ~x697 & ~x704 & ~x705 & ~x708 & ~x713 & ~x723 & ~x725 & ~x727 & ~x731 & ~x733 & ~x734 & ~x738 & ~x741 & ~x743 & ~x746 & ~x748 & ~x752 & ~x754 & ~x759 & ~x762 & ~x765 & ~x768 & ~x774 & ~x779 & ~x783;
assign c478 =  x375 &  x404 &  x409 &  x435 &  x463 & ~x12 & ~x14 & ~x17 & ~x33 & ~x41 & ~x47 & ~x49 & ~x56 & ~x59 & ~x63 & ~x69 & ~x80 & ~x85 & ~x88 & ~x116 & ~x120 & ~x121 & ~x138 & ~x143 & ~x145 & ~x151 & ~x158 & ~x159 & ~x186 & ~x197 & ~x201 & ~x207 & ~x284 & ~x305 & ~x306 & ~x310 & ~x336 & ~x341 & ~x368 & ~x393 & ~x394 & ~x418 & ~x420 & ~x445 & ~x478 & ~x479 & ~x504 & ~x552 & ~x558 & ~x566 & ~x569 & ~x580 & ~x588 & ~x596 & ~x611 & ~x621 & ~x622 & ~x624 & ~x636 & ~x638 & ~x639 & ~x642 & ~x651 & ~x673 & ~x677 & ~x680 & ~x693 & ~x701 & ~x706 & ~x707 & ~x710 & ~x713 & ~x722 & ~x727 & ~x734 & ~x764 & ~x767 & ~x775 & ~x779 & ~x780 & ~x781 & ~x783;
assign c480 =  x187 &  x215 &  x270 &  x298 &  x518 & ~x14 & ~x69 & ~x111 & ~x126 & ~x155 & ~x173 & ~x255 & ~x330 & ~x332 & ~x362 & ~x421 & ~x448 & ~x531 & ~x562 & ~x594 & ~x620 & ~x623 & ~x667 & ~x680 & ~x688 & ~x704 & ~x715 & ~x745 & ~x764 & ~x783;
assign c482 = ~x0 & ~x10 & ~x14 & ~x19 & ~x23 & ~x26 & ~x31 & ~x35 & ~x37 & ~x39 & ~x40 & ~x43 & ~x51 & ~x52 & ~x58 & ~x68 & ~x72 & ~x76 & ~x79 & ~x84 & ~x86 & ~x90 & ~x94 & ~x98 & ~x100 & ~x108 & ~x124 & ~x125 & ~x134 & ~x137 & ~x138 & ~x139 & ~x142 & ~x144 & ~x154 & ~x169 & ~x181 & ~x182 & ~x192 & ~x193 & ~x194 & ~x222 & ~x224 & ~x236 & ~x237 & ~x252 & ~x275 & ~x277 & ~x281 & ~x292 & ~x310 & ~x331 & ~x334 & ~x335 & ~x363 & ~x364 & ~x391 & ~x420 & ~x421 & ~x446 & ~x451 & ~x470 & ~x473 & ~x479 & ~x480 & ~x502 & ~x503 & ~x508 & ~x509 & ~x526 & ~x527 & ~x532 & ~x539 & ~x561 & ~x562 & ~x563 & ~x584 & ~x585 & ~x589 & ~x612 & ~x614 & ~x617 & ~x618 & ~x628 & ~x642 & ~x648 & ~x649 & ~x656 & ~x670 & ~x671 & ~x677 & ~x678 & ~x680 & ~x695 & ~x707 & ~x712 & ~x719 & ~x724 & ~x728 & ~x730 & ~x736 & ~x739 & ~x744 & ~x745 & ~x746 & ~x752 & ~x754 & ~x756 & ~x757 & ~x760 & ~x770 & ~x774;
assign c484 =  x374 &  x402 &  x406 & ~x3 & ~x5 & ~x6 & ~x8 & ~x16 & ~x17 & ~x18 & ~x20 & ~x23 & ~x25 & ~x26 & ~x28 & ~x30 & ~x31 & ~x34 & ~x40 & ~x43 & ~x44 & ~x45 & ~x47 & ~x49 & ~x53 & ~x57 & ~x59 & ~x69 & ~x72 & ~x77 & ~x82 & ~x83 & ~x90 & ~x93 & ~x94 & ~x96 & ~x97 & ~x98 & ~x100 & ~x101 & ~x104 & ~x106 & ~x118 & ~x119 & ~x121 & ~x127 & ~x129 & ~x137 & ~x138 & ~x140 & ~x147 & ~x148 & ~x149 & ~x155 & ~x167 & ~x169 & ~x171 & ~x172 & ~x176 & ~x195 & ~x196 & ~x201 & ~x211 & ~x224 & ~x225 & ~x226 & ~x228 & ~x253 & ~x254 & ~x255 & ~x276 & ~x280 & ~x283 & ~x304 & ~x305 & ~x306 & ~x307 & ~x311 & ~x332 & ~x335 & ~x362 & ~x365 & ~x366 & ~x390 & ~x420 & ~x422 & ~x423 & ~x424 & ~x444 & ~x447 & ~x450 & ~x471 & ~x475 & ~x476 & ~x477 & ~x498 & ~x500 & ~x501 & ~x505 & ~x506 & ~x507 & ~x510 & ~x525 & ~x532 & ~x537 & ~x540 & ~x551 & ~x553 & ~x554 & ~x558 & ~x560 & ~x562 & ~x566 & ~x581 & ~x586 & ~x589 & ~x592 & ~x611 & ~x614 & ~x620 & ~x643 & ~x647 & ~x667 & ~x668 & ~x671 & ~x699 & ~x704 & ~x707 & ~x709 & ~x718 & ~x722 & ~x725 & ~x726 & ~x734 & ~x736 & ~x748 & ~x752 & ~x757 & ~x759 & ~x769 & ~x770 & ~x776 & ~x779;
assign c486 =  x291 &  x352 & ~x31 & ~x32 & ~x54 & ~x56 & ~x94 & ~x97 & ~x102 & ~x127 & ~x147 & ~x183 & ~x224 & ~x246 & ~x255 & ~x259 & ~x266 & ~x286 & ~x294 & ~x301 & ~x420 & ~x445 & ~x529 & ~x579 & ~x671 & ~x698 & ~x705 & ~x740 & ~x742;
assign c488 =  x295 &  x436 & ~x6 & ~x11 & ~x25 & ~x34 & ~x37 & ~x45 & ~x50 & ~x61 & ~x74 & ~x91 & ~x96 & ~x101 & ~x106 & ~x108 & ~x123 & ~x130 & ~x145 & ~x153 & ~x165 & ~x190 & ~x208 & ~x209 & ~x218 & ~x222 & ~x236 & ~x244 & ~x264 & ~x274 & ~x282 & ~x308 & ~x333 & ~x338 & ~x362 & ~x367 & ~x391 & ~x419 & ~x421 & ~x423 & ~x508 & ~x555 & ~x556 & ~x568 & ~x582 & ~x591 & ~x611 & ~x614 & ~x622 & ~x680 & ~x699 & ~x712 & ~x723 & ~x725 & ~x732 & ~x738 & ~x758 & ~x762 & ~x770 & ~x775 & ~x779;
assign c490 =  x483 & ~x18 & ~x31 & ~x35 & ~x69 & ~x82 & ~x92 & ~x95 & ~x116 & ~x128 & ~x213 & ~x241 & ~x278 & ~x284 & ~x296 & ~x338 & ~x363 & ~x393 & ~x416 & ~x419 & ~x585 & ~x586 & ~x617 & ~x620 & ~x625 & ~x645 & ~x647 & ~x706 & ~x710 & ~x716 & ~x721 & ~x751 & ~x761 & ~x777;
assign c492 =  x196;
assign c494 =  x464 &  x466 &  x468 &  x491 & ~x5 & ~x14 & ~x44 & ~x50 & ~x52 & ~x59 & ~x60 & ~x64 & ~x65 & ~x67 & ~x74 & ~x75 & ~x93 & ~x95 & ~x100 & ~x104 & ~x105 & ~x196 & ~x252 & ~x283 & ~x284 & ~x329 & ~x336 & ~x357 & ~x366 & ~x389 & ~x392 & ~x444 & ~x445 & ~x554 & ~x555 & ~x558 & ~x588 & ~x591 & ~x596 & ~x617 & ~x622 & ~x697 & ~x723 & ~x725 & ~x735 & ~x741 & ~x744 & ~x748 & ~x752 & ~x764 & ~x777 & ~x783;
assign c496 =  x299 &  x354 &  x381 &  x409 & ~x1 & ~x5 & ~x6 & ~x15 & ~x17 & ~x24 & ~x29 & ~x30 & ~x40 & ~x47 & ~x48 & ~x50 & ~x55 & ~x67 & ~x74 & ~x79 & ~x82 & ~x83 & ~x88 & ~x93 & ~x96 & ~x98 & ~x101 & ~x103 & ~x115 & ~x119 & ~x127 & ~x142 & ~x143 & ~x146 & ~x167 & ~x170 & ~x185 & ~x193 & ~x203 & ~x224 & ~x229 & ~x231 & ~x240 & ~x250 & ~x251 & ~x252 & ~x257 & ~x283 & ~x303 & ~x304 & ~x307 & ~x311 & ~x334 & ~x340 & ~x363 & ~x390 & ~x391 & ~x416 & ~x449 & ~x474 & ~x502 & ~x529 & ~x559 & ~x564 & ~x585 & ~x593 & ~x594 & ~x595 & ~x619 & ~x622 & ~x668 & ~x670 & ~x677 & ~x679 & ~x680 & ~x698 & ~x701 & ~x705 & ~x707 & ~x708 & ~x717 & ~x720 & ~x728 & ~x729 & ~x731 & ~x732 & ~x733 & ~x735 & ~x737 & ~x738 & ~x740 & ~x748 & ~x752 & ~x759 & ~x763 & ~x767 & ~x769;
assign c498 =  x50;
assign c4100 =  x373 &  x438 & ~x1 & ~x6 & ~x13 & ~x18 & ~x24 & ~x26 & ~x39 & ~x41 & ~x53 & ~x56 & ~x61 & ~x62 & ~x67 & ~x98 & ~x99 & ~x108 & ~x119 & ~x127 & ~x141 & ~x165 & ~x195 & ~x196 & ~x211 & ~x238 & ~x251 & ~x254 & ~x330 & ~x361 & ~x363 & ~x366 & ~x389 & ~x390 & ~x417 & ~x422 & ~x448 & ~x449 & ~x474 & ~x504 & ~x553 & ~x564 & ~x582 & ~x586 & ~x587 & ~x589 & ~x590 & ~x596 & ~x609 & ~x672 & ~x679 & ~x698 & ~x699 & ~x700 & ~x716 & ~x728 & ~x735 & ~x738 & ~x739 & ~x742 & ~x750 & ~x757 & ~x765 & ~x775 & ~x780 & ~x781 & ~x782;
assign c4102 = ~x2 & ~x5 & ~x14 & ~x18 & ~x19 & ~x22 & ~x26 & ~x37 & ~x44 & ~x45 & ~x49 & ~x56 & ~x65 & ~x68 & ~x70 & ~x85 & ~x92 & ~x93 & ~x94 & ~x97 & ~x101 & ~x102 & ~x108 & ~x110 & ~x114 & ~x115 & ~x137 & ~x143 & ~x145 & ~x155 & ~x165 & ~x166 & ~x169 & ~x172 & ~x173 & ~x183 & ~x200 & ~x210 & ~x218 & ~x220 & ~x239 & ~x248 & ~x249 & ~x250 & ~x251 & ~x253 & ~x255 & ~x258 & ~x266 & ~x275 & ~x276 & ~x282 & ~x286 & ~x301 & ~x305 & ~x321 & ~x322 & ~x329 & ~x330 & ~x331 & ~x332 & ~x336 & ~x339 & ~x387 & ~x390 & ~x421 & ~x449 & ~x475 & ~x477 & ~x479 & ~x504 & ~x532 & ~x533 & ~x534 & ~x555 & ~x557 & ~x559 & ~x560 & ~x561 & ~x562 & ~x583 & ~x587 & ~x589 & ~x609 & ~x610 & ~x615 & ~x617 & ~x620 & ~x625 & ~x647 & ~x648 & ~x649 & ~x653 & ~x668 & ~x670 & ~x673 & ~x675 & ~x698 & ~x702 & ~x709 & ~x711 & ~x722 & ~x733 & ~x734 & ~x738 & ~x744 & ~x746 & ~x751 & ~x754 & ~x757 & ~x761 & ~x764 & ~x767 & ~x768 & ~x773 & ~x777;
assign c4104 = ~x25 & ~x35 & ~x49 & ~x57 & ~x58 & ~x80 & ~x104 & ~x151 & ~x195 & ~x197 & ~x208 & ~x253 & ~x255 & ~x264 & ~x320 & ~x360 & ~x365 & ~x393 & ~x445 & ~x542 & ~x544 & ~x560 & ~x570 & ~x584 & ~x585 & ~x624 & ~x642 & ~x653 & ~x654 & ~x655 & ~x714 & ~x728 & ~x737 & ~x749 & ~x767 & ~x781 & ~x783;
assign c4106 =  x431 & ~x12 & ~x18 & ~x23 & ~x27 & ~x29 & ~x45 & ~x46 & ~x49 & ~x63 & ~x73 & ~x81 & ~x89 & ~x101 & ~x102 & ~x106 & ~x117 & ~x123 & ~x130 & ~x136 & ~x137 & ~x139 & ~x143 & ~x188 & ~x205 & ~x206 & ~x222 & ~x234 & ~x254 & ~x280 & ~x308 & ~x334 & ~x362 & ~x367 & ~x388 & ~x393 & ~x394 & ~x420 & ~x475 & ~x478 & ~x510 & ~x526 & ~x534 & ~x535 & ~x558 & ~x564 & ~x565 & ~x566 & ~x574 & ~x589 & ~x611 & ~x613 & ~x619 & ~x630 & ~x643 & ~x646 & ~x647 & ~x657 & ~x667 & ~x670 & ~x671 & ~x672 & ~x685 & ~x686 & ~x687 & ~x688 & ~x698 & ~x702 & ~x712 & ~x716 & ~x737 & ~x739 & ~x740 & ~x746 & ~x753 & ~x755 & ~x763 & ~x776 & ~x781 & ~x782;
assign c4108 = ~x15 & ~x24 & ~x30 & ~x39 & ~x64 & ~x68 & ~x69 & ~x78 & ~x95 & ~x101 & ~x141 & ~x143 & ~x156 & ~x183 & ~x194 & ~x199 & ~x202 & ~x211 & ~x248 & ~x249 & ~x251 & ~x255 & ~x258 & ~x266 & ~x277 & ~x285 & ~x314 & ~x321 & ~x330 & ~x361 & ~x365 & ~x417 & ~x505 & ~x510 & ~x544 & ~x551 & ~x580 & ~x593 & ~x598 & ~x653 & ~x668 & ~x705 & ~x736 & ~x744 & ~x747 & ~x754 & ~x772 & ~x781;
assign c4110 =  x401 &  x402 & ~x2 & ~x7 & ~x17 & ~x43 & ~x63 & ~x65 & ~x76 & ~x78 & ~x84 & ~x85 & ~x88 & ~x94 & ~x99 & ~x110 & ~x124 & ~x131 & ~x134 & ~x149 & ~x158 & ~x161 & ~x162 & ~x178 & ~x223 & ~x241 & ~x243 & ~x255 & ~x269 & ~x270 & ~x284 & ~x285 & ~x297 & ~x333 & ~x335 & ~x386 & ~x392 & ~x420 & ~x424 & ~x445 & ~x472 & ~x476 & ~x478 & ~x497 & ~x531 & ~x558 & ~x560 & ~x565 & ~x579 & ~x585 & ~x591 & ~x641 & ~x643 & ~x664 & ~x702 & ~x703 & ~x717 & ~x724 & ~x733 & ~x750 & ~x751 & ~x760 & ~x767 & ~x770 & ~x772 & ~x778;
assign c4112 =  x214 &  x325 &  x374 & ~x11 & ~x31 & ~x34 & ~x55 & ~x69 & ~x71 & ~x82 & ~x83 & ~x85 & ~x87 & ~x121 & ~x141 & ~x145 & ~x146 & ~x163 & ~x171 & ~x174 & ~x191 & ~x194 & ~x198 & ~x228 & ~x231 & ~x251 & ~x275 & ~x277 & ~x280 & ~x282 & ~x284 & ~x300 & ~x301 & ~x307 & ~x308 & ~x311 & ~x314 & ~x337 & ~x356 & ~x364 & ~x394 & ~x396 & ~x450 & ~x474 & ~x528 & ~x553 & ~x555 & ~x558 & ~x563 & ~x582 & ~x588 & ~x616 & ~x622 & ~x672 & ~x681 & ~x683 & ~x684 & ~x705 & ~x713 & ~x720 & ~x723 & ~x726 & ~x763;
assign c4114 =  x534;
assign c4116 =  x463 &  x489 &  x490 &  x517 &  x544 &  x600 &  x627 & ~x3 & ~x4 & ~x5 & ~x7 & ~x10 & ~x11 & ~x12 & ~x13 & ~x15 & ~x17 & ~x21 & ~x53 & ~x57 & ~x58 & ~x61 & ~x64 & ~x66 & ~x67 & ~x68 & ~x72 & ~x74 & ~x76 & ~x77 & ~x78 & ~x84 & ~x86 & ~x92 & ~x95 & ~x96 & ~x97 & ~x99 & ~x100 & ~x107 & ~x112 & ~x114 & ~x115 & ~x118 & ~x119 & ~x120 & ~x126 & ~x127 & ~x134 & ~x135 & ~x136 & ~x137 & ~x138 & ~x139 & ~x140 & ~x141 & ~x147 & ~x148 & ~x167 & ~x170 & ~x171 & ~x175 & ~x177 & ~x195 & ~x198 & ~x200 & ~x203 & ~x223 & ~x224 & ~x225 & ~x226 & ~x227 & ~x229 & ~x232 & ~x254 & ~x255 & ~x256 & ~x259 & ~x280 & ~x282 & ~x284 & ~x310 & ~x335 & ~x338 & ~x341 & ~x365 & ~x366 & ~x369 & ~x392 & ~x393 & ~x424 & ~x444 & ~x445 & ~x446 & ~x450 & ~x451 & ~x452 & ~x471 & ~x473 & ~x478 & ~x500 & ~x502 & ~x503 & ~x504 & ~x507 & ~x508 & ~x527 & ~x528 & ~x530 & ~x532 & ~x537 & ~x540 & ~x541 & ~x542 & ~x554 & ~x556 & ~x559 & ~x561 & ~x562 & ~x563 & ~x564 & ~x566 & ~x568 & ~x569 & ~x576 & ~x581 & ~x584 & ~x586 & ~x587 & ~x592 & ~x593 & ~x594 & ~x604 & ~x607 & ~x611 & ~x613 & ~x614 & ~x616 & ~x617 & ~x618 & ~x619 & ~x621 & ~x624 & ~x632 & ~x636 & ~x638 & ~x640 & ~x642 & ~x644 & ~x660 & ~x661 & ~x663 & ~x673 & ~x674 & ~x675 & ~x676 & ~x689 & ~x691 & ~x695 & ~x696 & ~x697 & ~x699 & ~x700 & ~x701 & ~x703 & ~x704 & ~x705 & ~x708 & ~x713 & ~x717 & ~x721 & ~x723 & ~x724 & ~x725 & ~x727 & ~x729 & ~x732 & ~x738 & ~x740 & ~x742 & ~x743 & ~x747 & ~x748 & ~x750 & ~x752 & ~x756 & ~x759 & ~x760 & ~x768 & ~x773 & ~x774 & ~x778 & ~x781 & ~x782;
assign c4118 = ~x8 & ~x26 & ~x52 & ~x65 & ~x88 & ~x92 & ~x96 & ~x97 & ~x102 & ~x104 & ~x115 & ~x167 & ~x183 & ~x193 & ~x229 & ~x238 & ~x251 & ~x275 & ~x293 & ~x322 & ~x363 & ~x471 & ~x479 & ~x504 & ~x529 & ~x549 & ~x567 & ~x583 & ~x633 & ~x642 & ~x643 & ~x647 & ~x648 & ~x651 & ~x681 & ~x692 & ~x701 & ~x718 & ~x722;
assign c4120 =  x346 &  x463 &  x490 & ~x14 & ~x17 & ~x18 & ~x20 & ~x22 & ~x23 & ~x34 & ~x35 & ~x43 & ~x44 & ~x49 & ~x50 & ~x56 & ~x60 & ~x70 & ~x74 & ~x87 & ~x89 & ~x97 & ~x98 & ~x102 & ~x103 & ~x106 & ~x113 & ~x119 & ~x121 & ~x122 & ~x140 & ~x141 & ~x149 & ~x150 & ~x165 & ~x176 & ~x195 & ~x196 & ~x199 & ~x200 & ~x202 & ~x223 & ~x224 & ~x229 & ~x230 & ~x248 & ~x250 & ~x256 & ~x261 & ~x275 & ~x276 & ~x279 & ~x280 & ~x287 & ~x302 & ~x305 & ~x315 & ~x332 & ~x333 & ~x336 & ~x340 & ~x357 & ~x360 & ~x361 & ~x384 & ~x385 & ~x390 & ~x395 & ~x421 & ~x446 & ~x474 & ~x475 & ~x478 & ~x479 & ~x501 & ~x504 & ~x505 & ~x529 & ~x530 & ~x533 & ~x535 & ~x536 & ~x554 & ~x557 & ~x558 & ~x580 & ~x581 & ~x584 & ~x585 & ~x588 & ~x593 & ~x595 & ~x597 & ~x613 & ~x614 & ~x615 & ~x618 & ~x621 & ~x639 & ~x640 & ~x641 & ~x646 & ~x647 & ~x648 & ~x649 & ~x665 & ~x672 & ~x673 & ~x674 & ~x675 & ~x676 & ~x677 & ~x693 & ~x695 & ~x696 & ~x697 & ~x698 & ~x699 & ~x701 & ~x709 & ~x712 & ~x715 & ~x716 & ~x721 & ~x723 & ~x728 & ~x736 & ~x737 & ~x739 & ~x742 & ~x744 & ~x746 & ~x747 & ~x754 & ~x755 & ~x764 & ~x765 & ~x767 & ~x768 & ~x769 & ~x780;
assign c4122 = ~x14 & ~x15 & ~x17 & ~x25 & ~x29 & ~x30 & ~x31 & ~x33 & ~x34 & ~x40 & ~x47 & ~x48 & ~x52 & ~x54 & ~x60 & ~x62 & ~x64 & ~x66 & ~x67 & ~x71 & ~x72 & ~x74 & ~x75 & ~x76 & ~x77 & ~x79 & ~x80 & ~x91 & ~x94 & ~x98 & ~x100 & ~x108 & ~x111 & ~x112 & ~x113 & ~x120 & ~x126 & ~x140 & ~x141 & ~x144 & ~x145 & ~x146 & ~x147 & ~x148 & ~x154 & ~x163 & ~x170 & ~x172 & ~x181 & ~x182 & ~x196 & ~x199 & ~x209 & ~x220 & ~x223 & ~x224 & ~x225 & ~x230 & ~x237 & ~x245 & ~x251 & ~x252 & ~x253 & ~x257 & ~x265 & ~x272 & ~x274 & ~x277 & ~x279 & ~x283 & ~x301 & ~x303 & ~x310 & ~x311 & ~x333 & ~x335 & ~x388 & ~x391 & ~x392 & ~x397 & ~x417 & ~x418 & ~x419 & ~x422 & ~x441 & ~x499 & ~x507 & ~x525 & ~x527 & ~x528 & ~x533 & ~x534 & ~x555 & ~x557 & ~x558 & ~x560 & ~x564 & ~x581 & ~x585 & ~x587 & ~x589 & ~x591 & ~x593 & ~x627 & ~x647 & ~x651 & ~x669 & ~x670 & ~x672 & ~x681 & ~x682 & ~x694 & ~x698 & ~x706 & ~x708 & ~x710 & ~x724 & ~x725 & ~x731 & ~x732 & ~x735 & ~x736 & ~x740 & ~x745 & ~x747 & ~x748 & ~x750 & ~x753 & ~x755 & ~x760 & ~x768 & ~x770 & ~x772 & ~x777 & ~x780 & ~x782;
assign c4124 =  x346 &  x399 & ~x0 & ~x2 & ~x26 & ~x27 & ~x35 & ~x45 & ~x46 & ~x47 & ~x49 & ~x58 & ~x66 & ~x69 & ~x75 & ~x96 & ~x101 & ~x112 & ~x115 & ~x116 & ~x168 & ~x171 & ~x172 & ~x203 & ~x205 & ~x250 & ~x260 & ~x277 & ~x281 & ~x305 & ~x307 & ~x310 & ~x314 & ~x364 & ~x368 & ~x369 & ~x393 & ~x418 & ~x421 & ~x446 & ~x503 & ~x527 & ~x533 & ~x561 & ~x564 & ~x567 & ~x568 & ~x580 & ~x581 & ~x585 & ~x588 & ~x607 & ~x614 & ~x615 & ~x619 & ~x622 & ~x637 & ~x644 & ~x674 & ~x675 & ~x679 & ~x681 & ~x696 & ~x717 & ~x720 & ~x733 & ~x737 & ~x739 & ~x751 & ~x758 & ~x759 & ~x760 & ~x764 & ~x773 & ~x780 & ~x782;
assign c4126 =  x237 & ~x16 & ~x31 & ~x33 & ~x57 & ~x58 & ~x66 & ~x69 & ~x78 & ~x92 & ~x94 & ~x96 & ~x97 & ~x101 & ~x108 & ~x126 & ~x128 & ~x140 & ~x141 & ~x143 & ~x165 & ~x185 & ~x212 & ~x230 & ~x240 & ~x250 & ~x257 & ~x260 & ~x268 & ~x279 & ~x332 & ~x392 & ~x418 & ~x425 & ~x446 & ~x479 & ~x503 & ~x506 & ~x509 & ~x550 & ~x553 & ~x581 & ~x582 & ~x588 & ~x615 & ~x621 & ~x640 & ~x646 & ~x648 & ~x663 & ~x675 & ~x690 & ~x702 & ~x705 & ~x731 & ~x737 & ~x743 & ~x751 & ~x772 & ~x779;
assign c4128 =  x408 &  x409 & ~x27 & ~x37 & ~x67 & ~x93 & ~x104 & ~x112 & ~x113 & ~x122 & ~x138 & ~x140 & ~x151 & ~x152 & ~x180 & ~x219 & ~x235 & ~x236 & ~x253 & ~x277 & ~x291 & ~x309 & ~x310 & ~x366 & ~x497 & ~x513 & ~x536 & ~x537 & ~x539 & ~x671 & ~x680 & ~x703 & ~x766 & ~x781;
assign c4130 =  x427;
assign c4132 =  x465 & ~x12 & ~x26 & ~x33 & ~x38 & ~x49 & ~x68 & ~x69 & ~x82 & ~x83 & ~x86 & ~x88 & ~x90 & ~x95 & ~x97 & ~x99 & ~x102 & ~x121 & ~x123 & ~x128 & ~x129 & ~x132 & ~x137 & ~x138 & ~x141 & ~x147 & ~x148 & ~x173 & ~x192 & ~x193 & ~x194 & ~x195 & ~x219 & ~x220 & ~x253 & ~x277 & ~x285 & ~x303 & ~x307 & ~x308 & ~x309 & ~x339 & ~x362 & ~x365 & ~x366 & ~x368 & ~x396 & ~x418 & ~x446 & ~x447 & ~x453 & ~x477 & ~x478 & ~x480 & ~x505 & ~x508 & ~x532 & ~x534 & ~x539 & ~x555 & ~x556 & ~x560 & ~x566 & ~x577 & ~x581 & ~x583 & ~x606 & ~x613 & ~x619 & ~x620 & ~x623 & ~x636 & ~x646 & ~x648 & ~x652 & ~x665 & ~x666 & ~x667 & ~x672 & ~x673 & ~x690 & ~x691 & ~x695 & ~x698 & ~x701 & ~x702 & ~x704 & ~x709 & ~x710 & ~x711 & ~x713 & ~x716 & ~x722 & ~x729 & ~x733 & ~x740 & ~x741 & ~x742 & ~x744 & ~x746 & ~x750 & ~x751 & ~x757 & ~x761 & ~x765 & ~x768 & ~x774 & ~x776 & ~x778 & ~x780 & ~x782;
assign c4134 =  x292 &  x375 &  x492 & ~x2 & ~x6 & ~x8 & ~x13 & ~x19 & ~x20 & ~x23 & ~x30 & ~x31 & ~x44 & ~x45 & ~x46 & ~x48 & ~x49 & ~x53 & ~x59 & ~x61 & ~x76 & ~x81 & ~x85 & ~x98 & ~x101 & ~x106 & ~x109 & ~x112 & ~x114 & ~x118 & ~x123 & ~x127 & ~x135 & ~x140 & ~x142 & ~x146 & ~x150 & ~x161 & ~x162 & ~x175 & ~x176 & ~x178 & ~x193 & ~x195 & ~x202 & ~x203 & ~x221 & ~x225 & ~x227 & ~x230 & ~x234 & ~x252 & ~x256 & ~x258 & ~x260 & ~x277 & ~x283 & ~x285 & ~x288 & ~x309 & ~x311 & ~x313 & ~x328 & ~x333 & ~x334 & ~x335 & ~x339 & ~x365 & ~x389 & ~x391 & ~x393 & ~x396 & ~x416 & ~x420 & ~x421 & ~x451 & ~x479 & ~x507 & ~x508 & ~x530 & ~x531 & ~x532 & ~x534 & ~x537 & ~x556 & ~x557 & ~x561 & ~x570 & ~x571 & ~x584 & ~x585 & ~x586 & ~x589 & ~x593 & ~x610 & ~x613 & ~x616 & ~x622 & ~x626 & ~x650 & ~x651 & ~x652 & ~x654 & ~x670 & ~x674 & ~x679 & ~x692 & ~x695 & ~x696 & ~x705 & ~x706 & ~x709 & ~x710 & ~x712 & ~x714 & ~x720 & ~x723 & ~x728 & ~x729 & ~x739 & ~x742 & ~x748 & ~x754 & ~x756 & ~x757 & ~x759 & ~x773 & ~x780;
assign c4136 =  x588;
assign c4138 =  x485 &  x486 & ~x0 & ~x5 & ~x6 & ~x10 & ~x12 & ~x13 & ~x14 & ~x18 & ~x19 & ~x23 & ~x25 & ~x26 & ~x27 & ~x32 & ~x39 & ~x44 & ~x50 & ~x56 & ~x59 & ~x67 & ~x69 & ~x71 & ~x73 & ~x75 & ~x79 & ~x90 & ~x91 & ~x92 & ~x93 & ~x96 & ~x97 & ~x112 & ~x115 & ~x116 & ~x122 & ~x140 & ~x141 & ~x143 & ~x146 & ~x164 & ~x167 & ~x169 & ~x173 & ~x193 & ~x197 & ~x200 & ~x202 & ~x203 & ~x204 & ~x220 & ~x223 & ~x224 & ~x225 & ~x229 & ~x249 & ~x252 & ~x279 & ~x282 & ~x287 & ~x307 & ~x309 & ~x310 & ~x312 & ~x331 & ~x332 & ~x333 & ~x337 & ~x359 & ~x363 & ~x364 & ~x365 & ~x366 & ~x367 & ~x368 & ~x388 & ~x391 & ~x393 & ~x405 & ~x418 & ~x419 & ~x420 & ~x422 & ~x433 & ~x446 & ~x475 & ~x478 & ~x479 & ~x535 & ~x556 & ~x558 & ~x560 & ~x564 & ~x570 & ~x571 & ~x583 & ~x584 & ~x585 & ~x587 & ~x588 & ~x590 & ~x591 & ~x592 & ~x593 & ~x594 & ~x595 & ~x610 & ~x615 & ~x616 & ~x617 & ~x622 & ~x625 & ~x626 & ~x644 & ~x646 & ~x647 & ~x648 & ~x650 & ~x651 & ~x653 & ~x666 & ~x667 & ~x668 & ~x670 & ~x671 & ~x673 & ~x675 & ~x676 & ~x677 & ~x684 & ~x694 & ~x695 & ~x696 & ~x698 & ~x699 & ~x700 & ~x703 & ~x711 & ~x713 & ~x714 & ~x717 & ~x718 & ~x721 & ~x725 & ~x726 & ~x728 & ~x729 & ~x731 & ~x733 & ~x734 & ~x740 & ~x750 & ~x751 & ~x752 & ~x755 & ~x761 & ~x763 & ~x764 & ~x765 & ~x766 & ~x769 & ~x771 & ~x773 & ~x774 & ~x777 & ~x778 & ~x780 & ~x781;
assign c4140 =  x14;
assign c4142 =  x409 &  x430 & ~x3 & ~x10 & ~x15 & ~x16 & ~x30 & ~x41 & ~x65 & ~x70 & ~x83 & ~x85 & ~x96 & ~x97 & ~x98 & ~x100 & ~x106 & ~x112 & ~x114 & ~x126 & ~x128 & ~x129 & ~x132 & ~x133 & ~x136 & ~x156 & ~x168 & ~x171 & ~x172 & ~x184 & ~x199 & ~x212 & ~x239 & ~x267 & ~x281 & ~x310 & ~x333 & ~x361 & ~x367 & ~x390 & ~x473 & ~x478 & ~x498 & ~x503 & ~x507 & ~x525 & ~x529 & ~x533 & ~x556 & ~x562 & ~x592 & ~x593 & ~x594 & ~x639 & ~x641 & ~x642 & ~x643 & ~x672 & ~x673 & ~x699 & ~x709 & ~x720 & ~x733 & ~x743 & ~x746 & ~x750 & ~x756 & ~x758 & ~x759 & ~x764 & ~x765 & ~x777;
assign c4144 =  x643;
assign c4146 =  x408 &  x518 & ~x5 & ~x7 & ~x22 & ~x28 & ~x30 & ~x34 & ~x37 & ~x68 & ~x71 & ~x78 & ~x95 & ~x97 & ~x100 & ~x102 & ~x104 & ~x115 & ~x122 & ~x126 & ~x127 & ~x141 & ~x145 & ~x148 & ~x149 & ~x166 & ~x171 & ~x183 & ~x194 & ~x197 & ~x200 & ~x228 & ~x231 & ~x249 & ~x250 & ~x253 & ~x278 & ~x294 & ~x312 & ~x334 & ~x367 & ~x388 & ~x389 & ~x391 & ~x446 & ~x449 & ~x451 & ~x473 & ~x501 & ~x506 & ~x508 & ~x529 & ~x534 & ~x536 & ~x561 & ~x563 & ~x585 & ~x586 & ~x588 & ~x589 & ~x591 & ~x597 & ~x616 & ~x619 & ~x622 & ~x636 & ~x643 & ~x652 & ~x665 & ~x670 & ~x679 & ~x680 & ~x695 & ~x704 & ~x706 & ~x717 & ~x723 & ~x733 & ~x753 & ~x762 & ~x763 & ~x766 & ~x770 & ~x771;
assign c4148 =  x353 &  x435 & ~x18 & ~x21 & ~x32 & ~x37 & ~x39 & ~x52 & ~x56 & ~x67 & ~x69 & ~x80 & ~x125 & ~x127 & ~x141 & ~x148 & ~x166 & ~x169 & ~x185 & ~x198 & ~x200 & ~x240 & ~x258 & ~x259 & ~x267 & ~x277 & ~x286 & ~x310 & ~x311 & ~x322 & ~x364 & ~x369 & ~x391 & ~x425 & ~x452 & ~x475 & ~x480 & ~x505 & ~x532 & ~x536 & ~x540 & ~x552 & ~x565 & ~x567 & ~x583 & ~x612 & ~x614 & ~x621 & ~x634 & ~x640 & ~x646 & ~x665 & ~x672 & ~x699 & ~x716 & ~x717 & ~x737 & ~x743 & ~x747 & ~x757 & ~x774 & ~x775 & ~x777;
assign c4150 =  x464 & ~x0 & ~x2 & ~x5 & ~x6 & ~x14 & ~x17 & ~x24 & ~x25 & ~x26 & ~x27 & ~x33 & ~x34 & ~x38 & ~x41 & ~x49 & ~x61 & ~x63 & ~x64 & ~x67 & ~x75 & ~x77 & ~x78 & ~x86 & ~x87 & ~x96 & ~x97 & ~x102 & ~x103 & ~x104 & ~x105 & ~x114 & ~x122 & ~x129 & ~x133 & ~x140 & ~x141 & ~x145 & ~x148 & ~x166 & ~x167 & ~x170 & ~x172 & ~x178 & ~x188 & ~x194 & ~x195 & ~x199 & ~x207 & ~x223 & ~x224 & ~x251 & ~x253 & ~x277 & ~x279 & ~x282 & ~x283 & ~x284 & ~x306 & ~x333 & ~x337 & ~x339 & ~x357 & ~x359 & ~x363 & ~x393 & ~x417 & ~x422 & ~x423 & ~x447 & ~x448 & ~x449 & ~x450 & ~x453 & ~x478 & ~x480 & ~x502 & ~x509 & ~x513 & ~x525 & ~x526 & ~x528 & ~x531 & ~x532 & ~x537 & ~x540 & ~x556 & ~x557 & ~x567 & ~x573 & ~x583 & ~x588 & ~x591 & ~x593 & ~x600 & ~x602 & ~x613 & ~x619 & ~x621 & ~x627 & ~x629 & ~x639 & ~x640 & ~x641 & ~x643 & ~x644 & ~x658 & ~x669 & ~x674 & ~x675 & ~x683 & ~x684 & ~x697 & ~x706 & ~x707 & ~x711 & ~x714 & ~x724 & ~x730 & ~x731 & ~x737 & ~x744 & ~x746 & ~x747 & ~x750 & ~x753 & ~x754 & ~x759 & ~x763 & ~x765 & ~x766 & ~x768 & ~x771 & ~x773 & ~x774 & ~x781 & ~x783;
assign c4152 = ~x0 & ~x2 & ~x7 & ~x8 & ~x11 & ~x13 & ~x17 & ~x18 & ~x19 & ~x23 & ~x28 & ~x31 & ~x32 & ~x38 & ~x42 & ~x44 & ~x46 & ~x49 & ~x51 & ~x52 & ~x57 & ~x58 & ~x59 & ~x62 & ~x63 & ~x65 & ~x68 & ~x69 & ~x73 & ~x78 & ~x82 & ~x83 & ~x85 & ~x86 & ~x90 & ~x99 & ~x101 & ~x106 & ~x111 & ~x112 & ~x118 & ~x119 & ~x120 & ~x124 & ~x126 & ~x127 & ~x140 & ~x143 & ~x144 & ~x146 & ~x147 & ~x151 & ~x152 & ~x153 & ~x155 & ~x175 & ~x183 & ~x192 & ~x194 & ~x195 & ~x202 & ~x221 & ~x229 & ~x239 & ~x248 & ~x256 & ~x258 & ~x259 & ~x267 & ~x284 & ~x294 & ~x301 & ~x305 & ~x306 & ~x308 & ~x310 & ~x329 & ~x331 & ~x334 & ~x336 & ~x363 & ~x364 & ~x365 & ~x367 & ~x390 & ~x391 & ~x393 & ~x396 & ~x419 & ~x423 & ~x448 & ~x450 & ~x452 & ~x472 & ~x477 & ~x480 & ~x498 & ~x502 & ~x503 & ~x535 & ~x556 & ~x561 & ~x562 & ~x563 & ~x565 & ~x567 & ~x579 & ~x584 & ~x588 & ~x593 & ~x594 & ~x609 & ~x613 & ~x616 & ~x620 & ~x637 & ~x639 & ~x663 & ~x667 & ~x696 & ~x697 & ~x698 & ~x699 & ~x700 & ~x704 & ~x706 & ~x707 & ~x708 & ~x722 & ~x724 & ~x735 & ~x738 & ~x740 & ~x743 & ~x744 & ~x745 & ~x746 & ~x752 & ~x753 & ~x758 & ~x759 & ~x765 & ~x769 & ~x776 & ~x780 & ~x783;
assign c4154 =  x437 &  x466 & ~x12 & ~x36 & ~x58 & ~x73 & ~x89 & ~x91 & ~x98 & ~x134 & ~x154 & ~x182 & ~x210 & ~x266 & ~x294 & ~x322 & ~x334 & ~x475 & ~x500 & ~x505 & ~x508 & ~x529 & ~x562 & ~x564 & ~x591 & ~x598 & ~x627 & ~x655 & ~x656 & ~x674 & ~x683 & ~x697 & ~x705 & ~x707 & ~x710 & ~x741 & ~x779;
assign c4156 =  x243 & ~x0 & ~x3 & ~x5 & ~x6 & ~x29 & ~x33 & ~x34 & ~x36 & ~x44 & ~x52 & ~x56 & ~x58 & ~x63 & ~x65 & ~x69 & ~x70 & ~x76 & ~x80 & ~x81 & ~x82 & ~x85 & ~x90 & ~x101 & ~x110 & ~x116 & ~x121 & ~x122 & ~x137 & ~x158 & ~x167 & ~x168 & ~x171 & ~x192 & ~x213 & ~x222 & ~x226 & ~x227 & ~x228 & ~x229 & ~x249 & ~x252 & ~x268 & ~x276 & ~x277 & ~x281 & ~x282 & ~x303 & ~x304 & ~x308 & ~x309 & ~x313 & ~x332 & ~x333 & ~x338 & ~x363 & ~x364 & ~x368 & ~x388 & ~x389 & ~x390 & ~x392 & ~x418 & ~x420 & ~x502 & ~x505 & ~x531 & ~x563 & ~x615 & ~x618 & ~x630 & ~x641 & ~x642 & ~x643 & ~x645 & ~x647 & ~x649 & ~x670 & ~x671 & ~x679 & ~x686 & ~x697 & ~x700 & ~x704 & ~x706 & ~x712 & ~x713 & ~x716 & ~x717 & ~x719 & ~x728 & ~x733 & ~x736 & ~x740 & ~x747 & ~x748 & ~x756 & ~x757 & ~x758 & ~x760 & ~x766 & ~x773 & ~x775 & ~x777 & ~x779 & ~x782;
assign c4158 =  x315 &  x371 & ~x92 & ~x121 & ~x180 & ~x224 & ~x236 & ~x292 & ~x741;
assign c4160 =  x764;
assign c4162 =  x436 & ~x35 & ~x60 & ~x71 & ~x86 & ~x89 & ~x96 & ~x100 & ~x122 & ~x128 & ~x132 & ~x134 & ~x141 & ~x148 & ~x160 & ~x185 & ~x212 & ~x231 & ~x240 & ~x249 & ~x267 & ~x282 & ~x312 & ~x322 & ~x362 & ~x365 & ~x442 & ~x473 & ~x501 & ~x503 & ~x514 & ~x551 & ~x596 & ~x607 & ~x636 & ~x654 & ~x673 & ~x677 & ~x681 & ~x700 & ~x722 & ~x753 & ~x756 & ~x761 & ~x772;
assign c4164 =  x33;
assign c4166 =  x454 &  x455 &  x467 &  x468 &  x469 &  x489 &  x492;
assign c4168 =  x379 &  x435 & ~x36 & ~x37 & ~x53 & ~x55 & ~x66 & ~x69 & ~x70 & ~x73 & ~x85 & ~x88 & ~x95 & ~x97 & ~x105 & ~x115 & ~x122 & ~x126 & ~x127 & ~x133 & ~x136 & ~x138 & ~x139 & ~x140 & ~x145 & ~x147 & ~x154 & ~x169 & ~x172 & ~x174 & ~x182 & ~x189 & ~x191 & ~x199 & ~x200 & ~x216 & ~x226 & ~x238 & ~x251 & ~x253 & ~x256 & ~x259 & ~x272 & ~x277 & ~x279 & ~x284 & ~x299 & ~x300 & ~x304 & ~x305 & ~x306 & ~x307 & ~x313 & ~x314 & ~x367 & ~x448 & ~x474 & ~x477 & ~x501 & ~x530 & ~x534 & ~x539 & ~x558 & ~x563 & ~x587 & ~x590 & ~x607 & ~x614 & ~x618 & ~x620 & ~x638 & ~x639 & ~x641 & ~x645 & ~x647 & ~x648 & ~x671 & ~x676 & ~x691 & ~x693 & ~x721 & ~x727 & ~x740 & ~x761 & ~x766 & ~x768 & ~x771 & ~x773 & ~x777;
assign c4170 =  x372 &  x373 &  x412 &  x426 & ~x573;
assign c4172 =  x381 &  x403 &  x408 &  x460 & ~x20 & ~x36 & ~x41 & ~x57 & ~x68 & ~x71 & ~x72 & ~x78 & ~x85 & ~x86 & ~x94 & ~x106 & ~x117 & ~x122 & ~x124 & ~x156 & ~x166 & ~x176 & ~x184 & ~x212 & ~x225 & ~x284 & ~x445 & ~x446 & ~x523 & ~x527 & ~x539 & ~x567 & ~x579 & ~x591 & ~x605 & ~x606 & ~x749 & ~x773 & ~x781;
assign c4174 = ~x6 & ~x8 & ~x14 & ~x16 & ~x17 & ~x19 & ~x22 & ~x23 & ~x30 & ~x34 & ~x41 & ~x42 & ~x44 & ~x45 & ~x49 & ~x54 & ~x63 & ~x64 & ~x69 & ~x70 & ~x71 & ~x80 & ~x87 & ~x92 & ~x95 & ~x96 & ~x97 & ~x99 & ~x102 & ~x114 & ~x116 & ~x129 & ~x137 & ~x139 & ~x148 & ~x157 & ~x159 & ~x167 & ~x169 & ~x174 & ~x176 & ~x185 & ~x197 & ~x198 & ~x201 & ~x231 & ~x232 & ~x241 & ~x253 & ~x279 & ~x283 & ~x284 & ~x287 & ~x295 & ~x305 & ~x309 & ~x323 & ~x339 & ~x341 & ~x390 & ~x395 & ~x415 & ~x445 & ~x474 & ~x476 & ~x530 & ~x557 & ~x559 & ~x583 & ~x591 & ~x593 & ~x594 & ~x612 & ~x617 & ~x631 & ~x638 & ~x642 & ~x673 & ~x686 & ~x690 & ~x693 & ~x694 & ~x700 & ~x702 & ~x719 & ~x727 & ~x733 & ~x734 & ~x736 & ~x743 & ~x746 & ~x764 & ~x768 & ~x769 & ~x774 & ~x775 & ~x777 & ~x778;
assign c4176 =  x271 & ~x0 & ~x8 & ~x11 & ~x23 & ~x30 & ~x33 & ~x42 & ~x63 & ~x75 & ~x77 & ~x94 & ~x108 & ~x113 & ~x116 & ~x121 & ~x130 & ~x145 & ~x149 & ~x157 & ~x169 & ~x185 & ~x241 & ~x251 & ~x296 & ~x304 & ~x323 & ~x333 & ~x334 & ~x350 & ~x359 & ~x368 & ~x389 & ~x392 & ~x394 & ~x395 & ~x396 & ~x419 & ~x424 & ~x444 & ~x477 & ~x532 & ~x533 & ~x593 & ~x617 & ~x618 & ~x668 & ~x701 & ~x705 & ~x720 & ~x726 & ~x741 & ~x774 & ~x776 & ~x782;
assign c4178 =  x291 &  x347 &  x435 &  x464 &  x491 & ~x2 & ~x7 & ~x12 & ~x15 & ~x17 & ~x19 & ~x22 & ~x23 & ~x31 & ~x35 & ~x36 & ~x42 & ~x46 & ~x47 & ~x50 & ~x51 & ~x67 & ~x69 & ~x73 & ~x76 & ~x77 & ~x79 & ~x89 & ~x93 & ~x95 & ~x108 & ~x109 & ~x115 & ~x122 & ~x132 & ~x139 & ~x161 & ~x162 & ~x166 & ~x168 & ~x175 & ~x187 & ~x193 & ~x194 & ~x230 & ~x232 & ~x243 & ~x254 & ~x282 & ~x284 & ~x286 & ~x307 & ~x312 & ~x338 & ~x341 & ~x390 & ~x396 & ~x421 & ~x446 & ~x448 & ~x451 & ~x479 & ~x532 & ~x533 & ~x535 & ~x541 & ~x542 & ~x559 & ~x561 & ~x566 & ~x579 & ~x585 & ~x592 & ~x593 & ~x595 & ~x596 & ~x610 & ~x622 & ~x624 & ~x634 & ~x643 & ~x668 & ~x698 & ~x715 & ~x716 & ~x719 & ~x723 & ~x732 & ~x736 & ~x741 & ~x742 & ~x744 & ~x745 & ~x746 & ~x767 & ~x770 & ~x772 & ~x780 & ~x783;
assign c4180 =  x86;
assign c4182 = ~x4 & ~x10 & ~x12 & ~x13 & ~x15 & ~x16 & ~x20 & ~x24 & ~x25 & ~x28 & ~x29 & ~x31 & ~x34 & ~x37 & ~x40 & ~x42 & ~x43 & ~x44 & ~x58 & ~x61 & ~x63 & ~x64 & ~x70 & ~x71 & ~x72 & ~x74 & ~x75 & ~x83 & ~x87 & ~x88 & ~x89 & ~x90 & ~x92 & ~x93 & ~x94 & ~x95 & ~x96 & ~x101 & ~x105 & ~x107 & ~x115 & ~x116 & ~x117 & ~x118 & ~x121 & ~x122 & ~x123 & ~x125 & ~x126 & ~x128 & ~x129 & ~x130 & ~x131 & ~x141 & ~x146 & ~x148 & ~x152 & ~x156 & ~x164 & ~x166 & ~x167 & ~x170 & ~x174 & ~x175 & ~x176 & ~x177 & ~x178 & ~x184 & ~x185 & ~x194 & ~x198 & ~x199 & ~x212 & ~x222 & ~x223 & ~x226 & ~x227 & ~x228 & ~x230 & ~x231 & ~x232 & ~x240 & ~x255 & ~x277 & ~x278 & ~x303 & ~x304 & ~x307 & ~x309 & ~x310 & ~x311 & ~x312 & ~x313 & ~x314 & ~x315 & ~x334 & ~x339 & ~x360 & ~x362 & ~x388 & ~x389 & ~x390 & ~x392 & ~x395 & ~x416 & ~x417 & ~x420 & ~x422 & ~x423 & ~x425 & ~x441 & ~x443 & ~x444 & ~x445 & ~x446 & ~x448 & ~x451 & ~x470 & ~x476 & ~x480 & ~x498 & ~x505 & ~x508 & ~x510 & ~x532 & ~x534 & ~x537 & ~x538 & ~x541 & ~x552 & ~x554 & ~x555 & ~x557 & ~x558 & ~x561 & ~x562 & ~x583 & ~x588 & ~x589 & ~x592 & ~x594 & ~x596 & ~x607 & ~x611 & ~x612 & ~x613 & ~x614 & ~x615 & ~x621 & ~x638 & ~x642 & ~x649 & ~x652 & ~x666 & ~x668 & ~x670 & ~x673 & ~x674 & ~x676 & ~x677 & ~x678 & ~x694 & ~x698 & ~x703 & ~x704 & ~x706 & ~x708 & ~x718 & ~x720 & ~x721 & ~x722 & ~x723 & ~x727 & ~x729 & ~x730 & ~x733 & ~x735 & ~x740 & ~x741 & ~x742 & ~x745 & ~x746 & ~x747 & ~x751 & ~x754 & ~x755 & ~x756 & ~x760 & ~x763 & ~x764 & ~x766 & ~x768 & ~x769 & ~x770 & ~x771 & ~x772 & ~x773 & ~x775 & ~x776 & ~x779 & ~x780 & ~x783;
assign c4184 =  x243 &  x298 &  x465 & ~x1 & ~x7 & ~x12 & ~x25 & ~x28 & ~x32 & ~x34 & ~x44 & ~x55 & ~x59 & ~x66 & ~x67 & ~x68 & ~x85 & ~x86 & ~x87 & ~x91 & ~x95 & ~x97 & ~x99 & ~x100 & ~x101 & ~x109 & ~x112 & ~x116 & ~x127 & ~x128 & ~x141 & ~x156 & ~x166 & ~x184 & ~x196 & ~x198 & ~x200 & ~x239 & ~x251 & ~x253 & ~x267 & ~x277 & ~x303 & ~x338 & ~x450 & ~x478 & ~x504 & ~x507 & ~x532 & ~x533 & ~x534 & ~x555 & ~x559 & ~x586 & ~x591 & ~x593 & ~x612 & ~x621 & ~x643 & ~x646 & ~x647 & ~x669 & ~x673 & ~x674 & ~x723 & ~x725 & ~x729 & ~x730 & ~x732 & ~x734 & ~x736 & ~x739 & ~x741 & ~x742 & ~x743 & ~x745 & ~x749 & ~x751 & ~x768 & ~x771 & ~x778;
assign c4186 =  x403 &  x406 & ~x0 & ~x5 & ~x16 & ~x17 & ~x18 & ~x20 & ~x21 & ~x23 & ~x27 & ~x28 & ~x36 & ~x37 & ~x39 & ~x40 & ~x51 & ~x55 & ~x56 & ~x66 & ~x69 & ~x70 & ~x71 & ~x74 & ~x76 & ~x78 & ~x80 & ~x88 & ~x91 & ~x93 & ~x94 & ~x95 & ~x96 & ~x97 & ~x98 & ~x99 & ~x101 & ~x102 & ~x107 & ~x110 & ~x118 & ~x119 & ~x124 & ~x125 & ~x126 & ~x130 & ~x137 & ~x140 & ~x142 & ~x143 & ~x145 & ~x147 & ~x157 & ~x158 & ~x164 & ~x166 & ~x170 & ~x201 & ~x212 & ~x227 & ~x239 & ~x253 & ~x256 & ~x267 & ~x280 & ~x283 & ~x309 & ~x311 & ~x312 & ~x334 & ~x335 & ~x336 & ~x339 & ~x361 & ~x389 & ~x393 & ~x420 & ~x421 & ~x422 & ~x449 & ~x451 & ~x471 & ~x473 & ~x475 & ~x476 & ~x478 & ~x500 & ~x502 & ~x514 & ~x529 & ~x537 & ~x540 & ~x541 & ~x555 & ~x561 & ~x563 & ~x566 & ~x568 & ~x584 & ~x586 & ~x588 & ~x589 & ~x592 & ~x606 & ~x619 & ~x633 & ~x640 & ~x643 & ~x648 & ~x650 & ~x661 & ~x663 & ~x664 & ~x667 & ~x669 & ~x672 & ~x689 & ~x690 & ~x696 & ~x699 & ~x700 & ~x701 & ~x704 & ~x715 & ~x723 & ~x728 & ~x730 & ~x732 & ~x734 & ~x735 & ~x738 & ~x747 & ~x748 & ~x751 & ~x754 & ~x756 & ~x762 & ~x766 & ~x768 & ~x769 & ~x771 & ~x781;
assign c4188 = ~x9 & ~x33 & ~x34 & ~x42 & ~x53 & ~x54 & ~x60 & ~x64 & ~x65 & ~x72 & ~x78 & ~x90 & ~x94 & ~x95 & ~x100 & ~x105 & ~x122 & ~x127 & ~x128 & ~x133 & ~x134 & ~x139 & ~x152 & ~x166 & ~x168 & ~x172 & ~x175 & ~x177 & ~x186 & ~x208 & ~x258 & ~x277 & ~x281 & ~x282 & ~x286 & ~x307 & ~x311 & ~x313 & ~x334 & ~x337 & ~x338 & ~x360 & ~x365 & ~x367 & ~x389 & ~x391 & ~x394 & ~x416 & ~x421 & ~x446 & ~x449 & ~x451 & ~x470 & ~x479 & ~x499 & ~x500 & ~x502 & ~x509 & ~x526 & ~x530 & ~x532 & ~x540 & ~x552 & ~x554 & ~x557 & ~x593 & ~x594 & ~x604 & ~x610 & ~x618 & ~x640 & ~x646 & ~x663 & ~x674 & ~x689 & ~x692 & ~x700 & ~x721 & ~x723 & ~x728 & ~x729 & ~x732 & ~x737 & ~x738 & ~x739 & ~x741 & ~x742 & ~x743 & ~x745 & ~x750 & ~x762 & ~x782 & ~x783;
assign c4190 = ~x3 & ~x7 & ~x11 & ~x15 & ~x19 & ~x23 & ~x33 & ~x35 & ~x36 & ~x43 & ~x45 & ~x56 & ~x65 & ~x66 & ~x69 & ~x70 & ~x73 & ~x77 & ~x80 & ~x81 & ~x85 & ~x88 & ~x90 & ~x92 & ~x93 & ~x94 & ~x111 & ~x115 & ~x117 & ~x125 & ~x127 & ~x133 & ~x136 & ~x143 & ~x149 & ~x150 & ~x151 & ~x157 & ~x169 & ~x176 & ~x177 & ~x199 & ~x213 & ~x224 & ~x226 & ~x232 & ~x240 & ~x252 & ~x256 & ~x257 & ~x268 & ~x284 & ~x308 & ~x310 & ~x332 & ~x334 & ~x336 & ~x339 & ~x361 & ~x363 & ~x364 & ~x389 & ~x391 & ~x397 & ~x417 & ~x418 & ~x419 & ~x472 & ~x474 & ~x477 & ~x479 & ~x498 & ~x505 & ~x536 & ~x560 & ~x561 & ~x562 & ~x565 & ~x568 & ~x580 & ~x586 & ~x588 & ~x595 & ~x605 & ~x606 & ~x607 & ~x614 & ~x633 & ~x635 & ~x646 & ~x673 & ~x675 & ~x676 & ~x678 & ~x679 & ~x700 & ~x720 & ~x722 & ~x732 & ~x734 & ~x738 & ~x754 & ~x759 & ~x760 & ~x771 & ~x775 & ~x779 & ~x780 & ~x783;
assign c4192 =  x240 & ~x14 & ~x32 & ~x47 & ~x52 & ~x59 & ~x67 & ~x69 & ~x79 & ~x83 & ~x84 & ~x88 & ~x142 & ~x152 & ~x162 & ~x175 & ~x202 & ~x219 & ~x236 & ~x246 & ~x247 & ~x332 & ~x448 & ~x501 & ~x502 & ~x534 & ~x536 & ~x540 & ~x545 & ~x570 & ~x642 & ~x643 & ~x647 & ~x651 & ~x652 & ~x711 & ~x718 & ~x720 & ~x733 & ~x735 & ~x751 & ~x752 & ~x765 & ~x767 & ~x771 & ~x774;
assign c4194 =  x115;
assign c4196 = ~x2 & ~x5 & ~x9 & ~x13 & ~x14 & ~x17 & ~x21 & ~x28 & ~x34 & ~x38 & ~x40 & ~x45 & ~x50 & ~x56 & ~x57 & ~x64 & ~x66 & ~x69 & ~x70 & ~x71 & ~x73 & ~x74 & ~x75 & ~x76 & ~x86 & ~x90 & ~x93 & ~x95 & ~x97 & ~x103 & ~x110 & ~x113 & ~x114 & ~x121 & ~x128 & ~x131 & ~x134 & ~x138 & ~x139 & ~x146 & ~x154 & ~x167 & ~x169 & ~x172 & ~x182 & ~x191 & ~x192 & ~x195 & ~x201 & ~x221 & ~x226 & ~x227 & ~x250 & ~x251 & ~x255 & ~x256 & ~x266 & ~x277 & ~x278 & ~x280 & ~x312 & ~x313 & ~x331 & ~x333 & ~x337 & ~x338 & ~x339 & ~x359 & ~x366 & ~x368 & ~x389 & ~x390 & ~x392 & ~x395 & ~x396 & ~x415 & ~x416 & ~x418 & ~x419 & ~x421 & ~x426 & ~x443 & ~x447 & ~x449 & ~x452 & ~x473 & ~x479 & ~x495 & ~x496 & ~x500 & ~x501 & ~x507 & ~x510 & ~x526 & ~x530 & ~x533 & ~x542 & ~x543 & ~x555 & ~x556 & ~x558 & ~x561 & ~x563 & ~x569 & ~x570 & ~x571 & ~x586 & ~x589 & ~x594 & ~x597 & ~x608 & ~x610 & ~x611 & ~x618 & ~x620 & ~x621 & ~x623 & ~x636 & ~x639 & ~x640 & ~x642 & ~x645 & ~x651 & ~x664 & ~x668 & ~x669 & ~x671 & ~x672 & ~x676 & ~x677 & ~x694 & ~x708 & ~x719 & ~x720 & ~x721 & ~x732 & ~x734 & ~x739 & ~x741 & ~x743 & ~x744 & ~x745 & ~x748 & ~x751 & ~x755 & ~x757 & ~x767 & ~x768 & ~x772 & ~x776 & ~x778 & ~x781;
assign c4198 =  x756;
assign c4200 =  x375 & ~x2 & ~x3 & ~x6 & ~x10 & ~x13 & ~x15 & ~x18 & ~x20 & ~x23 & ~x26 & ~x29 & ~x30 & ~x35 & ~x39 & ~x45 & ~x50 & ~x52 & ~x64 & ~x71 & ~x72 & ~x73 & ~x77 & ~x87 & ~x89 & ~x93 & ~x96 & ~x97 & ~x99 & ~x105 & ~x106 & ~x107 & ~x114 & ~x117 & ~x118 & ~x133 & ~x147 & ~x164 & ~x172 & ~x175 & ~x192 & ~x194 & ~x195 & ~x197 & ~x198 & ~x199 & ~x201 & ~x205 & ~x220 & ~x221 & ~x224 & ~x227 & ~x245 & ~x247 & ~x248 & ~x249 & ~x252 & ~x255 & ~x256 & ~x257 & ~x258 & ~x274 & ~x277 & ~x278 & ~x280 & ~x281 & ~x283 & ~x284 & ~x286 & ~x287 & ~x288 & ~x307 & ~x308 & ~x311 & ~x333 & ~x336 & ~x338 & ~x360 & ~x362 & ~x364 & ~x369 & ~x391 & ~x393 & ~x394 & ~x419 & ~x422 & ~x449 & ~x452 & ~x453 & ~x470 & ~x475 & ~x477 & ~x479 & ~x481 & ~x498 & ~x503 & ~x525 & ~x526 & ~x556 & ~x557 & ~x562 & ~x563 & ~x572 & ~x590 & ~x591 & ~x592 & ~x600 & ~x616 & ~x628 & ~x640 & ~x641 & ~x644 & ~x647 & ~x654 & ~x655 & ~x665 & ~x672 & ~x673 & ~x677 & ~x679 & ~x680 & ~x690 & ~x694 & ~x695 & ~x712 & ~x713 & ~x716 & ~x717 & ~x719 & ~x720 & ~x723 & ~x732 & ~x733 & ~x735 & ~x738 & ~x739 & ~x741 & ~x743 & ~x744 & ~x745 & ~x750 & ~x751 & ~x753 & ~x756 & ~x761 & ~x764 & ~x765 & ~x766 & ~x769 & ~x771 & ~x773 & ~x774 & ~x777 & ~x783;
assign c4202 = ~x3 & ~x9 & ~x20 & ~x21 & ~x24 & ~x33 & ~x34 & ~x42 & ~x44 & ~x47 & ~x51 & ~x55 & ~x64 & ~x68 & ~x71 & ~x73 & ~x81 & ~x82 & ~x91 & ~x94 & ~x95 & ~x97 & ~x102 & ~x107 & ~x109 & ~x112 & ~x114 & ~x130 & ~x139 & ~x144 & ~x145 & ~x150 & ~x151 & ~x166 & ~x179 & ~x180 & ~x201 & ~x208 & ~x215 & ~x216 & ~x218 & ~x219 & ~x220 & ~x243 & ~x249 & ~x254 & ~x255 & ~x256 & ~x257 & ~x271 & ~x275 & ~x279 & ~x283 & ~x306 & ~x309 & ~x310 & ~x311 & ~x331 & ~x335 & ~x338 & ~x341 & ~x366 & ~x367 & ~x390 & ~x391 & ~x393 & ~x397 & ~x420 & ~x444 & ~x471 & ~x472 & ~x473 & ~x480 & ~x497 & ~x502 & ~x504 & ~x524 & ~x527 & ~x537 & ~x538 & ~x554 & ~x556 & ~x558 & ~x565 & ~x568 & ~x570 & ~x593 & ~x597 & ~x615 & ~x622 & ~x642 & ~x645 & ~x646 & ~x648 & ~x650 & ~x652 & ~x653 & ~x672 & ~x677 & ~x681 & ~x685 & ~x709 & ~x713 & ~x716 & ~x724 & ~x728 & ~x730 & ~x732 & ~x737 & ~x740 & ~x741 & ~x742 & ~x746 & ~x747 & ~x749 & ~x751 & ~x779 & ~x780;
assign c4204 =  x361;
assign c4206 =  x427 &  x430 &  x457 &  x458 &  x459 &  x460 &  x464 &  x465 &  x467 & ~x331 & ~x541 & ~x543;
assign c4208 =  x465 & ~x36 & ~x44 & ~x48 & ~x57 & ~x58 & ~x60 & ~x63 & ~x67 & ~x70 & ~x73 & ~x75 & ~x77 & ~x83 & ~x84 & ~x85 & ~x92 & ~x94 & ~x98 & ~x115 & ~x119 & ~x120 & ~x125 & ~x126 & ~x136 & ~x143 & ~x155 & ~x166 & ~x182 & ~x196 & ~x198 & ~x210 & ~x266 & ~x277 & ~x278 & ~x283 & ~x307 & ~x321 & ~x337 & ~x339 & ~x360 & ~x389 & ~x391 & ~x419 & ~x423 & ~x472 & ~x480 & ~x500 & ~x503 & ~x507 & ~x534 & ~x535 & ~x562 & ~x563 & ~x585 & ~x587 & ~x616 & ~x620 & ~x647 & ~x666 & ~x671 & ~x706 & ~x718 & ~x719 & ~x724 & ~x729 & ~x734 & ~x740 & ~x756 & ~x759 & ~x767 & ~x772 & ~x778 & ~x779 & ~x782;
assign c4210 = ~x2 & ~x3 & ~x4 & ~x7 & ~x12 & ~x13 & ~x16 & ~x17 & ~x18 & ~x20 & ~x27 & ~x29 & ~x30 & ~x34 & ~x35 & ~x38 & ~x39 & ~x41 & ~x44 & ~x48 & ~x50 & ~x55 & ~x58 & ~x65 & ~x68 & ~x69 & ~x70 & ~x71 & ~x72 & ~x76 & ~x78 & ~x82 & ~x83 & ~x85 & ~x88 & ~x92 & ~x94 & ~x99 & ~x109 & ~x112 & ~x115 & ~x121 & ~x129 & ~x130 & ~x134 & ~x135 & ~x138 & ~x140 & ~x153 & ~x164 & ~x166 & ~x171 & ~x172 & ~x173 & ~x181 & ~x200 & ~x219 & ~x223 & ~x226 & ~x237 & ~x253 & ~x254 & ~x264 & ~x277 & ~x279 & ~x280 & ~x307 & ~x310 & ~x311 & ~x333 & ~x339 & ~x360 & ~x363 & ~x365 & ~x366 & ~x368 & ~x388 & ~x389 & ~x417 & ~x419 & ~x421 & ~x424 & ~x443 & ~x448 & ~x449 & ~x450 & ~x451 & ~x472 & ~x474 & ~x500 & ~x501 & ~x502 & ~x512 & ~x514 & ~x515 & ~x535 & ~x543 & ~x562 & ~x568 & ~x569 & ~x570 & ~x583 & ~x585 & ~x587 & ~x589 & ~x594 & ~x595 & ~x597 & ~x609 & ~x611 & ~x612 & ~x615 & ~x616 & ~x622 & ~x636 & ~x639 & ~x644 & ~x647 & ~x648 & ~x649 & ~x652 & ~x665 & ~x666 & ~x671 & ~x672 & ~x675 & ~x677 & ~x678 & ~x693 & ~x694 & ~x695 & ~x696 & ~x707 & ~x708 & ~x710 & ~x718 & ~x720 & ~x724 & ~x725 & ~x738 & ~x740 & ~x751 & ~x767 & ~x769 & ~x772 & ~x774 & ~x775 & ~x777 & ~x779 & ~x783;
assign c4212 = ~x43 & ~x56 & ~x66 & ~x76 & ~x98 & ~x104 & ~x116 & ~x153 & ~x189 & ~x208 & ~x209 & ~x238 & ~x246 & ~x248 & ~x264 & ~x292 & ~x301 & ~x321 & ~x479 & ~x573 & ~x598 & ~x650 & ~x651 & ~x684 & ~x727;
assign c4214 =  x437 & ~x0 & ~x1 & ~x9 & ~x13 & ~x32 & ~x53 & ~x61 & ~x62 & ~x70 & ~x81 & ~x87 & ~x89 & ~x91 & ~x92 & ~x94 & ~x96 & ~x99 & ~x100 & ~x109 & ~x110 & ~x114 & ~x116 & ~x118 & ~x122 & ~x123 & ~x126 & ~x129 & ~x140 & ~x141 & ~x143 & ~x144 & ~x150 & ~x157 & ~x172 & ~x176 & ~x196 & ~x198 & ~x213 & ~x223 & ~x227 & ~x229 & ~x252 & ~x269 & ~x280 & ~x283 & ~x286 & ~x296 & ~x309 & ~x311 & ~x313 & ~x324 & ~x360 & ~x367 & ~x389 & ~x396 & ~x420 & ~x421 & ~x423 & ~x445 & ~x473 & ~x474 & ~x475 & ~x479 & ~x502 & ~x524 & ~x525 & ~x527 & ~x534 & ~x535 & ~x536 & ~x551 & ~x553 & ~x555 & ~x565 & ~x581 & ~x584 & ~x586 & ~x587 & ~x594 & ~x612 & ~x616 & ~x617 & ~x637 & ~x642 & ~x674 & ~x697 & ~x700 & ~x703 & ~x720 & ~x727 & ~x733 & ~x749 & ~x754 & ~x756 & ~x759 & ~x764 & ~x772 & ~x773 & ~x778;
assign c4216 =  x493 &  x521 &  x606 & ~x179 & ~x207 & ~x235;
assign c4218 =  x0;
assign c4220 = ~x2 & ~x3 & ~x7 & ~x25 & ~x27 & ~x34 & ~x38 & ~x42 & ~x44 & ~x47 & ~x49 & ~x51 & ~x58 & ~x62 & ~x68 & ~x72 & ~x77 & ~x92 & ~x97 & ~x102 & ~x112 & ~x139 & ~x143 & ~x155 & ~x183 & ~x196 & ~x197 & ~x209 & ~x210 & ~x224 & ~x227 & ~x237 & ~x238 & ~x250 & ~x254 & ~x265 & ~x303 & ~x304 & ~x306 & ~x321 & ~x331 & ~x390 & ~x392 & ~x421 & ~x444 & ~x448 & ~x449 & ~x503 & ~x530 & ~x558 & ~x561 & ~x562 & ~x563 & ~x568 & ~x573 & ~x589 & ~x592 & ~x614 & ~x618 & ~x619 & ~x624 & ~x628 & ~x641 & ~x656 & ~x668 & ~x669 & ~x678 & ~x701 & ~x705 & ~x721 & ~x722 & ~x723 & ~x728 & ~x729 & ~x737 & ~x743 & ~x744 & ~x745 & ~x746 & ~x747 & ~x749 & ~x754 & ~x769 & ~x774;
assign c4222 =  x466 & ~x0 & ~x3 & ~x8 & ~x9 & ~x10 & ~x14 & ~x16 & ~x17 & ~x19 & ~x20 & ~x21 & ~x29 & ~x31 & ~x36 & ~x37 & ~x39 & ~x43 & ~x44 & ~x45 & ~x47 & ~x49 & ~x50 & ~x53 & ~x54 & ~x56 & ~x61 & ~x62 & ~x66 & ~x71 & ~x74 & ~x75 & ~x76 & ~x77 & ~x78 & ~x81 & ~x85 & ~x88 & ~x89 & ~x90 & ~x91 & ~x101 & ~x107 & ~x109 & ~x112 & ~x139 & ~x144 & ~x146 & ~x166 & ~x168 & ~x173 & ~x196 & ~x197 & ~x198 & ~x199 & ~x219 & ~x220 & ~x223 & ~x224 & ~x226 & ~x227 & ~x249 & ~x252 & ~x254 & ~x278 & ~x304 & ~x306 & ~x310 & ~x332 & ~x334 & ~x336 & ~x337 & ~x339 & ~x361 & ~x367 & ~x394 & ~x395 & ~x419 & ~x422 & ~x445 & ~x447 & ~x448 & ~x475 & ~x476 & ~x477 & ~x479 & ~x502 & ~x504 & ~x507 & ~x529 & ~x533 & ~x534 & ~x536 & ~x554 & ~x555 & ~x557 & ~x558 & ~x559 & ~x561 & ~x562 & ~x564 & ~x574 & ~x587 & ~x588 & ~x596 & ~x597 & ~x600 & ~x601 & ~x614 & ~x617 & ~x619 & ~x621 & ~x625 & ~x627 & ~x628 & ~x629 & ~x641 & ~x642 & ~x645 & ~x647 & ~x649 & ~x650 & ~x658 & ~x659 & ~x670 & ~x673 & ~x675 & ~x676 & ~x677 & ~x678 & ~x681 & ~x682 & ~x685 & ~x688 & ~x693 & ~x695 & ~x701 & ~x709 & ~x712 & ~x715 & ~x718 & ~x719 & ~x721 & ~x728 & ~x729 & ~x732 & ~x733 & ~x734 & ~x735 & ~x738 & ~x741 & ~x742 & ~x744 & ~x751 & ~x752 & ~x754 & ~x755 & ~x763 & ~x767 & ~x771 & ~x777;
assign c4224 =  x401 &  x455 &  x456 &  x491 & ~x2 & ~x17 & ~x21 & ~x22 & ~x28 & ~x33 & ~x38 & ~x60 & ~x66 & ~x73 & ~x74 & ~x85 & ~x87 & ~x91 & ~x100 & ~x101 & ~x104 & ~x115 & ~x116 & ~x118 & ~x122 & ~x123 & ~x125 & ~x130 & ~x144 & ~x146 & ~x147 & ~x148 & ~x150 & ~x151 & ~x169 & ~x170 & ~x175 & ~x178 & ~x195 & ~x200 & ~x207 & ~x255 & ~x278 & ~x283 & ~x306 & ~x334 & ~x336 & ~x359 & ~x364 & ~x366 & ~x368 & ~x419 & ~x531 & ~x535 & ~x555 & ~x556 & ~x584 & ~x585 & ~x588 & ~x593 & ~x595 & ~x611 & ~x612 & ~x613 & ~x616 & ~x618 & ~x619 & ~x620 & ~x621 & ~x638 & ~x647 & ~x649 & ~x673 & ~x675 & ~x676 & ~x689 & ~x694 & ~x703 & ~x705 & ~x708 & ~x709 & ~x710 & ~x723 & ~x729 & ~x731 & ~x732 & ~x737 & ~x738 & ~x741 & ~x742 & ~x748 & ~x751 & ~x757 & ~x761 & ~x762 & ~x764 & ~x766 & ~x773 & ~x774 & ~x775 & ~x778 & ~x783;
assign c4226 =  x409 & ~x17 & ~x24 & ~x27 & ~x30 & ~x39 & ~x41 & ~x43 & ~x47 & ~x51 & ~x52 & ~x55 & ~x56 & ~x58 & ~x68 & ~x69 & ~x71 & ~x73 & ~x74 & ~x84 & ~x90 & ~x100 & ~x102 & ~x103 & ~x105 & ~x118 & ~x123 & ~x128 & ~x142 & ~x147 & ~x151 & ~x161 & ~x165 & ~x168 & ~x170 & ~x174 & ~x195 & ~x196 & ~x197 & ~x199 & ~x201 & ~x202 & ~x215 & ~x216 & ~x221 & ~x243 & ~x250 & ~x276 & ~x278 & ~x298 & ~x313 & ~x334 & ~x336 & ~x341 & ~x364 & ~x366 & ~x389 & ~x420 & ~x424 & ~x443 & ~x445 & ~x468 & ~x471 & ~x501 & ~x502 & ~x503 & ~x507 & ~x513 & ~x522 & ~x526 & ~x528 & ~x531 & ~x532 & ~x541 & ~x551 & ~x553 & ~x554 & ~x561 & ~x563 & ~x567 & ~x580 & ~x622 & ~x623 & ~x645 & ~x648 & ~x650 & ~x672 & ~x675 & ~x679 & ~x691 & ~x697 & ~x722 & ~x734 & ~x736 & ~x742 & ~x749 & ~x754 & ~x755 & ~x758 & ~x759 & ~x760 & ~x761 & ~x765 & ~x768;
assign c4228 = ~x1 & ~x2 & ~x5 & ~x8 & ~x9 & ~x10 & ~x13 & ~x15 & ~x17 & ~x18 & ~x19 & ~x20 & ~x21 & ~x23 & ~x24 & ~x27 & ~x32 & ~x34 & ~x35 & ~x36 & ~x37 & ~x38 & ~x44 & ~x45 & ~x46 & ~x48 & ~x51 & ~x52 & ~x54 & ~x55 & ~x58 & ~x60 & ~x64 & ~x67 & ~x69 & ~x70 & ~x71 & ~x73 & ~x75 & ~x76 & ~x78 & ~x79 & ~x81 & ~x82 & ~x83 & ~x84 & ~x86 & ~x89 & ~x92 & ~x96 & ~x97 & ~x100 & ~x102 & ~x106 & ~x110 & ~x113 & ~x114 & ~x115 & ~x118 & ~x120 & ~x128 & ~x135 & ~x136 & ~x139 & ~x140 & ~x141 & ~x145 & ~x146 & ~x147 & ~x155 & ~x156 & ~x163 & ~x166 & ~x169 & ~x170 & ~x172 & ~x173 & ~x183 & ~x194 & ~x195 & ~x200 & ~x211 & ~x222 & ~x229 & ~x239 & ~x249 & ~x250 & ~x251 & ~x253 & ~x254 & ~x255 & ~x256 & ~x267 & ~x280 & ~x281 & ~x283 & ~x285 & ~x309 & ~x312 & ~x322 & ~x333 & ~x334 & ~x336 & ~x337 & ~x338 & ~x340 & ~x350 & ~x361 & ~x362 & ~x364 & ~x367 & ~x388 & ~x391 & ~x392 & ~x393 & ~x394 & ~x414 & ~x417 & ~x418 & ~x421 & ~x424 & ~x443 & ~x446 & ~x447 & ~x448 & ~x451 & ~x452 & ~x453 & ~x472 & ~x474 & ~x475 & ~x476 & ~x477 & ~x499 & ~x500 & ~x501 & ~x504 & ~x506 & ~x507 & ~x530 & ~x532 & ~x533 & ~x535 & ~x536 & ~x562 & ~x564 & ~x583 & ~x584 & ~x586 & ~x587 & ~x589 & ~x590 & ~x593 & ~x595 & ~x613 & ~x614 & ~x615 & ~x620 & ~x621 & ~x641 & ~x642 & ~x643 & ~x644 & ~x646 & ~x651 & ~x652 & ~x668 & ~x669 & ~x670 & ~x672 & ~x673 & ~x674 & ~x675 & ~x677 & ~x678 & ~x679 & ~x682 & ~x683 & ~x697 & ~x701 & ~x702 & ~x703 & ~x704 & ~x705 & ~x706 & ~x708 & ~x712 & ~x717 & ~x718 & ~x722 & ~x728 & ~x729 & ~x730 & ~x731 & ~x738 & ~x739 & ~x740 & ~x741 & ~x742 & ~x743 & ~x744 & ~x745 & ~x749 & ~x750 & ~x751 & ~x755 & ~x756 & ~x758 & ~x760 & ~x761 & ~x764 & ~x773 & ~x774 & ~x783;
assign c4230 =  x83;
assign c4232 = ~x0 & ~x1 & ~x2 & ~x4 & ~x8 & ~x12 & ~x13 & ~x15 & ~x16 & ~x18 & ~x20 & ~x32 & ~x33 & ~x35 & ~x38 & ~x41 & ~x45 & ~x47 & ~x48 & ~x53 & ~x55 & ~x59 & ~x60 & ~x67 & ~x70 & ~x72 & ~x80 & ~x82 & ~x84 & ~x86 & ~x100 & ~x106 & ~x107 & ~x108 & ~x111 & ~x112 & ~x129 & ~x133 & ~x137 & ~x145 & ~x156 & ~x163 & ~x183 & ~x184 & ~x195 & ~x221 & ~x239 & ~x266 & ~x279 & ~x294 & ~x308 & ~x310 & ~x332 & ~x350 & ~x351 & ~x362 & ~x388 & ~x390 & ~x444 & ~x451 & ~x471 & ~x498 & ~x499 & ~x500 & ~x501 & ~x527 & ~x528 & ~x529 & ~x531 & ~x534 & ~x535 & ~x556 & ~x563 & ~x566 & ~x584 & ~x585 & ~x592 & ~x593 & ~x611 & ~x615 & ~x616 & ~x642 & ~x647 & ~x649 & ~x668 & ~x672 & ~x680 & ~x693 & ~x695 & ~x716 & ~x717 & ~x719 & ~x721 & ~x725 & ~x726 & ~x732 & ~x744 & ~x745 & ~x746 & ~x748 & ~x749 & ~x757 & ~x758 & ~x766 & ~x775;
assign c4234 =  x379 &  x406 & ~x17 & ~x29 & ~x51 & ~x55 & ~x84 & ~x85 & ~x99 & ~x101 & ~x125 & ~x129 & ~x148 & ~x157 & ~x172 & ~x212 & ~x267 & ~x335 & ~x341 & ~x366 & ~x388 & ~x392 & ~x511 & ~x539 & ~x548 & ~x551 & ~x567 & ~x576 & ~x588 & ~x620 & ~x661 & ~x668 & ~x707 & ~x729 & ~x746 & ~x759 & ~x773 & ~x775 & ~x776 & ~x779;
assign c4236 =  x26 &  x445;
assign c4238 =  x293 &  x409 &  x464 & ~x12 & ~x14 & ~x18 & ~x21 & ~x22 & ~x32 & ~x34 & ~x37 & ~x46 & ~x47 & ~x49 & ~x66 & ~x71 & ~x84 & ~x92 & ~x105 & ~x119 & ~x123 & ~x140 & ~x167 & ~x176 & ~x205 & ~x206 & ~x218 & ~x219 & ~x222 & ~x226 & ~x233 & ~x234 & ~x246 & ~x247 & ~x250 & ~x258 & ~x261 & ~x274 & ~x280 & ~x288 & ~x289 & ~x303 & ~x329 & ~x336 & ~x337 & ~x390 & ~x417 & ~x502 & ~x505 & ~x506 & ~x528 & ~x582 & ~x594 & ~x597 & ~x599 & ~x610 & ~x611 & ~x616 & ~x624 & ~x626 & ~x627 & ~x640 & ~x646 & ~x651 & ~x654 & ~x673 & ~x676 & ~x678 & ~x681 & ~x682 & ~x683 & ~x700 & ~x703 & ~x706 & ~x708 & ~x709 & ~x710 & ~x711 & ~x713 & ~x714 & ~x718 & ~x730 & ~x740 & ~x745 & ~x749 & ~x750 & ~x753 & ~x763 & ~x765 & ~x774 & ~x778 & ~x779;
assign c4240 =  x272 & ~x0 & ~x3 & ~x7 & ~x14 & ~x17 & ~x22 & ~x25 & ~x27 & ~x32 & ~x35 & ~x39 & ~x42 & ~x43 & ~x47 & ~x48 & ~x51 & ~x53 & ~x55 & ~x59 & ~x60 & ~x69 & ~x73 & ~x77 & ~x82 & ~x83 & ~x88 & ~x91 & ~x104 & ~x105 & ~x109 & ~x111 & ~x115 & ~x120 & ~x129 & ~x130 & ~x132 & ~x139 & ~x144 & ~x147 & ~x166 & ~x170 & ~x171 & ~x174 & ~x176 & ~x186 & ~x194 & ~x199 & ~x201 & ~x202 & ~x226 & ~x228 & ~x241 & ~x277 & ~x284 & ~x285 & ~x295 & ~x304 & ~x308 & ~x333 & ~x336 & ~x338 & ~x339 & ~x359 & ~x363 & ~x366 & ~x395 & ~x421 & ~x422 & ~x447 & ~x450 & ~x451 & ~x502 & ~x505 & ~x508 & ~x537 & ~x558 & ~x560 & ~x561 & ~x562 & ~x564 & ~x589 & ~x592 & ~x594 & ~x610 & ~x613 & ~x615 & ~x616 & ~x621 & ~x661 & ~x662 & ~x665 & ~x667 & ~x669 & ~x672 & ~x677 & ~x699 & ~x702 & ~x715 & ~x723 & ~x727 & ~x730 & ~x731 & ~x735 & ~x742 & ~x744 & ~x746 & ~x754 & ~x755 & ~x757 & ~x763 & ~x765 & ~x767 & ~x768 & ~x771 & ~x772 & ~x773 & ~x777 & ~x778;
assign c4242 =  x757;
assign c4244 =  x193 &  x640;
assign c4246 =  x356 &  x411 & ~x3 & ~x14 & ~x18 & ~x22 & ~x23 & ~x26 & ~x40 & ~x48 & ~x50 & ~x53 & ~x56 & ~x57 & ~x58 & ~x63 & ~x65 & ~x70 & ~x71 & ~x77 & ~x80 & ~x81 & ~x83 & ~x89 & ~x93 & ~x94 & ~x96 & ~x99 & ~x101 & ~x102 & ~x107 & ~x114 & ~x116 & ~x121 & ~x123 & ~x124 & ~x127 & ~x128 & ~x129 & ~x157 & ~x167 & ~x168 & ~x184 & ~x185 & ~x212 & ~x222 & ~x250 & ~x253 & ~x279 & ~x295 & ~x306 & ~x307 & ~x364 & ~x388 & ~x389 & ~x391 & ~x419 & ~x445 & ~x474 & ~x501 & ~x503 & ~x506 & ~x533 & ~x535 & ~x559 & ~x560 & ~x561 & ~x564 & ~x587 & ~x588 & ~x615 & ~x620 & ~x640 & ~x643 & ~x649 & ~x651 & ~x673 & ~x696 & ~x703 & ~x720 & ~x724 & ~x728 & ~x736 & ~x743 & ~x746 & ~x747 & ~x754 & ~x760 & ~x768 & ~x774 & ~x776 & ~x782;
assign c4248 =  x464 & ~x1 & ~x4 & ~x6 & ~x8 & ~x11 & ~x12 & ~x16 & ~x21 & ~x28 & ~x29 & ~x31 & ~x36 & ~x45 & ~x47 & ~x56 & ~x62 & ~x63 & ~x66 & ~x73 & ~x78 & ~x85 & ~x87 & ~x90 & ~x92 & ~x94 & ~x95 & ~x96 & ~x102 & ~x104 & ~x113 & ~x117 & ~x124 & ~x130 & ~x138 & ~x142 & ~x150 & ~x161 & ~x162 & ~x166 & ~x167 & ~x170 & ~x171 & ~x178 & ~x197 & ~x222 & ~x227 & ~x235 & ~x245 & ~x248 & ~x275 & ~x284 & ~x308 & ~x327 & ~x330 & ~x333 & ~x334 & ~x338 & ~x355 & ~x357 & ~x359 & ~x362 & ~x389 & ~x392 & ~x393 & ~x395 & ~x418 & ~x445 & ~x447 & ~x451 & ~x473 & ~x474 & ~x501 & ~x502 & ~x505 & ~x532 & ~x555 & ~x560 & ~x572 & ~x588 & ~x591 & ~x592 & ~x594 & ~x596 & ~x597 & ~x598 & ~x602 & ~x612 & ~x619 & ~x620 & ~x621 & ~x622 & ~x623 & ~x627 & ~x629 & ~x640 & ~x645 & ~x658 & ~x669 & ~x677 & ~x679 & ~x702 & ~x706 & ~x711 & ~x726 & ~x728 & ~x729 & ~x739 & ~x740 & ~x741 & ~x744 & ~x749 & ~x751 & ~x756 & ~x760 & ~x761 & ~x766 & ~x771 & ~x772 & ~x774 & ~x782 & ~x783;
assign c4250 =  x320 &  x347 &  x380 &  x408 &  x435 &  x462 & ~x3 & ~x29 & ~x39 & ~x52 & ~x55 & ~x65 & ~x76 & ~x79 & ~x80 & ~x127 & ~x144 & ~x151 & ~x171 & ~x176 & ~x177 & ~x179 & ~x195 & ~x201 & ~x202 & ~x232 & ~x253 & ~x257 & ~x314 & ~x362 & ~x364 & ~x367 & ~x395 & ~x398 & ~x453 & ~x521 & ~x524 & ~x552 & ~x565 & ~x567 & ~x575 & ~x576 & ~x591 & ~x612 & ~x616 & ~x630 & ~x668 & ~x686 & ~x689 & ~x690 & ~x691 & ~x705 & ~x707 & ~x722 & ~x732 & ~x736 & ~x752 & ~x760 & ~x772;
assign c4252 =  x465 &  x466 & ~x6 & ~x9 & ~x58 & ~x63 & ~x70 & ~x74 & ~x91 & ~x101 & ~x107 & ~x120 & ~x125 & ~x135 & ~x138 & ~x145 & ~x151 & ~x166 & ~x199 & ~x206 & ~x226 & ~x234 & ~x257 & ~x285 & ~x309 & ~x316 & ~x333 & ~x339 & ~x421 & ~x444 & ~x451 & ~x481 & ~x510 & ~x539 & ~x542 & ~x558 & ~x560 & ~x567 & ~x569 & ~x622 & ~x644 & ~x699 & ~x704 & ~x722 & ~x726 & ~x757 & ~x780;
assign c4254 =  x400 & ~x9 & ~x13 & ~x26 & ~x32 & ~x39 & ~x40 & ~x48 & ~x56 & ~x64 & ~x68 & ~x71 & ~x81 & ~x91 & ~x93 & ~x103 & ~x107 & ~x113 & ~x118 & ~x136 & ~x142 & ~x148 & ~x166 & ~x170 & ~x229 & ~x250 & ~x256 & ~x282 & ~x283 & ~x304 & ~x360 & ~x366 & ~x377 & ~x390 & ~x416 & ~x418 & ~x445 & ~x447 & ~x449 & ~x473 & ~x474 & ~x478 & ~x529 & ~x559 & ~x560 & ~x586 & ~x590 & ~x600 & ~x613 & ~x626 & ~x656 & ~x668 & ~x672 & ~x674 & ~x676 & ~x679 & ~x686 & ~x687 & ~x693 & ~x696 & ~x700 & ~x706 & ~x708 & ~x710 & ~x712 & ~x719 & ~x723 & ~x736 & ~x745 & ~x752 & ~x755 & ~x763 & ~x771;
assign c4256 =  x701;
assign c4258 =  x374 &  x457 &  x490 & ~x2 & ~x18 & ~x36 & ~x51 & ~x60 & ~x69 & ~x79 & ~x80 & ~x83 & ~x86 & ~x90 & ~x97 & ~x99 & ~x140 & ~x145 & ~x146 & ~x203 & ~x204 & ~x247 & ~x248 & ~x256 & ~x258 & ~x333 & ~x360 & ~x361 & ~x386 & ~x389 & ~x424 & ~x425 & ~x477 & ~x480 & ~x506 & ~x527 & ~x533 & ~x556 & ~x562 & ~x589 & ~x592 & ~x610 & ~x611 & ~x664 & ~x672 & ~x684 & ~x691 & ~x742 & ~x744 & ~x747 & ~x776 & ~x780;
assign c4260 =  x268 & ~x0 & ~x5 & ~x15 & ~x19 & ~x20 & ~x23 & ~x25 & ~x27 & ~x29 & ~x30 & ~x32 & ~x34 & ~x40 & ~x43 & ~x45 & ~x46 & ~x48 & ~x52 & ~x55 & ~x57 & ~x58 & ~x62 & ~x66 & ~x69 & ~x73 & ~x76 & ~x81 & ~x85 & ~x86 & ~x87 & ~x94 & ~x98 & ~x104 & ~x106 & ~x114 & ~x115 & ~x117 & ~x121 & ~x123 & ~x124 & ~x133 & ~x136 & ~x138 & ~x140 & ~x141 & ~x144 & ~x147 & ~x150 & ~x151 & ~x152 & ~x164 & ~x180 & ~x191 & ~x192 & ~x193 & ~x195 & ~x217 & ~x219 & ~x223 & ~x226 & ~x237 & ~x244 & ~x248 & ~x251 & ~x255 & ~x256 & ~x265 & ~x272 & ~x274 & ~x276 & ~x280 & ~x283 & ~x301 & ~x302 & ~x303 & ~x306 & ~x310 & ~x332 & ~x333 & ~x334 & ~x337 & ~x338 & ~x391 & ~x394 & ~x417 & ~x418 & ~x420 & ~x421 & ~x422 & ~x475 & ~x499 & ~x502 & ~x526 & ~x528 & ~x533 & ~x536 & ~x559 & ~x561 & ~x563 & ~x564 & ~x565 & ~x584 & ~x593 & ~x611 & ~x614 & ~x619 & ~x623 & ~x624 & ~x647 & ~x649 & ~x652 & ~x669 & ~x672 & ~x676 & ~x677 & ~x695 & ~x696 & ~x705 & ~x729 & ~x738 & ~x740 & ~x741 & ~x742 & ~x746 & ~x747 & ~x751 & ~x754 & ~x755 & ~x757 & ~x762 & ~x763 & ~x764 & ~x776 & ~x779 & ~x780 & ~x783;
assign c4262 =  x325 &  x353 &  x409 &  x436 &  x464 & ~x4 & ~x7 & ~x12 & ~x13 & ~x17 & ~x18 & ~x19 & ~x21 & ~x24 & ~x27 & ~x28 & ~x29 & ~x32 & ~x36 & ~x38 & ~x40 & ~x41 & ~x42 & ~x43 & ~x44 & ~x45 & ~x48 & ~x51 & ~x52 & ~x54 & ~x60 & ~x62 & ~x69 & ~x72 & ~x73 & ~x74 & ~x75 & ~x77 & ~x78 & ~x87 & ~x88 & ~x89 & ~x91 & ~x93 & ~x96 & ~x97 & ~x99 & ~x100 & ~x107 & ~x109 & ~x114 & ~x118 & ~x121 & ~x125 & ~x135 & ~x136 & ~x139 & ~x143 & ~x145 & ~x153 & ~x164 & ~x165 & ~x166 & ~x167 & ~x168 & ~x169 & ~x170 & ~x172 & ~x175 & ~x181 & ~x194 & ~x195 & ~x198 & ~x199 & ~x200 & ~x209 & ~x218 & ~x220 & ~x223 & ~x226 & ~x227 & ~x246 & ~x248 & ~x250 & ~x253 & ~x255 & ~x256 & ~x257 & ~x273 & ~x276 & ~x280 & ~x282 & ~x283 & ~x285 & ~x301 & ~x302 & ~x306 & ~x308 & ~x309 & ~x312 & ~x313 & ~x329 & ~x331 & ~x332 & ~x337 & ~x339 & ~x359 & ~x360 & ~x361 & ~x362 & ~x366 & ~x367 & ~x369 & ~x387 & ~x390 & ~x396 & ~x397 & ~x416 & ~x417 & ~x418 & ~x421 & ~x422 & ~x423 & ~x446 & ~x450 & ~x452 & ~x474 & ~x501 & ~x504 & ~x506 & ~x507 & ~x561 & ~x564 & ~x582 & ~x583 & ~x585 & ~x588 & ~x589 & ~x591 & ~x592 & ~x593 & ~x609 & ~x610 & ~x612 & ~x614 & ~x615 & ~x616 & ~x617 & ~x620 & ~x621 & ~x622 & ~x638 & ~x639 & ~x640 & ~x641 & ~x643 & ~x644 & ~x649 & ~x651 & ~x652 & ~x653 & ~x654 & ~x665 & ~x666 & ~x668 & ~x669 & ~x670 & ~x675 & ~x678 & ~x680 & ~x694 & ~x704 & ~x706 & ~x707 & ~x709 & ~x710 & ~x720 & ~x722 & ~x723 & ~x725 & ~x728 & ~x730 & ~x731 & ~x735 & ~x737 & ~x739 & ~x743 & ~x746 & ~x749 & ~x757 & ~x760 & ~x761 & ~x762 & ~x765 & ~x767 & ~x768 & ~x770 & ~x774 & ~x775 & ~x776 & ~x777 & ~x782 & ~x783;
assign c4264 =  x191;
assign c4266 =  x490 &  x491 & ~x1 & ~x5 & ~x6 & ~x11 & ~x19 & ~x21 & ~x25 & ~x26 & ~x27 & ~x31 & ~x35 & ~x38 & ~x41 & ~x47 & ~x51 & ~x53 & ~x54 & ~x60 & ~x64 & ~x67 & ~x71 & ~x74 & ~x78 & ~x79 & ~x81 & ~x84 & ~x89 & ~x90 & ~x91 & ~x92 & ~x93 & ~x100 & ~x109 & ~x110 & ~x116 & ~x119 & ~x123 & ~x137 & ~x138 & ~x142 & ~x145 & ~x165 & ~x167 & ~x168 & ~x176 & ~x178 & ~x197 & ~x199 & ~x200 & ~x201 & ~x202 & ~x203 & ~x218 & ~x226 & ~x228 & ~x230 & ~x231 & ~x246 & ~x247 & ~x251 & ~x254 & ~x257 & ~x258 & ~x259 & ~x274 & ~x276 & ~x284 & ~x288 & ~x306 & ~x311 & ~x314 & ~x315 & ~x334 & ~x335 & ~x338 & ~x341 & ~x342 & ~x358 & ~x362 & ~x367 & ~x385 & ~x388 & ~x391 & ~x392 & ~x397 & ~x449 & ~x505 & ~x528 & ~x534 & ~x554 & ~x558 & ~x560 & ~x563 & ~x581 & ~x584 & ~x587 & ~x590 & ~x592 & ~x595 & ~x599 & ~x610 & ~x615 & ~x621 & ~x622 & ~x644 & ~x646 & ~x653 & ~x665 & ~x672 & ~x674 & ~x692 & ~x695 & ~x703 & ~x710 & ~x715 & ~x719 & ~x728 & ~x732 & ~x738 & ~x739 & ~x740 & ~x741 & ~x743 & ~x746 & ~x747 & ~x750 & ~x751 & ~x752 & ~x755 & ~x757 & ~x760 & ~x762 & ~x764 & ~x767 & ~x772 & ~x777 & ~x780 & ~x783;
assign c4268 =  x401 &  x408 &  x436 & ~x0 & ~x6 & ~x11 & ~x13 & ~x16 & ~x19 & ~x22 & ~x23 & ~x24 & ~x26 & ~x31 & ~x36 & ~x37 & ~x38 & ~x39 & ~x42 & ~x43 & ~x44 & ~x45 & ~x47 & ~x49 & ~x52 & ~x54 & ~x60 & ~x62 & ~x66 & ~x67 & ~x72 & ~x75 & ~x77 & ~x81 & ~x85 & ~x89 & ~x94 & ~x98 & ~x104 & ~x105 & ~x107 & ~x109 & ~x110 & ~x115 & ~x116 & ~x118 & ~x120 & ~x121 & ~x122 & ~x123 & ~x130 & ~x139 & ~x141 & ~x142 & ~x145 & ~x146 & ~x147 & ~x161 & ~x166 & ~x169 & ~x173 & ~x174 & ~x195 & ~x196 & ~x200 & ~x205 & ~x223 & ~x249 & ~x250 & ~x251 & ~x252 & ~x254 & ~x256 & ~x275 & ~x276 & ~x277 & ~x284 & ~x285 & ~x304 & ~x306 & ~x307 & ~x309 & ~x311 & ~x329 & ~x335 & ~x337 & ~x338 & ~x365 & ~x394 & ~x395 & ~x416 & ~x417 & ~x418 & ~x419 & ~x423 & ~x444 & ~x445 & ~x446 & ~x447 & ~x450 & ~x451 & ~x473 & ~x501 & ~x527 & ~x530 & ~x531 & ~x533 & ~x536 & ~x537 & ~x554 & ~x556 & ~x558 & ~x561 & ~x563 & ~x580 & ~x582 & ~x583 & ~x584 & ~x585 & ~x586 & ~x588 & ~x589 & ~x590 & ~x594 & ~x609 & ~x610 & ~x613 & ~x616 & ~x619 & ~x639 & ~x641 & ~x646 & ~x649 & ~x657 & ~x667 & ~x669 & ~x670 & ~x671 & ~x675 & ~x686 & ~x695 & ~x697 & ~x699 & ~x705 & ~x706 & ~x709 & ~x713 & ~x714 & ~x717 & ~x722 & ~x725 & ~x727 & ~x728 & ~x729 & ~x730 & ~x731 & ~x732 & ~x734 & ~x735 & ~x738 & ~x743 & ~x748 & ~x750 & ~x753 & ~x755 & ~x758 & ~x759 & ~x767 & ~x768 & ~x771 & ~x775 & ~x783;
assign c4270 =  x271 & ~x15 & ~x23 & ~x41 & ~x42 & ~x88 & ~x92 & ~x103 & ~x114 & ~x116 & ~x157 & ~x167 & ~x172 & ~x185 & ~x221 & ~x225 & ~x227 & ~x241 & ~x258 & ~x281 & ~x311 & ~x313 & ~x323 & ~x330 & ~x332 & ~x333 & ~x334 & ~x360 & ~x367 & ~x418 & ~x477 & ~x505 & ~x530 & ~x561 & ~x592 & ~x595 & ~x610 & ~x616 & ~x621 & ~x647 & ~x663 & ~x735 & ~x737 & ~x740 & ~x747 & ~x752 & ~x762 & ~x765;
assign c4272 =  x727;
assign c4274 =  x217 &  x299 &  x455 &  x483;
assign c4276 =  x758;
assign c4278 =  x289 &  x316 &  x317 &  x465 &  x493 &  x521 & ~x9 & ~x34 & ~x42 & ~x53 & ~x59 & ~x74 & ~x78 & ~x82 & ~x93 & ~x94 & ~x95 & ~x99 & ~x104 & ~x113 & ~x115 & ~x116 & ~x144 & ~x166 & ~x193 & ~x195 & ~x249 & ~x250 & ~x253 & ~x280 & ~x303 & ~x306 & ~x320 & ~x331 & ~x333 & ~x334 & ~x337 & ~x420 & ~x421 & ~x452 & ~x530 & ~x535 & ~x556 & ~x560 & ~x562 & ~x581 & ~x583 & ~x613 & ~x617 & ~x639 & ~x640 & ~x641 & ~x642 & ~x668 & ~x672 & ~x678 & ~x683 & ~x704 & ~x711 & ~x712 & ~x713 & ~x719 & ~x720 & ~x739 & ~x741 & ~x745 & ~x746 & ~x750 & ~x759 & ~x761 & ~x778;
assign c4280 =  x279;
assign c4282 =  x723;
assign c4284 =  x438 & ~x6 & ~x12 & ~x20 & ~x21 & ~x22 & ~x23 & ~x25 & ~x26 & ~x33 & ~x35 & ~x39 & ~x48 & ~x50 & ~x58 & ~x69 & ~x74 & ~x79 & ~x83 & ~x86 & ~x97 & ~x108 & ~x117 & ~x118 & ~x127 & ~x155 & ~x194 & ~x211 & ~x222 & ~x239 & ~x267 & ~x276 & ~x322 & ~x366 & ~x390 & ~x393 & ~x449 & ~x533 & ~x534 & ~x563 & ~x588 & ~x601 & ~x618 & ~x640 & ~x641 & ~x657 & ~x666 & ~x667 & ~x668 & ~x670 & ~x675 & ~x678 & ~x686 & ~x720 & ~x740 & ~x745 & ~x746 & ~x755 & ~x760 & ~x766 & ~x777;
assign c4286 =  x273 &  x356 &  x372 &  x428 & ~x186 & ~x213 & ~x267 & ~x387 & ~x388;
assign c4288 = ~x16 & ~x18 & ~x19 & ~x21 & ~x22 & ~x29 & ~x34 & ~x36 & ~x43 & ~x48 & ~x49 & ~x54 & ~x57 & ~x68 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x104 & ~x105 & ~x115 & ~x116 & ~x118 & ~x123 & ~x128 & ~x134 & ~x139 & ~x140 & ~x144 & ~x150 & ~x160 & ~x161 & ~x174 & ~x200 & ~x201 & ~x206 & ~x219 & ~x223 & ~x256 & ~x271 & ~x305 & ~x310 & ~x337 & ~x360 & ~x362 & ~x367 & ~x369 & ~x388 & ~x394 & ~x417 & ~x421 & ~x423 & ~x477 & ~x505 & ~x526 & ~x528 & ~x533 & ~x543 & ~x557 & ~x567 & ~x568 & ~x569 & ~x582 & ~x584 & ~x597 & ~x611 & ~x615 & ~x617 & ~x622 & ~x627 & ~x644 & ~x671 & ~x681 & ~x687 & ~x698 & ~x702 & ~x709 & ~x712 & ~x714 & ~x715 & ~x716 & ~x719 & ~x720 & ~x721 & ~x724 & ~x731 & ~x760 & ~x769 & ~x777 & ~x780 & ~x781;
assign c4290 =  x504;
assign c4292 =  x396;
assign c4294 = ~x0 & ~x15 & ~x18 & ~x22 & ~x26 & ~x27 & ~x28 & ~x32 & ~x33 & ~x35 & ~x63 & ~x65 & ~x72 & ~x85 & ~x86 & ~x95 & ~x98 & ~x103 & ~x106 & ~x107 & ~x117 & ~x119 & ~x124 & ~x137 & ~x139 & ~x144 & ~x160 & ~x164 & ~x180 & ~x189 & ~x196 & ~x200 & ~x208 & ~x221 & ~x235 & ~x253 & ~x272 & ~x274 & ~x278 & ~x283 & ~x303 & ~x307 & ~x312 & ~x329 & ~x331 & ~x333 & ~x337 & ~x359 & ~x362 & ~x365 & ~x389 & ~x390 & ~x394 & ~x396 & ~x397 & ~x444 & ~x448 & ~x450 & ~x454 & ~x475 & ~x476 & ~x477 & ~x506 & ~x525 & ~x532 & ~x537 & ~x585 & ~x592 & ~x599 & ~x615 & ~x618 & ~x645 & ~x652 & ~x654 & ~x657 & ~x667 & ~x671 & ~x673 & ~x674 & ~x675 & ~x679 & ~x697 & ~x701 & ~x704 & ~x705 & ~x712 & ~x713 & ~x724 & ~x725 & ~x753 & ~x755 & ~x759 & ~x763 & ~x765 & ~x766 & ~x772 & ~x778;
assign c4296 =  x399 &  x426 &  x466 &  x491 &  x493 & ~x2 & ~x5 & ~x22 & ~x28 & ~x37 & ~x54 & ~x62 & ~x66 & ~x71 & ~x78 & ~x96 & ~x98 & ~x116 & ~x117 & ~x137 & ~x168 & ~x194 & ~x197 & ~x202 & ~x277 & ~x336 & ~x339 & ~x445 & ~x446 & ~x477 & ~x503 & ~x530 & ~x582 & ~x594 & ~x598 & ~x616 & ~x620 & ~x622 & ~x640 & ~x642 & ~x644 & ~x651 & ~x669 & ~x673 & ~x676 & ~x693 & ~x697 & ~x707 & ~x709 & ~x711 & ~x725 & ~x732 & ~x735 & ~x737 & ~x747 & ~x760 & ~x761 & ~x766;
assign c4298 =  x403 &  x434 & ~x4 & ~x5 & ~x8 & ~x9 & ~x24 & ~x30 & ~x42 & ~x43 & ~x63 & ~x64 & ~x66 & ~x69 & ~x73 & ~x80 & ~x85 & ~x87 & ~x89 & ~x94 & ~x106 & ~x111 & ~x116 & ~x119 & ~x122 & ~x124 & ~x125 & ~x126 & ~x127 & ~x135 & ~x136 & ~x144 & ~x146 & ~x154 & ~x156 & ~x196 & ~x199 & ~x211 & ~x222 & ~x230 & ~x231 & ~x248 & ~x257 & ~x274 & ~x302 & ~x314 & ~x328 & ~x330 & ~x334 & ~x336 & ~x394 & ~x450 & ~x474 & ~x497 & ~x502 & ~x503 & ~x510 & ~x549 & ~x551 & ~x555 & ~x557 & ~x559 & ~x562 & ~x565 & ~x567 & ~x580 & ~x584 & ~x585 & ~x594 & ~x606 & ~x621 & ~x638 & ~x648 & ~x663 & ~x665 & ~x675 & ~x690 & ~x692 & ~x701 & ~x717 & ~x722 & ~x728 & ~x731 & ~x732 & ~x733 & ~x734 & ~x736 & ~x737 & ~x739 & ~x740 & ~x748 & ~x749 & ~x752 & ~x753 & ~x764 & ~x766 & ~x772 & ~x781 & ~x782;
assign c41 =  x545 & ~x7 & ~x8 & ~x12 & ~x14 & ~x17 & ~x19 & ~x22 & ~x23 & ~x24 & ~x25 & ~x26 & ~x32 & ~x35 & ~x55 & ~x56 & ~x58 & ~x60 & ~x83 & ~x85 & ~x86 & ~x89 & ~x108 & ~x115 & ~x116 & ~x118 & ~x139 & ~x142 & ~x144 & ~x145 & ~x146 & ~x162 & ~x163 & ~x165 & ~x167 & ~x168 & ~x169 & ~x171 & ~x192 & ~x193 & ~x195 & ~x219 & ~x220 & ~x223 & ~x224 & ~x225 & ~x226 & ~x248 & ~x250 & ~x255 & ~x270 & ~x280 & ~x306 & ~x307 & ~x308 & ~x311 & ~x334 & ~x335 & ~x339 & ~x363 & ~x364 & ~x368 & ~x395 & ~x420 & ~x421 & ~x448 & ~x449 & ~x450 & ~x475 & ~x505 & ~x506 & ~x530 & ~x587 & ~x589 & ~x612 & ~x614 & ~x618 & ~x627 & ~x629 & ~x630 & ~x632 & ~x633 & ~x635 & ~x636 & ~x638 & ~x645 & ~x648 & ~x652 & ~x658 & ~x661 & ~x665 & ~x672 & ~x676 & ~x683 & ~x685 & ~x690 & ~x692 & ~x694 & ~x697 & ~x699 & ~x712 & ~x713 & ~x726 & ~x728 & ~x735 & ~x737 & ~x738 & ~x742 & ~x748 & ~x749 & ~x755 & ~x760 & ~x761 & ~x762 & ~x764 & ~x765 & ~x770 & ~x772 & ~x773 & ~x776 & ~x780 & ~x783;
assign c43 =  x569 & ~x439 & ~x465;
assign c45 =  x122;
assign c47 =  x407 & ~x27 & ~x30 & ~x163 & ~x247 & ~x268 & ~x269 & ~x271 & ~x369 & ~x624 & ~x642 & ~x657 & ~x661 & ~x687 & ~x692;
assign c49 = ~x0 & ~x2 & ~x4 & ~x5 & ~x6 & ~x8 & ~x9 & ~x12 & ~x13 & ~x15 & ~x16 & ~x17 & ~x18 & ~x20 & ~x21 & ~x22 & ~x23 & ~x24 & ~x26 & ~x27 & ~x28 & ~x30 & ~x32 & ~x33 & ~x34 & ~x35 & ~x36 & ~x37 & ~x38 & ~x39 & ~x42 & ~x44 & ~x45 & ~x46 & ~x48 & ~x50 & ~x51 & ~x52 & ~x53 & ~x54 & ~x55 & ~x56 & ~x58 & ~x62 & ~x63 & ~x64 & ~x65 & ~x67 & ~x68 & ~x70 & ~x71 & ~x72 & ~x73 & ~x74 & ~x76 & ~x77 & ~x78 & ~x80 & ~x82 & ~x85 & ~x86 & ~x87 & ~x88 & ~x89 & ~x90 & ~x91 & ~x94 & ~x95 & ~x98 & ~x99 & ~x100 & ~x101 & ~x102 & ~x103 & ~x105 & ~x108 & ~x110 & ~x112 & ~x114 & ~x116 & ~x117 & ~x118 & ~x119 & ~x120 & ~x121 & ~x122 & ~x123 & ~x124 & ~x125 & ~x126 & ~x127 & ~x128 & ~x129 & ~x130 & ~x131 & ~x132 & ~x133 & ~x134 & ~x135 & ~x136 & ~x137 & ~x138 & ~x139 & ~x143 & ~x144 & ~x146 & ~x147 & ~x148 & ~x149 & ~x151 & ~x152 & ~x154 & ~x155 & ~x157 & ~x158 & ~x159 & ~x160 & ~x161 & ~x162 & ~x163 & ~x164 & ~x165 & ~x166 & ~x167 & ~x168 & ~x169 & ~x170 & ~x171 & ~x172 & ~x173 & ~x174 & ~x176 & ~x177 & ~x178 & ~x179 & ~x180 & ~x181 & ~x183 & ~x184 & ~x185 & ~x187 & ~x191 & ~x192 & ~x193 & ~x194 & ~x195 & ~x196 & ~x197 & ~x198 & ~x199 & ~x200 & ~x202 & ~x203 & ~x204 & ~x221 & ~x222 & ~x223 & ~x224 & ~x225 & ~x226 & ~x228 & ~x229 & ~x250 & ~x252 & ~x253 & ~x255 & ~x256 & ~x278 & ~x279 & ~x281 & ~x282 & ~x307 & ~x308 & ~x309 & ~x311 & ~x333 & ~x334 & ~x335 & ~x337 & ~x361 & ~x363 & ~x364 & ~x391 & ~x392 & ~x393 & ~x394 & ~x417 & ~x418 & ~x419 & ~x420 & ~x421 & ~x422 & ~x423 & ~x424 & ~x446 & ~x447 & ~x448 & ~x449 & ~x450 & ~x473 & ~x474 & ~x475 & ~x476 & ~x477 & ~x478 & ~x479 & ~x500 & ~x501 & ~x502 & ~x503 & ~x504 & ~x505 & ~x506 & ~x507 & ~x528 & ~x529 & ~x531 & ~x532 & ~x535 & ~x536 & ~x537 & ~x553 & ~x556 & ~x557 & ~x558 & ~x559 & ~x560 & ~x561 & ~x562 & ~x563 & ~x564 & ~x565 & ~x566 & ~x580 & ~x581 & ~x583 & ~x584 & ~x585 & ~x586 & ~x588 & ~x590 & ~x591 & ~x592 & ~x594 & ~x595 & ~x597 & ~x598 & ~x608 & ~x610 & ~x611 & ~x612 & ~x613 & ~x615 & ~x616 & ~x618 & ~x619 & ~x620 & ~x622 & ~x623 & ~x624 & ~x625 & ~x636 & ~x637 & ~x638 & ~x640 & ~x641 & ~x642 & ~x643 & ~x647 & ~x648 & ~x650 & ~x665 & ~x667 & ~x668 & ~x669 & ~x670 & ~x672 & ~x673 & ~x676 & ~x677 & ~x678 & ~x679 & ~x692 & ~x693 & ~x694 & ~x695 & ~x697 & ~x699 & ~x700 & ~x701 & ~x702 & ~x703 & ~x704 & ~x720 & ~x723 & ~x725 & ~x726 & ~x727 & ~x728 & ~x729 & ~x730 & ~x732 & ~x734 & ~x742 & ~x748 & ~x749 & ~x753 & ~x754 & ~x755 & ~x756 & ~x757 & ~x758 & ~x760 & ~x761 & ~x762 & ~x763 & ~x764 & ~x768 & ~x769 & ~x773 & ~x775 & ~x776 & ~x777 & ~x778 & ~x779 & ~x780 & ~x781 & ~x782 & ~x783;
assign c411 =  x238 &  x712;
assign c413 = ~x15 & ~x46 & ~x76 & ~x97 & ~x106 & ~x187 & ~x195 & ~x222 & ~x223 & ~x226 & ~x335 & ~x358 & ~x385 & ~x401 & ~x402 & ~x404 & ~x415 & ~x419 & ~x420 & ~x426 & ~x441 & ~x473 & ~x507 & ~x509 & ~x528 & ~x581 & ~x617 & ~x641 & ~x764 & ~x766 & ~x768;
assign c415 =  x600 &  x602 & ~x4 & ~x25 & ~x58 & ~x112 & ~x114 & ~x134 & ~x225 & ~x281 & ~x283 & ~x307 & ~x341 & ~x364 & ~x370 & ~x388 & ~x399 & ~x426 & ~x427 & ~x561 & ~x592 & ~x615 & ~x711 & ~x721 & ~x732 & ~x747 & ~x756 & ~x766;
assign c417 = ~x3 & ~x5 & ~x11 & ~x14 & ~x15 & ~x17 & ~x24 & ~x27 & ~x32 & ~x43 & ~x47 & ~x48 & ~x49 & ~x51 & ~x57 & ~x58 & ~x61 & ~x67 & ~x80 & ~x82 & ~x84 & ~x88 & ~x89 & ~x110 & ~x111 & ~x120 & ~x136 & ~x139 & ~x146 & ~x171 & ~x176 & ~x195 & ~x197 & ~x199 & ~x205 & ~x252 & ~x256 & ~x279 & ~x307 & ~x309 & ~x338 & ~x340 & ~x341 & ~x342 & ~x361 & ~x365 & ~x389 & ~x391 & ~x393 & ~x395 & ~x409 & ~x415 & ~x437 & ~x465 & ~x471 & ~x476 & ~x501 & ~x504 & ~x527 & ~x532 & ~x533 & ~x535 & ~x553 & ~x560 & ~x581 & ~x586 & ~x587 & ~x590 & ~x591 & ~x607 & ~x610 & ~x612 & ~x613 & ~x617 & ~x635 & ~x637 & ~x642 & ~x647 & ~x664 & ~x665 & ~x671 & ~x673 & ~x674 & ~x677 & ~x692 & ~x694 & ~x701 & ~x708 & ~x709 & ~x710 & ~x712 & ~x714 & ~x716 & ~x717 & ~x718 & ~x722 & ~x724 & ~x725 & ~x726 & ~x727 & ~x731 & ~x736 & ~x741 & ~x743 & ~x748 & ~x749 & ~x753 & ~x759 & ~x762 & ~x763 & ~x767 & ~x768 & ~x769 & ~x771 & ~x772 & ~x773 & ~x778 & ~x779 & ~x780 & ~x782 & ~x783;
assign c419 = ~x24 & ~x31 & ~x34 & ~x38 & ~x40 & ~x43 & ~x44 & ~x59 & ~x73 & ~x74 & ~x79 & ~x85 & ~x96 & ~x97 & ~x103 & ~x104 & ~x105 & ~x106 & ~x111 & ~x114 & ~x117 & ~x142 & ~x143 & ~x150 & ~x166 & ~x167 & ~x168 & ~x173 & ~x177 & ~x192 & ~x194 & ~x199 & ~x219 & ~x222 & ~x249 & ~x251 & ~x255 & ~x307 & ~x338 & ~x361 & ~x374 & ~x393 & ~x402 & ~x403 & ~x444 & ~x451 & ~x456 & ~x506 & ~x533 & ~x537 & ~x562 & ~x581 & ~x591 & ~x608 & ~x621 & ~x622 & ~x639 & ~x647 & ~x672 & ~x675 & ~x677 & ~x679 & ~x698 & ~x699 & ~x700 & ~x707 & ~x736 & ~x740 & ~x752 & ~x766 & ~x770 & ~x774 & ~x775 & ~x777 & ~x783;
assign c421 =  x572 &  x575 & ~x4 & ~x17 & ~x89 & ~x145 & ~x160 & ~x214 & ~x273 & ~x657 & ~x690 & ~x702 & ~x711 & ~x736;
assign c423 =  x235 &  x236 &  x238 & ~x346;
assign c425 =  x206 &  x208 & ~x15 & ~x25 & ~x31 & ~x37 & ~x71 & ~x81 & ~x123 & ~x136 & ~x161 & ~x168 & ~x219 & ~x220 & ~x274 & ~x282 & ~x308 & ~x311 & ~x362 & ~x422 & ~x535 & ~x560 & ~x563 & ~x671 & ~x672 & ~x696 & ~x703 & ~x707 & ~x725 & ~x733 & ~x736 & ~x781;
assign c427 = ~x4 & ~x7 & ~x8 & ~x27 & ~x29 & ~x36 & ~x46 & ~x78 & ~x88 & ~x90 & ~x91 & ~x132 & ~x136 & ~x156 & ~x158 & ~x175 & ~x184 & ~x197 & ~x281 & ~x364 & ~x365 & ~x379 & ~x389 & ~x390 & ~x406 & ~x431 & ~x432 & ~x445 & ~x447 & ~x449 & ~x451 & ~x460 & ~x487 & ~x511 & ~x514 & ~x527 & ~x589 & ~x593 & ~x595 & ~x644 & ~x699 & ~x701 & ~x759 & ~x763 & ~x765 & ~x777 & ~x780;
assign c429 =  x570 &  x599 & ~x217 & ~x624;
assign c431 =  x236 &  x237 &  x238 & ~x4 & ~x18 & ~x38 & ~x41 & ~x45 & ~x50 & ~x53 & ~x67 & ~x68 & ~x88 & ~x91 & ~x97 & ~x103 & ~x119 & ~x122 & ~x125 & ~x137 & ~x142 & ~x170 & ~x221 & ~x223 & ~x229 & ~x257 & ~x284 & ~x305 & ~x307 & ~x331 & ~x340 & ~x356 & ~x362 & ~x393 & ~x411 & ~x419 & ~x420 & ~x421 & ~x422 & ~x427 & ~x439 & ~x468 & ~x477 & ~x483 & ~x497 & ~x503 & ~x523 & ~x553 & ~x561 & ~x579 & ~x586 & ~x591 & ~x595 & ~x607 & ~x610 & ~x616 & ~x621 & ~x623 & ~x639 & ~x644 & ~x645 & ~x665 & ~x667 & ~x728 & ~x753 & ~x758 & ~x772 & ~x774 & ~x778;
assign c433 = ~x11 & ~x22 & ~x51 & ~x54 & ~x77 & ~x106 & ~x133 & ~x135 & ~x136 & ~x169 & ~x171 & ~x179 & ~x180 & ~x195 & ~x197 & ~x219 & ~x226 & ~x227 & ~x279 & ~x348 & ~x366 & ~x398 & ~x427 & ~x450 & ~x451 & ~x502 & ~x647 & ~x663 & ~x693 & ~x713 & ~x729 & ~x741 & ~x751;
assign c435 = ~x11 & ~x19 & ~x24 & ~x51 & ~x111 & ~x167 & ~x168 & ~x171 & ~x172 & ~x222 & ~x257 & ~x279 & ~x286 & ~x313 & ~x337 & ~x341 & ~x348 & ~x357 & ~x399 & ~x400 & ~x470 & ~x500 & ~x559 & ~x561 & ~x578 & ~x580 & ~x668 & ~x687 & ~x704 & ~x715 & ~x720 & ~x746 & ~x775 & ~x777;
assign c437 =  x268 &  x327 & ~x78 & ~x181 & ~x258 & ~x369 & ~x423 & ~x526 & ~x531 & ~x618 & ~x637 & ~x642 & ~x651;
assign c439 =  x209 &  x211 &  x236 & ~x399 & ~x467 & ~x502;
assign c441 =  x524 & ~x0 & ~x247 & ~x248 & ~x297 & ~x299 & ~x425 & ~x452 & ~x533 & ~x615 & ~x746 & ~x754;
assign c443 =  x213 &  x214 &  x238 &  x328 & ~x47 & ~x86 & ~x113 & ~x121 & ~x152 & ~x180 & ~x504 & ~x733;
assign c445 =  x154 &  x179 & ~x135 & ~x219;
assign c447 =  x573 &  x575 & ~x48 & ~x52 & ~x86 & ~x166 & ~x169 & ~x189 & ~x191 & ~x192 & ~x269 & ~x270 & ~x275 & ~x278 & ~x390 & ~x533 & ~x634 & ~x655 & ~x668 & ~x670 & ~x691 & ~x704 & ~x734 & ~x762 & ~x771 & ~x782;
assign c449 =  x184 &  x185 & ~x267 & ~x268 & ~x269 & ~x293;
assign c451 =  x602 &  x624;
assign c453 =  x623 & ~x678;
assign c455 = ~x6 & ~x12 & ~x18 & ~x35 & ~x49 & ~x58 & ~x72 & ~x88 & ~x126 & ~x165 & ~x172 & ~x225 & ~x227 & ~x229 & ~x252 & ~x280 & ~x334 & ~x335 & ~x346 & ~x366 & ~x385 & ~x413 & ~x464 & ~x504 & ~x618 & ~x665 & ~x672 & ~x683 & ~x698 & ~x701 & ~x705 & ~x716 & ~x721 & ~x724 & ~x727 & ~x730 & ~x733 & ~x737 & ~x749 & ~x750 & ~x755 & ~x763 & ~x764;
assign c457 = ~x8 & ~x21 & ~x23 & ~x30 & ~x39 & ~x41 & ~x49 & ~x50 & ~x53 & ~x61 & ~x75 & ~x86 & ~x91 & ~x105 & ~x115 & ~x124 & ~x125 & ~x127 & ~x144 & ~x170 & ~x174 & ~x218 & ~x283 & ~x333 & ~x336 & ~x347 & ~x348 & ~x376 & ~x421 & ~x422 & ~x440 & ~x443 & ~x453 & ~x477 & ~x495 & ~x496 & ~x533 & ~x615 & ~x624 & ~x646 & ~x649 & ~x692 & ~x698 & ~x703 & ~x747 & ~x749 & ~x776 & ~x781;
assign c459 =  x209 &  x210 &  x211 & ~x18 & ~x20 & ~x28 & ~x30 & ~x38 & ~x46 & ~x47 & ~x53 & ~x70 & ~x114 & ~x140 & ~x153 & ~x172 & ~x227 & ~x246 & ~x252 & ~x275 & ~x276 & ~x313 & ~x330 & ~x335 & ~x364 & ~x368 & ~x369 & ~x387 & ~x391 & ~x392 & ~x393 & ~x395 & ~x397 & ~x413 & ~x414 & ~x415 & ~x440 & ~x441 & ~x448 & ~x454 & ~x482 & ~x496 & ~x499 & ~x504 & ~x511 & ~x558 & ~x583 & ~x596 & ~x614 & ~x669 & ~x680 & ~x702 & ~x708 & ~x710 & ~x762 & ~x763 & ~x774 & ~x775 & ~x779 & ~x781;
assign c461 =  x294 & ~x0 & ~x2 & ~x7 & ~x14 & ~x17 & ~x20 & ~x22 & ~x24 & ~x26 & ~x31 & ~x34 & ~x35 & ~x39 & ~x42 & ~x47 & ~x54 & ~x61 & ~x62 & ~x65 & ~x67 & ~x70 & ~x73 & ~x74 & ~x76 & ~x78 & ~x79 & ~x81 & ~x82 & ~x83 & ~x87 & ~x89 & ~x91 & ~x93 & ~x94 & ~x100 & ~x102 & ~x106 & ~x108 & ~x111 & ~x112 & ~x117 & ~x120 & ~x122 & ~x123 & ~x127 & ~x134 & ~x140 & ~x154 & ~x158 & ~x160 & ~x162 & ~x164 & ~x172 & ~x182 & ~x183 & ~x184 & ~x186 & ~x192 & ~x194 & ~x211 & ~x212 & ~x213 & ~x223 & ~x253 & ~x281 & ~x307 & ~x331 & ~x333 & ~x335 & ~x362 & ~x390 & ~x419 & ~x422 & ~x423 & ~x449 & ~x450 & ~x474 & ~x477 & ~x478 & ~x504 & ~x508 & ~x529 & ~x564 & ~x565 & ~x588 & ~x595 & ~x609 & ~x616 & ~x638 & ~x640 & ~x642 & ~x645 & ~x647 & ~x651 & ~x665 & ~x667 & ~x668 & ~x669 & ~x672 & ~x673 & ~x674 & ~x692 & ~x696 & ~x699 & ~x702 & ~x705 & ~x751 & ~x752 & ~x755 & ~x756 & ~x758 & ~x759 & ~x761 & ~x764 & ~x775 & ~x778 & ~x779 & ~x782;
assign c463 = ~x4 & ~x18 & ~x31 & ~x33 & ~x52 & ~x115 & ~x192 & ~x228 & ~x265 & ~x294 & ~x322 & ~x335 & ~x344 & ~x369 & ~x373 & ~x389 & ~x398 & ~x530 & ~x646 & ~x716;
assign c465 =  x155 & ~x237 & ~x267;
assign c467 = ~x13 & ~x15 & ~x16 & ~x24 & ~x33 & ~x36 & ~x46 & ~x60 & ~x65 & ~x70 & ~x76 & ~x81 & ~x82 & ~x92 & ~x101 & ~x113 & ~x115 & ~x136 & ~x168 & ~x197 & ~x199 & ~x223 & ~x282 & ~x308 & ~x310 & ~x338 & ~x353 & ~x355 & ~x365 & ~x380 & ~x383 & ~x389 & ~x412 & ~x423 & ~x440 & ~x447 & ~x448 & ~x480 & ~x503 & ~x536 & ~x559 & ~x611 & ~x617 & ~x619 & ~x620 & ~x639 & ~x672 & ~x673 & ~x692 & ~x722 & ~x726 & ~x728 & ~x773 & ~x778 & ~x779 & ~x781;
assign c469 =  x602 & ~x10 & ~x70 & ~x118 & ~x202 & ~x224 & ~x306 & ~x312 & ~x394 & ~x420 & ~x463 & ~x473 & ~x503 & ~x530 & ~x691 & ~x699 & ~x706 & ~x724 & ~x731 & ~x746;
assign c471 =  x714 &  x742;
assign c473 = ~x20 & ~x21 & ~x28 & ~x48 & ~x49 & ~x51 & ~x63 & ~x87 & ~x91 & ~x106 & ~x143 & ~x163 & ~x192 & ~x222 & ~x227 & ~x309 & ~x368 & ~x385 & ~x392 & ~x412 & ~x422 & ~x462 & ~x491 & ~x504 & ~x585 & ~x586 & ~x640 & ~x643 & ~x674 & ~x705 & ~x707 & ~x726 & ~x759 & ~x760 & ~x763;
assign c475 =  x236 & ~x8 & ~x60 & ~x76 & ~x101 & ~x106 & ~x113 & ~x129 & ~x165 & ~x167 & ~x188 & ~x217 & ~x257 & ~x274 & ~x275 & ~x284 & ~x313 & ~x375 & ~x414 & ~x417 & ~x423 & ~x471 & ~x482 & ~x511 & ~x542 & ~x563 & ~x570 & ~x593 & ~x677 & ~x763 & ~x775;
assign c477 =  x209 & ~x8 & ~x15 & ~x61 & ~x86 & ~x100 & ~x117 & ~x152 & ~x166 & ~x197 & ~x247 & ~x293 & ~x320 & ~x358 & ~x419 & ~x443 & ~x483 & ~x504 & ~x591 & ~x618 & ~x723 & ~x732;
assign c479 =  x178 & ~x274 & ~x346;
assign c481 =  x568 & ~x31 & ~x120 & ~x143 & ~x362 & ~x420 & ~x474 & ~x577 & ~x603 & ~x608 & ~x633 & ~x634 & ~x663 & ~x720 & ~x722;
assign c483 =  x188 & ~x297 & ~x298 & ~x314 & ~x496;
assign c485 =  x567 &  x597 & ~x1 & ~x34 & ~x53 & ~x138 & ~x167 & ~x204 & ~x232 & ~x340 & ~x528 & ~x532 & ~x563 & ~x664 & ~x665 & ~x674 & ~x681 & ~x712 & ~x744 & ~x745 & ~x750;
assign c487 =  x206 &  x208 &  x210 & ~x46 & ~x77 & ~x188 & ~x684;
assign c489 =  x262 & ~x76 & ~x101 & ~x248 & ~x274 & ~x401;
assign c491 = ~x32 & ~x56 & ~x70 & ~x100 & ~x101 & ~x140 & ~x191 & ~x197 & ~x364 & ~x371 & ~x399 & ~x408 & ~x419 & ~x428 & ~x504 & ~x639 & ~x641 & ~x702 & ~x730 & ~x762;
assign c493 =  x266 &  x546 &  x601 & ~x17 & ~x46 & ~x116 & ~x138 & ~x229 & ~x357 & ~x387 & ~x391 & ~x427 & ~x454 & ~x469 & ~x479 & ~x496 & ~x587 & ~x608;
assign c495 =  x577 &  x601 & ~x35 & ~x199 & ~x686;
assign c497 =  x181 &  x205;
assign c499 =  x580 &  x633;
assign c4101 =  x540 & ~x22 & ~x111 & ~x143 & ~x162 & ~x164 & ~x578 & ~x579 & ~x588 & ~x604 & ~x610 & ~x611 & ~x631 & ~x632 & ~x634 & ~x642 & ~x662 & ~x664 & ~x666 & ~x674 & ~x729 & ~x752 & ~x759 & ~x777;
assign c4103 =  x293 &  x294 &  x296 & ~x6 & ~x27 & ~x103 & ~x106 & ~x110 & ~x115 & ~x132 & ~x156 & ~x160 & ~x164 & ~x183 & ~x184 & ~x192 & ~x211 & ~x460 & ~x472 & ~x499 & ~x610;
assign c4105 = ~x0 & ~x2 & ~x7 & ~x22 & ~x27 & ~x28 & ~x33 & ~x54 & ~x80 & ~x86 & ~x94 & ~x98 & ~x118 & ~x141 & ~x144 & ~x194 & ~x198 & ~x199 & ~x200 & ~x203 & ~x224 & ~x250 & ~x379 & ~x380 & ~x382 & ~x383 & ~x419 & ~x421 & ~x422 & ~x473 & ~x477 & ~x502 & ~x507 & ~x532 & ~x533 & ~x560 & ~x643 & ~x698 & ~x729 & ~x742 & ~x765 & ~x770;
assign c4107 = ~x23 & ~x32 & ~x50 & ~x70 & ~x92 & ~x97 & ~x100 & ~x106 & ~x110 & ~x112 & ~x117 & ~x123 & ~x124 & ~x134 & ~x141 & ~x144 & ~x151 & ~x154 & ~x156 & ~x162 & ~x164 & ~x165 & ~x166 & ~x169 & ~x170 & ~x195 & ~x202 & ~x226 & ~x251 & ~x307 & ~x337 & ~x360 & ~x376 & ~x390 & ~x397 & ~x422 & ~x429 & ~x446 & ~x448 & ~x451 & ~x472 & ~x480 & ~x531 & ~x536 & ~x588 & ~x620 & ~x641 & ~x663 & ~x675 & ~x699 & ~x702 & ~x704 & ~x706 & ~x725 & ~x728 & ~x752 & ~x765 & ~x770;
assign c4109 =  x264 &  x288 &  x294 & ~x45 & ~x55 & ~x80 & ~x96 & ~x117 & ~x130 & ~x139 & ~x154 & ~x222 & ~x389 & ~x588 & ~x700 & ~x732;
assign c4111 =  x578 &  x601 & ~x391 & ~x395 & ~x452 & ~x561 & ~x697;
assign c4113 =  x239 &  x240 &  x270 & ~x8 & ~x11 & ~x16 & ~x20 & ~x26 & ~x29 & ~x34 & ~x35 & ~x39 & ~x41 & ~x42 & ~x46 & ~x47 & ~x49 & ~x52 & ~x56 & ~x64 & ~x68 & ~x77 & ~x83 & ~x85 & ~x87 & ~x97 & ~x100 & ~x105 & ~x106 & ~x120 & ~x124 & ~x127 & ~x130 & ~x135 & ~x137 & ~x139 & ~x140 & ~x141 & ~x148 & ~x151 & ~x155 & ~x157 & ~x174 & ~x176 & ~x194 & ~x197 & ~x198 & ~x201 & ~x224 & ~x225 & ~x230 & ~x231 & ~x254 & ~x256 & ~x259 & ~x277 & ~x278 & ~x280 & ~x283 & ~x284 & ~x309 & ~x311 & ~x360 & ~x361 & ~x368 & ~x369 & ~x387 & ~x388 & ~x394 & ~x397 & ~x414 & ~x420 & ~x421 & ~x424 & ~x425 & ~x445 & ~x454 & ~x473 & ~x505 & ~x526 & ~x534 & ~x555 & ~x559 & ~x562 & ~x563 & ~x583 & ~x585 & ~x586 & ~x610 & ~x612 & ~x619 & ~x639 & ~x641 & ~x644 & ~x668 & ~x671 & ~x698 & ~x700 & ~x701 & ~x702 & ~x727 & ~x731 & ~x733 & ~x754 & ~x758 & ~x760 & ~x766 & ~x768 & ~x771 & ~x773 & ~x774 & ~x777 & ~x778 & ~x782;
assign c4115 =  x179 &  x182 & ~x291;
assign c4117 =  x181 &  x182 & ~x292 & ~x293 & ~x397 & ~x468 & ~x562 & ~x777;
assign c4119 =  x739;
assign c4121 =  x40;
assign c4123 =  x261 &  x264 & ~x6 & ~x13 & ~x14 & ~x58 & ~x62 & ~x69 & ~x74 & ~x96 & ~x109 & ~x115 & ~x130 & ~x134 & ~x181 & ~x532 & ~x587 & ~x678 & ~x681 & ~x730 & ~x749 & ~x772;
assign c4125 = ~x0 & ~x1 & ~x6 & ~x8 & ~x10 & ~x15 & ~x19 & ~x21 & ~x28 & ~x30 & ~x44 & ~x46 & ~x52 & ~x59 & ~x62 & ~x64 & ~x76 & ~x82 & ~x85 & ~x88 & ~x110 & ~x112 & ~x113 & ~x115 & ~x116 & ~x132 & ~x133 & ~x136 & ~x137 & ~x140 & ~x142 & ~x166 & ~x167 & ~x173 & ~x189 & ~x190 & ~x196 & ~x199 & ~x200 & ~x216 & ~x217 & ~x219 & ~x221 & ~x222 & ~x227 & ~x243 & ~x250 & ~x269 & ~x271 & ~x272 & ~x273 & ~x274 & ~x275 & ~x276 & ~x280 & ~x281 & ~x284 & ~x295 & ~x299 & ~x300 & ~x302 & ~x306 & ~x310 & ~x329 & ~x333 & ~x339 & ~x360 & ~x367 & ~x392 & ~x393 & ~x398 & ~x423 & ~x424 & ~x450 & ~x452 & ~x453 & ~x477 & ~x480 & ~x503 & ~x507 & ~x531 & ~x533 & ~x536 & ~x537 & ~x563 & ~x565 & ~x566 & ~x567 & ~x585 & ~x591 & ~x612 & ~x613 & ~x614 & ~x617 & ~x622 & ~x639 & ~x642 & ~x651 & ~x665 & ~x669 & ~x674 & ~x676 & ~x677 & ~x681 & ~x682 & ~x685 & ~x696 & ~x699 & ~x704 & ~x710 & ~x711 & ~x717 & ~x725 & ~x727 & ~x731 & ~x733 & ~x738 & ~x749 & ~x752 & ~x755 & ~x758 & ~x759 & ~x760 & ~x761 & ~x764 & ~x768 & ~x769 & ~x772 & ~x773 & ~x775;
assign c4127 =  x209 &  x212 &  x409 & ~x347 & ~x442 & ~x478;
assign c4129 = ~x2 & ~x3 & ~x7 & ~x13 & ~x15 & ~x17 & ~x19 & ~x20 & ~x21 & ~x24 & ~x25 & ~x27 & ~x33 & ~x36 & ~x39 & ~x44 & ~x51 & ~x53 & ~x54 & ~x60 & ~x61 & ~x63 & ~x81 & ~x82 & ~x83 & ~x85 & ~x87 & ~x89 & ~x110 & ~x114 & ~x134 & ~x147 & ~x166 & ~x168 & ~x189 & ~x196 & ~x221 & ~x222 & ~x223 & ~x226 & ~x248 & ~x250 & ~x271 & ~x272 & ~x273 & ~x275 & ~x279 & ~x296 & ~x297 & ~x298 & ~x300 & ~x305 & ~x306 & ~x309 & ~x334 & ~x337 & ~x365 & ~x390 & ~x394 & ~x395 & ~x420 & ~x447 & ~x448 & ~x477 & ~x478 & ~x479 & ~x502 & ~x530 & ~x559 & ~x583 & ~x584 & ~x585 & ~x586 & ~x588 & ~x591 & ~x609 & ~x612 & ~x613 & ~x614 & ~x618 & ~x620 & ~x635 & ~x641 & ~x643 & ~x649 & ~x655 & ~x656 & ~x659 & ~x663 & ~x673 & ~x675 & ~x676 & ~x680 & ~x683 & ~x684 & ~x685 & ~x686 & ~x687 & ~x690 & ~x693 & ~x694 & ~x695 & ~x698 & ~x699 & ~x702 & ~x707 & ~x711 & ~x712 & ~x716 & ~x725 & ~x726 & ~x728 & ~x731 & ~x732 & ~x737 & ~x742 & ~x743 & ~x747 & ~x755 & ~x757 & ~x758 & ~x759 & ~x764 & ~x765 & ~x766 & ~x769 & ~x770 & ~x771 & ~x772 & ~x773 & ~x775 & ~x777 & ~x780 & ~x781;
assign c4131 =  x574 &  x600 & ~x381;
assign c4133 =  x122;
assign c4135 =  x178 &  x181;
assign c4137 =  x182 &  x206;
assign c4139 = ~x49 & ~x99 & ~x143 & ~x310 & ~x435 & ~x464 & ~x465 & ~x492 & ~x616 & ~x637 & ~x645 & ~x711 & ~x729 & ~x782;
assign c4141 = ~x52 & ~x67 & ~x99 & ~x164 & ~x198 & ~x254 & ~x295 & ~x335 & ~x367 & ~x369 & ~x393 & ~x394 & ~x414 & ~x421 & ~x425 & ~x456 & ~x467 & ~x513 & ~x523 & ~x560 & ~x614 & ~x647 & ~x701 & ~x732 & ~x747 & ~x762;
assign c4143 = ~x9 & ~x11 & ~x12 & ~x29 & ~x57 & ~x66 & ~x69 & ~x84 & ~x117 & ~x141 & ~x171 & ~x174 & ~x196 & ~x201 & ~x225 & ~x253 & ~x255 & ~x309 & ~x336 & ~x340 & ~x342 & ~x352 & ~x355 & ~x366 & ~x369 & ~x380 & ~x381 & ~x384 & ~x448 & ~x450 & ~x503 & ~x559 & ~x561 & ~x589 & ~x642 & ~x648 & ~x675 & ~x692 & ~x707 & ~x708 & ~x717 & ~x724 & ~x726 & ~x745 & ~x771;
assign c4145 =  x207 &  x211;
assign c4147 =  x266 & ~x76 & ~x436 & ~x646;
assign c4149 =  x571 & ~x22 & ~x50 & ~x139 & ~x217 & ~x218 & ~x246 & ~x276 & ~x297 & ~x305 & ~x340 & ~x508 & ~x531 & ~x560 & ~x652 & ~x674 & ~x683 & ~x703;
assign c4151 =  x543 &  x545 & ~x16 & ~x24 & ~x25 & ~x28 & ~x33 & ~x37 & ~x50 & ~x51 & ~x134 & ~x142 & ~x143 & ~x166 & ~x171 & ~x190 & ~x195 & ~x215 & ~x250 & ~x254 & ~x277 & ~x284 & ~x311 & ~x340 & ~x363 & ~x365 & ~x392 & ~x423 & ~x450 & ~x532 & ~x536 & ~x558 & ~x559 & ~x588 & ~x591 & ~x610 & ~x616 & ~x630 & ~x633 & ~x635 & ~x653 & ~x655 & ~x659 & ~x661 & ~x664 & ~x681 & ~x684 & ~x685 & ~x687 & ~x702 & ~x713 & ~x722 & ~x726 & ~x739 & ~x746 & ~x748 & ~x774 & ~x783;
assign c4153 =  x269 &  x293 & ~x12 & ~x14 & ~x50 & ~x80 & ~x107 & ~x116 & ~x154 & ~x161 & ~x173 & ~x183 & ~x186 & ~x194 & ~x252 & ~x388 & ~x470 & ~x474 & ~x488 & ~x534 & ~x585 & ~x588 & ~x673 & ~x697 & ~x724 & ~x758 & ~x783;
assign c4155 =  x241 &  x242 &  x266 & ~x0 & ~x4 & ~x5 & ~x7 & ~x9 & ~x10 & ~x14 & ~x16 & ~x18 & ~x19 & ~x27 & ~x29 & ~x30 & ~x31 & ~x33 & ~x34 & ~x36 & ~x41 & ~x54 & ~x55 & ~x61 & ~x64 & ~x65 & ~x66 & ~x67 & ~x70 & ~x71 & ~x77 & ~x78 & ~x81 & ~x84 & ~x85 & ~x89 & ~x97 & ~x102 & ~x107 & ~x109 & ~x110 & ~x112 & ~x114 & ~x115 & ~x117 & ~x119 & ~x121 & ~x122 & ~x123 & ~x125 & ~x127 & ~x138 & ~x139 & ~x143 & ~x144 & ~x147 & ~x149 & ~x151 & ~x153 & ~x154 & ~x155 & ~x156 & ~x164 & ~x175 & ~x176 & ~x177 & ~x178 & ~x179 & ~x180 & ~x181 & ~x195 & ~x196 & ~x197 & ~x200 & ~x224 & ~x226 & ~x227 & ~x256 & ~x277 & ~x278 & ~x283 & ~x285 & ~x304 & ~x307 & ~x311 & ~x333 & ~x341 & ~x359 & ~x361 & ~x362 & ~x363 & ~x364 & ~x365 & ~x388 & ~x389 & ~x394 & ~x395 & ~x415 & ~x416 & ~x418 & ~x420 & ~x423 & ~x424 & ~x441 & ~x442 & ~x452 & ~x453 & ~x468 & ~x469 & ~x470 & ~x471 & ~x472 & ~x476 & ~x478 & ~x479 & ~x480 & ~x481 & ~x495 & ~x496 & ~x498 & ~x501 & ~x502 & ~x504 & ~x506 & ~x510 & ~x524 & ~x528 & ~x529 & ~x532 & ~x555 & ~x557 & ~x559 & ~x560 & ~x579 & ~x580 & ~x583 & ~x587 & ~x607 & ~x610 & ~x634 & ~x635 & ~x639 & ~x640 & ~x642 & ~x644 & ~x648 & ~x664 & ~x674 & ~x692 & ~x693 & ~x699 & ~x701 & ~x704 & ~x705 & ~x718 & ~x719 & ~x723 & ~x725 & ~x728 & ~x729 & ~x731 & ~x733 & ~x742 & ~x743 & ~x745 & ~x746 & ~x757 & ~x758 & ~x767 & ~x771 & ~x773 & ~x778 & ~x780 & ~x781 & ~x782;
assign c4157 = ~x0 & ~x7 & ~x10 & ~x24 & ~x31 & ~x34 & ~x35 & ~x40 & ~x45 & ~x64 & ~x76 & ~x82 & ~x95 & ~x109 & ~x112 & ~x120 & ~x139 & ~x141 & ~x144 & ~x145 & ~x170 & ~x194 & ~x251 & ~x280 & ~x376 & ~x400 & ~x401 & ~x403 & ~x418 & ~x423 & ~x427 & ~x533 & ~x534 & ~x614 & ~x615 & ~x637 & ~x642 & ~x645 & ~x646 & ~x672 & ~x676 & ~x691 & ~x701 & ~x705 & ~x706 & ~x721 & ~x722 & ~x724 & ~x725 & ~x749 & ~x758 & ~x760 & ~x763 & ~x767 & ~x772 & ~x779 & ~x783;
assign c4159 =  x97 &  x544 &  x574;
assign c4161 =  x240 &  x243 & ~x20 & ~x26 & ~x34 & ~x57 & ~x60 & ~x72 & ~x73 & ~x84 & ~x107 & ~x112 & ~x132 & ~x134 & ~x147 & ~x179 & ~x202 & ~x282 & ~x336 & ~x363 & ~x420 & ~x422 & ~x453 & ~x468 & ~x470 & ~x479 & ~x481 & ~x497 & ~x504 & ~x523 & ~x524 & ~x525 & ~x557 & ~x578 & ~x580 & ~x582 & ~x636 & ~x644 & ~x676 & ~x695 & ~x698 & ~x728 & ~x740 & ~x752 & ~x765 & ~x775;
assign c4163 =  x212 &  x214 & ~x7 & ~x10 & ~x15 & ~x16 & ~x17 & ~x19 & ~x33 & ~x34 & ~x44 & ~x63 & ~x64 & ~x85 & ~x91 & ~x95 & ~x109 & ~x111 & ~x125 & ~x140 & ~x146 & ~x150 & ~x174 & ~x177 & ~x178 & ~x179 & ~x221 & ~x222 & ~x224 & ~x233 & ~x280 & ~x307 & ~x308 & ~x314 & ~x335 & ~x341 & ~x361 & ~x413 & ~x420 & ~x424 & ~x445 & ~x446 & ~x467 & ~x475 & ~x477 & ~x495 & ~x524 & ~x529 & ~x532 & ~x535 & ~x550 & ~x551 & ~x553 & ~x557 & ~x558 & ~x560 & ~x563 & ~x564 & ~x567 & ~x585 & ~x586 & ~x590 & ~x617 & ~x638 & ~x643 & ~x644 & ~x661 & ~x665 & ~x672 & ~x692 & ~x693 & ~x700 & ~x704 & ~x722 & ~x724 & ~x725 & ~x731 & ~x733 & ~x748 & ~x753 & ~x766 & ~x770 & ~x774;
assign c4165 =  x209 &  x211 &  x212 & ~x1 & ~x14 & ~x31 & ~x85 & ~x120 & ~x142 & ~x321 & ~x387 & ~x399 & ~x474 & ~x588 & ~x780 & ~x783;
assign c4167 =  x656 & ~x22 & ~x30 & ~x31 & ~x116 & ~x140 & ~x442 & ~x476 & ~x479 & ~x534 & ~x545 & ~x573;
assign c4169 =  x235 &  x236 & ~x32 & ~x79 & ~x179 & ~x386 & ~x495 & ~x496 & ~x497 & ~x663 & ~x722 & ~x733;
assign c4171 =  x235 &  x238 &  x261 &  x262 & ~x32 & ~x75 & ~x107 & ~x109 & ~x148 & ~x218 & ~x219 & ~x221 & ~x246 & ~x248 & ~x364 & ~x444 & ~x451 & ~x504 & ~x506 & ~x559 & ~x560 & ~x561 & ~x585 & ~x671 & ~x758;
assign c4173 =  x569 & ~x26 & ~x106 & ~x135 & ~x177 & ~x260 & ~x364 & ~x389 & ~x443 & ~x444 & ~x605 & ~x639 & ~x652 & ~x672 & ~x745 & ~x746 & ~x773;
assign c4175 = ~x19 & ~x74 & ~x79 & ~x87 & ~x105 & ~x112 & ~x144 & ~x146 & ~x169 & ~x264 & ~x305 & ~x333 & ~x336 & ~x338 & ~x361 & ~x402 & ~x416 & ~x418 & ~x427 & ~x429 & ~x430 & ~x440 & ~x449 & ~x502 & ~x530 & ~x556 & ~x618 & ~x619 & ~x636 & ~x645 & ~x695 & ~x699 & ~x716 & ~x727 & ~x738;
assign c4177 =  x238 & ~x36 & ~x58 & ~x93 & ~x165 & ~x318 & ~x320 & ~x559;
assign c4179 =  x566 &  x625;
assign c4181 =  x237 &  x239 &  x240 &  x241 &  x242 & ~x1 & ~x3 & ~x4 & ~x6 & ~x8 & ~x15 & ~x16 & ~x21 & ~x34 & ~x35 & ~x36 & ~x44 & ~x51 & ~x53 & ~x54 & ~x57 & ~x64 & ~x68 & ~x76 & ~x78 & ~x83 & ~x87 & ~x89 & ~x97 & ~x99 & ~x100 & ~x107 & ~x109 & ~x110 & ~x125 & ~x128 & ~x141 & ~x143 & ~x151 & ~x153 & ~x154 & ~x157 & ~x158 & ~x167 & ~x169 & ~x171 & ~x174 & ~x227 & ~x283 & ~x307 & ~x309 & ~x311 & ~x365 & ~x366 & ~x393 & ~x416 & ~x419 & ~x420 & ~x423 & ~x442 & ~x446 & ~x452 & ~x469 & ~x470 & ~x473 & ~x480 & ~x502 & ~x530 & ~x532 & ~x535 & ~x555 & ~x556 & ~x564 & ~x581 & ~x586 & ~x619 & ~x641 & ~x644 & ~x646 & ~x668 & ~x673 & ~x674 & ~x676 & ~x677 & ~x695 & ~x699 & ~x705 & ~x706 & ~x724 & ~x725 & ~x728 & ~x733 & ~x734 & ~x746 & ~x751 & ~x755 & ~x764 & ~x783;
assign c4183 =  x519 &  x570 & ~x25 & ~x36 & ~x61 & ~x81 & ~x111 & ~x140 & ~x163 & ~x168 & ~x169 & ~x201 & ~x223 & ~x229 & ~x233 & ~x451 & ~x534 & ~x535 & ~x629 & ~x630 & ~x632 & ~x635 & ~x657 & ~x660 & ~x661 & ~x687 & ~x710 & ~x781;
assign c4185 =  x211 &  x407 &  x408 & ~x6 & ~x8 & ~x120 & ~x138 & ~x160 & ~x168 & ~x205 & ~x245 & ~x332 & ~x344 & ~x359 & ~x390 & ~x398 & ~x421 & ~x455 & ~x495 & ~x496 & ~x528 & ~x560 & ~x639 & ~x667 & ~x720;
assign c4187 = ~x6 & ~x9 & ~x18 & ~x31 & ~x32 & ~x36 & ~x43 & ~x47 & ~x48 & ~x69 & ~x70 & ~x77 & ~x80 & ~x86 & ~x87 & ~x88 & ~x93 & ~x102 & ~x111 & ~x117 & ~x126 & ~x127 & ~x129 & ~x131 & ~x132 & ~x135 & ~x138 & ~x139 & ~x141 & ~x150 & ~x153 & ~x155 & ~x157 & ~x171 & ~x198 & ~x199 & ~x201 & ~x202 & ~x205 & ~x206 & ~x222 & ~x224 & ~x227 & ~x229 & ~x230 & ~x252 & ~x254 & ~x258 & ~x280 & ~x282 & ~x304 & ~x306 & ~x311 & ~x334 & ~x362 & ~x393 & ~x420 & ~x422 & ~x433 & ~x434 & ~x449 & ~x459 & ~x479 & ~x530 & ~x558 & ~x559 & ~x562 & ~x587 & ~x588 & ~x590 & ~x607 & ~x612 & ~x615 & ~x616 & ~x634 & ~x643 & ~x647 & ~x663 & ~x665 & ~x667 & ~x671 & ~x674 & ~x677 & ~x689 & ~x701 & ~x724 & ~x725 & ~x726 & ~x747 & ~x751 & ~x759 & ~x766 & ~x773 & ~x775 & ~x776 & ~x777 & ~x781 & ~x783;
assign c4189 =  x716 & ~x191;
assign c4191 =  x186 & ~x5 & ~x14 & ~x15 & ~x18 & ~x19 & ~x31 & ~x32 & ~x38 & ~x54 & ~x67 & ~x68 & ~x70 & ~x78 & ~x81 & ~x82 & ~x91 & ~x95 & ~x96 & ~x99 & ~x115 & ~x139 & ~x142 & ~x145 & ~x148 & ~x150 & ~x166 & ~x169 & ~x197 & ~x198 & ~x202 & ~x204 & ~x222 & ~x229 & ~x250 & ~x251 & ~x258 & ~x278 & ~x284 & ~x285 & ~x296 & ~x305 & ~x312 & ~x332 & ~x334 & ~x358 & ~x363 & ~x364 & ~x366 & ~x415 & ~x416 & ~x417 & ~x421 & ~x422 & ~x441 & ~x443 & ~x446 & ~x476 & ~x478 & ~x479 & ~x497 & ~x499 & ~x502 & ~x555 & ~x583 & ~x585 & ~x588 & ~x609 & ~x611 & ~x619 & ~x634 & ~x636 & ~x664 & ~x667 & ~x671 & ~x676 & ~x694 & ~x704 & ~x706 & ~x726 & ~x735 & ~x741 & ~x746 & ~x750 & ~x753 & ~x763 & ~x783;
assign c4193 =  x236 &  x238 & ~x18 & ~x30 & ~x54 & ~x99 & ~x102 & ~x106 & ~x113 & ~x147 & ~x159 & ~x173 & ~x195 & ~x197 & ~x230 & ~x231 & ~x256 & ~x306 & ~x332 & ~x387 & ~x394 & ~x421 & ~x439 & ~x495 & ~x506 & ~x526 & ~x543 & ~x552 & ~x583 & ~x609 & ~x616 & ~x669 & ~x768;
assign c4195 = ~x2 & ~x3 & ~x4 & ~x13 & ~x16 & ~x18 & ~x19 & ~x22 & ~x24 & ~x27 & ~x28 & ~x40 & ~x62 & ~x63 & ~x75 & ~x78 & ~x80 & ~x82 & ~x84 & ~x87 & ~x104 & ~x108 & ~x118 & ~x132 & ~x133 & ~x139 & ~x142 & ~x147 & ~x158 & ~x160 & ~x162 & ~x163 & ~x165 & ~x166 & ~x168 & ~x170 & ~x172 & ~x189 & ~x191 & ~x194 & ~x195 & ~x197 & ~x213 & ~x214 & ~x215 & ~x218 & ~x219 & ~x224 & ~x228 & ~x239 & ~x240 & ~x241 & ~x242 & ~x244 & ~x245 & ~x247 & ~x253 & ~x256 & ~x267 & ~x268 & ~x282 & ~x309 & ~x334 & ~x335 & ~x365 & ~x367 & ~x389 & ~x391 & ~x395 & ~x418 & ~x420 & ~x421 & ~x449 & ~x450 & ~x451 & ~x452 & ~x560 & ~x588 & ~x589 & ~x635 & ~x641 & ~x645 & ~x646 & ~x649 & ~x654 & ~x655 & ~x657 & ~x659 & ~x663 & ~x676 & ~x678 & ~x680 & ~x683 & ~x685 & ~x686 & ~x688 & ~x692 & ~x694 & ~x696 & ~x697 & ~x700 & ~x703 & ~x704 & ~x715 & ~x720 & ~x722 & ~x726 & ~x732 & ~x733 & ~x739 & ~x742 & ~x746 & ~x751 & ~x753 & ~x769 & ~x776 & ~x777 & ~x779 & ~x783;
assign c4197 =  x124;
assign c4199 =  x656 & ~x338 & ~x518;
assign c4201 = ~x5 & ~x9 & ~x17 & ~x27 & ~x32 & ~x33 & ~x43 & ~x55 & ~x59 & ~x63 & ~x64 & ~x67 & ~x68 & ~x71 & ~x74 & ~x83 & ~x89 & ~x91 & ~x100 & ~x101 & ~x106 & ~x112 & ~x117 & ~x135 & ~x138 & ~x142 & ~x147 & ~x168 & ~x220 & ~x222 & ~x278 & ~x308 & ~x333 & ~x334 & ~x363 & ~x394 & ~x407 & ~x447 & ~x462 & ~x474 & ~x477 & ~x487 & ~x501 & ~x502 & ~x508 & ~x515 & ~x532 & ~x543 & ~x562 & ~x584 & ~x590 & ~x591 & ~x615 & ~x618 & ~x639 & ~x640 & ~x643 & ~x647 & ~x649 & ~x667 & ~x668 & ~x671 & ~x673 & ~x674 & ~x675 & ~x695 & ~x701 & ~x705 & ~x706 & ~x708 & ~x724 & ~x738 & ~x754 & ~x755 & ~x756 & ~x761 & ~x762 & ~x768 & ~x779;
assign c4203 =  x327 & ~x3 & ~x6 & ~x19 & ~x42 & ~x66 & ~x74 & ~x85 & ~x101 & ~x115 & ~x121 & ~x128 & ~x146 & ~x147 & ~x150 & ~x155 & ~x157 & ~x159 & ~x160 & ~x162 & ~x163 & ~x172 & ~x250 & ~x256 & ~x281 & ~x305 & ~x308 & ~x336 & ~x348 & ~x368 & ~x388 & ~x415 & ~x424 & ~x469 & ~x498 & ~x501 & ~x507 & ~x530 & ~x532 & ~x535 & ~x560 & ~x562 & ~x569 & ~x588 & ~x614 & ~x642 & ~x671 & ~x696 & ~x703 & ~x704 & ~x752 & ~x754;
assign c4205 =  x539 & ~x40 & ~x66 & ~x80 & ~x82 & ~x88 & ~x150 & ~x151 & ~x152 & ~x207 & ~x253 & ~x365 & ~x445 & ~x451 & ~x527 & ~x581 & ~x635 & ~x662 & ~x665 & ~x717 & ~x727 & ~x736 & ~x738 & ~x750 & ~x766;
assign c4207 =  x182 &  x212 & ~x293;
assign c4209 =  x183 &  x184 &  x213 & ~x294 & ~x497;
assign c4211 =  x207 &  x233 & ~x519;
assign c4213 =  x660 & ~x9 & ~x14 & ~x20 & ~x64 & ~x110 & ~x169 & ~x336 & ~x338 & ~x364 & ~x387 & ~x396 & ~x416 & ~x427 & ~x453 & ~x455 & ~x547 & ~x561 & ~x617 & ~x676 & ~x775 & ~x779 & ~x782;
assign c4215 =  x630 &  x631 & ~x3 & ~x14 & ~x16 & ~x55 & ~x65 & ~x66 & ~x73 & ~x86 & ~x87 & ~x88 & ~x95 & ~x97 & ~x143 & ~x144 & ~x169 & ~x170 & ~x172 & ~x192 & ~x199 & ~x250 & ~x251 & ~x308 & ~x311 & ~x331 & ~x332 & ~x337 & ~x341 & ~x367 & ~x387 & ~x396 & ~x399 & ~x412 & ~x441 & ~x454 & ~x455 & ~x472 & ~x473 & ~x484 & ~x501 & ~x507 & ~x508 & ~x526 & ~x535 & ~x538 & ~x592 & ~x593 & ~x617 & ~x645 & ~x669 & ~x670 & ~x673 & ~x681 & ~x693 & ~x696 & ~x713 & ~x729 & ~x740 & ~x748 & ~x754 & ~x756 & ~x761 & ~x771 & ~x782 & ~x783;
assign c4217 = ~x0 & ~x8 & ~x18 & ~x28 & ~x41 & ~x49 & ~x70 & ~x72 & ~x77 & ~x91 & ~x114 & ~x134 & ~x192 & ~x257 & ~x279 & ~x282 & ~x292 & ~x314 & ~x316 & ~x319 & ~x336 & ~x339 & ~x345 & ~x359 & ~x363 & ~x413 & ~x440 & ~x469 & ~x534 & ~x535 & ~x556 & ~x586 & ~x619 & ~x664 & ~x674 & ~x675 & ~x710 & ~x712 & ~x735 & ~x773 & ~x777;
assign c4219 =  x549 & ~x198 & ~x275 & ~x353 & ~x390 & ~x396 & ~x476 & ~x661 & ~x674 & ~x694;
assign c4221 =  x215 &  x246 & ~x24 & ~x80 & ~x82 & ~x88 & ~x93 & ~x172 & ~x232 & ~x233 & ~x390 & ~x444 & ~x641 & ~x722 & ~x733 & ~x752;
assign c4223 = ~x10 & ~x28 & ~x29 & ~x34 & ~x46 & ~x50 & ~x52 & ~x57 & ~x62 & ~x75 & ~x88 & ~x110 & ~x111 & ~x119 & ~x121 & ~x135 & ~x170 & ~x200 & ~x220 & ~x221 & ~x332 & ~x377 & ~x404 & ~x425 & ~x429 & ~x455 & ~x477 & ~x484 & ~x505 & ~x512 & ~x530 & ~x537 & ~x553 & ~x554 & ~x593 & ~x608 & ~x610 & ~x613 & ~x620 & ~x668 & ~x670 & ~x705 & ~x722 & ~x730 & ~x775 & ~x779;
assign c4225 =  x208 &  x209 &  x210 & ~x85 & ~x153 & ~x273 & ~x397 & ~x416 & ~x442 & ~x732 & ~x770 & ~x775;
assign c4227 =  x600 & ~x9 & ~x12 & ~x16 & ~x20 & ~x22 & ~x26 & ~x37 & ~x39 & ~x47 & ~x80 & ~x81 & ~x84 & ~x85 & ~x112 & ~x113 & ~x117 & ~x118 & ~x140 & ~x168 & ~x169 & ~x172 & ~x197 & ~x279 & ~x335 & ~x362 & ~x365 & ~x392 & ~x396 & ~x421 & ~x422 & ~x445 & ~x473 & ~x490 & ~x500 & ~x501 & ~x586 & ~x589 & ~x590 & ~x614 & ~x641 & ~x642 & ~x691 & ~x693 & ~x694 & ~x699 & ~x719 & ~x728 & ~x734 & ~x736 & ~x743 & ~x747 & ~x749 & ~x765 & ~x766 & ~x770 & ~x772 & ~x774;
assign c4229 =  x156 &  x157 &  x568 & ~x499 & ~x767;
assign c4231 = ~x29 & ~x50 & ~x115 & ~x171 & ~x334 & ~x347 & ~x348 & ~x369 & ~x372 & ~x373 & ~x397 & ~x533 & ~x562 & ~x649 & ~x676 & ~x706 & ~x708 & ~x782;
assign c4233 = ~x0 & ~x4 & ~x10 & ~x15 & ~x17 & ~x19 & ~x20 & ~x32 & ~x36 & ~x44 & ~x47 & ~x49 & ~x53 & ~x54 & ~x55 & ~x61 & ~x66 & ~x68 & ~x69 & ~x77 & ~x78 & ~x79 & ~x80 & ~x82 & ~x83 & ~x92 & ~x93 & ~x102 & ~x109 & ~x113 & ~x116 & ~x121 & ~x134 & ~x135 & ~x136 & ~x140 & ~x142 & ~x146 & ~x149 & ~x161 & ~x162 & ~x169 & ~x196 & ~x197 & ~x223 & ~x233 & ~x260 & ~x281 & ~x282 & ~x308 & ~x315 & ~x343 & ~x360 & ~x365 & ~x366 & ~x384 & ~x386 & ~x388 & ~x392 & ~x395 & ~x403 & ~x415 & ~x420 & ~x421 & ~x424 & ~x439 & ~x440 & ~x445 & ~x467 & ~x469 & ~x470 & ~x476 & ~x477 & ~x478 & ~x479 & ~x480 & ~x494 & ~x507 & ~x522 & ~x557 & ~x587 & ~x588 & ~x589 & ~x591 & ~x614 & ~x617 & ~x618 & ~x635 & ~x638 & ~x641 & ~x643 & ~x647 & ~x648 & ~x649 & ~x669 & ~x676 & ~x680 & ~x705 & ~x713 & ~x718 & ~x719 & ~x720 & ~x724 & ~x728 & ~x729 & ~x732 & ~x734 & ~x736 & ~x747 & ~x749 & ~x751 & ~x754 & ~x756 & ~x767 & ~x776;
assign c4235 =  x541 & ~x8 & ~x9 & ~x30 & ~x171 & ~x260 & ~x281 & ~x282 & ~x288 & ~x311 & ~x315 & ~x318 & ~x342 & ~x390 & ~x612 & ~x613 & ~x632 & ~x641 & ~x657 & ~x658 & ~x662 & ~x684 & ~x685 & ~x713 & ~x747 & ~x772 & ~x778;
assign c4237 =  x182 &  x184 & ~x265;
assign c4239 = ~x1 & ~x2 & ~x7 & ~x25 & ~x30 & ~x32 & ~x46 & ~x49 & ~x51 & ~x52 & ~x53 & ~x61 & ~x74 & ~x79 & ~x106 & ~x137 & ~x142 & ~x144 & ~x172 & ~x202 & ~x220 & ~x255 & ~x256 & ~x280 & ~x283 & ~x311 & ~x313 & ~x335 & ~x339 & ~x340 & ~x363 & ~x386 & ~x387 & ~x388 & ~x392 & ~x395 & ~x415 & ~x437 & ~x443 & ~x444 & ~x447 & ~x450 & ~x452 & ~x454 & ~x456 & ~x465 & ~x475 & ~x506 & ~x535 & ~x536 & ~x560 & ~x562 & ~x563 & ~x586 & ~x587 & ~x615 & ~x636 & ~x637 & ~x642 & ~x647 & ~x666 & ~x686 & ~x689 & ~x690 & ~x692 & ~x695 & ~x700 & ~x702 & ~x704 & ~x710 & ~x713 & ~x715 & ~x722 & ~x733 & ~x734 & ~x737 & ~x741 & ~x747 & ~x750 & ~x753 & ~x763 & ~x765 & ~x769;
assign c4241 =  x185 &  x186 &  x215 & ~x10 & ~x16 & ~x22 & ~x26 & ~x28 & ~x31 & ~x32 & ~x43 & ~x46 & ~x52 & ~x61 & ~x62 & ~x64 & ~x70 & ~x80 & ~x81 & ~x90 & ~x94 & ~x96 & ~x98 & ~x99 & ~x110 & ~x115 & ~x119 & ~x124 & ~x126 & ~x135 & ~x141 & ~x146 & ~x148 & ~x151 & ~x169 & ~x170 & ~x172 & ~x173 & ~x174 & ~x177 & ~x193 & ~x194 & ~x199 & ~x200 & ~x203 & ~x221 & ~x227 & ~x229 & ~x230 & ~x253 & ~x257 & ~x258 & ~x277 & ~x279 & ~x281 & ~x286 & ~x287 & ~x308 & ~x337 & ~x340 & ~x365 & ~x366 & ~x369 & ~x396 & ~x419 & ~x441 & ~x446 & ~x470 & ~x471 & ~x474 & ~x496 & ~x498 & ~x502 & ~x525 & ~x526 & ~x528 & ~x530 & ~x555 & ~x561 & ~x562 & ~x581 & ~x583 & ~x587 & ~x590 & ~x615 & ~x643 & ~x662 & ~x665 & ~x667 & ~x669 & ~x670 & ~x671 & ~x673 & ~x676 & ~x695 & ~x696 & ~x699 & ~x700 & ~x705 & ~x721 & ~x722 & ~x723 & ~x726 & ~x727 & ~x743 & ~x747 & ~x748 & ~x751 & ~x752 & ~x753 & ~x756 & ~x757 & ~x759 & ~x761 & ~x765 & ~x766 & ~x767 & ~x773 & ~x774 & ~x775 & ~x779;
assign c4243 =  x180 &  x183 & ~x4 & ~x31 & ~x34 & ~x61 & ~x81 & ~x113 & ~x138 & ~x170 & ~x248 & ~x336 & ~x337 & ~x338 & ~x414 & ~x594 & ~x619 & ~x641 & ~x650 & ~x727 & ~x728 & ~x783;
assign c4245 =  x357 &  x514 & ~x47 & ~x111 & ~x164 & ~x220 & ~x275 & ~x276 & ~x446 & ~x530 & ~x582 & ~x609 & ~x610 & ~x637 & ~x681;
assign c4247 = ~x4 & ~x14 & ~x15 & ~x21 & ~x26 & ~x31 & ~x34 & ~x37 & ~x41 & ~x45 & ~x46 & ~x52 & ~x53 & ~x58 & ~x61 & ~x75 & ~x81 & ~x84 & ~x85 & ~x87 & ~x90 & ~x109 & ~x118 & ~x137 & ~x171 & ~x177 & ~x199 & ~x226 & ~x227 & ~x253 & ~x254 & ~x284 & ~x309 & ~x333 & ~x337 & ~x365 & ~x366 & ~x368 & ~x384 & ~x389 & ~x397 & ~x412 & ~x447 & ~x449 & ~x478 & ~x490 & ~x501 & ~x529 & ~x534 & ~x562 & ~x586 & ~x588 & ~x639 & ~x645 & ~x660 & ~x666 & ~x672 & ~x690 & ~x691 & ~x695 & ~x704 & ~x716 & ~x717 & ~x718 & ~x724 & ~x733 & ~x735 & ~x739 & ~x745 & ~x749 & ~x753 & ~x758 & ~x760 & ~x763;
assign c4249 = ~x14 & ~x16 & ~x25 & ~x45 & ~x59 & ~x71 & ~x82 & ~x88 & ~x91 & ~x103 & ~x109 & ~x118 & ~x193 & ~x198 & ~x222 & ~x223 & ~x252 & ~x277 & ~x306 & ~x365 & ~x390 & ~x461 & ~x462 & ~x464 & ~x475 & ~x479 & ~x480 & ~x501 & ~x502 & ~x517 & ~x589 & ~x590 & ~x638 & ~x645 & ~x646 & ~x648 & ~x692 & ~x697 & ~x698 & ~x703 & ~x738 & ~x753 & ~x774 & ~x779;
assign c4251 = ~x24 & ~x50 & ~x142 & ~x209 & ~x250 & ~x317 & ~x372 & ~x399 & ~x429 & ~x454 & ~x456 & ~x583 & ~x617 & ~x688 & ~x729 & ~x756 & ~x762;
assign c4253 =  x233 &  x235 &  x236 &  x237 & ~x13 & ~x536 & ~x734 & ~x770;
assign c4255 = ~x19 & ~x20 & ~x38 & ~x41 & ~x73 & ~x87 & ~x88 & ~x112 & ~x117 & ~x168 & ~x194 & ~x224 & ~x225 & ~x249 & ~x255 & ~x282 & ~x286 & ~x287 & ~x291 & ~x292 & ~x318 & ~x320 & ~x344 & ~x347 & ~x365 & ~x388 & ~x420 & ~x476 & ~x532 & ~x590 & ~x637 & ~x646 & ~x669 & ~x701 & ~x710 & ~x721 & ~x724 & ~x729 & ~x730 & ~x765 & ~x766 & ~x773 & ~x776 & ~x780 & ~x781;
assign c4257 =  x742;
assign c4259 =  x551 &  x576 & ~x215 & ~x240 & ~x241;
assign c4261 =  x238 &  x486 &  x487 & ~x412 & ~x441 & ~x468;
assign c4263 =  x571 & ~x1 & ~x2 & ~x51 & ~x136 & ~x217 & ~x246 & ~x248 & ~x275 & ~x340 & ~x593 & ~x614 & ~x653 & ~x683 & ~x684 & ~x708;
assign c4265 = ~x0 & ~x20 & ~x23 & ~x25 & ~x27 & ~x40 & ~x52 & ~x85 & ~x86 & ~x118 & ~x141 & ~x145 & ~x146 & ~x151 & ~x154 & ~x181 & ~x198 & ~x224 & ~x254 & ~x256 & ~x381 & ~x488 & ~x507 & ~x530 & ~x557 & ~x558 & ~x560 & ~x561 & ~x611 & ~x637 & ~x643 & ~x647 & ~x676 & ~x692 & ~x702 & ~x703 & ~x723 & ~x727 & ~x747 & ~x767 & ~x774;
assign c4267 =  x240 &  x241 &  x266 &  x300 & ~x7 & ~x26 & ~x55 & ~x57 & ~x62 & ~x68 & ~x80 & ~x85 & ~x86 & ~x95 & ~x116 & ~x117 & ~x122 & ~x144 & ~x148 & ~x152 & ~x166 & ~x169 & ~x191 & ~x195 & ~x306 & ~x417 & ~x446 & ~x450 & ~x479 & ~x500 & ~x585 & ~x615 & ~x673;
assign c4269 = ~x6 & ~x7 & ~x14 & ~x17 & ~x18 & ~x20 & ~x23 & ~x27 & ~x28 & ~x31 & ~x34 & ~x37 & ~x46 & ~x47 & ~x50 & ~x56 & ~x57 & ~x61 & ~x63 & ~x78 & ~x88 & ~x90 & ~x91 & ~x109 & ~x110 & ~x118 & ~x120 & ~x140 & ~x142 & ~x167 & ~x171 & ~x173 & ~x174 & ~x194 & ~x195 & ~x200 & ~x201 & ~x227 & ~x230 & ~x253 & ~x275 & ~x276 & ~x280 & ~x282 & ~x283 & ~x304 & ~x306 & ~x335 & ~x347 & ~x348 & ~x360 & ~x366 & ~x367 & ~x369 & ~x372 & ~x374 & ~x388 & ~x394 & ~x424 & ~x449 & ~x503 & ~x505 & ~x533 & ~x534 & ~x583 & ~x586 & ~x618 & ~x619 & ~x640 & ~x641 & ~x642 & ~x669 & ~x671 & ~x692 & ~x701 & ~x705 & ~x707 & ~x711 & ~x712 & ~x713 & ~x728 & ~x741 & ~x745 & ~x747 & ~x748 & ~x753 & ~x754 & ~x755 & ~x757 & ~x758 & ~x759 & ~x762 & ~x765;
assign c4271 = ~x2 & ~x43 & ~x44 & ~x75 & ~x109 & ~x136 & ~x144 & ~x194 & ~x201 & ~x225 & ~x252 & ~x311 & ~x334 & ~x338 & ~x355 & ~x356 & ~x382 & ~x383 & ~x394 & ~x396 & ~x400 & ~x409 & ~x410 & ~x417 & ~x423 & ~x428 & ~x437 & ~x438 & ~x439 & ~x466 & ~x468 & ~x479 & ~x505 & ~x507 & ~x558 & ~x559 & ~x562 & ~x564 & ~x592 & ~x619 & ~x640 & ~x642 & ~x668 & ~x676 & ~x693 & ~x700 & ~x704 & ~x717 & ~x732 & ~x735 & ~x750 & ~x759 & ~x781;
assign c4273 =  x208 &  x210 & ~x26 & ~x54 & ~x78 & ~x137 & ~x139 & ~x163 & ~x219 & ~x320 & ~x368 & ~x386 & ~x418 & ~x499 & ~x647 & ~x736 & ~x769 & ~x771;
assign c4275 =  x654 &  x655 & ~x26 & ~x84 & ~x141 & ~x223 & ~x516 & ~x543;
assign c4277 =  x293 & ~x17 & ~x69 & ~x100 & ~x112 & ~x130 & ~x139 & ~x143 & ~x148 & ~x158 & ~x168 & ~x183 & ~x184 & ~x190 & ~x222 & ~x251 & ~x279 & ~x280 & ~x307 & ~x363 & ~x365 & ~x367 & ~x390 & ~x431 & ~x432 & ~x446 & ~x450 & ~x505 & ~x508 & ~x540 & ~x668 & ~x693 & ~x697 & ~x701 & ~x706 & ~x728 & ~x754 & ~x758 & ~x765 & ~x766 & ~x767;
assign c4279 =  x433 & ~x27 & ~x43 & ~x91 & ~x108 & ~x136 & ~x143 & ~x149 & ~x163 & ~x219 & ~x223 & ~x250 & ~x340 & ~x347 & ~x371 & ~x372 & ~x389 & ~x473 & ~x476 & ~x556 & ~x561 & ~x611 & ~x666 & ~x709 & ~x744 & ~x750 & ~x782 & ~x783;
assign c4281 =  x237 &  x240 &  x270 & ~x0 & ~x11 & ~x37 & ~x43 & ~x47 & ~x67 & ~x80 & ~x85 & ~x86 & ~x90 & ~x107 & ~x122 & ~x127 & ~x132 & ~x151 & ~x154 & ~x157 & ~x158 & ~x159 & ~x165 & ~x191 & ~x251 & ~x282 & ~x309 & ~x363 & ~x394 & ~x414 & ~x415 & ~x447 & ~x528 & ~x529 & ~x532 & ~x559 & ~x564 & ~x567 & ~x569 & ~x587 & ~x597 & ~x598 & ~x619 & ~x622 & ~x647 & ~x648 & ~x673 & ~x700 & ~x769 & ~x779;
assign c4283 = ~x0 & ~x15 & ~x26 & ~x27 & ~x29 & ~x33 & ~x41 & ~x47 & ~x56 & ~x58 & ~x63 & ~x65 & ~x75 & ~x77 & ~x83 & ~x85 & ~x104 & ~x109 & ~x117 & ~x121 & ~x138 & ~x144 & ~x166 & ~x169 & ~x171 & ~x173 & ~x176 & ~x221 & ~x227 & ~x259 & ~x277 & ~x284 & ~x307 & ~x310 & ~x320 & ~x343 & ~x346 & ~x366 & ~x367 & ~x393 & ~x416 & ~x421 & ~x503 & ~x505 & ~x532 & ~x584 & ~x587 & ~x612 & ~x635 & ~x645 & ~x646 & ~x665 & ~x672 & ~x691 & ~x692 & ~x695 & ~x701 & ~x705 & ~x718 & ~x726 & ~x727 & ~x728 & ~x734 & ~x745 & ~x750 & ~x755 & ~x769 & ~x773;
assign c4285 =  x330;
assign c4287 = ~x8 & ~x11 & ~x15 & ~x17 & ~x20 & ~x21 & ~x22 & ~x25 & ~x28 & ~x32 & ~x35 & ~x42 & ~x46 & ~x54 & ~x59 & ~x69 & ~x70 & ~x72 & ~x77 & ~x79 & ~x80 & ~x85 & ~x104 & ~x107 & ~x108 & ~x111 & ~x112 & ~x113 & ~x117 & ~x118 & ~x119 & ~x135 & ~x137 & ~x140 & ~x151 & ~x152 & ~x153 & ~x162 & ~x163 & ~x166 & ~x169 & ~x177 & ~x178 & ~x182 & ~x193 & ~x198 & ~x201 & ~x204 & ~x207 & ~x224 & ~x229 & ~x231 & ~x232 & ~x250 & ~x256 & ~x257 & ~x283 & ~x309 & ~x313 & ~x360 & ~x385 & ~x389 & ~x419 & ~x422 & ~x439 & ~x440 & ~x444 & ~x452 & ~x469 & ~x473 & ~x475 & ~x476 & ~x488 & ~x496 & ~x502 & ~x506 & ~x552 & ~x560 & ~x564 & ~x565 & ~x578 & ~x580 & ~x606 & ~x613 & ~x618 & ~x633 & ~x638 & ~x642 & ~x643 & ~x644 & ~x659 & ~x660 & ~x661 & ~x664 & ~x669 & ~x670 & ~x688 & ~x689 & ~x692 & ~x705 & ~x715 & ~x718 & ~x720 & ~x722 & ~x727 & ~x728 & ~x750 & ~x760 & ~x761 & ~x764;
assign c4289 =  x183 &  x214 & ~x324;
assign c4291 =  x549 &  x600 & ~x11 & ~x41 & ~x48 & ~x141 & ~x314 & ~x555 & ~x663 & ~x683 & ~x702 & ~x740;
assign c4293 =  x236 &  x238 & ~x42 & ~x49 & ~x52 & ~x55 & ~x65 & ~x79 & ~x84 & ~x109 & ~x112 & ~x122 & ~x153 & ~x231 & ~x258 & ~x393 & ~x412 & ~x447 & ~x476 & ~x506 & ~x516 & ~x534 & ~x562 & ~x642 & ~x775;
assign c4295 =  x213 &  x214 &  x238 & ~x48 & ~x59 & ~x70 & ~x105 & ~x122 & ~x296 & ~x414 & ~x442 & ~x451 & ~x468 & ~x637 & ~x663 & ~x762;
assign c4297 =  x259 & ~x164 & ~x169 & ~x188 & ~x275 & ~x372 & ~x373 & ~x401 & ~x421 & ~x621;
assign c4299 =  x183 &  x184 &  x657 & ~x469 & ~x495;
assign c50 =  x207 &  x235 &  x263 &  x291 &  x319 &  x467 &  x495 & ~x0 & ~x9 & ~x19 & ~x23 & ~x25 & ~x31 & ~x33 & ~x34 & ~x36 & ~x46 & ~x47 & ~x53 & ~x60 & ~x70 & ~x77 & ~x86 & ~x93 & ~x115 & ~x117 & ~x118 & ~x119 & ~x120 & ~x135 & ~x137 & ~x144 & ~x148 & ~x168 & ~x169 & ~x172 & ~x192 & ~x196 & ~x197 & ~x224 & ~x229 & ~x250 & ~x274 & ~x283 & ~x284 & ~x285 & ~x305 & ~x307 & ~x311 & ~x329 & ~x332 & ~x334 & ~x341 & ~x342 & ~x359 & ~x363 & ~x396 & ~x397 & ~x417 & ~x422 & ~x428 & ~x429 & ~x444 & ~x445 & ~x447 & ~x449 & ~x450 & ~x474 & ~x475 & ~x476 & ~x478 & ~x500 & ~x503 & ~x504 & ~x505 & ~x529 & ~x531 & ~x533 & ~x534 & ~x555 & ~x557 & ~x561 & ~x585 & ~x591 & ~x610 & ~x614 & ~x617 & ~x641 & ~x642 & ~x643 & ~x645 & ~x671 & ~x674 & ~x694 & ~x697 & ~x698 & ~x703 & ~x705 & ~x706 & ~x715 & ~x717 & ~x719 & ~x721 & ~x725 & ~x733 & ~x734 & ~x736 & ~x744 & ~x746 & ~x747 & ~x748 & ~x752 & ~x753 & ~x754 & ~x756 & ~x761 & ~x765 & ~x767 & ~x769 & ~x770 & ~x771 & ~x772 & ~x778;
assign c52 = ~x0 & ~x3 & ~x6 & ~x13 & ~x16 & ~x22 & ~x28 & ~x30 & ~x31 & ~x33 & ~x34 & ~x36 & ~x38 & ~x43 & ~x46 & ~x50 & ~x52 & ~x53 & ~x54 & ~x56 & ~x57 & ~x58 & ~x61 & ~x62 & ~x63 & ~x64 & ~x69 & ~x70 & ~x73 & ~x77 & ~x78 & ~x83 & ~x85 & ~x87 & ~x89 & ~x91 & ~x92 & ~x93 & ~x94 & ~x108 & ~x110 & ~x112 & ~x116 & ~x118 & ~x119 & ~x135 & ~x136 & ~x137 & ~x144 & ~x146 & ~x147 & ~x167 & ~x170 & ~x173 & ~x195 & ~x196 & ~x198 & ~x200 & ~x218 & ~x219 & ~x225 & ~x226 & ~x227 & ~x240 & ~x241 & ~x243 & ~x244 & ~x245 & ~x246 & ~x249 & ~x252 & ~x255 & ~x257 & ~x267 & ~x269 & ~x270 & ~x272 & ~x273 & ~x274 & ~x275 & ~x276 & ~x277 & ~x278 & ~x299 & ~x300 & ~x301 & ~x307 & ~x329 & ~x333 & ~x334 & ~x338 & ~x361 & ~x362 & ~x363 & ~x390 & ~x391 & ~x392 & ~x395 & ~x396 & ~x417 & ~x419 & ~x424 & ~x445 & ~x449 & ~x451 & ~x460 & ~x461 & ~x462 & ~x474 & ~x476 & ~x478 & ~x479 & ~x480 & ~x482 & ~x486 & ~x487 & ~x488 & ~x489 & ~x490 & ~x503 & ~x507 & ~x531 & ~x534 & ~x535 & ~x559 & ~x560 & ~x561 & ~x562 & ~x584 & ~x590 & ~x611 & ~x613 & ~x615 & ~x642 & ~x643 & ~x646 & ~x647 & ~x664 & ~x666 & ~x667 & ~x672 & ~x675 & ~x676 & ~x677 & ~x678 & ~x680 & ~x687 & ~x688 & ~x689 & ~x691 & ~x692 & ~x693 & ~x694 & ~x696 & ~x699 & ~x701 & ~x702 & ~x703 & ~x704 & ~x709 & ~x710 & ~x712 & ~x714 & ~x715 & ~x716 & ~x718 & ~x719 & ~x720 & ~x722 & ~x723 & ~x724 & ~x728 & ~x730 & ~x732 & ~x733 & ~x735 & ~x739 & ~x741 & ~x743 & ~x745 & ~x748 & ~x750 & ~x751 & ~x752 & ~x753 & ~x754 & ~x755 & ~x756 & ~x758 & ~x760 & ~x762 & ~x765 & ~x768 & ~x773 & ~x774 & ~x775 & ~x776 & ~x778 & ~x780;
assign c54 =  x110;
assign c56 =  x347 &  x403 & ~x2 & ~x4 & ~x7 & ~x9 & ~x16 & ~x18 & ~x21 & ~x23 & ~x32 & ~x36 & ~x37 & ~x40 & ~x43 & ~x45 & ~x46 & ~x49 & ~x51 & ~x52 & ~x53 & ~x56 & ~x60 & ~x64 & ~x65 & ~x69 & ~x85 & ~x87 & ~x90 & ~x91 & ~x97 & ~x119 & ~x120 & ~x121 & ~x123 & ~x125 & ~x139 & ~x141 & ~x142 & ~x146 & ~x165 & ~x171 & ~x175 & ~x176 & ~x178 & ~x194 & ~x202 & ~x223 & ~x227 & ~x228 & ~x232 & ~x252 & ~x253 & ~x254 & ~x255 & ~x282 & ~x284 & ~x307 & ~x336 & ~x366 & ~x367 & ~x386 & ~x389 & ~x391 & ~x393 & ~x417 & ~x442 & ~x445 & ~x447 & ~x449 & ~x450 & ~x453 & ~x470 & ~x474 & ~x475 & ~x476 & ~x477 & ~x479 & ~x480 & ~x481 & ~x483 & ~x501 & ~x512 & ~x525 & ~x530 & ~x534 & ~x542 & ~x543 & ~x552 & ~x558 & ~x583 & ~x587 & ~x588 & ~x590 & ~x613 & ~x615 & ~x616 & ~x621 & ~x644 & ~x662 & ~x663 & ~x666 & ~x668 & ~x672 & ~x675 & ~x676 & ~x691 & ~x694 & ~x698 & ~x699 & ~x701 & ~x703 & ~x704 & ~x710 & ~x713 & ~x714 & ~x715 & ~x716 & ~x717 & ~x719 & ~x722 & ~x725 & ~x727 & ~x733 & ~x736 & ~x738 & ~x744 & ~x745 & ~x754 & ~x760 & ~x770 & ~x777 & ~x778 & ~x780 & ~x781;
assign c58 =  x755;
assign c510 =  x687;
assign c512 =  x314 &  x499;
assign c514 =  x45;
assign c516 = ~x0 & ~x1 & ~x3 & ~x20 & ~x31 & ~x35 & ~x48 & ~x79 & ~x94 & ~x106 & ~x120 & ~x141 & ~x145 & ~x165 & ~x169 & ~x173 & ~x174 & ~x197 & ~x203 & ~x226 & ~x227 & ~x251 & ~x260 & ~x274 & ~x282 & ~x287 & ~x294 & ~x295 & ~x297 & ~x298 & ~x300 & ~x301 & ~x308 & ~x313 & ~x314 & ~x327 & ~x328 & ~x329 & ~x330 & ~x337 & ~x357 & ~x360 & ~x387 & ~x394 & ~x398 & ~x428 & ~x444 & ~x479 & ~x500 & ~x518 & ~x519 & ~x529 & ~x531 & ~x532 & ~x545 & ~x557 & ~x564 & ~x610 & ~x613 & ~x615 & ~x647 & ~x648 & ~x663 & ~x665 & ~x668 & ~x670 & ~x673 & ~x676 & ~x678 & ~x694 & ~x705 & ~x710 & ~x717 & ~x739 & ~x742 & ~x751 & ~x753 & ~x758 & ~x759 & ~x762 & ~x764 & ~x765 & ~x766 & ~x775;
assign c518 =  x262 &  x290 & ~x0 & ~x4 & ~x5 & ~x6 & ~x7 & ~x8 & ~x9 & ~x12 & ~x17 & ~x18 & ~x20 & ~x21 & ~x22 & ~x23 & ~x24 & ~x28 & ~x29 & ~x30 & ~x33 & ~x37 & ~x38 & ~x39 & ~x41 & ~x42 & ~x45 & ~x47 & ~x48 & ~x50 & ~x51 & ~x52 & ~x53 & ~x54 & ~x56 & ~x57 & ~x59 & ~x64 & ~x67 & ~x69 & ~x74 & ~x75 & ~x76 & ~x79 & ~x80 & ~x87 & ~x91 & ~x94 & ~x105 & ~x106 & ~x107 & ~x110 & ~x114 & ~x118 & ~x138 & ~x141 & ~x142 & ~x147 & ~x165 & ~x166 & ~x167 & ~x168 & ~x169 & ~x171 & ~x173 & ~x191 & ~x196 & ~x198 & ~x199 & ~x202 & ~x216 & ~x220 & ~x221 & ~x226 & ~x227 & ~x230 & ~x250 & ~x257 & ~x258 & ~x276 & ~x277 & ~x285 & ~x302 & ~x303 & ~x304 & ~x305 & ~x306 & ~x333 & ~x337 & ~x339 & ~x341 & ~x360 & ~x361 & ~x363 & ~x364 & ~x368 & ~x370 & ~x371 & ~x388 & ~x392 & ~x393 & ~x394 & ~x395 & ~x396 & ~x397 & ~x416 & ~x421 & ~x423 & ~x427 & ~x428 & ~x445 & ~x446 & ~x457 & ~x472 & ~x473 & ~x477 & ~x478 & ~x486 & ~x487 & ~x488 & ~x489 & ~x507 & ~x517 & ~x527 & ~x528 & ~x532 & ~x534 & ~x555 & ~x561 & ~x586 & ~x587 & ~x588 & ~x590 & ~x614 & ~x615 & ~x616 & ~x619 & ~x640 & ~x643 & ~x648 & ~x650 & ~x667 & ~x669 & ~x673 & ~x676 & ~x679 & ~x693 & ~x695 & ~x699 & ~x702 & ~x703 & ~x705 & ~x706 & ~x708 & ~x710 & ~x712 & ~x717 & ~x719 & ~x720 & ~x723 & ~x725 & ~x726 & ~x730 & ~x733 & ~x736 & ~x740 & ~x741 & ~x742 & ~x745 & ~x746 & ~x749 & ~x750 & ~x752 & ~x753 & ~x756 & ~x757 & ~x759 & ~x760 & ~x761 & ~x763 & ~x774 & ~x779 & ~x780 & ~x781;
assign c520 =  x731;
assign c522 =  x21;
assign c524 = ~x104 & ~x135 & ~x164 & ~x213 & ~x215 & ~x217 & ~x237 & ~x238 & ~x307 & ~x411 & ~x522 & ~x523 & ~x549 & ~x562 & ~x650 & ~x708;
assign c526 = ~x0 & ~x3 & ~x17 & ~x18 & ~x21 & ~x38 & ~x44 & ~x67 & ~x70 & ~x90 & ~x102 & ~x105 & ~x106 & ~x109 & ~x112 & ~x113 & ~x117 & ~x120 & ~x125 & ~x134 & ~x136 & ~x141 & ~x158 & ~x160 & ~x166 & ~x194 & ~x200 & ~x201 & ~x203 & ~x223 & ~x250 & ~x280 & ~x283 & ~x285 & ~x338 & ~x339 & ~x350 & ~x351 & ~x352 & ~x382 & ~x388 & ~x416 & ~x417 & ~x418 & ~x419 & ~x440 & ~x451 & ~x467 & ~x469 & ~x472 & ~x477 & ~x500 & ~x564 & ~x582 & ~x586 & ~x641 & ~x666 & ~x674 & ~x675 & ~x704 & ~x724 & ~x733 & ~x747 & ~x749 & ~x761 & ~x778 & ~x783;
assign c528 =  x198;
assign c530 =  x216 & ~x5 & ~x6 & ~x14 & ~x18 & ~x21 & ~x36 & ~x44 & ~x48 & ~x56 & ~x63 & ~x64 & ~x66 & ~x75 & ~x78 & ~x88 & ~x98 & ~x108 & ~x109 & ~x121 & ~x122 & ~x126 & ~x135 & ~x149 & ~x197 & ~x203 & ~x225 & ~x228 & ~x275 & ~x285 & ~x298 & ~x299 & ~x300 & ~x329 & ~x338 & ~x356 & ~x359 & ~x368 & ~x386 & ~x392 & ~x414 & ~x445 & ~x451 & ~x473 & ~x498 & ~x500 & ~x504 & ~x530 & ~x533 & ~x556 & ~x584 & ~x667 & ~x670 & ~x671 & ~x674 & ~x693 & ~x701 & ~x719 & ~x720 & ~x726 & ~x733 & ~x743 & ~x750 & ~x751 & ~x754 & ~x757 & ~x763 & ~x764 & ~x766 & ~x768;
assign c532 =  x348 & ~x22 & ~x90 & ~x118 & ~x122 & ~x127 & ~x133 & ~x136 & ~x143 & ~x158 & ~x159 & ~x164 & ~x184 & ~x234 & ~x279 & ~x342 & ~x343 & ~x385 & ~x446 & ~x470 & ~x474 & ~x607 & ~x608 & ~x684 & ~x686 & ~x704 & ~x737 & ~x739 & ~x747;
assign c534 =  x265 & ~x13 & ~x14 & ~x27 & ~x29 & ~x48 & ~x67 & ~x69 & ~x76 & ~x83 & ~x84 & ~x122 & ~x123 & ~x124 & ~x141 & ~x178 & ~x205 & ~x206 & ~x253 & ~x280 & ~x285 & ~x300 & ~x305 & ~x308 & ~x330 & ~x388 & ~x414 & ~x457 & ~x459 & ~x474 & ~x478 & ~x498 & ~x527 & ~x533 & ~x555 & ~x561 & ~x583 & ~x608 & ~x616 & ~x617 & ~x633 & ~x639 & ~x646 & ~x666 & ~x695 & ~x713 & ~x714 & ~x739 & ~x743 & ~x748 & ~x756 & ~x762;
assign c536 =  x287 & ~x7 & ~x16 & ~x21 & ~x46 & ~x54 & ~x64 & ~x65 & ~x66 & ~x107 & ~x137 & ~x163 & ~x170 & ~x191 & ~x192 & ~x194 & ~x227 & ~x228 & ~x276 & ~x279 & ~x301 & ~x303 & ~x331 & ~x335 & ~x360 & ~x421 & ~x460 & ~x481 & ~x483 & ~x484 & ~x486 & ~x488 & ~x519 & ~x520 & ~x521 & ~x530 & ~x559 & ~x592 & ~x612 & ~x619 & ~x640 & ~x699 & ~x706 & ~x732 & ~x739 & ~x757 & ~x759 & ~x765 & ~x771 & ~x774;
assign c538 =  x275 & ~x386 & ~x387 & ~x415;
assign c540 = ~x9 & ~x10 & ~x22 & ~x30 & ~x34 & ~x37 & ~x50 & ~x52 & ~x54 & ~x56 & ~x70 & ~x85 & ~x95 & ~x96 & ~x100 & ~x107 & ~x108 & ~x121 & ~x123 & ~x126 & ~x134 & ~x139 & ~x140 & ~x141 & ~x143 & ~x165 & ~x170 & ~x201 & ~x202 & ~x223 & ~x229 & ~x256 & ~x284 & ~x308 & ~x311 & ~x323 & ~x324 & ~x328 & ~x337 & ~x339 & ~x352 & ~x353 & ~x354 & ~x362 & ~x368 & ~x382 & ~x394 & ~x414 & ~x421 & ~x423 & ~x473 & ~x474 & ~x505 & ~x514 & ~x530 & ~x533 & ~x536 & ~x540 & ~x543 & ~x544 & ~x557 & ~x563 & ~x564 & ~x583 & ~x585 & ~x591 & ~x615 & ~x639 & ~x640 & ~x670 & ~x674 & ~x675 & ~x693 & ~x701 & ~x707 & ~x726 & ~x735 & ~x751 & ~x755 & ~x758 & ~x759 & ~x770 & ~x782;
assign c542 =  x206 & ~x2 & ~x13 & ~x16 & ~x21 & ~x23 & ~x24 & ~x28 & ~x31 & ~x35 & ~x42 & ~x43 & ~x44 & ~x48 & ~x49 & ~x50 & ~x55 & ~x57 & ~x60 & ~x64 & ~x68 & ~x72 & ~x74 & ~x75 & ~x82 & ~x85 & ~x86 & ~x90 & ~x93 & ~x94 & ~x95 & ~x101 & ~x107 & ~x110 & ~x112 & ~x117 & ~x118 & ~x135 & ~x137 & ~x139 & ~x140 & ~x142 & ~x145 & ~x163 & ~x171 & ~x172 & ~x225 & ~x228 & ~x248 & ~x250 & ~x251 & ~x252 & ~x256 & ~x266 & ~x267 & ~x269 & ~x270 & ~x271 & ~x272 & ~x275 & ~x282 & ~x300 & ~x301 & ~x303 & ~x304 & ~x306 & ~x307 & ~x309 & ~x331 & ~x332 & ~x334 & ~x336 & ~x366 & ~x368 & ~x394 & ~x395 & ~x418 & ~x419 & ~x420 & ~x424 & ~x447 & ~x448 & ~x450 & ~x473 & ~x475 & ~x476 & ~x478 & ~x479 & ~x489 & ~x502 & ~x505 & ~x519 & ~x520 & ~x529 & ~x533 & ~x534 & ~x542 & ~x543 & ~x546 & ~x562 & ~x612 & ~x614 & ~x616 & ~x617 & ~x639 & ~x640 & ~x641 & ~x646 & ~x667 & ~x671 & ~x676 & ~x677 & ~x678 & ~x697 & ~x699 & ~x700 & ~x701 & ~x703 & ~x711 & ~x721 & ~x724 & ~x727 & ~x729 & ~x730 & ~x733 & ~x734 & ~x738 & ~x739 & ~x740 & ~x742 & ~x751 & ~x754 & ~x763 & ~x765 & ~x766 & ~x768 & ~x769 & ~x770 & ~x771 & ~x773 & ~x774 & ~x775 & ~x777;
assign c544 =  x297 &  x375 & ~x189 & ~x214 & ~x215 & ~x217 & ~x383 & ~x411;
assign c546 =  x668;
assign c548 =  x613;
assign c550 =  x323 &  x324 & ~x212 & ~x214 & ~x215 & ~x216 & ~x523;
assign c552 =  x271 & ~x10 & ~x57 & ~x118 & ~x121 & ~x155 & ~x159 & ~x186 & ~x188 & ~x202 & ~x258 & ~x355 & ~x357 & ~x361 & ~x368 & ~x386 & ~x416 & ~x449 & ~x651 & ~x695 & ~x727;
assign c554 =  x184 &  x208 & ~x4 & ~x5 & ~x6 & ~x9 & ~x12 & ~x13 & ~x22 & ~x26 & ~x27 & ~x30 & ~x31 & ~x33 & ~x39 & ~x40 & ~x41 & ~x42 & ~x43 & ~x47 & ~x50 & ~x51 & ~x53 & ~x55 & ~x56 & ~x58 & ~x59 & ~x63 & ~x64 & ~x67 & ~x69 & ~x70 & ~x74 & ~x75 & ~x79 & ~x81 & ~x86 & ~x88 & ~x89 & ~x91 & ~x93 & ~x107 & ~x109 & ~x110 & ~x111 & ~x113 & ~x115 & ~x118 & ~x119 & ~x120 & ~x141 & ~x143 & ~x144 & ~x145 & ~x147 & ~x163 & ~x166 & ~x167 & ~x173 & ~x193 & ~x194 & ~x196 & ~x199 & ~x200 & ~x219 & ~x220 & ~x225 & ~x228 & ~x240 & ~x241 & ~x242 & ~x243 & ~x244 & ~x247 & ~x250 & ~x251 & ~x270 & ~x272 & ~x273 & ~x274 & ~x276 & ~x279 & ~x280 & ~x303 & ~x304 & ~x305 & ~x308 & ~x310 & ~x313 & ~x334 & ~x336 & ~x338 & ~x360 & ~x361 & ~x362 & ~x363 & ~x365 & ~x366 & ~x368 & ~x389 & ~x392 & ~x393 & ~x397 & ~x416 & ~x418 & ~x420 & ~x421 & ~x422 & ~x444 & ~x447 & ~x448 & ~x451 & ~x452 & ~x453 & ~x454 & ~x472 & ~x474 & ~x475 & ~x480 & ~x483 & ~x501 & ~x528 & ~x529 & ~x531 & ~x532 & ~x533 & ~x557 & ~x560 & ~x561 & ~x585 & ~x588 & ~x591 & ~x613 & ~x615 & ~x617 & ~x618 & ~x619 & ~x637 & ~x640 & ~x642 & ~x644 & ~x646 & ~x648 & ~x649 & ~x665 & ~x666 & ~x670 & ~x671 & ~x672 & ~x673 & ~x674 & ~x690 & ~x691 & ~x692 & ~x693 & ~x697 & ~x699 & ~x702 & ~x704 & ~x711 & ~x715 & ~x716 & ~x718 & ~x726 & ~x727 & ~x732 & ~x733 & ~x734 & ~x735 & ~x737 & ~x739 & ~x742 & ~x745 & ~x746 & ~x749 & ~x753 & ~x756 & ~x758 & ~x759 & ~x760 & ~x762 & ~x763 & ~x764 & ~x766 & ~x767 & ~x768 & ~x770 & ~x772 & ~x773 & ~x774 & ~x778 & ~x781 & ~x782;
assign c556 =  x158 &  x187 & ~x0 & ~x1 & ~x5 & ~x6 & ~x7 & ~x8 & ~x9 & ~x11 & ~x12 & ~x13 & ~x14 & ~x16 & ~x18 & ~x19 & ~x21 & ~x22 & ~x23 & ~x24 & ~x25 & ~x27 & ~x28 & ~x31 & ~x32 & ~x33 & ~x34 & ~x35 & ~x36 & ~x38 & ~x39 & ~x41 & ~x42 & ~x43 & ~x44 & ~x45 & ~x47 & ~x49 & ~x50 & ~x52 & ~x53 & ~x56 & ~x58 & ~x59 & ~x60 & ~x62 & ~x64 & ~x65 & ~x66 & ~x67 & ~x68 & ~x69 & ~x70 & ~x71 & ~x72 & ~x74 & ~x75 & ~x76 & ~x77 & ~x81 & ~x84 & ~x85 & ~x86 & ~x87 & ~x88 & ~x89 & ~x90 & ~x91 & ~x92 & ~x93 & ~x94 & ~x95 & ~x96 & ~x97 & ~x98 & ~x100 & ~x101 & ~x102 & ~x103 & ~x104 & ~x105 & ~x106 & ~x107 & ~x108 & ~x109 & ~x110 & ~x111 & ~x112 & ~x113 & ~x115 & ~x116 & ~x118 & ~x119 & ~x121 & ~x138 & ~x139 & ~x140 & ~x141 & ~x143 & ~x144 & ~x145 & ~x147 & ~x166 & ~x168 & ~x169 & ~x170 & ~x172 & ~x173 & ~x174 & ~x193 & ~x194 & ~x196 & ~x197 & ~x199 & ~x200 & ~x219 & ~x223 & ~x224 & ~x225 & ~x226 & ~x227 & ~x228 & ~x229 & ~x242 & ~x243 & ~x244 & ~x245 & ~x247 & ~x248 & ~x249 & ~x250 & ~x251 & ~x256 & ~x271 & ~x272 & ~x273 & ~x274 & ~x275 & ~x277 & ~x278 & ~x279 & ~x280 & ~x281 & ~x282 & ~x283 & ~x284 & ~x285 & ~x300 & ~x301 & ~x302 & ~x303 & ~x304 & ~x305 & ~x308 & ~x310 & ~x311 & ~x313 & ~x331 & ~x332 & ~x333 & ~x334 & ~x335 & ~x336 & ~x339 & ~x340 & ~x360 & ~x362 & ~x363 & ~x364 & ~x366 & ~x367 & ~x387 & ~x390 & ~x391 & ~x392 & ~x393 & ~x394 & ~x395 & ~x396 & ~x416 & ~x417 & ~x418 & ~x419 & ~x421 & ~x422 & ~x423 & ~x424 & ~x425 & ~x444 & ~x445 & ~x446 & ~x447 & ~x450 & ~x474 & ~x475 & ~x477 & ~x479 & ~x501 & ~x503 & ~x504 & ~x505 & ~x506 & ~x528 & ~x530 & ~x532 & ~x533 & ~x534 & ~x535 & ~x556 & ~x557 & ~x558 & ~x559 & ~x562 & ~x563 & ~x585 & ~x586 & ~x587 & ~x588 & ~x589 & ~x590 & ~x591 & ~x611 & ~x613 & ~x614 & ~x615 & ~x616 & ~x617 & ~x618 & ~x639 & ~x640 & ~x641 & ~x643 & ~x644 & ~x645 & ~x646 & ~x647 & ~x648 & ~x649 & ~x665 & ~x666 & ~x667 & ~x669 & ~x670 & ~x671 & ~x672 & ~x673 & ~x674 & ~x675 & ~x678 & ~x692 & ~x694 & ~x695 & ~x696 & ~x697 & ~x698 & ~x699 & ~x700 & ~x701 & ~x702 & ~x703 & ~x704 & ~x705 & ~x706 & ~x707 & ~x712 & ~x713 & ~x714 & ~x718 & ~x719 & ~x720 & ~x721 & ~x723 & ~x724 & ~x727 & ~x731 & ~x732 & ~x733 & ~x734 & ~x737 & ~x739 & ~x741 & ~x742 & ~x743 & ~x744 & ~x746 & ~x747 & ~x748 & ~x749 & ~x750 & ~x751 & ~x752 & ~x753 & ~x754 & ~x755 & ~x756 & ~x758 & ~x759 & ~x760 & ~x761 & ~x762 & ~x764 & ~x765 & ~x766 & ~x767 & ~x768 & ~x770 & ~x771 & ~x773 & ~x774 & ~x775 & ~x776 & ~x777 & ~x778 & ~x779 & ~x780 & ~x781 & ~x782 & ~x783;
assign c558 = ~x1 & ~x2 & ~x7 & ~x8 & ~x10 & ~x11 & ~x13 & ~x14 & ~x15 & ~x16 & ~x17 & ~x18 & ~x19 & ~x20 & ~x22 & ~x23 & ~x25 & ~x27 & ~x29 & ~x30 & ~x31 & ~x32 & ~x35 & ~x36 & ~x37 & ~x38 & ~x39 & ~x42 & ~x43 & ~x44 & ~x46 & ~x47 & ~x48 & ~x50 & ~x51 & ~x54 & ~x55 & ~x56 & ~x58 & ~x59 & ~x60 & ~x61 & ~x64 & ~x67 & ~x71 & ~x72 & ~x73 & ~x74 & ~x78 & ~x79 & ~x80 & ~x81 & ~x82 & ~x83 & ~x84 & ~x88 & ~x89 & ~x90 & ~x92 & ~x93 & ~x94 & ~x97 & ~x98 & ~x99 & ~x100 & ~x101 & ~x105 & ~x107 & ~x108 & ~x109 & ~x110 & ~x111 & ~x112 & ~x113 & ~x114 & ~x115 & ~x137 & ~x138 & ~x139 & ~x140 & ~x141 & ~x142 & ~x143 & ~x144 & ~x145 & ~x146 & ~x164 & ~x165 & ~x168 & ~x169 & ~x171 & ~x172 & ~x192 & ~x198 & ~x199 & ~x200 & ~x221 & ~x222 & ~x223 & ~x224 & ~x225 & ~x227 & ~x228 & ~x247 & ~x249 & ~x251 & ~x253 & ~x255 & ~x256 & ~x277 & ~x278 & ~x284 & ~x293 & ~x294 & ~x295 & ~x296 & ~x297 & ~x298 & ~x299 & ~x300 & ~x301 & ~x302 & ~x305 & ~x306 & ~x308 & ~x309 & ~x310 & ~x334 & ~x335 & ~x336 & ~x337 & ~x339 & ~x360 & ~x362 & ~x363 & ~x366 & ~x367 & ~x389 & ~x390 & ~x391 & ~x392 & ~x393 & ~x394 & ~x395 & ~x418 & ~x419 & ~x420 & ~x421 & ~x422 & ~x446 & ~x447 & ~x449 & ~x480 & ~x492 & ~x502 & ~x503 & ~x504 & ~x507 & ~x517 & ~x518 & ~x519 & ~x520 & ~x529 & ~x532 & ~x536 & ~x545 & ~x558 & ~x562 & ~x563 & ~x585 & ~x587 & ~x588 & ~x589 & ~x590 & ~x591 & ~x613 & ~x615 & ~x616 & ~x618 & ~x619 & ~x620 & ~x622 & ~x645 & ~x646 & ~x649 & ~x666 & ~x667 & ~x668 & ~x670 & ~x671 & ~x672 & ~x675 & ~x689 & ~x693 & ~x694 & ~x695 & ~x698 & ~x700 & ~x702 & ~x703 & ~x705 & ~x706 & ~x707 & ~x708 & ~x709 & ~x710 & ~x712 & ~x714 & ~x717 & ~x718 & ~x721 & ~x722 & ~x727 & ~x728 & ~x730 & ~x731 & ~x732 & ~x733 & ~x734 & ~x736 & ~x737 & ~x739 & ~x742 & ~x743 & ~x746 & ~x751 & ~x752 & ~x755 & ~x756 & ~x758 & ~x759 & ~x761 & ~x763 & ~x764 & ~x765 & ~x766 & ~x767 & ~x768 & ~x771 & ~x773 & ~x774 & ~x775 & ~x776 & ~x777 & ~x779 & ~x781 & ~x783;
assign c560 = ~x14 & ~x26 & ~x44 & ~x48 & ~x59 & ~x72 & ~x79 & ~x82 & ~x98 & ~x116 & ~x122 & ~x139 & ~x148 & ~x149 & ~x151 & ~x155 & ~x168 & ~x171 & ~x178 & ~x202 & ~x232 & ~x236 & ~x255 & ~x257 & ~x259 & ~x282 & ~x284 & ~x286 & ~x308 & ~x311 & ~x343 & ~x369 & ~x397 & ~x414 & ~x442 & ~x445 & ~x458 & ~x478 & ~x524 & ~x530 & ~x531 & ~x534 & ~x588 & ~x609 & ~x642 & ~x661 & ~x670 & ~x671 & ~x690 & ~x699 & ~x712 & ~x713 & ~x714 & ~x720 & ~x722 & ~x737 & ~x742 & ~x762 & ~x765 & ~x766 & ~x781;
assign c562 = ~x6 & ~x14 & ~x22 & ~x33 & ~x36 & ~x51 & ~x54 & ~x64 & ~x74 & ~x75 & ~x83 & ~x101 & ~x115 & ~x117 & ~x132 & ~x135 & ~x145 & ~x148 & ~x156 & ~x158 & ~x159 & ~x161 & ~x162 & ~x163 & ~x174 & ~x183 & ~x184 & ~x185 & ~x186 & ~x187 & ~x210 & ~x211 & ~x212 & ~x222 & ~x228 & ~x231 & ~x255 & ~x258 & ~x280 & ~x285 & ~x287 & ~x288 & ~x308 & ~x314 & ~x364 & ~x365 & ~x383 & ~x392 & ~x393 & ~x412 & ~x413 & ~x415 & ~x441 & ~x474 & ~x476 & ~x496 & ~x556 & ~x590 & ~x591 & ~x611 & ~x612 & ~x638 & ~x640 & ~x661 & ~x663 & ~x668 & ~x695 & ~x696 & ~x698 & ~x717 & ~x719 & ~x732 & ~x736 & ~x740 & ~x741 & ~x742 & ~x743 & ~x747 & ~x753 & ~x758 & ~x772 & ~x782 & ~x783;
assign c564 =  x216 & ~x2 & ~x3 & ~x21 & ~x44 & ~x72 & ~x96 & ~x134 & ~x139 & ~x146 & ~x171 & ~x299 & ~x300 & ~x302 & ~x325 & ~x327 & ~x328 & ~x355 & ~x357 & ~x360 & ~x361 & ~x388 & ~x394 & ~x413 & ~x414 & ~x584 & ~x741 & ~x754 & ~x764 & ~x769;
assign c566 =  x177 &  x205 &  x206 &  x289 & ~x2 & ~x7 & ~x10 & ~x11 & ~x16 & ~x21 & ~x29 & ~x33 & ~x36 & ~x42 & ~x43 & ~x48 & ~x50 & ~x54 & ~x55 & ~x57 & ~x59 & ~x60 & ~x71 & ~x74 & ~x75 & ~x79 & ~x83 & ~x84 & ~x85 & ~x90 & ~x91 & ~x92 & ~x100 & ~x102 & ~x106 & ~x107 & ~x109 & ~x110 & ~x112 & ~x114 & ~x118 & ~x133 & ~x134 & ~x139 & ~x164 & ~x165 & ~x195 & ~x198 & ~x220 & ~x221 & ~x223 & ~x227 & ~x228 & ~x250 & ~x254 & ~x278 & ~x279 & ~x281 & ~x283 & ~x303 & ~x307 & ~x309 & ~x330 & ~x333 & ~x334 & ~x361 & ~x364 & ~x367 & ~x388 & ~x390 & ~x420 & ~x422 & ~x423 & ~x425 & ~x444 & ~x445 & ~x449 & ~x450 & ~x453 & ~x454 & ~x475 & ~x476 & ~x478 & ~x479 & ~x481 & ~x483 & ~x502 & ~x507 & ~x510 & ~x516 & ~x518 & ~x519 & ~x528 & ~x556 & ~x558 & ~x561 & ~x584 & ~x585 & ~x588 & ~x616 & ~x645 & ~x669 & ~x672 & ~x673 & ~x674 & ~x676 & ~x696 & ~x697 & ~x703 & ~x707 & ~x708 & ~x722 & ~x727 & ~x731 & ~x738 & ~x740 & ~x745 & ~x748 & ~x752 & ~x758 & ~x760 & ~x762 & ~x765 & ~x768 & ~x772 & ~x776 & ~x777 & ~x779 & ~x783;
assign c568 =  x169;
assign c570 =  x305;
assign c572 =  x20;
assign c574 =  x699;
assign c576 =  x232 &  x609 & ~x37 & ~x270 & ~x272 & ~x301 & ~x302 & ~x360 & ~x466 & ~x489 & ~x518 & ~x548 & ~x549;
assign c578 =  x627 & ~x0 & ~x8 & ~x20 & ~x21 & ~x24 & ~x26 & ~x27 & ~x41 & ~x43 & ~x44 & ~x45 & ~x48 & ~x51 & ~x56 & ~x68 & ~x73 & ~x75 & ~x79 & ~x82 & ~x84 & ~x87 & ~x91 & ~x93 & ~x94 & ~x109 & ~x112 & ~x116 & ~x120 & ~x140 & ~x150 & ~x167 & ~x177 & ~x197 & ~x201 & ~x203 & ~x220 & ~x222 & ~x223 & ~x225 & ~x243 & ~x244 & ~x246 & ~x247 & ~x249 & ~x250 & ~x252 & ~x268 & ~x269 & ~x270 & ~x271 & ~x277 & ~x278 & ~x279 & ~x282 & ~x286 & ~x298 & ~x299 & ~x312 & ~x328 & ~x330 & ~x331 & ~x332 & ~x333 & ~x335 & ~x336 & ~x343 & ~x357 & ~x362 & ~x365 & ~x370 & ~x395 & ~x416 & ~x418 & ~x420 & ~x421 & ~x424 & ~x443 & ~x447 & ~x448 & ~x450 & ~x454 & ~x455 & ~x456 & ~x457 & ~x471 & ~x475 & ~x501 & ~x502 & ~x506 & ~x532 & ~x557 & ~x560 & ~x581 & ~x584 & ~x608 & ~x609 & ~x615 & ~x634 & ~x636 & ~x641 & ~x644 & ~x647 & ~x663 & ~x668 & ~x670 & ~x671 & ~x675 & ~x689 & ~x693 & ~x699 & ~x703 & ~x704 & ~x707 & ~x708 & ~x711 & ~x715 & ~x722 & ~x725 & ~x726 & ~x730 & ~x731 & ~x732 & ~x741 & ~x742 & ~x743 & ~x745 & ~x748 & ~x755 & ~x756 & ~x757 & ~x763 & ~x770 & ~x774;
assign c580 =  x163 & ~x271 & ~x272;
assign c582 =  x214 & ~x0 & ~x1 & ~x2 & ~x4 & ~x5 & ~x6 & ~x8 & ~x12 & ~x13 & ~x14 & ~x15 & ~x16 & ~x18 & ~x21 & ~x22 & ~x23 & ~x26 & ~x29 & ~x30 & ~x34 & ~x38 & ~x39 & ~x40 & ~x43 & ~x47 & ~x49 & ~x50 & ~x51 & ~x53 & ~x54 & ~x55 & ~x56 & ~x60 & ~x61 & ~x62 & ~x63 & ~x65 & ~x68 & ~x69 & ~x70 & ~x71 & ~x72 & ~x75 & ~x80 & ~x83 & ~x84 & ~x85 & ~x87 & ~x88 & ~x89 & ~x93 & ~x97 & ~x100 & ~x103 & ~x105 & ~x106 & ~x107 & ~x108 & ~x112 & ~x114 & ~x115 & ~x116 & ~x122 & ~x124 & ~x125 & ~x126 & ~x127 & ~x135 & ~x138 & ~x143 & ~x144 & ~x145 & ~x164 & ~x167 & ~x169 & ~x173 & ~x175 & ~x193 & ~x194 & ~x196 & ~x201 & ~x202 & ~x223 & ~x226 & ~x251 & ~x253 & ~x256 & ~x278 & ~x286 & ~x297 & ~x299 & ~x300 & ~x301 & ~x305 & ~x306 & ~x311 & ~x312 & ~x313 & ~x327 & ~x331 & ~x334 & ~x339 & ~x340 & ~x341 & ~x356 & ~x358 & ~x359 & ~x360 & ~x362 & ~x363 & ~x364 & ~x366 & ~x385 & ~x390 & ~x393 & ~x395 & ~x396 & ~x397 & ~x398 & ~x413 & ~x417 & ~x423 & ~x443 & ~x446 & ~x448 & ~x450 & ~x470 & ~x472 & ~x475 & ~x477 & ~x499 & ~x502 & ~x503 & ~x504 & ~x505 & ~x526 & ~x531 & ~x558 & ~x560 & ~x562 & ~x582 & ~x583 & ~x584 & ~x585 & ~x586 & ~x590 & ~x610 & ~x614 & ~x615 & ~x617 & ~x640 & ~x641 & ~x642 & ~x646 & ~x647 & ~x668 & ~x669 & ~x670 & ~x675 & ~x677 & ~x695 & ~x699 & ~x703 & ~x704 & ~x720 & ~x721 & ~x722 & ~x725 & ~x728 & ~x730 & ~x734 & ~x736 & ~x742 & ~x743 & ~x746 & ~x747 & ~x749 & ~x750 & ~x751 & ~x755 & ~x757 & ~x759 & ~x761 & ~x762 & ~x767 & ~x768 & ~x770 & ~x776 & ~x778;
assign c584 =  x288 &  x344 &  x632 & ~x21 & ~x42 & ~x46 & ~x51 & ~x101 & ~x106 & ~x108 & ~x112 & ~x118 & ~x120 & ~x141 & ~x145 & ~x220 & ~x228 & ~x256 & ~x280 & ~x307 & ~x362 & ~x366 & ~x388 & ~x449 & ~x454 & ~x485 & ~x503 & ~x533 & ~x611 & ~x692 & ~x700 & ~x724 & ~x740 & ~x741 & ~x749 & ~x778;
assign c586 = ~x218 & ~x243 & ~x245 & ~x401 & ~x456 & ~x457 & ~x458 & ~x486;
assign c588 = ~x0 & ~x1 & ~x2 & ~x3 & ~x4 & ~x5 & ~x6 & ~x7 & ~x8 & ~x11 & ~x13 & ~x14 & ~x15 & ~x17 & ~x18 & ~x19 & ~x21 & ~x22 & ~x23 & ~x24 & ~x25 & ~x26 & ~x27 & ~x28 & ~x29 & ~x30 & ~x31 & ~x32 & ~x33 & ~x34 & ~x35 & ~x36 & ~x37 & ~x38 & ~x39 & ~x40 & ~x41 & ~x42 & ~x43 & ~x44 & ~x45 & ~x47 & ~x48 & ~x49 & ~x50 & ~x51 & ~x53 & ~x54 & ~x55 & ~x57 & ~x58 & ~x60 & ~x61 & ~x62 & ~x63 & ~x64 & ~x65 & ~x66 & ~x68 & ~x69 & ~x73 & ~x74 & ~x75 & ~x76 & ~x78 & ~x79 & ~x80 & ~x81 & ~x82 & ~x83 & ~x85 & ~x86 & ~x88 & ~x89 & ~x90 & ~x91 & ~x92 & ~x94 & ~x95 & ~x96 & ~x99 & ~x107 & ~x110 & ~x111 & ~x112 & ~x113 & ~x115 & ~x116 & ~x117 & ~x119 & ~x120 & ~x122 & ~x137 & ~x138 & ~x139 & ~x140 & ~x141 & ~x143 & ~x144 & ~x145 & ~x147 & ~x165 & ~x166 & ~x167 & ~x168 & ~x169 & ~x170 & ~x171 & ~x172 & ~x173 & ~x174 & ~x193 & ~x194 & ~x195 & ~x196 & ~x197 & ~x198 & ~x201 & ~x218 & ~x219 & ~x220 & ~x223 & ~x225 & ~x226 & ~x228 & ~x243 & ~x244 & ~x245 & ~x246 & ~x247 & ~x248 & ~x249 & ~x250 & ~x251 & ~x252 & ~x253 & ~x254 & ~x258 & ~x271 & ~x272 & ~x273 & ~x274 & ~x275 & ~x277 & ~x279 & ~x280 & ~x281 & ~x282 & ~x283 & ~x284 & ~x285 & ~x286 & ~x300 & ~x301 & ~x302 & ~x303 & ~x304 & ~x305 & ~x307 & ~x308 & ~x309 & ~x310 & ~x311 & ~x330 & ~x331 & ~x332 & ~x333 & ~x334 & ~x335 & ~x336 & ~x337 & ~x338 & ~x340 & ~x359 & ~x360 & ~x361 & ~x363 & ~x366 & ~x367 & ~x389 & ~x390 & ~x391 & ~x392 & ~x395 & ~x419 & ~x420 & ~x421 & ~x422 & ~x424 & ~x431 & ~x432 & ~x433 & ~x434 & ~x443 & ~x445 & ~x446 & ~x447 & ~x448 & ~x450 & ~x458 & ~x459 & ~x461 & ~x462 & ~x473 & ~x475 & ~x476 & ~x478 & ~x488 & ~x500 & ~x501 & ~x502 & ~x503 & ~x505 & ~x506 & ~x528 & ~x529 & ~x530 & ~x531 & ~x533 & ~x534 & ~x535 & ~x556 & ~x557 & ~x559 & ~x560 & ~x561 & ~x562 & ~x583 & ~x585 & ~x589 & ~x590 & ~x611 & ~x612 & ~x613 & ~x615 & ~x616 & ~x617 & ~x618 & ~x619 & ~x637 & ~x639 & ~x641 & ~x643 & ~x646 & ~x647 & ~x648 & ~x668 & ~x669 & ~x670 & ~x672 & ~x673 & ~x674 & ~x675 & ~x676 & ~x677 & ~x689 & ~x691 & ~x692 & ~x693 & ~x694 & ~x695 & ~x696 & ~x698 & ~x699 & ~x701 & ~x702 & ~x703 & ~x704 & ~x705 & ~x706 & ~x707 & ~x708 & ~x709 & ~x710 & ~x713 & ~x715 & ~x716 & ~x717 & ~x720 & ~x721 & ~x722 & ~x723 & ~x724 & ~x725 & ~x726 & ~x727 & ~x728 & ~x730 & ~x731 & ~x732 & ~x734 & ~x735 & ~x736 & ~x737 & ~x738 & ~x739 & ~x740 & ~x741 & ~x742 & ~x743 & ~x744 & ~x745 & ~x746 & ~x747 & ~x748 & ~x749 & ~x750 & ~x751 & ~x752 & ~x753 & ~x754 & ~x756 & ~x757 & ~x758 & ~x759 & ~x761 & ~x763 & ~x764 & ~x765 & ~x766 & ~x767 & ~x768 & ~x769 & ~x770 & ~x771 & ~x772 & ~x773 & ~x774 & ~x775 & ~x776 & ~x777 & ~x778 & ~x781 & ~x782 & ~x783;
assign c590 = ~x2 & ~x7 & ~x15 & ~x16 & ~x24 & ~x25 & ~x28 & ~x33 & ~x37 & ~x44 & ~x46 & ~x49 & ~x51 & ~x72 & ~x86 & ~x95 & ~x105 & ~x107 & ~x116 & ~x119 & ~x144 & ~x145 & ~x176 & ~x195 & ~x225 & ~x226 & ~x231 & ~x250 & ~x254 & ~x255 & ~x258 & ~x313 & ~x323 & ~x328 & ~x331 & ~x335 & ~x340 & ~x354 & ~x362 & ~x382 & ~x389 & ~x396 & ~x413 & ~x414 & ~x417 & ~x444 & ~x469 & ~x476 & ~x478 & ~x499 & ~x503 & ~x505 & ~x510 & ~x513 & ~x514 & ~x526 & ~x543 & ~x544 & ~x553 & ~x560 & ~x562 & ~x563 & ~x566 & ~x582 & ~x584 & ~x593 & ~x614 & ~x616 & ~x642 & ~x666 & ~x668 & ~x693 & ~x701 & ~x723 & ~x732 & ~x745 & ~x746 & ~x747 & ~x749 & ~x750 & ~x767 & ~x772 & ~x773 & ~x778;
assign c592 =  x203 &  x286 &  x314 &  x583;
assign c594 =  x295 &  x296 &  x297 & ~x98 & ~x154 & ~x159 & ~x165 & ~x187 & ~x285 & ~x313 & ~x356 & ~x388 & ~x413 & ~x472 & ~x498 & ~x554;
assign c596 =  x212 &  x236 &  x377 & ~x1 & ~x14 & ~x18 & ~x19 & ~x25 & ~x35 & ~x36 & ~x39 & ~x45 & ~x49 & ~x52 & ~x56 & ~x60 & ~x61 & ~x62 & ~x69 & ~x72 & ~x74 & ~x77 & ~x82 & ~x90 & ~x92 & ~x100 & ~x110 & ~x114 & ~x118 & ~x121 & ~x136 & ~x145 & ~x169 & ~x195 & ~x228 & ~x249 & ~x250 & ~x278 & ~x280 & ~x295 & ~x296 & ~x297 & ~x329 & ~x330 & ~x334 & ~x387 & ~x392 & ~x394 & ~x416 & ~x420 & ~x450 & ~x478 & ~x501 & ~x533 & ~x534 & ~x587 & ~x619 & ~x643 & ~x645 & ~x666 & ~x696 & ~x698 & ~x721 & ~x724 & ~x725 & ~x727 & ~x729 & ~x734 & ~x742 & ~x743 & ~x745 & ~x753 & ~x759 & ~x776 & ~x779 & ~x781 & ~x783;
assign c598 =  x272 & ~x7 & ~x11 & ~x65 & ~x101 & ~x128 & ~x133 & ~x158 & ~x353 & ~x355 & ~x356 & ~x383 & ~x413 & ~x441 & ~x554 & ~x586 & ~x780;
assign c5100 =  x265 &  x293 & ~x0 & ~x5 & ~x6 & ~x24 & ~x39 & ~x59 & ~x60 & ~x63 & ~x65 & ~x70 & ~x85 & ~x92 & ~x93 & ~x116 & ~x141 & ~x150 & ~x168 & ~x192 & ~x195 & ~x220 & ~x221 & ~x227 & ~x228 & ~x229 & ~x254 & ~x260 & ~x262 & ~x287 & ~x305 & ~x314 & ~x329 & ~x337 & ~x341 & ~x363 & ~x371 & ~x389 & ~x393 & ~x398 & ~x420 & ~x428 & ~x442 & ~x445 & ~x448 & ~x449 & ~x451 & ~x478 & ~x515 & ~x517 & ~x526 & ~x532 & ~x554 & ~x557 & ~x579 & ~x583 & ~x607 & ~x613 & ~x616 & ~x637 & ~x641 & ~x661 & ~x662 & ~x664 & ~x669 & ~x697 & ~x699 & ~x700 & ~x711 & ~x712 & ~x716 & ~x720 & ~x732 & ~x751 & ~x762 & ~x770 & ~x773 & ~x774 & ~x777;
assign c5102 =  x377 &  x379 & ~x3 & ~x8 & ~x19 & ~x33 & ~x36 & ~x40 & ~x41 & ~x43 & ~x48 & ~x49 & ~x50 & ~x52 & ~x58 & ~x63 & ~x64 & ~x66 & ~x67 & ~x73 & ~x78 & ~x91 & ~x92 & ~x111 & ~x113 & ~x137 & ~x138 & ~x140 & ~x143 & ~x145 & ~x165 & ~x167 & ~x169 & ~x170 & ~x174 & ~x193 & ~x198 & ~x227 & ~x228 & ~x250 & ~x266 & ~x267 & ~x268 & ~x269 & ~x276 & ~x278 & ~x279 & ~x282 & ~x297 & ~x298 & ~x300 & ~x301 & ~x302 & ~x305 & ~x334 & ~x336 & ~x339 & ~x390 & ~x392 & ~x396 & ~x418 & ~x422 & ~x447 & ~x459 & ~x461 & ~x462 & ~x476 & ~x479 & ~x490 & ~x504 & ~x506 & ~x559 & ~x560 & ~x561 & ~x587 & ~x588 & ~x614 & ~x643 & ~x645 & ~x667 & ~x668 & ~x670 & ~x694 & ~x696 & ~x697 & ~x699 & ~x705 & ~x713 & ~x717 & ~x718 & ~x720 & ~x722 & ~x728 & ~x729 & ~x736 & ~x738 & ~x739 & ~x749 & ~x750 & ~x762 & ~x764 & ~x769 & ~x775 & ~x776 & ~x778 & ~x781;
assign c5104 =  x215 & ~x0 & ~x2 & ~x5 & ~x6 & ~x17 & ~x20 & ~x25 & ~x31 & ~x35 & ~x36 & ~x39 & ~x51 & ~x54 & ~x61 & ~x67 & ~x71 & ~x74 & ~x82 & ~x86 & ~x94 & ~x96 & ~x101 & ~x103 & ~x107 & ~x113 & ~x119 & ~x122 & ~x130 & ~x131 & ~x136 & ~x144 & ~x170 & ~x226 & ~x257 & ~x279 & ~x281 & ~x282 & ~x296 & ~x299 & ~x301 & ~x331 & ~x339 & ~x357 & ~x358 & ~x366 & ~x368 & ~x392 & ~x395 & ~x418 & ~x422 & ~x445 & ~x472 & ~x500 & ~x502 & ~x504 & ~x544 & ~x563 & ~x587 & ~x590 & ~x613 & ~x614 & ~x641 & ~x646 & ~x648 & ~x669 & ~x675 & ~x699 & ~x700 & ~x725 & ~x726 & ~x729 & ~x731 & ~x742 & ~x744 & ~x747 & ~x751 & ~x752 & ~x756 & ~x779 & ~x780;
assign c5106 =  x597 &  x600 &  x601 &  x627 & ~x7 & ~x8 & ~x23 & ~x35 & ~x57 & ~x72 & ~x82 & ~x94 & ~x97 & ~x113 & ~x123 & ~x145 & ~x148 & ~x149 & ~x150 & ~x175 & ~x193 & ~x198 & ~x259 & ~x280 & ~x284 & ~x301 & ~x302 & ~x306 & ~x307 & ~x315 & ~x330 & ~x334 & ~x335 & ~x342 & ~x359 & ~x363 & ~x369 & ~x397 & ~x399 & ~x421 & ~x423 & ~x429 & ~x449 & ~x460 & ~x503 & ~x506 & ~x535 & ~x563 & ~x584 & ~x588 & ~x591 & ~x619 & ~x676 & ~x688 & ~x693 & ~x696 & ~x735 & ~x739 & ~x748 & ~x753 & ~x770 & ~x781;
assign c5108 =  x295;
assign c5110 =  x186 &  x210 &  x211 &  x236 &  x263 &  x346 &  x630 &  x632 & ~x7 & ~x8 & ~x15 & ~x30 & ~x37 & ~x41 & ~x44 & ~x56 & ~x58 & ~x60 & ~x61 & ~x65 & ~x67 & ~x73 & ~x85 & ~x96 & ~x115 & ~x228 & ~x248 & ~x277 & ~x279 & ~x330 & ~x331 & ~x336 & ~x360 & ~x387 & ~x388 & ~x450 & ~x476 & ~x479 & ~x510 & ~x511 & ~x529 & ~x584 & ~x614 & ~x669 & ~x716 & ~x722 & ~x730 & ~x731 & ~x741 & ~x755 & ~x759 & ~x760 & ~x782;
assign c5112 =  x209 &  x210 &  x236 &  x292 & ~x3 & ~x10 & ~x14 & ~x15 & ~x43 & ~x49 & ~x50 & ~x66 & ~x71 & ~x85 & ~x94 & ~x124 & ~x140 & ~x142 & ~x143 & ~x144 & ~x193 & ~x196 & ~x202 & ~x204 & ~x228 & ~x230 & ~x231 & ~x232 & ~x249 & ~x250 & ~x256 & ~x257 & ~x260 & ~x281 & ~x282 & ~x285 & ~x305 & ~x312 & ~x331 & ~x339 & ~x341 & ~x358 & ~x361 & ~x369 & ~x387 & ~x391 & ~x414 & ~x421 & ~x472 & ~x474 & ~x478 & ~x490 & ~x491 & ~x499 & ~x502 & ~x505 & ~x530 & ~x533 & ~x535 & ~x553 & ~x555 & ~x588 & ~x589 & ~x608 & ~x609 & ~x617 & ~x637 & ~x638 & ~x645 & ~x669 & ~x674 & ~x677 & ~x692 & ~x694 & ~x697 & ~x700 & ~x702 & ~x725 & ~x730 & ~x734 & ~x740 & ~x743 & ~x746 & ~x753 & ~x762 & ~x770 & ~x771 & ~x780;
assign c5114 = ~x7 & ~x11 & ~x21 & ~x37 & ~x40 & ~x44 & ~x48 & ~x56 & ~x72 & ~x74 & ~x76 & ~x81 & ~x84 & ~x91 & ~x92 & ~x145 & ~x146 & ~x170 & ~x200 & ~x226 & ~x227 & ~x228 & ~x250 & ~x253 & ~x276 & ~x277 & ~x280 & ~x281 & ~x294 & ~x296 & ~x298 & ~x301 & ~x324 & ~x325 & ~x327 & ~x330 & ~x335 & ~x357 & ~x360 & ~x361 & ~x365 & ~x389 & ~x415 & ~x419 & ~x447 & ~x472 & ~x478 & ~x499 & ~x501 & ~x513 & ~x515 & ~x516 & ~x545 & ~x547 & ~x557 & ~x560 & ~x613 & ~x617 & ~x643 & ~x646 & ~x669 & ~x671 & ~x677 & ~x697 & ~x698 & ~x723 & ~x726 & ~x727 & ~x729 & ~x738 & ~x741 & ~x749 & ~x754 & ~x756 & ~x758 & ~x759 & ~x761;
assign c5116 =  x209 &  x211 &  x212 & ~x3 & ~x10 & ~x12 & ~x17 & ~x23 & ~x26 & ~x34 & ~x35 & ~x36 & ~x41 & ~x43 & ~x46 & ~x47 & ~x50 & ~x51 & ~x53 & ~x54 & ~x55 & ~x56 & ~x60 & ~x62 & ~x63 & ~x64 & ~x65 & ~x71 & ~x76 & ~x82 & ~x83 & ~x88 & ~x89 & ~x91 & ~x92 & ~x95 & ~x96 & ~x98 & ~x99 & ~x104 & ~x105 & ~x108 & ~x111 & ~x112 & ~x115 & ~x118 & ~x120 & ~x128 & ~x136 & ~x138 & ~x140 & ~x141 & ~x142 & ~x166 & ~x168 & ~x172 & ~x173 & ~x193 & ~x199 & ~x200 & ~x223 & ~x224 & ~x226 & ~x253 & ~x255 & ~x276 & ~x277 & ~x279 & ~x280 & ~x297 & ~x298 & ~x300 & ~x301 & ~x302 & ~x309 & ~x328 & ~x329 & ~x332 & ~x333 & ~x357 & ~x361 & ~x387 & ~x390 & ~x418 & ~x419 & ~x421 & ~x444 & ~x446 & ~x450 & ~x453 & ~x473 & ~x476 & ~x477 & ~x480 & ~x504 & ~x505 & ~x509 & ~x517 & ~x518 & ~x519 & ~x528 & ~x529 & ~x530 & ~x533 & ~x534 & ~x536 & ~x546 & ~x556 & ~x558 & ~x561 & ~x585 & ~x587 & ~x588 & ~x592 & ~x611 & ~x621 & ~x639 & ~x640 & ~x641 & ~x644 & ~x647 & ~x648 & ~x650 & ~x672 & ~x674 & ~x678 & ~x679 & ~x694 & ~x696 & ~x699 & ~x700 & ~x701 & ~x703 & ~x704 & ~x710 & ~x720 & ~x721 & ~x726 & ~x727 & ~x730 & ~x737 & ~x738 & ~x741 & ~x744 & ~x752 & ~x753 & ~x754 & ~x757 & ~x762 & ~x765 & ~x771 & ~x776 & ~x780 & ~x782 & ~x783;
assign c5118 = ~x4 & ~x5 & ~x7 & ~x10 & ~x11 & ~x12 & ~x14 & ~x16 & ~x17 & ~x18 & ~x19 & ~x20 & ~x21 & ~x22 & ~x23 & ~x24 & ~x27 & ~x32 & ~x33 & ~x34 & ~x36 & ~x39 & ~x44 & ~x48 & ~x50 & ~x51 & ~x52 & ~x59 & ~x61 & ~x62 & ~x66 & ~x69 & ~x72 & ~x73 & ~x77 & ~x79 & ~x82 & ~x84 & ~x85 & ~x88 & ~x89 & ~x92 & ~x98 & ~x100 & ~x101 & ~x104 & ~x112 & ~x113 & ~x118 & ~x133 & ~x140 & ~x141 & ~x144 & ~x163 & ~x171 & ~x173 & ~x192 & ~x193 & ~x197 & ~x199 & ~x223 & ~x224 & ~x229 & ~x239 & ~x240 & ~x241 & ~x242 & ~x243 & ~x244 & ~x245 & ~x253 & ~x254 & ~x255 & ~x271 & ~x272 & ~x274 & ~x280 & ~x283 & ~x301 & ~x302 & ~x306 & ~x307 & ~x310 & ~x330 & ~x332 & ~x335 & ~x339 & ~x359 & ~x362 & ~x364 & ~x365 & ~x366 & ~x389 & ~x392 & ~x396 & ~x397 & ~x398 & ~x415 & ~x416 & ~x417 & ~x422 & ~x445 & ~x446 & ~x464 & ~x474 & ~x477 & ~x491 & ~x492 & ~x503 & ~x504 & ~x505 & ~x506 & ~x516 & ~x518 & ~x529 & ~x544 & ~x545 & ~x546 & ~x561 & ~x589 & ~x590 & ~x593 & ~x611 & ~x614 & ~x615 & ~x616 & ~x617 & ~x618 & ~x621 & ~x622 & ~x638 & ~x646 & ~x648 & ~x649 & ~x650 & ~x651 & ~x665 & ~x666 & ~x669 & ~x670 & ~x672 & ~x673 & ~x677 & ~x679 & ~x680 & ~x681 & ~x696 & ~x697 & ~x699 & ~x700 & ~x701 & ~x704 & ~x706 & ~x719 & ~x720 & ~x724 & ~x727 & ~x730 & ~x731 & ~x732 & ~x739 & ~x742 & ~x743 & ~x747 & ~x750 & ~x754 & ~x757 & ~x758 & ~x759 & ~x765 & ~x766 & ~x767 & ~x768 & ~x772 & ~x774 & ~x780 & ~x781 & ~x782 & ~x783;
assign c5120 =  x657 & ~x0 & ~x2 & ~x12 & ~x20 & ~x22 & ~x34 & ~x51 & ~x61 & ~x66 & ~x68 & ~x81 & ~x96 & ~x99 & ~x101 & ~x106 & ~x107 & ~x144 & ~x145 & ~x172 & ~x198 & ~x216 & ~x224 & ~x227 & ~x239 & ~x240 & ~x241 & ~x243 & ~x246 & ~x255 & ~x279 & ~x301 & ~x303 & ~x306 & ~x308 & ~x365 & ~x367 & ~x368 & ~x389 & ~x393 & ~x418 & ~x436 & ~x446 & ~x488 & ~x489 & ~x506 & ~x516 & ~x520 & ~x534 & ~x535 & ~x547 & ~x559 & ~x564 & ~x612 & ~x613 & ~x618 & ~x649 & ~x650 & ~x672 & ~x701 & ~x708 & ~x710 & ~x712 & ~x718 & ~x724 & ~x727 & ~x734 & ~x735 & ~x743 & ~x759 & ~x761 & ~x765 & ~x774;
assign c5122 = ~x1 & ~x2 & ~x3 & ~x5 & ~x9 & ~x11 & ~x12 & ~x14 & ~x16 & ~x17 & ~x21 & ~x22 & ~x25 & ~x28 & ~x29 & ~x30 & ~x31 & ~x32 & ~x33 & ~x36 & ~x37 & ~x38 & ~x39 & ~x41 & ~x42 & ~x45 & ~x48 & ~x49 & ~x54 & ~x57 & ~x58 & ~x62 & ~x63 & ~x64 & ~x65 & ~x66 & ~x69 & ~x70 & ~x77 & ~x79 & ~x80 & ~x81 & ~x88 & ~x89 & ~x90 & ~x92 & ~x93 & ~x109 & ~x110 & ~x113 & ~x114 & ~x115 & ~x116 & ~x117 & ~x118 & ~x119 & ~x120 & ~x137 & ~x139 & ~x140 & ~x141 & ~x143 & ~x145 & ~x147 & ~x165 & ~x166 & ~x168 & ~x169 & ~x171 & ~x193 & ~x194 & ~x196 & ~x198 & ~x199 & ~x200 & ~x220 & ~x225 & ~x227 & ~x228 & ~x243 & ~x244 & ~x246 & ~x249 & ~x250 & ~x252 & ~x255 & ~x256 & ~x257 & ~x259 & ~x267 & ~x268 & ~x270 & ~x272 & ~x275 & ~x276 & ~x277 & ~x279 & ~x280 & ~x281 & ~x283 & ~x285 & ~x297 & ~x298 & ~x299 & ~x300 & ~x301 & ~x302 & ~x303 & ~x304 & ~x307 & ~x311 & ~x312 & ~x328 & ~x330 & ~x333 & ~x336 & ~x337 & ~x340 & ~x359 & ~x361 & ~x362 & ~x363 & ~x365 & ~x368 & ~x387 & ~x388 & ~x391 & ~x394 & ~x395 & ~x397 & ~x415 & ~x416 & ~x417 & ~x418 & ~x422 & ~x423 & ~x443 & ~x444 & ~x445 & ~x446 & ~x447 & ~x448 & ~x449 & ~x451 & ~x452 & ~x459 & ~x471 & ~x473 & ~x474 & ~x477 & ~x478 & ~x485 & ~x489 & ~x490 & ~x500 & ~x504 & ~x506 & ~x528 & ~x529 & ~x530 & ~x534 & ~x535 & ~x536 & ~x555 & ~x556 & ~x557 & ~x561 & ~x584 & ~x585 & ~x590 & ~x591 & ~x612 & ~x616 & ~x619 & ~x638 & ~x639 & ~x640 & ~x641 & ~x644 & ~x647 & ~x664 & ~x668 & ~x671 & ~x672 & ~x673 & ~x674 & ~x676 & ~x677 & ~x692 & ~x694 & ~x695 & ~x696 & ~x697 & ~x699 & ~x701 & ~x702 & ~x705 & ~x707 & ~x708 & ~x711 & ~x712 & ~x717 & ~x718 & ~x721 & ~x724 & ~x726 & ~x727 & ~x728 & ~x730 & ~x732 & ~x734 & ~x735 & ~x739 & ~x740 & ~x741 & ~x742 & ~x745 & ~x747 & ~x748 & ~x750 & ~x754 & ~x757 & ~x760 & ~x761 & ~x762 & ~x763 & ~x765 & ~x767 & ~x770 & ~x772 & ~x774 & ~x776 & ~x778 & ~x780 & ~x781 & ~x783;
assign c5124 = ~x2 & ~x15 & ~x16 & ~x17 & ~x19 & ~x20 & ~x24 & ~x27 & ~x32 & ~x38 & ~x50 & ~x54 & ~x56 & ~x67 & ~x74 & ~x81 & ~x84 & ~x91 & ~x103 & ~x106 & ~x108 & ~x110 & ~x120 & ~x134 & ~x136 & ~x138 & ~x141 & ~x159 & ~x162 & ~x164 & ~x169 & ~x198 & ~x254 & ~x276 & ~x280 & ~x281 & ~x282 & ~x292 & ~x293 & ~x296 & ~x298 & ~x299 & ~x300 & ~x301 & ~x303 & ~x310 & ~x325 & ~x326 & ~x330 & ~x331 & ~x337 & ~x360 & ~x389 & ~x390 & ~x392 & ~x393 & ~x395 & ~x420 & ~x446 & ~x447 & ~x448 & ~x479 & ~x481 & ~x489 & ~x501 & ~x503 & ~x518 & ~x519 & ~x529 & ~x531 & ~x532 & ~x546 & ~x557 & ~x562 & ~x585 & ~x587 & ~x591 & ~x615 & ~x620 & ~x642 & ~x647 & ~x648 & ~x671 & ~x678 & ~x700 & ~x701 & ~x704 & ~x708 & ~x727 & ~x733 & ~x734 & ~x737 & ~x740 & ~x741 & ~x742 & ~x754 & ~x757 & ~x760 & ~x762 & ~x764 & ~x775 & ~x776 & ~x777 & ~x781 & ~x782;
assign c5126 = ~x0 & ~x5 & ~x6 & ~x7 & ~x15 & ~x20 & ~x26 & ~x27 & ~x28 & ~x31 & ~x32 & ~x37 & ~x40 & ~x43 & ~x44 & ~x48 & ~x55 & ~x56 & ~x61 & ~x72 & ~x73 & ~x77 & ~x78 & ~x81 & ~x85 & ~x89 & ~x90 & ~x95 & ~x97 & ~x99 & ~x101 & ~x103 & ~x105 & ~x106 & ~x107 & ~x110 & ~x111 & ~x113 & ~x114 & ~x115 & ~x116 & ~x117 & ~x120 & ~x122 & ~x123 & ~x142 & ~x147 & ~x167 & ~x169 & ~x172 & ~x173 & ~x175 & ~x178 & ~x195 & ~x196 & ~x198 & ~x199 & ~x205 & ~x226 & ~x251 & ~x258 & ~x282 & ~x287 & ~x298 & ~x299 & ~x300 & ~x301 & ~x302 & ~x307 & ~x311 & ~x328 & ~x329 & ~x330 & ~x332 & ~x339 & ~x340 & ~x362 & ~x364 & ~x365 & ~x367 & ~x370 & ~x385 & ~x389 & ~x393 & ~x395 & ~x415 & ~x423 & ~x424 & ~x425 & ~x443 & ~x444 & ~x451 & ~x471 & ~x473 & ~x476 & ~x498 & ~x499 & ~x502 & ~x503 & ~x504 & ~x528 & ~x529 & ~x530 & ~x531 & ~x532 & ~x533 & ~x553 & ~x554 & ~x558 & ~x560 & ~x581 & ~x588 & ~x589 & ~x610 & ~x613 & ~x635 & ~x637 & ~x638 & ~x639 & ~x642 & ~x643 & ~x645 & ~x646 & ~x666 & ~x669 & ~x670 & ~x671 & ~x675 & ~x688 & ~x693 & ~x694 & ~x695 & ~x700 & ~x701 & ~x702 & ~x704 & ~x708 & ~x709 & ~x714 & ~x723 & ~x724 & ~x725 & ~x726 & ~x732 & ~x733 & ~x734 & ~x739 & ~x741 & ~x742 & ~x749 & ~x751 & ~x752 & ~x753 & ~x756 & ~x761 & ~x763 & ~x770 & ~x772 & ~x773 & ~x774 & ~x777 & ~x779 & ~x781 & ~x782 & ~x783;
assign c5128 =  x187 &  x188 &  x210 &  x212 & ~x13 & ~x18 & ~x20 & ~x32 & ~x54 & ~x59 & ~x63 & ~x65 & ~x66 & ~x68 & ~x74 & ~x81 & ~x84 & ~x87 & ~x90 & ~x99 & ~x100 & ~x101 & ~x108 & ~x109 & ~x115 & ~x136 & ~x143 & ~x144 & ~x147 & ~x148 & ~x196 & ~x226 & ~x228 & ~x248 & ~x271 & ~x272 & ~x286 & ~x287 & ~x300 & ~x303 & ~x306 & ~x309 & ~x331 & ~x332 & ~x336 & ~x337 & ~x360 & ~x365 & ~x366 & ~x387 & ~x392 & ~x393 & ~x394 & ~x416 & ~x422 & ~x443 & ~x448 & ~x449 & ~x476 & ~x477 & ~x499 & ~x501 & ~x556 & ~x557 & ~x584 & ~x588 & ~x615 & ~x619 & ~x620 & ~x643 & ~x672 & ~x673 & ~x674 & ~x676 & ~x683 & ~x691 & ~x692 & ~x694 & ~x697 & ~x699 & ~x703 & ~x720 & ~x726 & ~x744 & ~x750 & ~x751 & ~x753 & ~x756 & ~x769 & ~x774 & ~x777;
assign c5130 =  x699;
assign c5132 =  x9;
assign c5134 = ~x2 & ~x3 & ~x13 & ~x39 & ~x40 & ~x44 & ~x69 & ~x71 & ~x90 & ~x97 & ~x110 & ~x123 & ~x124 & ~x125 & ~x138 & ~x139 & ~x146 & ~x150 & ~x151 & ~x174 & ~x179 & ~x201 & ~x205 & ~x207 & ~x223 & ~x252 & ~x261 & ~x262 & ~x284 & ~x288 & ~x311 & ~x337 & ~x356 & ~x364 & ~x441 & ~x445 & ~x457 & ~x487 & ~x488 & ~x497 & ~x502 & ~x530 & ~x552 & ~x562 & ~x579 & ~x590 & ~x592 & ~x605 & ~x613 & ~x614 & ~x621 & ~x634 & ~x637 & ~x647 & ~x660 & ~x662 & ~x686 & ~x706 & ~x707 & ~x708 & ~x711 & ~x715 & ~x717 & ~x724 & ~x734 & ~x736 & ~x739 & ~x740 & ~x742 & ~x743 & ~x744 & ~x764;
assign c5136 = ~x1 & ~x6 & ~x8 & ~x9 & ~x10 & ~x12 & ~x15 & ~x18 & ~x19 & ~x24 & ~x25 & ~x27 & ~x32 & ~x35 & ~x36 & ~x38 & ~x46 & ~x48 & ~x49 & ~x50 & ~x51 & ~x52 & ~x54 & ~x56 & ~x58 & ~x60 & ~x64 & ~x65 & ~x66 & ~x68 & ~x70 & ~x71 & ~x73 & ~x80 & ~x87 & ~x88 & ~x92 & ~x95 & ~x102 & ~x109 & ~x112 & ~x116 & ~x118 & ~x133 & ~x134 & ~x137 & ~x140 & ~x142 & ~x145 & ~x166 & ~x172 & ~x193 & ~x195 & ~x196 & ~x221 & ~x223 & ~x225 & ~x249 & ~x255 & ~x265 & ~x270 & ~x273 & ~x275 & ~x279 & ~x294 & ~x295 & ~x297 & ~x298 & ~x299 & ~x300 & ~x304 & ~x305 & ~x308 & ~x311 & ~x328 & ~x329 & ~x331 & ~x336 & ~x337 & ~x339 & ~x358 & ~x363 & ~x365 & ~x366 & ~x367 & ~x389 & ~x390 & ~x392 & ~x394 & ~x396 & ~x416 & ~x418 & ~x422 & ~x446 & ~x448 & ~x450 & ~x451 & ~x452 & ~x476 & ~x477 & ~x478 & ~x479 & ~x489 & ~x501 & ~x504 & ~x506 & ~x516 & ~x517 & ~x519 & ~x520 & ~x533 & ~x535 & ~x547 & ~x559 & ~x560 & ~x562 & ~x587 & ~x588 & ~x590 & ~x592 & ~x593 & ~x594 & ~x613 & ~x614 & ~x616 & ~x618 & ~x621 & ~x643 & ~x672 & ~x675 & ~x676 & ~x678 & ~x695 & ~x696 & ~x697 & ~x699 & ~x710 & ~x722 & ~x723 & ~x724 & ~x725 & ~x726 & ~x728 & ~x732 & ~x733 & ~x734 & ~x735 & ~x736 & ~x737 & ~x740 & ~x741 & ~x747 & ~x750 & ~x753 & ~x756 & ~x757 & ~x759 & ~x763 & ~x767 & ~x768 & ~x769 & ~x770 & ~x773 & ~x774 & ~x775 & ~x778 & ~x782 & ~x783;
assign c5138 =  x210 &  x211 & ~x5 & ~x7 & ~x18 & ~x20 & ~x21 & ~x25 & ~x28 & ~x32 & ~x33 & ~x35 & ~x37 & ~x45 & ~x46 & ~x56 & ~x64 & ~x65 & ~x72 & ~x77 & ~x83 & ~x85 & ~x87 & ~x102 & ~x108 & ~x124 & ~x129 & ~x135 & ~x144 & ~x146 & ~x147 & ~x164 & ~x165 & ~x167 & ~x169 & ~x170 & ~x175 & ~x198 & ~x199 & ~x224 & ~x227 & ~x230 & ~x252 & ~x274 & ~x284 & ~x285 & ~x296 & ~x309 & ~x326 & ~x327 & ~x328 & ~x331 & ~x334 & ~x337 & ~x356 & ~x361 & ~x364 & ~x367 & ~x368 & ~x385 & ~x388 & ~x390 & ~x391 & ~x442 & ~x445 & ~x448 & ~x452 & ~x477 & ~x482 & ~x502 & ~x503 & ~x504 & ~x509 & ~x517 & ~x528 & ~x532 & ~x561 & ~x588 & ~x591 & ~x611 & ~x613 & ~x615 & ~x620 & ~x642 & ~x671 & ~x675 & ~x676 & ~x702 & ~x724 & ~x727 & ~x735 & ~x736 & ~x738 & ~x744 & ~x751 & ~x762 & ~x763 & ~x769 & ~x772 & ~x773 & ~x774 & ~x780 & ~x781;
assign c5140 =  x164;
assign c5142 =  x204 &  x314 &  x346 &  x371 & ~x302;
assign c5144 =  x264 &  x292 & ~x2 & ~x4 & ~x11 & ~x15 & ~x18 & ~x29 & ~x36 & ~x38 & ~x42 & ~x45 & ~x47 & ~x51 & ~x59 & ~x61 & ~x65 & ~x70 & ~x75 & ~x80 & ~x83 & ~x91 & ~x95 & ~x98 & ~x103 & ~x106 & ~x117 & ~x118 & ~x119 & ~x122 & ~x125 & ~x139 & ~x165 & ~x166 & ~x168 & ~x174 & ~x196 & ~x202 & ~x204 & ~x255 & ~x259 & ~x283 & ~x285 & ~x286 & ~x307 & ~x310 & ~x311 & ~x336 & ~x340 & ~x364 & ~x367 & ~x387 & ~x396 & ~x397 & ~x398 & ~x413 & ~x422 & ~x441 & ~x444 & ~x445 & ~x448 & ~x475 & ~x476 & ~x481 & ~x515 & ~x531 & ~x542 & ~x554 & ~x555 & ~x556 & ~x581 & ~x588 & ~x590 & ~x608 & ~x611 & ~x612 & ~x617 & ~x619 & ~x637 & ~x640 & ~x641 & ~x643 & ~x645 & ~x646 & ~x648 & ~x665 & ~x666 & ~x667 & ~x675 & ~x678 & ~x689 & ~x690 & ~x692 & ~x695 & ~x700 & ~x701 & ~x702 & ~x703 & ~x708 & ~x709 & ~x716 & ~x717 & ~x719 & ~x724 & ~x725 & ~x738 & ~x740 & ~x742 & ~x743 & ~x745 & ~x746 & ~x752 & ~x753 & ~x757 & ~x759 & ~x764 & ~x766 & ~x767 & ~x770 & ~x783;
assign c5146 =  x270 &  x273 &  x374 & ~x159 & ~x257 & ~x385 & ~x387 & ~x453;
assign c5148 = ~x128 & ~x161 & ~x183 & ~x184 & ~x313 & ~x342 & ~x408 & ~x409 & ~x439 & ~x440 & ~x467 & ~x496 & ~x576 & ~x591 & ~x610 & ~x641 & ~x725 & ~x727 & ~x736;
assign c5150 =  x88;
assign c5152 =  x189 & ~x0 & ~x2 & ~x5 & ~x8 & ~x10 & ~x22 & ~x23 & ~x30 & ~x34 & ~x37 & ~x47 & ~x52 & ~x55 & ~x59 & ~x70 & ~x72 & ~x75 & ~x76 & ~x77 & ~x78 & ~x82 & ~x85 & ~x87 & ~x88 & ~x90 & ~x95 & ~x97 & ~x99 & ~x107 & ~x108 & ~x109 & ~x111 & ~x120 & ~x121 & ~x139 & ~x143 & ~x145 & ~x149 & ~x167 & ~x168 & ~x169 & ~x173 & ~x174 & ~x175 & ~x194 & ~x197 & ~x199 & ~x227 & ~x249 & ~x250 & ~x251 & ~x252 & ~x253 & ~x254 & ~x255 & ~x256 & ~x257 & ~x279 & ~x282 & ~x284 & ~x298 & ~x300 & ~x304 & ~x308 & ~x312 & ~x328 & ~x330 & ~x332 & ~x333 & ~x334 & ~x335 & ~x340 & ~x362 & ~x366 & ~x367 & ~x386 & ~x387 & ~x388 & ~x392 & ~x394 & ~x414 & ~x416 & ~x417 & ~x418 & ~x419 & ~x420 & ~x423 & ~x443 & ~x444 & ~x450 & ~x472 & ~x475 & ~x502 & ~x527 & ~x528 & ~x531 & ~x533 & ~x557 & ~x564 & ~x583 & ~x585 & ~x591 & ~x608 & ~x611 & ~x613 & ~x618 & ~x619 & ~x642 & ~x643 & ~x666 & ~x667 & ~x670 & ~x673 & ~x676 & ~x693 & ~x695 & ~x697 & ~x699 & ~x700 & ~x703 & ~x705 & ~x716 & ~x719 & ~x722 & ~x724 & ~x725 & ~x730 & ~x734 & ~x738 & ~x741 & ~x744 & ~x746 & ~x747 & ~x748 & ~x753 & ~x756 & ~x757 & ~x758 & ~x764 & ~x766 & ~x767 & ~x771 & ~x774 & ~x775 & ~x776 & ~x780 & ~x781;
assign c5154 = ~x1 & ~x5 & ~x9 & ~x21 & ~x26 & ~x30 & ~x33 & ~x35 & ~x37 & ~x42 & ~x46 & ~x47 & ~x49 & ~x52 & ~x53 & ~x59 & ~x65 & ~x76 & ~x79 & ~x82 & ~x84 & ~x85 & ~x90 & ~x91 & ~x93 & ~x96 & ~x98 & ~x99 & ~x101 & ~x103 & ~x104 & ~x105 & ~x110 & ~x118 & ~x121 & ~x124 & ~x138 & ~x140 & ~x143 & ~x144 & ~x147 & ~x166 & ~x195 & ~x198 & ~x200 & ~x229 & ~x252 & ~x283 & ~x308 & ~x311 & ~x312 & ~x322 & ~x323 & ~x334 & ~x338 & ~x353 & ~x357 & ~x366 & ~x368 & ~x383 & ~x384 & ~x387 & ~x393 & ~x394 & ~x397 & ~x415 & ~x423 & ~x424 & ~x441 & ~x443 & ~x454 & ~x471 & ~x498 & ~x499 & ~x504 & ~x527 & ~x534 & ~x543 & ~x560 & ~x561 & ~x564 & ~x570 & ~x597 & ~x614 & ~x617 & ~x642 & ~x645 & ~x648 & ~x649 & ~x668 & ~x671 & ~x677 & ~x695 & ~x702 & ~x703 & ~x725 & ~x735 & ~x736 & ~x737 & ~x738 & ~x739 & ~x745 & ~x752 & ~x754 & ~x759 & ~x760 & ~x761 & ~x769 & ~x770 & ~x771 & ~x779 & ~x782;
assign c5156 =  x289 &  x317 &  x345 &  x346 & ~x7 & ~x8 & ~x14 & ~x15 & ~x24 & ~x27 & ~x37 & ~x38 & ~x43 & ~x44 & ~x47 & ~x48 & ~x49 & ~x52 & ~x61 & ~x62 & ~x70 & ~x73 & ~x74 & ~x77 & ~x78 & ~x86 & ~x91 & ~x93 & ~x96 & ~x101 & ~x121 & ~x123 & ~x134 & ~x135 & ~x142 & ~x146 & ~x165 & ~x166 & ~x170 & ~x172 & ~x281 & ~x284 & ~x330 & ~x333 & ~x336 & ~x338 & ~x361 & ~x389 & ~x391 & ~x394 & ~x419 & ~x422 & ~x447 & ~x450 & ~x451 & ~x472 & ~x478 & ~x483 & ~x510 & ~x512 & ~x514 & ~x515 & ~x545 & ~x559 & ~x562 & ~x574 & ~x587 & ~x612 & ~x640 & ~x669 & ~x675 & ~x701 & ~x705 & ~x708 & ~x719 & ~x724 & ~x725 & ~x729 & ~x745 & ~x751 & ~x753 & ~x756 & ~x758 & ~x761 & ~x768 & ~x771 & ~x772 & ~x775 & ~x782;
assign c5158 =  x724;
assign c5160 =  x47;
assign c5162 =  x234 &  x262 &  x290 &  x632 & ~x3 & ~x4 & ~x5 & ~x26 & ~x32 & ~x37 & ~x39 & ~x40 & ~x41 & ~x47 & ~x48 & ~x51 & ~x53 & ~x54 & ~x58 & ~x60 & ~x62 & ~x67 & ~x72 & ~x75 & ~x78 & ~x81 & ~x83 & ~x88 & ~x89 & ~x100 & ~x102 & ~x103 & ~x104 & ~x109 & ~x112 & ~x115 & ~x117 & ~x140 & ~x145 & ~x146 & ~x164 & ~x194 & ~x221 & ~x225 & ~x245 & ~x247 & ~x249 & ~x255 & ~x269 & ~x272 & ~x274 & ~x277 & ~x279 & ~x283 & ~x300 & ~x302 & ~x303 & ~x304 & ~x305 & ~x308 & ~x309 & ~x311 & ~x330 & ~x332 & ~x334 & ~x337 & ~x340 & ~x363 & ~x365 & ~x389 & ~x391 & ~x392 & ~x418 & ~x445 & ~x448 & ~x449 & ~x450 & ~x455 & ~x464 & ~x473 & ~x474 & ~x475 & ~x476 & ~x500 & ~x501 & ~x504 & ~x507 & ~x518 & ~x520 & ~x528 & ~x529 & ~x533 & ~x534 & ~x556 & ~x562 & ~x583 & ~x588 & ~x611 & ~x612 & ~x614 & ~x615 & ~x641 & ~x642 & ~x648 & ~x666 & ~x667 & ~x668 & ~x671 & ~x691 & ~x705 & ~x706 & ~x717 & ~x725 & ~x726 & ~x728 & ~x731 & ~x736 & ~x741 & ~x742 & ~x744 & ~x747 & ~x748 & ~x750 & ~x751 & ~x760 & ~x763 & ~x768 & ~x769 & ~x774 & ~x775 & ~x780;
assign c5164 =  x196;
assign c5166 =  x185 & ~x2 & ~x3 & ~x4 & ~x8 & ~x9 & ~x11 & ~x12 & ~x13 & ~x18 & ~x19 & ~x20 & ~x21 & ~x23 & ~x24 & ~x25 & ~x26 & ~x27 & ~x28 & ~x30 & ~x31 & ~x35 & ~x36 & ~x37 & ~x38 & ~x41 & ~x42 & ~x43 & ~x46 & ~x48 & ~x49 & ~x50 & ~x51 & ~x53 & ~x54 & ~x55 & ~x57 & ~x58 & ~x59 & ~x60 & ~x62 & ~x63 & ~x64 & ~x65 & ~x66 & ~x67 & ~x70 & ~x72 & ~x73 & ~x74 & ~x75 & ~x76 & ~x77 & ~x78 & ~x79 & ~x80 & ~x81 & ~x83 & ~x85 & ~x86 & ~x88 & ~x90 & ~x92 & ~x94 & ~x95 & ~x105 & ~x106 & ~x108 & ~x109 & ~x110 & ~x112 & ~x115 & ~x118 & ~x121 & ~x122 & ~x135 & ~x137 & ~x139 & ~x140 & ~x141 & ~x142 & ~x145 & ~x147 & ~x148 & ~x149 & ~x164 & ~x165 & ~x166 & ~x167 & ~x170 & ~x175 & ~x176 & ~x192 & ~x197 & ~x199 & ~x200 & ~x201 & ~x202 & ~x203 & ~x220 & ~x221 & ~x222 & ~x223 & ~x225 & ~x226 & ~x229 & ~x231 & ~x244 & ~x248 & ~x253 & ~x255 & ~x258 & ~x270 & ~x271 & ~x272 & ~x274 & ~x275 & ~x276 & ~x277 & ~x281 & ~x284 & ~x285 & ~x298 & ~x299 & ~x300 & ~x301 & ~x302 & ~x305 & ~x306 & ~x307 & ~x308 & ~x310 & ~x311 & ~x312 & ~x313 & ~x328 & ~x330 & ~x331 & ~x332 & ~x334 & ~x336 & ~x337 & ~x339 & ~x342 & ~x358 & ~x359 & ~x360 & ~x363 & ~x365 & ~x366 & ~x367 & ~x368 & ~x370 & ~x385 & ~x386 & ~x387 & ~x388 & ~x389 & ~x390 & ~x391 & ~x392 & ~x393 & ~x394 & ~x398 & ~x414 & ~x417 & ~x419 & ~x420 & ~x421 & ~x422 & ~x423 & ~x424 & ~x425 & ~x442 & ~x444 & ~x445 & ~x447 & ~x449 & ~x450 & ~x453 & ~x455 & ~x470 & ~x471 & ~x472 & ~x474 & ~x475 & ~x476 & ~x477 & ~x478 & ~x479 & ~x481 & ~x483 & ~x499 & ~x500 & ~x502 & ~x503 & ~x505 & ~x510 & ~x512 & ~x526 & ~x530 & ~x532 & ~x533 & ~x536 & ~x538 & ~x539 & ~x541 & ~x554 & ~x556 & ~x557 & ~x558 & ~x559 & ~x560 & ~x562 & ~x582 & ~x583 & ~x584 & ~x585 & ~x586 & ~x587 & ~x588 & ~x589 & ~x590 & ~x609 & ~x610 & ~x611 & ~x613 & ~x616 & ~x617 & ~x619 & ~x639 & ~x641 & ~x643 & ~x644 & ~x646 & ~x647 & ~x648 & ~x662 & ~x664 & ~x666 & ~x667 & ~x671 & ~x672 & ~x674 & ~x675 & ~x677 & ~x692 & ~x693 & ~x694 & ~x695 & ~x698 & ~x699 & ~x700 & ~x704 & ~x705 & ~x706 & ~x708 & ~x711 & ~x712 & ~x713 & ~x714 & ~x715 & ~x717 & ~x720 & ~x721 & ~x723 & ~x725 & ~x726 & ~x730 & ~x732 & ~x736 & ~x738 & ~x742 & ~x746 & ~x747 & ~x750 & ~x753 & ~x754 & ~x755 & ~x756 & ~x758 & ~x759 & ~x763 & ~x764 & ~x765 & ~x766 & ~x767 & ~x768 & ~x770 & ~x771 & ~x774 & ~x777 & ~x778 & ~x779 & ~x782 & ~x783;
assign c5168 =  x276;
assign c5172 =  x155 & ~x7 & ~x25 & ~x112 & ~x245 & ~x267 & ~x268 & ~x269 & ~x271 & ~x328 & ~x335 & ~x360 & ~x424 & ~x452 & ~x484 & ~x486 & ~x487 & ~x669 & ~x676 & ~x739 & ~x767;
assign c5174 =  x324 & ~x3 & ~x15 & ~x18 & ~x77 & ~x96 & ~x97 & ~x111 & ~x119 & ~x161 & ~x198 & ~x202 & ~x214 & ~x222 & ~x240 & ~x260 & ~x362 & ~x386 & ~x399 & ~x445 & ~x504 & ~x556 & ~x651 & ~x668 & ~x701 & ~x706 & ~x707 & ~x709 & ~x715 & ~x739 & ~x759 & ~x763;
assign c5176 = ~x6 & ~x10 & ~x12 & ~x25 & ~x26 & ~x33 & ~x34 & ~x36 & ~x44 & ~x46 & ~x48 & ~x53 & ~x56 & ~x59 & ~x60 & ~x62 & ~x63 & ~x65 & ~x67 & ~x69 & ~x75 & ~x77 & ~x83 & ~x85 & ~x86 & ~x88 & ~x93 & ~x98 & ~x100 & ~x101 & ~x103 & ~x110 & ~x119 & ~x120 & ~x123 & ~x131 & ~x139 & ~x140 & ~x144 & ~x145 & ~x146 & ~x148 & ~x166 & ~x168 & ~x170 & ~x172 & ~x174 & ~x176 & ~x202 & ~x229 & ~x231 & ~x253 & ~x256 & ~x280 & ~x283 & ~x287 & ~x307 & ~x308 & ~x310 & ~x313 & ~x350 & ~x352 & ~x381 & ~x382 & ~x384 & ~x385 & ~x386 & ~x389 & ~x390 & ~x391 & ~x395 & ~x414 & ~x415 & ~x422 & ~x425 & ~x426 & ~x442 & ~x445 & ~x447 & ~x448 & ~x452 & ~x453 & ~x472 & ~x473 & ~x481 & ~x503 & ~x504 & ~x509 & ~x525 & ~x528 & ~x535 & ~x536 & ~x554 & ~x557 & ~x558 & ~x584 & ~x585 & ~x666 & ~x669 & ~x672 & ~x694 & ~x696 & ~x697 & ~x698 & ~x706 & ~x723 & ~x724 & ~x728 & ~x734 & ~x745 & ~x746 & ~x748 & ~x756 & ~x774 & ~x775 & ~x779 & ~x782;
assign c5178 =  x347 &  x372 & ~x18 & ~x62 & ~x63 & ~x69 & ~x114 & ~x117 & ~x281 & ~x283 & ~x408 & ~x409 & ~x437 & ~x450 & ~x482 & ~x483 & ~x484 & ~x534 & ~x535 & ~x560 & ~x563 & ~x618 & ~x758 & ~x770;
assign c5180 =  x238 &  x241 & ~x1 & ~x13 & ~x25 & ~x45 & ~x52 & ~x68 & ~x75 & ~x85 & ~x86 & ~x94 & ~x97 & ~x101 & ~x102 & ~x104 & ~x110 & ~x111 & ~x115 & ~x125 & ~x128 & ~x132 & ~x149 & ~x228 & ~x279 & ~x281 & ~x285 & ~x311 & ~x325 & ~x326 & ~x336 & ~x339 & ~x355 & ~x359 & ~x383 & ~x384 & ~x445 & ~x448 & ~x450 & ~x470 & ~x471 & ~x475 & ~x500 & ~x532 & ~x554 & ~x584 & ~x609 & ~x611 & ~x613 & ~x616 & ~x636 & ~x637 & ~x676 & ~x692 & ~x695 & ~x697 & ~x698 & ~x702 & ~x715 & ~x716 & ~x718 & ~x728 & ~x740 & ~x743 & ~x744 & ~x748 & ~x759 & ~x771 & ~x777 & ~x781 & ~x783;
assign c5182 =  x600 & ~x20 & ~x25 & ~x37 & ~x44 & ~x46 & ~x51 & ~x56 & ~x61 & ~x72 & ~x82 & ~x86 & ~x87 & ~x96 & ~x103 & ~x108 & ~x111 & ~x138 & ~x146 & ~x196 & ~x199 & ~x253 & ~x296 & ~x327 & ~x364 & ~x385 & ~x387 & ~x389 & ~x397 & ~x398 & ~x413 & ~x421 & ~x428 & ~x442 & ~x445 & ~x450 & ~x470 & ~x473 & ~x474 & ~x486 & ~x508 & ~x529 & ~x589 & ~x620 & ~x645 & ~x669 & ~x677 & ~x720 & ~x723 & ~x732 & ~x769;
assign c5184 = ~x4 & ~x7 & ~x8 & ~x18 & ~x27 & ~x32 & ~x33 & ~x35 & ~x36 & ~x40 & ~x45 & ~x54 & ~x55 & ~x68 & ~x76 & ~x88 & ~x89 & ~x91 & ~x98 & ~x103 & ~x117 & ~x122 & ~x128 & ~x138 & ~x141 & ~x155 & ~x157 & ~x167 & ~x173 & ~x175 & ~x185 & ~x187 & ~x197 & ~x201 & ~x203 & ~x230 & ~x250 & ~x252 & ~x257 & ~x258 & ~x280 & ~x284 & ~x309 & ~x313 & ~x337 & ~x340 & ~x354 & ~x357 & ~x359 & ~x362 & ~x385 & ~x386 & ~x416 & ~x418 & ~x424 & ~x446 & ~x448 & ~x449 & ~x471 & ~x475 & ~x501 & ~x503 & ~x527 & ~x529 & ~x531 & ~x532 & ~x562 & ~x584 & ~x586 & ~x611 & ~x613 & ~x616 & ~x617 & ~x644 & ~x669 & ~x697 & ~x698 & ~x703 & ~x704 & ~x707 & ~x708 & ~x710 & ~x719 & ~x730 & ~x738 & ~x740 & ~x748 & ~x753 & ~x754 & ~x760 & ~x769 & ~x770;
assign c5186 =  x155 & ~x1 & ~x2 & ~x12 & ~x14 & ~x15 & ~x18 & ~x20 & ~x24 & ~x25 & ~x26 & ~x28 & ~x33 & ~x34 & ~x36 & ~x37 & ~x42 & ~x43 & ~x51 & ~x56 & ~x62 & ~x72 & ~x73 & ~x77 & ~x85 & ~x88 & ~x89 & ~x91 & ~x92 & ~x94 & ~x95 & ~x110 & ~x114 & ~x139 & ~x140 & ~x142 & ~x144 & ~x162 & ~x166 & ~x169 & ~x173 & ~x190 & ~x191 & ~x200 & ~x223 & ~x224 & ~x225 & ~x240 & ~x243 & ~x244 & ~x251 & ~x252 & ~x269 & ~x270 & ~x272 & ~x273 & ~x274 & ~x276 & ~x277 & ~x285 & ~x302 & ~x303 & ~x304 & ~x309 & ~x327 & ~x329 & ~x334 & ~x336 & ~x339 & ~x340 & ~x341 & ~x358 & ~x359 & ~x362 & ~x363 & ~x366 & ~x387 & ~x388 & ~x389 & ~x393 & ~x394 & ~x396 & ~x415 & ~x418 & ~x419 & ~x420 & ~x422 & ~x423 & ~x444 & ~x445 & ~x448 & ~x473 & ~x474 & ~x475 & ~x478 & ~x485 & ~x500 & ~x501 & ~x504 & ~x506 & ~x515 & ~x516 & ~x517 & ~x529 & ~x556 & ~x559 & ~x563 & ~x592 & ~x593 & ~x613 & ~x614 & ~x643 & ~x644 & ~x669 & ~x670 & ~x671 & ~x676 & ~x679 & ~x691 & ~x692 & ~x697 & ~x703 & ~x704 & ~x706 & ~x708 & ~x713 & ~x719 & ~x721 & ~x724 & ~x729 & ~x732 & ~x733 & ~x737 & ~x744 & ~x746 & ~x749 & ~x750 & ~x752 & ~x761 & ~x762 & ~x763 & ~x766 & ~x767 & ~x768 & ~x769 & ~x772 & ~x773 & ~x774 & ~x778 & ~x780 & ~x782;
assign c5188 =  x141;
assign c5190 =  x192;
assign c5192 =  x24;
assign c5194 =  x260 &  x288 & ~x0 & ~x2 & ~x4 & ~x5 & ~x7 & ~x8 & ~x10 & ~x11 & ~x13 & ~x18 & ~x20 & ~x25 & ~x27 & ~x28 & ~x32 & ~x34 & ~x40 & ~x42 & ~x46 & ~x49 & ~x50 & ~x52 & ~x60 & ~x63 & ~x65 & ~x66 & ~x75 & ~x77 & ~x80 & ~x82 & ~x84 & ~x88 & ~x100 & ~x101 & ~x110 & ~x115 & ~x116 & ~x117 & ~x135 & ~x136 & ~x137 & ~x141 & ~x142 & ~x144 & ~x164 & ~x166 & ~x171 & ~x197 & ~x221 & ~x224 & ~x225 & ~x226 & ~x227 & ~x253 & ~x254 & ~x256 & ~x267 & ~x268 & ~x269 & ~x270 & ~x271 & ~x272 & ~x274 & ~x275 & ~x300 & ~x301 & ~x303 & ~x304 & ~x306 & ~x309 & ~x311 & ~x329 & ~x330 & ~x332 & ~x338 & ~x340 & ~x388 & ~x392 & ~x418 & ~x421 & ~x446 & ~x450 & ~x453 & ~x475 & ~x476 & ~x479 & ~x489 & ~x490 & ~x503 & ~x507 & ~x517 & ~x518 & ~x519 & ~x530 & ~x534 & ~x559 & ~x562 & ~x587 & ~x591 & ~x613 & ~x640 & ~x643 & ~x645 & ~x646 & ~x647 & ~x667 & ~x670 & ~x674 & ~x676 & ~x677 & ~x680 & ~x695 & ~x700 & ~x701 & ~x705 & ~x707 & ~x721 & ~x724 & ~x725 & ~x727 & ~x728 & ~x732 & ~x736 & ~x737 & ~x739 & ~x745 & ~x747 & ~x748 & ~x750 & ~x758 & ~x762 & ~x767 & ~x770 & ~x771 & ~x778 & ~x781;
assign c5196 =  x263 &  x290 &  x318 &  x347 & ~x0 & ~x3 & ~x5 & ~x6 & ~x8 & ~x10 & ~x15 & ~x20 & ~x21 & ~x23 & ~x24 & ~x32 & ~x33 & ~x40 & ~x41 & ~x49 & ~x54 & ~x56 & ~x57 & ~x59 & ~x63 & ~x69 & ~x72 & ~x73 & ~x74 & ~x80 & ~x82 & ~x88 & ~x92 & ~x100 & ~x101 & ~x102 & ~x103 & ~x105 & ~x107 & ~x108 & ~x109 & ~x116 & ~x119 & ~x120 & ~x121 & ~x135 & ~x138 & ~x140 & ~x145 & ~x164 & ~x165 & ~x168 & ~x173 & ~x174 & ~x176 & ~x194 & ~x201 & ~x203 & ~x230 & ~x251 & ~x252 & ~x254 & ~x256 & ~x258 & ~x281 & ~x283 & ~x286 & ~x305 & ~x306 & ~x309 & ~x313 & ~x330 & ~x358 & ~x359 & ~x361 & ~x365 & ~x367 & ~x369 & ~x390 & ~x391 & ~x395 & ~x423 & ~x424 & ~x427 & ~x448 & ~x455 & ~x472 & ~x473 & ~x488 & ~x499 & ~x500 & ~x501 & ~x506 & ~x514 & ~x517 & ~x518 & ~x528 & ~x532 & ~x535 & ~x563 & ~x582 & ~x588 & ~x590 & ~x591 & ~x610 & ~x617 & ~x640 & ~x643 & ~x644 & ~x647 & ~x664 & ~x666 & ~x669 & ~x676 & ~x700 & ~x702 & ~x709 & ~x717 & ~x719 & ~x720 & ~x726 & ~x732 & ~x733 & ~x740 & ~x742 & ~x762 & ~x764 & ~x765 & ~x769 & ~x773 & ~x774 & ~x777 & ~x780 & ~x781 & ~x783;
assign c5198 =  x626 & ~x0 & ~x11 & ~x30 & ~x50 & ~x75 & ~x117 & ~x143 & ~x164 & ~x190 & ~x195 & ~x215 & ~x217 & ~x224 & ~x241 & ~x244 & ~x266 & ~x272 & ~x427 & ~x449 & ~x478 & ~x529 & ~x611 & ~x644 & ~x674 & ~x688 & ~x714 & ~x718 & ~x719 & ~x735 & ~x737 & ~x783;
assign c5200 =  x599 &  x600 &  x601 & ~x2 & ~x5 & ~x12 & ~x15 & ~x21 & ~x23 & ~x25 & ~x30 & ~x31 & ~x32 & ~x34 & ~x35 & ~x36 & ~x38 & ~x44 & ~x48 & ~x56 & ~x58 & ~x62 & ~x65 & ~x66 & ~x67 & ~x68 & ~x70 & ~x81 & ~x85 & ~x93 & ~x110 & ~x114 & ~x140 & ~x143 & ~x168 & ~x170 & ~x174 & ~x198 & ~x222 & ~x224 & ~x228 & ~x247 & ~x248 & ~x254 & ~x267 & ~x268 & ~x269 & ~x270 & ~x273 & ~x274 & ~x275 & ~x282 & ~x284 & ~x300 & ~x304 & ~x312 & ~x329 & ~x330 & ~x339 & ~x357 & ~x358 & ~x362 & ~x363 & ~x365 & ~x369 & ~x387 & ~x390 & ~x392 & ~x394 & ~x396 & ~x398 & ~x400 & ~x416 & ~x417 & ~x421 & ~x427 & ~x428 & ~x429 & ~x443 & ~x445 & ~x447 & ~x448 & ~x450 & ~x457 & ~x458 & ~x459 & ~x472 & ~x476 & ~x478 & ~x502 & ~x504 & ~x533 & ~x558 & ~x560 & ~x562 & ~x591 & ~x613 & ~x617 & ~x619 & ~x642 & ~x643 & ~x665 & ~x668 & ~x674 & ~x675 & ~x682 & ~x683 & ~x685 & ~x691 & ~x694 & ~x695 & ~x696 & ~x708 & ~x711 & ~x713 & ~x715 & ~x721 & ~x724 & ~x726 & ~x729 & ~x737 & ~x746 & ~x750 & ~x753 & ~x756 & ~x758 & ~x763 & ~x767 & ~x775 & ~x776 & ~x777 & ~x781;
assign c5202 =  x242 & ~x3 & ~x8 & ~x10 & ~x20 & ~x25 & ~x31 & ~x35 & ~x41 & ~x47 & ~x54 & ~x64 & ~x70 & ~x71 & ~x75 & ~x84 & ~x85 & ~x89 & ~x90 & ~x100 & ~x107 & ~x114 & ~x119 & ~x127 & ~x129 & ~x143 & ~x146 & ~x148 & ~x150 & ~x157 & ~x174 & ~x201 & ~x259 & ~x312 & ~x325 & ~x326 & ~x328 & ~x329 & ~x330 & ~x332 & ~x336 & ~x355 & ~x360 & ~x361 & ~x384 & ~x390 & ~x391 & ~x395 & ~x396 & ~x414 & ~x416 & ~x417 & ~x441 & ~x444 & ~x445 & ~x450 & ~x451 & ~x475 & ~x499 & ~x500 & ~x501 & ~x502 & ~x503 & ~x526 & ~x528 & ~x529 & ~x534 & ~x562 & ~x584 & ~x590 & ~x612 & ~x647 & ~x670 & ~x672 & ~x673 & ~x677 & ~x694 & ~x696 & ~x719 & ~x722 & ~x723 & ~x728 & ~x737 & ~x740 & ~x746 & ~x755 & ~x764 & ~x765 & ~x771 & ~x774 & ~x775 & ~x776 & ~x778 & ~x779 & ~x781 & ~x783;
assign c5204 =  x46;
assign c5206 =  x179 & ~x0 & ~x2 & ~x5 & ~x11 & ~x13 & ~x19 & ~x22 & ~x26 & ~x27 & ~x28 & ~x32 & ~x33 & ~x36 & ~x37 & ~x44 & ~x45 & ~x50 & ~x51 & ~x52 & ~x53 & ~x55 & ~x56 & ~x57 & ~x58 & ~x63 & ~x64 & ~x65 & ~x67 & ~x68 & ~x69 & ~x81 & ~x83 & ~x84 & ~x86 & ~x89 & ~x90 & ~x91 & ~x93 & ~x94 & ~x104 & ~x105 & ~x107 & ~x109 & ~x111 & ~x112 & ~x113 & ~x114 & ~x116 & ~x134 & ~x137 & ~x139 & ~x140 & ~x142 & ~x144 & ~x164 & ~x166 & ~x167 & ~x168 & ~x171 & ~x192 & ~x195 & ~x196 & ~x198 & ~x200 & ~x218 & ~x221 & ~x222 & ~x225 & ~x226 & ~x227 & ~x244 & ~x245 & ~x249 & ~x250 & ~x251 & ~x252 & ~x254 & ~x265 & ~x266 & ~x267 & ~x268 & ~x269 & ~x270 & ~x272 & ~x273 & ~x277 & ~x278 & ~x280 & ~x282 & ~x298 & ~x299 & ~x300 & ~x301 & ~x302 & ~x303 & ~x311 & ~x329 & ~x330 & ~x332 & ~x334 & ~x335 & ~x338 & ~x339 & ~x360 & ~x361 & ~x364 & ~x367 & ~x388 & ~x389 & ~x392 & ~x394 & ~x395 & ~x418 & ~x420 & ~x425 & ~x446 & ~x447 & ~x449 & ~x450 & ~x474 & ~x475 & ~x477 & ~x502 & ~x503 & ~x506 & ~x507 & ~x508 & ~x518 & ~x532 & ~x535 & ~x536 & ~x537 & ~x545 & ~x546 & ~x547 & ~x557 & ~x559 & ~x560 & ~x584 & ~x589 & ~x590 & ~x592 & ~x593 & ~x615 & ~x616 & ~x617 & ~x618 & ~x619 & ~x621 & ~x639 & ~x640 & ~x641 & ~x642 & ~x643 & ~x645 & ~x649 & ~x651 & ~x665 & ~x666 & ~x669 & ~x670 & ~x674 & ~x676 & ~x679 & ~x680 & ~x681 & ~x692 & ~x695 & ~x697 & ~x698 & ~x699 & ~x701 & ~x702 & ~x703 & ~x705 & ~x708 & ~x710 & ~x711 & ~x723 & ~x725 & ~x727 & ~x728 & ~x729 & ~x730 & ~x733 & ~x734 & ~x736 & ~x737 & ~x738 & ~x739 & ~x740 & ~x741 & ~x746 & ~x747 & ~x749 & ~x752 & ~x753 & ~x754 & ~x755 & ~x758 & ~x759 & ~x760 & ~x764 & ~x765 & ~x768 & ~x771 & ~x772 & ~x773 & ~x775 & ~x779 & ~x780 & ~x781 & ~x783;
assign c5208 =  x733;
assign c5210 = ~x1 & ~x3 & ~x4 & ~x5 & ~x6 & ~x7 & ~x9 & ~x10 & ~x11 & ~x12 & ~x13 & ~x14 & ~x15 & ~x16 & ~x19 & ~x20 & ~x21 & ~x25 & ~x26 & ~x27 & ~x28 & ~x29 & ~x30 & ~x34 & ~x35 & ~x39 & ~x41 & ~x42 & ~x43 & ~x45 & ~x47 & ~x48 & ~x49 & ~x52 & ~x53 & ~x56 & ~x59 & ~x61 & ~x62 & ~x63 & ~x64 & ~x66 & ~x67 & ~x72 & ~x78 & ~x79 & ~x80 & ~x81 & ~x82 & ~x84 & ~x85 & ~x86 & ~x88 & ~x90 & ~x94 & ~x97 & ~x108 & ~x113 & ~x116 & ~x117 & ~x118 & ~x119 & ~x120 & ~x122 & ~x123 & ~x124 & ~x139 & ~x141 & ~x144 & ~x145 & ~x146 & ~x148 & ~x149 & ~x165 & ~x170 & ~x171 & ~x172 & ~x173 & ~x174 & ~x175 & ~x176 & ~x191 & ~x192 & ~x193 & ~x195 & ~x198 & ~x199 & ~x200 & ~x203 & ~x220 & ~x222 & ~x227 & ~x230 & ~x231 & ~x232 & ~x248 & ~x249 & ~x250 & ~x251 & ~x252 & ~x253 & ~x254 & ~x255 & ~x257 & ~x259 & ~x260 & ~x277 & ~x279 & ~x283 & ~x284 & ~x287 & ~x298 & ~x299 & ~x300 & ~x301 & ~x306 & ~x307 & ~x308 & ~x309 & ~x311 & ~x312 & ~x313 & ~x314 & ~x331 & ~x335 & ~x336 & ~x337 & ~x338 & ~x341 & ~x342 & ~x359 & ~x360 & ~x361 & ~x365 & ~x366 & ~x367 & ~x368 & ~x371 & ~x387 & ~x388 & ~x389 & ~x394 & ~x395 & ~x398 & ~x399 & ~x416 & ~x421 & ~x425 & ~x443 & ~x462 & ~x463 & ~x475 & ~x477 & ~x486 & ~x488 & ~x489 & ~x491 & ~x499 & ~x500 & ~x501 & ~x502 & ~x503 & ~x504 & ~x505 & ~x528 & ~x530 & ~x531 & ~x532 & ~x533 & ~x534 & ~x558 & ~x560 & ~x561 & ~x563 & ~x582 & ~x584 & ~x585 & ~x586 & ~x588 & ~x589 & ~x590 & ~x593 & ~x608 & ~x609 & ~x612 & ~x614 & ~x615 & ~x618 & ~x620 & ~x638 & ~x641 & ~x643 & ~x644 & ~x645 & ~x646 & ~x647 & ~x649 & ~x661 & ~x662 & ~x669 & ~x670 & ~x672 & ~x673 & ~x674 & ~x675 & ~x676 & ~x678 & ~x691 & ~x692 & ~x693 & ~x694 & ~x696 & ~x707 & ~x711 & ~x715 & ~x717 & ~x720 & ~x721 & ~x722 & ~x723 & ~x727 & ~x728 & ~x729 & ~x733 & ~x734 & ~x736 & ~x738 & ~x739 & ~x743 & ~x744 & ~x746 & ~x747 & ~x748 & ~x749 & ~x750 & ~x751 & ~x752 & ~x753 & ~x755 & ~x756 & ~x758 & ~x759 & ~x762 & ~x769 & ~x770 & ~x772 & ~x773 & ~x774 & ~x775 & ~x777 & ~x778 & ~x779 & ~x782 & ~x783;
assign c5212 =  x272 & ~x25 & ~x27 & ~x100 & ~x103 & ~x122 & ~x140 & ~x161 & ~x164 & ~x174 & ~x187 & ~x188 & ~x227 & ~x357 & ~x359 & ~x384 & ~x420 & ~x470 & ~x530 & ~x589 & ~x648 & ~x671 & ~x723 & ~x737 & ~x743;
assign c5214 =  x235 &  x263 &  x292 &  x656 & ~x15 & ~x18 & ~x25 & ~x70 & ~x74 & ~x75 & ~x94 & ~x103 & ~x116 & ~x120 & ~x148 & ~x171 & ~x228 & ~x229 & ~x231 & ~x247 & ~x272 & ~x283 & ~x340 & ~x341 & ~x366 & ~x387 & ~x423 & ~x446 & ~x450 & ~x474 & ~x476 & ~x477 & ~x518 & ~x533 & ~x534 & ~x558 & ~x559 & ~x582 & ~x584 & ~x586 & ~x589 & ~x616 & ~x636 & ~x637 & ~x644 & ~x666 & ~x668 & ~x676 & ~x691 & ~x730 & ~x744 & ~x755 & ~x783;
assign c5216 =  x314 &  x583;
assign c5218 =  x664 &  x690;
assign c5220 =  x135 & ~x401;
assign c5222 =  x263 &  x291 &  x319 &  x347 & ~x3 & ~x4 & ~x7 & ~x14 & ~x15 & ~x19 & ~x26 & ~x34 & ~x36 & ~x39 & ~x42 & ~x49 & ~x50 & ~x56 & ~x59 & ~x60 & ~x63 & ~x74 & ~x75 & ~x87 & ~x96 & ~x108 & ~x110 & ~x115 & ~x116 & ~x117 & ~x119 & ~x121 & ~x122 & ~x135 & ~x136 & ~x144 & ~x148 & ~x163 & ~x165 & ~x169 & ~x172 & ~x195 & ~x201 & ~x202 & ~x228 & ~x229 & ~x230 & ~x251 & ~x254 & ~x255 & ~x256 & ~x257 & ~x280 & ~x304 & ~x310 & ~x329 & ~x334 & ~x335 & ~x340 & ~x357 & ~x360 & ~x364 & ~x392 & ~x397 & ~x398 & ~x419 & ~x426 & ~x445 & ~x448 & ~x449 & ~x463 & ~x470 & ~x473 & ~x476 & ~x500 & ~x501 & ~x502 & ~x503 & ~x507 & ~x515 & ~x517 & ~x533 & ~x535 & ~x589 & ~x612 & ~x616 & ~x637 & ~x645 & ~x666 & ~x668 & ~x669 & ~x673 & ~x703 & ~x705 & ~x717 & ~x723 & ~x725 & ~x733 & ~x741 & ~x743 & ~x755 & ~x758 & ~x761 & ~x770 & ~x775 & ~x778 & ~x783;
assign c5224 =  x502;
assign c5226 =  x203 &  x344 &  x373 &  x526 & ~x269;
assign c5228 =  x656 & ~x0 & ~x2 & ~x4 & ~x5 & ~x6 & ~x10 & ~x17 & ~x18 & ~x20 & ~x23 & ~x25 & ~x27 & ~x31 & ~x32 & ~x43 & ~x44 & ~x45 & ~x47 & ~x49 & ~x51 & ~x52 & ~x53 & ~x54 & ~x56 & ~x59 & ~x61 & ~x68 & ~x71 & ~x73 & ~x75 & ~x78 & ~x80 & ~x81 & ~x82 & ~x83 & ~x88 & ~x89 & ~x93 & ~x94 & ~x95 & ~x96 & ~x97 & ~x98 & ~x99 & ~x101 & ~x102 & ~x103 & ~x104 & ~x109 & ~x113 & ~x114 & ~x115 & ~x117 & ~x119 & ~x120 & ~x121 & ~x135 & ~x136 & ~x137 & ~x139 & ~x140 & ~x142 & ~x143 & ~x146 & ~x147 & ~x164 & ~x168 & ~x170 & ~x171 & ~x173 & ~x193 & ~x194 & ~x195 & ~x197 & ~x200 & ~x201 & ~x219 & ~x221 & ~x225 & ~x227 & ~x228 & ~x230 & ~x239 & ~x240 & ~x241 & ~x242 & ~x243 & ~x244 & ~x245 & ~x246 & ~x247 & ~x250 & ~x252 & ~x253 & ~x254 & ~x255 & ~x272 & ~x274 & ~x279 & ~x280 & ~x281 & ~x282 & ~x301 & ~x302 & ~x308 & ~x330 & ~x331 & ~x332 & ~x333 & ~x336 & ~x337 & ~x339 & ~x360 & ~x363 & ~x364 & ~x392 & ~x396 & ~x397 & ~x420 & ~x423 & ~x424 & ~x446 & ~x447 & ~x448 & ~x473 & ~x501 & ~x502 & ~x503 & ~x507 & ~x529 & ~x530 & ~x531 & ~x532 & ~x556 & ~x557 & ~x558 & ~x559 & ~x562 & ~x583 & ~x589 & ~x590 & ~x610 & ~x612 & ~x613 & ~x614 & ~x618 & ~x637 & ~x639 & ~x640 & ~x642 & ~x644 & ~x645 & ~x665 & ~x666 & ~x667 & ~x668 & ~x672 & ~x676 & ~x677 & ~x680 & ~x690 & ~x691 & ~x694 & ~x695 & ~x698 & ~x703 & ~x704 & ~x706 & ~x713 & ~x716 & ~x718 & ~x721 & ~x722 & ~x725 & ~x726 & ~x733 & ~x734 & ~x736 & ~x737 & ~x739 & ~x742 & ~x744 & ~x746 & ~x748 & ~x750 & ~x752 & ~x754 & ~x755 & ~x758 & ~x759 & ~x760 & ~x761 & ~x762 & ~x764 & ~x766 & ~x767 & ~x768 & ~x771 & ~x772 & ~x773 & ~x776 & ~x781 & ~x783;
assign c5230 =  x232 &  x260 &  x288 &  x344 &  x497 &  x629 & ~x10 & ~x18 & ~x61 & ~x92 & ~x104 & ~x280 & ~x331 & ~x337 & ~x388 & ~x446 & ~x474 & ~x475 & ~x483 & ~x506 & ~x561 & ~x618 & ~x647 & ~x675 & ~x699 & ~x740 & ~x747 & ~x754 & ~x769;
assign c5232 = ~x75 & ~x104 & ~x125 & ~x127 & ~x153 & ~x157 & ~x158 & ~x206 & ~x224 & ~x225 & ~x234 & ~x262 & ~x314 & ~x381 & ~x386 & ~x387 & ~x467 & ~x468 & ~x526 & ~x535 & ~x618 & ~x636 & ~x719 & ~x723 & ~x732 & ~x738 & ~x773 & ~x778;
assign c5234 =  x178 &  x179 &  x206 &  x317 &  x606 &  x608 & ~x677;
assign c5236 =  x714 &  x717;
assign c5238 = ~x24 & ~x38 & ~x63 & ~x68 & ~x89 & ~x122 & ~x126 & ~x307 & ~x309 & ~x322 & ~x323 & ~x328 & ~x351 & ~x353 & ~x382 & ~x441 & ~x442 & ~x501 & ~x537 & ~x570 & ~x740 & ~x747 & ~x763;
assign c5240 =  x246 & ~x1 & ~x7 & ~x30 & ~x33 & ~x42 & ~x73 & ~x92 & ~x112 & ~x146 & ~x168 & ~x228 & ~x251 & ~x306 & ~x326 & ~x327 & ~x329 & ~x332 & ~x334 & ~x359 & ~x476 & ~x530 & ~x533 & ~x534 & ~x591 & ~x670 & ~x731 & ~x765 & ~x770;
assign c5242 =  x189 &  x190 &  x239 &  x240 & ~x33 & ~x40 & ~x69 & ~x172 & ~x224 & ~x226 & ~x307 & ~x329 & ~x330 & ~x331 & ~x365 & ~x394 & ~x478 & ~x668 & ~x671 & ~x728 & ~x736;
assign c5244 =  x304 &  x329 & ~x383;
assign c5246 = ~x2 & ~x3 & ~x7 & ~x11 & ~x17 & ~x20 & ~x22 & ~x24 & ~x27 & ~x32 & ~x39 & ~x41 & ~x47 & ~x51 & ~x55 & ~x59 & ~x62 & ~x69 & ~x73 & ~x75 & ~x82 & ~x92 & ~x97 & ~x101 & ~x102 & ~x104 & ~x108 & ~x109 & ~x112 & ~x121 & ~x125 & ~x128 & ~x131 & ~x136 & ~x137 & ~x150 & ~x167 & ~x170 & ~x171 & ~x172 & ~x174 & ~x177 & ~x178 & ~x197 & ~x199 & ~x201 & ~x202 & ~x203 & ~x229 & ~x231 & ~x232 & ~x250 & ~x256 & ~x258 & ~x282 & ~x283 & ~x286 & ~x307 & ~x310 & ~x311 & ~x335 & ~x336 & ~x339 & ~x351 & ~x353 & ~x355 & ~x365 & ~x366 & ~x381 & ~x382 & ~x383 & ~x385 & ~x386 & ~x389 & ~x391 & ~x392 & ~x396 & ~x422 & ~x423 & ~x425 & ~x440 & ~x442 & ~x443 & ~x445 & ~x446 & ~x452 & ~x471 & ~x475 & ~x497 & ~x498 & ~x500 & ~x501 & ~x524 & ~x530 & ~x531 & ~x533 & ~x553 & ~x562 & ~x587 & ~x588 & ~x611 & ~x614 & ~x618 & ~x636 & ~x638 & ~x643 & ~x648 & ~x664 & ~x665 & ~x671 & ~x674 & ~x675 & ~x676 & ~x677 & ~x678 & ~x689 & ~x690 & ~x697 & ~x698 & ~x706 & ~x707 & ~x715 & ~x718 & ~x726 & ~x729 & ~x734 & ~x735 & ~x742 & ~x744 & ~x751 & ~x753 & ~x768 & ~x770 & ~x774 & ~x777 & ~x781 & ~x783;
assign c5248 =  x520 & ~x11 & ~x103 & ~x124 & ~x131 & ~x175 & ~x254 & ~x311 & ~x323 & ~x328 & ~x381 & ~x383 & ~x385 & ~x439 & ~x442 & ~x525 & ~x695 & ~x737 & ~x759;
assign c5250 =  x268 & ~x10 & ~x13 & ~x16 & ~x22 & ~x25 & ~x30 & ~x43 & ~x55 & ~x66 & ~x82 & ~x84 & ~x107 & ~x130 & ~x134 & ~x141 & ~x143 & ~x147 & ~x160 & ~x173 & ~x176 & ~x184 & ~x255 & ~x279 & ~x282 & ~x334 & ~x354 & ~x356 & ~x367 & ~x387 & ~x411 & ~x416 & ~x419 & ~x424 & ~x448 & ~x468 & ~x498 & ~x555 & ~x610 & ~x615 & ~x621 & ~x672 & ~x675 & ~x702 & ~x704 & ~x722 & ~x733 & ~x736 & ~x763 & ~x781;
assign c5252 =  x316 &  x344 & ~x4 & ~x5 & ~x16 & ~x17 & ~x21 & ~x24 & ~x28 & ~x31 & ~x46 & ~x49 & ~x73 & ~x84 & ~x86 & ~x91 & ~x100 & ~x101 & ~x112 & ~x125 & ~x131 & ~x134 & ~x136 & ~x142 & ~x165 & ~x167 & ~x169 & ~x194 & ~x199 & ~x221 & ~x228 & ~x281 & ~x327 & ~x328 & ~x358 & ~x359 & ~x386 & ~x422 & ~x447 & ~x450 & ~x489 & ~x515 & ~x516 & ~x518 & ~x520 & ~x532 & ~x546 & ~x547 & ~x560 & ~x589 & ~x590 & ~x592 & ~x612 & ~x616 & ~x618 & ~x641 & ~x646 & ~x672 & ~x676 & ~x677 & ~x695 & ~x705 & ~x725 & ~x732 & ~x743 & ~x747 & ~x759 & ~x767 & ~x776;
assign c5254 =  x240 &  x243 & ~x6 & ~x36 & ~x60 & ~x63 & ~x64 & ~x78 & ~x117 & ~x135 & ~x172 & ~x177 & ~x201 & ~x326 & ~x333 & ~x337 & ~x356 & ~x357 & ~x365 & ~x386 & ~x413 & ~x414 & ~x422 & ~x447 & ~x479 & ~x553 & ~x671 & ~x739 & ~x761 & ~x762 & ~x778;
assign c5256 = ~x3 & ~x20 & ~x22 & ~x28 & ~x50 & ~x60 & ~x67 & ~x71 & ~x73 & ~x76 & ~x82 & ~x227 & ~x266 & ~x267 & ~x268 & ~x269 & ~x270 & ~x271 & ~x272 & ~x278 & ~x280 & ~x298 & ~x299 & ~x300 & ~x301 & ~x303 & ~x338 & ~x423 & ~x446 & ~x447 & ~x477 & ~x482 & ~x489 & ~x504 & ~x517 & ~x519 & ~x545 & ~x546 & ~x551 & ~x579 & ~x614 & ~x670 & ~x675 & ~x700 & ~x736 & ~x756 & ~x757 & ~x780;
assign c5258 =  x735;
assign c5260 =  x210 &  x213 &  x214 &  x215 &  x216 &  x237 & ~x2 & ~x5 & ~x16 & ~x19 & ~x22 & ~x27 & ~x35 & ~x36 & ~x39 & ~x41 & ~x50 & ~x52 & ~x57 & ~x58 & ~x61 & ~x62 & ~x66 & ~x69 & ~x76 & ~x87 & ~x91 & ~x94 & ~x100 & ~x106 & ~x109 & ~x111 & ~x121 & ~x136 & ~x171 & ~x193 & ~x199 & ~x227 & ~x228 & ~x253 & ~x254 & ~x277 & ~x278 & ~x329 & ~x330 & ~x332 & ~x337 & ~x338 & ~x362 & ~x363 & ~x389 & ~x393 & ~x394 & ~x422 & ~x423 & ~x445 & ~x447 & ~x448 & ~x450 & ~x516 & ~x529 & ~x531 & ~x545 & ~x546 & ~x557 & ~x561 & ~x563 & ~x587 & ~x591 & ~x640 & ~x641 & ~x643 & ~x646 & ~x676 & ~x701 & ~x719 & ~x723 & ~x724 & ~x735 & ~x736 & ~x739 & ~x740 & ~x742 & ~x747 & ~x756 & ~x759 & ~x763 & ~x765 & ~x766 & ~x768 & ~x773 & ~x774;
assign c5262 =  x224;
assign c5264 =  x267 &  x272 &  x293 & ~x158 & ~x159 & ~x384 & ~x386 & ~x678;
assign c5266 =  x184 & ~x0 & ~x3 & ~x4 & ~x6 & ~x8 & ~x9 & ~x10 & ~x12 & ~x13 & ~x15 & ~x17 & ~x20 & ~x21 & ~x24 & ~x28 & ~x30 & ~x31 & ~x32 & ~x34 & ~x35 & ~x36 & ~x37 & ~x40 & ~x45 & ~x48 & ~x50 & ~x52 & ~x53 & ~x54 & ~x55 & ~x57 & ~x60 & ~x62 & ~x63 & ~x65 & ~x66 & ~x68 & ~x69 & ~x70 & ~x71 & ~x72 & ~x73 & ~x76 & ~x77 & ~x81 & ~x82 & ~x83 & ~x85 & ~x87 & ~x89 & ~x91 & ~x93 & ~x94 & ~x95 & ~x100 & ~x106 & ~x111 & ~x112 & ~x113 & ~x116 & ~x117 & ~x118 & ~x120 & ~x134 & ~x136 & ~x138 & ~x139 & ~x140 & ~x141 & ~x142 & ~x166 & ~x167 & ~x169 & ~x170 & ~x172 & ~x173 & ~x194 & ~x195 & ~x196 & ~x197 & ~x198 & ~x199 & ~x201 & ~x220 & ~x223 & ~x224 & ~x226 & ~x227 & ~x246 & ~x247 & ~x251 & ~x252 & ~x253 & ~x255 & ~x268 & ~x269 & ~x270 & ~x271 & ~x272 & ~x273 & ~x274 & ~x275 & ~x277 & ~x278 & ~x279 & ~x282 & ~x283 & ~x300 & ~x303 & ~x304 & ~x305 & ~x307 & ~x309 & ~x310 & ~x311 & ~x330 & ~x331 & ~x332 & ~x333 & ~x335 & ~x337 & ~x359 & ~x360 & ~x361 & ~x363 & ~x389 & ~x392 & ~x395 & ~x417 & ~x419 & ~x421 & ~x445 & ~x446 & ~x447 & ~x448 & ~x449 & ~x450 & ~x475 & ~x476 & ~x477 & ~x479 & ~x486 & ~x487 & ~x488 & ~x501 & ~x503 & ~x504 & ~x505 & ~x509 & ~x510 & ~x529 & ~x533 & ~x534 & ~x538 & ~x557 & ~x558 & ~x560 & ~x561 & ~x562 & ~x585 & ~x586 & ~x588 & ~x590 & ~x591 & ~x614 & ~x618 & ~x619 & ~x640 & ~x642 & ~x643 & ~x645 & ~x667 & ~x668 & ~x671 & ~x672 & ~x674 & ~x675 & ~x695 & ~x696 & ~x699 & ~x700 & ~x701 & ~x704 & ~x706 & ~x707 & ~x708 & ~x710 & ~x711 & ~x713 & ~x714 & ~x716 & ~x719 & ~x720 & ~x721 & ~x722 & ~x723 & ~x725 & ~x726 & ~x728 & ~x730 & ~x733 & ~x734 & ~x737 & ~x739 & ~x740 & ~x742 & ~x743 & ~x744 & ~x745 & ~x747 & ~x748 & ~x749 & ~x750 & ~x756 & ~x759 & ~x763 & ~x764 & ~x765 & ~x766 & ~x768 & ~x769 & ~x771 & ~x772 & ~x774 & ~x779 & ~x781 & ~x782;
assign c5268 =  x326 &  x327 & ~x86 & ~x92 & ~x96 & ~x105 & ~x115 & ~x118 & ~x136 & ~x145 & ~x198 & ~x213 & ~x214 & ~x221 & ~x365 & ~x381 & ~x410 & ~x439 & ~x530 & ~x591 & ~x669 & ~x716 & ~x744 & ~x772;
assign c5270 = ~x2 & ~x7 & ~x8 & ~x11 & ~x22 & ~x27 & ~x28 & ~x29 & ~x30 & ~x33 & ~x35 & ~x42 & ~x43 & ~x44 & ~x49 & ~x50 & ~x56 & ~x58 & ~x59 & ~x60 & ~x62 & ~x69 & ~x76 & ~x77 & ~x83 & ~x85 & ~x86 & ~x91 & ~x94 & ~x96 & ~x104 & ~x105 & ~x106 & ~x108 & ~x110 & ~x111 & ~x115 & ~x120 & ~x125 & ~x136 & ~x140 & ~x143 & ~x144 & ~x172 & ~x173 & ~x195 & ~x197 & ~x200 & ~x201 & ~x202 & ~x223 & ~x225 & ~x227 & ~x228 & ~x230 & ~x252 & ~x253 & ~x278 & ~x280 & ~x308 & ~x313 & ~x339 & ~x341 & ~x365 & ~x368 & ~x394 & ~x395 & ~x397 & ~x417 & ~x422 & ~x424 & ~x425 & ~x434 & ~x435 & ~x438 & ~x444 & ~x446 & ~x447 & ~x448 & ~x464 & ~x465 & ~x466 & ~x477 & ~x479 & ~x494 & ~x499 & ~x521 & ~x522 & ~x526 & ~x528 & ~x529 & ~x533 & ~x534 & ~x555 & ~x556 & ~x560 & ~x564 & ~x583 & ~x584 & ~x610 & ~x615 & ~x619 & ~x641 & ~x644 & ~x645 & ~x664 & ~x666 & ~x667 & ~x669 & ~x673 & ~x674 & ~x675 & ~x692 & ~x694 & ~x701 & ~x702 & ~x703 & ~x704 & ~x706 & ~x716 & ~x717 & ~x718 & ~x722 & ~x724 & ~x729 & ~x730 & ~x731 & ~x749 & ~x750 & ~x751 & ~x755 & ~x759 & ~x761 & ~x764 & ~x765 & ~x771 & ~x773 & ~x775 & ~x779 & ~x783;
assign c5272 =  x188 &  x189 &  x213 &  x214 &  x216 & ~x273 & ~x274 & ~x300 & ~x303;
assign c5274 = ~x8 & ~x22 & ~x23 & ~x34 & ~x37 & ~x40 & ~x49 & ~x55 & ~x57 & ~x59 & ~x62 & ~x64 & ~x65 & ~x66 & ~x69 & ~x78 & ~x83 & ~x88 & ~x95 & ~x98 & ~x100 & ~x101 & ~x102 & ~x112 & ~x113 & ~x122 & ~x123 & ~x140 & ~x141 & ~x151 & ~x167 & ~x168 & ~x170 & ~x173 & ~x177 & ~x194 & ~x199 & ~x227 & ~x229 & ~x250 & ~x252 & ~x255 & ~x272 & ~x275 & ~x277 & ~x280 & ~x281 & ~x284 & ~x296 & ~x301 & ~x303 & ~x304 & ~x305 & ~x312 & ~x325 & ~x328 & ~x332 & ~x355 & ~x358 & ~x359 & ~x366 & ~x395 & ~x397 & ~x417 & ~x424 & ~x425 & ~x448 & ~x477 & ~x480 & ~x501 & ~x505 & ~x513 & ~x514 & ~x515 & ~x532 & ~x535 & ~x544 & ~x561 & ~x562 & ~x564 & ~x583 & ~x586 & ~x589 & ~x592 & ~x612 & ~x614 & ~x615 & ~x619 & ~x621 & ~x636 & ~x642 & ~x643 & ~x648 & ~x650 & ~x664 & ~x669 & ~x672 & ~x697 & ~x700 & ~x701 & ~x702 & ~x704 & ~x706 & ~x707 & ~x740 & ~x754 & ~x760 & ~x761 & ~x771 & ~x783;
assign c5276 =  x161 &  x162 & ~x18 & ~x23 & ~x24 & ~x41 & ~x52 & ~x59 & ~x68 & ~x97 & ~x118 & ~x119 & ~x170 & ~x202 & ~x225 & ~x245 & ~x247 & ~x249 & ~x250 & ~x271 & ~x272 & ~x275 & ~x301 & ~x302 & ~x330 & ~x418 & ~x694 & ~x750 & ~x781;
assign c5278 = ~x24 & ~x27 & ~x36 & ~x39 & ~x49 & ~x74 & ~x80 & ~x87 & ~x98 & ~x99 & ~x110 & ~x121 & ~x129 & ~x142 & ~x143 & ~x150 & ~x158 & ~x161 & ~x165 & ~x178 & ~x186 & ~x197 & ~x223 & ~x279 & ~x280 & ~x281 & ~x315 & ~x342 & ~x390 & ~x420 & ~x424 & ~x445 & ~x449 & ~x473 & ~x476 & ~x532 & ~x534 & ~x560 & ~x563 & ~x584 & ~x590 & ~x606 & ~x612 & ~x647 & ~x660 & ~x668 & ~x674 & ~x679 & ~x687 & ~x704 & ~x705 & ~x710 & ~x712 & ~x713 & ~x723 & ~x753 & ~x754 & ~x765 & ~x772;
assign c5280 =  x590;
assign c5282 = ~x2 & ~x18 & ~x24 & ~x26 & ~x30 & ~x34 & ~x35 & ~x39 & ~x40 & ~x42 & ~x43 & ~x49 & ~x50 & ~x69 & ~x72 & ~x76 & ~x79 & ~x89 & ~x90 & ~x109 & ~x120 & ~x138 & ~x139 & ~x142 & ~x146 & ~x147 & ~x193 & ~x198 & ~x199 & ~x222 & ~x224 & ~x225 & ~x250 & ~x255 & ~x257 & ~x266 & ~x267 & ~x268 & ~x271 & ~x273 & ~x278 & ~x282 & ~x295 & ~x296 & ~x298 & ~x302 & ~x304 & ~x330 & ~x335 & ~x338 & ~x357 & ~x362 & ~x363 & ~x390 & ~x418 & ~x423 & ~x425 & ~x426 & ~x450 & ~x456 & ~x457 & ~x474 & ~x479 & ~x500 & ~x501 & ~x505 & ~x506 & ~x516 & ~x517 & ~x518 & ~x519 & ~x531 & ~x532 & ~x561 & ~x586 & ~x589 & ~x611 & ~x614 & ~x617 & ~x639 & ~x665 & ~x673 & ~x691 & ~x695 & ~x699 & ~x706 & ~x714 & ~x716 & ~x719 & ~x721 & ~x722 & ~x723 & ~x732 & ~x736 & ~x739 & ~x742 & ~x749 & ~x753 & ~x754 & ~x762 & ~x771 & ~x775 & ~x778 & ~x779;
assign c5284 =  x218 &  x241 & ~x63 & ~x108 & ~x133 & ~x167 & ~x169 & ~x229 & ~x303 & ~x306 & ~x328 & ~x332 & ~x357 & ~x413 & ~x535 & ~x771;
assign c5286 =  x248;
assign c5288 =  x207 &  x235 &  x262 &  x318 & ~x7 & ~x9 & ~x17 & ~x19 & ~x20 & ~x25 & ~x27 & ~x33 & ~x37 & ~x41 & ~x46 & ~x57 & ~x60 & ~x61 & ~x70 & ~x71 & ~x86 & ~x88 & ~x89 & ~x93 & ~x97 & ~x99 & ~x100 & ~x104 & ~x105 & ~x110 & ~x118 & ~x120 & ~x144 & ~x148 & ~x166 & ~x169 & ~x170 & ~x173 & ~x174 & ~x192 & ~x198 & ~x200 & ~x202 & ~x219 & ~x220 & ~x222 & ~x226 & ~x229 & ~x251 & ~x254 & ~x274 & ~x281 & ~x298 & ~x299 & ~x301 & ~x309 & ~x330 & ~x331 & ~x335 & ~x336 & ~x337 & ~x339 & ~x362 & ~x365 & ~x368 & ~x390 & ~x391 & ~x397 & ~x417 & ~x419 & ~x427 & ~x443 & ~x445 & ~x446 & ~x453 & ~x454 & ~x455 & ~x471 & ~x474 & ~x478 & ~x501 & ~x502 & ~x505 & ~x506 & ~x517 & ~x529 & ~x531 & ~x534 & ~x558 & ~x559 & ~x560 & ~x584 & ~x586 & ~x587 & ~x588 & ~x589 & ~x590 & ~x614 & ~x616 & ~x640 & ~x644 & ~x646 & ~x689 & ~x694 & ~x700 & ~x701 & ~x704 & ~x716 & ~x720 & ~x721 & ~x722 & ~x724 & ~x733 & ~x734 & ~x738 & ~x747 & ~x748 & ~x749 & ~x750 & ~x756 & ~x757 & ~x768 & ~x772 & ~x780 & ~x781;
assign c5290 = ~x25 & ~x30 & ~x31 & ~x63 & ~x65 & ~x66 & ~x69 & ~x75 & ~x96 & ~x111 & ~x117 & ~x143 & ~x164 & ~x165 & ~x187 & ~x238 & ~x241 & ~x242 & ~x244 & ~x309 & ~x339 & ~x407 & ~x437 & ~x445 & ~x521 & ~x559 & ~x616 & ~x641 & ~x646 & ~x665 & ~x666 & ~x667 & ~x670 & ~x676 & ~x713 & ~x714 & ~x719 & ~x722 & ~x746 & ~x765;
assign c5292 =  x136;
assign c5294 =  x390;
assign c5296 = ~x1 & ~x2 & ~x12 & ~x15 & ~x17 & ~x19 & ~x20 & ~x31 & ~x32 & ~x40 & ~x44 & ~x48 & ~x50 & ~x56 & ~x57 & ~x59 & ~x60 & ~x62 & ~x65 & ~x68 & ~x69 & ~x82 & ~x86 & ~x89 & ~x107 & ~x111 & ~x116 & ~x118 & ~x120 & ~x136 & ~x139 & ~x141 & ~x148 & ~x164 & ~x192 & ~x197 & ~x222 & ~x224 & ~x249 & ~x251 & ~x277 & ~x282 & ~x294 & ~x295 & ~x296 & ~x302 & ~x310 & ~x327 & ~x328 & ~x330 & ~x338 & ~x339 & ~x357 & ~x361 & ~x363 & ~x391 & ~x394 & ~x415 & ~x423 & ~x458 & ~x461 & ~x462 & ~x477 & ~x488 & ~x491 & ~x502 & ~x505 & ~x533 & ~x557 & ~x558 & ~x559 & ~x561 & ~x586 & ~x588 & ~x589 & ~x614 & ~x615 & ~x620 & ~x643 & ~x647 & ~x650 & ~x668 & ~x670 & ~x675 & ~x679 & ~x681 & ~x682 & ~x685 & ~x694 & ~x701 & ~x703 & ~x717 & ~x725 & ~x726 & ~x727 & ~x729 & ~x737 & ~x742 & ~x745 & ~x750 & ~x759 & ~x761 & ~x772 & ~x773 & ~x776 & ~x778 & ~x780 & ~x782;
assign c5298 =  x216 &  x239 &  x240 & ~x3 & ~x4 & ~x7 & ~x8 & ~x12 & ~x18 & ~x23 & ~x35 & ~x37 & ~x50 & ~x53 & ~x56 & ~x65 & ~x75 & ~x77 & ~x82 & ~x84 & ~x85 & ~x86 & ~x87 & ~x90 & ~x91 & ~x98 & ~x100 & ~x107 & ~x111 & ~x113 & ~x115 & ~x126 & ~x131 & ~x132 & ~x223 & ~x250 & ~x256 & ~x273 & ~x274 & ~x276 & ~x277 & ~x282 & ~x283 & ~x306 & ~x307 & ~x308 & ~x328 & ~x329 & ~x336 & ~x357 & ~x389 & ~x391 & ~x392 & ~x393 & ~x421 & ~x451 & ~x474 & ~x476 & ~x504 & ~x505 & ~x507 & ~x529 & ~x556 & ~x559 & ~x561 & ~x586 & ~x587 & ~x643 & ~x644 & ~x672 & ~x698 & ~x699 & ~x701 & ~x721 & ~x726 & ~x727 & ~x729 & ~x730 & ~x754 & ~x758 & ~x759 & ~x761 & ~x762 & ~x764 & ~x765 & ~x771 & ~x777;
assign c51 =  x267 &  x294 & ~x1 & ~x4 & ~x8 & ~x9 & ~x12 & ~x13 & ~x19 & ~x20 & ~x21 & ~x23 & ~x31 & ~x33 & ~x35 & ~x36 & ~x37 & ~x48 & ~x53 & ~x55 & ~x61 & ~x64 & ~x65 & ~x68 & ~x72 & ~x73 & ~x77 & ~x86 & ~x89 & ~x102 & ~x105 & ~x111 & ~x113 & ~x117 & ~x131 & ~x133 & ~x134 & ~x136 & ~x144 & ~x159 & ~x167 & ~x168 & ~x170 & ~x171 & ~x172 & ~x187 & ~x188 & ~x189 & ~x217 & ~x218 & ~x220 & ~x223 & ~x244 & ~x245 & ~x246 & ~x247 & ~x251 & ~x253 & ~x254 & ~x271 & ~x273 & ~x275 & ~x279 & ~x281 & ~x298 & ~x301 & ~x304 & ~x306 & ~x328 & ~x329 & ~x331 & ~x333 & ~x338 & ~x362 & ~x365 & ~x392 & ~x393 & ~x396 & ~x397 & ~x423 & ~x454 & ~x474 & ~x501 & ~x505 & ~x510 & ~x511 & ~x531 & ~x559 & ~x560 & ~x565 & ~x585 & ~x588 & ~x591 & ~x592 & ~x611 & ~x614 & ~x638 & ~x673 & ~x693 & ~x706 & ~x710 & ~x721 & ~x728 & ~x732 & ~x735 & ~x741 & ~x751 & ~x753 & ~x756 & ~x767 & ~x774 & ~x776 & ~x777 & ~x779 & ~x780 & ~x782;
assign c53 =  x242 &  x270 &  x298 &  x325 & ~x13 & ~x15 & ~x22 & ~x28 & ~x34 & ~x39 & ~x40 & ~x61 & ~x62 & ~x66 & ~x71 & ~x83 & ~x86 & ~x95 & ~x96 & ~x104 & ~x108 & ~x136 & ~x138 & ~x142 & ~x192 & ~x194 & ~x196 & ~x218 & ~x226 & ~x248 & ~x252 & ~x274 & ~x275 & ~x276 & ~x278 & ~x282 & ~x302 & ~x333 & ~x335 & ~x359 & ~x362 & ~x364 & ~x415 & ~x417 & ~x446 & ~x447 & ~x449 & ~x476 & ~x503 & ~x557 & ~x588 & ~x616 & ~x641 & ~x642 & ~x669 & ~x696 & ~x704 & ~x705 & ~x750 & ~x751 & ~x757 & ~x761 & ~x766 & ~x771 & ~x779 & ~x782 & ~x783;
assign c55 =  x324 &  x351 & ~x9 & ~x11 & ~x16 & ~x33 & ~x43 & ~x68 & ~x78 & ~x87 & ~x102 & ~x103 & ~x167 & ~x225 & ~x247 & ~x249 & ~x255 & ~x275 & ~x276 & ~x278 & ~x327 & ~x331 & ~x354 & ~x362 & ~x364 & ~x427 & ~x444 & ~x483 & ~x532 & ~x558 & ~x614 & ~x621 & ~x641 & ~x671 & ~x700 & ~x741 & ~x751 & ~x769 & ~x781;
assign c57 =  x271 &  x299 &  x326 &  x353 & ~x16 & ~x22 & ~x24 & ~x31 & ~x35 & ~x37 & ~x40 & ~x45 & ~x51 & ~x66 & ~x92 & ~x95 & ~x102 & ~x105 & ~x106 & ~x115 & ~x116 & ~x140 & ~x174 & ~x221 & ~x223 & ~x249 & ~x281 & ~x282 & ~x303 & ~x333 & ~x359 & ~x363 & ~x424 & ~x451 & ~x473 & ~x584 & ~x589 & ~x700 & ~x701 & ~x703 & ~x722 & ~x726 & ~x728 & ~x735 & ~x744 & ~x753 & ~x776;
assign c59 =  x352 & ~x10 & ~x15 & ~x20 & ~x23 & ~x26 & ~x27 & ~x36 & ~x39 & ~x43 & ~x53 & ~x56 & ~x60 & ~x81 & ~x82 & ~x87 & ~x90 & ~x94 & ~x100 & ~x117 & ~x166 & ~x168 & ~x170 & ~x173 & ~x194 & ~x200 & ~x222 & ~x226 & ~x229 & ~x303 & ~x307 & ~x336 & ~x341 & ~x361 & ~x367 & ~x368 & ~x391 & ~x395 & ~x396 & ~x414 & ~x416 & ~x426 & ~x441 & ~x445 & ~x446 & ~x476 & ~x478 & ~x482 & ~x498 & ~x503 & ~x524 & ~x528 & ~x529 & ~x530 & ~x531 & ~x555 & ~x588 & ~x612 & ~x615 & ~x666 & ~x671 & ~x694 & ~x697 & ~x700 & ~x702 & ~x706 & ~x721 & ~x724 & ~x736 & ~x746 & ~x748 & ~x754 & ~x756 & ~x762 & ~x765;
assign c511 =  x96;
assign c513 =  x149 &  x350 & ~x260 & ~x286;
assign c515 =  x458 &  x514 &  x542 & ~x22 & ~x89 & ~x140 & ~x290 & ~x361 & ~x396 & ~x425 & ~x426 & ~x566 & ~x645 & ~x674 & ~x702 & ~x737 & ~x756 & ~x772;
assign c517 =  x350 & ~x59 & ~x66 & ~x159 & ~x275 & ~x371 & ~x384 & ~x509 & ~x511;
assign c519 =  x326 & ~x1 & ~x2 & ~x8 & ~x11 & ~x14 & ~x15 & ~x18 & ~x22 & ~x23 & ~x24 & ~x32 & ~x35 & ~x36 & ~x37 & ~x38 & ~x48 & ~x54 & ~x58 & ~x61 & ~x62 & ~x63 & ~x64 & ~x65 & ~x69 & ~x71 & ~x72 & ~x76 & ~x78 & ~x81 & ~x83 & ~x84 & ~x85 & ~x86 & ~x88 & ~x89 & ~x90 & ~x106 & ~x108 & ~x113 & ~x116 & ~x117 & ~x118 & ~x135 & ~x139 & ~x145 & ~x146 & ~x169 & ~x196 & ~x198 & ~x202 & ~x227 & ~x229 & ~x251 & ~x253 & ~x254 & ~x255 & ~x256 & ~x277 & ~x279 & ~x283 & ~x284 & ~x295 & ~x296 & ~x306 & ~x309 & ~x331 & ~x335 & ~x337 & ~x340 & ~x357 & ~x362 & ~x390 & ~x394 & ~x418 & ~x419 & ~x420 & ~x421 & ~x442 & ~x447 & ~x475 & ~x476 & ~x479 & ~x504 & ~x506 & ~x530 & ~x531 & ~x532 & ~x533 & ~x534 & ~x558 & ~x561 & ~x588 & ~x644 & ~x669 & ~x670 & ~x672 & ~x673 & ~x676 & ~x679 & ~x697 & ~x698 & ~x704 & ~x721 & ~x724 & ~x726 & ~x728 & ~x732 & ~x736 & ~x742 & ~x744 & ~x745 & ~x748 & ~x751 & ~x755 & ~x756 & ~x765 & ~x766 & ~x768 & ~x769 & ~x773 & ~x782;
assign c521 = ~x16 & ~x24 & ~x26 & ~x27 & ~x32 & ~x48 & ~x55 & ~x63 & ~x77 & ~x89 & ~x96 & ~x132 & ~x136 & ~x159 & ~x172 & ~x246 & ~x247 & ~x303 & ~x330 & ~x333 & ~x357 & ~x367 & ~x387 & ~x413 & ~x425 & ~x445 & ~x503 & ~x507 & ~x510 & ~x538 & ~x567 & ~x619 & ~x622 & ~x626 & ~x627 & ~x696 & ~x758 & ~x766;
assign c523 =  x297 &  x352 &  x380 & ~x6 & ~x10 & ~x27 & ~x34 & ~x80 & ~x103 & ~x112 & ~x114 & ~x116 & ~x169 & ~x191 & ~x220 & ~x248 & ~x274 & ~x303 & ~x305 & ~x310 & ~x360 & ~x363 & ~x415 & ~x416 & ~x418 & ~x443 & ~x474 & ~x504 & ~x539 & ~x583 & ~x668 & ~x673 & ~x696 & ~x704 & ~x727 & ~x758 & ~x774;
assign c525 =  x358 &  x455 &  x511;
assign c527 =  x434 & ~x1 & ~x34 & ~x37 & ~x52 & ~x68 & ~x103 & ~x109 & ~x141 & ~x194 & ~x254 & ~x279 & ~x304 & ~x331 & ~x412 & ~x440 & ~x441 & ~x481 & ~x529 & ~x647 & ~x743 & ~x751 & ~x759;
assign c529 =  x439 & ~x151 & ~x326 & ~x352 & ~x607;
assign c531 = ~x2 & ~x7 & ~x15 & ~x16 & ~x32 & ~x36 & ~x47 & ~x54 & ~x56 & ~x80 & ~x84 & ~x108 & ~x109 & ~x112 & ~x135 & ~x137 & ~x138 & ~x139 & ~x149 & ~x164 & ~x168 & ~x171 & ~x176 & ~x186 & ~x187 & ~x188 & ~x193 & ~x197 & ~x198 & ~x215 & ~x272 & ~x275 & ~x278 & ~x305 & ~x306 & ~x329 & ~x341 & ~x359 & ~x365 & ~x366 & ~x368 & ~x369 & ~x370 & ~x390 & ~x416 & ~x418 & ~x420 & ~x423 & ~x447 & ~x449 & ~x501 & ~x502 & ~x508 & ~x533 & ~x538 & ~x539 & ~x559 & ~x564 & ~x565 & ~x585 & ~x592 & ~x593 & ~x609 & ~x614 & ~x624 & ~x625 & ~x626 & ~x638 & ~x645 & ~x651 & ~x653 & ~x655 & ~x665 & ~x675 & ~x687 & ~x697 & ~x703 & ~x708 & ~x726 & ~x729 & ~x746 & ~x749 & ~x753 & ~x754 & ~x759 & ~x767 & ~x782;
assign c533 =  x439 & ~x30 & ~x36 & ~x38 & ~x65 & ~x71 & ~x85 & ~x86 & ~x96 & ~x126 & ~x137 & ~x188 & ~x189 & ~x193 & ~x196 & ~x222 & ~x245 & ~x247 & ~x261 & ~x281 & ~x331 & ~x361 & ~x500 & ~x535 & ~x538 & ~x644 & ~x675 & ~x678 & ~x701 & ~x709 & ~x762 & ~x765;
assign c535 =  x287 &  x296 & ~x346;
assign c537 = ~x0 & ~x6 & ~x7 & ~x15 & ~x22 & ~x32 & ~x34 & ~x36 & ~x44 & ~x52 & ~x59 & ~x61 & ~x88 & ~x90 & ~x91 & ~x92 & ~x111 & ~x117 & ~x137 & ~x141 & ~x170 & ~x175 & ~x201 & ~x225 & ~x226 & ~x228 & ~x252 & ~x325 & ~x351 & ~x389 & ~x405 & ~x406 & ~x417 & ~x418 & ~x450 & ~x459 & ~x473 & ~x476 & ~x477 & ~x479 & ~x487 & ~x535 & ~x589 & ~x641 & ~x646 & ~x677 & ~x695 & ~x701 & ~x705 & ~x706 & ~x707 & ~x724 & ~x729 & ~x730 & ~x740 & ~x748 & ~x751 & ~x763 & ~x768 & ~x770 & ~x771 & ~x772;
assign c539 =  x272 &  x328 & ~x22 & ~x37 & ~x46 & ~x48 & ~x90 & ~x111 & ~x136 & ~x138 & ~x166 & ~x173 & ~x278 & ~x304 & ~x305 & ~x307 & ~x332 & ~x451 & ~x476 & ~x533 & ~x554 & ~x611 & ~x613 & ~x641 & ~x642 & ~x702 & ~x706 & ~x724 & ~x728 & ~x742 & ~x746 & ~x783;
assign c541 =  x228;
assign c543 =  x269 &  x296 &  x351 & ~x0 & ~x8 & ~x15 & ~x18 & ~x27 & ~x29 & ~x30 & ~x33 & ~x48 & ~x52 & ~x73 & ~x85 & ~x99 & ~x101 & ~x133 & ~x136 & ~x138 & ~x164 & ~x171 & ~x195 & ~x198 & ~x201 & ~x226 & ~x246 & ~x248 & ~x254 & ~x274 & ~x301 & ~x303 & ~x304 & ~x305 & ~x308 & ~x336 & ~x356 & ~x365 & ~x389 & ~x390 & ~x396 & ~x421 & ~x446 & ~x472 & ~x474 & ~x480 & ~x499 & ~x530 & ~x534 & ~x557 & ~x559 & ~x563 & ~x588 & ~x592 & ~x613 & ~x614 & ~x697 & ~x701 & ~x718 & ~x728 & ~x729 & ~x735 & ~x737 & ~x744 & ~x750 & ~x769 & ~x773 & ~x774 & ~x777 & ~x779;
assign c545 =  x436 &  x489 &  x516 &  x517 & ~x3 & ~x4 & ~x20 & ~x33 & ~x63 & ~x222 & ~x365 & ~x449 & ~x536 & ~x621 & ~x642 & ~x760;
assign c547 =  x295 &  x323 &  x406 & ~x2 & ~x5 & ~x65 & ~x103 & ~x218 & ~x273 & ~x274 & ~x279 & ~x281 & ~x301 & ~x304 & ~x338 & ~x365 & ~x388 & ~x480 & ~x510 & ~x562 & ~x589 & ~x617 & ~x724 & ~x727 & ~x754 & ~x755 & ~x768 & ~x776 & ~x778;
assign c549 =  x516 &  x544 & ~x172 & ~x248 & ~x251 & ~x394 & ~x396 & ~x511 & ~x540 & ~x582 & ~x622 & ~x703;
assign c551 =  x456 &  x597 & ~x194 & ~x323 & ~x351 & ~x390 & ~x585 & ~x710 & ~x727 & ~x744;
assign c553 = ~x4 & ~x5 & ~x10 & ~x12 & ~x15 & ~x18 & ~x22 & ~x27 & ~x30 & ~x34 & ~x38 & ~x39 & ~x40 & ~x43 & ~x48 & ~x51 & ~x61 & ~x67 & ~x69 & ~x79 & ~x82 & ~x94 & ~x96 & ~x98 & ~x129 & ~x131 & ~x132 & ~x134 & ~x138 & ~x145 & ~x159 & ~x162 & ~x187 & ~x188 & ~x194 & ~x195 & ~x218 & ~x222 & ~x225 & ~x226 & ~x244 & ~x245 & ~x246 & ~x271 & ~x273 & ~x274 & ~x277 & ~x300 & ~x301 & ~x302 & ~x303 & ~x304 & ~x305 & ~x306 & ~x307 & ~x310 & ~x311 & ~x327 & ~x339 & ~x340 & ~x358 & ~x360 & ~x388 & ~x393 & ~x416 & ~x418 & ~x424 & ~x427 & ~x448 & ~x449 & ~x454 & ~x474 & ~x478 & ~x483 & ~x503 & ~x505 & ~x506 & ~x507 & ~x513 & ~x516 & ~x528 & ~x530 & ~x535 & ~x542 & ~x556 & ~x559 & ~x560 & ~x566 & ~x587 & ~x592 & ~x593 & ~x610 & ~x611 & ~x636 & ~x639 & ~x640 & ~x646 & ~x648 & ~x666 & ~x669 & ~x672 & ~x673 & ~x674 & ~x675 & ~x692 & ~x695 & ~x696 & ~x702 & ~x707 & ~x708 & ~x709 & ~x710 & ~x721 & ~x724 & ~x725 & ~x730 & ~x732 & ~x741 & ~x747 & ~x750 & ~x753 & ~x754 & ~x755 & ~x759 & ~x763 & ~x776 & ~x780;
assign c555 =  x300 &  x328 &  x383 & ~x8 & ~x39 & ~x45 & ~x48 & ~x49 & ~x56 & ~x73 & ~x74 & ~x89 & ~x117 & ~x138 & ~x338 & ~x360 & ~x361 & ~x389 & ~x421 & ~x447 & ~x449 & ~x502 & ~x504 & ~x616 & ~x669 & ~x674 & ~x693 & ~x697 & ~x726 & ~x728 & ~x729 & ~x730 & ~x748 & ~x749 & ~x752 & ~x753 & ~x758 & ~x773 & ~x775 & ~x779;
assign c557 =  x407 &  x433 &  x488 & ~x3 & ~x4 & ~x21 & ~x37 & ~x80 & ~x81 & ~x108 & ~x116 & ~x121 & ~x195 & ~x256 & ~x468 & ~x477 & ~x510 & ~x537 & ~x669 & ~x697 & ~x720 & ~x728 & ~x729 & ~x733;
assign c559 =  x501;
assign c561 =  x432 &  x459 &  x513 & ~x2 & ~x12 & ~x16 & ~x22 & ~x41 & ~x54 & ~x58 & ~x60 & ~x61 & ~x73 & ~x77 & ~x80 & ~x82 & ~x83 & ~x86 & ~x88 & ~x92 & ~x93 & ~x112 & ~x167 & ~x283 & ~x284 & ~x315 & ~x340 & ~x391 & ~x392 & ~x394 & ~x426 & ~x477 & ~x504 & ~x507 & ~x562 & ~x563 & ~x649 & ~x670 & ~x699 & ~x701 & ~x716 & ~x717 & ~x737 & ~x739 & ~x747 & ~x752 & ~x781;
assign c563 = ~x1 & ~x8 & ~x10 & ~x12 & ~x14 & ~x26 & ~x34 & ~x40 & ~x54 & ~x56 & ~x62 & ~x78 & ~x90 & ~x93 & ~x109 & ~x113 & ~x116 & ~x123 & ~x133 & ~x139 & ~x140 & ~x148 & ~x157 & ~x162 & ~x163 & ~x166 & ~x168 & ~x185 & ~x218 & ~x219 & ~x244 & ~x273 & ~x275 & ~x278 & ~x281 & ~x301 & ~x303 & ~x304 & ~x305 & ~x309 & ~x335 & ~x339 & ~x362 & ~x364 & ~x423 & ~x427 & ~x480 & ~x502 & ~x505 & ~x510 & ~x511 & ~x512 & ~x529 & ~x538 & ~x556 & ~x561 & ~x562 & ~x568 & ~x597 & ~x654 & ~x666 & ~x669 & ~x670 & ~x673 & ~x674 & ~x699 & ~x709 & ~x722 & ~x730 & ~x751 & ~x752 & ~x758 & ~x759 & ~x767 & ~x771 & ~x776;
assign c565 =  x486 &  x514 &  x542 & ~x2 & ~x4 & ~x18 & ~x27 & ~x33 & ~x34 & ~x46 & ~x47 & ~x50 & ~x57 & ~x61 & ~x67 & ~x110 & ~x113 & ~x138 & ~x162 & ~x168 & ~x195 & ~x196 & ~x200 & ~x226 & ~x227 & ~x249 & ~x253 & ~x254 & ~x255 & ~x257 & ~x276 & ~x360 & ~x364 & ~x390 & ~x394 & ~x395 & ~x423 & ~x504 & ~x532 & ~x533 & ~x556 & ~x559 & ~x565 & ~x583 & ~x587 & ~x589 & ~x616 & ~x621 & ~x635 & ~x637 & ~x645 & ~x650 & ~x668 & ~x690 & ~x691 & ~x695 & ~x700 & ~x702 & ~x713 & ~x719 & ~x720 & ~x726 & ~x729 & ~x734 & ~x740 & ~x772 & ~x773 & ~x778;
assign c567 = ~x18 & ~x20 & ~x33 & ~x34 & ~x44 & ~x45 & ~x53 & ~x57 & ~x69 & ~x71 & ~x74 & ~x76 & ~x83 & ~x96 & ~x97 & ~x110 & ~x126 & ~x128 & ~x158 & ~x160 & ~x163 & ~x165 & ~x195 & ~x214 & ~x243 & ~x270 & ~x271 & ~x272 & ~x280 & ~x299 & ~x304 & ~x332 & ~x333 & ~x338 & ~x419 & ~x425 & ~x483 & ~x484 & ~x511 & ~x514 & ~x528 & ~x529 & ~x562 & ~x564 & ~x565 & ~x585 & ~x589 & ~x594 & ~x612 & ~x619 & ~x641 & ~x643 & ~x666 & ~x674 & ~x678 & ~x696 & ~x705 & ~x706 & ~x710 & ~x713 & ~x731 & ~x735 & ~x741 & ~x766 & ~x770 & ~x777;
assign c569 =  x462 &  x487 &  x514 & ~x8 & ~x31 & ~x84 & ~x254 & ~x503 & ~x641 & ~x660 & ~x712 & ~x742;
assign c571 = ~x0 & ~x4 & ~x6 & ~x8 & ~x9 & ~x10 & ~x12 & ~x14 & ~x17 & ~x20 & ~x26 & ~x31 & ~x35 & ~x36 & ~x43 & ~x44 & ~x49 & ~x54 & ~x57 & ~x64 & ~x65 & ~x66 & ~x67 & ~x69 & ~x74 & ~x77 & ~x78 & ~x84 & ~x85 & ~x86 & ~x93 & ~x94 & ~x99 & ~x102 & ~x108 & ~x109 & ~x110 & ~x111 & ~x114 & ~x118 & ~x134 & ~x136 & ~x138 & ~x143 & ~x145 & ~x162 & ~x163 & ~x165 & ~x169 & ~x172 & ~x190 & ~x194 & ~x199 & ~x218 & ~x222 & ~x225 & ~x226 & ~x227 & ~x228 & ~x229 & ~x253 & ~x255 & ~x274 & ~x276 & ~x279 & ~x280 & ~x282 & ~x283 & ~x286 & ~x288 & ~x289 & ~x290 & ~x291 & ~x304 & ~x310 & ~x314 & ~x331 & ~x333 & ~x335 & ~x336 & ~x339 & ~x342 & ~x358 & ~x363 & ~x364 & ~x390 & ~x393 & ~x394 & ~x395 & ~x415 & ~x449 & ~x451 & ~x452 & ~x477 & ~x478 & ~x479 & ~x530 & ~x531 & ~x532 & ~x559 & ~x584 & ~x585 & ~x610 & ~x611 & ~x612 & ~x614 & ~x616 & ~x618 & ~x640 & ~x641 & ~x643 & ~x666 & ~x667 & ~x675 & ~x689 & ~x700 & ~x702 & ~x711 & ~x713 & ~x715 & ~x717 & ~x722 & ~x726 & ~x732 & ~x735 & ~x736 & ~x737 & ~x738 & ~x744 & ~x745 & ~x750 & ~x751 & ~x754 & ~x755 & ~x757 & ~x758 & ~x760 & ~x762 & ~x764 & ~x766 & ~x769 & ~x770 & ~x771 & ~x772 & ~x779 & ~x782;
assign c573 =  x434 &  x461 &  x488 &  x542 & ~x339 & ~x477 & ~x661 & ~x692 & ~x721 & ~x737;
assign c575 =  x355 &  x463 & ~x48 & ~x333 & ~x447 & ~x501 & ~x506 & ~x646 & ~x722;
assign c577 =  x357 & ~x85 & ~x323 & ~x376;
assign c579 =  x298 &  x354 & ~x330 & ~x333 & ~x358 & ~x598 & ~x625 & ~x651 & ~x775 & ~x779;
assign c581 =  x355 &  x409 & ~x104 & ~x138 & ~x306 & ~x324 & ~x351 & ~x366;
assign c583 = ~x6 & ~x32 & ~x44 & ~x65 & ~x73 & ~x87 & ~x94 & ~x101 & ~x131 & ~x135 & ~x157 & ~x159 & ~x160 & ~x162 & ~x186 & ~x215 & ~x216 & ~x246 & ~x272 & ~x273 & ~x303 & ~x304 & ~x339 & ~x346 & ~x347 & ~x359 & ~x388 & ~x451 & ~x505 & ~x506 & ~x507 & ~x563 & ~x589 & ~x619 & ~x643 & ~x735 & ~x760 & ~x771;
assign c585 =  x243 &  x271 & ~x5 & ~x8 & ~x139 & ~x193 & ~x194 & ~x220 & ~x229 & ~x247 & ~x254 & ~x257 & ~x292 & ~x474 & ~x558 & ~x585 & ~x637 & ~x715 & ~x718 & ~x723 & ~x756 & ~x764 & ~x766;
assign c587 = ~x0 & ~x3 & ~x9 & ~x12 & ~x15 & ~x19 & ~x20 & ~x23 & ~x31 & ~x42 & ~x80 & ~x83 & ~x89 & ~x92 & ~x95 & ~x107 & ~x109 & ~x112 & ~x113 & ~x117 & ~x119 & ~x120 & ~x122 & ~x135 & ~x143 & ~x146 & ~x162 & ~x163 & ~x164 & ~x166 & ~x168 & ~x176 & ~x177 & ~x178 & ~x188 & ~x189 & ~x190 & ~x192 & ~x196 & ~x200 & ~x204 & ~x205 & ~x217 & ~x218 & ~x227 & ~x248 & ~x249 & ~x254 & ~x276 & ~x304 & ~x306 & ~x331 & ~x332 & ~x360 & ~x364 & ~x367 & ~x389 & ~x391 & ~x393 & ~x418 & ~x420 & ~x446 & ~x449 & ~x451 & ~x452 & ~x473 & ~x476 & ~x480 & ~x503 & ~x504 & ~x506 & ~x507 & ~x509 & ~x559 & ~x586 & ~x589 & ~x590 & ~x591 & ~x592 & ~x595 & ~x608 & ~x618 & ~x620 & ~x621 & ~x623 & ~x624 & ~x625 & ~x626 & ~x627 & ~x636 & ~x644 & ~x646 & ~x649 & ~x655 & ~x663 & ~x668 & ~x669 & ~x672 & ~x681 & ~x690 & ~x696 & ~x701 & ~x708 & ~x709 & ~x710 & ~x717 & ~x728 & ~x735 & ~x740 & ~x746 & ~x749 & ~x751 & ~x762 & ~x763 & ~x775 & ~x776 & ~x778 & ~x780 & ~x781;
assign c589 =  x429 &  x457 &  x484 &  x540 & ~x0 & ~x18 & ~x20 & ~x22 & ~x30 & ~x52 & ~x58 & ~x59 & ~x79 & ~x80 & ~x84 & ~x87 & ~x112 & ~x137 & ~x141 & ~x142 & ~x144 & ~x147 & ~x165 & ~x166 & ~x167 & ~x168 & ~x194 & ~x197 & ~x199 & ~x221 & ~x227 & ~x249 & ~x283 & ~x284 & ~x307 & ~x313 & ~x335 & ~x337 & ~x361 & ~x367 & ~x370 & ~x389 & ~x398 & ~x416 & ~x425 & ~x453 & ~x500 & ~x505 & ~x506 & ~x535 & ~x561 & ~x587 & ~x615 & ~x616 & ~x646 & ~x663 & ~x674 & ~x686 & ~x705 & ~x707 & ~x712 & ~x713 & ~x725 & ~x730 & ~x738 & ~x751 & ~x753 & ~x761 & ~x762;
assign c591 =  x296 & ~x20 & ~x43 & ~x45 & ~x47 & ~x64 & ~x71 & ~x75 & ~x79 & ~x103 & ~x171 & ~x190 & ~x191 & ~x193 & ~x194 & ~x195 & ~x218 & ~x250 & ~x274 & ~x276 & ~x300 & ~x301 & ~x304 & ~x305 & ~x310 & ~x328 & ~x354 & ~x356 & ~x358 & ~x359 & ~x383 & ~x449 & ~x476 & ~x498 & ~x528 & ~x532 & ~x588 & ~x615 & ~x617 & ~x702 & ~x705 & ~x711 & ~x719 & ~x723 & ~x742 & ~x749 & ~x758 & ~x772 & ~x774 & ~x779 & ~x782;
assign c593 =  x454 & ~x226 & ~x351 & ~x377 & ~x405;
assign c595 = ~x0 & ~x1 & ~x4 & ~x6 & ~x8 & ~x10 & ~x15 & ~x18 & ~x23 & ~x31 & ~x32 & ~x35 & ~x47 & ~x61 & ~x80 & ~x81 & ~x100 & ~x104 & ~x111 & ~x114 & ~x129 & ~x132 & ~x134 & ~x135 & ~x137 & ~x139 & ~x160 & ~x166 & ~x168 & ~x172 & ~x187 & ~x189 & ~x194 & ~x198 & ~x199 & ~x215 & ~x255 & ~x261 & ~x273 & ~x274 & ~x279 & ~x284 & ~x285 & ~x300 & ~x302 & ~x303 & ~x306 & ~x312 & ~x327 & ~x330 & ~x332 & ~x341 & ~x343 & ~x363 & ~x364 & ~x367 & ~x371 & ~x388 & ~x389 & ~x398 & ~x421 & ~x443 & ~x445 & ~x447 & ~x448 & ~x449 & ~x474 & ~x481 & ~x486 & ~x498 & ~x506 & ~x537 & ~x561 & ~x565 & ~x587 & ~x615 & ~x622 & ~x639 & ~x643 & ~x644 & ~x645 & ~x646 & ~x668 & ~x669 & ~x678 & ~x704 & ~x708 & ~x718 & ~x720 & ~x729 & ~x738 & ~x745 & ~x747 & ~x750 & ~x754 & ~x772 & ~x773 & ~x782;
assign c597 = ~x28 & ~x37 & ~x38 & ~x43 & ~x48 & ~x52 & ~x70 & ~x74 & ~x91 & ~x99 & ~x102 & ~x103 & ~x108 & ~x111 & ~x112 & ~x113 & ~x120 & ~x140 & ~x160 & ~x161 & ~x217 & ~x220 & ~x255 & ~x264 & ~x289 & ~x291 & ~x301 & ~x304 & ~x306 & ~x316 & ~x317 & ~x332 & ~x337 & ~x360 & ~x389 & ~x396 & ~x397 & ~x428 & ~x446 & ~x453 & ~x472 & ~x474 & ~x480 & ~x481 & ~x498 & ~x533 & ~x648 & ~x670 & ~x672 & ~x692 & ~x725 & ~x727 & ~x728 & ~x737 & ~x756 & ~x766 & ~x777 & ~x780 & ~x783;
assign c599 =  x152 &  x153 &  x154 & ~x1 & ~x5 & ~x12 & ~x13 & ~x15 & ~x22 & ~x23 & ~x24 & ~x25 & ~x27 & ~x29 & ~x30 & ~x50 & ~x54 & ~x55 & ~x59 & ~x60 & ~x62 & ~x64 & ~x69 & ~x70 & ~x72 & ~x74 & ~x75 & ~x78 & ~x79 & ~x87 & ~x88 & ~x104 & ~x105 & ~x109 & ~x112 & ~x115 & ~x116 & ~x133 & ~x135 & ~x143 & ~x163 & ~x166 & ~x170 & ~x193 & ~x196 & ~x221 & ~x236 & ~x250 & ~x253 & ~x254 & ~x256 & ~x262 & ~x263 & ~x275 & ~x280 & ~x282 & ~x289 & ~x303 & ~x307 & ~x311 & ~x314 & ~x332 & ~x333 & ~x360 & ~x365 & ~x366 & ~x369 & ~x394 & ~x419 & ~x423 & ~x475 & ~x476 & ~x506 & ~x532 & ~x561 & ~x585 & ~x615 & ~x643 & ~x670 & ~x673 & ~x697 & ~x703 & ~x709 & ~x715 & ~x716 & ~x720 & ~x724 & ~x725 & ~x726 & ~x727 & ~x730 & ~x731 & ~x733 & ~x735 & ~x736 & ~x738 & ~x740 & ~x742 & ~x743 & ~x748 & ~x750 & ~x761 & ~x764 & ~x765 & ~x768 & ~x776 & ~x777 & ~x778;
assign c5101 =  x356 & ~x1 & ~x26 & ~x31 & ~x33 & ~x62 & ~x66 & ~x79 & ~x81 & ~x107 & ~x121 & ~x144 & ~x145 & ~x193 & ~x201 & ~x222 & ~x250 & ~x252 & ~x257 & ~x305 & ~x308 & ~x325 & ~x392 & ~x416 & ~x444 & ~x472 & ~x478 & ~x529 & ~x533 & ~x563 & ~x591 & ~x620 & ~x647 & ~x667 & ~x670 & ~x672 & ~x726 & ~x739 & ~x752 & ~x759 & ~x760;
assign c5103 =  x460 &  x516 &  x543 &  x544 & ~x2 & ~x10 & ~x122 & ~x192 & ~x338 & ~x451 & ~x481 & ~x482 & ~x642 & ~x719 & ~x770;
assign c5105 =  x356 &  x384 &  x411 &  x412;
assign c5107 =  x95;
assign c5109 =  x330 & ~x326;
assign c5111 =  x380 & ~x53 & ~x58 & ~x61 & ~x93 & ~x106 & ~x121 & ~x139 & ~x145 & ~x148 & ~x222 & ~x248 & ~x334 & ~x362 & ~x390 & ~x395 & ~x414 & ~x425 & ~x441 & ~x443 & ~x453 & ~x471 & ~x523 & ~x532 & ~x538 & ~x550 & ~x556 & ~x582 & ~x609 & ~x613 & ~x619 & ~x644 & ~x669 & ~x729 & ~x730 & ~x770 & ~x782 & ~x783;
assign c5113 =  x254;
assign c5115 =  x431 &  x486 & ~x31 & ~x39 & ~x43 & ~x52 & ~x57 & ~x73 & ~x82 & ~x85 & ~x113 & ~x116 & ~x137 & ~x141 & ~x228 & ~x369 & ~x370 & ~x373 & ~x399 & ~x427 & ~x474 & ~x477 & ~x481 & ~x619 & ~x644 & ~x648 & ~x674 & ~x695 & ~x704 & ~x728 & ~x737 & ~x739 & ~x743;
assign c5117 =  x270 &  x297 &  x324 & ~x22 & ~x51 & ~x87 & ~x104 & ~x106 & ~x110 & ~x116 & ~x136 & ~x141 & ~x164 & ~x172 & ~x173 & ~x200 & ~x219 & ~x247 & ~x249 & ~x254 & ~x279 & ~x303 & ~x329 & ~x355 & ~x364 & ~x365 & ~x448 & ~x449 & ~x451 & ~x505 & ~x583 & ~x584 & ~x588 & ~x642 & ~x644 & ~x668 & ~x671 & ~x674 & ~x690 & ~x704 & ~x721 & ~x723 & ~x743 & ~x747 & ~x750 & ~x760 & ~x772 & ~x778;
assign c5119 =  x402 &  x456 &  x457 &  x485 &  x513 &  x541 & ~x2 & ~x18 & ~x54 & ~x59 & ~x60 & ~x137 & ~x165 & ~x246 & ~x247 & ~x274 & ~x275 & ~x280 & ~x364 & ~x367 & ~x395 & ~x505 & ~x508 & ~x613 & ~x615 & ~x646 & ~x708 & ~x711 & ~x714 & ~x739 & ~x753 & ~x757 & ~x761 & ~x768 & ~x771;
assign c5121 = ~x5 & ~x6 & ~x25 & ~x26 & ~x68 & ~x71 & ~x77 & ~x79 & ~x81 & ~x83 & ~x91 & ~x98 & ~x100 & ~x107 & ~x113 & ~x127 & ~x133 & ~x150 & ~x160 & ~x192 & ~x199 & ~x218 & ~x219 & ~x225 & ~x251 & ~x253 & ~x275 & ~x303 & ~x369 & ~x390 & ~x402 & ~x456 & ~x477 & ~x483 & ~x505 & ~x508 & ~x511 & ~x537 & ~x539 & ~x556 & ~x584 & ~x620 & ~x623 & ~x710 & ~x711 & ~x727 & ~x729 & ~x731 & ~x736 & ~x769 & ~x777 & ~x782;
assign c5123 =  x353 & ~x1 & ~x6 & ~x29 & ~x32 & ~x34 & ~x35 & ~x37 & ~x39 & ~x46 & ~x47 & ~x52 & ~x57 & ~x58 & ~x63 & ~x73 & ~x78 & ~x80 & ~x84 & ~x96 & ~x107 & ~x108 & ~x110 & ~x113 & ~x115 & ~x120 & ~x124 & ~x140 & ~x142 & ~x144 & ~x150 & ~x167 & ~x195 & ~x198 & ~x225 & ~x250 & ~x307 & ~x310 & ~x322 & ~x332 & ~x333 & ~x338 & ~x367 & ~x384 & ~x388 & ~x412 & ~x416 & ~x446 & ~x473 & ~x530 & ~x531 & ~x562 & ~x589 & ~x639 & ~x675 & ~x698 & ~x699 & ~x700 & ~x702 & ~x724 & ~x728 & ~x733 & ~x735 & ~x742 & ~x761 & ~x770 & ~x772 & ~x774 & ~x779 & ~x783;
assign c5125 =  x426 &  x498;
assign c5127 =  x246 &  x358;
assign c5129 =  x297 & ~x5 & ~x7 & ~x8 & ~x11 & ~x14 & ~x19 & ~x25 & ~x28 & ~x33 & ~x34 & ~x46 & ~x52 & ~x53 & ~x63 & ~x64 & ~x66 & ~x67 & ~x76 & ~x79 & ~x82 & ~x83 & ~x86 & ~x88 & ~x94 & ~x95 & ~x104 & ~x108 & ~x138 & ~x139 & ~x143 & ~x164 & ~x166 & ~x168 & ~x198 & ~x200 & ~x248 & ~x249 & ~x255 & ~x274 & ~x275 & ~x276 & ~x279 & ~x280 & ~x293 & ~x301 & ~x303 & ~x304 & ~x305 & ~x307 & ~x309 & ~x310 & ~x330 & ~x335 & ~x339 & ~x366 & ~x369 & ~x385 & ~x390 & ~x395 & ~x398 & ~x425 & ~x448 & ~x452 & ~x477 & ~x500 & ~x506 & ~x507 & ~x530 & ~x557 & ~x585 & ~x613 & ~x639 & ~x646 & ~x665 & ~x668 & ~x674 & ~x693 & ~x694 & ~x697 & ~x699 & ~x725 & ~x728 & ~x733 & ~x734 & ~x744 & ~x750 & ~x751 & ~x754 & ~x760 & ~x764 & ~x777;
assign c5131 =  x299 &  x325 &  x326 &  x352 &  x379 & ~x2 & ~x4 & ~x5 & ~x8 & ~x16 & ~x21 & ~x23 & ~x25 & ~x26 & ~x27 & ~x28 & ~x31 & ~x33 & ~x37 & ~x44 & ~x47 & ~x51 & ~x52 & ~x56 & ~x60 & ~x64 & ~x65 & ~x87 & ~x88 & ~x95 & ~x106 & ~x118 & ~x139 & ~x165 & ~x170 & ~x171 & ~x197 & ~x198 & ~x199 & ~x222 & ~x224 & ~x249 & ~x253 & ~x254 & ~x275 & ~x277 & ~x280 & ~x304 & ~x305 & ~x310 & ~x331 & ~x332 & ~x334 & ~x360 & ~x362 & ~x363 & ~x367 & ~x389 & ~x390 & ~x394 & ~x417 & ~x419 & ~x422 & ~x446 & ~x449 & ~x475 & ~x476 & ~x503 & ~x505 & ~x530 & ~x531 & ~x613 & ~x640 & ~x643 & ~x673 & ~x675 & ~x694 & ~x697 & ~x699 & ~x702 & ~x704 & ~x713 & ~x715 & ~x716 & ~x724 & ~x728 & ~x732 & ~x734 & ~x738 & ~x743 & ~x748 & ~x750 & ~x753 & ~x754 & ~x755 & ~x756 & ~x757 & ~x758 & ~x759 & ~x761 & ~x773 & ~x778;
assign c5133 =  x493 & ~x10 & ~x31 & ~x48 & ~x71 & ~x84 & ~x122 & ~x151 & ~x153 & ~x161 & ~x162 & ~x198 & ~x200 & ~x246 & ~x247 & ~x275 & ~x335 & ~x420 & ~x501 & ~x511 & ~x567 & ~x625 & ~x644 & ~x670 & ~x702 & ~x727 & ~x733 & ~x760 & ~x776;
assign c5135 = ~x6 & ~x8 & ~x19 & ~x25 & ~x26 & ~x36 & ~x39 & ~x47 & ~x54 & ~x75 & ~x77 & ~x78 & ~x85 & ~x90 & ~x103 & ~x131 & ~x140 & ~x167 & ~x168 & ~x170 & ~x173 & ~x191 & ~x193 & ~x249 & ~x274 & ~x294 & ~x303 & ~x321 & ~x331 & ~x332 & ~x334 & ~x359 & ~x360 & ~x367 & ~x391 & ~x394 & ~x395 & ~x397 & ~x416 & ~x447 & ~x450 & ~x475 & ~x502 & ~x530 & ~x557 & ~x560 & ~x561 & ~x618 & ~x632 & ~x633 & ~x643 & ~x666 & ~x669 & ~x672 & ~x693 & ~x694 & ~x695 & ~x698 & ~x725 & ~x727 & ~x730 & ~x739 & ~x741 & ~x744 & ~x746 & ~x764 & ~x769;
assign c5137 =  x352 &  x435 & ~x568 & ~x626 & ~x756;
assign c5139 =  x388;
assign c5141 =  x272 &  x300 &  x327 & ~x3 & ~x4 & ~x19 & ~x25 & ~x51 & ~x52 & ~x53 & ~x64 & ~x65 & ~x79 & ~x81 & ~x86 & ~x87 & ~x92 & ~x102 & ~x105 & ~x138 & ~x142 & ~x146 & ~x166 & ~x170 & ~x172 & ~x193 & ~x194 & ~x224 & ~x249 & ~x255 & ~x303 & ~x305 & ~x331 & ~x334 & ~x365 & ~x367 & ~x419 & ~x475 & ~x477 & ~x533 & ~x557 & ~x669 & ~x674 & ~x701 & ~x714 & ~x715 & ~x724;
assign c5143 =  x455 & ~x11 & ~x20 & ~x33 & ~x50 & ~x57 & ~x66 & ~x92 & ~x114 & ~x164 & ~x193 & ~x194 & ~x352 & ~x378 & ~x379 & ~x590 & ~x613 & ~x614 & ~x619 & ~x638 & ~x644 & ~x673 & ~x686 & ~x689 & ~x692 & ~x693 & ~x699 & ~x702 & ~x708 & ~x710 & ~x734 & ~x735 & ~x740 & ~x751 & ~x758 & ~x759 & ~x763 & ~x777;
assign c5145 = ~x1 & ~x2 & ~x3 & ~x9 & ~x22 & ~x33 & ~x37 & ~x45 & ~x46 & ~x49 & ~x54 & ~x59 & ~x65 & ~x89 & ~x91 & ~x96 & ~x105 & ~x108 & ~x110 & ~x114 & ~x128 & ~x134 & ~x160 & ~x161 & ~x163 & ~x164 & ~x165 & ~x189 & ~x194 & ~x219 & ~x220 & ~x222 & ~x223 & ~x262 & ~x263 & ~x272 & ~x273 & ~x289 & ~x301 & ~x309 & ~x311 & ~x330 & ~x336 & ~x361 & ~x388 & ~x395 & ~x453 & ~x477 & ~x502 & ~x528 & ~x530 & ~x561 & ~x563 & ~x589 & ~x591 & ~x612 & ~x615 & ~x616 & ~x638 & ~x645 & ~x705 & ~x706 & ~x718 & ~x720 & ~x723 & ~x726 & ~x735 & ~x737 & ~x744 & ~x756 & ~x767 & ~x768 & ~x769 & ~x774;
assign c5147 =  x432 &  x514 & ~x61 & ~x225 & ~x374 & ~x588 & ~x639;
assign c5149 =  x384 & ~x324 & ~x351 & ~x378;
assign c5151 = ~x0 & ~x6 & ~x9 & ~x15 & ~x16 & ~x19 & ~x32 & ~x43 & ~x44 & ~x45 & ~x68 & ~x86 & ~x101 & ~x106 & ~x112 & ~x140 & ~x141 & ~x142 & ~x160 & ~x163 & ~x190 & ~x193 & ~x196 & ~x198 & ~x199 & ~x200 & ~x201 & ~x224 & ~x228 & ~x248 & ~x250 & ~x252 & ~x253 & ~x275 & ~x279 & ~x300 & ~x301 & ~x306 & ~x310 & ~x330 & ~x331 & ~x333 & ~x338 & ~x340 & ~x342 & ~x356 & ~x367 & ~x368 & ~x369 & ~x389 & ~x414 & ~x419 & ~x424 & ~x439 & ~x441 & ~x442 & ~x452 & ~x453 & ~x475 & ~x496 & ~x497 & ~x510 & ~x524 & ~x525 & ~x528 & ~x532 & ~x533 & ~x535 & ~x552 & ~x565 & ~x567 & ~x584 & ~x593 & ~x597 & ~x608 & ~x613 & ~x621 & ~x648 & ~x653 & ~x669 & ~x678 & ~x694 & ~x707 & ~x724 & ~x730 & ~x732 & ~x737 & ~x750 & ~x751 & ~x753 & ~x761 & ~x767 & ~x768 & ~x774 & ~x776 & ~x781 & ~x782;
assign c5153 =  x330 & ~x326;
assign c5155 = ~x34 & ~x52 & ~x57 & ~x113 & ~x115 & ~x129 & ~x138 & ~x145 & ~x187 & ~x248 & ~x276 & ~x303 & ~x397 & ~x482 & ~x509 & ~x534 & ~x567 & ~x585 & ~x587 & ~x591 & ~x618 & ~x625 & ~x638 & ~x646 & ~x654 & ~x702 & ~x709 & ~x778;
assign c5157 =  x354 & ~x58 & ~x61 & ~x569 & ~x620 & ~x650 & ~x699 & ~x703 & ~x749 & ~x777;
assign c5159 =  x551 & ~x237 & ~x249 & ~x279 & ~x290 & ~x291 & ~x317 & ~x588 & ~x698;
assign c5161 =  x302 &  x330;
assign c5163 =  x429 &  x457 &  x484 &  x512 & ~x3 & ~x16 & ~x22 & ~x43 & ~x49 & ~x114 & ~x175 & ~x195 & ~x221 & ~x232 & ~x233 & ~x246 & ~x253 & ~x258 & ~x286 & ~x287 & ~x336 & ~x451 & ~x614 & ~x619 & ~x635 & ~x650 & ~x667 & ~x678 & ~x688 & ~x689 & ~x694 & ~x698 & ~x703 & ~x711 & ~x718 & ~x730 & ~x733 & ~x761 & ~x779;
assign c5165 =  x429 &  x484 &  x599 & ~x7 & ~x8 & ~x10 & ~x14 & ~x16 & ~x20 & ~x25 & ~x27 & ~x34 & ~x39 & ~x46 & ~x48 & ~x50 & ~x57 & ~x59 & ~x61 & ~x62 & ~x63 & ~x81 & ~x86 & ~x88 & ~x89 & ~x94 & ~x96 & ~x138 & ~x140 & ~x141 & ~x147 & ~x165 & ~x171 & ~x191 & ~x254 & ~x255 & ~x276 & ~x277 & ~x282 & ~x308 & ~x310 & ~x334 & ~x335 & ~x340 & ~x365 & ~x392 & ~x396 & ~x417 & ~x418 & ~x420 & ~x445 & ~x450 & ~x475 & ~x501 & ~x503 & ~x532 & ~x559 & ~x584 & ~x585 & ~x588 & ~x589 & ~x591 & ~x611 & ~x613 & ~x614 & ~x616 & ~x617 & ~x619 & ~x641 & ~x643 & ~x645 & ~x675 & ~x678 & ~x681 & ~x693 & ~x694 & ~x703 & ~x705 & ~x711 & ~x713 & ~x719 & ~x721 & ~x730 & ~x735 & ~x736 & ~x737 & ~x738 & ~x740 & ~x746 & ~x764 & ~x771 & ~x773 & ~x780 & ~x783;
assign c5167 =  x213 &  x241 &  x268 & ~x59 & ~x103 & ~x108 & ~x110 & ~x190 & ~x218 & ~x237 & ~x245 & ~x246 & ~x249 & ~x263 & ~x331 & ~x336 & ~x502 & ~x588 & ~x673 & ~x701 & ~x707 & ~x711 & ~x716 & ~x767;
assign c5169 = ~x2 & ~x3 & ~x4 & ~x6 & ~x14 & ~x26 & ~x27 & ~x31 & ~x40 & ~x43 & ~x44 & ~x46 & ~x48 & ~x49 & ~x57 & ~x58 & ~x60 & ~x77 & ~x79 & ~x85 & ~x88 & ~x99 & ~x103 & ~x109 & ~x110 & ~x112 & ~x114 & ~x115 & ~x116 & ~x122 & ~x130 & ~x136 & ~x140 & ~x143 & ~x148 & ~x158 & ~x160 & ~x161 & ~x162 & ~x164 & ~x166 & ~x173 & ~x191 & ~x217 & ~x218 & ~x220 & ~x222 & ~x253 & ~x277 & ~x301 & ~x302 & ~x305 & ~x307 & ~x333 & ~x335 & ~x337 & ~x360 & ~x361 & ~x363 & ~x386 & ~x390 & ~x391 & ~x394 & ~x396 & ~x418 & ~x422 & ~x447 & ~x477 & ~x478 & ~x479 & ~x482 & ~x499 & ~x500 & ~x503 & ~x511 & ~x512 & ~x525 & ~x538 & ~x540 & ~x556 & ~x557 & ~x562 & ~x567 & ~x568 & ~x581 & ~x587 & ~x590 & ~x594 & ~x595 & ~x597 & ~x598 & ~x608 & ~x610 & ~x614 & ~x615 & ~x620 & ~x623 & ~x626 & ~x638 & ~x640 & ~x648 & ~x651 & ~x652 & ~x671 & ~x677 & ~x678 & ~x693 & ~x701 & ~x720 & ~x724 & ~x731 & ~x732 & ~x735 & ~x736 & ~x748 & ~x751 & ~x753 & ~x754 & ~x757 & ~x762;
assign c5171 =  x269 &  x297 &  x381 & ~x10 & ~x20 & ~x44 & ~x50 & ~x70 & ~x77 & ~x78 & ~x84 & ~x86 & ~x87 & ~x107 & ~x108 & ~x116 & ~x132 & ~x133 & ~x136 & ~x164 & ~x190 & ~x246 & ~x274 & ~x300 & ~x329 & ~x332 & ~x336 & ~x359 & ~x362 & ~x389 & ~x417 & ~x423 & ~x444 & ~x475 & ~x529 & ~x614 & ~x674 & ~x708 & ~x725 & ~x726 & ~x728 & ~x729 & ~x734 & ~x779;
assign c5173 = ~x1 & ~x5 & ~x17 & ~x23 & ~x26 & ~x30 & ~x36 & ~x39 & ~x48 & ~x55 & ~x62 & ~x65 & ~x77 & ~x85 & ~x86 & ~x90 & ~x102 & ~x105 & ~x107 & ~x108 & ~x142 & ~x148 & ~x161 & ~x167 & ~x185 & ~x189 & ~x197 & ~x216 & ~x242 & ~x247 & ~x272 & ~x275 & ~x277 & ~x303 & ~x308 & ~x331 & ~x334 & ~x365 & ~x418 & ~x422 & ~x449 & ~x450 & ~x477 & ~x479 & ~x563 & ~x566 & ~x568 & ~x596 & ~x611 & ~x613 & ~x626 & ~x658 & ~x680 & ~x692 & ~x706 & ~x714 & ~x715 & ~x752 & ~x758 & ~x774 & ~x776 & ~x779;
assign c5175 =  x200;
assign c5177 =  x242 &  x623 & ~x164 & ~x249 & ~x263 & ~x265 & ~x317;
assign c5179 =  x381 &  x408 &  x462 & ~x16 & ~x21 & ~x22 & ~x29 & ~x56 & ~x61 & ~x71 & ~x86 & ~x104 & ~x107 & ~x108 & ~x227 & ~x309 & ~x367 & ~x474 & ~x537 & ~x588 & ~x640 & ~x712 & ~x722 & ~x752 & ~x756 & ~x767;
assign c5181 =  x384 & ~x324 & ~x326 & ~x351 & ~x620;
assign c5183 =  x268 &  x295 &  x350 & ~x15 & ~x29 & ~x39 & ~x61 & ~x62 & ~x64 & ~x79 & ~x81 & ~x114 & ~x135 & ~x139 & ~x142 & ~x190 & ~x192 & ~x197 & ~x221 & ~x245 & ~x246 & ~x247 & ~x274 & ~x288 & ~x301 & ~x305 & ~x316 & ~x317 & ~x335 & ~x336 & ~x344 & ~x358 & ~x361 & ~x369 & ~x372 & ~x389 & ~x426 & ~x474 & ~x477 & ~x504 & ~x508 & ~x558 & ~x610 & ~x639 & ~x645 & ~x670 & ~x710 & ~x719 & ~x720 & ~x722 & ~x728 & ~x732 & ~x773;
assign c5185 = ~x0 & ~x130 & ~x277 & ~x347 & ~x477 & ~x510 & ~x564 & ~x627;
assign c5187 = ~x35 & ~x116 & ~x162 & ~x195 & ~x245 & ~x263 & ~x281 & ~x290 & ~x301 & ~x304 & ~x317 & ~x334 & ~x363 & ~x392 & ~x397 & ~x425 & ~x511 & ~x535 & ~x548 & ~x583 & ~x584 & ~x770 & ~x771;
assign c5189 =  x294 & ~x1 & ~x3 & ~x16 & ~x21 & ~x25 & ~x28 & ~x37 & ~x43 & ~x48 & ~x49 & ~x66 & ~x67 & ~x69 & ~x78 & ~x104 & ~x110 & ~x119 & ~x120 & ~x136 & ~x158 & ~x159 & ~x187 & ~x190 & ~x194 & ~x215 & ~x225 & ~x245 & ~x249 & ~x270 & ~x272 & ~x275 & ~x302 & ~x303 & ~x305 & ~x334 & ~x338 & ~x357 & ~x358 & ~x392 & ~x448 & ~x449 & ~x451 & ~x452 & ~x454 & ~x481 & ~x506 & ~x507 & ~x510 & ~x530 & ~x568 & ~x588 & ~x614 & ~x624 & ~x644 & ~x650 & ~x652 & ~x673 & ~x695 & ~x697 & ~x698 & ~x726 & ~x731 & ~x737 & ~x741 & ~x753 & ~x756 & ~x769 & ~x775 & ~x776 & ~x783;
assign c5191 =  x120;
assign c5193 =  x228;
assign c5195 =  x486 &  x513 & ~x21 & ~x28 & ~x48 & ~x51 & ~x121 & ~x137 & ~x163 & ~x248 & ~x255 & ~x283 & ~x285 & ~x286 & ~x304 & ~x362 & ~x398 & ~x419 & ~x453 & ~x503 & ~x508 & ~x589 & ~x591 & ~x636 & ~x642 & ~x645 & ~x676 & ~x686 & ~x689 & ~x712 & ~x717 & ~x721 & ~x740 & ~x777;
assign c5197 =  x175 & ~x372;
assign c5199 =  x382 &  x409 & ~x62 & ~x179 & ~x351 & ~x365 & ~x395 & ~x496 & ~x538 & ~x592 & ~x670;
assign c5201 =  x465 & ~x83 & ~x104 & ~x118 & ~x119 & ~x133 & ~x146 & ~x162 & ~x277 & ~x375 & ~x390 & ~x451 & ~x544 & ~x580 & ~x586 & ~x731 & ~x759;
assign c5203 =  x359;
assign c5205 =  x351 &  x379 &  x433 & ~x0 & ~x91 & ~x112 & ~x131 & ~x303 & ~x320 & ~x422 & ~x475 & ~x586 & ~x590 & ~x674 & ~x702 & ~x755;
assign c5207 =  x274 & ~x430;
assign c5209 =  x355 &  x383 &  x410 & ~x172 & ~x448 & ~x499 & ~x538 & ~x568;
assign c5211 =  x440 & ~x354 & ~x381 & ~x635;
assign c5213 = ~x45 & ~x76 & ~x108 & ~x168 & ~x188 & ~x192 & ~x275 & ~x291 & ~x317 & ~x369 & ~x392 & ~x414 & ~x428 & ~x456 & ~x473 & ~x478 & ~x567 & ~x611 & ~x695;
assign c5215 =  x414 & ~x324 & ~x378;
assign c5217 =  x355 & ~x8 & ~x11 & ~x23 & ~x26 & ~x29 & ~x34 & ~x53 & ~x54 & ~x62 & ~x71 & ~x79 & ~x83 & ~x91 & ~x96 & ~x108 & ~x120 & ~x137 & ~x142 & ~x253 & ~x279 & ~x281 & ~x304 & ~x331 & ~x337 & ~x358 & ~x360 & ~x367 & ~x386 & ~x389 & ~x413 & ~x415 & ~x420 & ~x443 & ~x450 & ~x469 & ~x498 & ~x504 & ~x509 & ~x510 & ~x586 & ~x616 & ~x646 & ~x647 & ~x668 & ~x703 & ~x725;
assign c5219 =  x95;
assign c5221 = ~x1 & ~x4 & ~x7 & ~x9 & ~x17 & ~x24 & ~x25 & ~x30 & ~x31 & ~x33 & ~x34 & ~x37 & ~x38 & ~x39 & ~x57 & ~x60 & ~x61 & ~x63 & ~x72 & ~x93 & ~x115 & ~x138 & ~x140 & ~x141 & ~x142 & ~x168 & ~x169 & ~x173 & ~x174 & ~x195 & ~x197 & ~x219 & ~x220 & ~x221 & ~x223 & ~x228 & ~x236 & ~x237 & ~x246 & ~x251 & ~x258 & ~x260 & ~x263 & ~x264 & ~x273 & ~x276 & ~x283 & ~x287 & ~x289 & ~x290 & ~x301 & ~x302 & ~x303 & ~x306 & ~x309 & ~x330 & ~x331 & ~x332 & ~x336 & ~x340 & ~x362 & ~x369 & ~x387 & ~x388 & ~x393 & ~x394 & ~x418 & ~x419 & ~x424 & ~x427 & ~x443 & ~x453 & ~x454 & ~x476 & ~x504 & ~x535 & ~x562 & ~x587 & ~x591 & ~x641 & ~x646 & ~x673 & ~x694 & ~x695 & ~x706 & ~x711 & ~x715 & ~x730 & ~x746 & ~x750 & ~x751 & ~x752 & ~x780;
assign c5223 =  x285 &  x550 & ~x628;
assign c5225 =  x383 & ~x45 & ~x132 & ~x159 & ~x179 & ~x206 & ~x215 & ~x363 & ~x444 & ~x451 & ~x480 & ~x501 & ~x504 & ~x554 & ~x594 & ~x614 & ~x618 & ~x651 & ~x671;
assign c5227 =  x295 &  x378 & ~x37 & ~x54 & ~x57 & ~x89 & ~x92 & ~x93 & ~x99 & ~x104 & ~x108 & ~x109 & ~x194 & ~x222 & ~x228 & ~x249 & ~x335 & ~x355 & ~x359 & ~x364 & ~x419 & ~x471 & ~x473 & ~x476 & ~x481 & ~x505 & ~x510 & ~x556 & ~x558 & ~x559 & ~x560 & ~x645 & ~x704 & ~x716 & ~x721 & ~x722 & ~x778;
assign c5229 =  x300 &  x327 &  x355 & ~x1 & ~x3 & ~x4 & ~x6 & ~x8 & ~x10 & ~x12 & ~x18 & ~x21 & ~x22 & ~x23 & ~x29 & ~x30 & ~x34 & ~x35 & ~x36 & ~x38 & ~x42 & ~x43 & ~x44 & ~x45 & ~x48 & ~x49 & ~x50 & ~x51 & ~x52 & ~x54 & ~x59 & ~x62 & ~x64 & ~x65 & ~x70 & ~x71 & ~x72 & ~x76 & ~x77 & ~x78 & ~x79 & ~x80 & ~x85 & ~x86 & ~x87 & ~x88 & ~x89 & ~x92 & ~x95 & ~x96 & ~x99 & ~x103 & ~x106 & ~x107 & ~x109 & ~x110 & ~x112 & ~x115 & ~x117 & ~x120 & ~x138 & ~x139 & ~x140 & ~x141 & ~x142 & ~x143 & ~x144 & ~x145 & ~x147 & ~x167 & ~x168 & ~x169 & ~x170 & ~x171 & ~x172 & ~x173 & ~x174 & ~x194 & ~x196 & ~x198 & ~x200 & ~x224 & ~x225 & ~x226 & ~x251 & ~x252 & ~x254 & ~x256 & ~x283 & ~x306 & ~x307 & ~x332 & ~x358 & ~x360 & ~x361 & ~x363 & ~x364 & ~x366 & ~x386 & ~x388 & ~x389 & ~x390 & ~x392 & ~x393 & ~x394 & ~x417 & ~x420 & ~x421 & ~x444 & ~x445 & ~x447 & ~x448 & ~x449 & ~x451 & ~x473 & ~x474 & ~x477 & ~x501 & ~x502 & ~x504 & ~x528 & ~x529 & ~x531 & ~x532 & ~x533 & ~x534 & ~x556 & ~x557 & ~x558 & ~x559 & ~x560 & ~x561 & ~x585 & ~x586 & ~x588 & ~x589 & ~x614 & ~x616 & ~x617 & ~x618 & ~x640 & ~x641 & ~x644 & ~x645 & ~x646 & ~x668 & ~x671 & ~x673 & ~x674 & ~x675 & ~x679 & ~x695 & ~x696 & ~x698 & ~x699 & ~x700 & ~x704 & ~x705 & ~x706 & ~x722 & ~x724 & ~x726 & ~x727 & ~x728 & ~x729 & ~x730 & ~x732 & ~x733 & ~x734 & ~x748 & ~x749 & ~x750 & ~x751 & ~x752 & ~x754 & ~x755 & ~x757 & ~x759 & ~x760 & ~x761 & ~x763 & ~x764 & ~x765 & ~x767 & ~x769 & ~x771 & ~x777 & ~x778 & ~x781 & ~x783;
assign c5231 =  x184 &  x241 &  x269 &  x296 & ~x12 & ~x20 & ~x47 & ~x57 & ~x64 & ~x67 & ~x101 & ~x102 & ~x106 & ~x136 & ~x140 & ~x145 & ~x170 & ~x218 & ~x272 & ~x275 & ~x338 & ~x358 & ~x359 & ~x450 & ~x476 & ~x537 & ~x672 & ~x699 & ~x702 & ~x704 & ~x739 & ~x740 & ~x753 & ~x761 & ~x763 & ~x764;
assign c5233 =  x431 &  x433 &  x459 &  x485 &  x486 &  x513 & ~x27 & ~x42 & ~x44 & ~x51 & ~x84 & ~x337 & ~x341 & ~x478 & ~x506 & ~x558 & ~x590 & ~x613 & ~x641 & ~x663 & ~x668 & ~x672 & ~x735 & ~x765 & ~x767;
assign c5235 =  x97;
assign c5237 =  x325 & ~x1 & ~x3 & ~x19 & ~x34 & ~x54 & ~x63 & ~x74 & ~x80 & ~x83 & ~x104 & ~x111 & ~x130 & ~x132 & ~x138 & ~x221 & ~x248 & ~x249 & ~x250 & ~x252 & ~x277 & ~x303 & ~x304 & ~x328 & ~x330 & ~x332 & ~x335 & ~x356 & ~x361 & ~x364 & ~x383 & ~x416 & ~x423 & ~x426 & ~x446 & ~x505 & ~x558 & ~x586 & ~x588 & ~x612 & ~x613 & ~x645 & ~x691 & ~x719 & ~x722 & ~x726 & ~x727 & ~x736 & ~x737 & ~x747 & ~x752 & ~x755 & ~x764;
assign c5239 =  x458 &  x486 & ~x37 & ~x203 & ~x213 & ~x242 & ~x276 & ~x503 & ~x641 & ~x658;
assign c5241 =  x187 &  x273 & ~x4 & ~x25 & ~x51 & ~x67 & ~x112 & ~x420 & ~x445 & ~x689 & ~x749;
assign c5243 =  x469 & ~x5 & ~x14 & ~x26 & ~x51 & ~x53 & ~x57 & ~x81 & ~x85 & ~x167 & ~x197 & ~x221 & ~x226 & ~x232 & ~x233 & ~x234 & ~x260 & ~x279 & ~x283 & ~x288 & ~x313 & ~x327 & ~x362 & ~x446 & ~x536 & ~x586 & ~x588 & ~x590 & ~x592 & ~x639 & ~x671 & ~x697 & ~x718 & ~x723 & ~x726 & ~x729;
assign c5245 =  x231 & ~x345;
assign c5247 =  x325 & ~x4 & ~x16 & ~x28 & ~x31 & ~x53 & ~x54 & ~x65 & ~x69 & ~x73 & ~x78 & ~x79 & ~x84 & ~x87 & ~x94 & ~x100 & ~x101 & ~x102 & ~x108 & ~x130 & ~x137 & ~x171 & ~x197 & ~x222 & ~x226 & ~x251 & ~x278 & ~x279 & ~x322 & ~x364 & ~x367 & ~x389 & ~x391 & ~x393 & ~x447 & ~x451 & ~x475 & ~x476 & ~x478 & ~x508 & ~x531 & ~x535 & ~x562 & ~x565 & ~x590 & ~x619 & ~x648 & ~x672 & ~x674 & ~x696 & ~x706 & ~x724 & ~x725 & ~x726 & ~x727 & ~x731 & ~x732 & ~x754 & ~x766 & ~x780 & ~x782;
assign c5249 =  x272 &  x329 & ~x174 & ~x304 & ~x749;
assign c5251 =  x705;
assign c5253 =  x463 & ~x63 & ~x255 & ~x629 & ~x640;
assign c5255 =  x270 &  x325 & ~x4 & ~x11 & ~x38 & ~x41 & ~x145 & ~x276 & ~x330 & ~x336 & ~x360 & ~x370 & ~x371 & ~x427 & ~x544 & ~x697 & ~x723 & ~x724 & ~x749;
assign c5257 =  x380 & ~x3 & ~x4 & ~x35 & ~x39 & ~x52 & ~x53 & ~x64 & ~x65 & ~x72 & ~x75 & ~x92 & ~x107 & ~x109 & ~x112 & ~x113 & ~x128 & ~x134 & ~x139 & ~x141 & ~x145 & ~x160 & ~x162 & ~x165 & ~x188 & ~x197 & ~x219 & ~x223 & ~x227 & ~x248 & ~x256 & ~x275 & ~x314 & ~x336 & ~x360 & ~x361 & ~x362 & ~x363 & ~x365 & ~x390 & ~x448 & ~x451 & ~x453 & ~x454 & ~x455 & ~x475 & ~x504 & ~x505 & ~x527 & ~x529 & ~x561 & ~x582 & ~x589 & ~x609 & ~x613 & ~x615 & ~x672 & ~x695 & ~x736 & ~x743 & ~x761 & ~x765 & ~x775 & ~x778 & ~x780;
assign c5259 =  x326 &  x407 & ~x2 & ~x8 & ~x11 & ~x18 & ~x25 & ~x27 & ~x52 & ~x64 & ~x71 & ~x91 & ~x108 & ~x141 & ~x194 & ~x225 & ~x253 & ~x276 & ~x281 & ~x331 & ~x394 & ~x477 & ~x481 & ~x502 & ~x504 & ~x528 & ~x560 & ~x584 & ~x585 & ~x611 & ~x616 & ~x618 & ~x673 & ~x687 & ~x749 & ~x757 & ~x771 & ~x777;
assign c5261 =  x303 &  x359 &  x415;
assign c5263 =  x458 &  x486 & ~x4 & ~x15 & ~x18 & ~x23 & ~x25 & ~x26 & ~x41 & ~x43 & ~x45 & ~x47 & ~x53 & ~x54 & ~x55 & ~x75 & ~x78 & ~x85 & ~x88 & ~x94 & ~x108 & ~x109 & ~x114 & ~x115 & ~x140 & ~x144 & ~x178 & ~x196 & ~x220 & ~x223 & ~x224 & ~x229 & ~x231 & ~x241 & ~x256 & ~x259 & ~x275 & ~x286 & ~x287 & ~x313 & ~x331 & ~x332 & ~x342 & ~x360 & ~x362 & ~x389 & ~x447 & ~x482 & ~x504 & ~x509 & ~x529 & ~x534 & ~x585 & ~x611 & ~x645 & ~x648 & ~x677 & ~x689 & ~x702 & ~x705 & ~x716 & ~x718 & ~x722 & ~x723 & ~x729 & ~x733 & ~x747 & ~x761 & ~x763 & ~x768;
assign c5265 =  x406 & ~x33 & ~x99 & ~x100 & ~x189 & ~x218 & ~x220 & ~x247 & ~x339 & ~x402 & ~x474 & ~x624 & ~x676;
assign c5267 =  x199;
assign c5269 =  x299 & ~x3 & ~x7 & ~x8 & ~x14 & ~x26 & ~x35 & ~x46 & ~x56 & ~x58 & ~x67 & ~x69 & ~x81 & ~x96 & ~x108 & ~x112 & ~x113 & ~x115 & ~x119 & ~x143 & ~x168 & ~x221 & ~x222 & ~x224 & ~x225 & ~x248 & ~x255 & ~x276 & ~x280 & ~x294 & ~x308 & ~x313 & ~x334 & ~x338 & ~x357 & ~x361 & ~x388 & ~x392 & ~x394 & ~x396 & ~x419 & ~x477 & ~x505 & ~x587 & ~x589 & ~x613 & ~x640 & ~x646 & ~x706 & ~x708 & ~x716 & ~x719 & ~x722 & ~x732 & ~x739 & ~x742 & ~x743 & ~x744 & ~x747 & ~x748 & ~x754 & ~x755 & ~x764 & ~x767 & ~x772;
assign c5271 =  x243 &  x271 &  x299 & ~x3 & ~x6 & ~x7 & ~x10 & ~x11 & ~x13 & ~x15 & ~x16 & ~x20 & ~x27 & ~x32 & ~x35 & ~x37 & ~x39 & ~x43 & ~x44 & ~x45 & ~x46 & ~x50 & ~x51 & ~x53 & ~x56 & ~x64 & ~x67 & ~x73 & ~x75 & ~x79 & ~x81 & ~x88 & ~x96 & ~x110 & ~x111 & ~x115 & ~x135 & ~x139 & ~x140 & ~x141 & ~x144 & ~x166 & ~x168 & ~x170 & ~x171 & ~x191 & ~x194 & ~x195 & ~x219 & ~x220 & ~x221 & ~x223 & ~x226 & ~x228 & ~x248 & ~x251 & ~x252 & ~x254 & ~x255 & ~x275 & ~x276 & ~x280 & ~x281 & ~x282 & ~x283 & ~x303 & ~x305 & ~x310 & ~x332 & ~x335 & ~x336 & ~x360 & ~x363 & ~x364 & ~x366 & ~x388 & ~x389 & ~x392 & ~x393 & ~x416 & ~x417 & ~x419 & ~x445 & ~x446 & ~x447 & ~x475 & ~x477 & ~x478 & ~x504 & ~x529 & ~x530 & ~x557 & ~x558 & ~x559 & ~x561 & ~x584 & ~x585 & ~x588 & ~x639 & ~x643 & ~x669 & ~x671 & ~x676 & ~x688 & ~x689 & ~x690 & ~x695 & ~x700 & ~x703 & ~x714 & ~x719 & ~x721 & ~x725 & ~x727 & ~x728 & ~x729 & ~x740 & ~x741 & ~x744 & ~x750 & ~x752 & ~x753 & ~x755 & ~x756 & ~x758 & ~x762 & ~x764 & ~x769 & ~x770 & ~x775 & ~x781 & ~x782 & ~x783;
assign c5273 =  x490 & ~x0 & ~x7 & ~x9 & ~x64 & ~x67 & ~x68 & ~x113 & ~x164 & ~x218 & ~x248 & ~x302 & ~x304 & ~x333 & ~x337 & ~x400 & ~x418 & ~x540 & ~x563 & ~x586 & ~x587 & ~x596 & ~x620 & ~x624 & ~x641 & ~x646 & ~x665 & ~x669 & ~x727;
assign c5275 =  x325 &  x408 & ~x7 & ~x16 & ~x63 & ~x85 & ~x104 & ~x112 & ~x141 & ~x172 & ~x201 & ~x223 & ~x251 & ~x304 & ~x305 & ~x308 & ~x332 & ~x337 & ~x385 & ~x420 & ~x530 & ~x543 & ~x585 & ~x694 & ~x696 & ~x774;
assign c5277 =  x329 & ~x47 & ~x332 & ~x348 & ~x531 & ~x557 & ~x612 & ~x617;
assign c5279 =  x270 & ~x6 & ~x7 & ~x8 & ~x9 & ~x11 & ~x15 & ~x17 & ~x22 & ~x23 & ~x57 & ~x66 & ~x68 & ~x70 & ~x71 & ~x86 & ~x104 & ~x105 & ~x106 & ~x107 & ~x109 & ~x117 & ~x118 & ~x132 & ~x133 & ~x134 & ~x135 & ~x140 & ~x142 & ~x145 & ~x166 & ~x174 & ~x222 & ~x224 & ~x229 & ~x247 & ~x251 & ~x255 & ~x267 & ~x293 & ~x305 & ~x308 & ~x363 & ~x388 & ~x446 & ~x477 & ~x502 & ~x504 & ~x531 & ~x532 & ~x559 & ~x560 & ~x588 & ~x589 & ~x613 & ~x614 & ~x618 & ~x643 & ~x644 & ~x645 & ~x646 & ~x670 & ~x673 & ~x677 & ~x700 & ~x703 & ~x726 & ~x728 & ~x729 & ~x733 & ~x748 & ~x749 & ~x756 & ~x757 & ~x759 & ~x762 & ~x763 & ~x765 & ~x779;
assign c5281 =  x359 &  x415 & ~x326;
assign c5283 =  x241 & ~x1 & ~x2 & ~x12 & ~x15 & ~x16 & ~x19 & ~x20 & ~x22 & ~x27 & ~x28 & ~x31 & ~x39 & ~x40 & ~x42 & ~x46 & ~x48 & ~x49 & ~x50 & ~x51 & ~x58 & ~x60 & ~x61 & ~x62 & ~x67 & ~x68 & ~x70 & ~x71 & ~x73 & ~x74 & ~x75 & ~x78 & ~x93 & ~x94 & ~x106 & ~x109 & ~x111 & ~x115 & ~x116 & ~x117 & ~x132 & ~x134 & ~x141 & ~x144 & ~x145 & ~x146 & ~x161 & ~x162 & ~x164 & ~x166 & ~x167 & ~x170 & ~x173 & ~x188 & ~x189 & ~x191 & ~x195 & ~x196 & ~x201 & ~x217 & ~x218 & ~x219 & ~x222 & ~x224 & ~x229 & ~x244 & ~x245 & ~x251 & ~x253 & ~x274 & ~x276 & ~x277 & ~x304 & ~x305 & ~x306 & ~x311 & ~x332 & ~x337 & ~x339 & ~x340 & ~x361 & ~x367 & ~x368 & ~x388 & ~x389 & ~x390 & ~x391 & ~x392 & ~x393 & ~x395 & ~x418 & ~x419 & ~x420 & ~x449 & ~x475 & ~x476 & ~x501 & ~x502 & ~x506 & ~x533 & ~x559 & ~x561 & ~x562 & ~x587 & ~x588 & ~x590 & ~x591 & ~x614 & ~x615 & ~x616 & ~x645 & ~x646 & ~x647 & ~x669 & ~x672 & ~x674 & ~x684 & ~x693 & ~x695 & ~x697 & ~x700 & ~x701 & ~x705 & ~x707 & ~x709 & ~x717 & ~x724 & ~x728 & ~x730 & ~x733 & ~x739 & ~x742 & ~x743 & ~x744 & ~x746 & ~x747 & ~x748 & ~x749 & ~x752 & ~x754 & ~x758 & ~x759 & ~x760 & ~x766 & ~x768 & ~x770 & ~x771 & ~x773 & ~x774 & ~x778 & ~x780 & ~x782;
assign c5285 =  x436 &  x463 & ~x19 & ~x30 & ~x34 & ~x40 & ~x52 & ~x55 & ~x59 & ~x60 & ~x97 & ~x105 & ~x136 & ~x141 & ~x169 & ~x178 & ~x225 & ~x255 & ~x307 & ~x308 & ~x333 & ~x336 & ~x388 & ~x392 & ~x419 & ~x449 & ~x470 & ~x474 & ~x494 & ~x500 & ~x501 & ~x510 & ~x511 & ~x526 & ~x536 & ~x555 & ~x558 & ~x560 & ~x565 & ~x585 & ~x614 & ~x616 & ~x623 & ~x640 & ~x643 & ~x695 & ~x697 & ~x703 & ~x704 & ~x751 & ~x761;
assign c5287 =  x273 &  x301 &  x328 & ~x304 & ~x332 & ~x361 & ~x618;
assign c5289 =  x294 &  x322 &  x378 & ~x85 & ~x98 & ~x137 & ~x160 & ~x218 & ~x274 & ~x275 & ~x280 & ~x299 & ~x302 & ~x339 & ~x389 & ~x391 & ~x418 & ~x423 & ~x427 & ~x445 & ~x446 & ~x450 & ~x482 & ~x483 & ~x512 & ~x559 & ~x561 & ~x612 & ~x642 & ~x650 & ~x670 & ~x703 & ~x725;
assign c5291 =  x382 & ~x158 & ~x186 & ~x225 & ~x248 & ~x280 & ~x421 & ~x473 & ~x481 & ~x527 & ~x538 & ~x540 & ~x553 & ~x558 & ~x565 & ~x591 & ~x614 & ~x616 & ~x625 & ~x653 & ~x755;
assign c5293 =  x399 & ~x17 & ~x349 & ~x376 & ~x403 & ~x431 & ~x754;
assign c5295 = ~x29 & ~x47 & ~x112 & ~x180 & ~x193 & ~x203 & ~x207 & ~x221 & ~x227 & ~x233 & ~x234 & ~x248 & ~x253 & ~x255 & ~x258 & ~x271 & ~x277 & ~x282 & ~x325 & ~x333 & ~x340 & ~x392 & ~x398 & ~x413 & ~x418 & ~x421 & ~x425 & ~x426 & ~x443 & ~x477 & ~x480 & ~x502 & ~x506 & ~x509 & ~x539 & ~x554 & ~x558 & ~x563 & ~x566 & ~x582 & ~x594 & ~x595 & ~x644 & ~x646 & ~x649 & ~x651 & ~x683 & ~x687 & ~x726 & ~x758 & ~x768;
assign c5297 =  x459 &  x487 &  x515 &  x543 & ~x0 & ~x10 & ~x11 & ~x12 & ~x15 & ~x20 & ~x27 & ~x33 & ~x35 & ~x37 & ~x44 & ~x50 & ~x51 & ~x54 & ~x68 & ~x79 & ~x84 & ~x107 & ~x109 & ~x136 & ~x138 & ~x139 & ~x142 & ~x143 & ~x145 & ~x163 & ~x164 & ~x170 & ~x171 & ~x172 & ~x175 & ~x176 & ~x191 & ~x197 & ~x198 & ~x200 & ~x220 & ~x221 & ~x224 & ~x227 & ~x247 & ~x248 & ~x276 & ~x307 & ~x330 & ~x331 & ~x340 & ~x358 & ~x366 & ~x386 & ~x388 & ~x389 & ~x395 & ~x396 & ~x423 & ~x446 & ~x452 & ~x453 & ~x509 & ~x531 & ~x556 & ~x565 & ~x590 & ~x646 & ~x648 & ~x649 & ~x665 & ~x673 & ~x679 & ~x682 & ~x683 & ~x684 & ~x696 & ~x707 & ~x709 & ~x714 & ~x720 & ~x735 & ~x739 & ~x744 & ~x763 & ~x775 & ~x777 & ~x778 & ~x782;
assign c5299 =  x388;
assign c60 =  x546 & ~x48 & ~x50 & ~x59 & ~x108 & ~x129 & ~x137 & ~x141 & ~x210 & ~x230 & ~x246 & ~x255 & ~x257 & ~x314 & ~x333 & ~x362 & ~x367 & ~x398 & ~x418 & ~x424 & ~x447 & ~x455 & ~x474 & ~x479 & ~x511 & ~x530 & ~x561 & ~x661 & ~x667 & ~x685 & ~x686 & ~x703 & ~x721 & ~x724 & ~x782;
assign c62 =  x235 & ~x2 & ~x7 & ~x12 & ~x15 & ~x19 & ~x35 & ~x64 & ~x67 & ~x83 & ~x138 & ~x145 & ~x169 & ~x217 & ~x221 & ~x267 & ~x268 & ~x278 & ~x307 & ~x335 & ~x337 & ~x349 & ~x424 & ~x478 & ~x535 & ~x585 & ~x590 & ~x615 & ~x651 & ~x652 & ~x657 & ~x666 & ~x672 & ~x673 & ~x677 & ~x691 & ~x737 & ~x740 & ~x755 & ~x756 & ~x758 & ~x782;
assign c64 = ~x5 & ~x6 & ~x12 & ~x15 & ~x16 & ~x17 & ~x18 & ~x26 & ~x29 & ~x30 & ~x32 & ~x34 & ~x38 & ~x43 & ~x54 & ~x56 & ~x65 & ~x76 & ~x80 & ~x107 & ~x115 & ~x118 & ~x131 & ~x133 & ~x135 & ~x136 & ~x137 & ~x140 & ~x143 & ~x163 & ~x165 & ~x169 & ~x170 & ~x174 & ~x186 & ~x187 & ~x197 & ~x198 & ~x202 & ~x203 & ~x216 & ~x219 & ~x227 & ~x228 & ~x229 & ~x231 & ~x240 & ~x241 & ~x242 & ~x247 & ~x253 & ~x254 & ~x257 & ~x267 & ~x282 & ~x307 & ~x311 & ~x331 & ~x336 & ~x337 & ~x339 & ~x363 & ~x367 & ~x370 & ~x447 & ~x449 & ~x452 & ~x476 & ~x478 & ~x503 & ~x504 & ~x505 & ~x529 & ~x558 & ~x562 & ~x563 & ~x564 & ~x583 & ~x584 & ~x585 & ~x586 & ~x587 & ~x592 & ~x607 & ~x609 & ~x620 & ~x621 & ~x636 & ~x642 & ~x645 & ~x648 & ~x649 & ~x654 & ~x657 & ~x658 & ~x659 & ~x661 & ~x670 & ~x672 & ~x676 & ~x683 & ~x688 & ~x690 & ~x693 & ~x697 & ~x702 & ~x709 & ~x710 & ~x712 & ~x714 & ~x719 & ~x720 & ~x726 & ~x735 & ~x737 & ~x738 & ~x740 & ~x743 & ~x744 & ~x746 & ~x748 & ~x753 & ~x763 & ~x764 & ~x765 & ~x771 & ~x773 & ~x776;
assign c66 =  x117;
assign c68 =  x428 & ~x2 & ~x4 & ~x17 & ~x18 & ~x38 & ~x43 & ~x50 & ~x51 & ~x60 & ~x62 & ~x63 & ~x73 & ~x75 & ~x80 & ~x90 & ~x115 & ~x139 & ~x141 & ~x142 & ~x146 & ~x166 & ~x168 & ~x193 & ~x197 & ~x214 & ~x225 & ~x248 & ~x256 & ~x279 & ~x281 & ~x282 & ~x294 & ~x304 & ~x308 & ~x334 & ~x337 & ~x341 & ~x355 & ~x360 & ~x389 & ~x390 & ~x394 & ~x422 & ~x425 & ~x448 & ~x454 & ~x481 & ~x502 & ~x505 & ~x509 & ~x561 & ~x565 & ~x566 & ~x588 & ~x591 & ~x593 & ~x612 & ~x617 & ~x621 & ~x640 & ~x643 & ~x671 & ~x682 & ~x686 & ~x688 & ~x690 & ~x699 & ~x701 & ~x702 & ~x712 & ~x715 & ~x720 & ~x726 & ~x738 & ~x742 & ~x744 & ~x755 & ~x762 & ~x766 & ~x775 & ~x779 & ~x783;
assign c610 =  x64;
assign c612 = ~x1 & ~x5 & ~x14 & ~x20 & ~x22 & ~x29 & ~x30 & ~x42 & ~x43 & ~x44 & ~x45 & ~x46 & ~x49 & ~x59 & ~x61 & ~x64 & ~x69 & ~x81 & ~x82 & ~x89 & ~x92 & ~x96 & ~x107 & ~x111 & ~x117 & ~x120 & ~x122 & ~x133 & ~x134 & ~x136 & ~x143 & ~x151 & ~x162 & ~x165 & ~x167 & ~x168 & ~x171 & ~x176 & ~x191 & ~x193 & ~x196 & ~x201 & ~x206 & ~x208 & ~x214 & ~x220 & ~x224 & ~x229 & ~x232 & ~x234 & ~x235 & ~x241 & ~x249 & ~x250 & ~x253 & ~x254 & ~x257 & ~x258 & ~x259 & ~x269 & ~x270 & ~x278 & ~x280 & ~x282 & ~x287 & ~x299 & ~x301 & ~x308 & ~x309 & ~x310 & ~x314 & ~x315 & ~x330 & ~x332 & ~x333 & ~x339 & ~x343 & ~x391 & ~x392 & ~x393 & ~x398 & ~x418 & ~x419 & ~x425 & ~x426 & ~x443 & ~x447 & ~x450 & ~x474 & ~x475 & ~x478 & ~x499 & ~x500 & ~x503 & ~x507 & ~x509 & ~x533 & ~x536 & ~x553 & ~x562 & ~x563 & ~x564 & ~x588 & ~x589 & ~x590 & ~x591 & ~x593 & ~x610 & ~x614 & ~x622 & ~x633 & ~x637 & ~x638 & ~x639 & ~x642 & ~x645 & ~x649 & ~x652 & ~x658 & ~x659 & ~x660 & ~x662 & ~x666 & ~x669 & ~x674 & ~x675 & ~x676 & ~x686 & ~x692 & ~x696 & ~x697 & ~x699 & ~x700 & ~x704 & ~x705 & ~x711 & ~x718 & ~x726 & ~x731 & ~x732 & ~x740 & ~x742 & ~x744 & ~x747 & ~x750 & ~x754 & ~x755 & ~x757 & ~x758 & ~x759 & ~x760 & ~x762 & ~x767 & ~x777 & ~x781;
assign c614 = ~x1 & ~x3 & ~x56 & ~x57 & ~x78 & ~x79 & ~x91 & ~x92 & ~x107 & ~x112 & ~x138 & ~x143 & ~x146 & ~x166 & ~x186 & ~x189 & ~x192 & ~x200 & ~x201 & ~x216 & ~x218 & ~x240 & ~x242 & ~x248 & ~x249 & ~x253 & ~x269 & ~x282 & ~x294 & ~x306 & ~x334 & ~x336 & ~x349 & ~x404 & ~x421 & ~x445 & ~x502 & ~x503 & ~x527 & ~x529 & ~x535 & ~x589 & ~x591 & ~x608 & ~x609 & ~x612 & ~x650 & ~x661 & ~x683 & ~x709 & ~x716 & ~x718 & ~x723 & ~x724 & ~x765 & ~x778;
assign c616 =  x518 &  x520 & ~x42 & ~x127 & ~x182 & ~x191 & ~x198 & ~x209 & ~x219 & ~x227 & ~x246 & ~x264 & ~x291 & ~x298 & ~x365 & ~x478 & ~x619 & ~x672 & ~x727 & ~x767 & ~x772;
assign c618 =  x4;
assign c620 =  x135 &  x161 &  x241 &  x294;
assign c622 =  x373 &  x401 &  x428 &  x456 &  x484 &  x575 &  x601 & ~x10 & ~x23 & ~x25 & ~x28 & ~x48 & ~x49 & ~x61 & ~x84 & ~x87 & ~x116 & ~x133 & ~x134 & ~x140 & ~x162 & ~x163 & ~x172 & ~x188 & ~x189 & ~x216 & ~x219 & ~x221 & ~x242 & ~x247 & ~x256 & ~x277 & ~x306 & ~x313 & ~x332 & ~x337 & ~x361 & ~x362 & ~x363 & ~x364 & ~x366 & ~x367 & ~x396 & ~x425 & ~x452 & ~x474 & ~x504 & ~x506 & ~x507 & ~x532 & ~x559 & ~x561 & ~x562 & ~x586 & ~x593 & ~x613 & ~x619 & ~x622 & ~x623 & ~x639 & ~x641 & ~x645 & ~x651 & ~x653 & ~x654 & ~x655 & ~x656 & ~x659 & ~x666 & ~x683 & ~x687 & ~x693 & ~x705 & ~x706 & ~x707 & ~x714 & ~x728 & ~x731 & ~x737 & ~x748 & ~x750 & ~x755 & ~x767 & ~x779;
assign c624 = ~x2 & ~x3 & ~x5 & ~x6 & ~x7 & ~x11 & ~x12 & ~x18 & ~x19 & ~x20 & ~x22 & ~x23 & ~x24 & ~x25 & ~x26 & ~x27 & ~x30 & ~x31 & ~x32 & ~x33 & ~x36 & ~x40 & ~x41 & ~x43 & ~x45 & ~x46 & ~x48 & ~x50 & ~x51 & ~x52 & ~x53 & ~x54 & ~x56 & ~x57 & ~x58 & ~x59 & ~x62 & ~x73 & ~x76 & ~x80 & ~x81 & ~x82 & ~x83 & ~x85 & ~x86 & ~x87 & ~x89 & ~x106 & ~x112 & ~x115 & ~x131 & ~x133 & ~x134 & ~x135 & ~x137 & ~x139 & ~x140 & ~x141 & ~x142 & ~x143 & ~x145 & ~x147 & ~x158 & ~x159 & ~x160 & ~x161 & ~x162 & ~x163 & ~x164 & ~x165 & ~x166 & ~x170 & ~x171 & ~x186 & ~x187 & ~x188 & ~x189 & ~x190 & ~x191 & ~x193 & ~x194 & ~x196 & ~x198 & ~x199 & ~x214 & ~x215 & ~x216 & ~x218 & ~x219 & ~x223 & ~x224 & ~x225 & ~x226 & ~x229 & ~x240 & ~x241 & ~x242 & ~x247 & ~x249 & ~x250 & ~x251 & ~x252 & ~x253 & ~x267 & ~x268 & ~x277 & ~x278 & ~x280 & ~x281 & ~x283 & ~x294 & ~x306 & ~x309 & ~x311 & ~x335 & ~x339 & ~x362 & ~x364 & ~x365 & ~x366 & ~x367 & ~x390 & ~x392 & ~x393 & ~x395 & ~x396 & ~x417 & ~x419 & ~x420 & ~x421 & ~x422 & ~x424 & ~x446 & ~x447 & ~x448 & ~x449 & ~x452 & ~x474 & ~x477 & ~x502 & ~x504 & ~x505 & ~x508 & ~x531 & ~x534 & ~x536 & ~x555 & ~x558 & ~x559 & ~x560 & ~x561 & ~x562 & ~x564 & ~x565 & ~x583 & ~x584 & ~x585 & ~x589 & ~x590 & ~x591 & ~x594 & ~x595 & ~x609 & ~x610 & ~x611 & ~x615 & ~x617 & ~x618 & ~x621 & ~x624 & ~x637 & ~x638 & ~x639 & ~x641 & ~x644 & ~x648 & ~x649 & ~x650 & ~x651 & ~x653 & ~x656 & ~x664 & ~x665 & ~x666 & ~x667 & ~x669 & ~x670 & ~x671 & ~x672 & ~x673 & ~x675 & ~x677 & ~x679 & ~x680 & ~x684 & ~x685 & ~x686 & ~x688 & ~x689 & ~x690 & ~x694 & ~x698 & ~x706 & ~x707 & ~x711 & ~x713 & ~x714 & ~x715 & ~x716 & ~x718 & ~x719 & ~x720 & ~x721 & ~x722 & ~x724 & ~x725 & ~x730 & ~x734 & ~x735 & ~x736 & ~x741 & ~x743 & ~x745 & ~x746 & ~x747 & ~x748 & ~x749 & ~x750 & ~x751 & ~x755 & ~x757 & ~x759 & ~x766 & ~x767 & ~x768 & ~x771 & ~x772 & ~x773 & ~x775 & ~x777 & ~x779 & ~x780 & ~x782 & ~x783;
assign c626 =  x132 &  x133 &  x186 &  x213 &  x214 &  x240 & ~x127 & ~x128 & ~x153 & ~x154 & ~x207 & ~x233 & ~x234 & ~x298;
assign c628 =  x489 &  x550 &  x571 & ~x95 & ~x97 & ~x150 & ~x206 & ~x207 & ~x234 & ~x300 & ~x636;
assign c630 =  x158 & ~x1 & ~x2 & ~x3 & ~x4 & ~x8 & ~x9 & ~x10 & ~x19 & ~x24 & ~x33 & ~x46 & ~x49 & ~x52 & ~x56 & ~x58 & ~x61 & ~x69 & ~x70 & ~x73 & ~x81 & ~x82 & ~x96 & ~x99 & ~x109 & ~x111 & ~x113 & ~x115 & ~x123 & ~x126 & ~x136 & ~x140 & ~x145 & ~x146 & ~x149 & ~x152 & ~x154 & ~x170 & ~x181 & ~x199 & ~x202 & ~x206 & ~x208 & ~x223 & ~x225 & ~x233 & ~x234 & ~x236 & ~x260 & ~x261 & ~x271 & ~x272 & ~x274 & ~x277 & ~x280 & ~x282 & ~x287 & ~x298 & ~x300 & ~x301 & ~x305 & ~x306 & ~x311 & ~x315 & ~x324 & ~x331 & ~x362 & ~x368 & ~x390 & ~x392 & ~x446 & ~x450 & ~x473 & ~x475 & ~x478 & ~x505 & ~x527 & ~x529 & ~x558 & ~x563 & ~x581 & ~x585 & ~x586 & ~x589 & ~x590 & ~x592 & ~x593 & ~x617 & ~x633 & ~x636 & ~x637 & ~x638 & ~x639 & ~x645 & ~x647 & ~x648 & ~x649 & ~x660 & ~x664 & ~x679 & ~x682 & ~x687 & ~x699 & ~x701 & ~x704 & ~x712 & ~x717 & ~x726 & ~x731 & ~x732 & ~x733 & ~x737 & ~x739 & ~x741 & ~x749 & ~x750 & ~x754 & ~x757 & ~x758;
assign c632 =  x188 &  x295 &  x321 &  x374 &  x375 &  x401 &  x429 &  x599 & ~x151 & ~x206 & ~x300 & ~x301 & ~x330 & ~x332 & ~x739;
assign c634 = ~x40 & ~x54 & ~x161 & ~x170 & ~x188 & ~x191 & ~x192 & ~x215 & ~x219 & ~x242 & ~x269 & ~x294 & ~x295 & ~x320 & ~x348 & ~x393 & ~x636 & ~x638 & ~x642 & ~x653 & ~x655 & ~x691 & ~x756 & ~x776;
assign c636 =  x643;
assign c638 = ~x1 & ~x3 & ~x4 & ~x5 & ~x8 & ~x11 & ~x13 & ~x14 & ~x16 & ~x17 & ~x18 & ~x20 & ~x21 & ~x22 & ~x23 & ~x26 & ~x28 & ~x31 & ~x32 & ~x33 & ~x34 & ~x38 & ~x40 & ~x44 & ~x46 & ~x47 & ~x49 & ~x50 & ~x51 & ~x54 & ~x58 & ~x59 & ~x61 & ~x66 & ~x67 & ~x68 & ~x77 & ~x78 & ~x81 & ~x83 & ~x86 & ~x87 & ~x88 & ~x92 & ~x93 & ~x107 & ~x110 & ~x111 & ~x113 & ~x114 & ~x116 & ~x118 & ~x121 & ~x136 & ~x138 & ~x139 & ~x140 & ~x141 & ~x142 & ~x146 & ~x149 & ~x162 & ~x163 & ~x170 & ~x171 & ~x172 & ~x173 & ~x174 & ~x175 & ~x176 & ~x190 & ~x191 & ~x193 & ~x194 & ~x195 & ~x197 & ~x199 & ~x200 & ~x201 & ~x202 & ~x217 & ~x218 & ~x219 & ~x220 & ~x221 & ~x223 & ~x224 & ~x225 & ~x226 & ~x228 & ~x230 & ~x244 & ~x247 & ~x250 & ~x252 & ~x253 & ~x254 & ~x257 & ~x268 & ~x269 & ~x271 & ~x272 & ~x281 & ~x283 & ~x285 & ~x294 & ~x295 & ~x297 & ~x298 & ~x301 & ~x302 & ~x304 & ~x308 & ~x309 & ~x324 & ~x333 & ~x337 & ~x339 & ~x350 & ~x362 & ~x364 & ~x365 & ~x368 & ~x390 & ~x391 & ~x392 & ~x393 & ~x395 & ~x421 & ~x422 & ~x423 & ~x446 & ~x447 & ~x448 & ~x449 & ~x450 & ~x475 & ~x506 & ~x508 & ~x529 & ~x530 & ~x533 & ~x535 & ~x536 & ~x556 & ~x557 & ~x558 & ~x559 & ~x560 & ~x562 & ~x563 & ~x564 & ~x565 & ~x583 & ~x584 & ~x586 & ~x589 & ~x590 & ~x591 & ~x592 & ~x611 & ~x612 & ~x614 & ~x615 & ~x617 & ~x619 & ~x620 & ~x621 & ~x637 & ~x638 & ~x639 & ~x642 & ~x643 & ~x644 & ~x647 & ~x648 & ~x649 & ~x650 & ~x652 & ~x661 & ~x668 & ~x670 & ~x671 & ~x672 & ~x673 & ~x676 & ~x680 & ~x681 & ~x682 & ~x683 & ~x684 & ~x689 & ~x691 & ~x693 & ~x694 & ~x695 & ~x696 & ~x697 & ~x698 & ~x700 & ~x703 & ~x706 & ~x708 & ~x710 & ~x711 & ~x713 & ~x714 & ~x715 & ~x716 & ~x717 & ~x719 & ~x720 & ~x722 & ~x723 & ~x724 & ~x726 & ~x729 & ~x733 & ~x736 & ~x739 & ~x742 & ~x753 & ~x754 & ~x755 & ~x756 & ~x757 & ~x758 & ~x760 & ~x761 & ~x766 & ~x767 & ~x770 & ~x772 & ~x773 & ~x774 & ~x776 & ~x777 & ~x779 & ~x783;
assign c640 =  x433 &  x440 &  x574 &  x575 &  x601 &  x602 & ~x11 & ~x13 & ~x16 & ~x18 & ~x31 & ~x33 & ~x35 & ~x39 & ~x42 & ~x43 & ~x44 & ~x51 & ~x59 & ~x64 & ~x76 & ~x77 & ~x78 & ~x79 & ~x81 & ~x85 & ~x87 & ~x88 & ~x92 & ~x93 & ~x116 & ~x117 & ~x119 & ~x137 & ~x139 & ~x141 & ~x142 & ~x148 & ~x166 & ~x168 & ~x171 & ~x172 & ~x195 & ~x199 & ~x202 & ~x220 & ~x221 & ~x222 & ~x230 & ~x254 & ~x259 & ~x277 & ~x280 & ~x283 & ~x285 & ~x310 & ~x311 & ~x339 & ~x364 & ~x367 & ~x390 & ~x394 & ~x421 & ~x444 & ~x448 & ~x473 & ~x474 & ~x476 & ~x506 & ~x507 & ~x532 & ~x563 & ~x592 & ~x616 & ~x621 & ~x622 & ~x646 & ~x647 & ~x651 & ~x656 & ~x657 & ~x675 & ~x676 & ~x684 & ~x687 & ~x688 & ~x689 & ~x690 & ~x692 & ~x702 & ~x704 & ~x707 & ~x710 & ~x712 & ~x714 & ~x718 & ~x719 & ~x721 & ~x729 & ~x737 & ~x739 & ~x747 & ~x750 & ~x751 & ~x757 & ~x765 & ~x766 & ~x774 & ~x776;
assign c642 =  x34;
assign c644 =  x375 &  x431 &  x459 & ~x3 & ~x11 & ~x13 & ~x17 & ~x18 & ~x25 & ~x39 & ~x40 & ~x57 & ~x58 & ~x66 & ~x76 & ~x82 & ~x85 & ~x112 & ~x139 & ~x143 & ~x164 & ~x167 & ~x171 & ~x173 & ~x177 & ~x190 & ~x196 & ~x215 & ~x221 & ~x227 & ~x229 & ~x230 & ~x243 & ~x251 & ~x272 & ~x285 & ~x297 & ~x302 & ~x306 & ~x308 & ~x311 & ~x336 & ~x359 & ~x360 & ~x372 & ~x398 & ~x425 & ~x427 & ~x445 & ~x504 & ~x505 & ~x526 & ~x532 & ~x533 & ~x534 & ~x536 & ~x556 & ~x558 & ~x565 & ~x566 & ~x589 & ~x593 & ~x637 & ~x647 & ~x650 & ~x653 & ~x665 & ~x666 & ~x670 & ~x677 & ~x679 & ~x684 & ~x694 & ~x695 & ~x715 & ~x721 & ~x723 & ~x729 & ~x732 & ~x733 & ~x738 & ~x744 & ~x746 & ~x753 & ~x760 & ~x762 & ~x768 & ~x769 & ~x773 & ~x778 & ~x780 & ~x782 & ~x783;
assign c646 =  x387 &  x426;
assign c648 =  x297 & ~x156 & ~x183 & ~x237 & ~x277 & ~x292 & ~x338 & ~x723 & ~x764;
assign c650 = ~x212 & ~x237 & ~x318 & ~x429 & ~x665;
assign c652 =  x600 &  x603 & ~x0 & ~x1 & ~x10 & ~x24 & ~x26 & ~x27 & ~x28 & ~x29 & ~x36 & ~x38 & ~x42 & ~x43 & ~x44 & ~x48 & ~x52 & ~x53 & ~x54 & ~x58 & ~x59 & ~x60 & ~x64 & ~x68 & ~x69 & ~x78 & ~x79 & ~x80 & ~x82 & ~x83 & ~x90 & ~x91 & ~x110 & ~x114 & ~x116 & ~x117 & ~x118 & ~x120 & ~x123 & ~x133 & ~x138 & ~x139 & ~x140 & ~x142 & ~x147 & ~x164 & ~x168 & ~x170 & ~x173 & ~x175 & ~x177 & ~x191 & ~x192 & ~x194 & ~x196 & ~x197 & ~x199 & ~x201 & ~x202 & ~x205 & ~x220 & ~x221 & ~x225 & ~x228 & ~x229 & ~x231 & ~x232 & ~x242 & ~x247 & ~x248 & ~x249 & ~x252 & ~x253 & ~x255 & ~x256 & ~x257 & ~x259 & ~x270 & ~x272 & ~x273 & ~x278 & ~x279 & ~x282 & ~x287 & ~x302 & ~x304 & ~x306 & ~x307 & ~x309 & ~x311 & ~x312 & ~x335 & ~x342 & ~x363 & ~x364 & ~x365 & ~x368 & ~x390 & ~x392 & ~x393 & ~x395 & ~x396 & ~x407 & ~x418 & ~x420 & ~x446 & ~x447 & ~x450 & ~x452 & ~x478 & ~x502 & ~x503 & ~x504 & ~x507 & ~x508 & ~x509 & ~x533 & ~x535 & ~x536 & ~x538 & ~x556 & ~x560 & ~x561 & ~x562 & ~x563 & ~x565 & ~x585 & ~x587 & ~x588 & ~x589 & ~x591 & ~x592 & ~x593 & ~x594 & ~x610 & ~x611 & ~x622 & ~x623 & ~x624 & ~x636 & ~x640 & ~x645 & ~x648 & ~x649 & ~x653 & ~x654 & ~x666 & ~x670 & ~x680 & ~x684 & ~x685 & ~x686 & ~x689 & ~x693 & ~x695 & ~x697 & ~x699 & ~x700 & ~x704 & ~x708 & ~x709 & ~x710 & ~x715 & ~x718 & ~x719 & ~x720 & ~x721 & ~x724 & ~x727 & ~x728 & ~x729 & ~x730 & ~x731 & ~x733 & ~x737 & ~x738 & ~x741 & ~x744 & ~x751 & ~x754 & ~x757 & ~x760 & ~x761 & ~x763 & ~x764 & ~x765 & ~x768 & ~x772 & ~x775 & ~x777 & ~x778 & ~x780;
assign c654 =  x88;
assign c656 =  x338;
assign c658 =  x320 &  x347 &  x429 &  x430 &  x457 &  x485 &  x513 &  x569 & ~x5 & ~x24 & ~x31 & ~x34 & ~x37 & ~x45 & ~x51 & ~x52 & ~x61 & ~x62 & ~x65 & ~x71 & ~x76 & ~x81 & ~x99 & ~x112 & ~x123 & ~x125 & ~x136 & ~x151 & ~x153 & ~x166 & ~x171 & ~x175 & ~x177 & ~x178 & ~x179 & ~x180 & ~x190 & ~x195 & ~x199 & ~x207 & ~x217 & ~x218 & ~x225 & ~x226 & ~x234 & ~x245 & ~x246 & ~x248 & ~x251 & ~x261 & ~x273 & ~x277 & ~x281 & ~x283 & ~x289 & ~x309 & ~x334 & ~x337 & ~x341 & ~x366 & ~x393 & ~x416 & ~x417 & ~x446 & ~x449 & ~x450 & ~x474 & ~x479 & ~x499 & ~x500 & ~x526 & ~x527 & ~x558 & ~x560 & ~x582 & ~x588 & ~x607 & ~x651 & ~x661 & ~x663 & ~x667 & ~x668 & ~x672 & ~x676 & ~x678 & ~x691 & ~x705 & ~x715 & ~x721 & ~x728 & ~x733 & ~x742 & ~x745 & ~x756 & ~x758 & ~x759 & ~x762 & ~x777 & ~x781;
assign c660 =  x295 &  x322 &  x570 & ~x236 & ~x238 & ~x265;
assign c662 = ~x15 & ~x32 & ~x56 & ~x190 & ~x195 & ~x231 & ~x232 & ~x299 & ~x324 & ~x328 & ~x361 & ~x385 & ~x421 & ~x485 & ~x498 & ~x536 & ~x584 & ~x598 & ~x636 & ~x718 & ~x758 & ~x766 & ~x783;
assign c664 =  x370 &  x398 &  x454 & ~x58 & ~x199 & ~x214 & ~x239 & ~x266 & ~x293 & ~x364 & ~x402 & ~x655 & ~x664 & ~x686;
assign c666 =  x156 &  x210 &  x293 &  x347 &  x375 &  x430 & ~x9 & ~x12 & ~x15 & ~x17 & ~x22 & ~x23 & ~x24 & ~x29 & ~x43 & ~x45 & ~x58 & ~x59 & ~x63 & ~x64 & ~x70 & ~x76 & ~x82 & ~x87 & ~x88 & ~x91 & ~x95 & ~x109 & ~x113 & ~x122 & ~x125 & ~x146 & ~x148 & ~x151 & ~x163 & ~x164 & ~x165 & ~x166 & ~x168 & ~x173 & ~x174 & ~x177 & ~x191 & ~x195 & ~x201 & ~x206 & ~x207 & ~x226 & ~x233 & ~x248 & ~x268 & ~x270 & ~x279 & ~x284 & ~x285 & ~x286 & ~x287 & ~x308 & ~x310 & ~x316 & ~x334 & ~x337 & ~x339 & ~x340 & ~x341 & ~x361 & ~x368 & ~x388 & ~x389 & ~x391 & ~x393 & ~x396 & ~x397 & ~x418 & ~x423 & ~x444 & ~x446 & ~x447 & ~x452 & ~x473 & ~x477 & ~x478 & ~x499 & ~x502 & ~x506 & ~x529 & ~x531 & ~x533 & ~x537 & ~x555 & ~x565 & ~x583 & ~x615 & ~x616 & ~x620 & ~x636 & ~x637 & ~x639 & ~x640 & ~x646 & ~x651 & ~x653 & ~x666 & ~x667 & ~x668 & ~x679 & ~x680 & ~x691 & ~x699 & ~x700 & ~x708 & ~x710 & ~x712 & ~x727 & ~x729 & ~x730 & ~x734 & ~x741 & ~x745 & ~x749 & ~x750 & ~x771 & ~x773 & ~x775 & ~x778 & ~x782 & ~x783;
assign c668 =  x401 &  x457 &  x514 &  x571 & ~x1 & ~x7 & ~x9 & ~x14 & ~x16 & ~x17 & ~x28 & ~x38 & ~x54 & ~x56 & ~x58 & ~x59 & ~x63 & ~x64 & ~x66 & ~x68 & ~x72 & ~x74 & ~x75 & ~x77 & ~x78 & ~x83 & ~x88 & ~x89 & ~x98 & ~x108 & ~x109 & ~x118 & ~x167 & ~x171 & ~x172 & ~x197 & ~x202 & ~x226 & ~x228 & ~x248 & ~x250 & ~x257 & ~x272 & ~x276 & ~x279 & ~x286 & ~x299 & ~x303 & ~x304 & ~x314 & ~x315 & ~x334 & ~x335 & ~x343 & ~x363 & ~x364 & ~x365 & ~x366 & ~x385 & ~x387 & ~x390 & ~x392 & ~x395 & ~x416 & ~x418 & ~x420 & ~x422 & ~x444 & ~x450 & ~x471 & ~x474 & ~x475 & ~x476 & ~x477 & ~x478 & ~x481 & ~x482 & ~x530 & ~x531 & ~x536 & ~x557 & ~x564 & ~x567 & ~x584 & ~x590 & ~x594 & ~x595 & ~x613 & ~x614 & ~x615 & ~x623 & ~x624 & ~x638 & ~x641 & ~x646 & ~x652 & ~x668 & ~x674 & ~x689 & ~x705 & ~x712 & ~x718 & ~x719 & ~x722 & ~x726 & ~x727 & ~x729 & ~x736 & ~x747 & ~x753 & ~x754 & ~x755 & ~x757 & ~x758 & ~x768 & ~x779 & ~x783;
assign c674 =  x134;
assign c676 =  x159 &  x239 &  x266 &  x293 &  x294 &  x320 &  x321 &  x348 &  x375 & ~x1 & ~x23 & ~x27 & ~x30 & ~x31 & ~x33 & ~x39 & ~x41 & ~x42 & ~x46 & ~x58 & ~x63 & ~x68 & ~x72 & ~x80 & ~x81 & ~x83 & ~x84 & ~x85 & ~x86 & ~x92 & ~x93 & ~x96 & ~x98 & ~x110 & ~x113 & ~x114 & ~x122 & ~x123 & ~x128 & ~x139 & ~x141 & ~x147 & ~x148 & ~x152 & ~x153 & ~x154 & ~x155 & ~x171 & ~x174 & ~x175 & ~x177 & ~x179 & ~x180 & ~x181 & ~x182 & ~x196 & ~x198 & ~x206 & ~x207 & ~x208 & ~x232 & ~x234 & ~x246 & ~x252 & ~x260 & ~x262 & ~x270 & ~x273 & ~x275 & ~x277 & ~x286 & ~x287 & ~x288 & ~x304 & ~x315 & ~x330 & ~x335 & ~x336 & ~x337 & ~x362 & ~x364 & ~x368 & ~x369 & ~x394 & ~x395 & ~x419 & ~x422 & ~x443 & ~x445 & ~x446 & ~x451 & ~x472 & ~x474 & ~x477 & ~x502 & ~x506 & ~x507 & ~x526 & ~x527 & ~x528 & ~x532 & ~x560 & ~x586 & ~x587 & ~x589 & ~x613 & ~x616 & ~x617 & ~x618 & ~x621 & ~x638 & ~x642 & ~x649 & ~x650 & ~x662 & ~x665 & ~x666 & ~x667 & ~x674 & ~x680 & ~x681 & ~x682 & ~x694 & ~x697 & ~x698 & ~x700 & ~x713 & ~x722 & ~x736 & ~x742 & ~x743 & ~x744 & ~x746 & ~x754 & ~x755 & ~x766 & ~x769 & ~x771 & ~x772 & ~x776 & ~x782;
assign c678 = ~x15 & ~x22 & ~x26 & ~x29 & ~x46 & ~x57 & ~x65 & ~x86 & ~x92 & ~x96 & ~x104 & ~x120 & ~x124 & ~x140 & ~x143 & ~x152 & ~x153 & ~x170 & ~x175 & ~x177 & ~x180 & ~x196 & ~x202 & ~x208 & ~x221 & ~x235 & ~x243 & ~x247 & ~x249 & ~x258 & ~x263 & ~x289 & ~x303 & ~x307 & ~x311 & ~x316 & ~x324 & ~x327 & ~x329 & ~x330 & ~x331 & ~x338 & ~x399 & ~x401 & ~x417 & ~x428 & ~x447 & ~x470 & ~x473 & ~x526 & ~x527 & ~x533 & ~x536 & ~x558 & ~x562 & ~x617 & ~x636 & ~x639 & ~x647 & ~x661 & ~x671 & ~x673 & ~x684 & ~x686 & ~x688 & ~x712 & ~x725 & ~x751 & ~x765 & ~x770;
assign c680 =  x543 & ~x19 & ~x20 & ~x30 & ~x40 & ~x46 & ~x47 & ~x49 & ~x51 & ~x62 & ~x65 & ~x69 & ~x70 & ~x90 & ~x135 & ~x136 & ~x168 & ~x169 & ~x192 & ~x203 & ~x244 & ~x253 & ~x271 & ~x274 & ~x285 & ~x298 & ~x301 & ~x302 & ~x324 & ~x326 & ~x327 & ~x330 & ~x334 & ~x339 & ~x350 & ~x388 & ~x448 & ~x533 & ~x537 & ~x559 & ~x561 & ~x564 & ~x612 & ~x614 & ~x621 & ~x645 & ~x670 & ~x676 & ~x680 & ~x681 & ~x689 & ~x690 & ~x693 & ~x698 & ~x700 & ~x706 & ~x727 & ~x741 & ~x743 & ~x751 & ~x769 & ~x770;
assign c682 =  x77;
assign c684 =  x321 & ~x48 & ~x87 & ~x90 & ~x124 & ~x139 & ~x164 & ~x181 & ~x254 & ~x269 & ~x297 & ~x316 & ~x341 & ~x351 & ~x387 & ~x478 & ~x479 & ~x498 & ~x582 & ~x596 & ~x635 & ~x653 & ~x663 & ~x692 & ~x781;
assign c686 =  x547 & ~x131 & ~x162 & ~x185 & ~x187 & ~x239 & ~x264 & ~x613 & ~x624 & ~x665;
assign c688 =  x431 &  x459 & ~x6 & ~x13 & ~x17 & ~x18 & ~x22 & ~x24 & ~x32 & ~x39 & ~x42 & ~x48 & ~x58 & ~x59 & ~x60 & ~x66 & ~x81 & ~x87 & ~x90 & ~x104 & ~x108 & ~x111 & ~x113 & ~x121 & ~x140 & ~x143 & ~x145 & ~x176 & ~x198 & ~x220 & ~x224 & ~x225 & ~x230 & ~x231 & ~x246 & ~x249 & ~x255 & ~x259 & ~x277 & ~x286 & ~x295 & ~x298 & ~x308 & ~x314 & ~x323 & ~x327 & ~x329 & ~x331 & ~x334 & ~x337 & ~x338 & ~x341 & ~x342 & ~x357 & ~x363 & ~x365 & ~x369 & ~x386 & ~x421 & ~x445 & ~x449 & ~x477 & ~x535 & ~x537 & ~x558 & ~x565 & ~x583 & ~x584 & ~x590 & ~x620 & ~x642 & ~x654 & ~x655 & ~x665 & ~x668 & ~x675 & ~x677 & ~x678 & ~x683 & ~x685 & ~x686 & ~x692 & ~x695 & ~x705 & ~x709 & ~x710 & ~x716 & ~x721 & ~x722 & ~x724 & ~x739 & ~x744 & ~x746 & ~x750 & ~x756 & ~x760 & ~x768 & ~x776 & ~x780 & ~x781;
assign c690 =  x701;
assign c692 =  x428 &  x517 &  x541 &  x545 & ~x201 & ~x269 & ~x297 & ~x305 & ~x341 & ~x618 & ~x715 & ~x718 & ~x725;
assign c694 =  x546 & ~x99 & ~x188 & ~x236 & ~x279 & ~x293 & ~x319 & ~x665 & ~x701;
assign c696 =  x388 & ~x246;
assign c698 =  x516 & ~x30 & ~x50 & ~x56 & ~x82 & ~x84 & ~x91 & ~x108 & ~x111 & ~x163 & ~x164 & ~x201 & ~x205 & ~x216 & ~x251 & ~x252 & ~x271 & ~x285 & ~x296 & ~x301 & ~x302 & ~x306 & ~x350 & ~x446 & ~x471 & ~x500 & ~x507 & ~x567 & ~x616 & ~x644 & ~x651 & ~x665 & ~x678 & ~x680 & ~x683 & ~x693 & ~x695 & ~x711 & ~x718 & ~x729 & ~x735 & ~x743 & ~x747;
assign c6100 = ~x17 & ~x28 & ~x60 & ~x106 & ~x111 & ~x132 & ~x137 & ~x165 & ~x188 & ~x214 & ~x215 & ~x216 & ~x239 & ~x293 & ~x294 & ~x305 & ~x307 & ~x314 & ~x349 & ~x501 & ~x614 & ~x645 & ~x658 & ~x667 & ~x718 & ~x734 & ~x745;
assign c6102 =  x545 &  x574 & ~x3 & ~x51 & ~x100 & ~x102 & ~x132 & ~x141 & ~x167 & ~x189 & ~x209 & ~x211 & ~x219 & ~x250 & ~x292 & ~x639 & ~x654 & ~x725;
assign c6104 =  x348 & ~x1 & ~x2 & ~x3 & ~x4 & ~x9 & ~x10 & ~x11 & ~x12 & ~x13 & ~x15 & ~x16 & ~x19 & ~x21 & ~x22 & ~x24 & ~x25 & ~x27 & ~x29 & ~x32 & ~x33 & ~x35 & ~x37 & ~x38 & ~x47 & ~x48 & ~x51 & ~x52 & ~x53 & ~x54 & ~x56 & ~x57 & ~x60 & ~x61 & ~x62 & ~x63 & ~x67 & ~x70 & ~x80 & ~x84 & ~x85 & ~x89 & ~x92 & ~x93 & ~x95 & ~x96 & ~x97 & ~x110 & ~x113 & ~x114 & ~x115 & ~x116 & ~x117 & ~x118 & ~x120 & ~x122 & ~x124 & ~x125 & ~x141 & ~x142 & ~x149 & ~x150 & ~x151 & ~x152 & ~x166 & ~x167 & ~x169 & ~x170 & ~x172 & ~x174 & ~x175 & ~x192 & ~x193 & ~x196 & ~x199 & ~x200 & ~x202 & ~x204 & ~x205 & ~x206 & ~x208 & ~x217 & ~x218 & ~x220 & ~x221 & ~x222 & ~x223 & ~x225 & ~x228 & ~x229 & ~x231 & ~x232 & ~x244 & ~x247 & ~x251 & ~x252 & ~x254 & ~x257 & ~x260 & ~x262 & ~x271 & ~x274 & ~x275 & ~x277 & ~x278 & ~x279 & ~x280 & ~x282 & ~x283 & ~x284 & ~x301 & ~x303 & ~x304 & ~x305 & ~x306 & ~x307 & ~x308 & ~x309 & ~x310 & ~x312 & ~x314 & ~x315 & ~x332 & ~x333 & ~x334 & ~x338 & ~x339 & ~x341 & ~x343 & ~x344 & ~x365 & ~x368 & ~x369 & ~x389 & ~x390 & ~x391 & ~x392 & ~x393 & ~x395 & ~x397 & ~x416 & ~x418 & ~x420 & ~x421 & ~x423 & ~x425 & ~x444 & ~x447 & ~x448 & ~x450 & ~x451 & ~x452 & ~x453 & ~x472 & ~x473 & ~x475 & ~x476 & ~x478 & ~x479 & ~x480 & ~x498 & ~x499 & ~x503 & ~x505 & ~x530 & ~x531 & ~x532 & ~x533 & ~x534 & ~x553 & ~x555 & ~x557 & ~x561 & ~x563 & ~x579 & ~x580 & ~x581 & ~x583 & ~x585 & ~x586 & ~x588 & ~x607 & ~x608 & ~x610 & ~x614 & ~x617 & ~x622 & ~x632 & ~x635 & ~x637 & ~x641 & ~x643 & ~x644 & ~x645 & ~x649 & ~x650 & ~x651 & ~x652 & ~x654 & ~x657 & ~x658 & ~x659 & ~x660 & ~x662 & ~x663 & ~x668 & ~x671 & ~x672 & ~x676 & ~x680 & ~x682 & ~x684 & ~x688 & ~x689 & ~x691 & ~x692 & ~x694 & ~x695 & ~x696 & ~x697 & ~x698 & ~x702 & ~x703 & ~x704 & ~x709 & ~x710 & ~x711 & ~x714 & ~x715 & ~x717 & ~x718 & ~x722 & ~x725 & ~x726 & ~x729 & ~x730 & ~x731 & ~x732 & ~x733 & ~x736 & ~x737 & ~x739 & ~x740 & ~x741 & ~x742 & ~x743 & ~x744 & ~x750 & ~x752 & ~x753 & ~x755 & ~x756 & ~x757 & ~x759 & ~x762 & ~x764 & ~x765 & ~x767 & ~x769 & ~x773 & ~x774 & ~x776 & ~x777 & ~x779 & ~x780 & ~x783;
assign c6106 =  x317 &  x373 &  x400 &  x428 &  x429 &  x485 &  x542 & ~x10 & ~x15 & ~x18 & ~x30 & ~x56 & ~x59 & ~x75 & ~x79 & ~x80 & ~x82 & ~x87 & ~x91 & ~x105 & ~x109 & ~x111 & ~x112 & ~x116 & ~x119 & ~x140 & ~x141 & ~x142 & ~x170 & ~x171 & ~x173 & ~x193 & ~x197 & ~x225 & ~x227 & ~x229 & ~x243 & ~x252 & ~x274 & ~x276 & ~x277 & ~x281 & ~x284 & ~x306 & ~x307 & ~x308 & ~x332 & ~x333 & ~x334 & ~x340 & ~x366 & ~x367 & ~x368 & ~x394 & ~x395 & ~x397 & ~x423 & ~x425 & ~x446 & ~x451 & ~x453 & ~x476 & ~x477 & ~x481 & ~x504 & ~x508 & ~x509 & ~x529 & ~x531 & ~x534 & ~x537 & ~x538 & ~x557 & ~x558 & ~x565 & ~x590 & ~x592 & ~x594 & ~x612 & ~x623 & ~x639 & ~x641 & ~x648 & ~x651 & ~x654 & ~x664 & ~x665 & ~x666 & ~x672 & ~x673 & ~x676 & ~x678 & ~x679 & ~x685 & ~x686 & ~x688 & ~x693 & ~x694 & ~x698 & ~x703 & ~x704 & ~x707 & ~x710 & ~x711 & ~x712 & ~x714 & ~x715 & ~x722 & ~x723 & ~x725 & ~x727 & ~x729 & ~x732 & ~x736 & ~x748 & ~x750 & ~x752 & ~x753 & ~x755 & ~x764 & ~x768;
assign c6108 =  x431 & ~x5 & ~x18 & ~x22 & ~x25 & ~x29 & ~x30 & ~x32 & ~x37 & ~x40 & ~x42 & ~x44 & ~x47 & ~x54 & ~x56 & ~x59 & ~x60 & ~x61 & ~x64 & ~x65 & ~x69 & ~x70 & ~x71 & ~x98 & ~x111 & ~x112 & ~x114 & ~x117 & ~x118 & ~x126 & ~x141 & ~x144 & ~x146 & ~x147 & ~x151 & ~x170 & ~x178 & ~x179 & ~x193 & ~x201 & ~x208 & ~x220 & ~x222 & ~x223 & ~x225 & ~x231 & ~x236 & ~x247 & ~x249 & ~x252 & ~x255 & ~x261 & ~x262 & ~x277 & ~x279 & ~x286 & ~x289 & ~x290 & ~x299 & ~x300 & ~x301 & ~x305 & ~x312 & ~x313 & ~x331 & ~x335 & ~x339 & ~x341 & ~x342 & ~x359 & ~x361 & ~x366 & ~x369 & ~x372 & ~x388 & ~x393 & ~x394 & ~x395 & ~x415 & ~x418 & ~x421 & ~x424 & ~x447 & ~x475 & ~x478 & ~x505 & ~x506 & ~x526 & ~x528 & ~x530 & ~x535 & ~x553 & ~x557 & ~x561 & ~x564 & ~x590 & ~x591 & ~x610 & ~x611 & ~x615 & ~x616 & ~x619 & ~x638 & ~x641 & ~x642 & ~x651 & ~x663 & ~x665 & ~x669 & ~x670 & ~x685 & ~x687 & ~x688 & ~x691 & ~x697 & ~x699 & ~x709 & ~x713 & ~x723 & ~x724 & ~x727 & ~x728 & ~x731 & ~x735 & ~x740 & ~x750 & ~x756 & ~x762 & ~x776 & ~x783;
assign c6110 =  x51;
assign c6112 =  x546 & ~x185 & ~x294 & ~x569 & ~x656;
assign c6114 =  x92;
assign c6116 =  x430 &  x457 &  x485 &  x513 &  x541 & ~x0 & ~x2 & ~x5 & ~x15 & ~x17 & ~x18 & ~x19 & ~x23 & ~x24 & ~x25 & ~x30 & ~x31 & ~x33 & ~x34 & ~x38 & ~x39 & ~x40 & ~x41 & ~x44 & ~x45 & ~x46 & ~x47 & ~x49 & ~x50 & ~x51 & ~x54 & ~x57 & ~x62 & ~x64 & ~x72 & ~x74 & ~x76 & ~x80 & ~x82 & ~x83 & ~x86 & ~x89 & ~x92 & ~x98 & ~x112 & ~x117 & ~x118 & ~x119 & ~x122 & ~x126 & ~x137 & ~x138 & ~x140 & ~x142 & ~x143 & ~x151 & ~x152 & ~x167 & ~x170 & ~x172 & ~x174 & ~x175 & ~x178 & ~x196 & ~x198 & ~x201 & ~x204 & ~x225 & ~x229 & ~x233 & ~x247 & ~x248 & ~x254 & ~x255 & ~x256 & ~x258 & ~x260 & ~x261 & ~x274 & ~x278 & ~x285 & ~x298 & ~x300 & ~x301 & ~x302 & ~x304 & ~x305 & ~x306 & ~x308 & ~x309 & ~x311 & ~x312 & ~x313 & ~x325 & ~x326 & ~x327 & ~x328 & ~x334 & ~x335 & ~x338 & ~x355 & ~x356 & ~x357 & ~x361 & ~x362 & ~x363 & ~x364 & ~x365 & ~x367 & ~x386 & ~x387 & ~x388 & ~x389 & ~x390 & ~x391 & ~x393 & ~x394 & ~x396 & ~x415 & ~x417 & ~x419 & ~x420 & ~x421 & ~x423 & ~x425 & ~x450 & ~x451 & ~x453 & ~x471 & ~x473 & ~x475 & ~x477 & ~x478 & ~x499 & ~x500 & ~x504 & ~x505 & ~x508 & ~x510 & ~x527 & ~x531 & ~x534 & ~x537 & ~x554 & ~x555 & ~x561 & ~x583 & ~x584 & ~x585 & ~x587 & ~x590 & ~x591 & ~x592 & ~x593 & ~x614 & ~x616 & ~x620 & ~x637 & ~x639 & ~x646 & ~x647 & ~x649 & ~x650 & ~x671 & ~x675 & ~x676 & ~x680 & ~x682 & ~x691 & ~x693 & ~x698 & ~x699 & ~x700 & ~x714 & ~x717 & ~x719 & ~x720 & ~x722 & ~x725 & ~x727 & ~x729 & ~x730 & ~x731 & ~x733 & ~x734 & ~x739 & ~x742 & ~x744 & ~x745 & ~x748 & ~x752 & ~x753 & ~x754 & ~x755 & ~x757 & ~x759 & ~x760 & ~x764 & ~x767 & ~x768 & ~x775 & ~x776 & ~x780;
assign c6118 =  x352 & ~x54 & ~x240 & ~x243 & ~x435 & ~x491;
assign c6120 =  x373 &  x429 &  x457 &  x569 & ~x0 & ~x2 & ~x13 & ~x17 & ~x23 & ~x24 & ~x27 & ~x29 & ~x34 & ~x55 & ~x60 & ~x62 & ~x65 & ~x75 & ~x84 & ~x90 & ~x94 & ~x107 & ~x111 & ~x121 & ~x135 & ~x144 & ~x145 & ~x149 & ~x162 & ~x168 & ~x170 & ~x176 & ~x194 & ~x218 & ~x219 & ~x242 & ~x243 & ~x244 & ~x246 & ~x247 & ~x253 & ~x269 & ~x275 & ~x281 & ~x303 & ~x306 & ~x307 & ~x308 & ~x312 & ~x339 & ~x366 & ~x390 & ~x392 & ~x445 & ~x448 & ~x449 & ~x473 & ~x475 & ~x478 & ~x506 & ~x529 & ~x534 & ~x557 & ~x562 & ~x566 & ~x585 & ~x592 & ~x593 & ~x594 & ~x621 & ~x638 & ~x641 & ~x648 & ~x650 & ~x652 & ~x653 & ~x680 & ~x681 & ~x686 & ~x688 & ~x689 & ~x690 & ~x693 & ~x695 & ~x708 & ~x716 & ~x718 & ~x719 & ~x721 & ~x722 & ~x724 & ~x726 & ~x733 & ~x736 & ~x749 & ~x753 & ~x757 & ~x760 & ~x762 & ~x779 & ~x782;
assign c6122 =  x460 &  x488 &  x523 &  x575 & ~x0 & ~x1 & ~x11 & ~x17 & ~x19 & ~x22 & ~x29 & ~x36 & ~x48 & ~x52 & ~x53 & ~x54 & ~x57 & ~x59 & ~x86 & ~x120 & ~x134 & ~x146 & ~x161 & ~x165 & ~x166 & ~x169 & ~x194 & ~x199 & ~x202 & ~x216 & ~x223 & ~x226 & ~x246 & ~x250 & ~x253 & ~x257 & ~x274 & ~x275 & ~x278 & ~x302 & ~x332 & ~x334 & ~x340 & ~x367 & ~x395 & ~x451 & ~x452 & ~x476 & ~x504 & ~x529 & ~x535 & ~x536 & ~x557 & ~x562 & ~x565 & ~x566 & ~x585 & ~x586 & ~x614 & ~x620 & ~x625 & ~x635 & ~x636 & ~x639 & ~x648 & ~x650 & ~x665 & ~x667 & ~x681 & ~x693 & ~x694 & ~x705 & ~x712 & ~x717 & ~x720 & ~x722 & ~x725 & ~x735 & ~x736 & ~x738 & ~x741 & ~x742 & ~x752 & ~x760 & ~x777 & ~x778 & ~x782;
assign c6124 =  x345 &  x400 &  x540 & ~x0 & ~x9 & ~x15 & ~x19 & ~x23 & ~x29 & ~x52 & ~x63 & ~x77 & ~x83 & ~x91 & ~x114 & ~x118 & ~x146 & ~x151 & ~x168 & ~x169 & ~x172 & ~x176 & ~x217 & ~x220 & ~x223 & ~x225 & ~x228 & ~x246 & ~x255 & ~x259 & ~x271 & ~x272 & ~x286 & ~x296 & ~x338 & ~x362 & ~x365 & ~x447 & ~x474 & ~x506 & ~x556 & ~x558 & ~x560 & ~x586 & ~x589 & ~x591 & ~x609 & ~x611 & ~x614 & ~x615 & ~x620 & ~x621 & ~x640 & ~x645 & ~x654 & ~x663 & ~x667 & ~x670 & ~x678 & ~x691 & ~x692 & ~x697 & ~x699 & ~x705 & ~x708 & ~x715 & ~x716 & ~x728 & ~x739 & ~x745 & ~x764 & ~x781;
assign c6126 =  x518 &  x546 & ~x0 & ~x1 & ~x8 & ~x9 & ~x13 & ~x14 & ~x22 & ~x28 & ~x38 & ~x42 & ~x73 & ~x78 & ~x85 & ~x92 & ~x111 & ~x117 & ~x136 & ~x138 & ~x139 & ~x141 & ~x168 & ~x190 & ~x192 & ~x196 & ~x197 & ~x200 & ~x202 & ~x203 & ~x218 & ~x219 & ~x220 & ~x224 & ~x243 & ~x245 & ~x246 & ~x250 & ~x258 & ~x275 & ~x278 & ~x279 & ~x298 & ~x303 & ~x324 & ~x334 & ~x350 & ~x393 & ~x451 & ~x474 & ~x475 & ~x477 & ~x479 & ~x502 & ~x556 & ~x560 & ~x563 & ~x586 & ~x593 & ~x613 & ~x614 & ~x621 & ~x652 & ~x653 & ~x654 & ~x655 & ~x666 & ~x676 & ~x687 & ~x689 & ~x693 & ~x694 & ~x698 & ~x705 & ~x708 & ~x716 & ~x721 & ~x729 & ~x732 & ~x737 & ~x739 & ~x749 & ~x751 & ~x758 & ~x762 & ~x764 & ~x765 & ~x766 & ~x767 & ~x768 & ~x773 & ~x775 & ~x780 & ~x782;
assign c6128 =  x460 & ~x28 & ~x45 & ~x80 & ~x97 & ~x115 & ~x145 & ~x180 & ~x234 & ~x245 & ~x248 & ~x256 & ~x274 & ~x299 & ~x319 & ~x327 & ~x337 & ~x355 & ~x384 & ~x455 & ~x474 & ~x481 & ~x499 & ~x634 & ~x637 & ~x657 & ~x667 & ~x670 & ~x679 & ~x743 & ~x748;
assign c6130 =  x428 &  x543 &  x544 &  x572 &  x573 & ~x1 & ~x10 & ~x13 & ~x18 & ~x19 & ~x20 & ~x50 & ~x57 & ~x89 & ~x115 & ~x118 & ~x139 & ~x142 & ~x168 & ~x193 & ~x198 & ~x222 & ~x223 & ~x225 & ~x227 & ~x268 & ~x270 & ~x281 & ~x285 & ~x301 & ~x306 & ~x307 & ~x309 & ~x335 & ~x368 & ~x418 & ~x446 & ~x448 & ~x504 & ~x507 & ~x534 & ~x561 & ~x648 & ~x679 & ~x685 & ~x689 & ~x701 & ~x703 & ~x732 & ~x736 & ~x745 & ~x747 & ~x749 & ~x759 & ~x762 & ~x776;
assign c6132 =  x376 &  x601 & ~x152 & ~x206 & ~x229 & ~x242 & ~x262 & ~x301 & ~x325 & ~x336 & ~x373 & ~x445 & ~x509 & ~x512 & ~x537 & ~x610 & ~x643;
assign c6134 =  x22;
assign c6136 =  x431 &  x459 & ~x1 & ~x7 & ~x8 & ~x10 & ~x13 & ~x14 & ~x16 & ~x21 & ~x22 & ~x29 & ~x30 & ~x32 & ~x33 & ~x40 & ~x43 & ~x44 & ~x45 & ~x51 & ~x52 & ~x53 & ~x54 & ~x55 & ~x57 & ~x60 & ~x61 & ~x62 & ~x64 & ~x72 & ~x73 & ~x77 & ~x78 & ~x82 & ~x84 & ~x88 & ~x89 & ~x90 & ~x95 & ~x96 & ~x105 & ~x107 & ~x108 & ~x111 & ~x112 & ~x116 & ~x117 & ~x119 & ~x120 & ~x121 & ~x122 & ~x133 & ~x137 & ~x141 & ~x142 & ~x143 & ~x146 & ~x150 & ~x151 & ~x191 & ~x194 & ~x196 & ~x200 & ~x201 & ~x202 & ~x214 & ~x218 & ~x222 & ~x224 & ~x225 & ~x229 & ~x230 & ~x242 & ~x243 & ~x250 & ~x251 & ~x252 & ~x257 & ~x258 & ~x259 & ~x270 & ~x275 & ~x279 & ~x282 & ~x283 & ~x284 & ~x285 & ~x286 & ~x287 & ~x288 & ~x289 & ~x300 & ~x301 & ~x305 & ~x309 & ~x312 & ~x315 & ~x316 & ~x333 & ~x335 & ~x336 & ~x339 & ~x340 & ~x357 & ~x360 & ~x361 & ~x362 & ~x364 & ~x368 & ~x369 & ~x372 & ~x388 & ~x390 & ~x392 & ~x395 & ~x397 & ~x416 & ~x419 & ~x421 & ~x422 & ~x424 & ~x445 & ~x448 & ~x452 & ~x476 & ~x481 & ~x500 & ~x506 & ~x529 & ~x535 & ~x537 & ~x556 & ~x558 & ~x559 & ~x563 & ~x566 & ~x583 & ~x584 & ~x589 & ~x590 & ~x591 & ~x594 & ~x609 & ~x612 & ~x615 & ~x618 & ~x622 & ~x637 & ~x638 & ~x639 & ~x640 & ~x646 & ~x647 & ~x653 & ~x669 & ~x672 & ~x673 & ~x674 & ~x678 & ~x679 & ~x681 & ~x683 & ~x686 & ~x688 & ~x694 & ~x696 & ~x698 & ~x702 & ~x706 & ~x708 & ~x711 & ~x712 & ~x714 & ~x717 & ~x719 & ~x720 & ~x721 & ~x722 & ~x727 & ~x731 & ~x740 & ~x744 & ~x747 & ~x748 & ~x750 & ~x751 & ~x753 & ~x757 & ~x758 & ~x760 & ~x772 & ~x774 & ~x775 & ~x777 & ~x778 & ~x779 & ~x780 & ~x781 & ~x783;
assign c6138 =  x376 &  x432 & ~x3 & ~x9 & ~x11 & ~x18 & ~x25 & ~x26 & ~x34 & ~x40 & ~x41 & ~x43 & ~x44 & ~x47 & ~x52 & ~x53 & ~x55 & ~x59 & ~x60 & ~x61 & ~x66 & ~x71 & ~x85 & ~x91 & ~x93 & ~x95 & ~x97 & ~x113 & ~x115 & ~x120 & ~x122 & ~x126 & ~x146 & ~x147 & ~x150 & ~x151 & ~x152 & ~x172 & ~x176 & ~x178 & ~x179 & ~x181 & ~x198 & ~x203 & ~x204 & ~x221 & ~x233 & ~x235 & ~x251 & ~x255 & ~x256 & ~x259 & ~x260 & ~x263 & ~x264 & ~x275 & ~x281 & ~x282 & ~x285 & ~x288 & ~x291 & ~x302 & ~x303 & ~x304 & ~x319 & ~x328 & ~x332 & ~x334 & ~x339 & ~x342 & ~x344 & ~x357 & ~x367 & ~x370 & ~x371 & ~x372 & ~x389 & ~x390 & ~x396 & ~x397 & ~x398 & ~x422 & ~x423 & ~x444 & ~x445 & ~x447 & ~x451 & ~x470 & ~x471 & ~x475 & ~x505 & ~x534 & ~x559 & ~x565 & ~x580 & ~x588 & ~x592 & ~x609 & ~x616 & ~x638 & ~x643 & ~x647 & ~x648 & ~x650 & ~x651 & ~x661 & ~x663 & ~x667 & ~x670 & ~x676 & ~x677 & ~x687 & ~x689 & ~x708 & ~x721 & ~x728 & ~x730 & ~x735 & ~x737 & ~x739 & ~x740 & ~x744 & ~x746 & ~x747 & ~x748 & ~x750 & ~x751 & ~x752 & ~x761 & ~x763 & ~x767 & ~x777 & ~x783;
assign c6140 =  x405 &  x431 &  x459 &  x600 & ~x2 & ~x5 & ~x17 & ~x23 & ~x33 & ~x34 & ~x40 & ~x54 & ~x60 & ~x70 & ~x83 & ~x90 & ~x92 & ~x95 & ~x123 & ~x153 & ~x180 & ~x196 & ~x207 & ~x208 & ~x222 & ~x223 & ~x225 & ~x255 & ~x260 & ~x275 & ~x277 & ~x303 & ~x315 & ~x316 & ~x394 & ~x444 & ~x448 & ~x449 & ~x472 & ~x479 & ~x500 & ~x508 & ~x527 & ~x559 & ~x579 & ~x589 & ~x614 & ~x616 & ~x633 & ~x647 & ~x649 & ~x665 & ~x668 & ~x675 & ~x677 & ~x681 & ~x692 & ~x694 & ~x707 & ~x708 & ~x714 & ~x715 & ~x718 & ~x730 & ~x736 & ~x737 & ~x739 & ~x750 & ~x757 & ~x762 & ~x769;
assign c6142 =  x215 &  x295 &  x456 & ~x211 & ~x236 & ~x262;
assign c6144 = ~x0 & ~x18 & ~x20 & ~x38 & ~x77 & ~x84 & ~x107 & ~x168 & ~x215 & ~x219 & ~x240 & ~x250 & ~x266 & ~x268 & ~x294 & ~x320 & ~x334 & ~x365 & ~x376 & ~x402 & ~x421 & ~x458 & ~x476 & ~x588 & ~x655 & ~x695 & ~x713 & ~x715 & ~x716 & ~x747 & ~x776;
assign c6146 =  x319 &  x346 &  x347 &  x401 &  x402 &  x429 &  x457 &  x513 &  x541 &  x569 &  x570 & ~x0 & ~x1 & ~x2 & ~x4 & ~x6 & ~x7 & ~x9 & ~x11 & ~x12 & ~x13 & ~x14 & ~x15 & ~x17 & ~x19 & ~x20 & ~x21 & ~x28 & ~x29 & ~x33 & ~x34 & ~x35 & ~x36 & ~x37 & ~x38 & ~x39 & ~x40 & ~x42 & ~x43 & ~x44 & ~x45 & ~x46 & ~x49 & ~x50 & ~x51 & ~x52 & ~x53 & ~x56 & ~x57 & ~x58 & ~x59 & ~x61 & ~x62 & ~x63 & ~x64 & ~x68 & ~x69 & ~x70 & ~x71 & ~x72 & ~x73 & ~x74 & ~x78 & ~x79 & ~x80 & ~x81 & ~x83 & ~x84 & ~x85 & ~x87 & ~x88 & ~x89 & ~x90 & ~x91 & ~x92 & ~x94 & ~x95 & ~x96 & ~x108 & ~x109 & ~x110 & ~x111 & ~x112 & ~x113 & ~x114 & ~x116 & ~x117 & ~x118 & ~x119 & ~x121 & ~x122 & ~x124 & ~x136 & ~x137 & ~x138 & ~x139 & ~x140 & ~x141 & ~x142 & ~x149 & ~x150 & ~x151 & ~x165 & ~x166 & ~x167 & ~x169 & ~x170 & ~x171 & ~x172 & ~x173 & ~x179 & ~x193 & ~x194 & ~x198 & ~x201 & ~x204 & ~x205 & ~x206 & ~x222 & ~x225 & ~x226 & ~x227 & ~x228 & ~x229 & ~x230 & ~x231 & ~x233 & ~x234 & ~x248 & ~x249 & ~x250 & ~x251 & ~x253 & ~x254 & ~x255 & ~x257 & ~x258 & ~x259 & ~x274 & ~x276 & ~x277 & ~x278 & ~x280 & ~x283 & ~x286 & ~x287 & ~x300 & ~x301 & ~x302 & ~x303 & ~x304 & ~x306 & ~x310 & ~x311 & ~x312 & ~x314 & ~x330 & ~x331 & ~x332 & ~x333 & ~x334 & ~x335 & ~x336 & ~x338 & ~x340 & ~x341 & ~x342 & ~x358 & ~x359 & ~x360 & ~x361 & ~x362 & ~x363 & ~x364 & ~x366 & ~x367 & ~x369 & ~x370 & ~x388 & ~x391 & ~x395 & ~x396 & ~x398 & ~x415 & ~x417 & ~x419 & ~x421 & ~x422 & ~x425 & ~x444 & ~x445 & ~x447 & ~x448 & ~x449 & ~x450 & ~x452 & ~x474 & ~x477 & ~x478 & ~x480 & ~x500 & ~x501 & ~x503 & ~x505 & ~x506 & ~x527 & ~x528 & ~x529 & ~x531 & ~x535 & ~x536 & ~x554 & ~x555 & ~x556 & ~x557 & ~x559 & ~x560 & ~x561 & ~x563 & ~x583 & ~x585 & ~x586 & ~x587 & ~x588 & ~x589 & ~x590 & ~x592 & ~x593 & ~x594 & ~x609 & ~x613 & ~x614 & ~x616 & ~x618 & ~x620 & ~x621 & ~x622 & ~x639 & ~x640 & ~x641 & ~x642 & ~x644 & ~x645 & ~x646 & ~x647 & ~x648 & ~x650 & ~x651 & ~x652 & ~x662 & ~x664 & ~x665 & ~x667 & ~x668 & ~x669 & ~x676 & ~x677 & ~x678 & ~x679 & ~x681 & ~x682 & ~x689 & ~x690 & ~x691 & ~x692 & ~x693 & ~x695 & ~x699 & ~x703 & ~x704 & ~x705 & ~x706 & ~x707 & ~x708 & ~x709 & ~x710 & ~x711 & ~x712 & ~x714 & ~x716 & ~x717 & ~x718 & ~x720 & ~x721 & ~x723 & ~x726 & ~x728 & ~x729 & ~x730 & ~x732 & ~x734 & ~x735 & ~x736 & ~x738 & ~x739 & ~x740 & ~x741 & ~x742 & ~x744 & ~x747 & ~x749 & ~x751 & ~x755 & ~x758 & ~x759 & ~x760 & ~x761 & ~x762 & ~x764 & ~x766 & ~x767 & ~x769 & ~x770 & ~x772 & ~x773 & ~x774 & ~x775 & ~x776 & ~x777 & ~x778 & ~x782 & ~x783;
assign c6148 =  x129 &  x157 &  x210 & ~x1 & ~x7 & ~x10 & ~x12 & ~x13 & ~x15 & ~x17 & ~x21 & ~x25 & ~x29 & ~x32 & ~x38 & ~x41 & ~x43 & ~x44 & ~x45 & ~x48 & ~x52 & ~x57 & ~x61 & ~x65 & ~x69 & ~x86 & ~x87 & ~x90 & ~x93 & ~x97 & ~x109 & ~x111 & ~x112 & ~x116 & ~x120 & ~x123 & ~x124 & ~x125 & ~x139 & ~x140 & ~x141 & ~x144 & ~x145 & ~x146 & ~x151 & ~x164 & ~x167 & ~x169 & ~x172 & ~x173 & ~x178 & ~x179 & ~x201 & ~x204 & ~x206 & ~x225 & ~x232 & ~x249 & ~x256 & ~x257 & ~x259 & ~x275 & ~x276 & ~x277 & ~x279 & ~x280 & ~x283 & ~x286 & ~x288 & ~x295 & ~x303 & ~x306 & ~x310 & ~x313 & ~x323 & ~x325 & ~x336 & ~x353 & ~x355 & ~x357 & ~x358 & ~x361 & ~x366 & ~x384 & ~x389 & ~x391 & ~x396 & ~x418 & ~x422 & ~x424 & ~x447 & ~x453 & ~x473 & ~x481 & ~x501 & ~x503 & ~x506 & ~x507 & ~x528 & ~x530 & ~x536 & ~x565 & ~x566 & ~x586 & ~x589 & ~x593 & ~x594 & ~x617 & ~x619 & ~x640 & ~x641 & ~x650 & ~x651 & ~x668 & ~x677 & ~x678 & ~x680 & ~x681 & ~x683 & ~x684 & ~x697 & ~x699 & ~x701 & ~x703 & ~x705 & ~x706 & ~x712 & ~x718 & ~x720 & ~x723 & ~x735 & ~x737 & ~x744 & ~x746 & ~x748 & ~x751 & ~x752 & ~x753 & ~x754 & ~x756 & ~x762 & ~x763 & ~x764 & ~x767 & ~x771 & ~x773 & ~x775 & ~x778;
assign c6150 =  x460 &  x487 & ~x13 & ~x20 & ~x21 & ~x23 & ~x26 & ~x33 & ~x43 & ~x49 & ~x65 & ~x70 & ~x85 & ~x106 & ~x110 & ~x120 & ~x147 & ~x150 & ~x176 & ~x203 & ~x204 & ~x217 & ~x259 & ~x275 & ~x277 & ~x296 & ~x331 & ~x356 & ~x358 & ~x360 & ~x413 & ~x416 & ~x418 & ~x419 & ~x442 & ~x477 & ~x484 & ~x506 & ~x528 & ~x625 & ~x655 & ~x685 & ~x691 & ~x707 & ~x722 & ~x728 & ~x738 & ~x740 & ~x745 & ~x764 & ~x773 & ~x774;
assign c6152 =  x458 &  x515 &  x543 &  x602 & ~x16 & ~x77 & ~x87 & ~x145 & ~x171 & ~x194 & ~x212 & ~x224 & ~x256 & ~x305 & ~x308 & ~x310 & ~x312 & ~x333 & ~x370 & ~x454 & ~x478 & ~x482 & ~x532 & ~x536 & ~x539 & ~x558 & ~x563 & ~x565 & ~x567 & ~x589 & ~x595 & ~x616 & ~x625 & ~x638 & ~x670 & ~x691 & ~x750 & ~x751 & ~x756;
assign c6154 =  x462 &  x495 &  x522 &  x547 &  x575 & ~x8 & ~x14 & ~x66 & ~x90 & ~x173 & ~x186 & ~x214 & ~x506 & ~x588 & ~x644 & ~x677 & ~x705 & ~x707 & ~x756 & ~x761;
assign c6156 =  x573 & ~x1 & ~x10 & ~x11 & ~x17 & ~x19 & ~x24 & ~x29 & ~x32 & ~x33 & ~x37 & ~x40 & ~x44 & ~x53 & ~x55 & ~x61 & ~x65 & ~x69 & ~x79 & ~x87 & ~x88 & ~x90 & ~x108 & ~x109 & ~x112 & ~x115 & ~x119 & ~x123 & ~x135 & ~x138 & ~x142 & ~x144 & ~x164 & ~x167 & ~x168 & ~x170 & ~x190 & ~x199 & ~x200 & ~x201 & ~x202 & ~x215 & ~x216 & ~x219 & ~x220 & ~x221 & ~x222 & ~x224 & ~x226 & ~x243 & ~x246 & ~x252 & ~x254 & ~x259 & ~x269 & ~x303 & ~x305 & ~x306 & ~x313 & ~x324 & ~x333 & ~x338 & ~x361 & ~x364 & ~x367 & ~x368 & ~x378 & ~x392 & ~x395 & ~x396 & ~x417 & ~x449 & ~x450 & ~x477 & ~x479 & ~x505 & ~x507 & ~x533 & ~x535 & ~x559 & ~x590 & ~x592 & ~x593 & ~x612 & ~x615 & ~x617 & ~x619 & ~x639 & ~x642 & ~x645 & ~x647 & ~x648 & ~x650 & ~x655 & ~x657 & ~x661 & ~x662 & ~x663 & ~x665 & ~x671 & ~x674 & ~x675 & ~x681 & ~x685 & ~x686 & ~x690 & ~x691 & ~x692 & ~x693 & ~x695 & ~x699 & ~x700 & ~x701 & ~x703 & ~x705 & ~x710 & ~x712 & ~x714 & ~x715 & ~x719 & ~x722 & ~x725 & ~x732 & ~x733 & ~x735 & ~x736 & ~x737 & ~x739 & ~x740 & ~x741 & ~x744 & ~x745 & ~x747 & ~x752 & ~x754 & ~x755 & ~x757 & ~x759 & ~x763 & ~x764 & ~x769;
assign c6158 =  x267 &  x321 & ~x7 & ~x10 & ~x33 & ~x52 & ~x54 & ~x63 & ~x70 & ~x71 & ~x96 & ~x97 & ~x110 & ~x117 & ~x121 & ~x122 & ~x125 & ~x126 & ~x142 & ~x144 & ~x145 & ~x153 & ~x177 & ~x181 & ~x190 & ~x199 & ~x202 & ~x218 & ~x222 & ~x227 & ~x236 & ~x245 & ~x249 & ~x263 & ~x271 & ~x272 & ~x275 & ~x276 & ~x280 & ~x289 & ~x298 & ~x305 & ~x308 & ~x313 & ~x324 & ~x338 & ~x365 & ~x368 & ~x391 & ~x393 & ~x418 & ~x423 & ~x446 & ~x504 & ~x530 & ~x557 & ~x559 & ~x562 & ~x563 & ~x583 & ~x584 & ~x587 & ~x609 & ~x615 & ~x631 & ~x632 & ~x639 & ~x657 & ~x680 & ~x689 & ~x692 & ~x703 & ~x716 & ~x722 & ~x729 & ~x732 & ~x735 & ~x739 & ~x762 & ~x764 & ~x767 & ~x773 & ~x776 & ~x778;
assign c6160 =  x407 & ~x137 & ~x189 & ~x214 & ~x240 & ~x268 & ~x405 & ~x669 & ~x759;
assign c6162 =  x574 & ~x47 & ~x60 & ~x61 & ~x76 & ~x78 & ~x89 & ~x119 & ~x143 & ~x144 & ~x159 & ~x160 & ~x163 & ~x190 & ~x213 & ~x217 & ~x228 & ~x229 & ~x248 & ~x257 & ~x339 & ~x362 & ~x418 & ~x502 & ~x508 & ~x557 & ~x560 & ~x619 & ~x624 & ~x627 & ~x656 & ~x662 & ~x663 & ~x673 & ~x674 & ~x677 & ~x686 & ~x718 & ~x722 & ~x738 & ~x743 & ~x770;
assign c6164 =  x357 &  x399 & ~x9 & ~x16 & ~x19 & ~x21 & ~x24 & ~x30 & ~x32 & ~x34 & ~x40 & ~x41 & ~x46 & ~x47 & ~x48 & ~x49 & ~x53 & ~x54 & ~x58 & ~x61 & ~x62 & ~x84 & ~x87 & ~x110 & ~x111 & ~x112 & ~x114 & ~x135 & ~x137 & ~x142 & ~x143 & ~x169 & ~x194 & ~x195 & ~x216 & ~x218 & ~x221 & ~x222 & ~x223 & ~x242 & ~x243 & ~x248 & ~x249 & ~x250 & ~x252 & ~x256 & ~x280 & ~x305 & ~x306 & ~x309 & ~x336 & ~x338 & ~x339 & ~x362 & ~x363 & ~x367 & ~x391 & ~x418 & ~x419 & ~x424 & ~x446 & ~x448 & ~x451 & ~x452 & ~x474 & ~x475 & ~x476 & ~x479 & ~x505 & ~x534 & ~x586 & ~x589 & ~x591 & ~x614 & ~x617 & ~x619 & ~x621 & ~x636 & ~x640 & ~x641 & ~x643 & ~x647 & ~x656 & ~x658 & ~x659 & ~x663 & ~x665 & ~x668 & ~x671 & ~x676 & ~x681 & ~x682 & ~x686 & ~x690 & ~x691 & ~x695 & ~x697 & ~x698 & ~x699 & ~x700 & ~x701 & ~x703 & ~x706 & ~x710 & ~x711 & ~x716 & ~x719 & ~x722 & ~x724 & ~x725 & ~x727 & ~x732 & ~x733 & ~x738 & ~x740 & ~x743 & ~x753 & ~x755 & ~x762 & ~x763 & ~x764 & ~x765 & ~x766 & ~x767 & ~x781 & ~x782;
assign c6166 =  x404 &  x432 &  x486 &  x514 &  x574 & ~x44 & ~x72 & ~x99 & ~x127 & ~x152 & ~x154 & ~x172 & ~x181 & ~x236 & ~x339 & ~x395 & ~x419 & ~x422 & ~x501 & ~x534 & ~x561 & ~x642 & ~x652 & ~x706;
assign c6168 =  x156 &  x236 &  x263 &  x318 &  x373 &  x401 &  x429 &  x457 &  x629 & ~x0 & ~x3 & ~x5 & ~x11 & ~x12 & ~x15 & ~x21 & ~x22 & ~x29 & ~x31 & ~x32 & ~x36 & ~x39 & ~x45 & ~x52 & ~x54 & ~x57 & ~x60 & ~x61 & ~x63 & ~x65 & ~x69 & ~x70 & ~x71 & ~x72 & ~x76 & ~x77 & ~x78 & ~x79 & ~x84 & ~x88 & ~x90 & ~x95 & ~x96 & ~x97 & ~x99 & ~x106 & ~x108 & ~x114 & ~x121 & ~x123 & ~x134 & ~x135 & ~x139 & ~x140 & ~x143 & ~x149 & ~x150 & ~x168 & ~x169 & ~x170 & ~x171 & ~x173 & ~x174 & ~x175 & ~x193 & ~x196 & ~x198 & ~x199 & ~x201 & ~x202 & ~x220 & ~x222 & ~x224 & ~x227 & ~x228 & ~x249 & ~x252 & ~x253 & ~x255 & ~x256 & ~x257 & ~x259 & ~x275 & ~x278 & ~x281 & ~x283 & ~x286 & ~x298 & ~x299 & ~x300 & ~x301 & ~x303 & ~x304 & ~x306 & ~x311 & ~x312 & ~x329 & ~x330 & ~x333 & ~x334 & ~x335 & ~x339 & ~x340 & ~x342 & ~x358 & ~x359 & ~x360 & ~x363 & ~x365 & ~x386 & ~x389 & ~x390 & ~x417 & ~x418 & ~x419 & ~x450 & ~x477 & ~x504 & ~x506 & ~x507 & ~x508 & ~x532 & ~x533 & ~x534 & ~x536 & ~x555 & ~x556 & ~x558 & ~x584 & ~x585 & ~x586 & ~x587 & ~x589 & ~x612 & ~x613 & ~x614 & ~x616 & ~x617 & ~x618 & ~x621 & ~x641 & ~x644 & ~x646 & ~x648 & ~x650 & ~x652 & ~x653 & ~x668 & ~x684 & ~x688 & ~x694 & ~x695 & ~x697 & ~x698 & ~x705 & ~x712 & ~x719 & ~x720 & ~x721 & ~x724 & ~x729 & ~x731 & ~x736 & ~x737 & ~x738 & ~x741 & ~x746 & ~x747 & ~x748 & ~x749 & ~x751 & ~x754 & ~x755 & ~x756 & ~x762 & ~x766 & ~x768 & ~x770 & ~x780 & ~x783;
assign c6170 =  x573 & ~x10 & ~x13 & ~x17 & ~x18 & ~x31 & ~x33 & ~x44 & ~x66 & ~x77 & ~x83 & ~x106 & ~x120 & ~x135 & ~x147 & ~x148 & ~x170 & ~x173 & ~x196 & ~x218 & ~x223 & ~x229 & ~x246 & ~x247 & ~x254 & ~x267 & ~x270 & ~x275 & ~x300 & ~x307 & ~x308 & ~x330 & ~x332 & ~x361 & ~x364 & ~x392 & ~x418 & ~x447 & ~x556 & ~x567 & ~x568 & ~x569 & ~x586 & ~x597 & ~x598 & ~x627 & ~x639 & ~x669 & ~x684 & ~x686 & ~x692 & ~x693 & ~x694 & ~x696 & ~x724 & ~x731 & ~x737 & ~x742 & ~x747 & ~x757 & ~x781 & ~x782 & ~x783;
assign c6172 =  x590;
assign c6174 =  x457 &  x631 & ~x0 & ~x1 & ~x3 & ~x4 & ~x5 & ~x7 & ~x8 & ~x10 & ~x11 & ~x16 & ~x17 & ~x19 & ~x27 & ~x29 & ~x35 & ~x37 & ~x40 & ~x41 & ~x42 & ~x43 & ~x48 & ~x54 & ~x57 & ~x63 & ~x65 & ~x66 & ~x69 & ~x70 & ~x77 & ~x79 & ~x80 & ~x81 & ~x88 & ~x90 & ~x105 & ~x106 & ~x107 & ~x109 & ~x112 & ~x115 & ~x116 & ~x117 & ~x119 & ~x138 & ~x143 & ~x144 & ~x147 & ~x148 & ~x149 & ~x167 & ~x168 & ~x170 & ~x173 & ~x195 & ~x199 & ~x200 & ~x202 & ~x225 & ~x227 & ~x228 & ~x231 & ~x240 & ~x256 & ~x268 & ~x270 & ~x279 & ~x283 & ~x295 & ~x297 & ~x299 & ~x302 & ~x307 & ~x308 & ~x309 & ~x312 & ~x327 & ~x330 & ~x341 & ~x359 & ~x360 & ~x365 & ~x368 & ~x369 & ~x389 & ~x392 & ~x394 & ~x396 & ~x418 & ~x422 & ~x446 & ~x449 & ~x450 & ~x451 & ~x452 & ~x474 & ~x475 & ~x476 & ~x478 & ~x480 & ~x505 & ~x507 & ~x508 & ~x509 & ~x529 & ~x534 & ~x535 & ~x537 & ~x558 & ~x560 & ~x562 & ~x563 & ~x565 & ~x588 & ~x589 & ~x592 & ~x613 & ~x616 & ~x617 & ~x640 & ~x641 & ~x643 & ~x653 & ~x666 & ~x669 & ~x670 & ~x671 & ~x674 & ~x675 & ~x676 & ~x678 & ~x681 & ~x682 & ~x683 & ~x684 & ~x685 & ~x689 & ~x691 & ~x693 & ~x697 & ~x699 & ~x701 & ~x704 & ~x705 & ~x706 & ~x719 & ~x722 & ~x724 & ~x725 & ~x726 & ~x729 & ~x732 & ~x733 & ~x735 & ~x740 & ~x741 & ~x743 & ~x744 & ~x746 & ~x750 & ~x751 & ~x754 & ~x755 & ~x756 & ~x761 & ~x763 & ~x764 & ~x765 & ~x766 & ~x767 & ~x768 & ~x770 & ~x772 & ~x773 & ~x774 & ~x776 & ~x778 & ~x780 & ~x782;
assign c6176 =  x573 & ~x10 & ~x19 & ~x32 & ~x34 & ~x35 & ~x38 & ~x45 & ~x50 & ~x91 & ~x185 & ~x197 & ~x198 & ~x201 & ~x228 & ~x238 & ~x239 & ~x285 & ~x292 & ~x305 & ~x531 & ~x585 & ~x593 & ~x644 & ~x663 & ~x668 & ~x688 & ~x692 & ~x723 & ~x724 & ~x739 & ~x748 & ~x755 & ~x771;
assign c6178 =  x102 &  x292 & ~x215;
assign c6180 =  x733;
assign c6182 =  x347 &  x374 &  x402 &  x457 &  x599 & ~x1 & ~x2 & ~x5 & ~x6 & ~x17 & ~x21 & ~x24 & ~x25 & ~x28 & ~x31 & ~x33 & ~x35 & ~x37 & ~x38 & ~x41 & ~x42 & ~x49 & ~x52 & ~x56 & ~x57 & ~x59 & ~x60 & ~x61 & ~x62 & ~x65 & ~x79 & ~x82 & ~x94 & ~x96 & ~x97 & ~x107 & ~x115 & ~x117 & ~x118 & ~x120 & ~x122 & ~x123 & ~x124 & ~x125 & ~x136 & ~x140 & ~x144 & ~x145 & ~x146 & ~x151 & ~x152 & ~x165 & ~x167 & ~x168 & ~x171 & ~x174 & ~x177 & ~x192 & ~x196 & ~x201 & ~x206 & ~x219 & ~x226 & ~x229 & ~x231 & ~x247 & ~x249 & ~x251 & ~x254 & ~x255 & ~x257 & ~x260 & ~x261 & ~x270 & ~x271 & ~x272 & ~x275 & ~x276 & ~x277 & ~x280 & ~x282 & ~x283 & ~x284 & ~x288 & ~x301 & ~x303 & ~x305 & ~x306 & ~x307 & ~x308 & ~x312 & ~x315 & ~x316 & ~x330 & ~x332 & ~x335 & ~x337 & ~x342 & ~x362 & ~x363 & ~x366 & ~x368 & ~x369 & ~x371 & ~x392 & ~x393 & ~x394 & ~x398 & ~x416 & ~x418 & ~x419 & ~x421 & ~x424 & ~x425 & ~x443 & ~x444 & ~x449 & ~x450 & ~x451 & ~x453 & ~x471 & ~x472 & ~x473 & ~x474 & ~x499 & ~x500 & ~x503 & ~x505 & ~x525 & ~x526 & ~x528 & ~x529 & ~x530 & ~x531 & ~x534 & ~x553 & ~x556 & ~x558 & ~x560 & ~x562 & ~x564 & ~x584 & ~x587 & ~x588 & ~x589 & ~x590 & ~x593 & ~x608 & ~x609 & ~x612 & ~x613 & ~x621 & ~x638 & ~x640 & ~x646 & ~x648 & ~x649 & ~x651 & ~x652 & ~x663 & ~x664 & ~x666 & ~x673 & ~x677 & ~x678 & ~x679 & ~x680 & ~x682 & ~x683 & ~x688 & ~x692 & ~x694 & ~x698 & ~x701 & ~x702 & ~x713 & ~x717 & ~x718 & ~x721 & ~x723 & ~x724 & ~x725 & ~x733 & ~x735 & ~x737 & ~x740 & ~x742 & ~x745 & ~x749 & ~x750 & ~x755 & ~x759 & ~x762 & ~x763 & ~x764 & ~x770 & ~x772 & ~x774 & ~x775 & ~x776 & ~x781;
assign c6184 = ~x3 & ~x4 & ~x7 & ~x12 & ~x13 & ~x15 & ~x17 & ~x18 & ~x20 & ~x21 & ~x31 & ~x40 & ~x42 & ~x47 & ~x48 & ~x53 & ~x55 & ~x62 & ~x69 & ~x80 & ~x85 & ~x91 & ~x96 & ~x97 & ~x106 & ~x108 & ~x112 & ~x113 & ~x115 & ~x120 & ~x121 & ~x134 & ~x135 & ~x141 & ~x145 & ~x147 & ~x151 & ~x161 & ~x164 & ~x168 & ~x170 & ~x172 & ~x174 & ~x175 & ~x180 & ~x187 & ~x188 & ~x193 & ~x202 & ~x205 & ~x207 & ~x221 & ~x228 & ~x233 & ~x242 & ~x246 & ~x247 & ~x248 & ~x251 & ~x254 & ~x257 & ~x261 & ~x262 & ~x276 & ~x281 & ~x288 & ~x306 & ~x310 & ~x316 & ~x331 & ~x334 & ~x336 & ~x338 & ~x339 & ~x340 & ~x359 & ~x370 & ~x387 & ~x388 & ~x395 & ~x397 & ~x417 & ~x419 & ~x421 & ~x423 & ~x443 & ~x444 & ~x446 & ~x450 & ~x473 & ~x479 & ~x499 & ~x502 & ~x503 & ~x526 & ~x527 & ~x534 & ~x553 & ~x554 & ~x560 & ~x561 & ~x563 & ~x587 & ~x589 & ~x590 & ~x592 & ~x594 & ~x606 & ~x607 & ~x612 & ~x621 & ~x633 & ~x636 & ~x638 & ~x639 & ~x640 & ~x646 & ~x648 & ~x649 & ~x651 & ~x652 & ~x653 & ~x654 & ~x655 & ~x656 & ~x657 & ~x658 & ~x660 & ~x661 & ~x662 & ~x664 & ~x668 & ~x674 & ~x678 & ~x683 & ~x685 & ~x686 & ~x689 & ~x690 & ~x700 & ~x701 & ~x702 & ~x705 & ~x708 & ~x710 & ~x712 & ~x715 & ~x716 & ~x720 & ~x721 & ~x723 & ~x725 & ~x727 & ~x729 & ~x736 & ~x740 & ~x741 & ~x744 & ~x747 & ~x756 & ~x763 & ~x764 & ~x765 & ~x770 & ~x776 & ~x778;
assign c6186 =  x110;
assign c6188 =  x517 & ~x17 & ~x84 & ~x141 & ~x168 & ~x190 & ~x200 & ~x228 & ~x267 & ~x278 & ~x420 & ~x424 & ~x507 & ~x532 & ~x593 & ~x612 & ~x617 & ~x630 & ~x632 & ~x660 & ~x746 & ~x754 & ~x758;
assign c6190 =  x353 &  x379 &  x385 & ~x22 & ~x30 & ~x84 & ~x188 & ~x215 & ~x217 & ~x218 & ~x248 & ~x256 & ~x340 & ~x480 & ~x643 & ~x651 & ~x658 & ~x659 & ~x661 & ~x663 & ~x664 & ~x675 & ~x725 & ~x730;
assign c6192 =  x320 &  x348 &  x402 &  x459 &  x600 & ~x6 & ~x8 & ~x20 & ~x21 & ~x32 & ~x40 & ~x48 & ~x52 & ~x53 & ~x60 & ~x62 & ~x74 & ~x87 & ~x92 & ~x111 & ~x138 & ~x151 & ~x167 & ~x168 & ~x175 & ~x179 & ~x190 & ~x191 & ~x194 & ~x204 & ~x219 & ~x223 & ~x224 & ~x232 & ~x234 & ~x246 & ~x253 & ~x254 & ~x255 & ~x270 & ~x286 & ~x289 & ~x302 & ~x303 & ~x308 & ~x311 & ~x334 & ~x338 & ~x396 & ~x417 & ~x424 & ~x451 & ~x477 & ~x499 & ~x501 & ~x505 & ~x506 & ~x508 & ~x535 & ~x552 & ~x557 & ~x558 & ~x563 & ~x564 & ~x593 & ~x621 & ~x640 & ~x663 & ~x664 & ~x667 & ~x671 & ~x677 & ~x725 & ~x730 & ~x740 & ~x744 & ~x748 & ~x762;
assign c6194 =  x99 & ~x25 & ~x103 & ~x121 & ~x130 & ~x132 & ~x158 & ~x172 & ~x186 & ~x187 & ~x213 & ~x230 & ~x242 & ~x248 & ~x284 & ~x695;
assign c6196 =  x346 &  x373 &  x401 &  x428 &  x455 &  x483 &  x511 &  x539 &  x544 &  x597 &  x599 & ~x26 & ~x42 & ~x72 & ~x125 & ~x126 & ~x153 & ~x275 & ~x305 & ~x332 & ~x366 & ~x449 & ~x502 & ~x508 & ~x558 & ~x561 & ~x586 & ~x593 & ~x644 & ~x650 & ~x662 & ~x698 & ~x711 & ~x777;
assign c6198 =  x458 &  x486 &  x514 &  x599 & ~x1 & ~x4 & ~x5 & ~x7 & ~x8 & ~x10 & ~x12 & ~x18 & ~x23 & ~x26 & ~x32 & ~x33 & ~x34 & ~x36 & ~x38 & ~x41 & ~x42 & ~x43 & ~x44 & ~x45 & ~x46 & ~x48 & ~x53 & ~x55 & ~x56 & ~x57 & ~x58 & ~x60 & ~x62 & ~x67 & ~x69 & ~x76 & ~x80 & ~x83 & ~x84 & ~x85 & ~x87 & ~x89 & ~x91 & ~x93 & ~x94 & ~x96 & ~x97 & ~x107 & ~x109 & ~x111 & ~x112 & ~x114 & ~x115 & ~x116 & ~x118 & ~x119 & ~x120 & ~x121 & ~x122 & ~x123 & ~x136 & ~x137 & ~x139 & ~x141 & ~x142 & ~x148 & ~x149 & ~x150 & ~x162 & ~x163 & ~x166 & ~x167 & ~x168 & ~x169 & ~x172 & ~x173 & ~x178 & ~x191 & ~x192 & ~x193 & ~x195 & ~x196 & ~x198 & ~x199 & ~x200 & ~x204 & ~x220 & ~x223 & ~x224 & ~x226 & ~x232 & ~x248 & ~x249 & ~x252 & ~x253 & ~x256 & ~x259 & ~x260 & ~x275 & ~x277 & ~x281 & ~x282 & ~x284 & ~x285 & ~x287 & ~x297 & ~x302 & ~x303 & ~x306 & ~x307 & ~x309 & ~x310 & ~x315 & ~x327 & ~x330 & ~x332 & ~x335 & ~x336 & ~x340 & ~x341 & ~x356 & ~x357 & ~x358 & ~x359 & ~x368 & ~x371 & ~x386 & ~x388 & ~x390 & ~x391 & ~x393 & ~x395 & ~x396 & ~x415 & ~x418 & ~x426 & ~x443 & ~x446 & ~x447 & ~x448 & ~x450 & ~x451 & ~x454 & ~x471 & ~x472 & ~x477 & ~x478 & ~x479 & ~x480 & ~x481 & ~x482 & ~x483 & ~x498 & ~x500 & ~x502 & ~x504 & ~x505 & ~x509 & ~x510 & ~x511 & ~x527 & ~x530 & ~x531 & ~x532 & ~x533 & ~x534 & ~x535 & ~x537 & ~x539 & ~x556 & ~x558 & ~x560 & ~x561 & ~x562 & ~x564 & ~x566 & ~x567 & ~x582 & ~x584 & ~x586 & ~x587 & ~x592 & ~x594 & ~x595 & ~x596 & ~x616 & ~x617 & ~x620 & ~x623 & ~x624 & ~x637 & ~x638 & ~x640 & ~x642 & ~x644 & ~x645 & ~x650 & ~x652 & ~x653 & ~x665 & ~x667 & ~x668 & ~x670 & ~x671 & ~x672 & ~x673 & ~x674 & ~x675 & ~x677 & ~x678 & ~x679 & ~x681 & ~x690 & ~x691 & ~x692 & ~x693 & ~x695 & ~x697 & ~x699 & ~x706 & ~x707 & ~x711 & ~x715 & ~x716 & ~x717 & ~x718 & ~x719 & ~x720 & ~x721 & ~x722 & ~x724 & ~x728 & ~x729 & ~x730 & ~x731 & ~x732 & ~x733 & ~x735 & ~x737 & ~x738 & ~x740 & ~x741 & ~x742 & ~x744 & ~x745 & ~x746 & ~x748 & ~x750 & ~x752 & ~x754 & ~x755 & ~x757 & ~x758 & ~x760 & ~x761 & ~x762 & ~x767 & ~x768 & ~x769 & ~x770 & ~x771 & ~x772 & ~x776 & ~x777 & ~x778 & ~x781 & ~x782 & ~x783;
assign c6200 =  x321 &  x349 &  x404 & ~x2 & ~x4 & ~x12 & ~x19 & ~x21 & ~x25 & ~x34 & ~x51 & ~x54 & ~x57 & ~x65 & ~x66 & ~x85 & ~x91 & ~x93 & ~x110 & ~x126 & ~x138 & ~x142 & ~x143 & ~x151 & ~x153 & ~x169 & ~x176 & ~x179 & ~x231 & ~x271 & ~x277 & ~x283 & ~x285 & ~x301 & ~x302 & ~x304 & ~x328 & ~x354 & ~x361 & ~x385 & ~x390 & ~x397 & ~x398 & ~x413 & ~x417 & ~x422 & ~x477 & ~x496 & ~x502 & ~x503 & ~x508 & ~x509 & ~x525 & ~x537 & ~x555 & ~x557 & ~x561 & ~x563 & ~x581 & ~x608 & ~x610 & ~x613 & ~x639 & ~x662 & ~x672 & ~x673 & ~x680 & ~x681 & ~x682 & ~x703 & ~x715 & ~x717 & ~x722 & ~x725 & ~x731 & ~x735 & ~x740 & ~x742 & ~x757 & ~x771;
assign c6202 =  x430 &  x486 &  x514 &  x515 &  x543 &  x572 & ~x0 & ~x4 & ~x7 & ~x8 & ~x9 & ~x11 & ~x14 & ~x18 & ~x21 & ~x25 & ~x26 & ~x27 & ~x28 & ~x29 & ~x31 & ~x32 & ~x37 & ~x39 & ~x40 & ~x43 & ~x45 & ~x49 & ~x52 & ~x53 & ~x54 & ~x58 & ~x59 & ~x68 & ~x71 & ~x72 & ~x74 & ~x76 & ~x80 & ~x82 & ~x83 & ~x86 & ~x93 & ~x94 & ~x97 & ~x102 & ~x105 & ~x107 & ~x108 & ~x110 & ~x111 & ~x112 & ~x113 & ~x115 & ~x117 & ~x120 & ~x138 & ~x141 & ~x144 & ~x146 & ~x147 & ~x148 & ~x163 & ~x165 & ~x170 & ~x174 & ~x196 & ~x198 & ~x199 & ~x201 & ~x227 & ~x247 & ~x248 & ~x249 & ~x251 & ~x254 & ~x256 & ~x275 & ~x280 & ~x283 & ~x285 & ~x287 & ~x303 & ~x305 & ~x306 & ~x307 & ~x311 & ~x312 & ~x313 & ~x331 & ~x332 & ~x337 & ~x338 & ~x343 & ~x360 & ~x361 & ~x364 & ~x365 & ~x368 & ~x371 & ~x386 & ~x387 & ~x388 & ~x389 & ~x390 & ~x391 & ~x392 & ~x394 & ~x398 & ~x420 & ~x422 & ~x426 & ~x427 & ~x443 & ~x444 & ~x448 & ~x449 & ~x450 & ~x454 & ~x471 & ~x472 & ~x473 & ~x475 & ~x479 & ~x498 & ~x501 & ~x502 & ~x503 & ~x506 & ~x507 & ~x511 & ~x529 & ~x531 & ~x534 & ~x537 & ~x538 & ~x539 & ~x555 & ~x557 & ~x559 & ~x563 & ~x564 & ~x565 & ~x567 & ~x581 & ~x582 & ~x583 & ~x585 & ~x587 & ~x588 & ~x589 & ~x594 & ~x596 & ~x615 & ~x617 & ~x619 & ~x620 & ~x622 & ~x625 & ~x636 & ~x637 & ~x638 & ~x644 & ~x645 & ~x651 & ~x662 & ~x665 & ~x666 & ~x667 & ~x668 & ~x669 & ~x672 & ~x675 & ~x676 & ~x677 & ~x678 & ~x679 & ~x682 & ~x688 & ~x691 & ~x699 & ~x701 & ~x707 & ~x709 & ~x714 & ~x715 & ~x722 & ~x723 & ~x726 & ~x727 & ~x730 & ~x732 & ~x733 & ~x736 & ~x744 & ~x749 & ~x750 & ~x752 & ~x754 & ~x757 & ~x758 & ~x759 & ~x760 & ~x763 & ~x765 & ~x770 & ~x773 & ~x774 & ~x775 & ~x777 & ~x778 & ~x779;
assign c6204 =  x578 & ~x9 & ~x77 & ~x78 & ~x144 & ~x155 & ~x236 & ~x277 & ~x390 & ~x536 & ~x559 & ~x565 & ~x651 & ~x661 & ~x665 & ~x739 & ~x752;
assign c6206 = ~x0 & ~x1 & ~x15 & ~x17 & ~x41 & ~x51 & ~x75 & ~x142 & ~x163 & ~x167 & ~x192 & ~x194 & ~x195 & ~x196 & ~x200 & ~x222 & ~x238 & ~x240 & ~x242 & ~x244 & ~x248 & ~x249 & ~x253 & ~x254 & ~x266 & ~x293 & ~x339 & ~x340 & ~x347 & ~x422 & ~x424 & ~x479 & ~x505 & ~x531 & ~x537 & ~x560 & ~x562 & ~x564 & ~x588 & ~x590 & ~x612 & ~x622 & ~x654 & ~x690 & ~x702 & ~x708 & ~x722 & ~x743 & ~x748 & ~x778;
assign c6208 =  x345 &  x428 &  x541 &  x578 &  x599 &  x600 &  x601 &  x602 & ~x8 & ~x10 & ~x13 & ~x16 & ~x19 & ~x26 & ~x39 & ~x46 & ~x52 & ~x54 & ~x55 & ~x56 & ~x64 & ~x67 & ~x79 & ~x82 & ~x106 & ~x107 & ~x114 & ~x115 & ~x116 & ~x119 & ~x138 & ~x139 & ~x143 & ~x145 & ~x164 & ~x165 & ~x192 & ~x193 & ~x218 & ~x223 & ~x224 & ~x227 & ~x228 & ~x229 & ~x230 & ~x243 & ~x246 & ~x251 & ~x274 & ~x278 & ~x282 & ~x285 & ~x303 & ~x308 & ~x310 & ~x331 & ~x336 & ~x338 & ~x339 & ~x360 & ~x361 & ~x392 & ~x393 & ~x394 & ~x421 & ~x422 & ~x446 & ~x477 & ~x479 & ~x503 & ~x530 & ~x563 & ~x564 & ~x583 & ~x588 & ~x589 & ~x614 & ~x616 & ~x636 & ~x640 & ~x641 & ~x648 & ~x652 & ~x653 & ~x654 & ~x663 & ~x673 & ~x674 & ~x675 & ~x679 & ~x681 & ~x685 & ~x687 & ~x694 & ~x695 & ~x697 & ~x698 & ~x701 & ~x706 & ~x709 & ~x713 & ~x717 & ~x721 & ~x722 & ~x724 & ~x729 & ~x730 & ~x731 & ~x734 & ~x740 & ~x741 & ~x743 & ~x747 & ~x754 & ~x757 & ~x760 & ~x762 & ~x768 & ~x773 & ~x776 & ~x780 & ~x783;
assign c6210 =  x720;
assign c6212 =  x209 & ~x212 & ~x268;
assign c6214 = ~x182 & ~x214 & ~x237 & ~x465 & ~x626 & ~x755 & ~x779;
assign c6216 =  x156 &  x600 & ~x0 & ~x8 & ~x15 & ~x16 & ~x17 & ~x20 & ~x24 & ~x27 & ~x28 & ~x30 & ~x31 & ~x32 & ~x33 & ~x37 & ~x38 & ~x41 & ~x44 & ~x45 & ~x49 & ~x58 & ~x63 & ~x65 & ~x66 & ~x69 & ~x70 & ~x71 & ~x77 & ~x82 & ~x87 & ~x89 & ~x91 & ~x93 & ~x95 & ~x96 & ~x97 & ~x104 & ~x107 & ~x109 & ~x110 & ~x111 & ~x118 & ~x123 & ~x124 & ~x125 & ~x135 & ~x136 & ~x139 & ~x140 & ~x145 & ~x146 & ~x149 & ~x150 & ~x151 & ~x167 & ~x171 & ~x172 & ~x173 & ~x176 & ~x177 & ~x178 & ~x193 & ~x194 & ~x205 & ~x222 & ~x227 & ~x229 & ~x232 & ~x251 & ~x252 & ~x254 & ~x257 & ~x258 & ~x259 & ~x269 & ~x270 & ~x276 & ~x281 & ~x296 & ~x298 & ~x302 & ~x304 & ~x310 & ~x312 & ~x313 & ~x314 & ~x324 & ~x325 & ~x326 & ~x327 & ~x328 & ~x331 & ~x332 & ~x334 & ~x336 & ~x340 & ~x342 & ~x354 & ~x355 & ~x360 & ~x365 & ~x367 & ~x369 & ~x387 & ~x389 & ~x390 & ~x393 & ~x397 & ~x418 & ~x420 & ~x421 & ~x422 & ~x423 & ~x442 & ~x446 & ~x448 & ~x449 & ~x450 & ~x476 & ~x478 & ~x501 & ~x503 & ~x507 & ~x530 & ~x558 & ~x560 & ~x564 & ~x565 & ~x566 & ~x584 & ~x586 & ~x591 & ~x592 & ~x612 & ~x614 & ~x615 & ~x616 & ~x617 & ~x618 & ~x622 & ~x623 & ~x624 & ~x625 & ~x626 & ~x647 & ~x654 & ~x667 & ~x673 & ~x681 & ~x684 & ~x689 & ~x690 & ~x695 & ~x696 & ~x701 & ~x702 & ~x703 & ~x704 & ~x707 & ~x710 & ~x711 & ~x714 & ~x717 & ~x722 & ~x724 & ~x725 & ~x726 & ~x731 & ~x733 & ~x735 & ~x738 & ~x741 & ~x752 & ~x754 & ~x758 & ~x760 & ~x762 & ~x763 & ~x764 & ~x765 & ~x766 & ~x768 & ~x770 & ~x774 & ~x777 & ~x780;
assign c6218 =  x126 &  x207 &  x570 & ~x1 & ~x14 & ~x21 & ~x29 & ~x33 & ~x56 & ~x60 & ~x65 & ~x79 & ~x132 & ~x134 & ~x135 & ~x170 & ~x173 & ~x175 & ~x192 & ~x222 & ~x230 & ~x248 & ~x267 & ~x271 & ~x273 & ~x294 & ~x305 & ~x311 & ~x312 & ~x333 & ~x334 & ~x393 & ~x418 & ~x419 & ~x421 & ~x424 & ~x478 & ~x479 & ~x530 & ~x537 & ~x562 & ~x566 & ~x584 & ~x595 & ~x611 & ~x653 & ~x666 & ~x683 & ~x685 & ~x692 & ~x707 & ~x719 & ~x722 & ~x742 & ~x762 & ~x767 & ~x778;
assign c6220 =  x140;
assign c6222 =  x159 &  x429 &  x457 &  x485 &  x513 &  x569 & ~x0 & ~x1 & ~x2 & ~x3 & ~x5 & ~x10 & ~x14 & ~x15 & ~x17 & ~x19 & ~x23 & ~x24 & ~x25 & ~x28 & ~x31 & ~x32 & ~x34 & ~x38 & ~x43 & ~x45 & ~x46 & ~x47 & ~x50 & ~x56 & ~x57 & ~x62 & ~x66 & ~x72 & ~x73 & ~x76 & ~x77 & ~x81 & ~x82 & ~x83 & ~x87 & ~x93 & ~x94 & ~x96 & ~x97 & ~x99 & ~x101 & ~x109 & ~x110 & ~x112 & ~x113 & ~x117 & ~x119 & ~x122 & ~x123 & ~x124 & ~x137 & ~x139 & ~x140 & ~x141 & ~x142 & ~x143 & ~x144 & ~x147 & ~x150 & ~x167 & ~x169 & ~x174 & ~x177 & ~x178 & ~x194 & ~x195 & ~x197 & ~x200 & ~x203 & ~x204 & ~x205 & ~x206 & ~x223 & ~x227 & ~x230 & ~x232 & ~x247 & ~x249 & ~x256 & ~x257 & ~x260 & ~x275 & ~x276 & ~x283 & ~x299 & ~x300 & ~x301 & ~x302 & ~x303 & ~x304 & ~x306 & ~x309 & ~x310 & ~x311 & ~x313 & ~x315 & ~x316 & ~x326 & ~x329 & ~x330 & ~x332 & ~x333 & ~x335 & ~x339 & ~x340 & ~x343 & ~x356 & ~x358 & ~x360 & ~x362 & ~x364 & ~x366 & ~x368 & ~x369 & ~x370 & ~x385 & ~x386 & ~x388 & ~x391 & ~x394 & ~x395 & ~x414 & ~x415 & ~x416 & ~x417 & ~x425 & ~x445 & ~x446 & ~x447 & ~x448 & ~x450 & ~x471 & ~x472 & ~x476 & ~x478 & ~x481 & ~x499 & ~x500 & ~x503 & ~x504 & ~x505 & ~x507 & ~x509 & ~x535 & ~x536 & ~x537 & ~x556 & ~x558 & ~x559 & ~x562 & ~x564 & ~x565 & ~x581 & ~x583 & ~x584 & ~x589 & ~x590 & ~x594 & ~x609 & ~x610 & ~x616 & ~x617 & ~x620 & ~x621 & ~x640 & ~x641 & ~x644 & ~x646 & ~x650 & ~x663 & ~x664 & ~x665 & ~x670 & ~x672 & ~x675 & ~x676 & ~x681 & ~x683 & ~x689 & ~x692 & ~x693 & ~x694 & ~x695 & ~x704 & ~x705 & ~x712 & ~x713 & ~x714 & ~x717 & ~x719 & ~x720 & ~x724 & ~x725 & ~x727 & ~x728 & ~x730 & ~x734 & ~x735 & ~x740 & ~x742 & ~x743 & ~x745 & ~x748 & ~x752 & ~x754 & ~x758 & ~x759 & ~x760 & ~x761 & ~x767 & ~x769 & ~x774 & ~x777 & ~x781 & ~x782 & ~x783;
assign c6224 =  x698;
assign c6226 =  x374 &  x457 &  x571 & ~x1 & ~x2 & ~x3 & ~x6 & ~x8 & ~x10 & ~x15 & ~x17 & ~x19 & ~x20 & ~x21 & ~x22 & ~x25 & ~x26 & ~x27 & ~x29 & ~x30 & ~x31 & ~x33 & ~x35 & ~x37 & ~x38 & ~x39 & ~x43 & ~x44 & ~x47 & ~x51 & ~x52 & ~x53 & ~x59 & ~x60 & ~x62 & ~x63 & ~x65 & ~x70 & ~x71 & ~x73 & ~x74 & ~x75 & ~x79 & ~x80 & ~x81 & ~x82 & ~x84 & ~x85 & ~x86 & ~x87 & ~x89 & ~x90 & ~x91 & ~x92 & ~x93 & ~x94 & ~x95 & ~x113 & ~x114 & ~x115 & ~x116 & ~x117 & ~x118 & ~x119 & ~x123 & ~x135 & ~x139 & ~x141 & ~x144 & ~x145 & ~x146 & ~x150 & ~x151 & ~x163 & ~x165 & ~x171 & ~x172 & ~x173 & ~x174 & ~x175 & ~x178 & ~x194 & ~x198 & ~x201 & ~x202 & ~x204 & ~x206 & ~x221 & ~x222 & ~x223 & ~x225 & ~x226 & ~x229 & ~x232 & ~x233 & ~x243 & ~x248 & ~x249 & ~x250 & ~x253 & ~x256 & ~x257 & ~x258 & ~x259 & ~x270 & ~x271 & ~x272 & ~x276 & ~x279 & ~x281 & ~x282 & ~x284 & ~x285 & ~x286 & ~x287 & ~x300 & ~x301 & ~x303 & ~x308 & ~x310 & ~x312 & ~x329 & ~x330 & ~x331 & ~x332 & ~x333 & ~x334 & ~x335 & ~x338 & ~x339 & ~x340 & ~x342 & ~x344 & ~x358 & ~x361 & ~x363 & ~x369 & ~x386 & ~x387 & ~x388 & ~x389 & ~x392 & ~x393 & ~x397 & ~x398 & ~x399 & ~x414 & ~x416 & ~x417 & ~x418 & ~x419 & ~x420 & ~x421 & ~x423 & ~x424 & ~x425 & ~x443 & ~x444 & ~x445 & ~x447 & ~x450 & ~x470 & ~x472 & ~x473 & ~x475 & ~x479 & ~x480 & ~x481 & ~x503 & ~x506 & ~x509 & ~x526 & ~x528 & ~x530 & ~x532 & ~x536 & ~x538 & ~x555 & ~x558 & ~x560 & ~x564 & ~x583 & ~x584 & ~x585 & ~x586 & ~x587 & ~x588 & ~x593 & ~x611 & ~x615 & ~x617 & ~x618 & ~x619 & ~x621 & ~x637 & ~x640 & ~x641 & ~x643 & ~x644 & ~x647 & ~x650 & ~x652 & ~x653 & ~x667 & ~x668 & ~x669 & ~x670 & ~x672 & ~x674 & ~x675 & ~x678 & ~x681 & ~x682 & ~x684 & ~x686 & ~x688 & ~x690 & ~x691 & ~x692 & ~x694 & ~x695 & ~x696 & ~x697 & ~x699 & ~x700 & ~x701 & ~x702 & ~x704 & ~x707 & ~x708 & ~x712 & ~x722 & ~x723 & ~x726 & ~x727 & ~x729 & ~x733 & ~x734 & ~x736 & ~x737 & ~x739 & ~x740 & ~x741 & ~x743 & ~x746 & ~x747 & ~x748 & ~x751 & ~x753 & ~x754 & ~x755 & ~x756 & ~x757 & ~x758 & ~x763 & ~x764 & ~x768 & ~x770 & ~x772 & ~x773 & ~x774 & ~x775 & ~x778 & ~x782 & ~x783;
assign c6228 =  x375 &  x403 &  x431 &  x516 &  x544 & ~x2 & ~x3 & ~x5 & ~x6 & ~x10 & ~x13 & ~x23 & ~x24 & ~x25 & ~x26 & ~x29 & ~x34 & ~x36 & ~x38 & ~x39 & ~x41 & ~x42 & ~x43 & ~x44 & ~x45 & ~x47 & ~x48 & ~x51 & ~x53 & ~x54 & ~x56 & ~x57 & ~x59 & ~x60 & ~x61 & ~x62 & ~x65 & ~x66 & ~x73 & ~x75 & ~x78 & ~x79 & ~x81 & ~x82 & ~x85 & ~x86 & ~x88 & ~x90 & ~x93 & ~x108 & ~x110 & ~x113 & ~x117 & ~x118 & ~x119 & ~x134 & ~x136 & ~x138 & ~x140 & ~x141 & ~x142 & ~x145 & ~x146 & ~x147 & ~x164 & ~x167 & ~x171 & ~x175 & ~x177 & ~x191 & ~x195 & ~x198 & ~x199 & ~x200 & ~x201 & ~x204 & ~x218 & ~x219 & ~x225 & ~x226 & ~x227 & ~x228 & ~x229 & ~x230 & ~x231 & ~x246 & ~x249 & ~x250 & ~x251 & ~x252 & ~x255 & ~x256 & ~x259 & ~x274 & ~x280 & ~x283 & ~x286 & ~x287 & ~x288 & ~x300 & ~x302 & ~x305 & ~x308 & ~x310 & ~x311 & ~x312 & ~x313 & ~x315 & ~x329 & ~x331 & ~x333 & ~x334 & ~x335 & ~x337 & ~x342 & ~x343 & ~x358 & ~x359 & ~x364 & ~x366 & ~x368 & ~x369 & ~x370 & ~x387 & ~x388 & ~x390 & ~x392 & ~x393 & ~x398 & ~x416 & ~x417 & ~x418 & ~x419 & ~x426 & ~x427 & ~x443 & ~x445 & ~x448 & ~x450 & ~x452 & ~x453 & ~x455 & ~x456 & ~x472 & ~x473 & ~x475 & ~x476 & ~x477 & ~x478 & ~x480 & ~x481 & ~x483 & ~x499 & ~x500 & ~x502 & ~x504 & ~x505 & ~x507 & ~x508 & ~x509 & ~x528 & ~x531 & ~x532 & ~x533 & ~x537 & ~x538 & ~x558 & ~x560 & ~x561 & ~x565 & ~x584 & ~x585 & ~x586 & ~x593 & ~x596 & ~x611 & ~x618 & ~x623 & ~x637 & ~x638 & ~x642 & ~x645 & ~x648 & ~x651 & ~x665 & ~x667 & ~x670 & ~x672 & ~x675 & ~x677 & ~x680 & ~x682 & ~x683 & ~x687 & ~x688 & ~x696 & ~x704 & ~x711 & ~x713 & ~x716 & ~x717 & ~x724 & ~x725 & ~x730 & ~x731 & ~x732 & ~x736 & ~x737 & ~x739 & ~x740 & ~x741 & ~x742 & ~x745 & ~x747 & ~x748 & ~x749 & ~x750 & ~x754 & ~x757 & ~x759 & ~x762 & ~x767 & ~x774 & ~x778 & ~x780;
assign c6230 =  x19;
assign c6232 =  x428 &  x468 & ~x0 & ~x4 & ~x5 & ~x7 & ~x8 & ~x9 & ~x21 & ~x27 & ~x33 & ~x38 & ~x39 & ~x46 & ~x54 & ~x60 & ~x62 & ~x65 & ~x66 & ~x67 & ~x78 & ~x91 & ~x92 & ~x110 & ~x116 & ~x118 & ~x119 & ~x122 & ~x123 & ~x141 & ~x143 & ~x145 & ~x164 & ~x167 & ~x168 & ~x169 & ~x175 & ~x201 & ~x219 & ~x220 & ~x229 & ~x231 & ~x241 & ~x246 & ~x248 & ~x249 & ~x251 & ~x256 & ~x269 & ~x271 & ~x279 & ~x281 & ~x301 & ~x312 & ~x331 & ~x337 & ~x341 & ~x361 & ~x366 & ~x394 & ~x397 & ~x415 & ~x418 & ~x419 & ~x444 & ~x446 & ~x472 & ~x474 & ~x478 & ~x480 & ~x501 & ~x507 & ~x530 & ~x532 & ~x533 & ~x536 & ~x537 & ~x557 & ~x558 & ~x561 & ~x562 & ~x565 & ~x584 & ~x587 & ~x591 & ~x593 & ~x613 & ~x618 & ~x623 & ~x624 & ~x640 & ~x641 & ~x642 & ~x644 & ~x646 & ~x647 & ~x649 & ~x671 & ~x678 & ~x680 & ~x681 & ~x684 & ~x692 & ~x693 & ~x696 & ~x706 & ~x708 & ~x710 & ~x711 & ~x713 & ~x716 & ~x719 & ~x720 & ~x721 & ~x722 & ~x728 & ~x736 & ~x745 & ~x756 & ~x762 & ~x764 & ~x772 & ~x774 & ~x777 & ~x782;
assign c6234 =  x517 &  x604 & ~x65 & ~x105 & ~x238 & ~x247 & ~x627 & ~x646 & ~x654 & ~x699;
assign c6236 =  x387 & ~x158 & ~x209;
assign c6238 = ~x0 & ~x2 & ~x3 & ~x4 & ~x6 & ~x7 & ~x9 & ~x10 & ~x11 & ~x12 & ~x13 & ~x14 & ~x16 & ~x17 & ~x18 & ~x19 & ~x20 & ~x21 & ~x22 & ~x23 & ~x24 & ~x26 & ~x28 & ~x29 & ~x30 & ~x33 & ~x34 & ~x36 & ~x37 & ~x41 & ~x42 & ~x43 & ~x44 & ~x45 & ~x49 & ~x50 & ~x51 & ~x52 & ~x53 & ~x54 & ~x55 & ~x56 & ~x57 & ~x59 & ~x60 & ~x61 & ~x62 & ~x64 & ~x65 & ~x68 & ~x69 & ~x75 & ~x77 & ~x78 & ~x79 & ~x80 & ~x82 & ~x85 & ~x86 & ~x87 & ~x89 & ~x90 & ~x91 & ~x92 & ~x95 & ~x105 & ~x106 & ~x107 & ~x108 & ~x109 & ~x110 & ~x111 & ~x113 & ~x114 & ~x115 & ~x118 & ~x122 & ~x123 & ~x134 & ~x136 & ~x139 & ~x140 & ~x142 & ~x143 & ~x145 & ~x146 & ~x148 & ~x149 & ~x163 & ~x166 & ~x167 & ~x172 & ~x173 & ~x175 & ~x176 & ~x177 & ~x178 & ~x189 & ~x190 & ~x191 & ~x192 & ~x193 & ~x194 & ~x195 & ~x196 & ~x197 & ~x200 & ~x201 & ~x202 & ~x203 & ~x204 & ~x205 & ~x206 & ~x216 & ~x217 & ~x219 & ~x220 & ~x221 & ~x224 & ~x225 & ~x226 & ~x227 & ~x229 & ~x231 & ~x232 & ~x234 & ~x242 & ~x243 & ~x244 & ~x245 & ~x246 & ~x249 & ~x250 & ~x251 & ~x252 & ~x253 & ~x256 & ~x257 & ~x259 & ~x261 & ~x274 & ~x276 & ~x281 & ~x282 & ~x288 & ~x289 & ~x304 & ~x305 & ~x307 & ~x309 & ~x310 & ~x315 & ~x332 & ~x333 & ~x339 & ~x341 & ~x342 & ~x343 & ~x344 & ~x360 & ~x361 & ~x362 & ~x364 & ~x365 & ~x366 & ~x368 & ~x369 & ~x388 & ~x389 & ~x390 & ~x391 & ~x392 & ~x393 & ~x396 & ~x398 & ~x415 & ~x418 & ~x420 & ~x423 & ~x424 & ~x425 & ~x426 & ~x447 & ~x448 & ~x449 & ~x451 & ~x452 & ~x473 & ~x474 & ~x475 & ~x476 & ~x480 & ~x481 & ~x500 & ~x502 & ~x505 & ~x507 & ~x508 & ~x527 & ~x528 & ~x529 & ~x531 & ~x534 & ~x535 & ~x537 & ~x554 & ~x555 & ~x556 & ~x558 & ~x559 & ~x560 & ~x563 & ~x564 & ~x582 & ~x583 & ~x587 & ~x590 & ~x592 & ~x607 & ~x610 & ~x612 & ~x614 & ~x615 & ~x616 & ~x617 & ~x618 & ~x620 & ~x635 & ~x636 & ~x637 & ~x639 & ~x642 & ~x647 & ~x648 & ~x651 & ~x652 & ~x656 & ~x657 & ~x658 & ~x659 & ~x660 & ~x661 & ~x662 & ~x663 & ~x664 & ~x667 & ~x668 & ~x669 & ~x670 & ~x671 & ~x672 & ~x674 & ~x675 & ~x677 & ~x680 & ~x683 & ~x684 & ~x685 & ~x686 & ~x688 & ~x691 & ~x693 & ~x695 & ~x697 & ~x698 & ~x700 & ~x701 & ~x704 & ~x705 & ~x707 & ~x708 & ~x709 & ~x710 & ~x711 & ~x712 & ~x713 & ~x714 & ~x715 & ~x716 & ~x717 & ~x718 & ~x719 & ~x720 & ~x721 & ~x722 & ~x723 & ~x724 & ~x725 & ~x728 & ~x736 & ~x737 & ~x738 & ~x741 & ~x744 & ~x747 & ~x748 & ~x749 & ~x751 & ~x752 & ~x754 & ~x755 & ~x756 & ~x759 & ~x762 & ~x763 & ~x764 & ~x765 & ~x771 & ~x772 & ~x773 & ~x775 & ~x777 & ~x780 & ~x781 & ~x782 & ~x783;
assign c6240 =  x574 & ~x39 & ~x54 & ~x94 & ~x161 & ~x186 & ~x238 & ~x282 & ~x368 & ~x392 & ~x480 & ~x651 & ~x655 & ~x662 & ~x686 & ~x694 & ~x717 & ~x718 & ~x726;
assign c6242 =  x132 &  x160 & ~x22 & ~x23 & ~x25 & ~x38 & ~x49 & ~x56 & ~x65 & ~x71 & ~x75 & ~x87 & ~x91 & ~x96 & ~x101 & ~x110 & ~x114 & ~x123 & ~x124 & ~x125 & ~x127 & ~x128 & ~x129 & ~x144 & ~x148 & ~x151 & ~x152 & ~x154 & ~x155 & ~x173 & ~x176 & ~x179 & ~x181 & ~x182 & ~x202 & ~x206 & ~x207 & ~x208 & ~x209 & ~x221 & ~x223 & ~x228 & ~x232 & ~x234 & ~x235 & ~x257 & ~x261 & ~x279 & ~x280 & ~x285 & ~x299 & ~x302 & ~x326 & ~x329 & ~x338 & ~x340 & ~x365 & ~x386 & ~x391 & ~x395 & ~x415 & ~x452 & ~x474 & ~x508 & ~x529 & ~x530 & ~x532 & ~x533 & ~x535 & ~x553 & ~x560 & ~x583 & ~x586 & ~x589 & ~x591 & ~x614 & ~x615 & ~x619 & ~x648 & ~x649 & ~x661 & ~x677 & ~x682 & ~x683 & ~x685 & ~x691 & ~x692 & ~x693 & ~x698 & ~x699 & ~x700 & ~x708 & ~x710 & ~x719 & ~x721 & ~x733 & ~x739 & ~x740 & ~x743 & ~x748 & ~x760 & ~x768 & ~x772 & ~x775 & ~x776;
assign c6244 =  x102 & ~x1 & ~x2 & ~x3 & ~x4 & ~x7 & ~x8 & ~x17 & ~x20 & ~x28 & ~x35 & ~x41 & ~x48 & ~x51 & ~x54 & ~x55 & ~x82 & ~x88 & ~x90 & ~x92 & ~x93 & ~x94 & ~x97 & ~x110 & ~x114 & ~x124 & ~x139 & ~x140 & ~x145 & ~x152 & ~x165 & ~x193 & ~x194 & ~x204 & ~x216 & ~x219 & ~x221 & ~x224 & ~x226 & ~x228 & ~x230 & ~x244 & ~x270 & ~x272 & ~x273 & ~x274 & ~x278 & ~x281 & ~x282 & ~x297 & ~x299 & ~x305 & ~x306 & ~x312 & ~x335 & ~x364 & ~x423 & ~x448 & ~x476 & ~x502 & ~x530 & ~x533 & ~x558 & ~x559 & ~x562 & ~x585 & ~x616 & ~x638 & ~x639 & ~x648 & ~x651 & ~x654 & ~x658 & ~x661 & ~x664 & ~x665 & ~x666 & ~x672 & ~x684 & ~x696 & ~x698 & ~x708 & ~x710 & ~x711 & ~x713 & ~x728 & ~x731 & ~x741 & ~x746 & ~x748 & ~x751 & ~x752 & ~x753 & ~x757 & ~x758 & ~x759 & ~x760 & ~x761 & ~x762 & ~x766 & ~x768 & ~x775;
assign c6246 =  x430 &  x576 &  x577 & ~x87 & ~x100 & ~x134 & ~x137 & ~x158 & ~x162 & ~x164 & ~x214 & ~x240 & ~x286 & ~x508 & ~x529 & ~x565 & ~x595 & ~x714 & ~x720 & ~x740 & ~x759 & ~x779;
assign c6248 =  x372 &  x373 &  x400 &  x427 &  x441 &  x573 &  x574 & ~x0 & ~x1 & ~x2 & ~x4 & ~x5 & ~x7 & ~x12 & ~x15 & ~x18 & ~x19 & ~x23 & ~x32 & ~x33 & ~x46 & ~x47 & ~x51 & ~x65 & ~x66 & ~x80 & ~x90 & ~x109 & ~x139 & ~x140 & ~x167 & ~x172 & ~x202 & ~x222 & ~x227 & ~x229 & ~x270 & ~x271 & ~x272 & ~x284 & ~x302 & ~x331 & ~x333 & ~x338 & ~x363 & ~x367 & ~x417 & ~x419 & ~x450 & ~x506 & ~x532 & ~x561 & ~x564 & ~x590 & ~x591 & ~x613 & ~x637 & ~x641 & ~x643 & ~x649 & ~x662 & ~x663 & ~x665 & ~x680 & ~x681 & ~x687 & ~x692 & ~x693 & ~x695 & ~x701 & ~x715 & ~x721 & ~x722 & ~x733 & ~x742 & ~x748 & ~x763 & ~x769 & ~x773 & ~x775 & ~x777 & ~x780;
assign c6250 = ~x7 & ~x14 & ~x19 & ~x26 & ~x31 & ~x37 & ~x38 & ~x40 & ~x56 & ~x58 & ~x64 & ~x67 & ~x81 & ~x84 & ~x85 & ~x115 & ~x116 & ~x121 & ~x125 & ~x126 & ~x134 & ~x140 & ~x149 & ~x173 & ~x190 & ~x192 & ~x196 & ~x206 & ~x220 & ~x224 & ~x225 & ~x235 & ~x236 & ~x244 & ~x250 & ~x252 & ~x259 & ~x263 & ~x271 & ~x272 & ~x279 & ~x281 & ~x289 & ~x298 & ~x299 & ~x310 & ~x317 & ~x324 & ~x332 & ~x337 & ~x358 & ~x359 & ~x397 & ~x442 & ~x446 & ~x451 & ~x454 & ~x482 & ~x498 & ~x504 & ~x509 & ~x525 & ~x530 & ~x532 & ~x555 & ~x560 & ~x561 & ~x589 & ~x593 & ~x608 & ~x611 & ~x614 & ~x621 & ~x635 & ~x637 & ~x649 & ~x650 & ~x651 & ~x667 & ~x672 & ~x674 & ~x677 & ~x678 & ~x684 & ~x688 & ~x690 & ~x695 & ~x697 & ~x702 & ~x706 & ~x708 & ~x710 & ~x711 & ~x720 & ~x745 & ~x749 & ~x753 & ~x757 & ~x764 & ~x765 & ~x768 & ~x773 & ~x780;
assign c6252 =  x292 &  x319 &  x346 &  x374 &  x375 &  x402 & ~x2 & ~x7 & ~x9 & ~x15 & ~x16 & ~x21 & ~x24 & ~x25 & ~x27 & ~x29 & ~x39 & ~x41 & ~x44 & ~x50 & ~x51 & ~x53 & ~x54 & ~x55 & ~x56 & ~x64 & ~x65 & ~x68 & ~x77 & ~x85 & ~x91 & ~x106 & ~x109 & ~x114 & ~x118 & ~x120 & ~x137 & ~x139 & ~x140 & ~x141 & ~x142 & ~x146 & ~x148 & ~x149 & ~x162 & ~x164 & ~x169 & ~x173 & ~x176 & ~x178 & ~x194 & ~x196 & ~x201 & ~x205 & ~x220 & ~x222 & ~x227 & ~x229 & ~x232 & ~x251 & ~x255 & ~x257 & ~x258 & ~x259 & ~x261 & ~x269 & ~x270 & ~x271 & ~x273 & ~x275 & ~x286 & ~x315 & ~x333 & ~x335 & ~x338 & ~x339 & ~x341 & ~x361 & ~x362 & ~x369 & ~x389 & ~x394 & ~x424 & ~x446 & ~x452 & ~x471 & ~x474 & ~x476 & ~x477 & ~x503 & ~x528 & ~x530 & ~x532 & ~x534 & ~x535 & ~x559 & ~x564 & ~x590 & ~x594 & ~x612 & ~x614 & ~x639 & ~x644 & ~x649 & ~x650 & ~x656 & ~x658 & ~x659 & ~x660 & ~x664 & ~x665 & ~x668 & ~x672 & ~x674 & ~x678 & ~x685 & ~x689 & ~x692 & ~x693 & ~x698 & ~x699 & ~x702 & ~x703 & ~x711 & ~x712 & ~x715 & ~x716 & ~x717 & ~x720 & ~x721 & ~x736 & ~x757 & ~x758 & ~x762 & ~x763 & ~x766 & ~x767 & ~x772 & ~x774 & ~x775 & ~x776 & ~x778 & ~x780 & ~x782 & ~x783;
assign c6254 =  x361;
assign c6256 =  x442 &  x603 & ~x183 & ~x263;
assign c6258 =  x337;
assign c6260 =  x294 &  x321 &  x348 &  x349 &  x375 &  x430 & ~x0 & ~x2 & ~x6 & ~x7 & ~x9 & ~x10 & ~x12 & ~x16 & ~x17 & ~x21 & ~x25 & ~x26 & ~x28 & ~x31 & ~x39 & ~x41 & ~x43 & ~x44 & ~x47 & ~x50 & ~x51 & ~x57 & ~x59 & ~x62 & ~x63 & ~x64 & ~x65 & ~x67 & ~x72 & ~x78 & ~x83 & ~x86 & ~x87 & ~x89 & ~x91 & ~x92 & ~x93 & ~x94 & ~x95 & ~x96 & ~x109 & ~x111 & ~x112 & ~x115 & ~x116 & ~x117 & ~x119 & ~x121 & ~x124 & ~x125 & ~x139 & ~x141 & ~x143 & ~x144 & ~x145 & ~x146 & ~x147 & ~x150 & ~x151 & ~x152 & ~x153 & ~x166 & ~x167 & ~x169 & ~x170 & ~x171 & ~x173 & ~x176 & ~x182 & ~x199 & ~x202 & ~x205 & ~x207 & ~x209 & ~x224 & ~x230 & ~x231 & ~x247 & ~x248 & ~x250 & ~x251 & ~x254 & ~x255 & ~x260 & ~x261 & ~x262 & ~x263 & ~x274 & ~x275 & ~x281 & ~x284 & ~x285 & ~x287 & ~x288 & ~x289 & ~x301 & ~x302 & ~x306 & ~x309 & ~x326 & ~x327 & ~x328 & ~x329 & ~x330 & ~x332 & ~x343 & ~x357 & ~x358 & ~x364 & ~x367 & ~x371 & ~x386 & ~x387 & ~x389 & ~x390 & ~x393 & ~x394 & ~x395 & ~x397 & ~x414 & ~x415 & ~x417 & ~x418 & ~x422 & ~x423 & ~x425 & ~x442 & ~x444 & ~x448 & ~x449 & ~x450 & ~x452 & ~x471 & ~x473 & ~x474 & ~x476 & ~x478 & ~x479 & ~x480 & ~x500 & ~x505 & ~x507 & ~x508 & ~x527 & ~x528 & ~x534 & ~x535 & ~x556 & ~x557 & ~x559 & ~x560 & ~x561 & ~x563 & ~x564 & ~x588 & ~x591 & ~x611 & ~x614 & ~x615 & ~x616 & ~x617 & ~x620 & ~x622 & ~x635 & ~x636 & ~x637 & ~x644 & ~x646 & ~x650 & ~x662 & ~x668 & ~x669 & ~x670 & ~x671 & ~x674 & ~x676 & ~x680 & ~x682 & ~x683 & ~x684 & ~x687 & ~x692 & ~x697 & ~x698 & ~x701 & ~x702 & ~x704 & ~x705 & ~x706 & ~x710 & ~x712 & ~x713 & ~x717 & ~x719 & ~x722 & ~x725 & ~x728 & ~x732 & ~x733 & ~x735 & ~x738 & ~x739 & ~x741 & ~x746 & ~x751 & ~x752 & ~x753 & ~x754 & ~x755 & ~x757 & ~x761 & ~x762 & ~x763 & ~x767 & ~x768 & ~x769 & ~x770 & ~x771 & ~x774 & ~x777 & ~x778 & ~x779 & ~x782 & ~x783;
assign c6262 =  x431 &  x487 & ~x8 & ~x11 & ~x12 & ~x19 & ~x32 & ~x33 & ~x35 & ~x41 & ~x45 & ~x48 & ~x49 & ~x55 & ~x56 & ~x59 & ~x64 & ~x66 & ~x69 & ~x77 & ~x80 & ~x82 & ~x87 & ~x88 & ~x92 & ~x94 & ~x95 & ~x106 & ~x110 & ~x111 & ~x116 & ~x117 & ~x122 & ~x123 & ~x136 & ~x137 & ~x140 & ~x162 & ~x165 & ~x171 & ~x172 & ~x177 & ~x179 & ~x190 & ~x198 & ~x202 & ~x218 & ~x220 & ~x223 & ~x225 & ~x231 & ~x234 & ~x242 & ~x243 & ~x244 & ~x245 & ~x246 & ~x247 & ~x253 & ~x254 & ~x255 & ~x269 & ~x270 & ~x271 & ~x272 & ~x275 & ~x276 & ~x279 & ~x287 & ~x289 & ~x298 & ~x301 & ~x302 & ~x303 & ~x304 & ~x305 & ~x310 & ~x328 & ~x329 & ~x330 & ~x331 & ~x333 & ~x334 & ~x336 & ~x340 & ~x360 & ~x369 & ~x372 & ~x386 & ~x387 & ~x389 & ~x391 & ~x394 & ~x398 & ~x400 & ~x401 & ~x414 & ~x418 & ~x421 & ~x425 & ~x426 & ~x428 & ~x446 & ~x447 & ~x449 & ~x450 & ~x452 & ~x454 & ~x456 & ~x472 & ~x475 & ~x476 & ~x479 & ~x480 & ~x481 & ~x483 & ~x508 & ~x527 & ~x537 & ~x538 & ~x555 & ~x558 & ~x562 & ~x563 & ~x565 & ~x567 & ~x583 & ~x585 & ~x593 & ~x594 & ~x612 & ~x613 & ~x614 & ~x616 & ~x617 & ~x621 & ~x622 & ~x623 & ~x625 & ~x636 & ~x644 & ~x650 & ~x651 & ~x662 & ~x667 & ~x669 & ~x670 & ~x680 & ~x682 & ~x690 & ~x691 & ~x694 & ~x695 & ~x700 & ~x702 & ~x703 & ~x704 & ~x708 & ~x714 & ~x716 & ~x717 & ~x721 & ~x723 & ~x724 & ~x726 & ~x729 & ~x731 & ~x732 & ~x738 & ~x740 & ~x746 & ~x751 & ~x752 & ~x754 & ~x755 & ~x757 & ~x760 & ~x766 & ~x767 & ~x768 & ~x769 & ~x773 & ~x776 & ~x777 & ~x778 & ~x779;
assign c6264 =  x571 & ~x18 & ~x30 & ~x31 & ~x36 & ~x47 & ~x49 & ~x59 & ~x60 & ~x76 & ~x84 & ~x90 & ~x110 & ~x113 & ~x135 & ~x155 & ~x189 & ~x191 & ~x195 & ~x210 & ~x217 & ~x220 & ~x229 & ~x237 & ~x255 & ~x257 & ~x305 & ~x309 & ~x363 & ~x419 & ~x445 & ~x476 & ~x530 & ~x560 & ~x565 & ~x621 & ~x623 & ~x661 & ~x706 & ~x707 & ~x717 & ~x739 & ~x744 & ~x759 & ~x760 & ~x771;
assign c6266 = ~x3 & ~x21 & ~x26 & ~x27 & ~x32 & ~x35 & ~x41 & ~x61 & ~x63 & ~x80 & ~x83 & ~x84 & ~x87 & ~x108 & ~x113 & ~x140 & ~x141 & ~x160 & ~x161 & ~x188 & ~x191 & ~x213 & ~x214 & ~x216 & ~x217 & ~x218 & ~x223 & ~x228 & ~x235 & ~x240 & ~x242 & ~x243 & ~x244 & ~x246 & ~x250 & ~x254 & ~x280 & ~x282 & ~x294 & ~x295 & ~x307 & ~x308 & ~x338 & ~x365 & ~x419 & ~x447 & ~x448 & ~x559 & ~x560 & ~x563 & ~x611 & ~x620 & ~x624 & ~x634 & ~x637 & ~x642 & ~x654 & ~x660 & ~x663 & ~x664 & ~x671 & ~x676 & ~x680 & ~x684 & ~x685 & ~x686 & ~x687 & ~x689 & ~x690 & ~x692 & ~x694 & ~x698 & ~x703 & ~x710 & ~x716 & ~x733 & ~x738 & ~x752 & ~x757 & ~x761 & ~x768 & ~x769 & ~x774 & ~x775;
assign c6268 =  x166;
assign c6270 =  x94 &  x344;
assign c6272 =  x157 &  x455 &  x483 & ~x16 & ~x25 & ~x30 & ~x31 & ~x46 & ~x50 & ~x62 & ~x67 & ~x73 & ~x82 & ~x88 & ~x96 & ~x97 & ~x115 & ~x124 & ~x125 & ~x138 & ~x140 & ~x141 & ~x149 & ~x151 & ~x152 & ~x166 & ~x170 & ~x176 & ~x177 & ~x193 & ~x194 & ~x196 & ~x200 & ~x203 & ~x227 & ~x229 & ~x252 & ~x256 & ~x257 & ~x258 & ~x270 & ~x271 & ~x272 & ~x274 & ~x283 & ~x285 & ~x297 & ~x300 & ~x303 & ~x308 & ~x309 & ~x322 & ~x324 & ~x326 & ~x332 & ~x338 & ~x340 & ~x360 & ~x361 & ~x365 & ~x392 & ~x417 & ~x419 & ~x421 & ~x424 & ~x444 & ~x506 & ~x507 & ~x560 & ~x562 & ~x563 & ~x589 & ~x592 & ~x618 & ~x621 & ~x622 & ~x623 & ~x642 & ~x643 & ~x644 & ~x649 & ~x651 & ~x666 & ~x670 & ~x672 & ~x677 & ~x681 & ~x686 & ~x687 & ~x689 & ~x691 & ~x699 & ~x702 & ~x705 & ~x706 & ~x708 & ~x718 & ~x725 & ~x733 & ~x735 & ~x737 & ~x738 & ~x744 & ~x747 & ~x748 & ~x751 & ~x753 & ~x755 & ~x761 & ~x762 & ~x763 & ~x764 & ~x768 & ~x774 & ~x782 & ~x783;
assign c6274 = ~x4 & ~x101 & ~x134 & ~x156 & ~x161 & ~x173 & ~x211 & ~x228 & ~x237 & ~x280 & ~x293 & ~x313 & ~x449 & ~x586 & ~x591 & ~x642 & ~x648 & ~x661 & ~x663 & ~x684 & ~x687 & ~x688 & ~x759 & ~x771 & ~x780;
assign c6276 =  x671;
assign c6278 =  x104 &  x131 &  x456;
assign c6280 =  x133 &  x240 & ~x113 & ~x124 & ~x181 & ~x273 & ~x326 & ~x327 & ~x329 & ~x330 & ~x359 & ~x413 & ~x609 & ~x661;
assign c6282 =  x13;
assign c6284 =  x3;
assign c6286 = ~x2 & ~x4 & ~x20 & ~x22 & ~x23 & ~x40 & ~x44 & ~x56 & ~x64 & ~x74 & ~x76 & ~x81 & ~x91 & ~x116 & ~x123 & ~x124 & ~x133 & ~x149 & ~x152 & ~x162 & ~x163 & ~x166 & ~x194 & ~x199 & ~x205 & ~x207 & ~x223 & ~x233 & ~x234 & ~x246 & ~x253 & ~x257 & ~x260 & ~x263 & ~x269 & ~x272 & ~x276 & ~x277 & ~x278 & ~x280 & ~x282 & ~x283 & ~x288 & ~x296 & ~x298 & ~x301 & ~x304 & ~x305 & ~x313 & ~x316 & ~x317 & ~x324 & ~x329 & ~x334 & ~x337 & ~x339 & ~x341 & ~x342 & ~x343 & ~x344 & ~x345 & ~x358 & ~x364 & ~x369 & ~x370 & ~x372 & ~x386 & ~x388 & ~x391 & ~x399 & ~x414 & ~x415 & ~x416 & ~x421 & ~x426 & ~x448 & ~x469 & ~x482 & ~x498 & ~x508 & ~x526 & ~x530 & ~x531 & ~x538 & ~x539 & ~x554 & ~x566 & ~x584 & ~x588 & ~x593 & ~x638 & ~x641 & ~x649 & ~x650 & ~x651 & ~x660 & ~x667 & ~x669 & ~x679 & ~x681 & ~x683 & ~x687 & ~x695 & ~x698 & ~x704 & ~x717 & ~x720 & ~x728 & ~x732 & ~x739 & ~x742 & ~x749 & ~x755 & ~x762 & ~x779 & ~x781;
assign c6288 =  x320 &  x517 & ~x10 & ~x19 & ~x34 & ~x53 & ~x70 & ~x84 & ~x89 & ~x144 & ~x189 & ~x216 & ~x218 & ~x223 & ~x226 & ~x227 & ~x246 & ~x257 & ~x315 & ~x333 & ~x342 & ~x391 & ~x470 & ~x481 & ~x554 & ~x590 & ~x635 & ~x637 & ~x659 & ~x689 & ~x694 & ~x704 & ~x709 & ~x710 & ~x719 & ~x725 & ~x726 & ~x765 & ~x770;
assign c6290 =  x399;
assign c6292 = ~x10 & ~x11 & ~x15 & ~x26 & ~x32 & ~x44 & ~x51 & ~x57 & ~x60 & ~x86 & ~x113 & ~x141 & ~x164 & ~x171 & ~x176 & ~x195 & ~x199 & ~x220 & ~x223 & ~x224 & ~x242 & ~x247 & ~x249 & ~x250 & ~x254 & ~x268 & ~x295 & ~x305 & ~x322 & ~x348 & ~x362 & ~x376 & ~x420 & ~x424 & ~x431 & ~x447 & ~x450 & ~x479 & ~x505 & ~x506 & ~x507 & ~x529 & ~x533 & ~x534 & ~x535 & ~x558 & ~x564 & ~x583 & ~x586 & ~x587 & ~x592 & ~x610 & ~x614 & ~x617 & ~x621 & ~x635 & ~x642 & ~x643 & ~x645 & ~x649 & ~x661 & ~x663 & ~x672 & ~x674 & ~x685 & ~x686 & ~x691 & ~x692 & ~x695 & ~x696 & ~x698 & ~x714 & ~x717 & ~x720 & ~x729 & ~x745 & ~x754 & ~x758 & ~x761 & ~x764 & ~x768;
assign c6294 =  x291 &  x318 &  x346 &  x401 &  x429 &  x484 &  x513 &  x541 &  x628 &  x629 & ~x2 & ~x6 & ~x10 & ~x13 & ~x14 & ~x23 & ~x25 & ~x29 & ~x34 & ~x36 & ~x39 & ~x40 & ~x41 & ~x42 & ~x43 & ~x45 & ~x46 & ~x47 & ~x49 & ~x53 & ~x55 & ~x56 & ~x58 & ~x60 & ~x61 & ~x67 & ~x69 & ~x71 & ~x72 & ~x74 & ~x79 & ~x83 & ~x89 & ~x91 & ~x92 & ~x93 & ~x96 & ~x97 & ~x99 & ~x106 & ~x107 & ~x108 & ~x109 & ~x111 & ~x112 & ~x113 & ~x114 & ~x116 & ~x121 & ~x123 & ~x139 & ~x141 & ~x142 & ~x143 & ~x144 & ~x146 & ~x148 & ~x149 & ~x150 & ~x171 & ~x178 & ~x196 & ~x197 & ~x198 & ~x201 & ~x203 & ~x204 & ~x205 & ~x222 & ~x223 & ~x224 & ~x226 & ~x227 & ~x229 & ~x230 & ~x248 & ~x249 & ~x250 & ~x253 & ~x254 & ~x259 & ~x269 & ~x270 & ~x274 & ~x276 & ~x277 & ~x278 & ~x281 & ~x284 & ~x285 & ~x287 & ~x302 & ~x303 & ~x305 & ~x307 & ~x309 & ~x310 & ~x311 & ~x315 & ~x330 & ~x334 & ~x336 & ~x337 & ~x359 & ~x360 & ~x361 & ~x364 & ~x366 & ~x367 & ~x387 & ~x389 & ~x391 & ~x394 & ~x397 & ~x418 & ~x422 & ~x423 & ~x424 & ~x425 & ~x445 & ~x446 & ~x448 & ~x449 & ~x451 & ~x453 & ~x474 & ~x480 & ~x505 & ~x506 & ~x508 & ~x528 & ~x529 & ~x535 & ~x554 & ~x557 & ~x562 & ~x563 & ~x582 & ~x584 & ~x585 & ~x586 & ~x589 & ~x591 & ~x592 & ~x593 & ~x594 & ~x609 & ~x610 & ~x611 & ~x613 & ~x615 & ~x618 & ~x622 & ~x638 & ~x639 & ~x641 & ~x644 & ~x645 & ~x647 & ~x648 & ~x651 & ~x663 & ~x666 & ~x669 & ~x671 & ~x673 & ~x674 & ~x676 & ~x677 & ~x678 & ~x679 & ~x682 & ~x684 & ~x691 & ~x694 & ~x696 & ~x698 & ~x700 & ~x705 & ~x707 & ~x710 & ~x715 & ~x717 & ~x718 & ~x719 & ~x721 & ~x726 & ~x727 & ~x731 & ~x733 & ~x734 & ~x736 & ~x737 & ~x738 & ~x739 & ~x741 & ~x746 & ~x749 & ~x750 & ~x752 & ~x757 & ~x765 & ~x766 & ~x769 & ~x770 & ~x771 & ~x774 & ~x775 & ~x777 & ~x778 & ~x781 & ~x783;
assign c6296 =  x131 &  x158 &  x185 & ~x28 & ~x46 & ~x50 & ~x60 & ~x66 & ~x116 & ~x120 & ~x139 & ~x148 & ~x149 & ~x150 & ~x152 & ~x153 & ~x178 & ~x179 & ~x207 & ~x221 & ~x223 & ~x230 & ~x234 & ~x246 & ~x247 & ~x273 & ~x274 & ~x275 & ~x276 & ~x301 & ~x303 & ~x330 & ~x354 & ~x357 & ~x358 & ~x379 & ~x388 & ~x450 & ~x476 & ~x477 & ~x590 & ~x610 & ~x621 & ~x622 & ~x638 & ~x640 & ~x648 & ~x649 & ~x663 & ~x686 & ~x697 & ~x708 & ~x741 & ~x744 & ~x746 & ~x748 & ~x764 & ~x781;
assign c6298 =  x374 &  x458 &  x486 &  x630 & ~x2 & ~x6 & ~x8 & ~x9 & ~x10 & ~x16 & ~x17 & ~x27 & ~x37 & ~x42 & ~x51 & ~x59 & ~x61 & ~x70 & ~x74 & ~x85 & ~x91 & ~x92 & ~x109 & ~x110 & ~x111 & ~x119 & ~x120 & ~x141 & ~x144 & ~x172 & ~x173 & ~x175 & ~x193 & ~x204 & ~x205 & ~x219 & ~x220 & ~x229 & ~x231 & ~x267 & ~x271 & ~x274 & ~x275 & ~x282 & ~x307 & ~x336 & ~x337 & ~x358 & ~x365 & ~x367 & ~x388 & ~x394 & ~x398 & ~x416 & ~x450 & ~x452 & ~x474 & ~x478 & ~x479 & ~x530 & ~x536 & ~x537 & ~x539 & ~x557 & ~x562 & ~x583 & ~x587 & ~x594 & ~x595 & ~x622 & ~x647 & ~x668 & ~x676 & ~x677 & ~x681 & ~x695 & ~x698 & ~x701 & ~x702 & ~x719 & ~x743 & ~x750 & ~x752 & ~x753 & ~x754 & ~x757 & ~x762 & ~x765 & ~x772 & ~x776 & ~x781;
assign c61 =  x234 & ~x2 & ~x13 & ~x29 & ~x32 & ~x50 & ~x53 & ~x59 & ~x66 & ~x75 & ~x81 & ~x94 & ~x95 & ~x106 & ~x117 & ~x118 & ~x139 & ~x140 & ~x167 & ~x172 & ~x194 & ~x222 & ~x226 & ~x283 & ~x310 & ~x339 & ~x359 & ~x373 & ~x422 & ~x423 & ~x477 & ~x479 & ~x503 & ~x534 & ~x559 & ~x561 & ~x563 & ~x587 & ~x640 & ~x644 & ~x646 & ~x691 & ~x694 & ~x711 & ~x714 & ~x717 & ~x749 & ~x751 & ~x752 & ~x771;
assign c63 =  x273 &  x301 & ~x0 & ~x5 & ~x6 & ~x7 & ~x8 & ~x25 & ~x28 & ~x35 & ~x38 & ~x40 & ~x41 & ~x42 & ~x44 & ~x48 & ~x50 & ~x53 & ~x57 & ~x68 & ~x70 & ~x74 & ~x78 & ~x79 & ~x84 & ~x85 & ~x90 & ~x93 & ~x94 & ~x96 & ~x103 & ~x106 & ~x114 & ~x115 & ~x117 & ~x118 & ~x120 & ~x122 & ~x124 & ~x142 & ~x166 & ~x168 & ~x169 & ~x170 & ~x173 & ~x177 & ~x196 & ~x197 & ~x199 & ~x201 & ~x230 & ~x251 & ~x255 & ~x280 & ~x306 & ~x308 & ~x311 & ~x337 & ~x338 & ~x362 & ~x365 & ~x417 & ~x419 & ~x421 & ~x448 & ~x474 & ~x477 & ~x506 & ~x533 & ~x534 & ~x558 & ~x560 & ~x583 & ~x584 & ~x609 & ~x611 & ~x638 & ~x664 & ~x665 & ~x670 & ~x671 & ~x676 & ~x678 & ~x691 & ~x693 & ~x696 & ~x697 & ~x700 & ~x705 & ~x717 & ~x718 & ~x724 & ~x729 & ~x731 & ~x741 & ~x744 & ~x747 & ~x751 & ~x754 & ~x755 & ~x759 & ~x765 & ~x770 & ~x775 & ~x776 & ~x779 & ~x783;
assign c65 = ~x46 & ~x48 & ~x58 & ~x84 & ~x92 & ~x96 & ~x228 & ~x251 & ~x305 & ~x312 & ~x335 & ~x420 & ~x455 & ~x456 & ~x485 & ~x515 & ~x516 & ~x517 & ~x645 & ~x719 & ~x722 & ~x733 & ~x737 & ~x762 & ~x774;
assign c67 =  x263 & ~x3 & ~x7 & ~x13 & ~x14 & ~x19 & ~x23 & ~x26 & ~x28 & ~x45 & ~x46 & ~x50 & ~x54 & ~x55 & ~x66 & ~x67 & ~x68 & ~x91 & ~x95 & ~x97 & ~x98 & ~x99 & ~x103 & ~x117 & ~x126 & ~x128 & ~x130 & ~x131 & ~x132 & ~x143 & ~x149 & ~x152 & ~x154 & ~x157 & ~x167 & ~x172 & ~x173 & ~x177 & ~x195 & ~x202 & ~x229 & ~x250 & ~x251 & ~x307 & ~x335 & ~x362 & ~x364 & ~x394 & ~x419 & ~x422 & ~x474 & ~x505 & ~x508 & ~x585 & ~x586 & ~x593 & ~x642 & ~x644 & ~x675 & ~x695 & ~x698 & ~x699 & ~x700 & ~x719 & ~x730 & ~x732 & ~x756 & ~x758 & ~x759 & ~x762 & ~x765 & ~x766 & ~x768;
assign c69 =  x123 & ~x26 & ~x290 & ~x316 & ~x387 & ~x561 & ~x589 & ~x716;
assign c611 = ~x5 & ~x6 & ~x8 & ~x9 & ~x11 & ~x12 & ~x14 & ~x15 & ~x18 & ~x19 & ~x20 & ~x24 & ~x25 & ~x28 & ~x30 & ~x36 & ~x38 & ~x46 & ~x48 & ~x51 & ~x52 & ~x55 & ~x63 & ~x69 & ~x72 & ~x75 & ~x80 & ~x81 & ~x82 & ~x84 & ~x86 & ~x87 & ~x90 & ~x92 & ~x96 & ~x98 & ~x99 & ~x105 & ~x110 & ~x112 & ~x114 & ~x121 & ~x128 & ~x131 & ~x134 & ~x139 & ~x140 & ~x144 & ~x167 & ~x193 & ~x197 & ~x198 & ~x201 & ~x225 & ~x226 & ~x250 & ~x256 & ~x277 & ~x308 & ~x310 & ~x337 & ~x338 & ~x340 & ~x347 & ~x363 & ~x365 & ~x394 & ~x445 & ~x446 & ~x447 & ~x448 & ~x449 & ~x450 & ~x451 & ~x477 & ~x480 & ~x504 & ~x506 & ~x532 & ~x535 & ~x560 & ~x562 & ~x565 & ~x566 & ~x586 & ~x588 & ~x596 & ~x613 & ~x618 & ~x619 & ~x620 & ~x646 & ~x648 & ~x649 & ~x653 & ~x654 & ~x669 & ~x678 & ~x695 & ~x700 & ~x704 & ~x705 & ~x709 & ~x711 & ~x714 & ~x717 & ~x718 & ~x723 & ~x733 & ~x738 & ~x748 & ~x751 & ~x756 & ~x758 & ~x762 & ~x764 & ~x770 & ~x771 & ~x778 & ~x779;
assign c613 =  x622;
assign c615 =  x152 &  x177 & ~x0 & ~x51 & ~x63 & ~x86 & ~x359 & ~x387 & ~x393 & ~x415 & ~x447 & ~x562 & ~x764;
assign c617 =  x325 & ~x0 & ~x1 & ~x4 & ~x6 & ~x7 & ~x8 & ~x12 & ~x14 & ~x18 & ~x25 & ~x28 & ~x36 & ~x37 & ~x40 & ~x47 & ~x48 & ~x57 & ~x78 & ~x79 & ~x82 & ~x83 & ~x86 & ~x91 & ~x93 & ~x108 & ~x111 & ~x112 & ~x113 & ~x118 & ~x120 & ~x138 & ~x139 & ~x146 & ~x165 & ~x168 & ~x169 & ~x170 & ~x172 & ~x191 & ~x195 & ~x196 & ~x197 & ~x199 & ~x203 & ~x219 & ~x231 & ~x232 & ~x246 & ~x249 & ~x254 & ~x278 & ~x306 & ~x309 & ~x315 & ~x336 & ~x337 & ~x341 & ~x342 & ~x358 & ~x362 & ~x368 & ~x369 & ~x383 & ~x384 & ~x386 & ~x390 & ~x412 & ~x419 & ~x424 & ~x439 & ~x441 & ~x448 & ~x449 & ~x477 & ~x478 & ~x501 & ~x503 & ~x505 & ~x506 & ~x508 & ~x534 & ~x535 & ~x587 & ~x617 & ~x618 & ~x619 & ~x641 & ~x642 & ~x645 & ~x648 & ~x663 & ~x666 & ~x669 & ~x670 & ~x671 & ~x673 & ~x675 & ~x680 & ~x682 & ~x693 & ~x694 & ~x696 & ~x698 & ~x703 & ~x706 & ~x714 & ~x719 & ~x720 & ~x723 & ~x727 & ~x728 & ~x729 & ~x732 & ~x733 & ~x736 & ~x738 & ~x740 & ~x741 & ~x742 & ~x746 & ~x747 & ~x751 & ~x753 & ~x756 & ~x763 & ~x764 & ~x766 & ~x768 & ~x769 & ~x773 & ~x774 & ~x777 & ~x779;
assign c619 =  x157 & ~x265 & ~x317;
assign c621 =  x271 & ~x66 & ~x94 & ~x96 & ~x112 & ~x147 & ~x165 & ~x176 & ~x363 & ~x419 & ~x601;
assign c623 =  x267 & ~x9 & ~x18 & ~x21 & ~x24 & ~x29 & ~x34 & ~x44 & ~x47 & ~x52 & ~x59 & ~x61 & ~x65 & ~x69 & ~x78 & ~x84 & ~x102 & ~x103 & ~x104 & ~x106 & ~x107 & ~x166 & ~x168 & ~x170 & ~x196 & ~x225 & ~x253 & ~x254 & ~x280 & ~x307 & ~x361 & ~x392 & ~x445 & ~x471 & ~x475 & ~x476 & ~x477 & ~x481 & ~x486 & ~x508 & ~x512 & ~x530 & ~x533 & ~x537 & ~x564 & ~x614 & ~x617 & ~x674 & ~x693 & ~x695 & ~x697 & ~x700 & ~x701 & ~x704 & ~x725 & ~x727 & ~x733 & ~x742 & ~x751 & ~x760 & ~x775 & ~x777 & ~x782;
assign c625 =  x538 & ~x105 & ~x117 & ~x138 & ~x195 & ~x253 & ~x260 & ~x434 & ~x697 & ~x699 & ~x702 & ~x729 & ~x730;
assign c627 =  x432 &  x434 &  x462 & ~x11 & ~x124 & ~x164 & ~x389 & ~x393 & ~x446 & ~x524 & ~x549 & ~x561 & ~x608 & ~x645 & ~x646 & ~x664;
assign c629 = ~x15 & ~x25 & ~x39 & ~x41 & ~x50 & ~x62 & ~x67 & ~x69 & ~x166 & ~x304 & ~x307 & ~x335 & ~x367 & ~x422 & ~x453 & ~x483 & ~x486 & ~x556 & ~x589 & ~x612 & ~x615 & ~x617 & ~x640 & ~x646 & ~x710 & ~x722 & ~x750 & ~x756 & ~x763 & ~x769 & ~x776;
assign c631 =  x610 & ~x290;
assign c633 =  x259 & ~x2 & ~x28 & ~x45 & ~x46 & ~x53 & ~x60 & ~x64 & ~x70 & ~x73 & ~x366 & ~x395 & ~x528 & ~x547 & ~x611 & ~x675 & ~x701 & ~x728 & ~x731 & ~x732 & ~x748;
assign c635 = ~x125 & ~x126 & ~x129 & ~x157 & ~x166 & ~x414 & ~x547 & ~x559 & ~x576 & ~x633;
assign c637 =  x213 & ~x9 & ~x20 & ~x32 & ~x35 & ~x41 & ~x55 & ~x61 & ~x102 & ~x114 & ~x131 & ~x144 & ~x169 & ~x172 & ~x278 & ~x434 & ~x435 & ~x586 & ~x587 & ~x590 & ~x616 & ~x619 & ~x673 & ~x678 & ~x702 & ~x714 & ~x731 & ~x740 & ~x741 & ~x744 & ~x750 & ~x770 & ~x771;
assign c639 =  x355 & ~x6 & ~x31 & ~x34 & ~x66 & ~x74 & ~x100 & ~x113 & ~x118 & ~x120 & ~x146 & ~x171 & ~x197 & ~x200 & ~x225 & ~x253 & ~x279 & ~x308 & ~x335 & ~x359 & ~x361 & ~x365 & ~x377 & ~x379 & ~x387 & ~x407 & ~x417 & ~x474 & ~x562 & ~x586 & ~x589 & ~x618 & ~x644 & ~x650 & ~x681 & ~x696 & ~x697 & ~x711 & ~x717 & ~x727 & ~x737 & ~x744 & ~x749 & ~x752 & ~x764 & ~x765 & ~x774;
assign c641 = ~x4 & ~x19 & ~x20 & ~x21 & ~x24 & ~x26 & ~x54 & ~x64 & ~x65 & ~x67 & ~x72 & ~x77 & ~x78 & ~x81 & ~x89 & ~x106 & ~x107 & ~x113 & ~x167 & ~x195 & ~x199 & ~x253 & ~x274 & ~x281 & ~x331 & ~x337 & ~x364 & ~x367 & ~x419 & ~x420 & ~x474 & ~x484 & ~x485 & ~x488 & ~x511 & ~x557 & ~x618 & ~x640 & ~x641 & ~x644 & ~x666 & ~x672 & ~x673 & ~x714 & ~x717 & ~x725 & ~x734 & ~x737 & ~x743 & ~x756 & ~x765 & ~x767;
assign c643 =  x239 & ~x393 & ~x485 & ~x497;
assign c645 = ~x1 & ~x3 & ~x8 & ~x10 & ~x26 & ~x61 & ~x105 & ~x110 & ~x112 & ~x132 & ~x141 & ~x272 & ~x283 & ~x287 & ~x316 & ~x319 & ~x320 & ~x332 & ~x343 & ~x359 & ~x370 & ~x397 & ~x453 & ~x656 & ~x673 & ~x676 & ~x698 & ~x703 & ~x705 & ~x755 & ~x759;
assign c647 =  x241 &  x298 &  x326 & ~x28 & ~x163 & ~x330 & ~x619 & ~x705 & ~x754;
assign c649 = ~x67 & ~x122 & ~x145 & ~x359 & ~x430 & ~x601;
assign c651 =  x272 & ~x63 & ~x166 & ~x322 & ~x325 & ~x337 & ~x350 & ~x379 & ~x446 & ~x478 & ~x503 & ~x658 & ~x659 & ~x660 & ~x698 & ~x765;
assign c653 =  x211 &  x212 &  x269 & ~x7 & ~x15 & ~x28 & ~x33 & ~x37 & ~x38 & ~x78 & ~x85 & ~x86 & ~x90 & ~x102 & ~x116 & ~x117 & ~x133 & ~x363 & ~x449 & ~x477 & ~x591 & ~x647 & ~x672 & ~x699 & ~x705 & ~x741 & ~x760 & ~x763 & ~x775 & ~x783;
assign c655 =  x185 & ~x101 & ~x159 & ~x237 & ~x266 & ~x341 & ~x421 & ~x422;
assign c657 =  x622;
assign c659 =  x272 &  x355 &  x382 & ~x5 & ~x9 & ~x36 & ~x42 & ~x43 & ~x49 & ~x52 & ~x60 & ~x63 & ~x66 & ~x69 & ~x83 & ~x90 & ~x94 & ~x115 & ~x145 & ~x168 & ~x171 & ~x332 & ~x358 & ~x365 & ~x387 & ~x418 & ~x707 & ~x736 & ~x746 & ~x759 & ~x761 & ~x762 & ~x765 & ~x768 & ~x778 & ~x779;
assign c661 = ~x48 & ~x60 & ~x92 & ~x105 & ~x111 & ~x117 & ~x137 & ~x139 & ~x140 & ~x144 & ~x172 & ~x198 & ~x224 & ~x253 & ~x278 & ~x332 & ~x336 & ~x340 & ~x420 & ~x428 & ~x449 & ~x455 & ~x456 & ~x457 & ~x486 & ~x492 & ~x493 & ~x504 & ~x563 & ~x675 & ~x676 & ~x681 & ~x691 & ~x708 & ~x724 & ~x735 & ~x739 & ~x741 & ~x773 & ~x779;
assign c663 =  x623 & ~x103 & ~x397;
assign c665 =  x653 & ~x132 & ~x512;
assign c667 =  x180 &  x571 &  x599 & ~x19 & ~x23 & ~x143 & ~x194 & ~x257 & ~x303 & ~x331 & ~x368 & ~x389 & ~x418 & ~x429 & ~x455 & ~x535 & ~x641 & ~x667 & ~x670 & ~x712 & ~x769;
assign c669 =  x290 & ~x13 & ~x56 & ~x120 & ~x149 & ~x372 & ~x400 & ~x401 & ~x402 & ~x473 & ~x504 & ~x734;
assign c671 = ~x2 & ~x61 & ~x63 & ~x76 & ~x89 & ~x108 & ~x109 & ~x117 & ~x142 & ~x165 & ~x166 & ~x253 & ~x280 & ~x338 & ~x359 & ~x360 & ~x366 & ~x386 & ~x447 & ~x505 & ~x506 & ~x547 & ~x548 & ~x562 & ~x564 & ~x576 & ~x581 & ~x588 & ~x591 & ~x608 & ~x618 & ~x632 & ~x637 & ~x646 & ~x648 & ~x649 & ~x680 & ~x681 & ~x697 & ~x700 & ~x712 & ~x723 & ~x730 & ~x743 & ~x754 & ~x757 & ~x761 & ~x782;
assign c673 =  x217 & ~x313 & ~x486 & ~x489;
assign c675 =  x213 &  x569 & ~x12 & ~x21 & ~x23 & ~x24 & ~x31 & ~x33 & ~x51 & ~x83 & ~x85 & ~x89 & ~x114 & ~x130 & ~x132 & ~x138 & ~x160 & ~x161 & ~x165 & ~x171 & ~x222 & ~x226 & ~x228 & ~x231 & ~x251 & ~x254 & ~x312 & ~x390 & ~x394 & ~x501 & ~x502 & ~x505 & ~x621 & ~x636 & ~x644 & ~x663 & ~x678 & ~x682 & ~x683 & ~x684 & ~x686 & ~x691 & ~x696 & ~x733 & ~x736 & ~x750 & ~x772 & ~x773 & ~x777;
assign c677 =  x241 & ~x24 & ~x32 & ~x43 & ~x114 & ~x131 & ~x133 & ~x135 & ~x249 & ~x306 & ~x369 & ~x504 & ~x618 & ~x633 & ~x634 & ~x659 & ~x668 & ~x674 & ~x694 & ~x703 & ~x709 & ~x713 & ~x715 & ~x725 & ~x741 & ~x761 & ~x781;
assign c679 =  x153 &  x625 & ~x313 & ~x646 & ~x781;
assign c681 = ~x31 & ~x90 & ~x138 & ~x192 & ~x294 & ~x322 & ~x343 & ~x345 & ~x363 & ~x386 & ~x388 & ~x448 & ~x471 & ~x529 & ~x685 & ~x699 & ~x728 & ~x743;
assign c683 =  x409 &  x491 & ~x129 & ~x154 & ~x553 & ~x571;
assign c685 =  x188 & ~x29 & ~x66 & ~x144 & ~x168 & ~x295 & ~x605 & ~x662 & ~x671 & ~x685;
assign c687 =  x438 &  x465 & ~x0 & ~x4 & ~x8 & ~x12 & ~x13 & ~x16 & ~x20 & ~x22 & ~x23 & ~x26 & ~x30 & ~x36 & ~x40 & ~x52 & ~x57 & ~x64 & ~x70 & ~x72 & ~x75 & ~x76 & ~x78 & ~x84 & ~x90 & ~x96 & ~x97 & ~x99 & ~x101 & ~x103 & ~x106 & ~x117 & ~x118 & ~x119 & ~x122 & ~x123 & ~x125 & ~x126 & ~x128 & ~x131 & ~x135 & ~x137 & ~x140 & ~x141 & ~x171 & ~x194 & ~x195 & ~x197 & ~x222 & ~x223 & ~x226 & ~x251 & ~x254 & ~x276 & ~x281 & ~x306 & ~x335 & ~x338 & ~x363 & ~x366 & ~x367 & ~x393 & ~x395 & ~x421 & ~x447 & ~x449 & ~x474 & ~x476 & ~x479 & ~x505 & ~x506 & ~x507 & ~x563 & ~x566 & ~x584 & ~x588 & ~x589 & ~x590 & ~x595 & ~x615 & ~x618 & ~x619 & ~x620 & ~x621 & ~x637 & ~x640 & ~x641 & ~x642 & ~x643 & ~x644 & ~x649 & ~x650 & ~x653 & ~x667 & ~x672 & ~x673 & ~x676 & ~x699 & ~x701 & ~x706 & ~x707 & ~x712 & ~x714 & ~x726 & ~x727 & ~x728 & ~x729 & ~x769 & ~x777 & ~x779 & ~x780;
assign c689 = ~x0 & ~x4 & ~x6 & ~x7 & ~x13 & ~x14 & ~x15 & ~x16 & ~x21 & ~x22 & ~x23 & ~x25 & ~x26 & ~x28 & ~x31 & ~x40 & ~x42 & ~x43 & ~x47 & ~x50 & ~x52 & ~x53 & ~x57 & ~x58 & ~x63 & ~x68 & ~x69 & ~x70 & ~x72 & ~x77 & ~x82 & ~x84 & ~x85 & ~x86 & ~x87 & ~x89 & ~x90 & ~x92 & ~x93 & ~x94 & ~x95 & ~x96 & ~x98 & ~x99 & ~x100 & ~x106 & ~x108 & ~x109 & ~x110 & ~x116 & ~x118 & ~x119 & ~x120 & ~x121 & ~x122 & ~x123 & ~x125 & ~x126 & ~x130 & ~x132 & ~x135 & ~x146 & ~x153 & ~x169 & ~x170 & ~x171 & ~x173 & ~x181 & ~x194 & ~x196 & ~x197 & ~x198 & ~x200 & ~x223 & ~x224 & ~x252 & ~x277 & ~x278 & ~x332 & ~x333 & ~x335 & ~x336 & ~x338 & ~x339 & ~x363 & ~x365 & ~x449 & ~x450 & ~x473 & ~x476 & ~x477 & ~x479 & ~x502 & ~x503 & ~x506 & ~x507 & ~x529 & ~x532 & ~x533 & ~x534 & ~x562 & ~x563 & ~x571 & ~x586 & ~x589 & ~x591 & ~x618 & ~x619 & ~x620 & ~x645 & ~x647 & ~x670 & ~x671 & ~x676 & ~x680 & ~x695 & ~x699 & ~x700 & ~x703 & ~x706 & ~x709 & ~x723 & ~x730 & ~x734 & ~x735 & ~x736 & ~x738 & ~x749 & ~x750 & ~x751 & ~x757 & ~x760 & ~x762 & ~x764 & ~x769 & ~x773 & ~x776 & ~x777 & ~x779 & ~x780 & ~x782;
assign c691 = ~x35 & ~x39 & ~x54 & ~x57 & ~x59 & ~x98 & ~x99 & ~x123 & ~x359 & ~x364 & ~x437 & ~x446 & ~x485 & ~x486 & ~x528 & ~x586 & ~x643 & ~x727 & ~x750;
assign c693 = ~x6 & ~x17 & ~x27 & ~x32 & ~x57 & ~x70 & ~x135 & ~x141 & ~x144 & ~x154 & ~x163 & ~x165 & ~x184 & ~x198 & ~x280 & ~x310 & ~x394 & ~x557 & ~x575 & ~x576 & ~x602 & ~x604 & ~x605 & ~x619 & ~x629 & ~x632 & ~x695 & ~x717 & ~x728 & ~x757 & ~x758 & ~x774;
assign c695 =  x352 &  x380 & ~x195 & ~x201 & ~x252 & ~x278 & ~x370 & ~x371 & ~x466 & ~x496 & ~x508 & ~x701 & ~x757 & ~x760;
assign c697 =  x269 & ~x121 & ~x122 & ~x570;
assign c699 =  x656 & ~x5 & ~x21 & ~x64 & ~x66 & ~x103 & ~x128 & ~x136 & ~x254 & ~x541 & ~x675 & ~x679 & ~x736 & ~x778;
assign c6101 = ~x7 & ~x10 & ~x17 & ~x24 & ~x26 & ~x28 & ~x32 & ~x33 & ~x40 & ~x44 & ~x49 & ~x57 & ~x60 & ~x61 & ~x72 & ~x74 & ~x85 & ~x91 & ~x93 & ~x104 & ~x106 & ~x107 & ~x120 & ~x121 & ~x123 & ~x126 & ~x128 & ~x133 & ~x144 & ~x146 & ~x155 & ~x176 & ~x177 & ~x178 & ~x201 & ~x255 & ~x280 & ~x363 & ~x367 & ~x392 & ~x450 & ~x472 & ~x514 & ~x557 & ~x589 & ~x590 & ~x591 & ~x610 & ~x615 & ~x619 & ~x647 & ~x663 & ~x670 & ~x705 & ~x707 & ~x715 & ~x717 & ~x718 & ~x721 & ~x723 & ~x728 & ~x744 & ~x755 & ~x783;
assign c6103 = ~x1 & ~x5 & ~x17 & ~x24 & ~x27 & ~x36 & ~x50 & ~x54 & ~x63 & ~x68 & ~x78 & ~x79 & ~x111 & ~x256 & ~x336 & ~x358 & ~x361 & ~x425 & ~x442 & ~x444 & ~x457 & ~x459 & ~x475 & ~x477 & ~x488 & ~x560 & ~x643 & ~x647 & ~x721 & ~x726 & ~x741;
assign c6105 =  x302 & ~x73 & ~x352 & ~x353 & ~x378 & ~x379 & ~x380 & ~x408 & ~x677 & ~x715 & ~x750 & ~x769 & ~x778;
assign c6107 = ~x21 & ~x49 & ~x84 & ~x116 & ~x168 & ~x199 & ~x282 & ~x287 & ~x313 & ~x342 & ~x344 & ~x404 & ~x429 & ~x508 & ~x615 & ~x617 & ~x661 & ~x720 & ~x723 & ~x740;
assign c6109 =  x275 & ~x96 & ~x120 & ~x121 & ~x125 & ~x606;
assign c6111 =  x214 &  x270 & ~x5 & ~x21 & ~x33 & ~x38 & ~x39 & ~x47 & ~x48 & ~x57 & ~x94 & ~x121 & ~x134 & ~x140 & ~x168 & ~x203 & ~x249 & ~x363 & ~x365 & ~x366 & ~x474 & ~x476 & ~x504 & ~x559 & ~x562 & ~x616 & ~x632 & ~x639 & ~x664 & ~x674 & ~x691 & ~x697 & ~x747 & ~x756 & ~x765 & ~x768;
assign c6113 =  x184 & ~x54 & ~x74 & ~x81 & ~x91 & ~x93 & ~x118 & ~x168 & ~x198 & ~x336 & ~x491 & ~x514 & ~x533 & ~x645 & ~x744 & ~x754;
assign c6115 =  x325 &  x408 & ~x2 & ~x4 & ~x5 & ~x10 & ~x14 & ~x19 & ~x20 & ~x23 & ~x25 & ~x32 & ~x38 & ~x42 & ~x43 & ~x48 & ~x50 & ~x51 & ~x53 & ~x58 & ~x59 & ~x62 & ~x76 & ~x77 & ~x86 & ~x91 & ~x92 & ~x106 & ~x108 & ~x110 & ~x114 & ~x116 & ~x136 & ~x137 & ~x138 & ~x140 & ~x142 & ~x165 & ~x166 & ~x167 & ~x169 & ~x172 & ~x224 & ~x228 & ~x229 & ~x254 & ~x255 & ~x281 & ~x283 & ~x285 & ~x308 & ~x309 & ~x311 & ~x313 & ~x335 & ~x340 & ~x359 & ~x362 & ~x363 & ~x364 & ~x384 & ~x386 & ~x395 & ~x412 & ~x414 & ~x420 & ~x451 & ~x479 & ~x502 & ~x503 & ~x531 & ~x535 & ~x588 & ~x616 & ~x643 & ~x648 & ~x664 & ~x670 & ~x673 & ~x692 & ~x697 & ~x698 & ~x699 & ~x701 & ~x704 & ~x706 & ~x707 & ~x715 & ~x719 & ~x720 & ~x721 & ~x728 & ~x731 & ~x734 & ~x736 & ~x738 & ~x741 & ~x742 & ~x744 & ~x746 & ~x748 & ~x749 & ~x750 & ~x751 & ~x754 & ~x757 & ~x758 & ~x760 & ~x761 & ~x764 & ~x765 & ~x768 & ~x774 & ~x778 & ~x779 & ~x782 & ~x783;
assign c6117 =  x214 & ~x29 & ~x107 & ~x132 & ~x405 & ~x491;
assign c6119 =  x556;
assign c6121 = ~x9 & ~x19 & ~x22 & ~x47 & ~x56 & ~x70 & ~x99 & ~x100 & ~x157 & ~x162 & ~x171 & ~x186 & ~x191 & ~x218 & ~x254 & ~x343 & ~x356 & ~x383 & ~x385 & ~x649 & ~x654 & ~x669 & ~x690 & ~x709 & ~x768 & ~x771;
assign c6123 =  x206 &  x207 &  x208 &  x230;
assign c6125 =  x275 & ~x11 & ~x121 & ~x126 & ~x313 & ~x475 & ~x701 & ~x748;
assign c6127 =  x208 & ~x1 & ~x100 & ~x162 & ~x423 & ~x438 & ~x544 & ~x667 & ~x680 & ~x691 & ~x716;
assign c6129 = ~x45 & ~x62 & ~x92 & ~x118 & ~x126 & ~x167 & ~x249 & ~x541 & ~x544 & ~x567 & ~x571 & ~x599 & ~x615 & ~x640 & ~x642 & ~x645 & ~x720 & ~x729;
assign c6131 =  x296 & ~x1 & ~x5 & ~x9 & ~x15 & ~x18 & ~x24 & ~x26 & ~x34 & ~x54 & ~x65 & ~x73 & ~x74 & ~x77 & ~x78 & ~x80 & ~x81 & ~x85 & ~x89 & ~x104 & ~x116 & ~x131 & ~x133 & ~x134 & ~x138 & ~x139 & ~x144 & ~x159 & ~x160 & ~x162 & ~x163 & ~x165 & ~x170 & ~x171 & ~x194 & ~x195 & ~x198 & ~x218 & ~x221 & ~x224 & ~x226 & ~x251 & ~x253 & ~x254 & ~x278 & ~x302 & ~x307 & ~x308 & ~x309 & ~x329 & ~x335 & ~x362 & ~x364 & ~x366 & ~x384 & ~x388 & ~x390 & ~x398 & ~x417 & ~x418 & ~x421 & ~x447 & ~x448 & ~x451 & ~x475 & ~x480 & ~x503 & ~x504 & ~x507 & ~x532 & ~x534 & ~x586 & ~x614 & ~x619 & ~x641 & ~x650 & ~x680 & ~x683 & ~x690 & ~x698 & ~x705 & ~x709 & ~x715 & ~x718 & ~x726 & ~x731 & ~x734 & ~x735 & ~x744 & ~x753 & ~x755 & ~x756 & ~x757 & ~x763 & ~x766 & ~x769 & ~x770 & ~x774;
assign c6133 = ~x17 & ~x21 & ~x26 & ~x33 & ~x44 & ~x50 & ~x69 & ~x70 & ~x74 & ~x77 & ~x81 & ~x91 & ~x95 & ~x96 & ~x106 & ~x109 & ~x111 & ~x113 & ~x123 & ~x136 & ~x166 & ~x167 & ~x168 & ~x169 & ~x191 & ~x192 & ~x198 & ~x219 & ~x250 & ~x278 & ~x282 & ~x307 & ~x336 & ~x363 & ~x367 & ~x391 & ~x421 & ~x476 & ~x479 & ~x505 & ~x530 & ~x532 & ~x533 & ~x543 & ~x544 & ~x555 & ~x556 & ~x568 & ~x569 & ~x570 & ~x581 & ~x611 & ~x613 & ~x615 & ~x617 & ~x673 & ~x703 & ~x722 & ~x728 & ~x729 & ~x733 & ~x735 & ~x750 & ~x752 & ~x757 & ~x768;
assign c6135 =  x324 & ~x4 & ~x6 & ~x11 & ~x13 & ~x22 & ~x23 & ~x24 & ~x25 & ~x26 & ~x33 & ~x44 & ~x60 & ~x62 & ~x67 & ~x68 & ~x69 & ~x70 & ~x74 & ~x75 & ~x77 & ~x81 & ~x82 & ~x86 & ~x87 & ~x89 & ~x91 & ~x113 & ~x118 & ~x135 & ~x139 & ~x142 & ~x146 & ~x164 & ~x170 & ~x171 & ~x191 & ~x196 & ~x197 & ~x244 & ~x275 & ~x276 & ~x286 & ~x310 & ~x313 & ~x334 & ~x338 & ~x355 & ~x357 & ~x360 & ~x364 & ~x369 & ~x383 & ~x385 & ~x386 & ~x416 & ~x418 & ~x424 & ~x479 & ~x505 & ~x530 & ~x531 & ~x532 & ~x535 & ~x563 & ~x587 & ~x589 & ~x638 & ~x639 & ~x642 & ~x644 & ~x645 & ~x665 & ~x668 & ~x673 & ~x675 & ~x676 & ~x680 & ~x694 & ~x698 & ~x699 & ~x700 & ~x701 & ~x709 & ~x710 & ~x718 & ~x723 & ~x725 & ~x738 & ~x739 & ~x742 & ~x745 & ~x749 & ~x751 & ~x752 & ~x754 & ~x769 & ~x770 & ~x771 & ~x775 & ~x782;
assign c6137 =  x241 &  x298 &  x326 & ~x91 & ~x563 & ~x674 & ~x727;
assign c6139 =  x178 &  x661 & ~x93 & ~x363 & ~x679 & ~x727;
assign c6141 =  x152 & ~x18 & ~x62 & ~x114 & ~x116 & ~x220 & ~x223 & ~x225 & ~x254 & ~x282 & ~x287 & ~x291 & ~x304 & ~x316 & ~x334 & ~x341 & ~x343 & ~x344 & ~x346 & ~x372 & ~x392 & ~x741 & ~x744 & ~x769;
assign c6143 = ~x12 & ~x91 & ~x97 & ~x110 & ~x136 & ~x194 & ~x442 & ~x455 & ~x481 & ~x513 & ~x514 & ~x529 & ~x560 & ~x582 & ~x645 & ~x700 & ~x706 & ~x730 & ~x743 & ~x775;
assign c6145 =  x577 &  x628 & ~x9 & ~x25 & ~x30 & ~x36 & ~x106 & ~x113 & ~x118 & ~x163 & ~x278 & ~x396 & ~x404 & ~x405 & ~x408 & ~x461 & ~x462 & ~x464 & ~x489 & ~x531 & ~x645 & ~x673 & ~x679 & ~x734 & ~x764 & ~x778 & ~x780;
assign c6147 =  x376 & ~x2 & ~x5 & ~x8 & ~x34 & ~x35 & ~x40 & ~x48 & ~x49 & ~x60 & ~x65 & ~x68 & ~x69 & ~x72 & ~x77 & ~x78 & ~x85 & ~x86 & ~x88 & ~x91 & ~x106 & ~x116 & ~x254 & ~x282 & ~x386 & ~x392 & ~x415 & ~x451 & ~x458 & ~x460 & ~x461 & ~x476 & ~x478 & ~x530 & ~x531 & ~x583 & ~x590 & ~x639 & ~x699 & ~x706 & ~x720 & ~x765 & ~x772;
assign c6149 =  x622;
assign c6151 =  x434 & ~x2 & ~x9 & ~x27 & ~x29 & ~x34 & ~x61 & ~x77 & ~x80 & ~x86 & ~x103 & ~x115 & ~x137 & ~x143 & ~x144 & ~x172 & ~x200 & ~x249 & ~x370 & ~x385 & ~x386 & ~x393 & ~x413 & ~x421 & ~x436 & ~x438 & ~x439 & ~x440 & ~x454 & ~x465 & ~x470 & ~x473 & ~x494 & ~x505 & ~x506 & ~x532 & ~x555 & ~x640 & ~x643 & ~x664 & ~x673 & ~x687 & ~x688 & ~x701 & ~x721 & ~x723 & ~x727 & ~x763 & ~x765;
assign c6153 =  x327 &  x464 & ~x17 & ~x37 & ~x47 & ~x60 & ~x62 & ~x88 & ~x142 & ~x168 & ~x194 & ~x228 & ~x278 & ~x293 & ~x306 & ~x311 & ~x331 & ~x358 & ~x359 & ~x386 & ~x387 & ~x533 & ~x589 & ~x641 & ~x707 & ~x736 & ~x738 & ~x749 & ~x759;
assign c6155 =  x301 & ~x14 & ~x80 & ~x106 & ~x195 & ~x225 & ~x352 & ~x353 & ~x382 & ~x393 & ~x460 & ~x462 & ~x463 & ~x504 & ~x559 & ~x560 & ~x678 & ~x722 & ~x772;
assign c6157 =  x215 &  x243 &  x271 &  x355 & ~x21 & ~x51 & ~x59 & ~x83 & ~x672 & ~x690 & ~x767;
assign c6159 = ~x38 & ~x55 & ~x78 & ~x89 & ~x94 & ~x100 & ~x125 & ~x126 & ~x138 & ~x165 & ~x304 & ~x349 & ~x363 & ~x446 & ~x472 & ~x523 & ~x530 & ~x551 & ~x580 & ~x606 & ~x616 & ~x675 & ~x699 & ~x704 & ~x735 & ~x762 & ~x764 & ~x768 & ~x774;
assign c6161 = ~x2 & ~x3 & ~x9 & ~x20 & ~x53 & ~x59 & ~x63 & ~x79 & ~x81 & ~x84 & ~x87 & ~x111 & ~x114 & ~x133 & ~x201 & ~x223 & ~x226 & ~x228 & ~x229 & ~x250 & ~x350 & ~x351 & ~x406 & ~x407 & ~x408 & ~x409 & ~x419 & ~x433 & ~x434 & ~x436 & ~x437 & ~x445 & ~x447 & ~x448 & ~x451 & ~x463 & ~x473 & ~x488 & ~x490 & ~x583 & ~x590 & ~x670 & ~x671 & ~x677 & ~x695 & ~x722 & ~x724 & ~x729 & ~x730 & ~x746 & ~x750 & ~x751 & ~x753 & ~x758 & ~x779;
assign c6163 =  x299 &  x355 & ~x9 & ~x11 & ~x38 & ~x48 & ~x111 & ~x119 & ~x224 & ~x279 & ~x308 & ~x311 & ~x378 & ~x380 & ~x445 & ~x674 & ~x676 & ~x703 & ~x723 & ~x742;
assign c6165 =  x300 &  x328 &  x383 & ~x5 & ~x47 & ~x102 & ~x115 & ~x305 & ~x324 & ~x325 & ~x388 & ~x473 & ~x479 & ~x641 & ~x668 & ~x700 & ~x743 & ~x747;
assign c6167 =  x295 & ~x11 & ~x217 & ~x283 & ~x356 & ~x464 & ~x466 & ~x475 & ~x492 & ~x621 & ~x705;
assign c6169 = ~x0 & ~x4 & ~x20 & ~x29 & ~x33 & ~x43 & ~x51 & ~x54 & ~x61 & ~x70 & ~x71 & ~x72 & ~x89 & ~x91 & ~x102 & ~x165 & ~x166 & ~x197 & ~x279 & ~x335 & ~x358 & ~x360 & ~x426 & ~x444 & ~x446 & ~x447 & ~x451 & ~x452 & ~x455 & ~x485 & ~x486 & ~x500 & ~x506 & ~x532 & ~x586 & ~x591 & ~x649 & ~x666 & ~x679 & ~x694 & ~x701 & ~x710 & ~x712 & ~x727 & ~x746 & ~x777;
assign c6171 = ~x5 & ~x9 & ~x10 & ~x11 & ~x13 & ~x14 & ~x15 & ~x16 & ~x19 & ~x20 & ~x21 & ~x22 & ~x23 & ~x24 & ~x29 & ~x31 & ~x32 & ~x33 & ~x34 & ~x35 & ~x36 & ~x38 & ~x40 & ~x42 & ~x50 & ~x51 & ~x52 & ~x55 & ~x56 & ~x57 & ~x58 & ~x59 & ~x65 & ~x66 & ~x69 & ~x72 & ~x74 & ~x75 & ~x79 & ~x81 & ~x82 & ~x87 & ~x89 & ~x91 & ~x92 & ~x93 & ~x94 & ~x95 & ~x102 & ~x103 & ~x104 & ~x106 & ~x110 & ~x111 & ~x112 & ~x114 & ~x115 & ~x116 & ~x120 & ~x132 & ~x133 & ~x134 & ~x137 & ~x139 & ~x140 & ~x141 & ~x142 & ~x143 & ~x144 & ~x145 & ~x146 & ~x160 & ~x163 & ~x165 & ~x166 & ~x167 & ~x168 & ~x169 & ~x170 & ~x171 & ~x173 & ~x188 & ~x189 & ~x190 & ~x192 & ~x195 & ~x199 & ~x200 & ~x201 & ~x217 & ~x218 & ~x219 & ~x220 & ~x221 & ~x222 & ~x223 & ~x225 & ~x226 & ~x227 & ~x248 & ~x249 & ~x253 & ~x254 & ~x277 & ~x278 & ~x280 & ~x281 & ~x282 & ~x304 & ~x305 & ~x307 & ~x309 & ~x310 & ~x311 & ~x335 & ~x337 & ~x338 & ~x340 & ~x361 & ~x364 & ~x365 & ~x377 & ~x390 & ~x391 & ~x393 & ~x394 & ~x395 & ~x403 & ~x404 & ~x405 & ~x406 & ~x419 & ~x420 & ~x421 & ~x423 & ~x446 & ~x448 & ~x474 & ~x475 & ~x476 & ~x477 & ~x478 & ~x501 & ~x503 & ~x504 & ~x506 & ~x508 & ~x530 & ~x531 & ~x532 & ~x534 & ~x535 & ~x536 & ~x559 & ~x562 & ~x563 & ~x565 & ~x585 & ~x589 & ~x590 & ~x591 & ~x592 & ~x613 & ~x614 & ~x616 & ~x617 & ~x619 & ~x620 & ~x622 & ~x624 & ~x640 & ~x642 & ~x643 & ~x644 & ~x647 & ~x648 & ~x653 & ~x668 & ~x671 & ~x672 & ~x673 & ~x676 & ~x678 & ~x679 & ~x681 & ~x682 & ~x684 & ~x695 & ~x698 & ~x699 & ~x701 & ~x702 & ~x703 & ~x704 & ~x705 & ~x708 & ~x709 & ~x710 & ~x711 & ~x713 & ~x717 & ~x719 & ~x720 & ~x723 & ~x725 & ~x726 & ~x727 & ~x728 & ~x731 & ~x732 & ~x733 & ~x738 & ~x741 & ~x742 & ~x743 & ~x744 & ~x745 & ~x746 & ~x748 & ~x750 & ~x752 & ~x753 & ~x754 & ~x755 & ~x756 & ~x758 & ~x759 & ~x760 & ~x761 & ~x762 & ~x763 & ~x765 & ~x767 & ~x768 & ~x771 & ~x774 & ~x775 & ~x776 & ~x779 & ~x780 & ~x783;
assign c6173 =  x328 &  x541 & ~x12 & ~x56 & ~x81 & ~x85 & ~x87 & ~x164 & ~x193 & ~x225 & ~x352 & ~x433 & ~x463 & ~x654 & ~x679;
assign c6175 = ~x56 & ~x59 & ~x62 & ~x67 & ~x447 & ~x453 & ~x455 & ~x456 & ~x485 & ~x499 & ~x514 & ~x516 & ~x776;
assign c6177 = ~x2 & ~x5 & ~x12 & ~x33 & ~x34 & ~x35 & ~x41 & ~x46 & ~x51 & ~x68 & ~x77 & ~x83 & ~x91 & ~x92 & ~x93 & ~x97 & ~x104 & ~x132 & ~x137 & ~x142 & ~x166 & ~x224 & ~x278 & ~x281 & ~x360 & ~x392 & ~x422 & ~x450 & ~x531 & ~x539 & ~x540 & ~x542 & ~x544 & ~x564 & ~x571 & ~x588 & ~x618 & ~x641 & ~x645 & ~x672 & ~x674 & ~x677 & ~x680 & ~x727 & ~x759 & ~x765 & ~x768 & ~x779 & ~x780 & ~x783;
assign c6179 = ~x10 & ~x25 & ~x27 & ~x33 & ~x70 & ~x87 & ~x101 & ~x103 & ~x105 & ~x118 & ~x312 & ~x422 & ~x425 & ~x428 & ~x437 & ~x457 & ~x464 & ~x494 & ~x586 & ~x587 & ~x615 & ~x646 & ~x665 & ~x670 & ~x685 & ~x757;
assign c6181 =  x468 &  x495 & ~x18 & ~x40 & ~x78 & ~x106 & ~x144 & ~x168 & ~x169 & ~x381 & ~x409 & ~x502 & ~x582 & ~x591 & ~x612 & ~x671 & ~x689 & ~x705 & ~x726 & ~x739 & ~x741 & ~x743 & ~x747 & ~x757 & ~x768;
assign c6183 =  x206 &  x633 &  x660 & ~x38 & ~x93 & ~x101 & ~x391;
assign c6185 =  x508;
assign c6187 =  x181 & ~x6 & ~x12 & ~x13 & ~x26 & ~x30 & ~x36 & ~x46 & ~x49 & ~x54 & ~x57 & ~x59 & ~x73 & ~x75 & ~x76 & ~x79 & ~x85 & ~x86 & ~x87 & ~x98 & ~x112 & ~x133 & ~x135 & ~x142 & ~x161 & ~x196 & ~x226 & ~x247 & ~x253 & ~x256 & ~x273 & ~x277 & ~x302 & ~x308 & ~x316 & ~x318 & ~x330 & ~x345 & ~x358 & ~x364 & ~x391 & ~x395 & ~x396 & ~x419 & ~x441 & ~x448 & ~x476 & ~x478 & ~x480 & ~x504 & ~x507 & ~x535 & ~x560 & ~x561 & ~x563 & ~x564 & ~x586 & ~x587 & ~x588 & ~x590 & ~x649 & ~x673 & ~x677 & ~x679 & ~x705 & ~x706 & ~x709 & ~x713 & ~x730 & ~x740 & ~x743 & ~x745 & ~x750 & ~x753 & ~x755 & ~x767 & ~x772 & ~x777 & ~x778;
assign c6189 =  x234 &  x577 & ~x327 & ~x516 & ~x700;
assign c6191 = ~x7 & ~x11 & ~x13 & ~x17 & ~x26 & ~x31 & ~x41 & ~x44 & ~x46 & ~x47 & ~x50 & ~x51 & ~x59 & ~x65 & ~x66 & ~x72 & ~x74 & ~x76 & ~x80 & ~x83 & ~x91 & ~x95 & ~x98 & ~x107 & ~x110 & ~x111 & ~x112 & ~x114 & ~x115 & ~x119 & ~x120 & ~x122 & ~x167 & ~x171 & ~x193 & ~x194 & ~x200 & ~x201 & ~x221 & ~x225 & ~x250 & ~x255 & ~x277 & ~x279 & ~x301 & ~x304 & ~x308 & ~x310 & ~x336 & ~x337 & ~x338 & ~x341 & ~x363 & ~x393 & ~x397 & ~x418 & ~x425 & ~x472 & ~x476 & ~x479 & ~x505 & ~x508 & ~x525 & ~x528 & ~x532 & ~x535 & ~x565 & ~x571 & ~x591 & ~x617 & ~x619 & ~x620 & ~x626 & ~x641 & ~x652 & ~x671 & ~x674 & ~x676 & ~x677 & ~x679 & ~x693 & ~x694 & ~x696 & ~x698 & ~x699 & ~x709 & ~x712 & ~x720 & ~x729 & ~x730 & ~x751 & ~x757 & ~x758 & ~x767 & ~x770 & ~x773 & ~x775 & ~x781;
assign c6193 =  x268 & ~x13 & ~x17 & ~x18 & ~x19 & ~x24 & ~x26 & ~x42 & ~x79 & ~x95 & ~x101 & ~x103 & ~x105 & ~x138 & ~x144 & ~x161 & ~x162 & ~x278 & ~x283 & ~x310 & ~x364 & ~x387 & ~x503 & ~x518 & ~x589 & ~x639 & ~x646 & ~x665 & ~x667 & ~x675 & ~x696 & ~x698 & ~x704 & ~x706 & ~x727 & ~x732 & ~x744 & ~x751 & ~x764 & ~x767 & ~x779;
assign c6195 =  x212 &  x268 &  x297 & ~x0 & ~x14 & ~x26 & ~x29 & ~x55 & ~x56 & ~x100 & ~x102 & ~x104 & ~x132 & ~x170 & ~x282 & ~x333 & ~x528 & ~x533 & ~x591 & ~x643 & ~x675 & ~x726 & ~x728 & ~x730;
assign c6197 =  x328 &  x384 & ~x19 & ~x31 & ~x37 & ~x118 & ~x136 & ~x141 & ~x145 & ~x170 & ~x227 & ~x278 & ~x351 & ~x420 & ~x443 & ~x476 & ~x560 & ~x672 & ~x675 & ~x691 & ~x722 & ~x737 & ~x741 & ~x743 & ~x759 & ~x766;
assign c6199 = ~x61 & ~x68 & ~x81 & ~x100 & ~x306 & ~x511 & ~x514 & ~x516 & ~x531 & ~x541 & ~x588 & ~x737;
assign c6201 =  x432 &  x435 &  x458 & ~x6 & ~x9 & ~x12 & ~x25 & ~x50 & ~x66 & ~x79 & ~x100 & ~x108 & ~x137 & ~x142 & ~x164 & ~x197 & ~x199 & ~x230 & ~x287 & ~x306 & ~x309 & ~x364 & ~x369 & ~x419 & ~x470 & ~x479 & ~x501 & ~x534 & ~x551 & ~x555 & ~x563 & ~x583 & ~x588 & ~x590 & ~x614 & ~x638 & ~x640 & ~x641 & ~x648 & ~x720 & ~x739 & ~x752 & ~x758 & ~x771;
assign c6203 =  x567 & ~x0 & ~x7 & ~x27 & ~x28 & ~x37 & ~x39 & ~x48 & ~x51 & ~x60 & ~x66 & ~x76 & ~x77 & ~x79 & ~x83 & ~x86 & ~x107 & ~x108 & ~x110 & ~x138 & ~x143 & ~x145 & ~x197 & ~x199 & ~x220 & ~x225 & ~x248 & ~x286 & ~x312 & ~x314 & ~x315 & ~x338 & ~x341 & ~x364 & ~x392 & ~x400 & ~x413 & ~x417 & ~x420 & ~x421 & ~x475 & ~x506 & ~x531 & ~x533 & ~x586 & ~x616 & ~x644 & ~x648 & ~x675 & ~x691 & ~x697 & ~x706 & ~x719 & ~x726 & ~x729 & ~x730 & ~x734 & ~x736 & ~x737 & ~x748 & ~x760 & ~x766 & ~x769 & ~x772 & ~x779 & ~x781;
assign c6205 =  x239 & ~x4 & ~x7 & ~x13 & ~x25 & ~x41 & ~x47 & ~x51 & ~x60 & ~x76 & ~x78 & ~x84 & ~x99 & ~x103 & ~x104 & ~x105 & ~x106 & ~x107 & ~x128 & ~x133 & ~x136 & ~x137 & ~x157 & ~x158 & ~x252 & ~x274 & ~x328 & ~x365 & ~x394 & ~x417 & ~x420 & ~x445 & ~x502 & ~x536 & ~x588 & ~x593 & ~x619 & ~x640 & ~x666 & ~x670 & ~x671 & ~x673 & ~x675 & ~x678 & ~x681 & ~x689 & ~x690 & ~x691 & ~x693 & ~x702 & ~x706 & ~x718 & ~x720 & ~x724 & ~x730 & ~x737 & ~x743 & ~x745 & ~x746 & ~x770 & ~x779 & ~x781;
assign c6207 = ~x15 & ~x16 & ~x34 & ~x71 & ~x73 & ~x75 & ~x113 & ~x114 & ~x127 & ~x129 & ~x172 & ~x256 & ~x348 & ~x349 & ~x360 & ~x414 & ~x415 & ~x449 & ~x559 & ~x562 & ~x573 & ~x591 & ~x600 & ~x697 & ~x743 & ~x751 & ~x783;
assign c6209 = ~x15 & ~x21 & ~x25 & ~x31 & ~x33 & ~x38 & ~x89 & ~x90 & ~x91 & ~x101 & ~x104 & ~x107 & ~x109 & ~x132 & ~x134 & ~x137 & ~x140 & ~x158 & ~x160 & ~x169 & ~x172 & ~x189 & ~x198 & ~x214 & ~x217 & ~x222 & ~x244 & ~x247 & ~x253 & ~x255 & ~x256 & ~x278 & ~x305 & ~x330 & ~x331 & ~x337 & ~x338 & ~x340 & ~x341 & ~x358 & ~x363 & ~x364 & ~x383 & ~x387 & ~x392 & ~x394 & ~x411 & ~x412 & ~x413 & ~x438 & ~x448 & ~x478 & ~x479 & ~x507 & ~x508 & ~x533 & ~x537 & ~x565 & ~x620 & ~x624 & ~x645 & ~x679 & ~x684 & ~x699 & ~x702 & ~x703 & ~x713 & ~x720 & ~x726 & ~x745 & ~x747 & ~x749 & ~x752 & ~x759 & ~x762 & ~x763 & ~x770;
assign c6211 =  x238 &  x380 & ~x29 & ~x33 & ~x96 & ~x98 & ~x114 & ~x127 & ~x130 & ~x156 & ~x620 & ~x705;
assign c6213 =  x456 & ~x38 & ~x74 & ~x79 & ~x96 & ~x121 & ~x125 & ~x127 & ~x149 & ~x154 & ~x155 & ~x173 & ~x201 & ~x225 & ~x309 & ~x418 & ~x502 & ~x504 & ~x505 & ~x560 & ~x566 & ~x569 & ~x595 & ~x624 & ~x741 & ~x755 & ~x756 & ~x758 & ~x765 & ~x769 & ~x770;
assign c6215 = ~x129 & ~x130 & ~x227 & ~x500 & ~x547 & ~x572 & ~x573 & ~x574;
assign c6217 =  x654 & ~x34 & ~x41 & ~x69 & ~x70 & ~x73 & ~x77 & ~x85 & ~x103 & ~x135 & ~x195 & ~x283 & ~x365 & ~x448 & ~x451 & ~x556 & ~x606 & ~x727 & ~x739 & ~x780;
assign c6219 =  x269 & ~x35 & ~x40 & ~x43 & ~x44 & ~x68 & ~x75 & ~x78 & ~x135 & ~x163 & ~x164 & ~x226 & ~x275 & ~x301 & ~x363 & ~x423 & ~x559 & ~x575 & ~x619 & ~x697 & ~x709 & ~x750 & ~x769;
assign c6221 =  x295 & ~x27 & ~x74 & ~x88 & ~x158 & ~x161 & ~x169 & ~x298 & ~x301 & ~x327 & ~x372 & ~x374 & ~x448 & ~x668 & ~x680 & ~x708 & ~x728;
assign c6223 =  x406 & ~x6 & ~x7 & ~x8 & ~x10 & ~x18 & ~x19 & ~x20 & ~x25 & ~x34 & ~x37 & ~x38 & ~x41 & ~x48 & ~x49 & ~x51 & ~x52 & ~x53 & ~x57 & ~x64 & ~x67 & ~x76 & ~x78 & ~x83 & ~x88 & ~x100 & ~x105 & ~x110 & ~x115 & ~x135 & ~x140 & ~x144 & ~x164 & ~x166 & ~x190 & ~x191 & ~x196 & ~x197 & ~x199 & ~x225 & ~x228 & ~x253 & ~x279 & ~x307 & ~x309 & ~x310 & ~x313 & ~x328 & ~x337 & ~x340 & ~x341 & ~x342 & ~x355 & ~x361 & ~x365 & ~x382 & ~x383 & ~x387 & ~x394 & ~x397 & ~x399 & ~x400 & ~x410 & ~x412 & ~x414 & ~x417 & ~x420 & ~x428 & ~x443 & ~x450 & ~x452 & ~x469 & ~x470 & ~x471 & ~x474 & ~x480 & ~x505 & ~x506 & ~x563 & ~x589 & ~x622 & ~x649 & ~x650 & ~x668 & ~x695 & ~x702 & ~x703 & ~x707 & ~x719 & ~x723 & ~x725 & ~x731 & ~x736 & ~x742 & ~x743 & ~x744 & ~x754 & ~x757 & ~x759 & ~x761 & ~x763 & ~x769 & ~x771 & ~x772 & ~x782;
assign c6225 =  x269 & ~x8 & ~x9 & ~x11 & ~x17 & ~x20 & ~x30 & ~x33 & ~x41 & ~x44 & ~x60 & ~x62 & ~x68 & ~x76 & ~x92 & ~x110 & ~x112 & ~x113 & ~x116 & ~x142 & ~x160 & ~x161 & ~x168 & ~x171 & ~x189 & ~x199 & ~x226 & ~x278 & ~x279 & ~x312 & ~x329 & ~x335 & ~x337 & ~x356 & ~x368 & ~x386 & ~x417 & ~x419 & ~x421 & ~x422 & ~x444 & ~x451 & ~x530 & ~x533 & ~x587 & ~x614 & ~x623 & ~x666 & ~x674 & ~x677 & ~x697 & ~x698 & ~x705 & ~x709 & ~x711 & ~x724 & ~x725 & ~x728 & ~x743 & ~x750 & ~x761;
assign c6227 =  x217 & ~x5 & ~x9 & ~x23 & ~x24 & ~x35 & ~x38 & ~x39 & ~x45 & ~x61 & ~x83 & ~x89 & ~x94 & ~x106 & ~x119 & ~x120 & ~x144 & ~x145 & ~x167 & ~x250 & ~x280 & ~x283 & ~x296 & ~x305 & ~x306 & ~x307 & ~x308 & ~x339 & ~x446 & ~x528 & ~x557 & ~x561 & ~x585 & ~x587 & ~x588 & ~x614 & ~x618 & ~x658 & ~x659 & ~x699 & ~x701 & ~x728 & ~x729 & ~x737 & ~x747 & ~x748 & ~x749 & ~x751 & ~x769 & ~x777;
assign c6229 = ~x7 & ~x25 & ~x30 & ~x36 & ~x38 & ~x49 & ~x51 & ~x52 & ~x60 & ~x62 & ~x66 & ~x76 & ~x79 & ~x88 & ~x97 & ~x104 & ~x106 & ~x142 & ~x162 & ~x198 & ~x227 & ~x252 & ~x306 & ~x310 & ~x335 & ~x337 & ~x339 & ~x359 & ~x360 & ~x364 & ~x445 & ~x448 & ~x449 & ~x452 & ~x500 & ~x506 & ~x507 & ~x532 & ~x534 & ~x536 & ~x559 & ~x563 & ~x564 & ~x571 & ~x572 & ~x573 & ~x591 & ~x595 & ~x599 & ~x617 & ~x623 & ~x644 & ~x650 & ~x653 & ~x702 & ~x704 & ~x737 & ~x740 & ~x741 & ~x742 & ~x753 & ~x754;
assign c6231 = ~x3 & ~x9 & ~x30 & ~x42 & ~x45 & ~x48 & ~x56 & ~x66 & ~x70 & ~x80 & ~x82 & ~x97 & ~x99 & ~x102 & ~x103 & ~x120 & ~x122 & ~x124 & ~x135 & ~x137 & ~x145 & ~x152 & ~x197 & ~x199 & ~x223 & ~x339 & ~x363 & ~x392 & ~x394 & ~x418 & ~x473 & ~x475 & ~x496 & ~x497 & ~x520 & ~x521 & ~x523 & ~x524 & ~x530 & ~x533 & ~x552 & ~x560 & ~x561 & ~x579 & ~x604 & ~x632 & ~x634 & ~x638 & ~x640 & ~x659 & ~x671 & ~x678 & ~x711 & ~x725 & ~x732 & ~x754 & ~x760 & ~x764;
assign c6233 =  x568 & ~x81 & ~x351 & ~x352 & ~x378 & ~x405 & ~x408 & ~x461 & ~x464 & ~x490 & ~x491 & ~x779;
assign c6235 = ~x22 & ~x64 & ~x70 & ~x75 & ~x93 & ~x126 & ~x159 & ~x167 & ~x225 & ~x249 & ~x364 & ~x366 & ~x390 & ~x477 & ~x480 & ~x506 & ~x512 & ~x517 & ~x564 & ~x615 & ~x697 & ~x721 & ~x741 & ~x743 & ~x749 & ~x753 & ~x773;
assign c6237 = ~x6 & ~x7 & ~x54 & ~x65 & ~x72 & ~x73 & ~x90 & ~x94 & ~x97 & ~x100 & ~x140 & ~x142 & ~x144 & ~x180 & ~x194 & ~x201 & ~x252 & ~x309 & ~x416 & ~x446 & ~x535 & ~x539 & ~x542 & ~x543 & ~x561 & ~x563 & ~x645 & ~x668 & ~x704 & ~x755 & ~x766;
assign c6239 =  x570 & ~x24 & ~x33 & ~x76 & ~x77 & ~x109 & ~x143 & ~x164 & ~x232 & ~x285 & ~x310 & ~x361 & ~x413 & ~x468 & ~x476 & ~x486 & ~x620 & ~x657 & ~x717 & ~x722;
assign c6241 =  x245 &  x273 &  x355 & ~x23 & ~x29 & ~x41 & ~x59 & ~x69 & ~x73 & ~x97 & ~x197 & ~x253 & ~x446 & ~x590 & ~x615 & ~x672 & ~x721 & ~x741 & ~x748 & ~x755 & ~x759;
assign c6243 = ~x3 & ~x15 & ~x43 & ~x58 & ~x81 & ~x110 & ~x111 & ~x112 & ~x114 & ~x121 & ~x148 & ~x150 & ~x175 & ~x227 & ~x284 & ~x286 & ~x288 & ~x394 & ~x429 & ~x442 & ~x459 & ~x460 & ~x473 & ~x475 & ~x558 & ~x560 & ~x561 & ~x585 & ~x614 & ~x703 & ~x708 & ~x713 & ~x757 & ~x766 & ~x770 & ~x776 & ~x781;
assign c6245 = ~x0 & ~x1 & ~x6 & ~x8 & ~x10 & ~x18 & ~x27 & ~x28 & ~x32 & ~x43 & ~x47 & ~x55 & ~x57 & ~x60 & ~x65 & ~x77 & ~x78 & ~x87 & ~x92 & ~x108 & ~x136 & ~x143 & ~x165 & ~x171 & ~x173 & ~x192 & ~x194 & ~x200 & ~x201 & ~x251 & ~x310 & ~x360 & ~x365 & ~x367 & ~x368 & ~x388 & ~x416 & ~x419 & ~x421 & ~x422 & ~x423 & ~x445 & ~x446 & ~x450 & ~x451 & ~x472 & ~x478 & ~x547 & ~x556 & ~x558 & ~x561 & ~x562 & ~x587 & ~x589 & ~x602 & ~x615 & ~x617 & ~x618 & ~x619 & ~x630 & ~x631 & ~x645 & ~x650 & ~x670 & ~x672 & ~x674 & ~x678 & ~x679 & ~x681 & ~x694 & ~x698 & ~x702 & ~x705 & ~x709 & ~x726 & ~x728 & ~x731 & ~x735 & ~x736 & ~x738 & ~x739 & ~x740 & ~x746 & ~x753 & ~x755 & ~x762 & ~x763 & ~x764 & ~x765 & ~x766 & ~x775 & ~x777 & ~x783;
assign c6247 =  x213 & ~x15 & ~x16 & ~x18 & ~x24 & ~x48 & ~x51 & ~x63 & ~x75 & ~x77 & ~x85 & ~x89 & ~x90 & ~x93 & ~x101 & ~x102 & ~x104 & ~x120 & ~x133 & ~x199 & ~x200 & ~x201 & ~x222 & ~x252 & ~x253 & ~x279 & ~x309 & ~x311 & ~x312 & ~x335 & ~x337 & ~x338 & ~x339 & ~x362 & ~x363 & ~x364 & ~x390 & ~x419 & ~x424 & ~x448 & ~x489 & ~x532 & ~x558 & ~x564 & ~x585 & ~x637 & ~x642 & ~x665 & ~x667 & ~x686 & ~x692 & ~x696 & ~x700 & ~x730 & ~x735 & ~x739 & ~x742 & ~x747 & ~x764 & ~x767 & ~x771 & ~x772 & ~x777 & ~x780;
assign c6249 = ~x57 & ~x77 & ~x84 & ~x94 & ~x110 & ~x116 & ~x119 & ~x123 & ~x172 & ~x175 & ~x201 & ~x220 & ~x225 & ~x228 & ~x281 & ~x388 & ~x421 & ~x443 & ~x474 & ~x478 & ~x570 & ~x587 & ~x598 & ~x600 & ~x633 & ~x655 & ~x700 & ~x708 & ~x722 & ~x736 & ~x739 & ~x741 & ~x761 & ~x765;
assign c6251 =  x187 &  x215 &  x271 & ~x630;
assign c6253 =  x461 &  x462 & ~x68 & ~x70 & ~x94 & ~x113 & ~x117 & ~x543 & ~x570 & ~x590 & ~x699 & ~x727;
assign c6255 = ~x0 & ~x1 & ~x8 & ~x11 & ~x15 & ~x16 & ~x17 & ~x21 & ~x24 & ~x26 & ~x29 & ~x31 & ~x33 & ~x34 & ~x35 & ~x40 & ~x42 & ~x57 & ~x66 & ~x67 & ~x78 & ~x80 & ~x81 & ~x91 & ~x103 & ~x108 & ~x109 & ~x112 & ~x115 & ~x132 & ~x137 & ~x138 & ~x139 & ~x140 & ~x142 & ~x144 & ~x160 & ~x161 & ~x164 & ~x167 & ~x168 & ~x169 & ~x172 & ~x193 & ~x195 & ~x196 & ~x202 & ~x223 & ~x226 & ~x252 & ~x254 & ~x281 & ~x331 & ~x334 & ~x337 & ~x356 & ~x357 & ~x360 & ~x361 & ~x384 & ~x386 & ~x391 & ~x393 & ~x395 & ~x411 & ~x412 & ~x414 & ~x422 & ~x425 & ~x451 & ~x452 & ~x477 & ~x478 & ~x479 & ~x502 & ~x504 & ~x508 & ~x529 & ~x532 & ~x560 & ~x587 & ~x588 & ~x589 & ~x593 & ~x612 & ~x616 & ~x618 & ~x636 & ~x643 & ~x650 & ~x651 & ~x656 & ~x657 & ~x658 & ~x669 & ~x693 & ~x694 & ~x695 & ~x696 & ~x697 & ~x700 & ~x705 & ~x707 & ~x720 & ~x725 & ~x728 & ~x729 & ~x730 & ~x732 & ~x738 & ~x739 & ~x740 & ~x745 & ~x748 & ~x753 & ~x754 & ~x762 & ~x763 & ~x777 & ~x780 & ~x781;
assign c6257 =  x577 &  x598 & ~x13 & ~x17 & ~x34 & ~x51 & ~x58 & ~x61 & ~x66 & ~x67 & ~x70 & ~x76 & ~x83 & ~x89 & ~x93 & ~x104 & ~x112 & ~x117 & ~x173 & ~x199 & ~x278 & ~x284 & ~x308 & ~x312 & ~x361 & ~x363 & ~x365 & ~x436 & ~x460 & ~x464 & ~x473 & ~x474 & ~x486 & ~x487 & ~x489 & ~x490 & ~x530 & ~x532 & ~x559 & ~x560 & ~x585 & ~x587 & ~x589 & ~x590 & ~x591 & ~x611 & ~x619 & ~x620 & ~x639 & ~x647 & ~x666 & ~x667 & ~x670 & ~x685 & ~x695 & ~x700 & ~x702 & ~x708 & ~x718 & ~x723 & ~x729 & ~x734 & ~x735 & ~x745 & ~x749 & ~x752 & ~x761 & ~x762 & ~x765 & ~x782;
assign c6259 =  x653 & ~x138 & ~x166;
assign c6261 =  x185 &  x351 & ~x22 & ~x26 & ~x69 & ~x103 & ~x105 & ~x111 & ~x225 & ~x254 & ~x340 & ~x401 & ~x706 & ~x735 & ~x766;
assign c6263 =  x181 &  x654 & ~x47 & ~x100 & ~x367 & ~x425 & ~x724;
assign c6265 = ~x2 & ~x4 & ~x5 & ~x10 & ~x16 & ~x33 & ~x34 & ~x35 & ~x37 & ~x44 & ~x45 & ~x53 & ~x59 & ~x63 & ~x66 & ~x76 & ~x77 & ~x89 & ~x95 & ~x97 & ~x100 & ~x101 & ~x105 & ~x122 & ~x126 & ~x127 & ~x130 & ~x131 & ~x133 & ~x137 & ~x140 & ~x163 & ~x169 & ~x170 & ~x171 & ~x172 & ~x175 & ~x177 & ~x195 & ~x227 & ~x231 & ~x255 & ~x257 & ~x287 & ~x336 & ~x364 & ~x390 & ~x474 & ~x499 & ~x501 & ~x507 & ~x523 & ~x526 & ~x552 & ~x554 & ~x555 & ~x557 & ~x563 & ~x578 & ~x580 & ~x583 & ~x586 & ~x607 & ~x608 & ~x615 & ~x619 & ~x621 & ~x635 & ~x647 & ~x677 & ~x704 & ~x722 & ~x723 & ~x724 & ~x729 & ~x733 & ~x743 & ~x750 & ~x766 & ~x775 & ~x776;
assign c6267 =  x540 & ~x0 & ~x2 & ~x6 & ~x10 & ~x11 & ~x13 & ~x23 & ~x24 & ~x25 & ~x26 & ~x32 & ~x35 & ~x39 & ~x45 & ~x51 & ~x54 & ~x58 & ~x74 & ~x85 & ~x86 & ~x88 & ~x108 & ~x109 & ~x114 & ~x134 & ~x136 & ~x138 & ~x139 & ~x141 & ~x163 & ~x165 & ~x166 & ~x169 & ~x173 & ~x199 & ~x223 & ~x226 & ~x246 & ~x248 & ~x251 & ~x252 & ~x277 & ~x279 & ~x307 & ~x310 & ~x311 & ~x314 & ~x338 & ~x340 & ~x360 & ~x363 & ~x368 & ~x369 & ~x370 & ~x372 & ~x395 & ~x399 & ~x401 & ~x416 & ~x420 & ~x422 & ~x424 & ~x426 & ~x447 & ~x452 & ~x478 & ~x502 & ~x504 & ~x560 & ~x589 & ~x613 & ~x640 & ~x642 & ~x643 & ~x671 & ~x672 & ~x673 & ~x675 & ~x676 & ~x677 & ~x680 & ~x682 & ~x686 & ~x688 & ~x693 & ~x694 & ~x702 & ~x704 & ~x710 & ~x714 & ~x733 & ~x740 & ~x746 & ~x752 & ~x757 & ~x758 & ~x759 & ~x763 & ~x764 & ~x770 & ~x772 & ~x776 & ~x779 & ~x781 & ~x783;
assign c6269 =  x326 &  x354 & ~x8 & ~x21 & ~x22 & ~x27 & ~x32 & ~x39 & ~x43 & ~x50 & ~x52 & ~x54 & ~x57 & ~x61 & ~x66 & ~x67 & ~x70 & ~x89 & ~x99 & ~x107 & ~x109 & ~x110 & ~x195 & ~x197 & ~x198 & ~x223 & ~x224 & ~x227 & ~x249 & ~x283 & ~x284 & ~x305 & ~x307 & ~x323 & ~x339 & ~x360 & ~x363 & ~x367 & ~x385 & ~x414 & ~x415 & ~x417 & ~x421 & ~x474 & ~x479 & ~x499 & ~x501 & ~x505 & ~x529 & ~x530 & ~x531 & ~x557 & ~x587 & ~x644 & ~x648 & ~x676 & ~x682 & ~x706 & ~x708 & ~x714 & ~x721 & ~x729 & ~x733 & ~x736 & ~x737 & ~x739 & ~x743 & ~x757 & ~x778;
assign c6271 =  x269 &  x297 &  x325 &  x409 & ~x13 & ~x103 & ~x274 & ~x644 & ~x783;
assign c6273 =  x127 &  x159;
assign c6275 =  x274 &  x302 & ~x15 & ~x19 & ~x21 & ~x24 & ~x25 & ~x32 & ~x38 & ~x48 & ~x51 & ~x55 & ~x60 & ~x69 & ~x86 & ~x136 & ~x146 & ~x174 & ~x175 & ~x200 & ~x225 & ~x252 & ~x255 & ~x256 & ~x284 & ~x306 & ~x309 & ~x336 & ~x352 & ~x353 & ~x367 & ~x389 & ~x394 & ~x422 & ~x445 & ~x449 & ~x450 & ~x475 & ~x528 & ~x531 & ~x535 & ~x556 & ~x560 & ~x614 & ~x672 & ~x687 & ~x708 & ~x722 & ~x729 & ~x760 & ~x770 & ~x773 & ~x775 & ~x777 & ~x782;
assign c6277 =  x749;
assign c6279 = ~x1 & ~x20 & ~x67 & ~x104 & ~x222 & ~x337 & ~x419 & ~x510 & ~x516 & ~x533 & ~x541 & ~x543 & ~x620 & ~x731 & ~x760 & ~x779;
assign c6281 =  x242 & ~x11 & ~x13 & ~x18 & ~x21 & ~x30 & ~x34 & ~x35 & ~x36 & ~x45 & ~x56 & ~x57 & ~x62 & ~x66 & ~x73 & ~x75 & ~x77 & ~x81 & ~x84 & ~x85 & ~x89 & ~x92 & ~x104 & ~x106 & ~x110 & ~x111 & ~x116 & ~x119 & ~x120 & ~x122 & ~x135 & ~x136 & ~x137 & ~x141 & ~x143 & ~x145 & ~x147 & ~x161 & ~x163 & ~x164 & ~x165 & ~x168 & ~x169 & ~x175 & ~x177 & ~x194 & ~x201 & ~x223 & ~x225 & ~x226 & ~x251 & ~x257 & ~x310 & ~x311 & ~x335 & ~x336 & ~x368 & ~x424 & ~x447 & ~x448 & ~x450 & ~x474 & ~x477 & ~x481 & ~x496 & ~x497 & ~x507 & ~x523 & ~x525 & ~x529 & ~x532 & ~x558 & ~x562 & ~x565 & ~x592 & ~x612 & ~x616 & ~x617 & ~x639 & ~x640 & ~x649 & ~x675 & ~x676 & ~x694 & ~x700 & ~x705 & ~x728 & ~x740 & ~x743 & ~x751 & ~x759 & ~x762 & ~x774 & ~x775 & ~x778 & ~x781 & ~x783;
assign c6283 =  x328 & ~x5 & ~x20 & ~x22 & ~x30 & ~x32 & ~x47 & ~x55 & ~x58 & ~x60 & ~x62 & ~x65 & ~x67 & ~x68 & ~x77 & ~x79 & ~x83 & ~x93 & ~x94 & ~x96 & ~x121 & ~x190 & ~x196 & ~x198 & ~x199 & ~x252 & ~x307 & ~x361 & ~x378 & ~x407 & ~x408 & ~x434 & ~x435 & ~x476 & ~x534 & ~x587 & ~x590 & ~x614 & ~x640 & ~x642 & ~x643 & ~x651 & ~x670 & ~x676 & ~x698 & ~x703 & ~x735 & ~x736 & ~x748 & ~x749 & ~x750 & ~x751 & ~x760 & ~x763 & ~x768 & ~x772 & ~x776 & ~x779;
assign c6285 =  x154 & ~x12 & ~x14 & ~x21 & ~x41 & ~x50 & ~x74 & ~x111 & ~x138 & ~x143 & ~x226 & ~x255 & ~x256 & ~x257 & ~x280 & ~x281 & ~x287 & ~x303 & ~x347 & ~x363 & ~x372 & ~x398 & ~x450 & ~x557 & ~x589 & ~x694 & ~x711 & ~x749 & ~x772;
assign c6287 =  x289 &  x656 & ~x12 & ~x13 & ~x18 & ~x30 & ~x32 & ~x38 & ~x49 & ~x60 & ~x69 & ~x70 & ~x71 & ~x79 & ~x91 & ~x92 & ~x93 & ~x98 & ~x101 & ~x102 & ~x147 & ~x200 & ~x201 & ~x202 & ~x229 & ~x279 & ~x281 & ~x306 & ~x336 & ~x338 & ~x364 & ~x421 & ~x455 & ~x480 & ~x504 & ~x506 & ~x537 & ~x591 & ~x593 & ~x613 & ~x642 & ~x644 & ~x666 & ~x678 & ~x705 & ~x722 & ~x728 & ~x732 & ~x739 & ~x772 & ~x776 & ~x777 & ~x781;
assign c6289 =  x151 & ~x0 & ~x8 & ~x11 & ~x24 & ~x56 & ~x70 & ~x77 & ~x131 & ~x304 & ~x339 & ~x367 & ~x426 & ~x427 & ~x429 & ~x474 & ~x475 & ~x476 & ~x686 & ~x692 & ~x696 & ~x752 & ~x758 & ~x766 & ~x767 & ~x779 & ~x781;
assign c6291 =  x185 & ~x458 & ~x488;
assign c6293 =  x233 & ~x457 & ~x482 & ~x483 & ~x484 & ~x512;
assign c6295 =  x402 & ~x11 & ~x23 & ~x29 & ~x53 & ~x58 & ~x67 & ~x70 & ~x74 & ~x85 & ~x106 & ~x112 & ~x137 & ~x281 & ~x332 & ~x333 & ~x335 & ~x365 & ~x389 & ~x421 & ~x423 & ~x472 & ~x475 & ~x476 & ~x486 & ~x488 & ~x513 & ~x677 & ~x698 & ~x704 & ~x707 & ~x720 & ~x759 & ~x775;
assign c6297 =  x298 & ~x320 & ~x321 & ~x442;
assign c6299 =  x299 &  x354 & ~x3 & ~x5 & ~x17 & ~x20 & ~x43 & ~x59 & ~x66 & ~x73 & ~x74 & ~x79 & ~x84 & ~x90 & ~x94 & ~x97 & ~x99 & ~x112 & ~x139 & ~x143 & ~x167 & ~x221 & ~x226 & ~x255 & ~x279 & ~x281 & ~x305 & ~x330 & ~x335 & ~x336 & ~x357 & ~x362 & ~x387 & ~x389 & ~x416 & ~x418 & ~x448 & ~x477 & ~x478 & ~x504 & ~x587 & ~x616 & ~x618 & ~x620 & ~x649 & ~x670 & ~x697 & ~x709 & ~x712 & ~x713 & ~x717 & ~x736 & ~x741 & ~x742 & ~x747 & ~x760 & ~x766 & ~x768 & ~x772 & ~x779 & ~x780;
assign c70 =  x231 &  x265 &  x266 &  x492 &  x520 &  x547 & ~x5 & ~x12 & ~x17 & ~x33 & ~x42 & ~x61 & ~x68 & ~x80 & ~x95 & ~x97 & ~x118 & ~x154 & ~x193 & ~x221 & ~x250 & ~x309 & ~x339 & ~x362 & ~x390 & ~x393 & ~x395 & ~x421 & ~x473 & ~x477 & ~x500 & ~x504 & ~x510 & ~x527 & ~x528 & ~x532 & ~x539 & ~x559 & ~x565 & ~x567 & ~x591 & ~x616 & ~x621 & ~x622 & ~x671 & ~x672 & ~x696 & ~x700 & ~x735 & ~x760 & ~x779;
assign c72 = ~x12 & ~x23 & ~x33 & ~x48 & ~x55 & ~x74 & ~x77 & ~x83 & ~x90 & ~x91 & ~x102 & ~x110 & ~x112 & ~x122 & ~x124 & ~x126 & ~x138 & ~x144 & ~x145 & ~x156 & ~x161 & ~x176 & ~x178 & ~x200 & ~x281 & ~x307 & ~x334 & ~x350 & ~x360 & ~x363 & ~x377 & ~x386 & ~x387 & ~x397 & ~x415 & ~x416 & ~x433 & ~x440 & ~x446 & ~x451 & ~x453 & ~x459 & ~x468 & ~x471 & ~x472 & ~x477 & ~x486 & ~x498 & ~x506 & ~x512 & ~x526 & ~x529 & ~x531 & ~x537 & ~x565 & ~x567 & ~x589 & ~x591 & ~x594 & ~x605 & ~x620 & ~x636 & ~x662 & ~x670 & ~x672 & ~x696 & ~x700 & ~x702 & ~x721 & ~x726 & ~x729 & ~x732 & ~x735 & ~x744 & ~x748 & ~x762 & ~x764 & ~x769 & ~x783;
assign c74 =  x206 &  x464 &  x574 &  x602 & ~x7 & ~x24 & ~x25 & ~x28 & ~x32 & ~x35 & ~x39 & ~x42 & ~x56 & ~x57 & ~x62 & ~x67 & ~x71 & ~x73 & ~x77 & ~x92 & ~x94 & ~x96 & ~x97 & ~x103 & ~x104 & ~x105 & ~x107 & ~x112 & ~x114 & ~x118 & ~x119 & ~x122 & ~x123 & ~x124 & ~x125 & ~x128 & ~x148 & ~x153 & ~x163 & ~x167 & ~x169 & ~x170 & ~x197 & ~x228 & ~x279 & ~x309 & ~x333 & ~x348 & ~x349 & ~x359 & ~x360 & ~x362 & ~x365 & ~x367 & ~x389 & ~x391 & ~x392 & ~x394 & ~x416 & ~x420 & ~x424 & ~x447 & ~x474 & ~x501 & ~x502 & ~x508 & ~x531 & ~x533 & ~x554 & ~x562 & ~x565 & ~x579 & ~x581 & ~x582 & ~x592 & ~x597 & ~x607 & ~x611 & ~x616 & ~x619 & ~x620 & ~x623 & ~x633 & ~x634 & ~x638 & ~x639 & ~x644 & ~x647 & ~x649 & ~x652 & ~x653 & ~x662 & ~x674 & ~x681 & ~x701 & ~x703 & ~x716 & ~x719 & ~x725 & ~x726 & ~x731 & ~x734 & ~x739 & ~x748 & ~x749 & ~x750 & ~x752 & ~x762 & ~x773 & ~x775 & ~x777;
assign c76 =  x300 & ~x184 & ~x456 & ~x604 & ~x658 & ~x659;
assign c78 =  x238 &  x464 &  x492 &  x576 &  x632 & ~x15 & ~x22 & ~x23 & ~x24 & ~x25 & ~x28 & ~x38 & ~x39 & ~x44 & ~x45 & ~x49 & ~x53 & ~x59 & ~x87 & ~x100 & ~x110 & ~x111 & ~x118 & ~x120 & ~x121 & ~x126 & ~x128 & ~x135 & ~x142 & ~x154 & ~x155 & ~x161 & ~x162 & ~x166 & ~x223 & ~x226 & ~x245 & ~x250 & ~x273 & ~x300 & ~x308 & ~x328 & ~x331 & ~x333 & ~x348 & ~x356 & ~x362 & ~x376 & ~x384 & ~x385 & ~x390 & ~x391 & ~x396 & ~x416 & ~x417 & ~x419 & ~x425 & ~x448 & ~x474 & ~x475 & ~x478 & ~x501 & ~x510 & ~x556 & ~x557 & ~x565 & ~x567 & ~x590 & ~x594 & ~x595 & ~x597 & ~x598 & ~x611 & ~x612 & ~x616 & ~x623 & ~x624 & ~x628 & ~x629 & ~x645 & ~x653 & ~x656 & ~x665 & ~x666 & ~x668 & ~x676 & ~x684 & ~x693 & ~x696 & ~x702 & ~x706 & ~x722 & ~x730 & ~x740 & ~x741 & ~x742 & ~x748 & ~x759 & ~x765 & ~x767 & ~x769 & ~x776;
assign c710 =  x240 &  x263 &  x264 &  x266 &  x435 &  x490 &  x601 &  x656 & ~x7 & ~x11 & ~x15 & ~x17 & ~x23 & ~x27 & ~x31 & ~x35 & ~x38 & ~x62 & ~x75 & ~x77 & ~x80 & ~x97 & ~x110 & ~x119 & ~x121 & ~x126 & ~x129 & ~x130 & ~x132 & ~x137 & ~x158 & ~x159 & ~x161 & ~x163 & ~x169 & ~x249 & ~x250 & ~x252 & ~x255 & ~x278 & ~x280 & ~x282 & ~x283 & ~x306 & ~x337 & ~x342 & ~x363 & ~x366 & ~x390 & ~x395 & ~x398 & ~x419 & ~x425 & ~x446 & ~x472 & ~x474 & ~x479 & ~x480 & ~x536 & ~x537 & ~x555 & ~x559 & ~x561 & ~x566 & ~x567 & ~x568 & ~x582 & ~x583 & ~x586 & ~x592 & ~x596 & ~x606 & ~x639 & ~x643 & ~x648 & ~x678 & ~x690 & ~x692 & ~x693 & ~x694 & ~x697 & ~x700 & ~x705 & ~x721 & ~x722 & ~x729 & ~x737 & ~x750 & ~x757 & ~x762 & ~x763 & ~x764 & ~x765 & ~x780;
assign c712 =  x561 &  x726;
assign c714 =  x236 &  x240 &  x241 &  x269 &  x325 &  x409 &  x437 & ~x6 & ~x9 & ~x10 & ~x15 & ~x26 & ~x31 & ~x38 & ~x42 & ~x46 & ~x49 & ~x54 & ~x55 & ~x56 & ~x59 & ~x61 & ~x63 & ~x66 & ~x70 & ~x71 & ~x74 & ~x86 & ~x94 & ~x105 & ~x114 & ~x135 & ~x139 & ~x141 & ~x144 & ~x145 & ~x155 & ~x156 & ~x162 & ~x163 & ~x165 & ~x195 & ~x251 & ~x275 & ~x277 & ~x281 & ~x282 & ~x330 & ~x331 & ~x333 & ~x337 & ~x396 & ~x397 & ~x446 & ~x451 & ~x476 & ~x477 & ~x507 & ~x508 & ~x513 & ~x530 & ~x531 & ~x532 & ~x533 & ~x535 & ~x556 & ~x581 & ~x582 & ~x586 & ~x589 & ~x590 & ~x591 & ~x595 & ~x611 & ~x614 & ~x616 & ~x635 & ~x644 & ~x650 & ~x663 & ~x671 & ~x698 & ~x700 & ~x723 & ~x724 & ~x733 & ~x735 & ~x751 & ~x760 & ~x764 & ~x767 & ~x772 & ~x775 & ~x776 & ~x782;
assign c716 =  x559;
assign c718 =  x300 & ~x54 & ~x59 & ~x133 & ~x163 & ~x284 & ~x376 & ~x402 & ~x427 & ~x509 & ~x510 & ~x603 & ~x604 & ~x646 & ~x732;
assign c720 =  x679;
assign c722 =  x266 &  x267 &  x440 & ~x0 & ~x2 & ~x3 & ~x4 & ~x6 & ~x7 & ~x11 & ~x12 & ~x13 & ~x15 & ~x16 & ~x17 & ~x20 & ~x24 & ~x27 & ~x28 & ~x33 & ~x35 & ~x36 & ~x37 & ~x43 & ~x44 & ~x46 & ~x48 & ~x50 & ~x51 & ~x53 & ~x54 & ~x55 & ~x57 & ~x59 & ~x63 & ~x65 & ~x74 & ~x76 & ~x79 & ~x80 & ~x85 & ~x86 & ~x87 & ~x88 & ~x89 & ~x92 & ~x96 & ~x100 & ~x107 & ~x110 & ~x116 & ~x119 & ~x121 & ~x122 & ~x124 & ~x125 & ~x126 & ~x127 & ~x128 & ~x130 & ~x132 & ~x134 & ~x137 & ~x139 & ~x142 & ~x144 & ~x156 & ~x158 & ~x159 & ~x161 & ~x165 & ~x166 & ~x167 & ~x168 & ~x170 & ~x186 & ~x188 & ~x190 & ~x191 & ~x194 & ~x219 & ~x221 & ~x222 & ~x225 & ~x226 & ~x251 & ~x277 & ~x279 & ~x281 & ~x304 & ~x305 & ~x308 & ~x310 & ~x332 & ~x334 & ~x336 & ~x337 & ~x362 & ~x367 & ~x368 & ~x387 & ~x388 & ~x389 & ~x390 & ~x393 & ~x423 & ~x446 & ~x447 & ~x448 & ~x473 & ~x477 & ~x479 & ~x501 & ~x502 & ~x506 & ~x529 & ~x531 & ~x532 & ~x535 & ~x554 & ~x555 & ~x556 & ~x560 & ~x569 & ~x570 & ~x582 & ~x583 & ~x584 & ~x585 & ~x587 & ~x595 & ~x610 & ~x611 & ~x612 & ~x613 & ~x614 & ~x617 & ~x618 & ~x620 & ~x622 & ~x623 & ~x626 & ~x639 & ~x643 & ~x644 & ~x648 & ~x651 & ~x652 & ~x653 & ~x654 & ~x665 & ~x667 & ~x675 & ~x678 & ~x693 & ~x695 & ~x698 & ~x700 & ~x702 & ~x703 & ~x705 & ~x706 & ~x709 & ~x720 & ~x721 & ~x728 & ~x735 & ~x737 & ~x749 & ~x751 & ~x752 & ~x756 & ~x760 & ~x761 & ~x770 & ~x771 & ~x772 & ~x774 & ~x775 & ~x776 & ~x778 & ~x779 & ~x782;
assign c724 =  x261 & ~x6 & ~x13 & ~x18 & ~x19 & ~x26 & ~x30 & ~x34 & ~x38 & ~x43 & ~x44 & ~x45 & ~x48 & ~x53 & ~x59 & ~x60 & ~x61 & ~x63 & ~x64 & ~x66 & ~x70 & ~x71 & ~x79 & ~x86 & ~x88 & ~x93 & ~x106 & ~x115 & ~x116 & ~x120 & ~x129 & ~x133 & ~x134 & ~x145 & ~x148 & ~x150 & ~x152 & ~x161 & ~x163 & ~x166 & ~x168 & ~x171 & ~x179 & ~x180 & ~x192 & ~x193 & ~x197 & ~x223 & ~x224 & ~x276 & ~x314 & ~x337 & ~x339 & ~x342 & ~x343 & ~x344 & ~x346 & ~x361 & ~x387 & ~x419 & ~x422 & ~x424 & ~x446 & ~x447 & ~x473 & ~x475 & ~x477 & ~x507 & ~x509 & ~x526 & ~x530 & ~x532 & ~x537 & ~x558 & ~x565 & ~x567 & ~x585 & ~x609 & ~x613 & ~x614 & ~x615 & ~x619 & ~x621 & ~x623 & ~x639 & ~x642 & ~x643 & ~x644 & ~x645 & ~x648 & ~x649 & ~x650 & ~x668 & ~x670 & ~x671 & ~x673 & ~x694 & ~x698 & ~x700 & ~x702 & ~x704 & ~x724 & ~x727 & ~x728 & ~x729 & ~x750 & ~x751 & ~x753 & ~x766 & ~x775 & ~x777 & ~x779;
assign c726 =  x268 &  x296 &  x410 & ~x0 & ~x4 & ~x5 & ~x7 & ~x14 & ~x15 & ~x16 & ~x22 & ~x23 & ~x24 & ~x29 & ~x33 & ~x34 & ~x36 & ~x44 & ~x48 & ~x52 & ~x55 & ~x60 & ~x68 & ~x79 & ~x85 & ~x101 & ~x104 & ~x111 & ~x115 & ~x120 & ~x121 & ~x127 & ~x131 & ~x155 & ~x157 & ~x161 & ~x162 & ~x166 & ~x169 & ~x190 & ~x194 & ~x225 & ~x248 & ~x278 & ~x333 & ~x335 & ~x370 & ~x373 & ~x394 & ~x416 & ~x417 & ~x420 & ~x421 & ~x450 & ~x473 & ~x480 & ~x501 & ~x504 & ~x541 & ~x554 & ~x556 & ~x559 & ~x560 & ~x561 & ~x564 & ~x589 & ~x609 & ~x611 & ~x620 & ~x621 & ~x622 & ~x624 & ~x648 & ~x652 & ~x667 & ~x671 & ~x672 & ~x695 & ~x696 & ~x700 & ~x708 & ~x720 & ~x723 & ~x727 & ~x730 & ~x735 & ~x736 & ~x737 & ~x748 & ~x753 & ~x757 & ~x775 & ~x783;
assign c728 =  x257 &  x262 & ~x122 & ~x181 & ~x554 & ~x558 & ~x622 & ~x644;
assign c730 =  x676;
assign c732 =  x209 &  x516 &  x599 & ~x104 & ~x168 & ~x250 & ~x313 & ~x317 & ~x318 & ~x331 & ~x391 & ~x445 & ~x475 & ~x594 & ~x603 & ~x609 & ~x614 & ~x647 & ~x659 & ~x662 & ~x663 & ~x687 & ~x688 & ~x691 & ~x714 & ~x719 & ~x728 & ~x741 & ~x766;
assign c734 =  x437 &  x463 & ~x3 & ~x7 & ~x8 & ~x9 & ~x10 & ~x11 & ~x13 & ~x18 & ~x19 & ~x20 & ~x21 & ~x26 & ~x32 & ~x33 & ~x37 & ~x39 & ~x40 & ~x41 & ~x43 & ~x47 & ~x48 & ~x49 & ~x50 & ~x52 & ~x55 & ~x56 & ~x59 & ~x61 & ~x64 & ~x65 & ~x68 & ~x71 & ~x75 & ~x78 & ~x82 & ~x83 & ~x86 & ~x89 & ~x90 & ~x91 & ~x92 & ~x94 & ~x95 & ~x97 & ~x99 & ~x101 & ~x104 & ~x105 & ~x109 & ~x110 & ~x111 & ~x118 & ~x119 & ~x120 & ~x122 & ~x130 & ~x132 & ~x133 & ~x136 & ~x138 & ~x139 & ~x141 & ~x161 & ~x162 & ~x163 & ~x164 & ~x166 & ~x168 & ~x171 & ~x172 & ~x189 & ~x190 & ~x191 & ~x192 & ~x193 & ~x221 & ~x224 & ~x225 & ~x250 & ~x253 & ~x254 & ~x255 & ~x275 & ~x276 & ~x278 & ~x279 & ~x281 & ~x282 & ~x303 & ~x305 & ~x307 & ~x310 & ~x331 & ~x334 & ~x336 & ~x340 & ~x345 & ~x348 & ~x349 & ~x360 & ~x361 & ~x362 & ~x364 & ~x365 & ~x367 & ~x369 & ~x370 & ~x372 & ~x374 & ~x376 & ~x377 & ~x387 & ~x388 & ~x390 & ~x393 & ~x422 & ~x423 & ~x446 & ~x448 & ~x451 & ~x474 & ~x477 & ~x479 & ~x480 & ~x501 & ~x502 & ~x503 & ~x505 & ~x508 & ~x528 & ~x533 & ~x534 & ~x535 & ~x537 & ~x556 & ~x558 & ~x560 & ~x564 & ~x566 & ~x567 & ~x569 & ~x590 & ~x593 & ~x594 & ~x597 & ~x607 & ~x609 & ~x613 & ~x614 & ~x619 & ~x620 & ~x623 & ~x624 & ~x635 & ~x638 & ~x643 & ~x644 & ~x645 & ~x647 & ~x649 & ~x650 & ~x664 & ~x667 & ~x668 & ~x669 & ~x671 & ~x672 & ~x677 & ~x678 & ~x695 & ~x699 & ~x700 & ~x706 & ~x707 & ~x717 & ~x718 & ~x721 & ~x722 & ~x725 & ~x727 & ~x731 & ~x733 & ~x745 & ~x748 & ~x751 & ~x756 & ~x758 & ~x759 & ~x762 & ~x764 & ~x767 & ~x768 & ~x774 & ~x775 & ~x778 & ~x781;
assign c736 =  x54;
assign c738 = ~x17 & ~x25 & ~x37 & ~x63 & ~x75 & ~x86 & ~x92 & ~x93 & ~x95 & ~x96 & ~x107 & ~x121 & ~x122 & ~x125 & ~x127 & ~x128 & ~x136 & ~x143 & ~x158 & ~x160 & ~x225 & ~x311 & ~x341 & ~x377 & ~x403 & ~x424 & ~x458 & ~x473 & ~x474 & ~x509 & ~x521 & ~x532 & ~x535 & ~x536 & ~x585 & ~x602 & ~x619 & ~x673 & ~x771 & ~x772 & ~x781;
assign c740 = ~x7 & ~x10 & ~x11 & ~x12 & ~x15 & ~x23 & ~x24 & ~x26 & ~x28 & ~x36 & ~x39 & ~x40 & ~x55 & ~x56 & ~x57 & ~x58 & ~x62 & ~x64 & ~x65 & ~x68 & ~x69 & ~x76 & ~x79 & ~x87 & ~x90 & ~x94 & ~x97 & ~x99 & ~x104 & ~x109 & ~x118 & ~x129 & ~x136 & ~x138 & ~x139 & ~x140 & ~x143 & ~x152 & ~x168 & ~x193 & ~x197 & ~x224 & ~x226 & ~x249 & ~x252 & ~x303 & ~x309 & ~x310 & ~x332 & ~x333 & ~x337 & ~x338 & ~x351 & ~x368 & ~x378 & ~x379 & ~x388 & ~x396 & ~x405 & ~x418 & ~x423 & ~x434 & ~x447 & ~x451 & ~x475 & ~x488 & ~x502 & ~x515 & ~x516 & ~x528 & ~x542 & ~x543 & ~x555 & ~x558 & ~x560 & ~x561 & ~x564 & ~x569 & ~x582 & ~x586 & ~x591 & ~x595 & ~x596 & ~x598 & ~x608 & ~x618 & ~x621 & ~x625 & ~x626 & ~x637 & ~x639 & ~x647 & ~x650 & ~x651 & ~x673 & ~x680 & ~x700 & ~x703 & ~x708 & ~x723 & ~x726 & ~x732 & ~x745 & ~x747 & ~x748 & ~x754 & ~x758 & ~x765 & ~x767 & ~x768 & ~x775 & ~x782;
assign c742 =  x367;
assign c744 =  x242 & ~x9 & ~x20 & ~x47 & ~x78 & ~x80 & ~x121 & ~x161 & ~x313 & ~x336 & ~x350 & ~x376 & ~x391 & ~x403 & ~x404 & ~x410 & ~x426 & ~x429 & ~x440 & ~x446 & ~x502 & ~x532 & ~x578 & ~x585 & ~x635 & ~x688 & ~x717 & ~x722 & ~x770;
assign c746 =  x282;
assign c748 =  x321 &  x322 & ~x5 & ~x15 & ~x26 & ~x29 & ~x57 & ~x61 & ~x68 & ~x94 & ~x107 & ~x114 & ~x115 & ~x130 & ~x133 & ~x134 & ~x140 & ~x152 & ~x153 & ~x154 & ~x156 & ~x160 & ~x162 & ~x170 & ~x172 & ~x173 & ~x174 & ~x176 & ~x177 & ~x178 & ~x181 & ~x194 & ~x195 & ~x197 & ~x207 & ~x209 & ~x210 & ~x211 & ~x219 & ~x221 & ~x222 & ~x236 & ~x238 & ~x249 & ~x278 & ~x306 & ~x361 & ~x363 & ~x390 & ~x417 & ~x420 & ~x444 & ~x446 & ~x447 & ~x448 & ~x476 & ~x477 & ~x499 & ~x500 & ~x513 & ~x567 & ~x585 & ~x586 & ~x594 & ~x595 & ~x611 & ~x617 & ~x620 & ~x638 & ~x667 & ~x669 & ~x673 & ~x675 & ~x704 & ~x753 & ~x757 & ~x760 & ~x761 & ~x764 & ~x765 & ~x767 & ~x768;
assign c752 =  x227;
assign c754 = ~x6 & ~x11 & ~x14 & ~x19 & ~x27 & ~x30 & ~x31 & ~x32 & ~x37 & ~x38 & ~x50 & ~x51 & ~x52 & ~x57 & ~x58 & ~x62 & ~x66 & ~x69 & ~x89 & ~x94 & ~x99 & ~x103 & ~x113 & ~x114 & ~x118 & ~x120 & ~x127 & ~x131 & ~x135 & ~x146 & ~x149 & ~x150 & ~x158 & ~x161 & ~x165 & ~x169 & ~x173 & ~x175 & ~x197 & ~x205 & ~x219 & ~x227 & ~x250 & ~x252 & ~x283 & ~x304 & ~x305 & ~x333 & ~x337 & ~x361 & ~x362 & ~x363 & ~x391 & ~x394 & ~x401 & ~x403 & ~x417 & ~x423 & ~x429 & ~x431 & ~x449 & ~x474 & ~x478 & ~x485 & ~x505 & ~x512 & ~x527 & ~x531 & ~x533 & ~x535 & ~x541 & ~x556 & ~x561 & ~x563 & ~x567 & ~x568 & ~x585 & ~x589 & ~x595 & ~x596 & ~x613 & ~x614 & ~x619 & ~x621 & ~x622 & ~x637 & ~x638 & ~x642 & ~x643 & ~x645 & ~x656 & ~x665 & ~x669 & ~x698 & ~x701 & ~x733 & ~x739 & ~x742 & ~x743 & ~x751 & ~x753 & ~x754 & ~x756 & ~x763 & ~x767 & ~x771 & ~x773 & ~x774 & ~x776 & ~x779;
assign c756 = ~x1 & ~x7 & ~x8 & ~x23 & ~x26 & ~x27 & ~x30 & ~x31 & ~x32 & ~x41 & ~x42 & ~x46 & ~x51 & ~x54 & ~x55 & ~x58 & ~x70 & ~x71 & ~x72 & ~x73 & ~x77 & ~x83 & ~x89 & ~x90 & ~x91 & ~x94 & ~x98 & ~x99 & ~x104 & ~x108 & ~x109 & ~x125 & ~x126 & ~x133 & ~x136 & ~x139 & ~x141 & ~x145 & ~x147 & ~x150 & ~x154 & ~x157 & ~x159 & ~x160 & ~x161 & ~x163 & ~x169 & ~x177 & ~x178 & ~x191 & ~x193 & ~x194 & ~x199 & ~x222 & ~x223 & ~x224 & ~x225 & ~x249 & ~x251 & ~x253 & ~x254 & ~x279 & ~x312 & ~x335 & ~x337 & ~x363 & ~x364 & ~x366 & ~x378 & ~x379 & ~x389 & ~x406 & ~x420 & ~x434 & ~x445 & ~x449 & ~x461 & ~x472 & ~x474 & ~x486 & ~x498 & ~x500 & ~x502 & ~x503 & ~x505 & ~x515 & ~x528 & ~x529 & ~x539 & ~x541 & ~x555 & ~x557 & ~x558 & ~x567 & ~x568 & ~x569 & ~x570 & ~x584 & ~x588 & ~x590 & ~x593 & ~x595 & ~x607 & ~x611 & ~x613 & ~x614 & ~x616 & ~x623 & ~x638 & ~x642 & ~x644 & ~x649 & ~x650 & ~x664 & ~x666 & ~x679 & ~x694 & ~x696 & ~x700 & ~x701 & ~x725 & ~x727 & ~x732 & ~x733 & ~x734 & ~x744 & ~x747 & ~x748 & ~x758 & ~x760 & ~x765 & ~x766 & ~x768 & ~x769 & ~x771 & ~x773 & ~x775 & ~x777 & ~x783;
assign c758 =  x436 &  x437 & ~x0 & ~x1 & ~x4 & ~x5 & ~x6 & ~x8 & ~x11 & ~x12 & ~x14 & ~x15 & ~x17 & ~x18 & ~x20 & ~x21 & ~x23 & ~x25 & ~x28 & ~x29 & ~x31 & ~x34 & ~x35 & ~x37 & ~x39 & ~x41 & ~x42 & ~x45 & ~x46 & ~x49 & ~x51 & ~x52 & ~x53 & ~x56 & ~x58 & ~x59 & ~x62 & ~x65 & ~x67 & ~x69 & ~x70 & ~x72 & ~x74 & ~x76 & ~x78 & ~x82 & ~x85 & ~x92 & ~x94 & ~x96 & ~x97 & ~x98 & ~x109 & ~x110 & ~x116 & ~x118 & ~x120 & ~x122 & ~x123 & ~x124 & ~x125 & ~x126 & ~x128 & ~x129 & ~x130 & ~x135 & ~x136 & ~x138 & ~x141 & ~x144 & ~x157 & ~x158 & ~x160 & ~x163 & ~x164 & ~x165 & ~x169 & ~x170 & ~x171 & ~x192 & ~x193 & ~x195 & ~x197 & ~x198 & ~x199 & ~x221 & ~x226 & ~x227 & ~x251 & ~x254 & ~x277 & ~x280 & ~x281 & ~x283 & ~x306 & ~x307 & ~x309 & ~x310 & ~x313 & ~x314 & ~x316 & ~x317 & ~x318 & ~x319 & ~x321 & ~x331 & ~x332 & ~x333 & ~x334 & ~x336 & ~x337 & ~x342 & ~x359 & ~x361 & ~x363 & ~x366 & ~x367 & ~x368 & ~x369 & ~x371 & ~x390 & ~x391 & ~x392 & ~x418 & ~x419 & ~x425 & ~x426 & ~x445 & ~x446 & ~x447 & ~x451 & ~x452 & ~x472 & ~x479 & ~x480 & ~x497 & ~x500 & ~x501 & ~x503 & ~x506 & ~x507 & ~x508 & ~x524 & ~x526 & ~x528 & ~x534 & ~x535 & ~x536 & ~x537 & ~x555 & ~x556 & ~x558 & ~x559 & ~x562 & ~x563 & ~x578 & ~x581 & ~x592 & ~x594 & ~x609 & ~x610 & ~x611 & ~x612 & ~x613 & ~x615 & ~x616 & ~x617 & ~x619 & ~x620 & ~x635 & ~x639 & ~x640 & ~x641 & ~x643 & ~x645 & ~x649 & ~x663 & ~x664 & ~x665 & ~x667 & ~x668 & ~x670 & ~x671 & ~x673 & ~x674 & ~x698 & ~x700 & ~x705 & ~x720 & ~x721 & ~x728 & ~x733 & ~x735 & ~x737 & ~x744 & ~x745 & ~x746 & ~x747 & ~x748 & ~x749 & ~x751 & ~x752 & ~x758 & ~x760 & ~x761 & ~x764 & ~x769 & ~x773 & ~x774 & ~x775 & ~x776 & ~x779 & ~x781 & ~x783;
assign c760 =  x736;
assign c762 =  x233 &  x234 &  x236 &  x237 &  x262 &  x263 &  x264 &  x266 &  x267 &  x464 &  x519 & ~x0 & ~x3 & ~x22 & ~x25 & ~x34 & ~x39 & ~x41 & ~x55 & ~x62 & ~x66 & ~x71 & ~x77 & ~x81 & ~x106 & ~x115 & ~x126 & ~x139 & ~x142 & ~x144 & ~x146 & ~x151 & ~x152 & ~x154 & ~x155 & ~x156 & ~x157 & ~x169 & ~x182 & ~x221 & ~x223 & ~x277 & ~x331 & ~x333 & ~x335 & ~x340 & ~x367 & ~x449 & ~x473 & ~x501 & ~x504 & ~x508 & ~x530 & ~x532 & ~x585 & ~x596 & ~x607 & ~x608 & ~x610 & ~x617 & ~x618 & ~x620 & ~x622 & ~x639 & ~x644 & ~x650 & ~x671 & ~x679 & ~x680 & ~x691 & ~x697 & ~x701 & ~x722 & ~x728 & ~x732 & ~x734 & ~x746 & ~x752 & ~x756 & ~x774;
assign c764 =  x267 &  x410 &  x544 &  x653;
assign c766 =  x271 & ~x8 & ~x31 & ~x39 & ~x47 & ~x64 & ~x72 & ~x79 & ~x82 & ~x85 & ~x90 & ~x101 & ~x102 & ~x107 & ~x111 & ~x114 & ~x126 & ~x130 & ~x141 & ~x142 & ~x147 & ~x155 & ~x156 & ~x157 & ~x161 & ~x167 & ~x197 & ~x199 & ~x200 & ~x221 & ~x306 & ~x361 & ~x362 & ~x378 & ~x388 & ~x389 & ~x404 & ~x415 & ~x416 & ~x421 & ~x422 & ~x432 & ~x451 & ~x458 & ~x482 & ~x486 & ~x501 & ~x508 & ~x531 & ~x582 & ~x585 & ~x589 & ~x610 & ~x614 & ~x619 & ~x638 & ~x642 & ~x643 & ~x673 & ~x674 & ~x695 & ~x725 & ~x729 & ~x740 & ~x745 & ~x754 & ~x780 & ~x781;
assign c768 =  x227;
assign c770 =  x15;
assign c772 =  x243 &  x269 &  x270 &  x271 &  x490 &  x572 & ~x13 & ~x47 & ~x77 & ~x113 & ~x122 & ~x127 & ~x133 & ~x198 & ~x199 & ~x378 & ~x539 & ~x553 & ~x621 & ~x635 & ~x721 & ~x746 & ~x760;
assign c774 =  x268 &  x433 &  x438 &  x440 & ~x569 & ~x598;
assign c776 =  x260 &  x268 &  x289 &  x290 &  x292 &  x463 &  x491 &  x519 & ~x48 & ~x55 & ~x71 & ~x104 & ~x111 & ~x113 & ~x121 & ~x123 & ~x145 & ~x151 & ~x152 & ~x164 & ~x248 & ~x250 & ~x304 & ~x311 & ~x359 & ~x419 & ~x420 & ~x536 & ~x564 & ~x622 & ~x704 & ~x777;
assign c778 =  x293 &  x294 & ~x0 & ~x9 & ~x16 & ~x28 & ~x38 & ~x42 & ~x44 & ~x45 & ~x48 & ~x61 & ~x68 & ~x71 & ~x83 & ~x84 & ~x123 & ~x125 & ~x126 & ~x129 & ~x138 & ~x141 & ~x144 & ~x154 & ~x156 & ~x157 & ~x164 & ~x174 & ~x183 & ~x185 & ~x194 & ~x208 & ~x209 & ~x211 & ~x212 & ~x220 & ~x224 & ~x392 & ~x403 & ~x419 & ~x421 & ~x424 & ~x472 & ~x474 & ~x476 & ~x502 & ~x527 & ~x529 & ~x532 & ~x538 & ~x565 & ~x582 & ~x593 & ~x619 & ~x643 & ~x701 & ~x723 & ~x729 & ~x773 & ~x779 & ~x782;
assign c780 = ~x0 & ~x2 & ~x4 & ~x6 & ~x9 & ~x11 & ~x12 & ~x13 & ~x16 & ~x21 & ~x22 & ~x23 & ~x30 & ~x35 & ~x38 & ~x39 & ~x41 & ~x42 & ~x43 & ~x46 & ~x47 & ~x48 & ~x50 & ~x53 & ~x56 & ~x57 & ~x58 & ~x60 & ~x64 & ~x65 & ~x73 & ~x78 & ~x79 & ~x81 & ~x82 & ~x86 & ~x89 & ~x93 & ~x94 & ~x97 & ~x101 & ~x104 & ~x106 & ~x107 & ~x108 & ~x109 & ~x118 & ~x121 & ~x122 & ~x123 & ~x124 & ~x129 & ~x133 & ~x138 & ~x141 & ~x149 & ~x150 & ~x151 & ~x156 & ~x157 & ~x158 & ~x159 & ~x160 & ~x162 & ~x165 & ~x166 & ~x170 & ~x174 & ~x180 & ~x190 & ~x194 & ~x198 & ~x200 & ~x220 & ~x247 & ~x304 & ~x305 & ~x307 & ~x308 & ~x335 & ~x336 & ~x337 & ~x338 & ~x363 & ~x364 & ~x365 & ~x378 & ~x390 & ~x391 & ~x406 & ~x416 & ~x417 & ~x419 & ~x421 & ~x432 & ~x433 & ~x434 & ~x444 & ~x446 & ~x448 & ~x449 & ~x458 & ~x473 & ~x476 & ~x485 & ~x501 & ~x505 & ~x506 & ~x513 & ~x514 & ~x527 & ~x528 & ~x532 & ~x533 & ~x534 & ~x535 & ~x542 & ~x557 & ~x562 & ~x563 & ~x569 & ~x570 & ~x582 & ~x585 & ~x586 & ~x587 & ~x588 & ~x595 & ~x597 & ~x598 & ~x611 & ~x612 & ~x613 & ~x619 & ~x624 & ~x625 & ~x638 & ~x639 & ~x640 & ~x643 & ~x667 & ~x669 & ~x670 & ~x671 & ~x673 & ~x674 & ~x694 & ~x695 & ~x697 & ~x698 & ~x702 & ~x704 & ~x705 & ~x722 & ~x723 & ~x724 & ~x725 & ~x730 & ~x731 & ~x733 & ~x734 & ~x738 & ~x751 & ~x756 & ~x760 & ~x778 & ~x780 & ~x781 & ~x783;
assign c782 =  x265 & ~x15 & ~x21 & ~x23 & ~x38 & ~x41 & ~x46 & ~x50 & ~x53 & ~x63 & ~x81 & ~x86 & ~x137 & ~x141 & ~x147 & ~x154 & ~x223 & ~x225 & ~x279 & ~x309 & ~x333 & ~x359 & ~x365 & ~x376 & ~x377 & ~x391 & ~x393 & ~x415 & ~x430 & ~x431 & ~x444 & ~x456 & ~x496 & ~x510 & ~x524 & ~x555 & ~x579 & ~x608 & ~x609 & ~x614 & ~x618 & ~x665 & ~x695 & ~x738 & ~x744 & ~x760 & ~x781;
assign c784 =  x316 &  x317 &  x318 &  x319 & ~x53 & ~x183 & ~x210 & ~x431 & ~x558 & ~x582;
assign c786 =  x229 &  x230;
assign c788 =  x436 &  x464 & ~x0 & ~x2 & ~x4 & ~x6 & ~x7 & ~x8 & ~x9 & ~x12 & ~x13 & ~x15 & ~x24 & ~x27 & ~x30 & ~x34 & ~x39 & ~x41 & ~x42 & ~x44 & ~x45 & ~x50 & ~x54 & ~x55 & ~x56 & ~x57 & ~x60 & ~x61 & ~x67 & ~x69 & ~x70 & ~x71 & ~x73 & ~x77 & ~x78 & ~x81 & ~x89 & ~x92 & ~x96 & ~x98 & ~x99 & ~x106 & ~x111 & ~x112 & ~x117 & ~x120 & ~x121 & ~x122 & ~x127 & ~x128 & ~x129 & ~x130 & ~x131 & ~x132 & ~x135 & ~x138 & ~x141 & ~x161 & ~x163 & ~x166 & ~x168 & ~x169 & ~x171 & ~x172 & ~x191 & ~x196 & ~x199 & ~x219 & ~x220 & ~x221 & ~x225 & ~x226 & ~x246 & ~x247 & ~x249 & ~x250 & ~x251 & ~x253 & ~x274 & ~x275 & ~x276 & ~x277 & ~x279 & ~x301 & ~x302 & ~x307 & ~x311 & ~x328 & ~x329 & ~x330 & ~x331 & ~x332 & ~x335 & ~x337 & ~x338 & ~x339 & ~x348 & ~x355 & ~x358 & ~x360 & ~x364 & ~x368 & ~x373 & ~x374 & ~x375 & ~x377 & ~x383 & ~x389 & ~x391 & ~x393 & ~x394 & ~x395 & ~x396 & ~x397 & ~x418 & ~x422 & ~x425 & ~x450 & ~x473 & ~x474 & ~x476 & ~x500 & ~x501 & ~x502 & ~x503 & ~x504 & ~x509 & ~x527 & ~x530 & ~x531 & ~x534 & ~x536 & ~x538 & ~x540 & ~x557 & ~x560 & ~x563 & ~x564 & ~x566 & ~x567 & ~x568 & ~x569 & ~x570 & ~x571 & ~x582 & ~x584 & ~x588 & ~x589 & ~x594 & ~x595 & ~x608 & ~x609 & ~x612 & ~x614 & ~x615 & ~x616 & ~x622 & ~x623 & ~x624 & ~x626 & ~x627 & ~x636 & ~x637 & ~x639 & ~x641 & ~x644 & ~x646 & ~x647 & ~x649 & ~x650 & ~x666 & ~x667 & ~x668 & ~x669 & ~x670 & ~x671 & ~x672 & ~x673 & ~x674 & ~x677 & ~x679 & ~x680 & ~x681 & ~x693 & ~x695 & ~x696 & ~x707 & ~x708 & ~x709 & ~x722 & ~x724 & ~x728 & ~x729 & ~x731 & ~x732 & ~x733 & ~x738 & ~x747 & ~x748 & ~x759 & ~x763 & ~x764 & ~x767 & ~x770 & ~x776 & ~x779 & ~x783;
assign c790 = ~x0 & ~x7 & ~x10 & ~x13 & ~x15 & ~x21 & ~x24 & ~x29 & ~x34 & ~x35 & ~x37 & ~x38 & ~x39 & ~x51 & ~x52 & ~x53 & ~x55 & ~x56 & ~x69 & ~x72 & ~x73 & ~x75 & ~x76 & ~x79 & ~x82 & ~x83 & ~x87 & ~x94 & ~x95 & ~x97 & ~x98 & ~x99 & ~x100 & ~x102 & ~x104 & ~x108 & ~x109 & ~x110 & ~x111 & ~x113 & ~x116 & ~x117 & ~x124 & ~x126 & ~x128 & ~x131 & ~x133 & ~x136 & ~x143 & ~x144 & ~x149 & ~x151 & ~x154 & ~x155 & ~x161 & ~x163 & ~x167 & ~x169 & ~x174 & ~x177 & ~x179 & ~x180 & ~x183 & ~x186 & ~x187 & ~x188 & ~x193 & ~x212 & ~x222 & ~x223 & ~x250 & ~x251 & ~x280 & ~x306 & ~x307 & ~x309 & ~x363 & ~x365 & ~x391 & ~x393 & ~x407 & ~x417 & ~x420 & ~x433 & ~x434 & ~x444 & ~x445 & ~x450 & ~x460 & ~x461 & ~x462 & ~x473 & ~x474 & ~x476 & ~x488 & ~x490 & ~x499 & ~x500 & ~x501 & ~x502 & ~x516 & ~x517 & ~x518 & ~x532 & ~x535 & ~x545 & ~x557 & ~x558 & ~x562 & ~x567 & ~x568 & ~x571 & ~x572 & ~x583 & ~x584 & ~x590 & ~x595 & ~x597 & ~x598 & ~x599 & ~x600 & ~x619 & ~x620 & ~x623 & ~x626 & ~x639 & ~x641 & ~x642 & ~x647 & ~x649 & ~x653 & ~x670 & ~x677 & ~x694 & ~x695 & ~x698 & ~x703 & ~x704 & ~x705 & ~x708 & ~x710 & ~x724 & ~x725 & ~x726 & ~x727 & ~x728 & ~x729 & ~x731 & ~x737 & ~x754 & ~x755 & ~x759 & ~x762 & ~x766 & ~x767 & ~x775;
assign c792 = ~x3 & ~x5 & ~x34 & ~x39 & ~x54 & ~x59 & ~x71 & ~x72 & ~x79 & ~x117 & ~x122 & ~x127 & ~x147 & ~x201 & ~x220 & ~x255 & ~x257 & ~x307 & ~x308 & ~x322 & ~x350 & ~x378 & ~x405 & ~x422 & ~x432 & ~x443 & ~x448 & ~x467 & ~x481 & ~x498 & ~x500 & ~x511 & ~x531 & ~x539 & ~x583 & ~x610 & ~x614 & ~x689 & ~x691 & ~x749 & ~x752 & ~x764 & ~x770;
assign c794 =  x237 & ~x4 & ~x10 & ~x13 & ~x14 & ~x17 & ~x20 & ~x21 & ~x25 & ~x30 & ~x33 & ~x35 & ~x39 & ~x42 & ~x43 & ~x49 & ~x54 & ~x65 & ~x67 & ~x70 & ~x73 & ~x74 & ~x79 & ~x82 & ~x87 & ~x90 & ~x94 & ~x97 & ~x105 & ~x108 & ~x109 & ~x123 & ~x125 & ~x126 & ~x129 & ~x132 & ~x133 & ~x138 & ~x139 & ~x140 & ~x141 & ~x149 & ~x152 & ~x153 & ~x155 & ~x158 & ~x161 & ~x162 & ~x166 & ~x170 & ~x172 & ~x173 & ~x174 & ~x195 & ~x223 & ~x253 & ~x282 & ~x286 & ~x302 & ~x303 & ~x304 & ~x307 & ~x309 & ~x312 & ~x313 & ~x315 & ~x317 & ~x319 & ~x320 & ~x330 & ~x338 & ~x340 & ~x347 & ~x363 & ~x368 & ~x369 & ~x372 & ~x386 & ~x387 & ~x389 & ~x390 & ~x396 & ~x397 & ~x415 & ~x417 & ~x420 & ~x423 & ~x445 & ~x452 & ~x453 & ~x476 & ~x481 & ~x498 & ~x501 & ~x502 & ~x503 & ~x504 & ~x507 & ~x525 & ~x529 & ~x534 & ~x538 & ~x555 & ~x560 & ~x561 & ~x581 & ~x582 & ~x586 & ~x588 & ~x591 & ~x593 & ~x609 & ~x610 & ~x613 & ~x615 & ~x619 & ~x649 & ~x663 & ~x664 & ~x669 & ~x671 & ~x673 & ~x674 & ~x678 & ~x690 & ~x691 & ~x698 & ~x703 & ~x720 & ~x724 & ~x734 & ~x735 & ~x738 & ~x740 & ~x746 & ~x747 & ~x749 & ~x758 & ~x759 & ~x773 & ~x780 & ~x782;
assign c796 = ~x18 & ~x19 & ~x31 & ~x40 & ~x46 & ~x50 & ~x73 & ~x84 & ~x88 & ~x100 & ~x102 & ~x104 & ~x105 & ~x108 & ~x129 & ~x132 & ~x135 & ~x150 & ~x155 & ~x159 & ~x161 & ~x166 & ~x168 & ~x177 & ~x178 & ~x184 & ~x185 & ~x219 & ~x221 & ~x222 & ~x226 & ~x254 & ~x337 & ~x418 & ~x432 & ~x448 & ~x478 & ~x487 & ~x492 & ~x532 & ~x538 & ~x542 & ~x565 & ~x566 & ~x602 & ~x612 & ~x638 & ~x645 & ~x651 & ~x667 & ~x672 & ~x702 & ~x737 & ~x751 & ~x753 & ~x767 & ~x769 & ~x771 & ~x783;
assign c798 = ~x1 & ~x4 & ~x6 & ~x9 & ~x10 & ~x15 & ~x17 & ~x20 & ~x21 & ~x24 & ~x27 & ~x28 & ~x29 & ~x31 & ~x34 & ~x36 & ~x38 & ~x39 & ~x42 & ~x44 & ~x45 & ~x49 & ~x50 & ~x51 & ~x54 & ~x58 & ~x64 & ~x65 & ~x66 & ~x70 & ~x73 & ~x79 & ~x81 & ~x83 & ~x86 & ~x88 & ~x91 & ~x93 & ~x94 & ~x96 & ~x103 & ~x105 & ~x106 & ~x107 & ~x108 & ~x111 & ~x112 & ~x113 & ~x117 & ~x118 & ~x119 & ~x122 & ~x125 & ~x126 & ~x128 & ~x137 & ~x138 & ~x139 & ~x140 & ~x141 & ~x142 & ~x145 & ~x148 & ~x149 & ~x151 & ~x153 & ~x154 & ~x155 & ~x158 & ~x161 & ~x164 & ~x166 & ~x167 & ~x168 & ~x174 & ~x178 & ~x184 & ~x185 & ~x190 & ~x191 & ~x192 & ~x193 & ~x197 & ~x222 & ~x223 & ~x224 & ~x225 & ~x252 & ~x277 & ~x279 & ~x282 & ~x306 & ~x333 & ~x334 & ~x335 & ~x336 & ~x337 & ~x364 & ~x389 & ~x391 & ~x393 & ~x415 & ~x416 & ~x420 & ~x432 & ~x433 & ~x434 & ~x443 & ~x448 & ~x449 & ~x450 & ~x460 & ~x461 & ~x472 & ~x473 & ~x474 & ~x475 & ~x477 & ~x479 & ~x487 & ~x488 & ~x499 & ~x500 & ~x503 & ~x505 & ~x506 & ~x514 & ~x515 & ~x516 & ~x517 & ~x527 & ~x529 & ~x531 & ~x532 & ~x542 & ~x543 & ~x544 & ~x555 & ~x564 & ~x565 & ~x566 & ~x567 & ~x570 & ~x571 & ~x583 & ~x584 & ~x589 & ~x591 & ~x592 & ~x593 & ~x594 & ~x595 & ~x596 & ~x598 & ~x611 & ~x620 & ~x623 & ~x624 & ~x625 & ~x641 & ~x647 & ~x649 & ~x650 & ~x651 & ~x652 & ~x668 & ~x672 & ~x677 & ~x678 & ~x679 & ~x696 & ~x698 & ~x700 & ~x704 & ~x705 & ~x711 & ~x724 & ~x727 & ~x731 & ~x739 & ~x741 & ~x746 & ~x752 & ~x753 & ~x754 & ~x755 & ~x758 & ~x759 & ~x761 & ~x763 & ~x764 & ~x766 & ~x770 & ~x773 & ~x775 & ~x780;
assign c7100 = ~x6 & ~x8 & ~x10 & ~x12 & ~x27 & ~x30 & ~x33 & ~x35 & ~x43 & ~x45 & ~x49 & ~x58 & ~x60 & ~x61 & ~x69 & ~x84 & ~x94 & ~x97 & ~x98 & ~x100 & ~x101 & ~x106 & ~x107 & ~x110 & ~x111 & ~x113 & ~x114 & ~x119 & ~x121 & ~x126 & ~x136 & ~x141 & ~x144 & ~x145 & ~x151 & ~x152 & ~x154 & ~x155 & ~x158 & ~x159 & ~x161 & ~x167 & ~x192 & ~x194 & ~x198 & ~x222 & ~x226 & ~x252 & ~x254 & ~x275 & ~x281 & ~x284 & ~x290 & ~x305 & ~x309 & ~x310 & ~x315 & ~x319 & ~x321 & ~x329 & ~x334 & ~x335 & ~x339 & ~x340 & ~x343 & ~x349 & ~x360 & ~x362 & ~x363 & ~x364 & ~x370 & ~x373 & ~x386 & ~x387 & ~x390 & ~x395 & ~x400 & ~x415 & ~x420 & ~x421 & ~x448 & ~x451 & ~x503 & ~x504 & ~x507 & ~x508 & ~x527 & ~x528 & ~x533 & ~x551 & ~x558 & ~x560 & ~x582 & ~x583 & ~x584 & ~x585 & ~x588 & ~x595 & ~x597 & ~x606 & ~x607 & ~x608 & ~x610 & ~x611 & ~x612 & ~x614 & ~x615 & ~x618 & ~x622 & ~x623 & ~x634 & ~x636 & ~x638 & ~x639 & ~x645 & ~x652 & ~x662 & ~x668 & ~x675 & ~x676 & ~x677 & ~x678 & ~x679 & ~x691 & ~x693 & ~x695 & ~x699 & ~x710 & ~x718 & ~x721 & ~x722 & ~x733 & ~x735 & ~x752 & ~x754 & ~x757 & ~x758 & ~x762 & ~x775 & ~x776 & ~x779 & ~x780;
assign c7102 = ~x10 & ~x12 & ~x22 & ~x29 & ~x43 & ~x60 & ~x69 & ~x71 & ~x75 & ~x80 & ~x82 & ~x85 & ~x92 & ~x93 & ~x104 & ~x109 & ~x119 & ~x122 & ~x127 & ~x130 & ~x141 & ~x150 & ~x166 & ~x169 & ~x189 & ~x211 & ~x221 & ~x225 & ~x307 & ~x360 & ~x363 & ~x403 & ~x405 & ~x424 & ~x428 & ~x430 & ~x455 & ~x457 & ~x483 & ~x505 & ~x509 & ~x526 & ~x529 & ~x555 & ~x556 & ~x561 & ~x581 & ~x588 & ~x613 & ~x615 & ~x643 & ~x645 & ~x672 & ~x693 & ~x697 & ~x726 & ~x751 & ~x754 & ~x771 & ~x780;
assign c7104 =  x355 & ~x0 & ~x10 & ~x12 & ~x15 & ~x17 & ~x22 & ~x23 & ~x25 & ~x32 & ~x33 & ~x36 & ~x41 & ~x45 & ~x50 & ~x55 & ~x61 & ~x64 & ~x65 & ~x67 & ~x68 & ~x69 & ~x70 & ~x72 & ~x82 & ~x85 & ~x86 & ~x87 & ~x88 & ~x89 & ~x91 & ~x93 & ~x94 & ~x95 & ~x99 & ~x100 & ~x102 & ~x104 & ~x106 & ~x114 & ~x115 & ~x119 & ~x120 & ~x121 & ~x124 & ~x125 & ~x133 & ~x143 & ~x147 & ~x148 & ~x149 & ~x160 & ~x163 & ~x164 & ~x167 & ~x171 & ~x173 & ~x175 & ~x190 & ~x191 & ~x192 & ~x199 & ~x200 & ~x203 & ~x204 & ~x205 & ~x220 & ~x223 & ~x226 & ~x249 & ~x251 & ~x253 & ~x254 & ~x278 & ~x280 & ~x304 & ~x306 & ~x307 & ~x308 & ~x311 & ~x332 & ~x333 & ~x337 & ~x360 & ~x364 & ~x365 & ~x388 & ~x389 & ~x392 & ~x405 & ~x417 & ~x422 & ~x432 & ~x433 & ~x445 & ~x447 & ~x460 & ~x473 & ~x474 & ~x477 & ~x487 & ~x488 & ~x499 & ~x501 & ~x505 & ~x514 & ~x515 & ~x529 & ~x531 & ~x532 & ~x534 & ~x536 & ~x562 & ~x563 & ~x565 & ~x569 & ~x583 & ~x584 & ~x585 & ~x586 & ~x590 & ~x593 & ~x594 & ~x597 & ~x613 & ~x614 & ~x616 & ~x619 & ~x624 & ~x643 & ~x644 & ~x645 & ~x646 & ~x670 & ~x673 & ~x674 & ~x691 & ~x699 & ~x701 & ~x703 & ~x707 & ~x723 & ~x726 & ~x748 & ~x754 & ~x756 & ~x759 & ~x760 & ~x763 & ~x765 & ~x767 & ~x771 & ~x773 & ~x776 & ~x780 & ~x782;
assign c7106 =  x292 &  x293 & ~x0 & ~x3 & ~x4 & ~x10 & ~x15 & ~x20 & ~x22 & ~x29 & ~x31 & ~x33 & ~x35 & ~x44 & ~x45 & ~x46 & ~x47 & ~x49 & ~x56 & ~x60 & ~x61 & ~x66 & ~x67 & ~x68 & ~x69 & ~x75 & ~x82 & ~x84 & ~x88 & ~x91 & ~x92 & ~x93 & ~x95 & ~x96 & ~x104 & ~x107 & ~x111 & ~x114 & ~x117 & ~x118 & ~x119 & ~x120 & ~x124 & ~x128 & ~x130 & ~x133 & ~x135 & ~x136 & ~x140 & ~x149 & ~x152 & ~x153 & ~x154 & ~x155 & ~x159 & ~x160 & ~x170 & ~x181 & ~x194 & ~x199 & ~x219 & ~x224 & ~x226 & ~x247 & ~x252 & ~x282 & ~x304 & ~x309 & ~x330 & ~x332 & ~x335 & ~x337 & ~x339 & ~x364 & ~x365 & ~x397 & ~x400 & ~x447 & ~x448 & ~x450 & ~x475 & ~x476 & ~x502 & ~x504 & ~x509 & ~x527 & ~x528 & ~x531 & ~x537 & ~x538 & ~x543 & ~x552 & ~x553 & ~x555 & ~x556 & ~x557 & ~x568 & ~x569 & ~x571 & ~x581 & ~x583 & ~x586 & ~x591 & ~x592 & ~x594 & ~x598 & ~x608 & ~x611 & ~x612 & ~x613 & ~x615 & ~x625 & ~x627 & ~x637 & ~x641 & ~x642 & ~x650 & ~x651 & ~x652 & ~x653 & ~x654 & ~x655 & ~x666 & ~x671 & ~x672 & ~x677 & ~x681 & ~x697 & ~x701 & ~x702 & ~x705 & ~x706 & ~x707 & ~x708 & ~x722 & ~x723 & ~x726 & ~x731 & ~x732 & ~x734 & ~x745 & ~x754 & ~x755 & ~x756 & ~x759 & ~x776 & ~x777 & ~x778 & ~x779 & ~x783;
assign c7108 =  x778;
assign c7110 =  x290 & ~x5 & ~x6 & ~x9 & ~x16 & ~x22 & ~x28 & ~x32 & ~x33 & ~x51 & ~x52 & ~x56 & ~x64 & ~x66 & ~x67 & ~x68 & ~x71 & ~x73 & ~x74 & ~x75 & ~x76 & ~x80 & ~x82 & ~x83 & ~x84 & ~x93 & ~x95 & ~x108 & ~x116 & ~x118 & ~x125 & ~x135 & ~x138 & ~x139 & ~x140 & ~x143 & ~x144 & ~x147 & ~x150 & ~x153 & ~x154 & ~x160 & ~x161 & ~x162 & ~x181 & ~x182 & ~x183 & ~x191 & ~x193 & ~x195 & ~x196 & ~x225 & ~x252 & ~x277 & ~x278 & ~x305 & ~x307 & ~x309 & ~x331 & ~x332 & ~x335 & ~x361 & ~x377 & ~x388 & ~x390 & ~x392 & ~x404 & ~x405 & ~x406 & ~x415 & ~x416 & ~x420 & ~x421 & ~x432 & ~x443 & ~x445 & ~x446 & ~x448 & ~x450 & ~x460 & ~x471 & ~x488 & ~x498 & ~x499 & ~x501 & ~x502 & ~x503 & ~x514 & ~x515 & ~x534 & ~x536 & ~x542 & ~x543 & ~x555 & ~x558 & ~x566 & ~x567 & ~x569 & ~x570 & ~x583 & ~x585 & ~x586 & ~x589 & ~x593 & ~x594 & ~x595 & ~x596 & ~x616 & ~x620 & ~x624 & ~x639 & ~x641 & ~x643 & ~x645 & ~x652 & ~x667 & ~x697 & ~x698 & ~x699 & ~x703 & ~x705 & ~x706 & ~x725 & ~x728 & ~x738 & ~x757 & ~x758 & ~x772 & ~x779 & ~x780 & ~x781;
assign c7112 =  x294 &  x295 &  x297 &  x298 &  x325 &  x353 & ~x3 & ~x6 & ~x9 & ~x11 & ~x15 & ~x18 & ~x19 & ~x21 & ~x38 & ~x40 & ~x41 & ~x42 & ~x43 & ~x46 & ~x48 & ~x50 & ~x62 & ~x67 & ~x74 & ~x86 & ~x90 & ~x91 & ~x96 & ~x97 & ~x99 & ~x103 & ~x105 & ~x107 & ~x111 & ~x116 & ~x117 & ~x118 & ~x124 & ~x125 & ~x129 & ~x130 & ~x136 & ~x147 & ~x149 & ~x153 & ~x154 & ~x159 & ~x160 & ~x167 & ~x168 & ~x170 & ~x184 & ~x185 & ~x191 & ~x194 & ~x197 & ~x250 & ~x251 & ~x252 & ~x253 & ~x305 & ~x309 & ~x360 & ~x389 & ~x392 & ~x394 & ~x418 & ~x423 & ~x444 & ~x477 & ~x478 & ~x480 & ~x507 & ~x530 & ~x565 & ~x566 & ~x567 & ~x588 & ~x589 & ~x612 & ~x648 & ~x668 & ~x671 & ~x675 & ~x690 & ~x694 & ~x723 & ~x724 & ~x730 & ~x733 & ~x747 & ~x751 & ~x756 & ~x759 & ~x769 & ~x777 & ~x780 & ~x781;
assign c7114 = ~x0 & ~x2 & ~x13 & ~x16 & ~x27 & ~x32 & ~x34 & ~x65 & ~x67 & ~x84 & ~x85 & ~x87 & ~x88 & ~x91 & ~x96 & ~x107 & ~x108 & ~x118 & ~x122 & ~x129 & ~x131 & ~x138 & ~x161 & ~x162 & ~x198 & ~x201 & ~x310 & ~x322 & ~x349 & ~x362 & ~x365 & ~x392 & ~x393 & ~x405 & ~x418 & ~x431 & ~x444 & ~x459 & ~x471 & ~x482 & ~x484 & ~x486 & ~x487 & ~x497 & ~x528 & ~x530 & ~x537 & ~x555 & ~x559 & ~x562 & ~x564 & ~x584 & ~x588 & ~x594 & ~x609 & ~x610 & ~x637 & ~x661 & ~x692 & ~x701 & ~x725 & ~x734 & ~x751 & ~x757 & ~x764 & ~x783;
assign c7116 = ~x0 & ~x3 & ~x4 & ~x5 & ~x6 & ~x7 & ~x9 & ~x11 & ~x13 & ~x19 & ~x25 & ~x27 & ~x29 & ~x30 & ~x33 & ~x35 & ~x37 & ~x41 & ~x45 & ~x48 & ~x50 & ~x51 & ~x57 & ~x58 & ~x60 & ~x63 & ~x66 & ~x71 & ~x75 & ~x82 & ~x83 & ~x86 & ~x91 & ~x93 & ~x94 & ~x108 & ~x109 & ~x111 & ~x112 & ~x116 & ~x120 & ~x121 & ~x122 & ~x123 & ~x124 & ~x126 & ~x130 & ~x137 & ~x140 & ~x142 & ~x146 & ~x164 & ~x166 & ~x167 & ~x190 & ~x191 & ~x195 & ~x200 & ~x217 & ~x219 & ~x225 & ~x227 & ~x247 & ~x254 & ~x280 & ~x322 & ~x333 & ~x338 & ~x339 & ~x349 & ~x359 & ~x389 & ~x393 & ~x419 & ~x432 & ~x433 & ~x445 & ~x446 & ~x451 & ~x460 & ~x500 & ~x504 & ~x505 & ~x511 & ~x512 & ~x528 & ~x530 & ~x531 & ~x538 & ~x544 & ~x556 & ~x557 & ~x564 & ~x566 & ~x582 & ~x585 & ~x587 & ~x593 & ~x595 & ~x596 & ~x598 & ~x614 & ~x615 & ~x619 & ~x622 & ~x626 & ~x643 & ~x645 & ~x646 & ~x649 & ~x651 & ~x652 & ~x655 & ~x670 & ~x671 & ~x673 & ~x674 & ~x675 & ~x678 & ~x694 & ~x696 & ~x703 & ~x708 & ~x728 & ~x729 & ~x730 & ~x731 & ~x732 & ~x735 & ~x737 & ~x754 & ~x756 & ~x759 & ~x760 & ~x761 & ~x763 & ~x769 & ~x772 & ~x775 & ~x778;
assign c7118 =  x164;
assign c7120 =  x346 & ~x26 & ~x30 & ~x91 & ~x102 & ~x117 & ~x124 & ~x132 & ~x146 & ~x149 & ~x150 & ~x164 & ~x172 & ~x178 & ~x198 & ~x202 & ~x227 & ~x281 & ~x364 & ~x365 & ~x377 & ~x405 & ~x415 & ~x417 & ~x419 & ~x441 & ~x450 & ~x460 & ~x476 & ~x484 & ~x498 & ~x510 & ~x527 & ~x538 & ~x566 & ~x580 & ~x587 & ~x592 & ~x595 & ~x639 & ~x642 & ~x662 & ~x672 & ~x719 & ~x722 & ~x759 & ~x763 & ~x770 & ~x773 & ~x775;
assign c7122 =  x237 &  x238 &  x437 & ~x9 & ~x10 & ~x31 & ~x34 & ~x36 & ~x38 & ~x39 & ~x50 & ~x53 & ~x54 & ~x63 & ~x68 & ~x74 & ~x86 & ~x90 & ~x97 & ~x104 & ~x125 & ~x128 & ~x132 & ~x136 & ~x138 & ~x142 & ~x143 & ~x162 & ~x165 & ~x194 & ~x195 & ~x198 & ~x199 & ~x279 & ~x284 & ~x304 & ~x342 & ~x360 & ~x361 & ~x367 & ~x378 & ~x405 & ~x417 & ~x419 & ~x421 & ~x434 & ~x446 & ~x450 & ~x451 & ~x468 & ~x470 & ~x473 & ~x475 & ~x498 & ~x510 & ~x524 & ~x543 & ~x551 & ~x558 & ~x571 & ~x580 & ~x596 & ~x607 & ~x611 & ~x612 & ~x622 & ~x669 & ~x674 & ~x679 & ~x692 & ~x704 & ~x729 & ~x730 & ~x731 & ~x749 & ~x751 & ~x760 & ~x778 & ~x780;
assign c7124 =  x44;
assign c7126 = ~x15 & ~x19 & ~x21 & ~x25 & ~x28 & ~x29 & ~x32 & ~x46 & ~x56 & ~x58 & ~x59 & ~x61 & ~x80 & ~x89 & ~x93 & ~x98 & ~x99 & ~x110 & ~x124 & ~x132 & ~x136 & ~x138 & ~x145 & ~x147 & ~x148 & ~x149 & ~x152 & ~x156 & ~x160 & ~x168 & ~x170 & ~x171 & ~x173 & ~x195 & ~x219 & ~x223 & ~x224 & ~x225 & ~x279 & ~x303 & ~x342 & ~x365 & ~x378 & ~x392 & ~x398 & ~x405 & ~x406 & ~x433 & ~x447 & ~x449 & ~x451 & ~x460 & ~x461 & ~x470 & ~x473 & ~x477 & ~x479 & ~x480 & ~x482 & ~x488 & ~x507 & ~x524 & ~x529 & ~x553 & ~x554 & ~x570 & ~x580 & ~x581 & ~x592 & ~x597 & ~x598 & ~x610 & ~x612 & ~x620 & ~x640 & ~x643 & ~x648 & ~x651 & ~x664 & ~x672 & ~x677 & ~x723 & ~x727 & ~x754 & ~x755 & ~x762;
assign c7128 = ~x8 & ~x14 & ~x19 & ~x22 & ~x28 & ~x38 & ~x42 & ~x46 & ~x47 & ~x48 & ~x52 & ~x53 & ~x56 & ~x60 & ~x66 & ~x68 & ~x73 & ~x75 & ~x82 & ~x84 & ~x85 & ~x86 & ~x87 & ~x88 & ~x90 & ~x91 & ~x99 & ~x102 & ~x105 & ~x112 & ~x125 & ~x127 & ~x134 & ~x142 & ~x146 & ~x150 & ~x153 & ~x167 & ~x170 & ~x175 & ~x220 & ~x221 & ~x224 & ~x251 & ~x253 & ~x280 & ~x283 & ~x303 & ~x310 & ~x333 & ~x365 & ~x377 & ~x405 & ~x417 & ~x419 & ~x420 & ~x421 & ~x432 & ~x443 & ~x448 & ~x449 & ~x459 & ~x461 & ~x471 & ~x476 & ~x478 & ~x487 & ~x488 & ~x506 & ~x525 & ~x532 & ~x534 & ~x535 & ~x539 & ~x542 & ~x543 & ~x553 & ~x556 & ~x557 & ~x562 & ~x565 & ~x582 & ~x585 & ~x587 & ~x589 & ~x590 & ~x591 & ~x594 & ~x617 & ~x618 & ~x642 & ~x645 & ~x646 & ~x647 & ~x666 & ~x669 & ~x675 & ~x677 & ~x680 & ~x696 & ~x700 & ~x702 & ~x703 & ~x705 & ~x707 & ~x708 & ~x715 & ~x729 & ~x734 & ~x760 & ~x761 & ~x763 & ~x768 & ~x770;
assign c7130 =  x240 &  x464 &  x520 & ~x2 & ~x6 & ~x16 & ~x19 & ~x27 & ~x36 & ~x44 & ~x48 & ~x49 & ~x67 & ~x70 & ~x73 & ~x83 & ~x90 & ~x116 & ~x121 & ~x131 & ~x133 & ~x136 & ~x139 & ~x160 & ~x161 & ~x224 & ~x275 & ~x316 & ~x317 & ~x319 & ~x334 & ~x343 & ~x363 & ~x369 & ~x371 & ~x372 & ~x374 & ~x375 & ~x386 & ~x391 & ~x397 & ~x414 & ~x443 & ~x451 & ~x452 & ~x473 & ~x476 & ~x479 & ~x508 & ~x532 & ~x536 & ~x560 & ~x582 & ~x588 & ~x593 & ~x611 & ~x620 & ~x622 & ~x624 & ~x625 & ~x626 & ~x641 & ~x643 & ~x645 & ~x647 & ~x652 & ~x655 & ~x665 & ~x666 & ~x675 & ~x678 & ~x680 & ~x682 & ~x683 & ~x694 & ~x705 & ~x730 & ~x737 & ~x747 & ~x756 & ~x757 & ~x758 & ~x759 & ~x762 & ~x763 & ~x766;
assign c7132 =  x339;
assign c7134 =  x208 &  x209 &  x352 &  x435 & ~x6 & ~x17 & ~x23 & ~x25 & ~x26 & ~x27 & ~x33 & ~x36 & ~x48 & ~x57 & ~x65 & ~x74 & ~x75 & ~x89 & ~x92 & ~x94 & ~x101 & ~x105 & ~x112 & ~x113 & ~x119 & ~x125 & ~x128 & ~x134 & ~x145 & ~x146 & ~x147 & ~x168 & ~x174 & ~x196 & ~x200 & ~x220 & ~x229 & ~x249 & ~x273 & ~x274 & ~x284 & ~x285 & ~x292 & ~x293 & ~x300 & ~x302 & ~x321 & ~x339 & ~x349 & ~x389 & ~x396 & ~x418 & ~x422 & ~x443 & ~x444 & ~x447 & ~x451 & ~x481 & ~x513 & ~x528 & ~x536 & ~x562 & ~x577 & ~x593 & ~x605 & ~x611 & ~x636 & ~x639 & ~x640 & ~x650 & ~x661 & ~x667 & ~x668 & ~x676 & ~x697 & ~x701 & ~x710 & ~x721 & ~x725 & ~x740 & ~x743 & ~x749 & ~x758 & ~x772 & ~x775 & ~x777;
assign c7136 = ~x13 & ~x28 & ~x37 & ~x46 & ~x57 & ~x61 & ~x68 & ~x76 & ~x77 & ~x80 & ~x102 & ~x106 & ~x110 & ~x114 & ~x122 & ~x134 & ~x155 & ~x157 & ~x171 & ~x196 & ~x219 & ~x277 & ~x278 & ~x287 & ~x303 & ~x305 & ~x331 & ~x336 & ~x340 & ~x358 & ~x359 & ~x360 & ~x362 & ~x364 & ~x377 & ~x391 & ~x392 & ~x405 & ~x433 & ~x448 & ~x457 & ~x461 & ~x480 & ~x513 & ~x530 & ~x536 & ~x551 & ~x552 & ~x569 & ~x585 & ~x593 & ~x594 & ~x614 & ~x615 & ~x617 & ~x641 & ~x661 & ~x689 & ~x721 & ~x734 & ~x747 & ~x753 & ~x769 & ~x774 & ~x782;
assign c7138 =  x207 &  x461 &  x517 & ~x4 & ~x7 & ~x9 & ~x14 & ~x15 & ~x22 & ~x23 & ~x24 & ~x45 & ~x51 & ~x53 & ~x58 & ~x59 & ~x68 & ~x69 & ~x72 & ~x74 & ~x75 & ~x78 & ~x79 & ~x80 & ~x81 & ~x89 & ~x97 & ~x106 & ~x108 & ~x113 & ~x122 & ~x124 & ~x125 & ~x127 & ~x130 & ~x132 & ~x141 & ~x143 & ~x144 & ~x158 & ~x161 & ~x164 & ~x170 & ~x191 & ~x192 & ~x195 & ~x200 & ~x224 & ~x230 & ~x246 & ~x250 & ~x254 & ~x255 & ~x277 & ~x292 & ~x302 & ~x306 & ~x307 & ~x308 & ~x312 & ~x315 & ~x317 & ~x318 & ~x329 & ~x330 & ~x331 & ~x334 & ~x337 & ~x339 & ~x340 & ~x360 & ~x361 & ~x362 & ~x363 & ~x366 & ~x371 & ~x389 & ~x390 & ~x392 & ~x395 & ~x415 & ~x417 & ~x420 & ~x448 & ~x449 & ~x476 & ~x479 & ~x506 & ~x526 & ~x528 & ~x531 & ~x532 & ~x535 & ~x538 & ~x551 & ~x563 & ~x581 & ~x585 & ~x587 & ~x588 & ~x589 & ~x590 & ~x591 & ~x592 & ~x606 & ~x612 & ~x615 & ~x616 & ~x621 & ~x636 & ~x639 & ~x647 & ~x663 & ~x667 & ~x669 & ~x673 & ~x674 & ~x675 & ~x676 & ~x678 & ~x692 & ~x700 & ~x701 & ~x708 & ~x716 & ~x720 & ~x721 & ~x723 & ~x724 & ~x733 & ~x744 & ~x767 & ~x780 & ~x781 & ~x783;
assign c7140 =  x435 & ~x0 & ~x11 & ~x14 & ~x20 & ~x24 & ~x30 & ~x34 & ~x40 & ~x49 & ~x54 & ~x56 & ~x57 & ~x60 & ~x92 & ~x93 & ~x96 & ~x99 & ~x100 & ~x108 & ~x111 & ~x124 & ~x135 & ~x158 & ~x160 & ~x163 & ~x165 & ~x167 & ~x170 & ~x173 & ~x203 & ~x222 & ~x250 & ~x305 & ~x308 & ~x342 & ~x350 & ~x387 & ~x390 & ~x397 & ~x404 & ~x420 & ~x431 & ~x445 & ~x452 & ~x455 & ~x472 & ~x496 & ~x503 & ~x509 & ~x534 & ~x563 & ~x564 & ~x566 & ~x577 & ~x579 & ~x587 & ~x589 & ~x591 & ~x609 & ~x610 & ~x619 & ~x634 & ~x636 & ~x643 & ~x646 & ~x664 & ~x671 & ~x672 & ~x693 & ~x717 & ~x724 & ~x743 & ~x750 & ~x752 & ~x753 & ~x766 & ~x772 & ~x779;
assign c7142 =  x738;
assign c7144 =  x380 &  x461 &  x489 & ~x4 & ~x5 & ~x7 & ~x8 & ~x18 & ~x32 & ~x36 & ~x72 & ~x84 & ~x87 & ~x89 & ~x91 & ~x96 & ~x101 & ~x104 & ~x128 & ~x142 & ~x145 & ~x147 & ~x160 & ~x162 & ~x163 & ~x170 & ~x226 & ~x228 & ~x250 & ~x252 & ~x254 & ~x256 & ~x282 & ~x283 & ~x284 & ~x308 & ~x309 & ~x311 & ~x312 & ~x339 & ~x340 & ~x347 & ~x349 & ~x350 & ~x367 & ~x368 & ~x372 & ~x375 & ~x376 & ~x395 & ~x397 & ~x422 & ~x452 & ~x476 & ~x478 & ~x500 & ~x503 & ~x504 & ~x531 & ~x534 & ~x556 & ~x576 & ~x577 & ~x578 & ~x603 & ~x604 & ~x605 & ~x606 & ~x616 & ~x619 & ~x634 & ~x644 & ~x645 & ~x646 & ~x663 & ~x687 & ~x688 & ~x701 & ~x702 & ~x703 & ~x716 & ~x722 & ~x727 & ~x739 & ~x745 & ~x747 & ~x748 & ~x750 & ~x766 & ~x772 & ~x774 & ~x775 & ~x776 & ~x778 & ~x781;
assign c7146 =  x269 &  x407 &  x462 &  x489 &  x545 &  x572 &  x628 &  x683 & ~x8 & ~x18 & ~x25 & ~x28 & ~x58 & ~x72 & ~x80 & ~x85 & ~x86 & ~x89 & ~x91 & ~x115 & ~x157 & ~x158 & ~x160 & ~x162 & ~x171 & ~x304 & ~x338 & ~x362 & ~x366 & ~x367 & ~x450 & ~x478 & ~x501 & ~x502 & ~x528 & ~x538 & ~x560 & ~x561 & ~x562 & ~x576 & ~x579 & ~x593 & ~x607 & ~x616 & ~x635 & ~x646 & ~x661 & ~x664 & ~x670 & ~x688 & ~x689 & ~x703 & ~x722 & ~x734 & ~x754 & ~x757 & ~x763 & ~x767 & ~x770 & ~x779;
assign c7148 = ~x6 & ~x9 & ~x23 & ~x26 & ~x36 & ~x38 & ~x42 & ~x43 & ~x45 & ~x70 & ~x74 & ~x87 & ~x92 & ~x104 & ~x110 & ~x125 & ~x127 & ~x133 & ~x134 & ~x143 & ~x162 & ~x166 & ~x169 & ~x221 & ~x223 & ~x248 & ~x277 & ~x305 & ~x309 & ~x310 & ~x319 & ~x321 & ~x322 & ~x333 & ~x334 & ~x346 & ~x350 & ~x359 & ~x364 & ~x368 & ~x375 & ~x376 & ~x404 & ~x405 & ~x418 & ~x429 & ~x431 & ~x447 & ~x450 & ~x452 & ~x455 & ~x471 & ~x473 & ~x478 & ~x481 & ~x506 & ~x533 & ~x561 & ~x562 & ~x563 & ~x567 & ~x592 & ~x607 & ~x609 & ~x614 & ~x618 & ~x636 & ~x661 & ~x666 & ~x670 & ~x692 & ~x695 & ~x700 & ~x701 & ~x725 & ~x726 & ~x732 & ~x744 & ~x746 & ~x749 & ~x766 & ~x769 & ~x771 & ~x774 & ~x776 & ~x783;
assign c7150 =  x87;
assign c7152 =  x705;
assign c7154 =  x708;
assign c7156 =  x259 &  x289 & ~x4 & ~x7 & ~x8 & ~x9 & ~x11 & ~x13 & ~x17 & ~x19 & ~x20 & ~x27 & ~x28 & ~x30 & ~x31 & ~x39 & ~x43 & ~x45 & ~x48 & ~x49 & ~x54 & ~x56 & ~x57 & ~x59 & ~x61 & ~x64 & ~x65 & ~x66 & ~x72 & ~x73 & ~x78 & ~x80 & ~x81 & ~x83 & ~x87 & ~x88 & ~x89 & ~x93 & ~x95 & ~x97 & ~x98 & ~x102 & ~x105 & ~x109 & ~x111 & ~x114 & ~x116 & ~x120 & ~x121 & ~x124 & ~x125 & ~x129 & ~x132 & ~x136 & ~x139 & ~x141 & ~x142 & ~x145 & ~x146 & ~x147 & ~x149 & ~x151 & ~x153 & ~x154 & ~x155 & ~x156 & ~x157 & ~x161 & ~x165 & ~x166 & ~x192 & ~x193 & ~x195 & ~x222 & ~x247 & ~x250 & ~x276 & ~x278 & ~x305 & ~x307 & ~x308 & ~x330 & ~x339 & ~x358 & ~x359 & ~x361 & ~x365 & ~x366 & ~x367 & ~x376 & ~x377 & ~x387 & ~x389 & ~x417 & ~x418 & ~x421 & ~x422 & ~x447 & ~x449 & ~x473 & ~x474 & ~x478 & ~x480 & ~x500 & ~x501 & ~x505 & ~x533 & ~x534 & ~x536 & ~x537 & ~x538 & ~x555 & ~x557 & ~x558 & ~x562 & ~x566 & ~x568 & ~x569 & ~x571 & ~x583 & ~x584 & ~x585 & ~x587 & ~x588 & ~x589 & ~x591 & ~x592 & ~x594 & ~x597 & ~x598 & ~x599 & ~x614 & ~x616 & ~x618 & ~x622 & ~x623 & ~x626 & ~x639 & ~x641 & ~x646 & ~x648 & ~x652 & ~x665 & ~x666 & ~x667 & ~x671 & ~x679 & ~x681 & ~x696 & ~x702 & ~x703 & ~x704 & ~x709 & ~x710 & ~x728 & ~x734 & ~x750 & ~x752 & ~x754 & ~x755 & ~x758 & ~x760 & ~x762 & ~x765 & ~x769 & ~x774 & ~x776 & ~x779 & ~x780 & ~x781 & ~x782;
assign c7158 =  x240 &  x261 & ~x12 & ~x14 & ~x22 & ~x26 & ~x31 & ~x34 & ~x38 & ~x47 & ~x53 & ~x57 & ~x59 & ~x64 & ~x73 & ~x77 & ~x85 & ~x92 & ~x93 & ~x94 & ~x99 & ~x101 & ~x102 & ~x103 & ~x107 & ~x108 & ~x110 & ~x118 & ~x120 & ~x128 & ~x129 & ~x130 & ~x137 & ~x139 & ~x140 & ~x141 & ~x147 & ~x150 & ~x153 & ~x154 & ~x159 & ~x225 & ~x249 & ~x251 & ~x277 & ~x283 & ~x305 & ~x306 & ~x307 & ~x311 & ~x335 & ~x338 & ~x339 & ~x359 & ~x360 & ~x361 & ~x369 & ~x375 & ~x376 & ~x385 & ~x390 & ~x394 & ~x397 & ~x420 & ~x425 & ~x450 & ~x451 & ~x473 & ~x479 & ~x501 & ~x531 & ~x533 & ~x536 & ~x549 & ~x550 & ~x554 & ~x563 & ~x577 & ~x578 & ~x581 & ~x582 & ~x585 & ~x588 & ~x610 & ~x613 & ~x616 & ~x618 & ~x622 & ~x639 & ~x642 & ~x645 & ~x664 & ~x691 & ~x692 & ~x696 & ~x701 & ~x702 & ~x720 & ~x724 & ~x731 & ~x733 & ~x738 & ~x748 & ~x753 & ~x756 & ~x767 & ~x771 & ~x773 & ~x779 & ~x780;
assign c7160 =  x259 &  x463 &  x519 & ~x2 & ~x8 & ~x32 & ~x41 & ~x46 & ~x56 & ~x58 & ~x76 & ~x86 & ~x88 & ~x95 & ~x101 & ~x110 & ~x114 & ~x121 & ~x134 & ~x137 & ~x152 & ~x161 & ~x217 & ~x274 & ~x275 & ~x301 & ~x336 & ~x338 & ~x367 & ~x368 & ~x389 & ~x394 & ~x395 & ~x417 & ~x418 & ~x420 & ~x450 & ~x506 & ~x527 & ~x528 & ~x532 & ~x534 & ~x536 & ~x553 & ~x556 & ~x566 & ~x580 & ~x582 & ~x584 & ~x586 & ~x598 & ~x606 & ~x610 & ~x625 & ~x635 & ~x646 & ~x664 & ~x667 & ~x669 & ~x672 & ~x674 & ~x678 & ~x699 & ~x727 & ~x730 & ~x733 & ~x734 & ~x750 & ~x761 & ~x781;
assign c7162 =  x145;
assign c7164 =  x285 & ~x156 & ~x398 & ~x420 & ~x543 & ~x554;
assign c7166 =  x340;
assign c7168 = ~x0 & ~x2 & ~x10 & ~x12 & ~x18 & ~x19 & ~x21 & ~x23 & ~x24 & ~x26 & ~x32 & ~x33 & ~x35 & ~x36 & ~x38 & ~x42 & ~x43 & ~x44 & ~x46 & ~x51 & ~x57 & ~x65 & ~x72 & ~x74 & ~x75 & ~x76 & ~x77 & ~x79 & ~x81 & ~x84 & ~x85 & ~x86 & ~x88 & ~x90 & ~x92 & ~x94 & ~x96 & ~x97 & ~x98 & ~x101 & ~x107 & ~x112 & ~x113 & ~x114 & ~x115 & ~x117 & ~x123 & ~x124 & ~x125 & ~x127 & ~x128 & ~x129 & ~x131 & ~x134 & ~x136 & ~x137 & ~x141 & ~x143 & ~x145 & ~x146 & ~x147 & ~x150 & ~x155 & ~x158 & ~x160 & ~x161 & ~x162 & ~x165 & ~x166 & ~x167 & ~x171 & ~x175 & ~x187 & ~x188 & ~x191 & ~x192 & ~x220 & ~x222 & ~x247 & ~x249 & ~x251 & ~x253 & ~x275 & ~x276 & ~x279 & ~x280 & ~x282 & ~x307 & ~x308 & ~x309 & ~x332 & ~x333 & ~x335 & ~x363 & ~x367 & ~x377 & ~x378 & ~x391 & ~x393 & ~x405 & ~x406 & ~x417 & ~x432 & ~x444 & ~x446 & ~x448 & ~x449 & ~x451 & ~x452 & ~x471 & ~x472 & ~x473 & ~x475 & ~x480 & ~x487 & ~x489 & ~x499 & ~x500 & ~x501 & ~x502 & ~x503 & ~x505 & ~x506 & ~x508 & ~x514 & ~x515 & ~x527 & ~x529 & ~x530 & ~x531 & ~x534 & ~x535 & ~x537 & ~x538 & ~x541 & ~x542 & ~x555 & ~x556 & ~x561 & ~x563 & ~x565 & ~x567 & ~x568 & ~x570 & ~x581 & ~x583 & ~x585 & ~x588 & ~x590 & ~x591 & ~x592 & ~x595 & ~x596 & ~x597 & ~x611 & ~x612 & ~x613 & ~x618 & ~x621 & ~x623 & ~x639 & ~x641 & ~x644 & ~x645 & ~x652 & ~x654 & ~x667 & ~x671 & ~x672 & ~x674 & ~x675 & ~x680 & ~x681 & ~x694 & ~x697 & ~x700 & ~x703 & ~x705 & ~x708 & ~x729 & ~x730 & ~x733 & ~x734 & ~x738 & ~x739 & ~x740 & ~x749 & ~x759 & ~x761 & ~x762 & ~x763 & ~x766 & ~x767 & ~x769 & ~x772 & ~x777 & ~x779 & ~x782 & ~x783;
assign c7170 =  x389;
assign c7172 =  x236 & ~x1 & ~x5 & ~x13 & ~x14 & ~x15 & ~x25 & ~x43 & ~x45 & ~x56 & ~x59 & ~x60 & ~x63 & ~x65 & ~x69 & ~x72 & ~x77 & ~x78 & ~x82 & ~x83 & ~x84 & ~x86 & ~x91 & ~x92 & ~x99 & ~x103 & ~x113 & ~x117 & ~x119 & ~x120 & ~x121 & ~x123 & ~x124 & ~x125 & ~x129 & ~x132 & ~x133 & ~x134 & ~x135 & ~x139 & ~x141 & ~x142 & ~x145 & ~x147 & ~x152 & ~x154 & ~x161 & ~x163 & ~x164 & ~x173 & ~x190 & ~x192 & ~x195 & ~x197 & ~x198 & ~x201 & ~x227 & ~x251 & ~x254 & ~x280 & ~x281 & ~x282 & ~x285 & ~x303 & ~x305 & ~x310 & ~x311 & ~x312 & ~x314 & ~x318 & ~x319 & ~x330 & ~x333 & ~x335 & ~x336 & ~x345 & ~x346 & ~x359 & ~x363 & ~x365 & ~x366 & ~x368 & ~x391 & ~x395 & ~x397 & ~x419 & ~x422 & ~x445 & ~x447 & ~x448 & ~x451 & ~x452 & ~x453 & ~x455 & ~x477 & ~x479 & ~x482 & ~x498 & ~x500 & ~x501 & ~x503 & ~x507 & ~x523 & ~x538 & ~x539 & ~x549 & ~x553 & ~x554 & ~x555 & ~x566 & ~x579 & ~x582 & ~x589 & ~x594 & ~x605 & ~x606 & ~x608 & ~x609 & ~x612 & ~x619 & ~x620 & ~x639 & ~x641 & ~x645 & ~x646 & ~x648 & ~x664 & ~x668 & ~x690 & ~x695 & ~x697 & ~x702 & ~x730 & ~x731 & ~x732 & ~x734 & ~x735 & ~x736 & ~x742 & ~x745 & ~x746 & ~x750 & ~x755 & ~x757 & ~x758 & ~x759 & ~x761 & ~x770 & ~x771 & ~x774 & ~x777 & ~x782;
assign c7174 =  x678;
assign c7176 =  x65;
assign c7178 =  x205 &  x491 &  x546 & ~x3 & ~x95 & ~x104 & ~x134 & ~x162 & ~x189 & ~x255 & ~x278 & ~x347 & ~x392 & ~x395 & ~x421 & ~x422 & ~x527 & ~x559 & ~x582 & ~x598 & ~x640 & ~x644 & ~x645 & ~x651 & ~x679 & ~x690 & ~x704 & ~x722 & ~x744;
assign c7180 =  x265 &  x267 &  x268 &  x296 & ~x44 & ~x54 & ~x70 & ~x74 & ~x86 & ~x145 & ~x152 & ~x159 & ~x182 & ~x209 & ~x251 & ~x333 & ~x370 & ~x371 & ~x373 & ~x398 & ~x399 & ~x502 & ~x503 & ~x510 & ~x584 & ~x590 & ~x636 & ~x642 & ~x703 & ~x777 & ~x781;
assign c7182 =  x269 & ~x1 & ~x19 & ~x26 & ~x33 & ~x34 & ~x37 & ~x43 & ~x44 & ~x46 & ~x47 & ~x76 & ~x92 & ~x109 & ~x117 & ~x138 & ~x155 & ~x157 & ~x158 & ~x162 & ~x167 & ~x198 & ~x219 & ~x256 & ~x274 & ~x310 & ~x311 & ~x313 & ~x334 & ~x342 & ~x346 & ~x357 & ~x359 & ~x362 & ~x373 & ~x393 & ~x419 & ~x423 & ~x449 & ~x455 & ~x501 & ~x508 & ~x510 & ~x524 & ~x550 & ~x555 & ~x576 & ~x579 & ~x583 & ~x594 & ~x595 & ~x612 & ~x618 & ~x639 & ~x640 & ~x665 & ~x666 & ~x671 & ~x681 & ~x688 & ~x689 & ~x723 & ~x747 & ~x753 & ~x756 & ~x759 & ~x770 & ~x772 & ~x783;
assign c7184 =  x279;
assign c7186 = ~x1 & ~x6 & ~x11 & ~x20 & ~x26 & ~x28 & ~x30 & ~x49 & ~x50 & ~x61 & ~x69 & ~x94 & ~x95 & ~x99 & ~x105 & ~x111 & ~x126 & ~x130 & ~x198 & ~x201 & ~x254 & ~x323 & ~x333 & ~x339 & ~x340 & ~x349 & ~x350 & ~x358 & ~x361 & ~x364 & ~x367 & ~x375 & ~x376 & ~x395 & ~x400 & ~x402 & ~x403 & ~x427 & ~x447 & ~x450 & ~x451 & ~x455 & ~x468 & ~x479 & ~x480 & ~x526 & ~x528 & ~x531 & ~x534 & ~x551 & ~x552 & ~x553 & ~x559 & ~x560 & ~x589 & ~x632 & ~x633 & ~x636 & ~x637 & ~x643 & ~x659 & ~x686 & ~x690 & ~x691 & ~x699 & ~x722 & ~x776 & ~x777;
assign c7188 =  x310;
assign c7190 = ~x0 & ~x2 & ~x3 & ~x5 & ~x8 & ~x16 & ~x17 & ~x19 & ~x25 & ~x34 & ~x35 & ~x49 & ~x50 & ~x52 & ~x54 & ~x57 & ~x60 & ~x65 & ~x74 & ~x78 & ~x79 & ~x81 & ~x84 & ~x85 & ~x87 & ~x89 & ~x106 & ~x111 & ~x116 & ~x117 & ~x118 & ~x120 & ~x144 & ~x146 & ~x161 & ~x169 & ~x174 & ~x193 & ~x200 & ~x227 & ~x228 & ~x252 & ~x276 & ~x280 & ~x281 & ~x282 & ~x285 & ~x304 & ~x315 & ~x317 & ~x319 & ~x321 & ~x330 & ~x332 & ~x337 & ~x338 & ~x341 & ~x345 & ~x346 & ~x350 & ~x360 & ~x361 & ~x371 & ~x388 & ~x390 & ~x392 & ~x394 & ~x399 & ~x414 & ~x421 & ~x427 & ~x451 & ~x477 & ~x501 & ~x506 & ~x524 & ~x527 & ~x530 & ~x531 & ~x532 & ~x551 & ~x553 & ~x554 & ~x561 & ~x565 & ~x567 & ~x576 & ~x577 & ~x579 & ~x588 & ~x590 & ~x592 & ~x607 & ~x608 & ~x609 & ~x615 & ~x617 & ~x621 & ~x632 & ~x633 & ~x639 & ~x641 & ~x645 & ~x666 & ~x667 & ~x668 & ~x672 & ~x687 & ~x689 & ~x690 & ~x694 & ~x695 & ~x702 & ~x720 & ~x727 & ~x734 & ~x744 & ~x750 & ~x752 & ~x753 & ~x758 & ~x762 & ~x767 & ~x771 & ~x773 & ~x778 & ~x781;
assign c7192 =  x206 &  x235 &  x521 & ~x2 & ~x4 & ~x11 & ~x12 & ~x13 & ~x14 & ~x20 & ~x37 & ~x44 & ~x53 & ~x59 & ~x67 & ~x68 & ~x73 & ~x76 & ~x87 & ~x92 & ~x102 & ~x109 & ~x110 & ~x138 & ~x152 & ~x166 & ~x220 & ~x337 & ~x340 & ~x347 & ~x349 & ~x367 & ~x376 & ~x424 & ~x432 & ~x443 & ~x505 & ~x531 & ~x559 & ~x560 & ~x562 & ~x584 & ~x586 & ~x621 & ~x666 & ~x667 & ~x671 & ~x673 & ~x680 & ~x700 & ~x701 & ~x751 & ~x757 & ~x760;
assign c7194 = ~x0 & ~x1 & ~x2 & ~x4 & ~x5 & ~x6 & ~x13 & ~x17 & ~x19 & ~x22 & ~x25 & ~x28 & ~x30 & ~x33 & ~x41 & ~x42 & ~x43 & ~x45 & ~x48 & ~x55 & ~x57 & ~x59 & ~x60 & ~x63 & ~x69 & ~x72 & ~x75 & ~x80 & ~x81 & ~x82 & ~x83 & ~x86 & ~x87 & ~x88 & ~x93 & ~x94 & ~x98 & ~x99 & ~x100 & ~x101 & ~x102 & ~x104 & ~x105 & ~x106 & ~x109 & ~x111 & ~x112 & ~x113 & ~x116 & ~x121 & ~x124 & ~x131 & ~x135 & ~x142 & ~x144 & ~x146 & ~x147 & ~x148 & ~x150 & ~x153 & ~x154 & ~x155 & ~x158 & ~x159 & ~x161 & ~x169 & ~x170 & ~x172 & ~x189 & ~x191 & ~x192 & ~x195 & ~x196 & ~x198 & ~x219 & ~x220 & ~x224 & ~x225 & ~x249 & ~x278 & ~x279 & ~x281 & ~x284 & ~x304 & ~x306 & ~x308 & ~x310 & ~x311 & ~x332 & ~x333 & ~x335 & ~x338 & ~x349 & ~x350 & ~x360 & ~x362 & ~x364 & ~x365 & ~x366 & ~x368 & ~x377 & ~x379 & ~x389 & ~x391 & ~x392 & ~x394 & ~x395 & ~x406 & ~x416 & ~x419 & ~x420 & ~x423 & ~x424 & ~x433 & ~x434 & ~x445 & ~x446 & ~x448 & ~x452 & ~x461 & ~x471 & ~x472 & ~x475 & ~x478 & ~x488 & ~x500 & ~x506 & ~x528 & ~x534 & ~x544 & ~x555 & ~x558 & ~x563 & ~x566 & ~x567 & ~x582 & ~x584 & ~x586 & ~x590 & ~x591 & ~x594 & ~x596 & ~x599 & ~x610 & ~x612 & ~x613 & ~x614 & ~x615 & ~x620 & ~x622 & ~x624 & ~x625 & ~x626 & ~x639 & ~x640 & ~x645 & ~x646 & ~x654 & ~x667 & ~x670 & ~x671 & ~x673 & ~x674 & ~x676 & ~x677 & ~x678 & ~x681 & ~x682 & ~x696 & ~x698 & ~x700 & ~x705 & ~x723 & ~x725 & ~x727 & ~x732 & ~x734 & ~x736 & ~x737 & ~x738 & ~x751 & ~x752 & ~x754 & ~x760 & ~x762 & ~x764 & ~x766 & ~x767 & ~x771 & ~x779 & ~x780;
assign c7196 =  x325 & ~x2 & ~x4 & ~x7 & ~x9 & ~x10 & ~x17 & ~x18 & ~x28 & ~x32 & ~x44 & ~x45 & ~x55 & ~x56 & ~x62 & ~x67 & ~x80 & ~x83 & ~x87 & ~x89 & ~x92 & ~x94 & ~x95 & ~x103 & ~x106 & ~x107 & ~x108 & ~x112 & ~x113 & ~x117 & ~x119 & ~x127 & ~x129 & ~x140 & ~x141 & ~x142 & ~x144 & ~x147 & ~x150 & ~x159 & ~x160 & ~x163 & ~x170 & ~x171 & ~x189 & ~x190 & ~x191 & ~x192 & ~x221 & ~x224 & ~x226 & ~x248 & ~x249 & ~x252 & ~x276 & ~x281 & ~x315 & ~x316 & ~x337 & ~x362 & ~x366 & ~x389 & ~x390 & ~x418 & ~x423 & ~x425 & ~x427 & ~x445 & ~x447 & ~x449 & ~x452 & ~x454 & ~x455 & ~x473 & ~x477 & ~x479 & ~x480 & ~x494 & ~x503 & ~x504 & ~x506 & ~x533 & ~x535 & ~x553 & ~x555 & ~x564 & ~x575 & ~x579 & ~x580 & ~x583 & ~x584 & ~x587 & ~x588 & ~x590 & ~x603 & ~x612 & ~x613 & ~x614 & ~x632 & ~x635 & ~x646 & ~x664 & ~x667 & ~x671 & ~x672 & ~x675 & ~x691 & ~x698 & ~x703 & ~x706 & ~x722 & ~x726 & ~x728 & ~x741 & ~x742 & ~x751 & ~x753 & ~x757 & ~x762 & ~x764 & ~x765 & ~x775 & ~x776 & ~x778 & ~x779 & ~x782;
assign c7198 =  x729;
assign c7200 = ~x14 & ~x15 & ~x19 & ~x24 & ~x25 & ~x29 & ~x32 & ~x34 & ~x36 & ~x37 & ~x39 & ~x44 & ~x46 & ~x47 & ~x53 & ~x59 & ~x63 & ~x67 & ~x82 & ~x83 & ~x88 & ~x89 & ~x95 & ~x96 & ~x97 & ~x100 & ~x102 & ~x109 & ~x117 & ~x119 & ~x125 & ~x127 & ~x131 & ~x138 & ~x143 & ~x148 & ~x149 & ~x153 & ~x154 & ~x156 & ~x158 & ~x160 & ~x162 & ~x175 & ~x178 & ~x185 & ~x190 & ~x191 & ~x197 & ~x208 & ~x210 & ~x211 & ~x212 & ~x221 & ~x222 & ~x226 & ~x246 & ~x253 & ~x277 & ~x303 & ~x335 & ~x336 & ~x362 & ~x364 & ~x394 & ~x396 & ~x421 & ~x445 & ~x450 & ~x452 & ~x473 & ~x476 & ~x502 & ~x506 & ~x508 & ~x509 & ~x510 & ~x514 & ~x532 & ~x536 & ~x537 & ~x539 & ~x543 & ~x554 & ~x555 & ~x568 & ~x586 & ~x587 & ~x588 & ~x597 & ~x598 & ~x611 & ~x614 & ~x617 & ~x619 & ~x623 & ~x626 & ~x638 & ~x644 & ~x645 & ~x646 & ~x652 & ~x672 & ~x677 & ~x694 & ~x700 & ~x701 & ~x723 & ~x730 & ~x734 & ~x753 & ~x754 & ~x758 & ~x760 & ~x761 & ~x762 & ~x768 & ~x769 & ~x772 & ~x781;
assign c7202 =  x328 & ~x29 & ~x37 & ~x55 & ~x65 & ~x91 & ~x95 & ~x156 & ~x157 & ~x160 & ~x192 & ~x279 & ~x362 & ~x378 & ~x422 & ~x432 & ~x445 & ~x446 & ~x481 & ~x485 & ~x486 & ~x504 & ~x511 & ~x512 & ~x532 & ~x578 & ~x584 & ~x605 & ~x616 & ~x618 & ~x641 & ~x644 & ~x725 & ~x756 & ~x757;
assign c7204 =  x270 &  x295 &  x296 & ~x4 & ~x29 & ~x69 & ~x72 & ~x92 & ~x103 & ~x108 & ~x120 & ~x124 & ~x128 & ~x136 & ~x140 & ~x144 & ~x155 & ~x158 & ~x161 & ~x170 & ~x184 & ~x186 & ~x192 & ~x196 & ~x249 & ~x276 & ~x305 & ~x337 & ~x344 & ~x361 & ~x391 & ~x426 & ~x448 & ~x449 & ~x471 & ~x507 & ~x525 & ~x526 & ~x552 & ~x559 & ~x579 & ~x613 & ~x636 & ~x641 & ~x643 & ~x644 & ~x663 & ~x671 & ~x689 & ~x716 & ~x723 & ~x745 & ~x749 & ~x756 & ~x767 & ~x769;
assign c7206 =  x644;
assign c7208 =  x310;
assign c7210 =  x492 & ~x1 & ~x2 & ~x5 & ~x8 & ~x11 & ~x17 & ~x18 & ~x20 & ~x22 & ~x25 & ~x27 & ~x48 & ~x56 & ~x57 & ~x68 & ~x70 & ~x73 & ~x74 & ~x77 & ~x86 & ~x90 & ~x94 & ~x102 & ~x105 & ~x107 & ~x110 & ~x114 & ~x116 & ~x117 & ~x121 & ~x127 & ~x133 & ~x134 & ~x140 & ~x141 & ~x142 & ~x190 & ~x193 & ~x194 & ~x195 & ~x219 & ~x220 & ~x223 & ~x225 & ~x247 & ~x252 & ~x253 & ~x276 & ~x282 & ~x311 & ~x321 & ~x332 & ~x337 & ~x339 & ~x360 & ~x363 & ~x368 & ~x376 & ~x377 & ~x386 & ~x387 & ~x389 & ~x396 & ~x402 & ~x423 & ~x426 & ~x429 & ~x444 & ~x445 & ~x448 & ~x452 & ~x454 & ~x455 & ~x472 & ~x478 & ~x480 & ~x500 & ~x503 & ~x504 & ~x506 & ~x509 & ~x527 & ~x528 & ~x538 & ~x558 & ~x560 & ~x581 & ~x583 & ~x587 & ~x588 & ~x589 & ~x597 & ~x598 & ~x609 & ~x614 & ~x617 & ~x618 & ~x621 & ~x622 & ~x669 & ~x676 & ~x678 & ~x680 & ~x681 & ~x700 & ~x703 & ~x705 & ~x719 & ~x720 & ~x721 & ~x726 & ~x727 & ~x728 & ~x731 & ~x733 & ~x737 & ~x739 & ~x740 & ~x749 & ~x755 & ~x762 & ~x766 & ~x771 & ~x772 & ~x774 & ~x778 & ~x781 & ~x782;
assign c7212 =  x707;
assign c7214 =  x232 &  x233 & ~x0 & ~x2 & ~x3 & ~x5 & ~x6 & ~x7 & ~x15 & ~x16 & ~x18 & ~x19 & ~x28 & ~x29 & ~x31 & ~x33 & ~x36 & ~x38 & ~x39 & ~x42 & ~x48 & ~x51 & ~x52 & ~x54 & ~x55 & ~x56 & ~x60 & ~x63 & ~x67 & ~x72 & ~x73 & ~x74 & ~x77 & ~x78 & ~x82 & ~x86 & ~x87 & ~x88 & ~x90 & ~x92 & ~x99 & ~x101 & ~x106 & ~x111 & ~x114 & ~x116 & ~x118 & ~x122 & ~x125 & ~x126 & ~x127 & ~x128 & ~x131 & ~x132 & ~x134 & ~x138 & ~x141 & ~x145 & ~x146 & ~x148 & ~x149 & ~x150 & ~x151 & ~x154 & ~x156 & ~x159 & ~x160 & ~x162 & ~x163 & ~x164 & ~x166 & ~x167 & ~x168 & ~x169 & ~x170 & ~x171 & ~x176 & ~x177 & ~x178 & ~x179 & ~x191 & ~x192 & ~x195 & ~x197 & ~x198 & ~x219 & ~x222 & ~x225 & ~x248 & ~x275 & ~x276 & ~x278 & ~x280 & ~x282 & ~x283 & ~x307 & ~x310 & ~x331 & ~x332 & ~x333 & ~x335 & ~x336 & ~x338 & ~x339 & ~x340 & ~x341 & ~x363 & ~x388 & ~x390 & ~x392 & ~x394 & ~x395 & ~x423 & ~x425 & ~x447 & ~x448 & ~x449 & ~x450 & ~x451 & ~x452 & ~x476 & ~x477 & ~x502 & ~x504 & ~x505 & ~x506 & ~x507 & ~x508 & ~x531 & ~x532 & ~x536 & ~x537 & ~x539 & ~x556 & ~x558 & ~x559 & ~x562 & ~x565 & ~x566 & ~x567 & ~x570 & ~x571 & ~x579 & ~x580 & ~x581 & ~x582 & ~x584 & ~x585 & ~x587 & ~x589 & ~x590 & ~x593 & ~x594 & ~x595 & ~x598 & ~x607 & ~x609 & ~x610 & ~x611 & ~x612 & ~x614 & ~x615 & ~x616 & ~x618 & ~x621 & ~x625 & ~x636 & ~x637 & ~x640 & ~x645 & ~x648 & ~x652 & ~x664 & ~x667 & ~x670 & ~x673 & ~x675 & ~x677 & ~x678 & ~x680 & ~x681 & ~x690 & ~x695 & ~x698 & ~x699 & ~x700 & ~x703 & ~x706 & ~x718 & ~x722 & ~x724 & ~x733 & ~x735 & ~x736 & ~x752 & ~x757 & ~x758 & ~x760 & ~x762 & ~x770 & ~x773 & ~x774 & ~x781;
assign c7216 = ~x5 & ~x13 & ~x18 & ~x44 & ~x52 & ~x54 & ~x61 & ~x67 & ~x78 & ~x81 & ~x85 & ~x93 & ~x98 & ~x107 & ~x120 & ~x129 & ~x135 & ~x137 & ~x139 & ~x148 & ~x160 & ~x163 & ~x169 & ~x181 & ~x184 & ~x207 & ~x211 & ~x220 & ~x221 & ~x225 & ~x305 & ~x308 & ~x309 & ~x363 & ~x429 & ~x488 & ~x499 & ~x507 & ~x514 & ~x533 & ~x537 & ~x543 & ~x556 & ~x569 & ~x598 & ~x612 & ~x625 & ~x627 & ~x645 & ~x649 & ~x650 & ~x651 & ~x668 & ~x679 & ~x698 & ~x701 & ~x703 & ~x723 & ~x751 & ~x763 & ~x783;
assign c7218 =  x209 &  x268 &  x572 &  x683 & ~x141 & ~x577 & ~x631 & ~x687;
assign c7220 =  x410 &  x492 & ~x13 & ~x14 & ~x42 & ~x46 & ~x59 & ~x73 & ~x77 & ~x86 & ~x108 & ~x125 & ~x129 & ~x169 & ~x191 & ~x198 & ~x199 & ~x221 & ~x229 & ~x276 & ~x310 & ~x336 & ~x337 & ~x378 & ~x391 & ~x405 & ~x443 & ~x460 & ~x472 & ~x486 & ~x505 & ~x514 & ~x515 & ~x534 & ~x541 & ~x542 & ~x561 & ~x567 & ~x568 & ~x581 & ~x584 & ~x610 & ~x611 & ~x614 & ~x621 & ~x645 & ~x646 & ~x665 & ~x672 & ~x673 & ~x675 & ~x702 & ~x725 & ~x734 & ~x743 & ~x749 & ~x750 & ~x769 & ~x770 & ~x773 & ~x774;
assign c7224 =  x464 & ~x4 & ~x10 & ~x13 & ~x14 & ~x21 & ~x27 & ~x28 & ~x33 & ~x35 & ~x37 & ~x44 & ~x45 & ~x49 & ~x50 & ~x51 & ~x52 & ~x53 & ~x55 & ~x59 & ~x61 & ~x67 & ~x68 & ~x72 & ~x76 & ~x78 & ~x84 & ~x85 & ~x87 & ~x93 & ~x94 & ~x98 & ~x101 & ~x104 & ~x105 & ~x107 & ~x109 & ~x111 & ~x116 & ~x117 & ~x119 & ~x122 & ~x126 & ~x129 & ~x132 & ~x134 & ~x135 & ~x136 & ~x141 & ~x142 & ~x145 & ~x157 & ~x158 & ~x160 & ~x161 & ~x164 & ~x194 & ~x195 & ~x218 & ~x221 & ~x223 & ~x224 & ~x225 & ~x247 & ~x252 & ~x253 & ~x281 & ~x300 & ~x302 & ~x303 & ~x304 & ~x311 & ~x313 & ~x328 & ~x330 & ~x347 & ~x348 & ~x349 & ~x361 & ~x364 & ~x375 & ~x376 & ~x392 & ~x394 & ~x396 & ~x401 & ~x417 & ~x422 & ~x424 & ~x425 & ~x443 & ~x444 & ~x447 & ~x452 & ~x471 & ~x476 & ~x477 & ~x481 & ~x499 & ~x502 & ~x508 & ~x527 & ~x533 & ~x536 & ~x555 & ~x564 & ~x565 & ~x566 & ~x587 & ~x606 & ~x609 & ~x634 & ~x640 & ~x641 & ~x649 & ~x663 & ~x670 & ~x671 & ~x678 & ~x680 & ~x690 & ~x693 & ~x695 & ~x701 & ~x702 & ~x708 & ~x710 & ~x718 & ~x726 & ~x727 & ~x730 & ~x735 & ~x747 & ~x755 & ~x758 & ~x761 & ~x762 & ~x763 & ~x765 & ~x766 & ~x767 & ~x770 & ~x773 & ~x780;
assign c7226 =  x235 & ~x3 & ~x10 & ~x12 & ~x13 & ~x15 & ~x33 & ~x43 & ~x44 & ~x48 & ~x58 & ~x75 & ~x93 & ~x105 & ~x125 & ~x134 & ~x136 & ~x143 & ~x160 & ~x166 & ~x169 & ~x192 & ~x196 & ~x197 & ~x220 & ~x228 & ~x248 & ~x254 & ~x284 & ~x307 & ~x318 & ~x319 & ~x321 & ~x332 & ~x342 & ~x343 & ~x363 & ~x366 & ~x369 & ~x370 & ~x372 & ~x392 & ~x446 & ~x447 & ~x473 & ~x504 & ~x508 & ~x530 & ~x534 & ~x559 & ~x581 & ~x586 & ~x594 & ~x606 & ~x612 & ~x613 & ~x616 & ~x621 & ~x632 & ~x635 & ~x642 & ~x664 & ~x674 & ~x675 & ~x689 & ~x694 & ~x703 & ~x721 & ~x722 & ~x729 & ~x730 & ~x735 & ~x736 & ~x741 & ~x747 & ~x755 & ~x780;
assign c7228 =  x316 &  x317 &  x318 & ~x19 & ~x180 & ~x183 & ~x205 & ~x209 & ~x212 & ~x499 & ~x540 & ~x555 & ~x595;
assign c7230 =  x264 &  x294 &  x295 & ~x5 & ~x6 & ~x12 & ~x16 & ~x19 & ~x22 & ~x23 & ~x24 & ~x26 & ~x27 & ~x30 & ~x31 & ~x36 & ~x37 & ~x38 & ~x43 & ~x46 & ~x49 & ~x50 & ~x52 & ~x54 & ~x59 & ~x62 & ~x67 & ~x70 & ~x72 & ~x73 & ~x76 & ~x77 & ~x82 & ~x86 & ~x88 & ~x90 & ~x91 & ~x98 & ~x101 & ~x107 & ~x108 & ~x109 & ~x113 & ~x115 & ~x119 & ~x120 & ~x122 & ~x124 & ~x126 & ~x131 & ~x136 & ~x137 & ~x142 & ~x143 & ~x145 & ~x146 & ~x149 & ~x165 & ~x167 & ~x169 & ~x170 & ~x172 & ~x188 & ~x190 & ~x195 & ~x196 & ~x219 & ~x220 & ~x224 & ~x226 & ~x227 & ~x250 & ~x255 & ~x275 & ~x278 & ~x279 & ~x282 & ~x305 & ~x310 & ~x332 & ~x333 & ~x341 & ~x368 & ~x388 & ~x390 & ~x391 & ~x446 & ~x447 & ~x449 & ~x450 & ~x474 & ~x475 & ~x477 & ~x478 & ~x479 & ~x501 & ~x504 & ~x506 & ~x515 & ~x529 & ~x530 & ~x540 & ~x541 & ~x542 & ~x563 & ~x564 & ~x565 & ~x569 & ~x570 & ~x583 & ~x589 & ~x591 & ~x592 & ~x593 & ~x595 & ~x596 & ~x597 & ~x598 & ~x599 & ~x608 & ~x613 & ~x614 & ~x622 & ~x625 & ~x636 & ~x639 & ~x641 & ~x642 & ~x645 & ~x646 & ~x648 & ~x650 & ~x652 & ~x653 & ~x654 & ~x673 & ~x677 & ~x692 & ~x695 & ~x696 & ~x698 & ~x720 & ~x723 & ~x724 & ~x725 & ~x727 & ~x728 & ~x733 & ~x735 & ~x736 & ~x739 & ~x740 & ~x745 & ~x751 & ~x753 & ~x754 & ~x761 & ~x763 & ~x764 & ~x765 & ~x768 & ~x771 & ~x781;
assign c7232 =  x233 &  x266 &  x631 &  x715 & ~x663;
assign c7234 = ~x0 & ~x4 & ~x5 & ~x9 & ~x11 & ~x12 & ~x14 & ~x15 & ~x17 & ~x18 & ~x19 & ~x21 & ~x22 & ~x28 & ~x36 & ~x37 & ~x40 & ~x41 & ~x43 & ~x47 & ~x52 & ~x54 & ~x57 & ~x59 & ~x61 & ~x66 & ~x68 & ~x70 & ~x72 & ~x74 & ~x78 & ~x89 & ~x91 & ~x92 & ~x95 & ~x97 & ~x98 & ~x100 & ~x102 & ~x103 & ~x108 & ~x109 & ~x110 & ~x112 & ~x117 & ~x118 & ~x120 & ~x124 & ~x128 & ~x131 & ~x133 & ~x136 & ~x140 & ~x153 & ~x156 & ~x158 & ~x165 & ~x169 & ~x171 & ~x194 & ~x196 & ~x200 & ~x201 & ~x219 & ~x226 & ~x227 & ~x253 & ~x276 & ~x277 & ~x279 & ~x281 & ~x303 & ~x304 & ~x310 & ~x311 & ~x330 & ~x339 & ~x349 & ~x359 & ~x362 & ~x363 & ~x366 & ~x377 & ~x385 & ~x388 & ~x389 & ~x405 & ~x413 & ~x414 & ~x417 & ~x432 & ~x433 & ~x443 & ~x444 & ~x446 & ~x447 & ~x450 & ~x460 & ~x473 & ~x474 & ~x479 & ~x497 & ~x500 & ~x504 & ~x509 & ~x515 & ~x526 & ~x531 & ~x537 & ~x559 & ~x561 & ~x563 & ~x581 & ~x584 & ~x588 & ~x590 & ~x592 & ~x614 & ~x615 & ~x619 & ~x637 & ~x650 & ~x666 & ~x669 & ~x671 & ~x675 & ~x677 & ~x680 & ~x692 & ~x695 & ~x696 & ~x701 & ~x705 & ~x706 & ~x720 & ~x721 & ~x726 & ~x735 & ~x737 & ~x738 & ~x741 & ~x748 & ~x750 & ~x752 & ~x764 & ~x772 & ~x774 & ~x775 & ~x776;
assign c7236 = ~x10 & ~x16 & ~x33 & ~x35 & ~x43 & ~x55 & ~x59 & ~x67 & ~x78 & ~x84 & ~x95 & ~x97 & ~x101 & ~x105 & ~x124 & ~x131 & ~x138 & ~x143 & ~x153 & ~x155 & ~x166 & ~x167 & ~x195 & ~x196 & ~x249 & ~x255 & ~x257 & ~x275 & ~x276 & ~x278 & ~x284 & ~x322 & ~x360 & ~x376 & ~x377 & ~x385 & ~x386 & ~x405 & ~x420 & ~x432 & ~x444 & ~x445 & ~x459 & ~x470 & ~x499 & ~x502 & ~x515 & ~x556 & ~x586 & ~x617 & ~x624 & ~x641 & ~x670 & ~x702 & ~x705 & ~x723 & ~x733 & ~x755 & ~x761 & ~x779;
assign c7238 =  x267 &  x294 &  x295 &  x323 &  x437 &  x438 & ~x4 & ~x14 & ~x18 & ~x22 & ~x25 & ~x26 & ~x31 & ~x33 & ~x57 & ~x68 & ~x82 & ~x83 & ~x100 & ~x112 & ~x127 & ~x136 & ~x140 & ~x151 & ~x153 & ~x166 & ~x186 & ~x250 & ~x282 & ~x334 & ~x335 & ~x336 & ~x360 & ~x390 & ~x450 & ~x478 & ~x502 & ~x529 & ~x531 & ~x536 & ~x540 & ~x541 & ~x554 & ~x563 & ~x566 & ~x580 & ~x583 & ~x588 & ~x597 & ~x624 & ~x648 & ~x649 & ~x665 & ~x667 & ~x668 & ~x693 & ~x702 & ~x731 & ~x733 & ~x736 & ~x743 & ~x744 & ~x745 & ~x749 & ~x762 & ~x763 & ~x768 & ~x771 & ~x776;
assign c7240 =  x262 &  x264 &  x265 &  x266 & ~x7 & ~x21 & ~x27 & ~x37 & ~x41 & ~x56 & ~x73 & ~x78 & ~x81 & ~x85 & ~x90 & ~x92 & ~x93 & ~x98 & ~x101 & ~x110 & ~x111 & ~x115 & ~x118 & ~x122 & ~x128 & ~x134 & ~x142 & ~x144 & ~x147 & ~x156 & ~x161 & ~x190 & ~x191 & ~x193 & ~x195 & ~x220 & ~x224 & ~x249 & ~x276 & ~x305 & ~x308 & ~x359 & ~x365 & ~x376 & ~x388 & ~x393 & ~x403 & ~x404 & ~x421 & ~x431 & ~x477 & ~x478 & ~x501 & ~x502 & ~x506 & ~x508 & ~x528 & ~x544 & ~x555 & ~x570 & ~x571 & ~x572 & ~x582 & ~x591 & ~x596 & ~x597 & ~x612 & ~x615 & ~x621 & ~x637 & ~x638 & ~x640 & ~x650 & ~x666 & ~x671 & ~x673 & ~x674 & ~x679 & ~x681 & ~x694 & ~x695 & ~x702 & ~x706 & ~x727 & ~x735 & ~x736 & ~x740 & ~x753 & ~x759 & ~x763 & ~x767 & ~x781;
assign c7242 =  x496 &  x689;
assign c7244 =  x478;
assign c7246 =  x460 &  x463 &  x464 & ~x0 & ~x11 & ~x14 & ~x21 & ~x24 & ~x26 & ~x28 & ~x29 & ~x30 & ~x48 & ~x60 & ~x84 & ~x93 & ~x95 & ~x98 & ~x113 & ~x120 & ~x132 & ~x190 & ~x193 & ~x196 & ~x220 & ~x255 & ~x257 & ~x274 & ~x276 & ~x281 & ~x303 & ~x304 & ~x311 & ~x316 & ~x335 & ~x339 & ~x341 & ~x345 & ~x347 & ~x349 & ~x365 & ~x399 & ~x420 & ~x425 & ~x448 & ~x472 & ~x476 & ~x505 & ~x506 & ~x508 & ~x509 & ~x556 & ~x564 & ~x567 & ~x569 & ~x587 & ~x590 & ~x596 & ~x619 & ~x620 & ~x625 & ~x637 & ~x651 & ~x665 & ~x668 & ~x680 & ~x693 & ~x697 & ~x721 & ~x725 & ~x749 & ~x752 & ~x766 & ~x767;
assign c7248 =  x208 &  x296 &  x461 &  x462 & ~x2 & ~x5 & ~x6 & ~x11 & ~x13 & ~x14 & ~x18 & ~x32 & ~x34 & ~x57 & ~x60 & ~x64 & ~x75 & ~x78 & ~x81 & ~x87 & ~x93 & ~x101 & ~x110 & ~x114 & ~x121 & ~x123 & ~x125 & ~x126 & ~x132 & ~x135 & ~x169 & ~x172 & ~x191 & ~x254 & ~x299 & ~x303 & ~x315 & ~x326 & ~x334 & ~x338 & ~x341 & ~x347 & ~x348 & ~x360 & ~x366 & ~x368 & ~x422 & ~x504 & ~x529 & ~x536 & ~x539 & ~x540 & ~x561 & ~x566 & ~x591 & ~x594 & ~x638 & ~x642 & ~x649 & ~x668 & ~x691 & ~x694 & ~x698 & ~x704 & ~x749 & ~x752 & ~x764 & ~x769 & ~x770 & ~x771 & ~x777 & ~x778;
assign c7250 =  x256 &  x285;
assign c7252 =  x209 &  x239 &  x241 &  x324 &  x489 &  x516 & ~x224 & ~x450 & ~x520 & ~x576 & ~x603 & ~x606 & ~x659 & ~x770;
assign c7254 =  x337;
assign c7256 =  x77;
assign c7258 = ~x1 & ~x3 & ~x4 & ~x7 & ~x15 & ~x19 & ~x25 & ~x28 & ~x33 & ~x37 & ~x39 & ~x41 & ~x45 & ~x47 & ~x49 & ~x50 & ~x66 & ~x68 & ~x75 & ~x78 & ~x82 & ~x83 & ~x88 & ~x89 & ~x98 & ~x101 & ~x104 & ~x109 & ~x111 & ~x118 & ~x121 & ~x126 & ~x127 & ~x134 & ~x144 & ~x146 & ~x154 & ~x156 & ~x160 & ~x166 & ~x169 & ~x173 & ~x182 & ~x183 & ~x185 & ~x187 & ~x195 & ~x198 & ~x204 & ~x223 & ~x225 & ~x226 & ~x229 & ~x253 & ~x278 & ~x281 & ~x305 & ~x334 & ~x336 & ~x337 & ~x364 & ~x365 & ~x379 & ~x389 & ~x405 & ~x406 & ~x418 & ~x423 & ~x479 & ~x486 & ~x500 & ~x501 & ~x504 & ~x505 & ~x507 & ~x513 & ~x535 & ~x541 & ~x542 & ~x555 & ~x569 & ~x587 & ~x588 & ~x589 & ~x592 & ~x597 & ~x613 & ~x614 & ~x617 & ~x618 & ~x639 & ~x696 & ~x697 & ~x698 & ~x723 & ~x725 & ~x729 & ~x732 & ~x733 & ~x755 & ~x757 & ~x758 & ~x759 & ~x760 & ~x767 & ~x769 & ~x773 & ~x778 & ~x779 & ~x780 & ~x781 & ~x782;
assign c7260 =  x319 & ~x149 & ~x180 & ~x181 & ~x216 & ~x432 & ~x569 & ~x571 & ~x624;
assign c7262 =  x236 &  x239 &  x264 &  x352 & ~x2 & ~x3 & ~x4 & ~x7 & ~x9 & ~x12 & ~x30 & ~x51 & ~x55 & ~x56 & ~x59 & ~x71 & ~x72 & ~x80 & ~x88 & ~x89 & ~x98 & ~x100 & ~x107 & ~x121 & ~x129 & ~x130 & ~x138 & ~x151 & ~x154 & ~x155 & ~x158 & ~x160 & ~x163 & ~x167 & ~x195 & ~x220 & ~x276 & ~x277 & ~x281 & ~x282 & ~x284 & ~x304 & ~x310 & ~x312 & ~x313 & ~x328 & ~x333 & ~x337 & ~x359 & ~x364 & ~x367 & ~x374 & ~x393 & ~x418 & ~x422 & ~x447 & ~x475 & ~x480 & ~x501 & ~x503 & ~x504 & ~x507 & ~x530 & ~x536 & ~x537 & ~x565 & ~x583 & ~x596 & ~x613 & ~x614 & ~x616 & ~x618 & ~x645 & ~x668 & ~x724 & ~x725 & ~x731 & ~x737 & ~x745 & ~x750 & ~x751 & ~x755 & ~x771 & ~x777 & ~x778;
assign c7264 =  x319 &  x322 &  x411 & ~x3 & ~x8 & ~x12 & ~x17 & ~x21 & ~x23 & ~x26 & ~x35 & ~x36 & ~x39 & ~x40 & ~x43 & ~x44 & ~x45 & ~x46 & ~x49 & ~x50 & ~x57 & ~x66 & ~x67 & ~x70 & ~x74 & ~x79 & ~x80 & ~x88 & ~x91 & ~x105 & ~x108 & ~x109 & ~x111 & ~x122 & ~x127 & ~x131 & ~x134 & ~x136 & ~x138 & ~x139 & ~x140 & ~x141 & ~x142 & ~x149 & ~x151 & ~x153 & ~x154 & ~x156 & ~x159 & ~x160 & ~x163 & ~x167 & ~x183 & ~x184 & ~x190 & ~x191 & ~x194 & ~x195 & ~x213 & ~x249 & ~x252 & ~x277 & ~x278 & ~x279 & ~x280 & ~x306 & ~x361 & ~x363 & ~x365 & ~x391 & ~x418 & ~x445 & ~x475 & ~x478 & ~x502 & ~x503 & ~x506 & ~x527 & ~x528 & ~x533 & ~x538 & ~x556 & ~x591 & ~x595 & ~x615 & ~x622 & ~x639 & ~x642 & ~x670 & ~x672 & ~x679 & ~x701 & ~x724 & ~x728 & ~x731 & ~x743 & ~x751 & ~x752 & ~x753 & ~x759 & ~x761 & ~x764 & ~x768 & ~x771 & ~x777 & ~x779 & ~x780 & ~x783;
assign c7266 = ~x3 & ~x4 & ~x6 & ~x8 & ~x9 & ~x11 & ~x13 & ~x15 & ~x20 & ~x25 & ~x28 & ~x31 & ~x32 & ~x36 & ~x38 & ~x43 & ~x44 & ~x48 & ~x49 & ~x51 & ~x55 & ~x56 & ~x57 & ~x59 & ~x60 & ~x66 & ~x75 & ~x79 & ~x81 & ~x82 & ~x84 & ~x88 & ~x89 & ~x90 & ~x92 & ~x95 & ~x96 & ~x99 & ~x104 & ~x106 & ~x109 & ~x110 & ~x111 & ~x112 & ~x116 & ~x117 & ~x118 & ~x119 & ~x121 & ~x125 & ~x127 & ~x135 & ~x139 & ~x140 & ~x142 & ~x143 & ~x149 & ~x153 & ~x154 & ~x157 & ~x160 & ~x162 & ~x163 & ~x165 & ~x166 & ~x168 & ~x169 & ~x170 & ~x171 & ~x192 & ~x193 & ~x196 & ~x221 & ~x247 & ~x248 & ~x250 & ~x254 & ~x280 & ~x281 & ~x282 & ~x283 & ~x306 & ~x307 & ~x334 & ~x335 & ~x337 & ~x338 & ~x339 & ~x350 & ~x359 & ~x364 & ~x366 & ~x378 & ~x389 & ~x393 & ~x395 & ~x405 & ~x406 & ~x416 & ~x433 & ~x434 & ~x445 & ~x457 & ~x460 & ~x472 & ~x473 & ~x474 & ~x475 & ~x477 & ~x479 & ~x480 & ~x481 & ~x486 & ~x488 & ~x500 & ~x501 & ~x506 & ~x508 & ~x510 & ~x513 & ~x527 & ~x530 & ~x531 & ~x535 & ~x537 & ~x555 & ~x558 & ~x560 & ~x562 & ~x564 & ~x566 & ~x584 & ~x590 & ~x612 & ~x617 & ~x618 & ~x620 & ~x621 & ~x623 & ~x638 & ~x642 & ~x643 & ~x646 & ~x647 & ~x650 & ~x667 & ~x671 & ~x696 & ~x697 & ~x698 & ~x703 & ~x706 & ~x722 & ~x725 & ~x727 & ~x728 & ~x734 & ~x735 & ~x736 & ~x752 & ~x755 & ~x756 & ~x757 & ~x760 & ~x762 & ~x765 & ~x766 & ~x767 & ~x770 & ~x771 & ~x772 & ~x778 & ~x780;
assign c7268 =  x765;
assign c7270 =  x231;
assign c7272 =  x206 &  x519 & ~x3 & ~x23 & ~x24 & ~x25 & ~x28 & ~x42 & ~x48 & ~x49 & ~x51 & ~x55 & ~x61 & ~x65 & ~x71 & ~x75 & ~x76 & ~x78 & ~x83 & ~x84 & ~x86 & ~x100 & ~x102 & ~x111 & ~x113 & ~x114 & ~x123 & ~x126 & ~x127 & ~x134 & ~x136 & ~x141 & ~x143 & ~x158 & ~x161 & ~x165 & ~x168 & ~x171 & ~x194 & ~x198 & ~x199 & ~x221 & ~x222 & ~x224 & ~x225 & ~x248 & ~x252 & ~x254 & ~x256 & ~x278 & ~x281 & ~x283 & ~x304 & ~x306 & ~x309 & ~x313 & ~x314 & ~x332 & ~x333 & ~x334 & ~x337 & ~x339 & ~x348 & ~x357 & ~x361 & ~x362 & ~x367 & ~x394 & ~x396 & ~x397 & ~x416 & ~x422 & ~x423 & ~x425 & ~x451 & ~x475 & ~x478 & ~x480 & ~x481 & ~x509 & ~x525 & ~x533 & ~x535 & ~x556 & ~x559 & ~x561 & ~x569 & ~x586 & ~x591 & ~x606 & ~x608 & ~x609 & ~x613 & ~x622 & ~x623 & ~x635 & ~x636 & ~x638 & ~x640 & ~x642 & ~x645 & ~x646 & ~x650 & ~x651 & ~x663 & ~x664 & ~x666 & ~x670 & ~x696 & ~x702 & ~x705 & ~x707 & ~x711 & ~x718 & ~x720 & ~x724 & ~x727 & ~x737 & ~x746 & ~x750 & ~x753 & ~x759 & ~x771 & ~x773 & ~x778 & ~x779 & ~x780 & ~x783;
assign c7274 = ~x2 & ~x7 & ~x8 & ~x18 & ~x21 & ~x22 & ~x23 & ~x24 & ~x29 & ~x31 & ~x43 & ~x44 & ~x45 & ~x49 & ~x53 & ~x55 & ~x57 & ~x63 & ~x64 & ~x67 & ~x68 & ~x69 & ~x71 & ~x72 & ~x75 & ~x81 & ~x83 & ~x86 & ~x90 & ~x91 & ~x93 & ~x94 & ~x96 & ~x99 & ~x101 & ~x105 & ~x106 & ~x111 & ~x112 & ~x113 & ~x118 & ~x119 & ~x120 & ~x124 & ~x127 & ~x131 & ~x137 & ~x143 & ~x147 & ~x148 & ~x149 & ~x150 & ~x153 & ~x155 & ~x156 & ~x159 & ~x160 & ~x162 & ~x170 & ~x176 & ~x177 & ~x178 & ~x179 & ~x182 & ~x183 & ~x189 & ~x191 & ~x196 & ~x198 & ~x209 & ~x223 & ~x224 & ~x226 & ~x250 & ~x251 & ~x277 & ~x304 & ~x306 & ~x333 & ~x334 & ~x391 & ~x417 & ~x431 & ~x445 & ~x449 & ~x474 & ~x476 & ~x486 & ~x487 & ~x502 & ~x515 & ~x530 & ~x531 & ~x532 & ~x533 & ~x534 & ~x541 & ~x543 & ~x554 & ~x555 & ~x567 & ~x569 & ~x570 & ~x571 & ~x572 & ~x582 & ~x589 & ~x590 & ~x591 & ~x596 & ~x597 & ~x598 & ~x599 & ~x611 & ~x614 & ~x616 & ~x620 & ~x624 & ~x625 & ~x626 & ~x627 & ~x638 & ~x639 & ~x642 & ~x646 & ~x653 & ~x654 & ~x655 & ~x666 & ~x668 & ~x674 & ~x677 & ~x679 & ~x680 & ~x701 & ~x705 & ~x708 & ~x710 & ~x724 & ~x725 & ~x727 & ~x729 & ~x730 & ~x731 & ~x732 & ~x734 & ~x736 & ~x738 & ~x754 & ~x762 & ~x764 & ~x781 & ~x782;
assign c7276 =  x261 &  x263 &  x266 & ~x0 & ~x4 & ~x12 & ~x18 & ~x22 & ~x26 & ~x29 & ~x38 & ~x39 & ~x40 & ~x49 & ~x60 & ~x64 & ~x74 & ~x79 & ~x86 & ~x99 & ~x109 & ~x125 & ~x126 & ~x128 & ~x138 & ~x143 & ~x151 & ~x152 & ~x158 & ~x165 & ~x196 & ~x248 & ~x280 & ~x283 & ~x306 & ~x307 & ~x311 & ~x334 & ~x388 & ~x395 & ~x404 & ~x432 & ~x433 & ~x446 & ~x500 & ~x506 & ~x507 & ~x528 & ~x544 & ~x556 & ~x557 & ~x566 & ~x572 & ~x582 & ~x583 & ~x585 & ~x614 & ~x639 & ~x642 & ~x652 & ~x671 & ~x672 & ~x697 & ~x698 & ~x706 & ~x707 & ~x723 & ~x725 & ~x729 & ~x730 & ~x739 & ~x755 & ~x761 & ~x762 & ~x763 & ~x766 & ~x775 & ~x780 & ~x783;
assign c7278 =  x701;
assign c7280 =  x516 &  x678 & ~x404;
assign c7282 = ~x1 & ~x3 & ~x7 & ~x13 & ~x14 & ~x33 & ~x34 & ~x44 & ~x45 & ~x47 & ~x51 & ~x53 & ~x63 & ~x95 & ~x96 & ~x108 & ~x112 & ~x113 & ~x123 & ~x127 & ~x131 & ~x132 & ~x133 & ~x136 & ~x140 & ~x143 & ~x146 & ~x147 & ~x151 & ~x153 & ~x155 & ~x158 & ~x164 & ~x167 & ~x174 & ~x177 & ~x179 & ~x180 & ~x185 & ~x187 & ~x188 & ~x191 & ~x197 & ~x214 & ~x223 & ~x333 & ~x363 & ~x388 & ~x391 & ~x433 & ~x435 & ~x446 & ~x460 & ~x461 & ~x472 & ~x473 & ~x479 & ~x502 & ~x507 & ~x515 & ~x535 & ~x539 & ~x567 & ~x568 & ~x585 & ~x588 & ~x591 & ~x595 & ~x610 & ~x614 & ~x640 & ~x642 & ~x647 & ~x651 & ~x698 & ~x745 & ~x751 & ~x768 & ~x771 & ~x783;
assign c7284 =  x236 &  x435 & ~x2 & ~x3 & ~x4 & ~x7 & ~x9 & ~x10 & ~x13 & ~x17 & ~x21 & ~x22 & ~x24 & ~x26 & ~x27 & ~x30 & ~x31 & ~x44 & ~x45 & ~x58 & ~x61 & ~x66 & ~x67 & ~x77 & ~x83 & ~x89 & ~x105 & ~x110 & ~x115 & ~x119 & ~x123 & ~x128 & ~x132 & ~x136 & ~x137 & ~x140 & ~x150 & ~x159 & ~x167 & ~x169 & ~x171 & ~x172 & ~x190 & ~x199 & ~x220 & ~x221 & ~x223 & ~x227 & ~x249 & ~x254 & ~x277 & ~x278 & ~x280 & ~x281 & ~x282 & ~x307 & ~x314 & ~x320 & ~x336 & ~x340 & ~x345 & ~x349 & ~x358 & ~x366 & ~x370 & ~x371 & ~x394 & ~x426 & ~x444 & ~x445 & ~x451 & ~x501 & ~x503 & ~x509 & ~x527 & ~x528 & ~x533 & ~x557 & ~x565 & ~x577 & ~x581 & ~x584 & ~x587 & ~x594 & ~x608 & ~x611 & ~x616 & ~x618 & ~x619 & ~x620 & ~x621 & ~x633 & ~x634 & ~x645 & ~x646 & ~x661 & ~x662 & ~x666 & ~x667 & ~x669 & ~x671 & ~x678 & ~x688 & ~x699 & ~x706 & ~x707 & ~x717 & ~x723 & ~x726 & ~x734 & ~x744 & ~x764 & ~x769 & ~x770 & ~x773 & ~x781;
assign c7286 =  x239 &  x241 & ~x1 & ~x2 & ~x11 & ~x20 & ~x22 & ~x26 & ~x47 & ~x49 & ~x50 & ~x51 & ~x53 & ~x55 & ~x59 & ~x68 & ~x78 & ~x79 & ~x81 & ~x86 & ~x90 & ~x91 & ~x92 & ~x94 & ~x102 & ~x106 & ~x110 & ~x113 & ~x125 & ~x128 & ~x130 & ~x131 & ~x141 & ~x142 & ~x145 & ~x146 & ~x167 & ~x172 & ~x194 & ~x196 & ~x199 & ~x223 & ~x227 & ~x229 & ~x250 & ~x251 & ~x252 & ~x283 & ~x284 & ~x308 & ~x313 & ~x322 & ~x331 & ~x333 & ~x335 & ~x339 & ~x340 & ~x342 & ~x350 & ~x358 & ~x359 & ~x364 & ~x367 & ~x385 & ~x386 & ~x394 & ~x396 & ~x423 & ~x448 & ~x450 & ~x498 & ~x499 & ~x501 & ~x502 & ~x506 & ~x508 & ~x529 & ~x534 & ~x556 & ~x585 & ~x592 & ~x593 & ~x609 & ~x610 & ~x615 & ~x632 & ~x639 & ~x640 & ~x647 & ~x666 & ~x668 & ~x673 & ~x676 & ~x688 & ~x692 & ~x695 & ~x697 & ~x699 & ~x700 & ~x701 & ~x702 & ~x720 & ~x723 & ~x731 & ~x734 & ~x740 & ~x742 & ~x743 & ~x745 & ~x751 & ~x763 & ~x772 & ~x776 & ~x777 & ~x780 & ~x783;
assign c7288 =  x6;
assign c7290 = ~x5 & ~x7 & ~x19 & ~x21 & ~x25 & ~x26 & ~x33 & ~x43 & ~x44 & ~x47 & ~x50 & ~x54 & ~x71 & ~x73 & ~x78 & ~x79 & ~x81 & ~x83 & ~x86 & ~x87 & ~x95 & ~x99 & ~x101 & ~x103 & ~x104 & ~x108 & ~x110 & ~x111 & ~x116 & ~x119 & ~x120 & ~x121 & ~x123 & ~x124 & ~x126 & ~x127 & ~x129 & ~x137 & ~x138 & ~x141 & ~x161 & ~x165 & ~x173 & ~x175 & ~x176 & ~x177 & ~x190 & ~x219 & ~x220 & ~x225 & ~x251 & ~x253 & ~x255 & ~x278 & ~x280 & ~x284 & ~x309 & ~x313 & ~x338 & ~x339 & ~x349 & ~x350 & ~x365 & ~x367 & ~x376 & ~x395 & ~x404 & ~x422 & ~x447 & ~x448 & ~x450 & ~x453 & ~x456 & ~x473 & ~x481 & ~x498 & ~x503 & ~x505 & ~x507 & ~x527 & ~x535 & ~x537 & ~x553 & ~x556 & ~x559 & ~x565 & ~x587 & ~x590 & ~x614 & ~x615 & ~x663 & ~x671 & ~x675 & ~x692 & ~x693 & ~x728 & ~x733 & ~x738 & ~x741 & ~x747 & ~x750 & ~x755 & ~x758 & ~x765 & ~x777 & ~x780 & ~x783;
assign c7294 =  x214 &  x298 &  x462 &  x463 &  x490 &  x544 & ~x19 & ~x50 & ~x57 & ~x63 & ~x101 & ~x121 & ~x192 & ~x311 & ~x350 & ~x377 & ~x393 & ~x395 & ~x454 & ~x482 & ~x535 & ~x561 & ~x605 & ~x608 & ~x635 & ~x661 & ~x692 & ~x702 & ~x716 & ~x740 & ~x775;
assign c7296 =  x206 & ~x2 & ~x3 & ~x6 & ~x7 & ~x9 & ~x12 & ~x13 & ~x14 & ~x15 & ~x16 & ~x17 & ~x19 & ~x20 & ~x21 & ~x22 & ~x23 & ~x24 & ~x29 & ~x32 & ~x34 & ~x35 & ~x37 & ~x39 & ~x49 & ~x50 & ~x52 & ~x53 & ~x57 & ~x59 & ~x62 & ~x63 & ~x64 & ~x65 & ~x69 & ~x72 & ~x75 & ~x76 & ~x77 & ~x79 & ~x80 & ~x81 & ~x82 & ~x85 & ~x86 & ~x92 & ~x97 & ~x100 & ~x101 & ~x102 & ~x104 & ~x105 & ~x110 & ~x112 & ~x115 & ~x116 & ~x117 & ~x119 & ~x120 & ~x122 & ~x123 & ~x125 & ~x127 & ~x129 & ~x131 & ~x133 & ~x138 & ~x139 & ~x140 & ~x144 & ~x145 & ~x146 & ~x160 & ~x165 & ~x167 & ~x192 & ~x194 & ~x196 & ~x197 & ~x198 & ~x220 & ~x221 & ~x226 & ~x250 & ~x252 & ~x253 & ~x257 & ~x258 & ~x275 & ~x277 & ~x278 & ~x287 & ~x288 & ~x289 & ~x291 & ~x303 & ~x304 & ~x305 & ~x306 & ~x317 & ~x332 & ~x333 & ~x334 & ~x335 & ~x337 & ~x339 & ~x344 & ~x370 & ~x391 & ~x396 & ~x416 & ~x417 & ~x418 & ~x424 & ~x425 & ~x447 & ~x451 & ~x452 & ~x470 & ~x473 & ~x476 & ~x478 & ~x480 & ~x481 & ~x499 & ~x501 & ~x505 & ~x524 & ~x525 & ~x527 & ~x528 & ~x534 & ~x538 & ~x539 & ~x549 & ~x551 & ~x554 & ~x557 & ~x558 & ~x562 & ~x577 & ~x578 & ~x580 & ~x581 & ~x587 & ~x591 & ~x604 & ~x607 & ~x608 & ~x609 & ~x610 & ~x614 & ~x616 & ~x619 & ~x620 & ~x622 & ~x632 & ~x635 & ~x638 & ~x641 & ~x642 & ~x644 & ~x645 & ~x660 & ~x663 & ~x666 & ~x669 & ~x671 & ~x673 & ~x674 & ~x675 & ~x688 & ~x689 & ~x695 & ~x696 & ~x697 & ~x698 & ~x699 & ~x700 & ~x702 & ~x703 & ~x705 & ~x706 & ~x717 & ~x718 & ~x720 & ~x721 & ~x724 & ~x734 & ~x735 & ~x743 & ~x744 & ~x746 & ~x749 & ~x750 & ~x751 & ~x758 & ~x759 & ~x760 & ~x762 & ~x766 & ~x768 & ~x770 & ~x779 & ~x781 & ~x783;
assign c7298 =  x210 &  x571 &  x653 & ~x127 & ~x577 & ~x658 & ~x675;
assign c71 =  x211 &  x578 & ~x547;
assign c73 =  x604 &  x627 &  x628 & ~x4 & ~x14 & ~x18 & ~x23 & ~x27 & ~x33 & ~x45 & ~x85 & ~x115 & ~x140 & ~x142 & ~x171 & ~x252 & ~x387 & ~x444 & ~x446 & ~x503 & ~x505 & ~x534 & ~x557 & ~x563 & ~x616 & ~x640 & ~x642 & ~x672 & ~x700 & ~x710 & ~x729 & ~x731 & ~x748 & ~x776 & ~x778;
assign c75 =  x549 & ~x0 & ~x4 & ~x9 & ~x11 & ~x12 & ~x17 & ~x29 & ~x31 & ~x33 & ~x34 & ~x37 & ~x46 & ~x48 & ~x54 & ~x55 & ~x57 & ~x59 & ~x74 & ~x79 & ~x80 & ~x91 & ~x107 & ~x134 & ~x143 & ~x144 & ~x147 & ~x165 & ~x169 & ~x173 & ~x174 & ~x193 & ~x195 & ~x199 & ~x224 & ~x229 & ~x250 & ~x255 & ~x256 & ~x281 & ~x306 & ~x308 & ~x312 & ~x336 & ~x339 & ~x365 & ~x366 & ~x367 & ~x368 & ~x389 & ~x390 & ~x394 & ~x419 & ~x446 & ~x448 & ~x449 & ~x473 & ~x475 & ~x476 & ~x477 & ~x478 & ~x503 & ~x533 & ~x534 & ~x562 & ~x581 & ~x587 & ~x589 & ~x590 & ~x591 & ~x612 & ~x615 & ~x618 & ~x619 & ~x639 & ~x640 & ~x642 & ~x648 & ~x666 & ~x667 & ~x668 & ~x673 & ~x674 & ~x675 & ~x686 & ~x687 & ~x688 & ~x689 & ~x694 & ~x696 & ~x699 & ~x700 & ~x703 & ~x704 & ~x715 & ~x716 & ~x719 & ~x725 & ~x727 & ~x736 & ~x737 & ~x738 & ~x741 & ~x746 & ~x753 & ~x754 & ~x755 & ~x756 & ~x758 & ~x766 & ~x770 & ~x774 & ~x776 & ~x777;
assign c77 =  x160;
assign c79 =  x429 & ~x87 & ~x210 & ~x237 & ~x264 & ~x480 & ~x587 & ~x617 & ~x742 & ~x781;
assign c711 =  x565;
assign c713 =  x484 & ~x6 & ~x19 & ~x55 & ~x97 & ~x144 & ~x198 & ~x203 & ~x222 & ~x228 & ~x233 & ~x253 & ~x308 & ~x313 & ~x649 & ~x650 & ~x710 & ~x713 & ~x714 & ~x719 & ~x766 & ~x769 & ~x777;
assign c715 =  x527;
assign c717 =  x346 &  x374 &  x405 & ~x13 & ~x47 & ~x82 & ~x134 & ~x170 & ~x195 & ~x196 & ~x222 & ~x226 & ~x228 & ~x282 & ~x340 & ~x396 & ~x416 & ~x473 & ~x482 & ~x497 & ~x498 & ~x561 & ~x704 & ~x763;
assign c719 =  x582;
assign c721 =  x596 & ~x17 & ~x54 & ~x63 & ~x85 & ~x91 & ~x113 & ~x137 & ~x139 & ~x202 & ~x227 & ~x309 & ~x361 & ~x528 & ~x638 & ~x667 & ~x677 & ~x679 & ~x750 & ~x762;
assign c723 =  x597 &  x598 & ~x9 & ~x23 & ~x45 & ~x47 & ~x50 & ~x52 & ~x69 & ~x78 & ~x81 & ~x137 & ~x138 & ~x160 & ~x277 & ~x283 & ~x310 & ~x478 & ~x564 & ~x641 & ~x648 & ~x679 & ~x681 & ~x693 & ~x695 & ~x707 & ~x716 & ~x729 & ~x743 & ~x749 & ~x753 & ~x762 & ~x767 & ~x774;
assign c725 =  x432 & ~x15 & ~x22 & ~x38 & ~x84 & ~x95 & ~x174 & ~x178 & ~x230 & ~x231 & ~x247 & ~x285 & ~x323 & ~x420 & ~x423 & ~x447 & ~x485 & ~x505 & ~x539 & ~x552 & ~x596 & ~x650 & ~x666 & ~x698 & ~x699 & ~x783;
assign c727 =  x127;
assign c729 =  x666;
assign c733 =  x317 &  x373 & ~x18 & ~x19 & ~x22 & ~x27 & ~x31 & ~x32 & ~x38 & ~x58 & ~x61 & ~x65 & ~x68 & ~x78 & ~x81 & ~x96 & ~x98 & ~x107 & ~x113 & ~x122 & ~x128 & ~x165 & ~x172 & ~x199 & ~x229 & ~x230 & ~x231 & ~x232 & ~x251 & ~x259 & ~x284 & ~x307 & ~x309 & ~x321 & ~x332 & ~x334 & ~x341 & ~x342 & ~x361 & ~x368 & ~x369 & ~x395 & ~x397 & ~x415 & ~x424 & ~x479 & ~x495 & ~x553 & ~x561 & ~x606 & ~x618 & ~x637 & ~x639 & ~x664 & ~x673 & ~x695 & ~x750 & ~x757;
assign c735 =  x514 & ~x7 & ~x12 & ~x30 & ~x51 & ~x52 & ~x54 & ~x57 & ~x58 & ~x60 & ~x76 & ~x93 & ~x95 & ~x139 & ~x148 & ~x195 & ~x253 & ~x277 & ~x305 & ~x306 & ~x361 & ~x365 & ~x420 & ~x475 & ~x531 & ~x590 & ~x615 & ~x618 & ~x622 & ~x628 & ~x651 & ~x653 & ~x656 & ~x658 & ~x659 & ~x682 & ~x683 & ~x684 & ~x686 & ~x691 & ~x701 & ~x703 & ~x706 & ~x707 & ~x708 & ~x714 & ~x730 & ~x731 & ~x736 & ~x740 & ~x741 & ~x743 & ~x747 & ~x748 & ~x755 & ~x767;
assign c737 =  x378 & ~x5 & ~x13 & ~x19 & ~x22 & ~x35 & ~x57 & ~x68 & ~x74 & ~x75 & ~x77 & ~x102 & ~x107 & ~x116 & ~x141 & ~x228 & ~x250 & ~x251 & ~x256 & ~x283 & ~x312 & ~x313 & ~x360 & ~x364 & ~x368 & ~x369 & ~x392 & ~x413 & ~x424 & ~x426 & ~x451 & ~x453 & ~x454 & ~x462 & ~x531 & ~x544 & ~x585 & ~x615 & ~x616 & ~x639 & ~x675 & ~x698 & ~x753 & ~x766 & ~x776;
assign c739 =  x428 &  x485 &  x487 & ~x232 & ~x233;
assign c741 =  x434 & ~x0 & ~x23 & ~x32 & ~x63 & ~x84 & ~x126 & ~x197 & ~x282 & ~x307 & ~x501 & ~x531 & ~x562 & ~x599 & ~x600 & ~x602 & ~x671 & ~x679 & ~x708 & ~x723 & ~x773;
assign c743 =  x400 &  x457 &  x486;
assign c745 = ~x9 & ~x16 & ~x26 & ~x30 & ~x35 & ~x40 & ~x77 & ~x86 & ~x114 & ~x128 & ~x139 & ~x167 & ~x196 & ~x229 & ~x257 & ~x277 & ~x286 & ~x310 & ~x609 & ~x643 & ~x686 & ~x704 & ~x708 & ~x709 & ~x714 & ~x732 & ~x740 & ~x768 & ~x770 & ~x777;
assign c747 = ~x20 & ~x32 & ~x143 & ~x297 & ~x329 & ~x340 & ~x548 & ~x574 & ~x614 & ~x680 & ~x705 & ~x744 & ~x755 & ~x777;
assign c749 =  x399 & ~x2 & ~x68 & ~x130 & ~x143 & ~x227 & ~x253 & ~x266 & ~x346 & ~x418 & ~x563 & ~x620 & ~x628 & ~x671 & ~x702 & ~x725;
assign c751 =  x126;
assign c753 =  x350 &  x351 & ~x13 & ~x26 & ~x48 & ~x61 & ~x136 & ~x306 & ~x330 & ~x342 & ~x361 & ~x367 & ~x386 & ~x387 & ~x421 & ~x425 & ~x449 & ~x482 & ~x499 & ~x517 & ~x585 & ~x589 & ~x741 & ~x742 & ~x772;
assign c755 =  x327 &  x432 & ~x47 & ~x50 & ~x96 & ~x112 & ~x172 & ~x199 & ~x254 & ~x320 & ~x334 & ~x441 & ~x442 & ~x706 & ~x772;
assign c757 =  x181 &  x182 &  x208 &  x210 &  x609;
assign c759 =  x546 & ~x13 & ~x21 & ~x22 & ~x23 & ~x24 & ~x30 & ~x32 & ~x41 & ~x53 & ~x58 & ~x60 & ~x78 & ~x87 & ~x112 & ~x115 & ~x135 & ~x138 & ~x141 & ~x144 & ~x164 & ~x169 & ~x171 & ~x174 & ~x188 & ~x197 & ~x225 & ~x226 & ~x228 & ~x250 & ~x253 & ~x278 & ~x282 & ~x333 & ~x336 & ~x337 & ~x338 & ~x361 & ~x362 & ~x364 & ~x366 & ~x367 & ~x391 & ~x395 & ~x420 & ~x423 & ~x448 & ~x477 & ~x503 & ~x530 & ~x533 & ~x535 & ~x558 & ~x586 & ~x587 & ~x615 & ~x644 & ~x645 & ~x654 & ~x655 & ~x675 & ~x677 & ~x679 & ~x680 & ~x681 & ~x684 & ~x685 & ~x687 & ~x689 & ~x699 & ~x705 & ~x707 & ~x708 & ~x709 & ~x710 & ~x714 & ~x716 & ~x720 & ~x723 & ~x727 & ~x732 & ~x733 & ~x735 & ~x737 & ~x742 & ~x743 & ~x745 & ~x751 & ~x758 & ~x760 & ~x761 & ~x762 & ~x763 & ~x767 & ~x768 & ~x781;
assign c761 =  x346 &  x374 &  x432 & ~x231 & ~x314;
assign c763 = ~x145 & ~x160 & ~x177 & ~x302 & ~x318 & ~x353 & ~x420 & ~x586 & ~x647 & ~x660 & ~x678 & ~x683 & ~x685 & ~x708;
assign c765 =  x370 &  x458;
assign c767 =  x182 &  x348 & ~x6 & ~x32 & ~x37 & ~x39 & ~x84 & ~x94 & ~x313 & ~x338 & ~x340 & ~x456 & ~x471 & ~x481 & ~x501 & ~x669 & ~x721 & ~x763;
assign c769 =  x401 &  x458 &  x489 & ~x34 & ~x350 & ~x723;
assign c771 =  x344 &  x372 &  x430 &  x431 &  x432 & ~x470;
assign c773 =  x576 & ~x44 & ~x45 & ~x56 & ~x65 & ~x66 & ~x87 & ~x92 & ~x93 & ~x109 & ~x111 & ~x133 & ~x140 & ~x142 & ~x145 & ~x147 & ~x164 & ~x199 & ~x201 & ~x202 & ~x281 & ~x283 & ~x305 & ~x309 & ~x337 & ~x366 & ~x389 & ~x410 & ~x420 & ~x439 & ~x445 & ~x446 & ~x448 & ~x449 & ~x466 & ~x467 & ~x476 & ~x477 & ~x494 & ~x529 & ~x531 & ~x556 & ~x561 & ~x587 & ~x615 & ~x617 & ~x642 & ~x648 & ~x649 & ~x663 & ~x667 & ~x675 & ~x676 & ~x690 & ~x695 & ~x701 & ~x704 & ~x722 & ~x736 & ~x742 & ~x746 & ~x751 & ~x758 & ~x769 & ~x771 & ~x777 & ~x782;
assign c775 =  x372 &  x406 & ~x177 & ~x561;
assign c777 =  x211 &  x349 & ~x7 & ~x16 & ~x43 & ~x80 & ~x94 & ~x113 & ~x142 & ~x177 & ~x196 & ~x229 & ~x247 & ~x253 & ~x280 & ~x314 & ~x339 & ~x359 & ~x365 & ~x389 & ~x397 & ~x415 & ~x424 & ~x452 & ~x458 & ~x459 & ~x504 & ~x559 & ~x669 & ~x697 & ~x700 & ~x705 & ~x740 & ~x748;
assign c779 =  x432 &  x607;
assign c781 =  x405 &  x603 & ~x231 & ~x385 & ~x386 & ~x412 & ~x413 & ~x687 & ~x688 & ~x704;
assign c783 =  x426 & ~x65 & ~x685 & ~x686 & ~x688 & ~x707 & ~x745;
assign c785 =  x462 & ~x11 & ~x12 & ~x15 & ~x19 & ~x38 & ~x63 & ~x64 & ~x92 & ~x108 & ~x111 & ~x124 & ~x145 & ~x148 & ~x153 & ~x167 & ~x173 & ~x174 & ~x175 & ~x180 & ~x197 & ~x199 & ~x203 & ~x205 & ~x208 & ~x219 & ~x225 & ~x235 & ~x261 & ~x286 & ~x307 & ~x343 & ~x365 & ~x367 & ~x370 & ~x385 & ~x386 & ~x390 & ~x392 & ~x415 & ~x448 & ~x449 & ~x475 & ~x527 & ~x552 & ~x568 & ~x584 & ~x608 & ~x610 & ~x612 & ~x622 & ~x633 & ~x640 & ~x641 & ~x647 & ~x652 & ~x653 & ~x663 & ~x664 & ~x666 & ~x669 & ~x671 & ~x692 & ~x699 & ~x730 & ~x756 & ~x765 & ~x772 & ~x774;
assign c787 = ~x18 & ~x29 & ~x71 & ~x92 & ~x119 & ~x177 & ~x205 & ~x223 & ~x269 & ~x307 & ~x315 & ~x344 & ~x388 & ~x402 & ~x411 & ~x429 & ~x450 & ~x458 & ~x485 & ~x487 & ~x499 & ~x514 & ~x635 & ~x727 & ~x743 & ~x772 & ~x780;
assign c789 =  x319 &  x375 &  x403 & ~x313 & ~x413;
assign c791 =  x264 &  x433 & ~x20 & ~x49 & ~x90 & ~x193 & ~x257 & ~x296 & ~x334 & ~x535 & ~x586 & ~x635 & ~x675 & ~x724 & ~x755 & ~x772;
assign c793 =  x372 &  x400 &  x458 &  x459 &  x460 & ~x23 & ~x178 & ~x202 & ~x753;
assign c795 =  x625 & ~x2 & ~x21 & ~x77 & ~x79 & ~x82 & ~x116 & ~x137 & ~x284 & ~x437 & ~x473 & ~x529 & ~x677 & ~x707 & ~x708 & ~x709 & ~x710 & ~x723 & ~x731 & ~x738 & ~x748;
assign c797 = ~x7 & ~x8 & ~x26 & ~x42 & ~x60 & ~x63 & ~x68 & ~x70 & ~x83 & ~x141 & ~x148 & ~x151 & ~x164 & ~x177 & ~x179 & ~x204 & ~x207 & ~x225 & ~x230 & ~x231 & ~x289 & ~x298 & ~x309 & ~x311 & ~x344 & ~x354 & ~x365 & ~x410 & ~x411 & ~x418 & ~x484 & ~x495 & ~x522 & ~x533 & ~x535 & ~x539 & ~x540 & ~x565 & ~x578 & ~x633 & ~x640 & ~x691 & ~x718 & ~x728 & ~x755;
assign c799 = ~x263 & ~x298 & ~x326 & ~x338 & ~x422 & ~x433 & ~x464 & ~x710 & ~x774;
assign c7101 =  x377 & ~x10 & ~x30 & ~x40 & ~x47 & ~x59 & ~x65 & ~x70 & ~x79 & ~x86 & ~x99 & ~x115 & ~x194 & ~x222 & ~x251 & ~x281 & ~x339 & ~x357 & ~x384 & ~x415 & ~x425 & ~x443 & ~x444 & ~x454 & ~x485 & ~x487 & ~x512 & ~x513 & ~x531 & ~x532 & ~x544 & ~x545 & ~x555 & ~x614 & ~x618 & ~x667 & ~x720 & ~x722 & ~x724 & ~x749 & ~x754;
assign c7103 =  x542 & ~x18 & ~x25 & ~x32 & ~x36 & ~x38 & ~x47 & ~x51 & ~x83 & ~x85 & ~x105 & ~x106 & ~x136 & ~x137 & ~x162 & ~x166 & ~x171 & ~x186 & ~x194 & ~x196 & ~x198 & ~x222 & ~x225 & ~x248 & ~x251 & ~x308 & ~x335 & ~x337 & ~x363 & ~x391 & ~x392 & ~x420 & ~x474 & ~x475 & ~x532 & ~x534 & ~x535 & ~x588 & ~x616 & ~x619 & ~x620 & ~x621 & ~x640 & ~x644 & ~x648 & ~x649 & ~x651 & ~x652 & ~x653 & ~x656 & ~x658 & ~x660 & ~x661 & ~x662 & ~x667 & ~x668 & ~x669 & ~x670 & ~x671 & ~x676 & ~x682 & ~x687 & ~x694 & ~x703 & ~x705 & ~x708 & ~x709 & ~x713 & ~x720 & ~x738 & ~x739 & ~x740 & ~x741 & ~x745 & ~x747 & ~x760 & ~x762 & ~x764 & ~x765 & ~x776 & ~x777 & ~x782;
assign c7105 =  x511 & ~x81 & ~x230 & ~x660 & ~x684 & ~x686 & ~x715 & ~x758;
assign c7107 =  x628 & ~x8 & ~x22 & ~x40 & ~x41 & ~x43 & ~x70 & ~x87 & ~x92 & ~x101 & ~x103 & ~x109 & ~x111 & ~x135 & ~x144 & ~x166 & ~x195 & ~x196 & ~x197 & ~x307 & ~x310 & ~x364 & ~x367 & ~x399 & ~x416 & ~x419 & ~x426 & ~x448 & ~x481 & ~x483 & ~x517 & ~x616 & ~x645 & ~x697 & ~x712 & ~x715 & ~x718 & ~x724 & ~x728 & ~x730 & ~x735 & ~x737 & ~x739 & ~x744 & ~x765 & ~x774;
assign c7109 =  x352 &  x353 &  x379 & ~x2 & ~x6 & ~x12 & ~x24 & ~x27 & ~x38 & ~x40 & ~x42 & ~x47 & ~x50 & ~x58 & ~x59 & ~x60 & ~x65 & ~x66 & ~x67 & ~x68 & ~x70 & ~x72 & ~x80 & ~x83 & ~x86 & ~x90 & ~x93 & ~x96 & ~x99 & ~x100 & ~x103 & ~x106 & ~x114 & ~x128 & ~x129 & ~x130 & ~x139 & ~x145 & ~x158 & ~x172 & ~x173 & ~x174 & ~x177 & ~x191 & ~x193 & ~x194 & ~x199 & ~x222 & ~x224 & ~x225 & ~x226 & ~x227 & ~x253 & ~x276 & ~x277 & ~x305 & ~x308 & ~x311 & ~x313 & ~x332 & ~x335 & ~x359 & ~x361 & ~x364 & ~x365 & ~x368 & ~x370 & ~x386 & ~x395 & ~x396 & ~x398 & ~x400 & ~x411 & ~x412 & ~x416 & ~x419 & ~x420 & ~x423 & ~x425 & ~x428 & ~x441 & ~x445 & ~x449 & ~x453 & ~x454 & ~x471 & ~x479 & ~x481 & ~x495 & ~x498 & ~x499 & ~x501 & ~x507 & ~x529 & ~x534 & ~x538 & ~x554 & ~x559 & ~x560 & ~x563 & ~x587 & ~x593 & ~x614 & ~x618 & ~x641 & ~x644 & ~x670 & ~x674 & ~x697 & ~x700 & ~x704 & ~x720 & ~x731 & ~x732 & ~x739 & ~x742 & ~x746 & ~x747 & ~x750 & ~x751 & ~x752 & ~x754 & ~x755 & ~x759 & ~x763 & ~x765 & ~x766 & ~x768 & ~x769 & ~x770 & ~x773 & ~x776 & ~x777;
assign c7111 =  x458 & ~x2 & ~x3 & ~x5 & ~x11 & ~x15 & ~x16 & ~x20 & ~x23 & ~x40 & ~x64 & ~x67 & ~x76 & ~x80 & ~x104 & ~x107 & ~x117 & ~x130 & ~x132 & ~x134 & ~x140 & ~x146 & ~x149 & ~x161 & ~x167 & ~x168 & ~x196 & ~x228 & ~x232 & ~x247 & ~x253 & ~x280 & ~x282 & ~x306 & ~x313 & ~x322 & ~x323 & ~x324 & ~x337 & ~x366 & ~x390 & ~x392 & ~x444 & ~x445 & ~x447 & ~x482 & ~x501 & ~x505 & ~x536 & ~x583 & ~x618 & ~x619 & ~x620 & ~x675 & ~x702 & ~x704 & ~x723 & ~x727 & ~x737 & ~x738 & ~x743 & ~x749 & ~x751 & ~x765 & ~x766 & ~x769 & ~x774 & ~x776;
assign c7113 =  x485 & ~x6 & ~x32 & ~x38 & ~x48 & ~x61 & ~x68 & ~x83 & ~x87 & ~x135 & ~x172 & ~x200 & ~x364 & ~x394 & ~x446 & ~x587 & ~x641 & ~x657 & ~x660 & ~x680 & ~x683 & ~x699 & ~x703 & ~x714 & ~x731;
assign c7115 =  x185 & ~x62 & ~x208 & ~x263 & ~x686;
assign c7117 =  x208 & ~x20 & ~x26 & ~x34 & ~x47 & ~x69 & ~x84 & ~x104 & ~x105 & ~x137 & ~x142 & ~x172 & ~x177 & ~x178 & ~x199 & ~x201 & ~x203 & ~x256 & ~x283 & ~x285 & ~x312 & ~x332 & ~x337 & ~x338 & ~x339 & ~x346 & ~x360 & ~x395 & ~x413 & ~x414 & ~x415 & ~x418 & ~x468 & ~x533 & ~x536 & ~x561 & ~x583 & ~x591 & ~x592 & ~x597 & ~x599 & ~x608 & ~x609 & ~x695 & ~x736 & ~x752 & ~x761 & ~x769 & ~x782;
assign c7119 =  x433 &  x578;
assign c7121 = ~x6 & ~x8 & ~x9 & ~x10 & ~x32 & ~x34 & ~x42 & ~x45 & ~x63 & ~x66 & ~x77 & ~x79 & ~x89 & ~x100 & ~x107 & ~x113 & ~x116 & ~x120 & ~x122 & ~x137 & ~x144 & ~x145 & ~x146 & ~x148 & ~x153 & ~x169 & ~x174 & ~x179 & ~x181 & ~x198 & ~x206 & ~x207 & ~x208 & ~x223 & ~x225 & ~x226 & ~x228 & ~x229 & ~x235 & ~x236 & ~x253 & ~x255 & ~x256 & ~x261 & ~x263 & ~x284 & ~x288 & ~x290 & ~x310 & ~x314 & ~x318 & ~x333 & ~x334 & ~x335 & ~x338 & ~x341 & ~x345 & ~x365 & ~x367 & ~x369 & ~x371 & ~x372 & ~x385 & ~x387 & ~x391 & ~x394 & ~x396 & ~x397 & ~x416 & ~x440 & ~x441 & ~x450 & ~x452 & ~x469 & ~x471 & ~x477 & ~x480 & ~x497 & ~x501 & ~x504 & ~x505 & ~x528 & ~x529 & ~x530 & ~x534 & ~x535 & ~x555 & ~x556 & ~x558 & ~x564 & ~x585 & ~x588 & ~x607 & ~x613 & ~x614 & ~x642 & ~x646 & ~x651 & ~x669 & ~x670 & ~x671 & ~x692 & ~x694 & ~x712 & ~x717 & ~x719 & ~x722 & ~x729 & ~x730 & ~x739 & ~x741 & ~x749 & ~x754 & ~x760 & ~x770 & ~x771 & ~x772 & ~x776 & ~x783;
assign c7123 =  x347 & ~x0 & ~x3 & ~x6 & ~x16 & ~x38 & ~x40 & ~x51 & ~x55 & ~x62 & ~x65 & ~x71 & ~x117 & ~x141 & ~x280 & ~x301 & ~x326 & ~x359 & ~x388 & ~x392 & ~x396 & ~x419 & ~x446 & ~x481 & ~x537 & ~x556 & ~x640 & ~x646 & ~x669 & ~x670 & ~x671 & ~x692 & ~x694 & ~x735 & ~x737 & ~x746 & ~x747 & ~x766 & ~x768 & ~x770 & ~x775 & ~x778;
assign c7125 = ~x4 & ~x7 & ~x14 & ~x16 & ~x18 & ~x19 & ~x20 & ~x23 & ~x30 & ~x32 & ~x33 & ~x40 & ~x42 & ~x43 & ~x44 & ~x47 & ~x49 & ~x52 & ~x55 & ~x56 & ~x58 & ~x62 & ~x63 & ~x64 & ~x72 & ~x73 & ~x78 & ~x79 & ~x80 & ~x84 & ~x89 & ~x91 & ~x95 & ~x97 & ~x106 & ~x109 & ~x115 & ~x119 & ~x121 & ~x123 & ~x124 & ~x134 & ~x135 & ~x136 & ~x137 & ~x144 & ~x145 & ~x146 & ~x149 & ~x150 & ~x151 & ~x154 & ~x164 & ~x167 & ~x170 & ~x171 & ~x172 & ~x176 & ~x179 & ~x193 & ~x194 & ~x199 & ~x201 & ~x202 & ~x223 & ~x226 & ~x227 & ~x228 & ~x231 & ~x233 & ~x250 & ~x251 & ~x252 & ~x253 & ~x254 & ~x260 & ~x277 & ~x284 & ~x285 & ~x287 & ~x301 & ~x307 & ~x308 & ~x309 & ~x310 & ~x313 & ~x316 & ~x317 & ~x332 & ~x333 & ~x337 & ~x339 & ~x340 & ~x341 & ~x389 & ~x390 & ~x391 & ~x393 & ~x418 & ~x419 & ~x420 & ~x421 & ~x423 & ~x443 & ~x453 & ~x473 & ~x477 & ~x478 & ~x500 & ~x502 & ~x504 & ~x525 & ~x527 & ~x529 & ~x531 & ~x534 & ~x555 & ~x556 & ~x557 & ~x560 & ~x562 & ~x579 & ~x580 & ~x582 & ~x584 & ~x587 & ~x588 & ~x589 & ~x590 & ~x591 & ~x609 & ~x610 & ~x612 & ~x613 & ~x618 & ~x633 & ~x635 & ~x639 & ~x647 & ~x663 & ~x666 & ~x669 & ~x671 & ~x675 & ~x676 & ~x696 & ~x697 & ~x698 & ~x699 & ~x700 & ~x703 & ~x704 & ~x705 & ~x706 & ~x707 & ~x708 & ~x709 & ~x710 & ~x711 & ~x712 & ~x713 & ~x714 & ~x718 & ~x719 & ~x720 & ~x722 & ~x727 & ~x731 & ~x733 & ~x734 & ~x735 & ~x736 & ~x737 & ~x739 & ~x740 & ~x741 & ~x746 & ~x748 & ~x752 & ~x755 & ~x756 & ~x760 & ~x763 & ~x764 & ~x765 & ~x766 & ~x767 & ~x769 & ~x770 & ~x771 & ~x773 & ~x774 & ~x778 & ~x780 & ~x781 & ~x783;
assign c7127 =  x209 &  x262 & ~x6 & ~x14 & ~x19 & ~x20 & ~x33 & ~x54 & ~x61 & ~x63 & ~x66 & ~x71 & ~x73 & ~x81 & ~x82 & ~x86 & ~x88 & ~x96 & ~x97 & ~x106 & ~x109 & ~x119 & ~x122 & ~x135 & ~x138 & ~x144 & ~x149 & ~x150 & ~x162 & ~x176 & ~x198 & ~x199 & ~x203 & ~x204 & ~x221 & ~x222 & ~x225 & ~x230 & ~x231 & ~x232 & ~x250 & ~x281 & ~x308 & ~x311 & ~x312 & ~x361 & ~x363 & ~x424 & ~x471 & ~x499 & ~x505 & ~x530 & ~x562 & ~x590 & ~x609 & ~x611 & ~x612 & ~x639 & ~x640 & ~x641 & ~x666 & ~x697 & ~x701 & ~x704 & ~x726 & ~x731 & ~x743 & ~x747 & ~x758 & ~x763 & ~x767 & ~x772 & ~x783;
assign c7129 =  x511 & ~x233 & ~x261 & ~x325 & ~x688;
assign c7131 = ~x30 & ~x43 & ~x60 & ~x62 & ~x170 & ~x254 & ~x327 & ~x357 & ~x418 & ~x445 & ~x461 & ~x491 & ~x640 & ~x646 & ~x691 & ~x717 & ~x730 & ~x742 & ~x745 & ~x765 & ~x768 & ~x772;
assign c7133 =  x206 &  x580 & ~x548;
assign c7135 =  x188;
assign c7137 =  x182 &  x663;
assign c7139 = ~x20 & ~x63 & ~x101 & ~x178 & ~x190 & ~x256 & ~x267 & ~x295 & ~x304 & ~x358 & ~x387 & ~x391 & ~x444 & ~x466 & ~x494 & ~x506 & ~x534 & ~x557 & ~x647 & ~x679 & ~x698 & ~x702 & ~x708 & ~x755 & ~x765 & ~x772;
assign c7141 =  x548 & ~x22 & ~x41 & ~x82 & ~x92 & ~x96 & ~x101 & ~x113 & ~x163 & ~x169 & ~x172 & ~x177 & ~x203 & ~x228 & ~x250 & ~x254 & ~x303 & ~x330 & ~x331 & ~x362 & ~x363 & ~x365 & ~x393 & ~x414 & ~x423 & ~x440 & ~x442 & ~x445 & ~x447 & ~x466 & ~x469 & ~x470 & ~x477 & ~x495 & ~x550 & ~x555 & ~x564 & ~x620 & ~x673 & ~x697 & ~x700 & ~x722 & ~x759 & ~x777;
assign c7143 =  x377 & ~x8 & ~x19 & ~x40 & ~x110 & ~x136 & ~x267 & ~x305 & ~x360 & ~x385 & ~x440 & ~x453 & ~x588 & ~x638 & ~x669;
assign c7145 =  x607 & ~x414;
assign c7147 = ~x20 & ~x21 & ~x23 & ~x44 & ~x54 & ~x59 & ~x84 & ~x87 & ~x88 & ~x90 & ~x101 & ~x113 & ~x131 & ~x134 & ~x136 & ~x137 & ~x145 & ~x177 & ~x195 & ~x197 & ~x205 & ~x228 & ~x271 & ~x279 & ~x281 & ~x305 & ~x331 & ~x333 & ~x339 & ~x357 & ~x358 & ~x384 & ~x390 & ~x412 & ~x413 & ~x418 & ~x420 & ~x423 & ~x439 & ~x443 & ~x451 & ~x476 & ~x481 & ~x505 & ~x506 & ~x559 & ~x588 & ~x589 & ~x591 & ~x641 & ~x644 & ~x645 & ~x646 & ~x673 & ~x674 & ~x684 & ~x686 & ~x691 & ~x700 & ~x704 & ~x714 & ~x720 & ~x729 & ~x742 & ~x745 & ~x754 & ~x771 & ~x774 & ~x780 & ~x782;
assign c7149 =  x349 & ~x457 & ~x517;
assign c7151 = ~x11 & ~x25 & ~x37 & ~x45 & ~x116 & ~x154 & ~x155 & ~x169 & ~x182 & ~x183 & ~x193 & ~x197 & ~x199 & ~x211 & ~x223 & ~x249 & ~x251 & ~x266 & ~x282 & ~x294 & ~x320 & ~x321 & ~x347 & ~x362 & ~x366 & ~x367 & ~x390 & ~x473 & ~x558 & ~x616 & ~x638 & ~x667 & ~x669 & ~x694 & ~x699 & ~x702 & ~x703 & ~x705 & ~x711 & ~x723 & ~x728 & ~x737 & ~x738 & ~x739 & ~x756 & ~x758 & ~x765 & ~x779 & ~x783;
assign c7153 = ~x13 & ~x14 & ~x22 & ~x27 & ~x30 & ~x36 & ~x40 & ~x44 & ~x46 & ~x51 & ~x59 & ~x62 & ~x72 & ~x77 & ~x125 & ~x134 & ~x163 & ~x175 & ~x195 & ~x196 & ~x200 & ~x222 & ~x223 & ~x229 & ~x256 & ~x257 & ~x277 & ~x283 & ~x284 & ~x311 & ~x312 & ~x337 & ~x338 & ~x339 & ~x340 & ~x362 & ~x364 & ~x368 & ~x369 & ~x389 & ~x394 & ~x419 & ~x478 & ~x501 & ~x562 & ~x587 & ~x588 & ~x589 & ~x591 & ~x612 & ~x613 & ~x619 & ~x620 & ~x644 & ~x645 & ~x647 & ~x656 & ~x660 & ~x679 & ~x681 & ~x686 & ~x704 & ~x711 & ~x714 & ~x722 & ~x724 & ~x731 & ~x748 & ~x752 & ~x753 & ~x754 & ~x761 & ~x773;
assign c7155 =  x237 &  x291 &  x462 & ~x73 & ~x144 & ~x175 & ~x180 & ~x204 & ~x229 & ~x230 & ~x295 & ~x418 & ~x444 & ~x445 & ~x449 & ~x643 & ~x672 & ~x690;
assign c7157 = ~x28 & ~x119 & ~x179 & ~x235 & ~x271 & ~x280 & ~x286 & ~x309 & ~x318 & ~x329 & ~x358 & ~x403 & ~x410 & ~x411 & ~x412 & ~x465 & ~x466 & ~x678 & ~x687 & ~x691 & ~x727;
assign c7159 =  x271 &  x377 &  x405 & ~x2 & ~x47 & ~x67 & ~x73 & ~x98 & ~x101 & ~x138 & ~x283 & ~x369 & ~x416 & ~x469 & ~x668 & ~x696 & ~x704 & ~x754;
assign c7161 = ~x21 & ~x28 & ~x72 & ~x183 & ~x237 & ~x239 & ~x293 & ~x321 & ~x322 & ~x349 & ~x367 & ~x395 & ~x423 & ~x448 & ~x506 & ~x561 & ~x666 & ~x674 & ~x675 & ~x697 & ~x709 & ~x719 & ~x743 & ~x770;
assign c7163 =  x608;
assign c7165 =  x602 & ~x9 & ~x24 & ~x38 & ~x55 & ~x93 & ~x106 & ~x116 & ~x168 & ~x201 & ~x222 & ~x227 & ~x258 & ~x284 & ~x346 & ~x368 & ~x389 & ~x424 & ~x457 & ~x528 & ~x532 & ~x555 & ~x639 & ~x673 & ~x674 & ~x686 & ~x719 & ~x758 & ~x767 & ~x769 & ~x771;
assign c7167 =  x459 & ~x8 & ~x13 & ~x25 & ~x47 & ~x59 & ~x64 & ~x70 & ~x82 & ~x140 & ~x144 & ~x152 & ~x171 & ~x206 & ~x232 & ~x255 & ~x256 & ~x260 & ~x323 & ~x333 & ~x350 & ~x365 & ~x377 & ~x420 & ~x443 & ~x450 & ~x532 & ~x537 & ~x592 & ~x594 & ~x722 & ~x726 & ~x729 & ~x731 & ~x738 & ~x744;
assign c7169 =  x379 &  x491 & ~x1 & ~x8 & ~x10 & ~x11 & ~x17 & ~x19 & ~x24 & ~x25 & ~x31 & ~x38 & ~x41 & ~x43 & ~x54 & ~x56 & ~x59 & ~x60 & ~x66 & ~x67 & ~x72 & ~x74 & ~x76 & ~x78 & ~x80 & ~x81 & ~x87 & ~x89 & ~x90 & ~x92 & ~x94 & ~x101 & ~x103 & ~x105 & ~x108 & ~x110 & ~x118 & ~x133 & ~x140 & ~x148 & ~x149 & ~x150 & ~x175 & ~x176 & ~x178 & ~x192 & ~x194 & ~x198 & ~x199 & ~x203 & ~x205 & ~x206 & ~x221 & ~x231 & ~x249 & ~x255 & ~x259 & ~x277 & ~x279 & ~x281 & ~x282 & ~x287 & ~x288 & ~x304 & ~x314 & ~x316 & ~x333 & ~x334 & ~x339 & ~x343 & ~x357 & ~x359 & ~x362 & ~x366 & ~x385 & ~x390 & ~x392 & ~x393 & ~x398 & ~x411 & ~x413 & ~x414 & ~x417 & ~x423 & ~x426 & ~x429 & ~x442 & ~x448 & ~x451 & ~x457 & ~x458 & ~x466 & ~x473 & ~x476 & ~x477 & ~x481 & ~x482 & ~x484 & ~x485 & ~x486 & ~x494 & ~x497 & ~x504 & ~x507 & ~x508 & ~x510 & ~x513 & ~x523 & ~x532 & ~x540 & ~x554 & ~x558 & ~x580 & ~x581 & ~x583 & ~x588 & ~x589 & ~x592 & ~x606 & ~x608 & ~x609 & ~x610 & ~x611 & ~x615 & ~x637 & ~x642 & ~x643 & ~x649 & ~x670 & ~x672 & ~x675 & ~x689 & ~x695 & ~x697 & ~x701 & ~x717 & ~x725 & ~x728 & ~x731 & ~x741 & ~x742 & ~x743 & ~x745 & ~x747 & ~x751 & ~x753 & ~x756 & ~x759 & ~x760 & ~x765 & ~x766 & ~x768 & ~x769 & ~x772 & ~x782;
assign c7171 =  x568 & ~x87 & ~x121 & ~x309 & ~x380 & ~x637 & ~x648 & ~x705;
assign c7173 =  x323 & ~x7 & ~x9 & ~x13 & ~x22 & ~x24 & ~x27 & ~x36 & ~x42 & ~x47 & ~x49 & ~x63 & ~x64 & ~x66 & ~x85 & ~x95 & ~x96 & ~x110 & ~x112 & ~x134 & ~x137 & ~x138 & ~x151 & ~x165 & ~x167 & ~x171 & ~x178 & ~x192 & ~x198 & ~x204 & ~x206 & ~x207 & ~x219 & ~x220 & ~x223 & ~x227 & ~x230 & ~x246 & ~x247 & ~x248 & ~x259 & ~x262 & ~x276 & ~x283 & ~x286 & ~x301 & ~x303 & ~x310 & ~x317 & ~x337 & ~x339 & ~x344 & ~x356 & ~x367 & ~x372 & ~x375 & ~x392 & ~x396 & ~x402 & ~x412 & ~x413 & ~x417 & ~x425 & ~x429 & ~x439 & ~x442 & ~x445 & ~x452 & ~x466 & ~x467 & ~x470 & ~x477 & ~x493 & ~x506 & ~x535 & ~x581 & ~x609 & ~x612 & ~x616 & ~x634 & ~x636 & ~x638 & ~x650 & ~x666 & ~x674 & ~x692 & ~x699 & ~x707 & ~x718 & ~x719 & ~x734 & ~x735 & ~x739 & ~x755 & ~x759 & ~x763 & ~x768 & ~x774 & ~x776 & ~x779;
assign c7175 = ~x2 & ~x7 & ~x14 & ~x15 & ~x25 & ~x36 & ~x42 & ~x53 & ~x64 & ~x73 & ~x79 & ~x92 & ~x99 & ~x105 & ~x109 & ~x112 & ~x144 & ~x163 & ~x171 & ~x178 & ~x187 & ~x191 & ~x199 & ~x214 & ~x224 & ~x327 & ~x333 & ~x345 & ~x357 & ~x369 & ~x383 & ~x384 & ~x395 & ~x412 & ~x421 & ~x441 & ~x475 & ~x476 & ~x493 & ~x532 & ~x559 & ~x566 & ~x588 & ~x619 & ~x645 & ~x706 & ~x708 & ~x712 & ~x719 & ~x744 & ~x748 & ~x755 & ~x777 & ~x783;
assign c7177 = ~x0 & ~x1 & ~x7 & ~x12 & ~x17 & ~x19 & ~x22 & ~x29 & ~x30 & ~x31 & ~x32 & ~x35 & ~x37 & ~x40 & ~x41 & ~x54 & ~x59 & ~x62 & ~x63 & ~x66 & ~x74 & ~x81 & ~x85 & ~x86 & ~x87 & ~x89 & ~x92 & ~x93 & ~x97 & ~x102 & ~x116 & ~x117 & ~x128 & ~x130 & ~x132 & ~x134 & ~x136 & ~x137 & ~x145 & ~x147 & ~x148 & ~x162 & ~x165 & ~x169 & ~x170 & ~x173 & ~x174 & ~x176 & ~x177 & ~x191 & ~x192 & ~x200 & ~x201 & ~x218 & ~x222 & ~x224 & ~x227 & ~x229 & ~x248 & ~x252 & ~x253 & ~x257 & ~x276 & ~x280 & ~x284 & ~x306 & ~x309 & ~x332 & ~x366 & ~x386 & ~x389 & ~x392 & ~x396 & ~x414 & ~x415 & ~x422 & ~x440 & ~x441 & ~x442 & ~x447 & ~x449 & ~x470 & ~x472 & ~x473 & ~x479 & ~x480 & ~x481 & ~x483 & ~x496 & ~x498 & ~x501 & ~x504 & ~x510 & ~x512 & ~x518 & ~x528 & ~x529 & ~x533 & ~x534 & ~x535 & ~x538 & ~x539 & ~x544 & ~x554 & ~x555 & ~x556 & ~x558 & ~x559 & ~x562 & ~x565 & ~x572 & ~x583 & ~x584 & ~x585 & ~x594 & ~x595 & ~x610 & ~x614 & ~x616 & ~x618 & ~x620 & ~x637 & ~x645 & ~x665 & ~x676 & ~x677 & ~x693 & ~x699 & ~x702 & ~x703 & ~x722 & ~x725 & ~x728 & ~x735 & ~x750 & ~x754 & ~x756 & ~x759 & ~x760 & ~x764 & ~x766 & ~x772 & ~x777 & ~x779 & ~x783;
assign c7179 =  x553 & ~x71 & ~x126 & ~x168 & ~x290 & ~x291 & ~x535 & ~x750 & ~x761;
assign c7181 =  x210 &  x550 & ~x8 & ~x13 & ~x24 & ~x55 & ~x77 & ~x78 & ~x106 & ~x137 & ~x172 & ~x174 & ~x253 & ~x280 & ~x332 & ~x339 & ~x389 & ~x532 & ~x587 & ~x689 & ~x693 & ~x714 & ~x718 & ~x719 & ~x725 & ~x741 & ~x758;
assign c7183 =  x153 &  x347;
assign c7185 = ~x20 & ~x41 & ~x82 & ~x84 & ~x101 & ~x183 & ~x239 & ~x281 & ~x294 & ~x311 & ~x351 & ~x390 & ~x587 & ~x592 & ~x701 & ~x770;
assign c7187 = ~x0 & ~x9 & ~x11 & ~x17 & ~x22 & ~x23 & ~x24 & ~x26 & ~x27 & ~x33 & ~x35 & ~x36 & ~x37 & ~x39 & ~x43 & ~x48 & ~x51 & ~x55 & ~x59 & ~x61 & ~x62 & ~x65 & ~x66 & ~x67 & ~x69 & ~x77 & ~x78 & ~x81 & ~x82 & ~x84 & ~x89 & ~x93 & ~x97 & ~x112 & ~x116 & ~x118 & ~x127 & ~x128 & ~x130 & ~x133 & ~x134 & ~x135 & ~x138 & ~x139 & ~x141 & ~x142 & ~x144 & ~x145 & ~x147 & ~x149 & ~x164 & ~x166 & ~x167 & ~x169 & ~x171 & ~x172 & ~x173 & ~x174 & ~x192 & ~x203 & ~x204 & ~x205 & ~x222 & ~x226 & ~x231 & ~x250 & ~x251 & ~x253 & ~x255 & ~x258 & ~x260 & ~x287 & ~x303 & ~x305 & ~x310 & ~x311 & ~x312 & ~x314 & ~x334 & ~x337 & ~x358 & ~x360 & ~x363 & ~x367 & ~x369 & ~x384 & ~x386 & ~x388 & ~x389 & ~x392 & ~x394 & ~x395 & ~x397 & ~x413 & ~x414 & ~x415 & ~x422 & ~x423 & ~x425 & ~x443 & ~x451 & ~x452 & ~x470 & ~x474 & ~x475 & ~x482 & ~x496 & ~x501 & ~x502 & ~x504 & ~x506 & ~x507 & ~x511 & ~x524 & ~x527 & ~x533 & ~x534 & ~x538 & ~x543 & ~x553 & ~x560 & ~x561 & ~x566 & ~x578 & ~x581 & ~x583 & ~x586 & ~x606 & ~x608 & ~x609 & ~x612 & ~x614 & ~x617 & ~x618 & ~x634 & ~x639 & ~x641 & ~x662 & ~x664 & ~x665 & ~x672 & ~x673 & ~x676 & ~x689 & ~x698 & ~x700 & ~x701 & ~x702 & ~x703 & ~x707 & ~x718 & ~x725 & ~x731 & ~x733 & ~x734 & ~x736 & ~x737 & ~x743 & ~x747 & ~x749 & ~x751 & ~x754 & ~x755 & ~x757 & ~x758 & ~x764 & ~x768 & ~x772;
assign c7189 =  x405 & ~x4 & ~x162 & ~x174 & ~x414 & ~x439 & ~x516 & ~x534 & ~x563;
assign c7191 =  x345 &  x404 &  x406 & ~x118 & ~x471;
assign c7193 =  x373 &  x458 &  x462 & ~x377;
assign c7195 =  x461 & ~x18 & ~x22 & ~x43 & ~x44 & ~x58 & ~x69 & ~x77 & ~x112 & ~x115 & ~x136 & ~x166 & ~x195 & ~x227 & ~x232 & ~x251 & ~x255 & ~x259 & ~x280 & ~x284 & ~x285 & ~x351 & ~x364 & ~x396 & ~x397 & ~x421 & ~x448 & ~x504 & ~x530 & ~x534 & ~x565 & ~x652 & ~x677 & ~x695 & ~x707 & ~x709 & ~x722 & ~x730 & ~x745 & ~x752 & ~x764;
assign c7197 =  x373 &  x430 &  x461 & ~x172 & ~x257 & ~x391 & ~x762;
assign c7199 =  x156 &  x654;
assign c7201 =  x578 &  x656;
assign c7203 = ~x2 & ~x3 & ~x5 & ~x6 & ~x10 & ~x13 & ~x16 & ~x26 & ~x31 & ~x35 & ~x40 & ~x43 & ~x45 & ~x51 & ~x52 & ~x53 & ~x54 & ~x56 & ~x58 & ~x65 & ~x71 & ~x74 & ~x90 & ~x91 & ~x103 & ~x105 & ~x110 & ~x116 & ~x121 & ~x138 & ~x149 & ~x150 & ~x166 & ~x168 & ~x169 & ~x170 & ~x172 & ~x179 & ~x180 & ~x181 & ~x191 & ~x202 & ~x203 & ~x221 & ~x223 & ~x231 & ~x233 & ~x251 & ~x252 & ~x254 & ~x256 & ~x258 & ~x259 & ~x260 & ~x276 & ~x281 & ~x283 & ~x284 & ~x285 & ~x286 & ~x306 & ~x307 & ~x313 & ~x321 & ~x333 & ~x335 & ~x338 & ~x340 & ~x359 & ~x361 & ~x363 & ~x388 & ~x390 & ~x391 & ~x392 & ~x415 & ~x419 & ~x424 & ~x439 & ~x443 & ~x445 & ~x449 & ~x452 & ~x474 & ~x476 & ~x477 & ~x480 & ~x495 & ~x510 & ~x523 & ~x529 & ~x530 & ~x532 & ~x536 & ~x537 & ~x538 & ~x541 & ~x566 & ~x580 & ~x581 & ~x583 & ~x584 & ~x586 & ~x587 & ~x588 & ~x589 & ~x598 & ~x609 & ~x622 & ~x624 & ~x635 & ~x640 & ~x644 & ~x653 & ~x662 & ~x663 & ~x666 & ~x667 & ~x670 & ~x676 & ~x680 & ~x691 & ~x695 & ~x697 & ~x698 & ~x720 & ~x721 & ~x728 & ~x730 & ~x731 & ~x732 & ~x751 & ~x757 & ~x759 & ~x769 & ~x775 & ~x782;
assign c7205 =  x123;
assign c7207 =  x634 & ~x250 & ~x252 & ~x469 & ~x506;
assign c7209 =  x488 &  x578 & ~x203 & ~x538;
assign c7211 =  x372 &  x400 &  x460 & ~x441;
assign c7213 =  x158 & ~x151;
assign c7215 =  x455 &  x551;
assign c7217 =  x318 &  x375 &  x404 & ~x59 & ~x94 & ~x258 & ~x457 & ~x481 & ~x510 & ~x563 & ~x728 & ~x769;
assign c7219 =  x568 & ~x271;
assign c7221 =  x566 & ~x123 & ~x313;
assign c7223 =  x606 & ~x1 & ~x45 & ~x65 & ~x341 & ~x451 & ~x528;
assign c7225 =  x405 & ~x8 & ~x18 & ~x20 & ~x22 & ~x25 & ~x28 & ~x31 & ~x33 & ~x38 & ~x40 & ~x44 & ~x46 & ~x56 & ~x58 & ~x59 & ~x61 & ~x65 & ~x66 & ~x71 & ~x73 & ~x76 & ~x79 & ~x80 & ~x92 & ~x100 & ~x101 & ~x106 & ~x109 & ~x111 & ~x113 & ~x114 & ~x117 & ~x120 & ~x123 & ~x124 & ~x127 & ~x129 & ~x131 & ~x138 & ~x143 & ~x145 & ~x148 & ~x149 & ~x150 & ~x152 & ~x163 & ~x167 & ~x170 & ~x171 & ~x173 & ~x178 & ~x193 & ~x194 & ~x198 & ~x200 & ~x223 & ~x225 & ~x229 & ~x250 & ~x252 & ~x256 & ~x279 & ~x283 & ~x284 & ~x305 & ~x310 & ~x313 & ~x331 & ~x332 & ~x339 & ~x340 & ~x358 & ~x359 & ~x362 & ~x363 & ~x368 & ~x387 & ~x388 & ~x389 & ~x392 & ~x396 & ~x411 & ~x417 & ~x421 & ~x424 & ~x425 & ~x441 & ~x442 & ~x452 & ~x453 & ~x475 & ~x477 & ~x479 & ~x480 & ~x484 & ~x496 & ~x504 & ~x508 & ~x511 & ~x527 & ~x529 & ~x533 & ~x555 & ~x560 & ~x564 & ~x580 & ~x584 & ~x585 & ~x608 & ~x613 & ~x616 & ~x619 & ~x637 & ~x643 & ~x646 & ~x647 & ~x666 & ~x669 & ~x670 & ~x671 & ~x693 & ~x696 & ~x699 & ~x733 & ~x738 & ~x747 & ~x750 & ~x757 & ~x759 & ~x760 & ~x766 & ~x770 & ~x774 & ~x778 & ~x779 & ~x781;
assign c7227 =  x570 & ~x15 & ~x23 & ~x29 & ~x37 & ~x48 & ~x52 & ~x58 & ~x60 & ~x65 & ~x70 & ~x74 & ~x83 & ~x84 & ~x105 & ~x108 & ~x196 & ~x227 & ~x229 & ~x251 & ~x277 & ~x367 & ~x418 & ~x419 & ~x476 & ~x503 & ~x558 & ~x614 & ~x641 & ~x648 & ~x651 & ~x652 & ~x653 & ~x667 & ~x677 & ~x684 & ~x692 & ~x693 & ~x700 & ~x702 & ~x707 & ~x709 & ~x710 & ~x711 & ~x714 & ~x715 & ~x718 & ~x723 & ~x730 & ~x733 & ~x735 & ~x751 & ~x755 & ~x778 & ~x780;
assign c7229 =  x581;
assign c7231 =  x574 & ~x31 & ~x64 & ~x133 & ~x178 & ~x197 & ~x199 & ~x205 & ~x231 & ~x258 & ~x268 & ~x269 & ~x311 & ~x342 & ~x387 & ~x451 & ~x473 & ~x480 & ~x530 & ~x555 & ~x614 & ~x636 & ~x698 & ~x743;
assign c7233 =  x372 &  x405 & ~x12 & ~x80 & ~x358 & ~x418 & ~x480;
assign c7235 = ~x6 & ~x16 & ~x36 & ~x39 & ~x43 & ~x44 & ~x45 & ~x55 & ~x63 & ~x67 & ~x71 & ~x74 & ~x75 & ~x78 & ~x79 & ~x82 & ~x103 & ~x111 & ~x118 & ~x120 & ~x121 & ~x142 & ~x143 & ~x144 & ~x148 & ~x169 & ~x171 & ~x172 & ~x174 & ~x175 & ~x195 & ~x224 & ~x228 & ~x282 & ~x283 & ~x297 & ~x305 & ~x306 & ~x308 & ~x309 & ~x323 & ~x324 & ~x335 & ~x341 & ~x357 & ~x359 & ~x360 & ~x364 & ~x365 & ~x366 & ~x369 & ~x387 & ~x390 & ~x414 & ~x415 & ~x419 & ~x422 & ~x441 & ~x445 & ~x449 & ~x467 & ~x468 & ~x471 & ~x480 & ~x482 & ~x495 & ~x496 & ~x497 & ~x498 & ~x499 & ~x524 & ~x527 & ~x536 & ~x559 & ~x562 & ~x565 & ~x585 & ~x586 & ~x589 & ~x616 & ~x641 & ~x645 & ~x676 & ~x694 & ~x703 & ~x720 & ~x723 & ~x725 & ~x726 & ~x728 & ~x729 & ~x743 & ~x749 & ~x756 & ~x759 & ~x761 & ~x764 & ~x780;
assign c7237 = ~x7 & ~x17 & ~x29 & ~x31 & ~x51 & ~x60 & ~x73 & ~x76 & ~x77 & ~x84 & ~x119 & ~x132 & ~x146 & ~x159 & ~x219 & ~x226 & ~x253 & ~x274 & ~x275 & ~x283 & ~x290 & ~x309 & ~x317 & ~x333 & ~x508 & ~x592 & ~x594 & ~x615 & ~x660 & ~x677 & ~x680 & ~x681 & ~x682 & ~x683 & ~x685 & ~x686 & ~x687 & ~x708 & ~x711 & ~x712 & ~x726 & ~x741 & ~x748 & ~x749 & ~x778;
assign c7239 = ~x9 & ~x15 & ~x18 & ~x23 & ~x25 & ~x26 & ~x27 & ~x29 & ~x36 & ~x41 & ~x42 & ~x43 & ~x44 & ~x46 & ~x48 & ~x50 & ~x51 & ~x60 & ~x68 & ~x75 & ~x76 & ~x81 & ~x82 & ~x83 & ~x86 & ~x97 & ~x98 & ~x104 & ~x113 & ~x114 & ~x126 & ~x135 & ~x142 & ~x145 & ~x149 & ~x163 & ~x164 & ~x165 & ~x168 & ~x175 & ~x180 & ~x181 & ~x195 & ~x205 & ~x232 & ~x233 & ~x235 & ~x250 & ~x257 & ~x261 & ~x280 & ~x281 & ~x282 & ~x284 & ~x288 & ~x309 & ~x310 & ~x312 & ~x317 & ~x327 & ~x328 & ~x357 & ~x359 & ~x363 & ~x365 & ~x367 & ~x369 & ~x391 & ~x397 & ~x416 & ~x417 & ~x421 & ~x422 & ~x424 & ~x444 & ~x447 & ~x475 & ~x478 & ~x479 & ~x507 & ~x525 & ~x527 & ~x528 & ~x529 & ~x531 & ~x533 & ~x556 & ~x557 & ~x559 & ~x579 & ~x582 & ~x584 & ~x590 & ~x609 & ~x610 & ~x612 & ~x613 & ~x614 & ~x618 & ~x619 & ~x641 & ~x644 & ~x645 & ~x674 & ~x688 & ~x689 & ~x691 & ~x700 & ~x702 & ~x705 & ~x711 & ~x713 & ~x714 & ~x718 & ~x719 & ~x721 & ~x722 & ~x723 & ~x726 & ~x730 & ~x731 & ~x732 & ~x746 & ~x750 & ~x753 & ~x756 & ~x757 & ~x774 & ~x776 & ~x777;
assign c7241 =  x122;
assign c7243 =  x317 & ~x0 & ~x3 & ~x11 & ~x17 & ~x19 & ~x23 & ~x52 & ~x56 & ~x57 & ~x75 & ~x81 & ~x88 & ~x102 & ~x109 & ~x137 & ~x168 & ~x173 & ~x191 & ~x201 & ~x252 & ~x255 & ~x257 & ~x258 & ~x259 & ~x293 & ~x301 & ~x313 & ~x334 & ~x335 & ~x338 & ~x340 & ~x341 & ~x369 & ~x391 & ~x393 & ~x467 & ~x480 & ~x494 & ~x495 & ~x496 & ~x502 & ~x522 & ~x527 & ~x551 & ~x591 & ~x676 & ~x677 & ~x695 & ~x708 & ~x750 & ~x761 & ~x762 & ~x769 & ~x770;
assign c7245 =  x160;
assign c7247 =  x292 & ~x30 & ~x70 & ~x232 & ~x345 & ~x458;
assign c7249 =  x372 &  x428 &  x459 & ~x203 & ~x375 & ~x395 & ~x423 & ~x510 & ~x706 & ~x755;
assign c7251 =  x182 &  x605 & ~x2 & ~x17 & ~x23 & ~x45 & ~x55 & ~x56 & ~x67 & ~x78 & ~x79 & ~x105 & ~x107 & ~x116 & ~x132 & ~x137 & ~x141 & ~x145 & ~x166 & ~x193 & ~x197 & ~x342 & ~x369 & ~x394 & ~x395 & ~x423 & ~x448 & ~x451 & ~x531 & ~x561 & ~x564 & ~x674 & ~x690 & ~x695 & ~x704 & ~x717 & ~x727 & ~x732 & ~x744 & ~x755 & ~x758 & ~x773;
assign c7253 =  x212 &  x376 &  x377 & ~x251 & ~x340 & ~x396 & ~x414 & ~x425 & ~x528 & ~x532 & ~x698;
assign c7255 =  x524 & ~x2 & ~x220 & ~x325 & ~x392 & ~x479 & ~x709 & ~x715 & ~x716 & ~x717;
assign c7257 =  x405 & ~x10 & ~x15 & ~x23 & ~x25 & ~x32 & ~x35 & ~x38 & ~x44 & ~x47 & ~x74 & ~x81 & ~x95 & ~x102 & ~x118 & ~x122 & ~x125 & ~x141 & ~x144 & ~x146 & ~x155 & ~x162 & ~x163 & ~x168 & ~x200 & ~x202 & ~x223 & ~x334 & ~x339 & ~x362 & ~x363 & ~x367 & ~x390 & ~x413 & ~x416 & ~x441 & ~x442 & ~x443 & ~x461 & ~x480 & ~x508 & ~x532 & ~x563 & ~x613 & ~x668 & ~x671 & ~x675 & ~x696 & ~x698 & ~x701 & ~x729 & ~x730 & ~x754;
assign c7259 =  x659 &  x660 & ~x23 & ~x25 & ~x105 & ~x108 & ~x168 & ~x194 & ~x226 & ~x447 & ~x502 & ~x504 & ~x558 & ~x575 & ~x668 & ~x675 & ~x716 & ~x719 & ~x721 & ~x727 & ~x743 & ~x744;
assign c7261 =  x399 &  x456 &  x486;
assign c7263 = ~x34 & ~x97 & ~x207 & ~x218 & ~x234 & ~x317 & ~x327 & ~x339 & ~x372 & ~x385 & ~x412 & ~x438 & ~x466 & ~x683 & ~x712;
assign c7265 =  x461 &  x577 & ~x14 & ~x39 & ~x67 & ~x86 & ~x98 & ~x99 & ~x133 & ~x175 & ~x176 & ~x201 & ~x220 & ~x225 & ~x229 & ~x254 & ~x305 & ~x339 & ~x443 & ~x448 & ~x471 & ~x764 & ~x771;
assign c7267 =  x543 & ~x9 & ~x19 & ~x27 & ~x37 & ~x39 & ~x53 & ~x54 & ~x68 & ~x81 & ~x85 & ~x104 & ~x106 & ~x109 & ~x110 & ~x114 & ~x117 & ~x118 & ~x137 & ~x142 & ~x163 & ~x167 & ~x170 & ~x171 & ~x196 & ~x219 & ~x223 & ~x253 & ~x306 & ~x308 & ~x310 & ~x334 & ~x339 & ~x361 & ~x366 & ~x391 & ~x392 & ~x394 & ~x421 & ~x447 & ~x451 & ~x453 & ~x537 & ~x561 & ~x585 & ~x587 & ~x589 & ~x616 & ~x617 & ~x618 & ~x643 & ~x648 & ~x651 & ~x656 & ~x658 & ~x667 & ~x678 & ~x681 & ~x687 & ~x696 & ~x707 & ~x711 & ~x714 & ~x716 & ~x717 & ~x737 & ~x742 & ~x746 & ~x753 & ~x754 & ~x757 & ~x767 & ~x769 & ~x779 & ~x781;
assign c7269 =  x548 & ~x12 & ~x25 & ~x27 & ~x41 & ~x53 & ~x59 & ~x60 & ~x62 & ~x63 & ~x66 & ~x76 & ~x81 & ~x84 & ~x85 & ~x88 & ~x111 & ~x121 & ~x136 & ~x137 & ~x138 & ~x139 & ~x144 & ~x146 & ~x162 & ~x169 & ~x174 & ~x177 & ~x190 & ~x216 & ~x220 & ~x228 & ~x231 & ~x251 & ~x256 & ~x283 & ~x293 & ~x312 & ~x313 & ~x330 & ~x334 & ~x337 & ~x391 & ~x423 & ~x451 & ~x475 & ~x477 & ~x504 & ~x535 & ~x566 & ~x587 & ~x588 & ~x594 & ~x636 & ~x665 & ~x674 & ~x677 & ~x726 & ~x729 & ~x732 & ~x737 & ~x738 & ~x750 & ~x753 & ~x754 & ~x757 & ~x759 & ~x765 & ~x773 & ~x774 & ~x776 & ~x777 & ~x778;
assign c7271 =  x404 &  x519 & ~x99 & ~x110 & ~x138 & ~x225 & ~x284 & ~x294 & ~x312 & ~x472 & ~x534 & ~x696 & ~x738 & ~x762;
assign c7273 =  x573 & ~x235 & ~x290 & ~x317 & ~x383 & ~x396 & ~x685 & ~x709 & ~x739;
assign c7275 =  x487 & ~x32 & ~x40 & ~x95 & ~x116 & ~x257 & ~x269 & ~x296 & ~x419 & ~x526 & ~x739;
assign c7277 =  x455 &  x513 &  x515;
assign c7279 =  x608 & ~x711;
assign c7281 = ~x1 & ~x10 & ~x15 & ~x25 & ~x26 & ~x30 & ~x31 & ~x33 & ~x36 & ~x39 & ~x44 & ~x46 & ~x47 & ~x56 & ~x57 & ~x61 & ~x65 & ~x67 & ~x71 & ~x80 & ~x92 & ~x94 & ~x104 & ~x105 & ~x106 & ~x116 & ~x117 & ~x131 & ~x137 & ~x139 & ~x141 & ~x167 & ~x169 & ~x176 & ~x177 & ~x185 & ~x195 & ~x197 & ~x204 & ~x229 & ~x230 & ~x242 & ~x255 & ~x257 & ~x258 & ~x270 & ~x278 & ~x279 & ~x280 & ~x281 & ~x283 & ~x306 & ~x309 & ~x316 & ~x336 & ~x338 & ~x341 & ~x344 & ~x364 & ~x367 & ~x368 & ~x395 & ~x411 & ~x425 & ~x452 & ~x475 & ~x507 & ~x508 & ~x509 & ~x529 & ~x532 & ~x533 & ~x534 & ~x580 & ~x581 & ~x590 & ~x591 & ~x614 & ~x644 & ~x649 & ~x663 & ~x664 & ~x665 & ~x698 & ~x702 & ~x704 & ~x705 & ~x714 & ~x716 & ~x717 & ~x725 & ~x728 & ~x734 & ~x737 & ~x739 & ~x742 & ~x753 & ~x756 & ~x760 & ~x762 & ~x763 & ~x767 & ~x774 & ~x775 & ~x780;
assign c7283 =  x375 &  x408 & ~x89 & ~x276 & ~x386 & ~x596;
assign c7285 = ~x7 & ~x12 & ~x15 & ~x17 & ~x24 & ~x27 & ~x34 & ~x36 & ~x39 & ~x43 & ~x51 & ~x54 & ~x59 & ~x61 & ~x64 & ~x66 & ~x78 & ~x98 & ~x104 & ~x121 & ~x124 & ~x125 & ~x133 & ~x139 & ~x140 & ~x143 & ~x153 & ~x172 & ~x177 & ~x193 & ~x203 & ~x207 & ~x208 & ~x226 & ~x235 & ~x254 & ~x258 & ~x279 & ~x283 & ~x284 & ~x285 & ~x287 & ~x289 & ~x314 & ~x317 & ~x333 & ~x339 & ~x394 & ~x411 & ~x412 & ~x420 & ~x421 & ~x424 & ~x438 & ~x445 & ~x446 & ~x467 & ~x470 & ~x475 & ~x478 & ~x480 & ~x492 & ~x495 & ~x498 & ~x500 & ~x501 & ~x523 & ~x528 & ~x530 & ~x531 & ~x553 & ~x557 & ~x565 & ~x582 & ~x584 & ~x608 & ~x613 & ~x614 & ~x617 & ~x618 & ~x621 & ~x634 & ~x640 & ~x642 & ~x646 & ~x647 & ~x649 & ~x650 & ~x665 & ~x668 & ~x676 & ~x699 & ~x700 & ~x704 & ~x711 & ~x714 & ~x720 & ~x722 & ~x723 & ~x725 & ~x734 & ~x738 & ~x740 & ~x742 & ~x750 & ~x771 & ~x774 & ~x775 & ~x778;
assign c7287 =  x344 &  x430 &  x432 & ~x66 & ~x507 & ~x508;
assign c7289 =  x373 &  x430 &  x460 & ~x498;
assign c7291 =  x374 &  x433 & ~x112 & ~x441 & ~x731;
assign c7293 =  x348 &  x376 &  x406 & ~x5 & ~x58 & ~x398 & ~x439 & ~x443 & ~x470;
assign c7295 =  x595 & ~x648 & ~x678 & ~x718;
assign c7297 =  x376 & ~x16 & ~x21 & ~x24 & ~x25 & ~x31 & ~x39 & ~x46 & ~x49 & ~x59 & ~x65 & ~x69 & ~x86 & ~x88 & ~x91 & ~x92 & ~x94 & ~x101 & ~x103 & ~x106 & ~x121 & ~x136 & ~x137 & ~x138 & ~x142 & ~x147 & ~x162 & ~x173 & ~x194 & ~x195 & ~x228 & ~x254 & ~x281 & ~x284 & ~x305 & ~x306 & ~x311 & ~x338 & ~x339 & ~x369 & ~x389 & ~x397 & ~x412 & ~x413 & ~x421 & ~x429 & ~x430 & ~x440 & ~x448 & ~x458 & ~x460 & ~x469 & ~x470 & ~x472 & ~x499 & ~x507 & ~x528 & ~x529 & ~x530 & ~x536 & ~x541 & ~x553 & ~x554 & ~x558 & ~x560 & ~x586 & ~x608 & ~x613 & ~x614 & ~x619 & ~x637 & ~x645 & ~x646 & ~x666 & ~x669 & ~x671 & ~x675 & ~x692 & ~x693 & ~x695 & ~x696 & ~x698 & ~x700 & ~x705 & ~x723 & ~x732 & ~x749 & ~x760 & ~x766 & ~x769;
assign c7299 =  x596 &  x601 & ~x94 & ~x199 & ~x310 & ~x747 & ~x754 & ~x782;
assign c80 = ~x26 & ~x60 & ~x72 & ~x105 & ~x117 & ~x136 & ~x165 & ~x216 & ~x266 & ~x385 & ~x402 & ~x426 & ~x447 & ~x478 & ~x484 & ~x498 & ~x501 & ~x527 & ~x581 & ~x596 & ~x653 & ~x664 & ~x669 & ~x675 & ~x711 & ~x726 & ~x742 & ~x772;
assign c82 =  x183 &  x288 &  x404 & ~x8 & ~x16 & ~x59 & ~x65 & ~x85 & ~x103 & ~x107 & ~x116 & ~x136 & ~x160 & ~x166 & ~x172 & ~x193 & ~x199 & ~x253 & ~x256 & ~x282 & ~x364 & ~x366 & ~x368 & ~x369 & ~x388 & ~x445 & ~x475 & ~x536 & ~x618 & ~x620 & ~x713 & ~x720 & ~x729 & ~x732 & ~x734 & ~x738 & ~x743 & ~x756 & ~x765 & ~x772 & ~x775;
assign c84 =  x270 &  x349 &  x629 & ~x85 & ~x97 & ~x222 & ~x268 & ~x593 & ~x594 & ~x678;
assign c86 =  x492 &  x629 & ~x149 & ~x150 & ~x438 & ~x546 & ~x623;
assign c88 =  x406 &  x486 &  x513 &  x626 & ~x543;
assign c810 =  x349 &  x628 & ~x39 & ~x63 & ~x74 & ~x142 & ~x192 & ~x346 & ~x374 & ~x416 & ~x483 & ~x559 & ~x565 & ~x623 & ~x666 & ~x734 & ~x755 & ~x756 & ~x762 & ~x783;
assign c812 =  x699;
assign c814 =  x113;
assign c816 =  x154 &  x179 &  x205 &  x287 &  x430 & ~x52 & ~x99 & ~x529;
assign c818 =  x379 &  x540 &  x623;
assign c820 =  x545 &  x578 &  x660 & ~x470 & ~x471;
assign c822 =  x301 &  x380 &  x458 & ~x5 & ~x8 & ~x15 & ~x16 & ~x28 & ~x41 & ~x69 & ~x74 & ~x83 & ~x87 & ~x88 & ~x96 & ~x98 & ~x117 & ~x120 & ~x121 & ~x148 & ~x149 & ~x163 & ~x173 & ~x194 & ~x198 & ~x200 & ~x224 & ~x250 & ~x253 & ~x255 & ~x310 & ~x362 & ~x387 & ~x394 & ~x415 & ~x425 & ~x443 & ~x444 & ~x452 & ~x453 & ~x472 & ~x502 & ~x528 & ~x530 & ~x533 & ~x557 & ~x559 & ~x562 & ~x564 & ~x612 & ~x615 & ~x641 & ~x646 & ~x697 & ~x699 & ~x729 & ~x760 & ~x766;
assign c824 =  x3;
assign c826 =  x476;
assign c828 =  x750;
assign c830 =  x404 &  x458 &  x485 &  x512 & ~x5 & ~x12 & ~x44 & ~x53 & ~x56 & ~x61 & ~x75 & ~x79 & ~x101 & ~x120 & ~x121 & ~x123 & ~x145 & ~x146 & ~x163 & ~x228 & ~x251 & ~x279 & ~x338 & ~x362 & ~x367 & ~x477 & ~x482 & ~x501 & ~x515 & ~x560 & ~x564 & ~x613 & ~x616 & ~x641 & ~x642 & ~x675 & ~x695 & ~x696 & ~x719 & ~x729 & ~x749 & ~x760 & ~x763 & ~x776;
assign c832 =  x328 &  x657 & ~x270 & ~x452;
assign c834 =  x279;
assign c836 =  x316 &  x404 &  x433 &  x490 &  x606 & ~x682;
assign c838 =  x180 & ~x8 & ~x45 & ~x169 & ~x256 & ~x293 & ~x313 & ~x334 & ~x482 & ~x513 & ~x539 & ~x553 & ~x585 & ~x589 & ~x596 & ~x612 & ~x653 & ~x711 & ~x768;
assign c840 =  x319 & ~x17 & ~x53 & ~x118 & ~x135 & ~x281 & ~x293 & ~x360 & ~x372 & ~x373 & ~x439 & ~x474 & ~x479 & ~x480 & ~x527 & ~x538 & ~x638 & ~x649 & ~x712 & ~x723 & ~x733;
assign c842 =  x514 & ~x6 & ~x20 & ~x34 & ~x119 & ~x152 & ~x179 & ~x308 & ~x427 & ~x508 & ~x538 & ~x704 & ~x742 & ~x757 & ~x778;
assign c844 =  x292 &  x349 & ~x1 & ~x72 & ~x138 & ~x193 & ~x199 & ~x346 & ~x365 & ~x525 & ~x575 & ~x591 & ~x619 & ~x675 & ~x708 & ~x728 & ~x739 & ~x745 & ~x763 & ~x764 & ~x775 & ~x777 & ~x783;
assign c846 = ~x25 & ~x28 & ~x29 & ~x68 & ~x75 & ~x164 & ~x174 & ~x179 & ~x201 & ~x206 & ~x219 & ~x220 & ~x228 & ~x239 & ~x248 & ~x278 & ~x281 & ~x288 & ~x311 & ~x364 & ~x393 & ~x398 & ~x399 & ~x426 & ~x427 & ~x448 & ~x466 & ~x467 & ~x475 & ~x480 & ~x482 & ~x531 & ~x536 & ~x539 & ~x552 & ~x595 & ~x607 & ~x610 & ~x614 & ~x623 & ~x651 & ~x652 & ~x665 & ~x672 & ~x700 & ~x704 & ~x708 & ~x710 & ~x717 & ~x739 & ~x743 & ~x746 & ~x768;
assign c848 =  x345 &  x375 &  x433 &  x461 & ~x19 & ~x20 & ~x47 & ~x54 & ~x77 & ~x89 & ~x97 & ~x159 & ~x169 & ~x365 & ~x391 & ~x399 & ~x428 & ~x565 & ~x705 & ~x708 & ~x761;
assign c850 =  x314 &  x372 &  x403 &  x433 & ~x426;
assign c852 =  x273 &  x353 & ~x23 & ~x25 & ~x47 & ~x172 & ~x256 & ~x387 & ~x410 & ~x416 & ~x425 & ~x555 & ~x615 & ~x640 & ~x649 & ~x679 & ~x758 & ~x770;
assign c854 =  x478;
assign c856 =  x617;
assign c858 =  x543 & ~x20 & ~x88 & ~x98 & ~x151 & ~x355 & ~x416 & ~x450 & ~x471 & ~x485 & ~x509 & ~x531 & ~x540 & ~x541 & ~x545 & ~x567 & ~x594 & ~x623 & ~x624 & ~x671 & ~x742 & ~x782;
assign c860 =  x449;
assign c862 =  x264 &  x353 & ~x315 & ~x385 & ~x437 & ~x495 & ~x633 & ~x739 & ~x755;
assign c864 =  x379 &  x403 &  x457 &  x512 &  x656 & ~x2 & ~x5 & ~x7 & ~x8 & ~x11 & ~x12 & ~x15 & ~x18 & ~x19 & ~x24 & ~x28 & ~x31 & ~x32 & ~x38 & ~x46 & ~x50 & ~x54 & ~x55 & ~x60 & ~x64 & ~x66 & ~x71 & ~x73 & ~x75 & ~x76 & ~x79 & ~x80 & ~x83 & ~x86 & ~x87 & ~x90 & ~x93 & ~x97 & ~x98 & ~x102 & ~x105 & ~x109 & ~x113 & ~x134 & ~x135 & ~x137 & ~x140 & ~x143 & ~x144 & ~x163 & ~x167 & ~x192 & ~x194 & ~x195 & ~x199 & ~x201 & ~x223 & ~x224 & ~x225 & ~x251 & ~x252 & ~x253 & ~x255 & ~x279 & ~x281 & ~x283 & ~x304 & ~x309 & ~x334 & ~x361 & ~x362 & ~x365 & ~x389 & ~x390 & ~x396 & ~x418 & ~x420 & ~x422 & ~x451 & ~x474 & ~x476 & ~x479 & ~x504 & ~x506 & ~x531 & ~x532 & ~x533 & ~x562 & ~x585 & ~x589 & ~x641 & ~x643 & ~x645 & ~x668 & ~x669 & ~x672 & ~x675 & ~x693 & ~x701 & ~x708 & ~x709 & ~x710 & ~x711 & ~x712 & ~x715 & ~x718 & ~x723 & ~x724 & ~x726 & ~x728 & ~x736 & ~x740 & ~x744 & ~x745 & ~x748 & ~x752 & ~x756 & ~x757 & ~x762 & ~x765 & ~x768 & ~x771 & ~x773 & ~x776 & ~x778 & ~x781 & ~x782;
assign c866 =  x304 &  x358;
assign c868 =  x291 &  x462 &  x516 &  x544 & ~x17 & ~x18 & ~x24 & ~x35 & ~x43 & ~x47 & ~x52 & ~x67 & ~x69 & ~x72 & ~x77 & ~x87 & ~x92 & ~x98 & ~x102 & ~x104 & ~x114 & ~x119 & ~x135 & ~x142 & ~x143 & ~x146 & ~x149 & ~x168 & ~x169 & ~x171 & ~x172 & ~x200 & ~x202 & ~x221 & ~x225 & ~x227 & ~x281 & ~x309 & ~x311 & ~x336 & ~x366 & ~x368 & ~x392 & ~x398 & ~x413 & ~x418 & ~x421 & ~x423 & ~x445 & ~x451 & ~x467 & ~x468 & ~x471 & ~x472 & ~x480 & ~x483 & ~x499 & ~x501 & ~x510 & ~x511 & ~x512 & ~x532 & ~x535 & ~x536 & ~x554 & ~x560 & ~x587 & ~x609 & ~x616 & ~x618 & ~x621 & ~x649 & ~x667 & ~x673 & ~x675 & ~x678 & ~x697 & ~x701 & ~x703 & ~x705 & ~x706 & ~x709 & ~x710 & ~x718 & ~x721 & ~x728 & ~x754 & ~x757 & ~x765 & ~x766 & ~x767 & ~x773 & ~x777;
assign c870 =  x351 &  x457 &  x484 & ~x8 & ~x10 & ~x16 & ~x18 & ~x21 & ~x24 & ~x31 & ~x32 & ~x35 & ~x40 & ~x41 & ~x43 & ~x45 & ~x50 & ~x51 & ~x52 & ~x58 & ~x62 & ~x66 & ~x68 & ~x71 & ~x79 & ~x93 & ~x102 & ~x103 & ~x104 & ~x106 & ~x112 & ~x117 & ~x118 & ~x120 & ~x140 & ~x144 & ~x165 & ~x167 & ~x171 & ~x173 & ~x223 & ~x255 & ~x280 & ~x283 & ~x306 & ~x310 & ~x366 & ~x368 & ~x390 & ~x396 & ~x397 & ~x420 & ~x479 & ~x488 & ~x505 & ~x531 & ~x557 & ~x560 & ~x577 & ~x584 & ~x586 & ~x588 & ~x619 & ~x640 & ~x641 & ~x642 & ~x646 & ~x666 & ~x667 & ~x673 & ~x674 & ~x676 & ~x678 & ~x694 & ~x695 & ~x697 & ~x704 & ~x711 & ~x719 & ~x721 & ~x723 & ~x740 & ~x741 & ~x742 & ~x750 & ~x752 & ~x754 & ~x759 & ~x761 & ~x763 & ~x765 & ~x771 & ~x781;
assign c872 =  x153 & ~x5 & ~x12 & ~x26 & ~x27 & ~x38 & ~x48 & ~x50 & ~x51 & ~x60 & ~x61 & ~x64 & ~x72 & ~x75 & ~x89 & ~x90 & ~x96 & ~x99 & ~x100 & ~x103 & ~x111 & ~x121 & ~x131 & ~x141 & ~x145 & ~x147 & ~x159 & ~x160 & ~x164 & ~x172 & ~x173 & ~x174 & ~x193 & ~x194 & ~x199 & ~x200 & ~x201 & ~x210 & ~x249 & ~x255 & ~x279 & ~x304 & ~x361 & ~x364 & ~x389 & ~x394 & ~x418 & ~x421 & ~x474 & ~x479 & ~x491 & ~x530 & ~x532 & ~x593 & ~x620 & ~x642 & ~x643 & ~x645 & ~x649 & ~x668 & ~x676 & ~x694 & ~x699 & ~x708 & ~x714 & ~x716 & ~x718 & ~x720 & ~x723 & ~x726 & ~x740 & ~x743 & ~x744 & ~x745 & ~x752 & ~x753 & ~x759 & ~x762 & ~x774 & ~x776 & ~x779;
assign c874 =  x158 &  x237 &  x435 & ~x241 & ~x539;
assign c876 =  x587;
assign c878 =  x542 &  x569 &  x682;
assign c880 =  x7;
assign c882 =  x317 &  x375 &  x405 &  x434 & ~x10 & ~x12 & ~x16 & ~x22 & ~x25 & ~x35 & ~x37 & ~x39 & ~x53 & ~x72 & ~x75 & ~x84 & ~x94 & ~x97 & ~x106 & ~x163 & ~x172 & ~x193 & ~x196 & ~x219 & ~x225 & ~x251 & ~x274 & ~x278 & ~x313 & ~x330 & ~x359 & ~x367 & ~x371 & ~x385 & ~x400 & ~x413 & ~x414 & ~x422 & ~x426 & ~x428 & ~x443 & ~x444 & ~x451 & ~x509 & ~x510 & ~x526 & ~x530 & ~x555 & ~x564 & ~x584 & ~x590 & ~x613 & ~x643 & ~x668 & ~x702 & ~x709 & ~x710 & ~x733 & ~x740 & ~x759 & ~x775 & ~x780;
assign c884 =  x287 &  x374 & ~x10 & ~x11 & ~x17 & ~x21 & ~x33 & ~x36 & ~x37 & ~x40 & ~x42 & ~x51 & ~x74 & ~x77 & ~x92 & ~x93 & ~x97 & ~x113 & ~x133 & ~x137 & ~x139 & ~x145 & ~x163 & ~x172 & ~x195 & ~x199 & ~x218 & ~x339 & ~x392 & ~x397 & ~x398 & ~x399 & ~x451 & ~x505 & ~x557 & ~x563 & ~x590 & ~x641 & ~x644 & ~x645 & ~x669 & ~x670 & ~x671 & ~x699 & ~x702 & ~x725 & ~x729 & ~x730 & ~x733 & ~x734 & ~x738 & ~x739 & ~x745 & ~x746 & ~x760 & ~x774 & ~x779;
assign c886 =  x392;
assign c888 =  x431 &  x458 &  x513 &  x597 &  x626 & ~x4 & ~x5 & ~x19 & ~x20 & ~x30 & ~x38 & ~x39 & ~x41 & ~x56 & ~x72 & ~x79 & ~x85 & ~x94 & ~x95 & ~x96 & ~x103 & ~x105 & ~x109 & ~x110 & ~x114 & ~x119 & ~x135 & ~x144 & ~x164 & ~x166 & ~x167 & ~x174 & ~x197 & ~x225 & ~x307 & ~x308 & ~x309 & ~x311 & ~x312 & ~x332 & ~x333 & ~x335 & ~x336 & ~x338 & ~x367 & ~x420 & ~x474 & ~x479 & ~x505 & ~x506 & ~x529 & ~x544 & ~x558 & ~x561 & ~x584 & ~x593 & ~x612 & ~x613 & ~x615 & ~x640 & ~x641 & ~x642 & ~x645 & ~x647 & ~x648 & ~x649 & ~x651 & ~x705 & ~x723 & ~x744 & ~x747 & ~x752 & ~x753 & ~x763 & ~x765 & ~x776 & ~x779 & ~x781;
assign c890 =  x378 &  x437 &  x466 &  x488 &  x516 & ~x1 & ~x5 & ~x13 & ~x25 & ~x30 & ~x45 & ~x49 & ~x81 & ~x169 & ~x170 & ~x225 & ~x305 & ~x414 & ~x457 & ~x504 & ~x508 & ~x589 & ~x612 & ~x700 & ~x733 & ~x737 & ~x754 & ~x765 & ~x773;
assign c892 =  x356 &  x407 & ~x1 & ~x24 & ~x69 & ~x73 & ~x103 & ~x139 & ~x200 & ~x223 & ~x229 & ~x282 & ~x340 & ~x452 & ~x504 & ~x507 & ~x520 & ~x547 & ~x558 & ~x664 & ~x698 & ~x705 & ~x733 & ~x740 & ~x769 & ~x782;
assign c894 =  x572 &  x600 &  x660 & ~x15 & ~x16 & ~x21 & ~x28 & ~x31 & ~x38 & ~x40 & ~x43 & ~x56 & ~x57 & ~x63 & ~x66 & ~x70 & ~x73 & ~x78 & ~x83 & ~x84 & ~x86 & ~x87 & ~x88 & ~x91 & ~x99 & ~x100 & ~x101 & ~x117 & ~x120 & ~x130 & ~x137 & ~x139 & ~x140 & ~x143 & ~x159 & ~x169 & ~x172 & ~x173 & ~x196 & ~x220 & ~x222 & ~x226 & ~x249 & ~x250 & ~x254 & ~x277 & ~x283 & ~x304 & ~x306 & ~x309 & ~x332 & ~x335 & ~x338 & ~x360 & ~x364 & ~x365 & ~x366 & ~x385 & ~x386 & ~x393 & ~x396 & ~x398 & ~x415 & ~x419 & ~x420 & ~x441 & ~x443 & ~x445 & ~x473 & ~x482 & ~x499 & ~x504 & ~x508 & ~x509 & ~x512 & ~x527 & ~x539 & ~x540 & ~x559 & ~x569 & ~x584 & ~x586 & ~x591 & ~x610 & ~x616 & ~x621 & ~x622 & ~x641 & ~x642 & ~x643 & ~x645 & ~x648 & ~x650 & ~x651 & ~x652 & ~x665 & ~x667 & ~x671 & ~x674 & ~x710 & ~x711 & ~x717 & ~x720 & ~x722 & ~x723 & ~x728 & ~x734 & ~x735 & ~x737 & ~x738 & ~x740 & ~x742 & ~x751 & ~x761 & ~x763 & ~x766 & ~x768 & ~x769 & ~x776;
assign c896 =  x263 &  x377 &  x659 & ~x197 & ~x237;
assign c898 =  x184 &  x489 &  x659 & ~x2 & ~x5 & ~x15 & ~x53 & ~x119 & ~x120 & ~x229 & ~x253 & ~x309 & ~x314 & ~x333 & ~x360 & ~x387 & ~x389 & ~x398 & ~x415 & ~x419 & ~x423 & ~x425 & ~x445 & ~x485 & ~x486 & ~x509 & ~x566 & ~x583 & ~x596 & ~x609 & ~x618 & ~x650 & ~x675 & ~x678 & ~x704 & ~x732 & ~x733 & ~x742 & ~x749 & ~x755 & ~x762 & ~x780;
assign c8100 =  x459 &  x595 & ~x0 & ~x7 & ~x8 & ~x14 & ~x15 & ~x20 & ~x22 & ~x26 & ~x27 & ~x34 & ~x37 & ~x44 & ~x48 & ~x50 & ~x52 & ~x55 & ~x56 & ~x63 & ~x64 & ~x68 & ~x73 & ~x76 & ~x85 & ~x86 & ~x88 & ~x89 & ~x91 & ~x96 & ~x99 & ~x101 & ~x102 & ~x105 & ~x108 & ~x112 & ~x113 & ~x118 & ~x120 & ~x121 & ~x122 & ~x123 & ~x138 & ~x139 & ~x145 & ~x146 & ~x147 & ~x173 & ~x195 & ~x200 & ~x203 & ~x230 & ~x257 & ~x279 & ~x287 & ~x334 & ~x336 & ~x339 & ~x343 & ~x365 & ~x390 & ~x420 & ~x421 & ~x425 & ~x446 & ~x447 & ~x450 & ~x451 & ~x452 & ~x475 & ~x497 & ~x499 & ~x505 & ~x507 & ~x508 & ~x525 & ~x526 & ~x534 & ~x535 & ~x536 & ~x551 & ~x558 & ~x561 & ~x579 & ~x580 & ~x581 & ~x584 & ~x585 & ~x589 & ~x590 & ~x606 & ~x609 & ~x615 & ~x617 & ~x632 & ~x634 & ~x635 & ~x636 & ~x638 & ~x663 & ~x668 & ~x672 & ~x673 & ~x687 & ~x703 & ~x715 & ~x718 & ~x734 & ~x749 & ~x758 & ~x764 & ~x769 & ~x771 & ~x772 & ~x774 & ~x776 & ~x779 & ~x781 & ~x782;
assign c8102 =  x658 & ~x0 & ~x10 & ~x18 & ~x23 & ~x25 & ~x31 & ~x32 & ~x36 & ~x39 & ~x53 & ~x56 & ~x58 & ~x65 & ~x71 & ~x73 & ~x75 & ~x84 & ~x99 & ~x115 & ~x134 & ~x142 & ~x163 & ~x174 & ~x190 & ~x192 & ~x194 & ~x226 & ~x251 & ~x254 & ~x304 & ~x307 & ~x313 & ~x314 & ~x334 & ~x335 & ~x439 & ~x474 & ~x480 & ~x496 & ~x498 & ~x504 & ~x525 & ~x558 & ~x582 & ~x602 & ~x646 & ~x671 & ~x675 & ~x678 & ~x699 & ~x705 & ~x706 & ~x710 & ~x714 & ~x718 & ~x722 & ~x729 & ~x740 & ~x743 & ~x745 & ~x757 & ~x758 & ~x762 & ~x765 & ~x766 & ~x769 & ~x770 & ~x774;
assign c8104 =  x541 &  x654 & ~x0 & ~x40 & ~x76 & ~x80 & ~x101 & ~x172 & ~x337 & ~x369 & ~x475 & ~x572 & ~x589 & ~x590 & ~x618 & ~x637;
assign c8106 =  x404 &  x433 &  x461 & ~x1 & ~x2 & ~x3 & ~x7 & ~x13 & ~x15 & ~x16 & ~x21 & ~x22 & ~x24 & ~x25 & ~x26 & ~x29 & ~x31 & ~x36 & ~x41 & ~x44 & ~x47 & ~x48 & ~x49 & ~x54 & ~x55 & ~x58 & ~x63 & ~x68 & ~x74 & ~x77 & ~x82 & ~x83 & ~x85 & ~x88 & ~x89 & ~x93 & ~x95 & ~x96 & ~x101 & ~x102 & ~x107 & ~x108 & ~x109 & ~x115 & ~x135 & ~x138 & ~x139 & ~x141 & ~x144 & ~x146 & ~x147 & ~x163 & ~x165 & ~x169 & ~x171 & ~x190 & ~x191 & ~x192 & ~x193 & ~x196 & ~x197 & ~x202 & ~x219 & ~x225 & ~x226 & ~x227 & ~x251 & ~x253 & ~x254 & ~x278 & ~x280 & ~x283 & ~x284 & ~x305 & ~x308 & ~x322 & ~x331 & ~x336 & ~x359 & ~x365 & ~x370 & ~x388 & ~x395 & ~x396 & ~x416 & ~x418 & ~x419 & ~x420 & ~x422 & ~x425 & ~x426 & ~x441 & ~x442 & ~x446 & ~x448 & ~x450 & ~x453 & ~x456 & ~x458 & ~x469 & ~x470 & ~x472 & ~x480 & ~x484 & ~x499 & ~x501 & ~x503 & ~x504 & ~x507 & ~x509 & ~x510 & ~x512 & ~x528 & ~x533 & ~x536 & ~x537 & ~x539 & ~x540 & ~x556 & ~x557 & ~x559 & ~x582 & ~x583 & ~x586 & ~x587 & ~x589 & ~x591 & ~x594 & ~x612 & ~x613 & ~x614 & ~x620 & ~x622 & ~x640 & ~x642 & ~x645 & ~x646 & ~x647 & ~x648 & ~x649 & ~x650 & ~x668 & ~x674 & ~x675 & ~x677 & ~x679 & ~x698 & ~x702 & ~x708 & ~x723 & ~x733 & ~x734 & ~x741 & ~x744 & ~x752 & ~x756 & ~x757 & ~x758 & ~x760 & ~x762 & ~x763 & ~x766 & ~x767 & ~x770 & ~x771 & ~x773 & ~x781 & ~x783;
assign c8108 =  x289 &  x376 & ~x4 & ~x6 & ~x20 & ~x75 & ~x83 & ~x90 & ~x95 & ~x98 & ~x102 & ~x111 & ~x134 & ~x164 & ~x189 & ~x193 & ~x194 & ~x257 & ~x315 & ~x334 & ~x368 & ~x394 & ~x400 & ~x451 & ~x477 & ~x509 & ~x528 & ~x534 & ~x559 & ~x619 & ~x672 & ~x680 & ~x681 & ~x691 & ~x699 & ~x701 & ~x713 & ~x721 & ~x727 & ~x733 & ~x750 & ~x756 & ~x780;
assign c8110 =  x324 &  x434 & ~x66 & ~x117 & ~x329 & ~x365 & ~x408 & ~x409 & ~x410 & ~x411 & ~x439 & ~x441 & ~x499 & ~x589 & ~x624 & ~x625 & ~x679 & ~x709;
assign c8112 =  x461 &  x515 &  x542 & ~x324 & ~x484 & ~x509 & ~x523;
assign c8114 =  x348 &  x405 & ~x34 & ~x37 & ~x55 & ~x63 & ~x123 & ~x137 & ~x169 & ~x195 & ~x252 & ~x257 & ~x266 & ~x374 & ~x399 & ~x443 & ~x536 & ~x564 & ~x611 & ~x646 & ~x666 & ~x718;
assign c8116 =  x303 &  x408 &  x486;
assign c8118 =  x353 &  x376 &  x377 &  x430 &  x457 &  x484 &  x626 & ~x4 & ~x6 & ~x11 & ~x15 & ~x16 & ~x17 & ~x18 & ~x23 & ~x32 & ~x33 & ~x34 & ~x35 & ~x39 & ~x45 & ~x52 & ~x53 & ~x54 & ~x56 & ~x58 & ~x59 & ~x61 & ~x62 & ~x73 & ~x75 & ~x81 & ~x84 & ~x87 & ~x93 & ~x97 & ~x101 & ~x103 & ~x104 & ~x105 & ~x106 & ~x107 & ~x108 & ~x110 & ~x113 & ~x114 & ~x137 & ~x139 & ~x171 & ~x196 & ~x199 & ~x250 & ~x252 & ~x253 & ~x255 & ~x277 & ~x278 & ~x309 & ~x310 & ~x311 & ~x332 & ~x337 & ~x338 & ~x340 & ~x361 & ~x368 & ~x386 & ~x389 & ~x395 & ~x398 & ~x399 & ~x415 & ~x419 & ~x423 & ~x424 & ~x425 & ~x443 & ~x444 & ~x445 & ~x448 & ~x451 & ~x452 & ~x473 & ~x502 & ~x529 & ~x533 & ~x556 & ~x558 & ~x563 & ~x585 & ~x586 & ~x587 & ~x589 & ~x591 & ~x615 & ~x645 & ~x646 & ~x667 & ~x670 & ~x671 & ~x673 & ~x674 & ~x676 & ~x694 & ~x700 & ~x704 & ~x709 & ~x712 & ~x713 & ~x715 & ~x717 & ~x719 & ~x722 & ~x724 & ~x725 & ~x729 & ~x730 & ~x733 & ~x738 & ~x743 & ~x748 & ~x753 & ~x754 & ~x756 & ~x758 & ~x764 & ~x767 & ~x774 & ~x779 & ~x780;
assign c8120 =  x431 &  x663;
assign c8122 =  x355 &  x403 &  x656 &  x657 & ~x453 & ~x547 & ~x548;
assign c8124 =  x355 &  x381 & ~x23 & ~x29 & ~x39 & ~x41 & ~x46 & ~x60 & ~x61 & ~x77 & ~x80 & ~x84 & ~x86 & ~x93 & ~x102 & ~x105 & ~x114 & ~x123 & ~x124 & ~x148 & ~x176 & ~x279 & ~x298 & ~x334 & ~x392 & ~x398 & ~x444 & ~x448 & ~x452 & ~x501 & ~x502 & ~x508 & ~x529 & ~x556 & ~x557 & ~x559 & ~x589 & ~x615 & ~x619 & ~x639 & ~x646 & ~x648 & ~x666 & ~x674 & ~x696 & ~x707 & ~x735 & ~x736 & ~x739 & ~x745 & ~x760;
assign c8126 =  x344 &  x460 &  x544 &  x660 & ~x618;
assign c8128 =  x462 &  x515 & ~x39 & ~x46 & ~x54 & ~x59 & ~x61 & ~x64 & ~x86 & ~x91 & ~x93 & ~x113 & ~x139 & ~x142 & ~x285 & ~x337 & ~x425 & ~x427 & ~x445 & ~x456 & ~x469 & ~x479 & ~x481 & ~x494 & ~x495 & ~x499 & ~x509 & ~x532 & ~x535 & ~x537 & ~x551 & ~x557 & ~x578 & ~x585 & ~x588 & ~x619 & ~x634 & ~x638 & ~x645 & ~x661 & ~x664 & ~x666 & ~x667 & ~x670 & ~x706 & ~x707 & ~x722 & ~x731 & ~x750 & ~x762 & ~x769 & ~x775;
assign c8130 =  x291 &  x320 &  x349 & ~x6 & ~x11 & ~x35 & ~x49 & ~x62 & ~x68 & ~x69 & ~x72 & ~x73 & ~x74 & ~x79 & ~x83 & ~x85 & ~x87 & ~x102 & ~x106 & ~x117 & ~x118 & ~x119 & ~x133 & ~x134 & ~x136 & ~x140 & ~x144 & ~x163 & ~x172 & ~x197 & ~x198 & ~x222 & ~x227 & ~x254 & ~x284 & ~x344 & ~x345 & ~x358 & ~x359 & ~x361 & ~x362 & ~x384 & ~x389 & ~x390 & ~x391 & ~x392 & ~x399 & ~x413 & ~x420 & ~x423 & ~x425 & ~x475 & ~x500 & ~x502 & ~x532 & ~x559 & ~x589 & ~x615 & ~x622 & ~x644 & ~x680 & ~x692 & ~x694 & ~x695 & ~x698 & ~x702 & ~x705 & ~x710 & ~x719 & ~x721 & ~x724 & ~x733 & ~x734 & ~x742 & ~x744 & ~x745 & ~x753 & ~x769 & ~x776;
assign c8132 =  x516 &  x543 &  x685 & ~x32 & ~x43 & ~x46 & ~x63 & ~x74 & ~x85 & ~x89 & ~x92 & ~x132 & ~x140 & ~x144 & ~x200 & ~x227 & ~x252 & ~x530 & ~x533 & ~x557 & ~x561 & ~x648 & ~x670 & ~x678 & ~x703 & ~x726 & ~x739;
assign c8134 = ~x2 & ~x13 & ~x14 & ~x17 & ~x27 & ~x29 & ~x30 & ~x38 & ~x48 & ~x50 & ~x61 & ~x65 & ~x68 & ~x73 & ~x80 & ~x85 & ~x106 & ~x117 & ~x131 & ~x133 & ~x141 & ~x143 & ~x148 & ~x160 & ~x166 & ~x172 & ~x173 & ~x190 & ~x191 & ~x199 & ~x223 & ~x225 & ~x226 & ~x228 & ~x250 & ~x254 & ~x282 & ~x306 & ~x336 & ~x362 & ~x389 & ~x398 & ~x400 & ~x419 & ~x422 & ~x423 & ~x440 & ~x449 & ~x453 & ~x469 & ~x481 & ~x482 & ~x502 & ~x507 & ~x532 & ~x535 & ~x558 & ~x560 & ~x566 & ~x573 & ~x581 & ~x616 & ~x617 & ~x618 & ~x624 & ~x625 & ~x647 & ~x652 & ~x677 & ~x681 & ~x694 & ~x697 & ~x702 & ~x709 & ~x717 & ~x725 & ~x733 & ~x742 & ~x744 & ~x749 & ~x759 & ~x766 & ~x767 & ~x768 & ~x769 & ~x774 & ~x780 & ~x782;
assign c8136 =  x261 &  x318 &  x348 & ~x14 & ~x29 & ~x31 & ~x55 & ~x63 & ~x84 & ~x98 & ~x112 & ~x114 & ~x119 & ~x168 & ~x198 & ~x312 & ~x335 & ~x338 & ~x372 & ~x471 & ~x584 & ~x611 & ~x613 & ~x642 & ~x644 & ~x645 & ~x648 & ~x649 & ~x680 & ~x708 & ~x711 & ~x713 & ~x720 & ~x723 & ~x726 & ~x727 & ~x730 & ~x733 & ~x735 & ~x743 & ~x750 & ~x772 & ~x775 & ~x777;
assign c8138 =  x299 &  x408 &  x656 &  x657 & ~x3 & ~x9 & ~x15 & ~x23 & ~x24 & ~x30 & ~x32 & ~x39 & ~x46 & ~x52 & ~x56 & ~x58 & ~x59 & ~x61 & ~x63 & ~x71 & ~x78 & ~x83 & ~x95 & ~x100 & ~x101 & ~x103 & ~x105 & ~x112 & ~x114 & ~x133 & ~x137 & ~x144 & ~x145 & ~x165 & ~x168 & ~x169 & ~x170 & ~x171 & ~x172 & ~x173 & ~x175 & ~x176 & ~x199 & ~x201 & ~x202 & ~x226 & ~x229 & ~x256 & ~x276 & ~x278 & ~x284 & ~x305 & ~x306 & ~x310 & ~x335 & ~x340 & ~x361 & ~x364 & ~x365 & ~x367 & ~x368 & ~x390 & ~x394 & ~x396 & ~x397 & ~x417 & ~x419 & ~x422 & ~x446 & ~x450 & ~x452 & ~x453 & ~x477 & ~x479 & ~x481 & ~x502 & ~x505 & ~x506 & ~x509 & ~x529 & ~x530 & ~x531 & ~x532 & ~x537 & ~x559 & ~x562 & ~x586 & ~x587 & ~x588 & ~x593 & ~x611 & ~x612 & ~x619 & ~x621 & ~x622 & ~x638 & ~x641 & ~x646 & ~x648 & ~x667 & ~x671 & ~x675 & ~x676 & ~x677 & ~x679 & ~x696 & ~x699 & ~x704 & ~x706 & ~x712 & ~x714 & ~x721 & ~x733 & ~x739 & ~x742 & ~x744 & ~x746 & ~x755 & ~x757 & ~x759 & ~x772 & ~x774 & ~x776 & ~x780 & ~x782 & ~x783;
assign c8140 =  x116;
assign c8142 =  x540 &  x568 & ~x29 & ~x71 & ~x78 & ~x81 & ~x97 & ~x99 & ~x142 & ~x308 & ~x309 & ~x333 & ~x364 & ~x426 & ~x507 & ~x509 & ~x562 & ~x563 & ~x570 & ~x583 & ~x665 & ~x668 & ~x699 & ~x701 & ~x727 & ~x731 & ~x780;
assign c8144 =  x43;
assign c8146 =  x332;
assign c8148 =  x279;
assign c8150 =  x152 &  x402 &  x403 & ~x549 & ~x687;
assign c8152 =  x10;
assign c8154 =  x265 &  x407 &  x460 &  x487 &  x569 & ~x30 & ~x33 & ~x148 & ~x205 & ~x418 & ~x428 & ~x429 & ~x448 & ~x450 & ~x482 & ~x497 & ~x606 & ~x607 & ~x615 & ~x676 & ~x777;
assign c8156 =  x464 &  x572 &  x631 &  x658 & ~x1 & ~x3 & ~x5 & ~x7 & ~x8 & ~x10 & ~x12 & ~x21 & ~x27 & ~x30 & ~x33 & ~x47 & ~x49 & ~x52 & ~x53 & ~x55 & ~x61 & ~x66 & ~x67 & ~x68 & ~x70 & ~x72 & ~x79 & ~x82 & ~x90 & ~x91 & ~x94 & ~x98 & ~x101 & ~x111 & ~x118 & ~x119 & ~x122 & ~x140 & ~x141 & ~x142 & ~x150 & ~x168 & ~x169 & ~x176 & ~x177 & ~x194 & ~x195 & ~x197 & ~x200 & ~x220 & ~x222 & ~x250 & ~x252 & ~x253 & ~x255 & ~x277 & ~x281 & ~x306 & ~x311 & ~x333 & ~x334 & ~x337 & ~x388 & ~x395 & ~x419 & ~x421 & ~x422 & ~x425 & ~x439 & ~x440 & ~x447 & ~x469 & ~x470 & ~x473 & ~x476 & ~x478 & ~x482 & ~x483 & ~x498 & ~x500 & ~x508 & ~x510 & ~x511 & ~x529 & ~x538 & ~x539 & ~x558 & ~x559 & ~x562 & ~x566 & ~x569 & ~x582 & ~x586 & ~x590 & ~x592 & ~x595 & ~x597 & ~x611 & ~x614 & ~x616 & ~x617 & ~x639 & ~x642 & ~x647 & ~x651 & ~x670 & ~x672 & ~x680 & ~x690 & ~x692 & ~x698 & ~x699 & ~x701 & ~x706 & ~x707 & ~x716 & ~x717 & ~x721 & ~x726 & ~x732 & ~x734 & ~x736 & ~x737 & ~x743 & ~x745 & ~x751 & ~x752 & ~x754 & ~x756 & ~x758 & ~x760 & ~x761 & ~x771 & ~x772 & ~x781 & ~x782 & ~x783;
assign c8158 =  x695;
assign c8160 =  x461 &  x516 & ~x0 & ~x6 & ~x11 & ~x17 & ~x19 & ~x21 & ~x23 & ~x43 & ~x46 & ~x47 & ~x48 & ~x49 & ~x52 & ~x57 & ~x67 & ~x74 & ~x76 & ~x80 & ~x81 & ~x87 & ~x88 & ~x91 & ~x94 & ~x98 & ~x106 & ~x112 & ~x115 & ~x121 & ~x134 & ~x140 & ~x143 & ~x165 & ~x166 & ~x167 & ~x169 & ~x192 & ~x194 & ~x198 & ~x221 & ~x224 & ~x251 & ~x252 & ~x253 & ~x257 & ~x280 & ~x282 & ~x294 & ~x305 & ~x306 & ~x331 & ~x335 & ~x336 & ~x339 & ~x360 & ~x361 & ~x366 & ~x388 & ~x395 & ~x396 & ~x397 & ~x417 & ~x425 & ~x448 & ~x449 & ~x452 & ~x455 & ~x456 & ~x470 & ~x474 & ~x475 & ~x482 & ~x484 & ~x485 & ~x501 & ~x504 & ~x508 & ~x511 & ~x513 & ~x528 & ~x529 & ~x531 & ~x533 & ~x535 & ~x539 & ~x555 & ~x561 & ~x565 & ~x566 & ~x568 & ~x583 & ~x584 & ~x585 & ~x586 & ~x588 & ~x590 & ~x591 & ~x595 & ~x609 & ~x610 & ~x614 & ~x615 & ~x616 & ~x618 & ~x620 & ~x636 & ~x637 & ~x638 & ~x643 & ~x645 & ~x647 & ~x648 & ~x663 & ~x665 & ~x667 & ~x669 & ~x671 & ~x672 & ~x673 & ~x675 & ~x694 & ~x700 & ~x706 & ~x707 & ~x709 & ~x719 & ~x720 & ~x721 & ~x724 & ~x726 & ~x728 & ~x734 & ~x735 & ~x736 & ~x737 & ~x742 & ~x743 & ~x747 & ~x753 & ~x759 & ~x761 & ~x769 & ~x770 & ~x773 & ~x774 & ~x778 & ~x781 & ~x782 & ~x783;
assign c8162 =  x214 &  x264 &  x292 &  x405 & ~x17 & ~x35 & ~x71 & ~x78 & ~x105 & ~x117 & ~x122 & ~x134 & ~x171 & ~x226 & ~x282 & ~x312 & ~x337 & ~x366 & ~x372 & ~x374 & ~x427 & ~x447 & ~x472 & ~x477 & ~x504 & ~x507 & ~x552 & ~x556 & ~x559 & ~x620 & ~x640 & ~x664 & ~x675 & ~x692 & ~x693 & ~x696 & ~x757 & ~x758 & ~x766 & ~x778;
assign c8164 =  x542 & ~x0 & ~x9 & ~x17 & ~x25 & ~x27 & ~x28 & ~x31 & ~x35 & ~x38 & ~x41 & ~x45 & ~x51 & ~x52 & ~x55 & ~x57 & ~x58 & ~x63 & ~x65 & ~x68 & ~x69 & ~x70 & ~x71 & ~x74 & ~x78 & ~x82 & ~x83 & ~x87 & ~x88 & ~x90 & ~x99 & ~x108 & ~x109 & ~x112 & ~x114 & ~x117 & ~x125 & ~x134 & ~x138 & ~x139 & ~x164 & ~x170 & ~x171 & ~x173 & ~x201 & ~x223 & ~x224 & ~x225 & ~x226 & ~x248 & ~x278 & ~x282 & ~x308 & ~x311 & ~x331 & ~x340 & ~x357 & ~x362 & ~x365 & ~x366 & ~x387 & ~x388 & ~x395 & ~x412 & ~x420 & ~x439 & ~x442 & ~x443 & ~x444 & ~x456 & ~x469 & ~x478 & ~x480 & ~x497 & ~x498 & ~x501 & ~x507 & ~x509 & ~x527 & ~x534 & ~x536 & ~x558 & ~x561 & ~x572 & ~x585 & ~x586 & ~x592 & ~x594 & ~x611 & ~x612 & ~x615 & ~x620 & ~x639 & ~x642 & ~x643 & ~x645 & ~x646 & ~x649 & ~x650 & ~x669 & ~x670 & ~x671 & ~x675 & ~x678 & ~x692 & ~x697 & ~x702 & ~x705 & ~x706 & ~x717 & ~x719 & ~x720 & ~x722 & ~x725 & ~x728 & ~x732 & ~x733 & ~x737 & ~x738 & ~x741 & ~x743 & ~x746 & ~x750 & ~x753 & ~x761 & ~x769 & ~x771 & ~x774 & ~x775 & ~x777 & ~x782;
assign c8166 =  x185 &  x654 & ~x152 & ~x204 & ~x258 & ~x268 & ~x467 & ~x468 & ~x523 & ~x533 & ~x620 & ~x632;
assign c8168 =  x577 & ~x1 & ~x3 & ~x5 & ~x6 & ~x7 & ~x20 & ~x22 & ~x27 & ~x28 & ~x33 & ~x36 & ~x40 & ~x43 & ~x45 & ~x51 & ~x65 & ~x69 & ~x79 & ~x83 & ~x84 & ~x86 & ~x89 & ~x97 & ~x99 & ~x104 & ~x106 & ~x111 & ~x113 & ~x117 & ~x131 & ~x163 & ~x164 & ~x167 & ~x170 & ~x191 & ~x200 & ~x220 & ~x225 & ~x229 & ~x248 & ~x249 & ~x255 & ~x274 & ~x281 & ~x284 & ~x307 & ~x337 & ~x338 & ~x362 & ~x366 & ~x394 & ~x396 & ~x413 & ~x416 & ~x426 & ~x430 & ~x441 & ~x448 & ~x484 & ~x498 & ~x508 & ~x513 & ~x525 & ~x527 & ~x530 & ~x531 & ~x533 & ~x534 & ~x535 & ~x536 & ~x537 & ~x539 & ~x558 & ~x560 & ~x563 & ~x589 & ~x591 & ~x607 & ~x613 & ~x636 & ~x648 & ~x650 & ~x651 & ~x652 & ~x663 & ~x678 & ~x698 & ~x699 & ~x705 & ~x707 & ~x709 & ~x718 & ~x725 & ~x732 & ~x736 & ~x742 & ~x745 & ~x746 & ~x748 & ~x758 & ~x763 & ~x765 & ~x771 & ~x773 & ~x774 & ~x776;
assign c8170 =  x726;
assign c8172 =  x380 &  x434 & ~x3 & ~x7 & ~x9 & ~x11 & ~x13 & ~x22 & ~x25 & ~x33 & ~x34 & ~x36 & ~x44 & ~x47 & ~x53 & ~x54 & ~x57 & ~x62 & ~x63 & ~x66 & ~x68 & ~x78 & ~x79 & ~x85 & ~x95 & ~x96 & ~x97 & ~x98 & ~x111 & ~x115 & ~x119 & ~x121 & ~x122 & ~x137 & ~x150 & ~x171 & ~x172 & ~x173 & ~x194 & ~x197 & ~x202 & ~x204 & ~x223 & ~x224 & ~x231 & ~x252 & ~x277 & ~x280 & ~x282 & ~x283 & ~x296 & ~x340 & ~x342 & ~x360 & ~x363 & ~x365 & ~x370 & ~x385 & ~x392 & ~x414 & ~x415 & ~x420 & ~x422 & ~x440 & ~x450 & ~x452 & ~x453 & ~x467 & ~x474 & ~x495 & ~x497 & ~x498 & ~x502 & ~x507 & ~x525 & ~x531 & ~x536 & ~x551 & ~x559 & ~x582 & ~x586 & ~x587 & ~x591 & ~x608 & ~x609 & ~x610 & ~x638 & ~x640 & ~x648 & ~x663 & ~x676 & ~x678 & ~x680 & ~x692 & ~x694 & ~x698 & ~x701 & ~x704 & ~x709 & ~x712 & ~x713 & ~x725 & ~x729 & ~x730 & ~x732 & ~x733 & ~x739 & ~x756 & ~x759 & ~x762 & ~x763 & ~x765 & ~x769 & ~x770 & ~x771 & ~x776 & ~x779;
assign c8174 =  x13;
assign c8176 =  x317 &  x403 &  x432 &  x514 &  x570 & ~x30 & ~x50 & ~x98 & ~x100 & ~x529 & ~x612 & ~x744 & ~x783;
assign c8178 =  x392;
assign c8180 =  x317 &  x433 &  x489 & ~x7 & ~x24 & ~x75 & ~x76 & ~x116 & ~x123 & ~x278 & ~x368 & ~x385 & ~x387 & ~x415 & ~x416 & ~x418 & ~x425 & ~x428 & ~x454 & ~x456 & ~x474 & ~x478 & ~x483 & ~x507 & ~x509 & ~x513 & ~x529 & ~x539 & ~x640 & ~x675 & ~x698 & ~x708 & ~x724 & ~x726 & ~x738 & ~x748 & ~x757 & ~x778;
assign c8182 =  x392;
assign c8184 =  x345 &  x404 & ~x43 & ~x146 & ~x171 & ~x339 & ~x391 & ~x428 & ~x568 & ~x617 & ~x621 & ~x624 & ~x675 & ~x680 & ~x682 & ~x745;
assign c8186 =  x350 &  x658 & ~x51 & ~x61 & ~x105 & ~x108 & ~x229 & ~x373 & ~x385 & ~x387 & ~x394 & ~x510 & ~x565 & ~x568 & ~x574 & ~x595 & ~x644 & ~x651 & ~x728 & ~x744;
assign c8188 =  x316 &  x346 &  x376 & ~x265;
assign c8190 =  x436 &  x460 & ~x38 & ~x87 & ~x96 & ~x353 & ~x444 & ~x479 & ~x521 & ~x549 & ~x557 & ~x759;
assign c8192 =  x350 &  x353 &  x378 & ~x15 & ~x21 & ~x25 & ~x32 & ~x34 & ~x44 & ~x53 & ~x59 & ~x60 & ~x69 & ~x76 & ~x80 & ~x91 & ~x104 & ~x105 & ~x119 & ~x122 & ~x139 & ~x140 & ~x141 & ~x142 & ~x171 & ~x202 & ~x228 & ~x286 & ~x309 & ~x314 & ~x335 & ~x336 & ~x340 & ~x365 & ~x373 & ~x374 & ~x386 & ~x397 & ~x442 & ~x449 & ~x450 & ~x470 & ~x472 & ~x478 & ~x479 & ~x528 & ~x531 & ~x554 & ~x555 & ~x559 & ~x563 & ~x583 & ~x608 & ~x619 & ~x620 & ~x633 & ~x635 & ~x636 & ~x637 & ~x642 & ~x645 & ~x646 & ~x663 & ~x665 & ~x677 & ~x678 & ~x679 & ~x689 & ~x702 & ~x709 & ~x716 & ~x730 & ~x736 & ~x745 & ~x746 & ~x755 & ~x764 & ~x766 & ~x778 & ~x781;
assign c8194 =  x262 &  x291 &  x320 &  x349 &  x379 & ~x9 & ~x16 & ~x22 & ~x23 & ~x27 & ~x30 & ~x32 & ~x64 & ~x72 & ~x73 & ~x82 & ~x83 & ~x90 & ~x98 & ~x117 & ~x135 & ~x142 & ~x143 & ~x144 & ~x255 & ~x256 & ~x278 & ~x305 & ~x316 & ~x339 & ~x345 & ~x363 & ~x373 & ~x389 & ~x390 & ~x398 & ~x400 & ~x415 & ~x426 & ~x445 & ~x449 & ~x471 & ~x475 & ~x500 & ~x506 & ~x528 & ~x529 & ~x558 & ~x587 & ~x590 & ~x591 & ~x616 & ~x641 & ~x642 & ~x644 & ~x648 & ~x668 & ~x670 & ~x671 & ~x678 & ~x697 & ~x706 & ~x708 & ~x718 & ~x723 & ~x726 & ~x743 & ~x744 & ~x748 & ~x753 & ~x757 & ~x761 & ~x762 & ~x770 & ~x776 & ~x778;
assign c8196 = ~x4 & ~x10 & ~x23 & ~x24 & ~x28 & ~x35 & ~x38 & ~x48 & ~x67 & ~x70 & ~x80 & ~x82 & ~x88 & ~x94 & ~x96 & ~x100 & ~x102 & ~x118 & ~x120 & ~x131 & ~x138 & ~x139 & ~x196 & ~x199 & ~x218 & ~x220 & ~x227 & ~x229 & ~x231 & ~x331 & ~x355 & ~x363 & ~x374 & ~x390 & ~x395 & ~x396 & ~x414 & ~x415 & ~x421 & ~x426 & ~x447 & ~x448 & ~x450 & ~x452 & ~x453 & ~x469 & ~x473 & ~x479 & ~x504 & ~x512 & ~x534 & ~x546 & ~x555 & ~x557 & ~x562 & ~x587 & ~x617 & ~x618 & ~x623 & ~x639 & ~x642 & ~x668 & ~x690 & ~x693 & ~x696 & ~x697 & ~x702 & ~x706 & ~x712 & ~x725 & ~x729 & ~x733 & ~x745 & ~x751 & ~x753 & ~x762 & ~x768 & ~x770 & ~x772 & ~x774 & ~x779;
assign c8198 =  x180 &  x181 &  x314 &  x432 & ~x31 & ~x44 & ~x114 & ~x747 & ~x759;
assign c8200 =  x317 & ~x1 & ~x12 & ~x16 & ~x30 & ~x32 & ~x33 & ~x36 & ~x38 & ~x43 & ~x44 & ~x46 & ~x54 & ~x67 & ~x68 & ~x70 & ~x79 & ~x81 & ~x82 & ~x84 & ~x86 & ~x87 & ~x88 & ~x92 & ~x94 & ~x96 & ~x97 & ~x106 & ~x108 & ~x109 & ~x112 & ~x113 & ~x115 & ~x116 & ~x119 & ~x138 & ~x161 & ~x166 & ~x167 & ~x169 & ~x199 & ~x221 & ~x225 & ~x252 & ~x256 & ~x278 & ~x281 & ~x291 & ~x334 & ~x335 & ~x362 & ~x365 & ~x367 & ~x398 & ~x399 & ~x400 & ~x420 & ~x421 & ~x473 & ~x474 & ~x477 & ~x479 & ~x510 & ~x529 & ~x530 & ~x535 & ~x561 & ~x564 & ~x588 & ~x589 & ~x612 & ~x616 & ~x619 & ~x647 & ~x674 & ~x676 & ~x679 & ~x698 & ~x701 & ~x702 & ~x703 & ~x722 & ~x723 & ~x725 & ~x731 & ~x732 & ~x734 & ~x741 & ~x744 & ~x746 & ~x748 & ~x749 & ~x750 & ~x754 & ~x758 & ~x760 & ~x761 & ~x766 & ~x770 & ~x772 & ~x773 & ~x774 & ~x780;
assign c8202 =  x28;
assign c8204 =  x308;
assign c8206 =  x514 &  x542 &  x655 & ~x71 & ~x87 & ~x96 & ~x223 & ~x337 & ~x338 & ~x511 & ~x535 & ~x600 & ~x718 & ~x722 & ~x768;
assign c8208 =  x406 &  x515 &  x547 & ~x457 & ~x545;
assign c8210 =  x517 &  x544 &  x657 & ~x11 & ~x26 & ~x27 & ~x30 & ~x39 & ~x111 & ~x121 & ~x124 & ~x203 & ~x255 & ~x256 & ~x294 & ~x306 & ~x308 & ~x369 & ~x441 & ~x447 & ~x484 & ~x485 & ~x501 & ~x525 & ~x559 & ~x580 & ~x585 & ~x593 & ~x636 & ~x668 & ~x703;
assign c8212 =  x515 &  x570 & ~x19 & ~x30 & ~x40 & ~x42 & ~x44 & ~x55 & ~x99 & ~x114 & ~x129 & ~x134 & ~x140 & ~x141 & ~x144 & ~x146 & ~x283 & ~x362 & ~x417 & ~x423 & ~x471 & ~x528 & ~x529 & ~x531 & ~x545 & ~x554 & ~x555 & ~x585 & ~x611 & ~x635 & ~x636 & ~x645 & ~x650 & ~x676 & ~x689 & ~x693 & ~x705 & ~x730 & ~x742 & ~x744 & ~x772;
assign c8214 =  x47;
assign c8216 =  x377 &  x404 &  x512 & ~x14 & ~x18 & ~x23 & ~x47 & ~x48 & ~x53 & ~x66 & ~x69 & ~x74 & ~x75 & ~x82 & ~x92 & ~x94 & ~x109 & ~x113 & ~x121 & ~x134 & ~x137 & ~x141 & ~x168 & ~x196 & ~x221 & ~x229 & ~x335 & ~x342 & ~x395 & ~x446 & ~x504 & ~x505 & ~x528 & ~x533 & ~x542 & ~x560 & ~x587 & ~x589 & ~x590 & ~x610 & ~x615 & ~x647 & ~x668 & ~x719 & ~x720 & ~x721 & ~x747 & ~x748 & ~x780;
assign c8218 =  x434 &  x486 &  x540 &  x653 & ~x65 & ~x75 & ~x203 & ~x279 & ~x363 & ~x388 & ~x479 & ~x502 & ~x508 & ~x559 & ~x563 & ~x586 & ~x587 & ~x613 & ~x721 & ~x767 & ~x774 & ~x781;
assign c8220 =  x76;
assign c8222 =  x321 &  x350 &  x379 &  x406 & ~x1 & ~x3 & ~x20 & ~x28 & ~x29 & ~x32 & ~x40 & ~x45 & ~x54 & ~x58 & ~x73 & ~x81 & ~x95 & ~x100 & ~x110 & ~x145 & ~x239 & ~x310 & ~x366 & ~x391 & ~x453 & ~x528 & ~x555 & ~x557 & ~x562 & ~x583 & ~x613 & ~x707 & ~x712 & ~x719 & ~x723 & ~x728 & ~x732 & ~x737 & ~x750 & ~x751 & ~x773;
assign c8224 =  x364;
assign c8226 =  x302 &  x380 &  x407 & ~x464;
assign c8228 =  x655 & ~x3 & ~x23 & ~x29 & ~x30 & ~x45 & ~x50 & ~x54 & ~x69 & ~x72 & ~x80 & ~x81 & ~x82 & ~x86 & ~x87 & ~x98 & ~x120 & ~x136 & ~x147 & ~x168 & ~x174 & ~x277 & ~x278 & ~x280 & ~x281 & ~x305 & ~x339 & ~x367 & ~x389 & ~x391 & ~x395 & ~x445 & ~x448 & ~x451 & ~x521 & ~x522 & ~x531 & ~x561 & ~x563 & ~x572 & ~x591 & ~x613 & ~x620 & ~x640 & ~x641 & ~x691 & ~x699 & ~x702 & ~x713 & ~x715 & ~x734 & ~x739 & ~x774 & ~x779;
assign c8230 =  x531;
assign c8232 =  x463 &  x633 & ~x19 & ~x29 & ~x57 & ~x105 & ~x254 & ~x292 & ~x309 & ~x508 & ~x538 & ~x592 & ~x614 & ~x684 & ~x718 & ~x742;
assign c8234 =  x489 &  x660 & ~x1 & ~x3 & ~x10 & ~x17 & ~x20 & ~x26 & ~x27 & ~x34 & ~x37 & ~x39 & ~x46 & ~x47 & ~x48 & ~x49 & ~x51 & ~x57 & ~x58 & ~x62 & ~x67 & ~x68 & ~x70 & ~x78 & ~x79 & ~x80 & ~x86 & ~x88 & ~x90 & ~x93 & ~x95 & ~x96 & ~x97 & ~x99 & ~x101 & ~x104 & ~x106 & ~x108 & ~x109 & ~x111 & ~x112 & ~x113 & ~x116 & ~x118 & ~x119 & ~x126 & ~x127 & ~x133 & ~x135 & ~x136 & ~x137 & ~x138 & ~x139 & ~x140 & ~x141 & ~x143 & ~x144 & ~x146 & ~x162 & ~x165 & ~x167 & ~x171 & ~x172 & ~x191 & ~x193 & ~x196 & ~x197 & ~x220 & ~x223 & ~x226 & ~x228 & ~x248 & ~x250 & ~x251 & ~x252 & ~x253 & ~x278 & ~x279 & ~x280 & ~x306 & ~x309 & ~x310 & ~x312 & ~x333 & ~x338 & ~x340 & ~x359 & ~x361 & ~x363 & ~x366 & ~x368 & ~x385 & ~x386 & ~x389 & ~x393 & ~x394 & ~x395 & ~x417 & ~x418 & ~x419 & ~x424 & ~x425 & ~x444 & ~x447 & ~x450 & ~x451 & ~x474 & ~x475 & ~x476 & ~x482 & ~x486 & ~x500 & ~x501 & ~x503 & ~x504 & ~x505 & ~x507 & ~x509 & ~x511 & ~x512 & ~x513 & ~x533 & ~x537 & ~x539 & ~x541 & ~x542 & ~x559 & ~x562 & ~x563 & ~x564 & ~x565 & ~x568 & ~x569 & ~x588 & ~x589 & ~x593 & ~x597 & ~x611 & ~x615 & ~x617 & ~x620 & ~x622 & ~x624 & ~x639 & ~x640 & ~x642 & ~x643 & ~x647 & ~x649 & ~x651 & ~x652 & ~x654 & ~x668 & ~x669 & ~x670 & ~x673 & ~x676 & ~x677 & ~x678 & ~x680 & ~x707 & ~x709 & ~x710 & ~x711 & ~x712 & ~x727 & ~x730 & ~x737 & ~x741 & ~x752 & ~x767 & ~x769 & ~x774 & ~x775 & ~x778 & ~x779;
assign c8236 =  x152 &  x154 &  x233 &  x322 & ~x26 & ~x30 & ~x70 & ~x98 & ~x174 & ~x195 & ~x229 & ~x369 & ~x587 & ~x702;
assign c8238 =  x328 &  x405 & ~x285 & ~x297 & ~x401;
assign c8240 =  x503;
assign c8242 =  x156 &  x235 &  x322 & ~x26 & ~x43 & ~x95 & ~x113 & ~x164 & ~x170 & ~x231 & ~x286 & ~x364 & ~x420 & ~x498 & ~x503 & ~x526 & ~x545 & ~x556 & ~x740 & ~x757 & ~x767 & ~x775;
assign c8244 =  x734;
assign c8246 =  x343 &  x460 & ~x0 & ~x7 & ~x8 & ~x10 & ~x25 & ~x30 & ~x31 & ~x32 & ~x34 & ~x37 & ~x40 & ~x43 & ~x53 & ~x56 & ~x64 & ~x65 & ~x69 & ~x76 & ~x77 & ~x84 & ~x85 & ~x89 & ~x95 & ~x96 & ~x97 & ~x108 & ~x111 & ~x113 & ~x119 & ~x120 & ~x133 & ~x138 & ~x141 & ~x143 & ~x147 & ~x163 & ~x164 & ~x169 & ~x193 & ~x221 & ~x222 & ~x251 & ~x255 & ~x280 & ~x283 & ~x335 & ~x336 & ~x337 & ~x366 & ~x367 & ~x388 & ~x394 & ~x396 & ~x422 & ~x454 & ~x455 & ~x505 & ~x509 & ~x511 & ~x535 & ~x557 & ~x560 & ~x561 & ~x562 & ~x564 & ~x584 & ~x590 & ~x617 & ~x619 & ~x643 & ~x648 & ~x651 & ~x679 & ~x680 & ~x698 & ~x711 & ~x720 & ~x722 & ~x723 & ~x728 & ~x734 & ~x735 & ~x742 & ~x746 & ~x770 & ~x779;
assign c8248 =  x375 &  x434 & ~x0 & ~x8 & ~x9 & ~x10 & ~x12 & ~x13 & ~x15 & ~x19 & ~x21 & ~x22 & ~x23 & ~x25 & ~x26 & ~x29 & ~x30 & ~x31 & ~x32 & ~x35 & ~x36 & ~x37 & ~x38 & ~x39 & ~x41 & ~x42 & ~x43 & ~x46 & ~x49 & ~x50 & ~x51 & ~x54 & ~x55 & ~x57 & ~x58 & ~x59 & ~x61 & ~x67 & ~x71 & ~x72 & ~x75 & ~x76 & ~x79 & ~x83 & ~x85 & ~x86 & ~x87 & ~x94 & ~x97 & ~x98 & ~x99 & ~x100 & ~x107 & ~x114 & ~x115 & ~x116 & ~x119 & ~x122 & ~x136 & ~x139 & ~x141 & ~x144 & ~x145 & ~x146 & ~x167 & ~x169 & ~x170 & ~x171 & ~x174 & ~x194 & ~x196 & ~x197 & ~x199 & ~x200 & ~x220 & ~x222 & ~x224 & ~x226 & ~x228 & ~x229 & ~x248 & ~x251 & ~x253 & ~x256 & ~x276 & ~x277 & ~x279 & ~x280 & ~x304 & ~x305 & ~x306 & ~x307 & ~x334 & ~x335 & ~x336 & ~x337 & ~x349 & ~x361 & ~x367 & ~x388 & ~x389 & ~x390 & ~x391 & ~x396 & ~x398 & ~x399 & ~x418 & ~x419 & ~x421 & ~x423 & ~x425 & ~x426 & ~x427 & ~x429 & ~x430 & ~x442 & ~x443 & ~x444 & ~x445 & ~x451 & ~x453 & ~x454 & ~x455 & ~x457 & ~x470 & ~x471 & ~x472 & ~x479 & ~x480 & ~x483 & ~x498 & ~x499 & ~x500 & ~x501 & ~x505 & ~x508 & ~x510 & ~x511 & ~x528 & ~x529 & ~x530 & ~x532 & ~x536 & ~x538 & ~x554 & ~x555 & ~x556 & ~x557 & ~x559 & ~x560 & ~x561 & ~x562 & ~x563 & ~x564 & ~x583 & ~x584 & ~x585 & ~x586 & ~x591 & ~x592 & ~x614 & ~x616 & ~x618 & ~x639 & ~x641 & ~x642 & ~x643 & ~x645 & ~x646 & ~x648 & ~x668 & ~x669 & ~x670 & ~x676 & ~x678 & ~x695 & ~x697 & ~x702 & ~x703 & ~x705 & ~x708 & ~x709 & ~x721 & ~x722 & ~x724 & ~x731 & ~x733 & ~x736 & ~x737 & ~x738 & ~x742 & ~x743 & ~x744 & ~x745 & ~x746 & ~x748 & ~x749 & ~x758 & ~x761 & ~x763 & ~x765 & ~x766 & ~x769 & ~x770 & ~x772 & ~x774 & ~x775 & ~x779 & ~x780 & ~x782;
assign c8250 =  x159 &  x183 &  x462 &  x655;
assign c8252 =  x434 &  x629 & ~x26 & ~x33 & ~x34 & ~x48 & ~x55 & ~x56 & ~x57 & ~x71 & ~x72 & ~x76 & ~x77 & ~x83 & ~x107 & ~x111 & ~x114 & ~x120 & ~x121 & ~x123 & ~x140 & ~x143 & ~x172 & ~x175 & ~x201 & ~x205 & ~x225 & ~x230 & ~x248 & ~x254 & ~x279 & ~x280 & ~x282 & ~x314 & ~x336 & ~x338 & ~x339 & ~x362 & ~x365 & ~x368 & ~x388 & ~x396 & ~x416 & ~x424 & ~x441 & ~x446 & ~x473 & ~x476 & ~x481 & ~x484 & ~x496 & ~x499 & ~x501 & ~x526 & ~x530 & ~x531 & ~x534 & ~x551 & ~x552 & ~x564 & ~x578 & ~x581 & ~x588 & ~x611 & ~x617 & ~x641 & ~x647 & ~x660 & ~x670 & ~x674 & ~x703 & ~x721 & ~x725 & ~x732 & ~x751 & ~x753 & ~x768 & ~x772;
assign c8254 =  x142;
assign c8256 =  x53;
assign c8258 =  x410 & ~x8 & ~x15 & ~x25 & ~x26 & ~x47 & ~x55 & ~x57 & ~x67 & ~x70 & ~x75 & ~x78 & ~x79 & ~x85 & ~x95 & ~x100 & ~x119 & ~x122 & ~x134 & ~x137 & ~x145 & ~x167 & ~x169 & ~x177 & ~x221 & ~x229 & ~x252 & ~x255 & ~x257 & ~x284 & ~x325 & ~x352 & ~x353 & ~x362 & ~x424 & ~x476 & ~x480 & ~x494 & ~x495 & ~x497 & ~x499 & ~x504 & ~x505 & ~x525 & ~x551 & ~x557 & ~x580 & ~x585 & ~x610 & ~x614 & ~x616 & ~x618 & ~x648 & ~x672 & ~x673 & ~x697 & ~x702 & ~x705 & ~x721 & ~x727 & ~x731 & ~x733 & ~x735 & ~x743 & ~x744 & ~x765 & ~x771 & ~x782;
assign c8260 =  x353 &  x380 &  x407 & ~x57 & ~x70 & ~x72 & ~x80 & ~x82 & ~x90 & ~x110 & ~x112 & ~x114 & ~x146 & ~x251 & ~x254 & ~x258 & ~x269 & ~x309 & ~x397 & ~x398 & ~x410 & ~x414 & ~x416 & ~x419 & ~x427 & ~x439 & ~x444 & ~x453 & ~x472 & ~x475 & ~x503 & ~x507 & ~x525 & ~x582 & ~x584 & ~x592 & ~x609 & ~x666 & ~x678 & ~x691 & ~x702 & ~x707 & ~x728 & ~x734 & ~x753;
assign c8262 =  x357 & ~x55 & ~x89 & ~x327 & ~x494 & ~x524;
assign c8264 =  x588;
assign c8266 =  x17;
assign c8268 =  x459 &  x460 & ~x7 & ~x10 & ~x20 & ~x38 & ~x42 & ~x43 & ~x46 & ~x50 & ~x59 & ~x62 & ~x68 & ~x72 & ~x75 & ~x99 & ~x128 & ~x139 & ~x147 & ~x164 & ~x169 & ~x171 & ~x176 & ~x197 & ~x306 & ~x338 & ~x340 & ~x396 & ~x422 & ~x426 & ~x427 & ~x448 & ~x451 & ~x480 & ~x502 & ~x520 & ~x522 & ~x549 & ~x561 & ~x562 & ~x616 & ~x646 & ~x667 & ~x670 & ~x675 & ~x719 & ~x733 & ~x743 & ~x748 & ~x751 & ~x757 & ~x766 & ~x773;
assign c8270 =  x81;
assign c8272 =  x211 &  x431 & ~x155 & ~x429 & ~x576;
assign c8274 =  x406 &  x433 &  x486 & ~x70 & ~x150 & ~x177 & ~x428 & ~x543 & ~x555 & ~x607 & ~x675;
assign c8276 =  x290 &  x405 &  x408 &  x544 &  x631 & ~x7 & ~x18 & ~x29 & ~x31 & ~x32 & ~x41 & ~x44 & ~x60 & ~x76 & ~x88 & ~x91 & ~x93 & ~x98 & ~x105 & ~x108 & ~x117 & ~x138 & ~x142 & ~x144 & ~x162 & ~x225 & ~x253 & ~x282 & ~x310 & ~x312 & ~x363 & ~x414 & ~x416 & ~x417 & ~x445 & ~x449 & ~x451 & ~x477 & ~x510 & ~x528 & ~x530 & ~x536 & ~x584 & ~x587 & ~x590 & ~x666 & ~x668 & ~x669 & ~x696 & ~x721 & ~x726 & ~x753 & ~x755 & ~x775 & ~x782;
assign c8278 =  x382 &  x433 & ~x2 & ~x14 & ~x17 & ~x18 & ~x23 & ~x25 & ~x26 & ~x33 & ~x35 & ~x38 & ~x41 & ~x44 & ~x47 & ~x65 & ~x68 & ~x69 & ~x71 & ~x80 & ~x90 & ~x91 & ~x95 & ~x107 & ~x109 & ~x111 & ~x143 & ~x149 & ~x168 & ~x170 & ~x171 & ~x172 & ~x196 & ~x197 & ~x199 & ~x201 & ~x202 & ~x204 & ~x229 & ~x231 & ~x259 & ~x280 & ~x283 & ~x285 & ~x308 & ~x312 & ~x313 & ~x339 & ~x340 & ~x362 & ~x363 & ~x371 & ~x388 & ~x390 & ~x392 & ~x397 & ~x399 & ~x401 & ~x416 & ~x417 & ~x421 & ~x422 & ~x425 & ~x439 & ~x451 & ~x453 & ~x469 & ~x473 & ~x474 & ~x524 & ~x530 & ~x552 & ~x556 & ~x582 & ~x586 & ~x591 & ~x608 & ~x609 & ~x610 & ~x617 & ~x635 & ~x639 & ~x640 & ~x642 & ~x667 & ~x675 & ~x692 & ~x693 & ~x705 & ~x714 & ~x717 & ~x722 & ~x723 & ~x727 & ~x733 & ~x735 & ~x739 & ~x748 & ~x751 & ~x758 & ~x768 & ~x771 & ~x773 & ~x777 & ~x782;
assign c8280 =  x226;
assign c8282 =  x379 &  x405 &  x431 &  x485 & ~x8 & ~x15 & ~x20 & ~x36 & ~x51 & ~x65 & ~x73 & ~x79 & ~x80 & ~x117 & ~x123 & ~x306 & ~x360 & ~x362 & ~x385 & ~x399 & ~x441 & ~x453 & ~x475 & ~x481 & ~x516 & ~x589 & ~x614 & ~x636 & ~x700 & ~x702 & ~x707 & ~x713 & ~x746;
assign c8284 =  x384 &  x410 & ~x325 & ~x326 & ~x494 & ~x551;
assign c8286 =  x763;
assign c8288 =  x32;
assign c8290 =  x53;
assign c8292 =  x545 &  x607 & ~x283 & ~x333 & ~x511 & ~x514 & ~x569 & ~x615 & ~x625 & ~x677 & ~x759 & ~x762 & ~x777;
assign c8294 =  x290 &  x349 & ~x1 & ~x7 & ~x14 & ~x61 & ~x69 & ~x70 & ~x78 & ~x83 & ~x88 & ~x108 & ~x109 & ~x111 & ~x171 & ~x224 & ~x227 & ~x237 & ~x250 & ~x276 & ~x279 & ~x285 & ~x303 & ~x333 & ~x344 & ~x370 & ~x399 & ~x446 & ~x475 & ~x533 & ~x558 & ~x587 & ~x590 & ~x615 & ~x642 & ~x643 & ~x677 & ~x680 & ~x700 & ~x708 & ~x739 & ~x742 & ~x765;
assign c8296 =  x89;
assign c8298 =  x434 & ~x0 & ~x1 & ~x5 & ~x16 & ~x24 & ~x26 & ~x27 & ~x28 & ~x33 & ~x41 & ~x50 & ~x53 & ~x56 & ~x59 & ~x62 & ~x63 & ~x76 & ~x80 & ~x90 & ~x98 & ~x100 & ~x101 & ~x107 & ~x108 & ~x114 & ~x122 & ~x123 & ~x131 & ~x134 & ~x136 & ~x137 & ~x140 & ~x144 & ~x150 & ~x169 & ~x172 & ~x173 & ~x176 & ~x177 & ~x192 & ~x193 & ~x195 & ~x203 & ~x223 & ~x226 & ~x232 & ~x253 & ~x257 & ~x259 & ~x277 & ~x281 & ~x295 & ~x304 & ~x305 & ~x310 & ~x334 & ~x336 & ~x339 & ~x341 & ~x361 & ~x365 & ~x369 & ~x370 & ~x396 & ~x417 & ~x420 & ~x422 & ~x424 & ~x441 & ~x449 & ~x452 & ~x456 & ~x472 & ~x479 & ~x482 & ~x485 & ~x498 & ~x504 & ~x509 & ~x525 & ~x528 & ~x529 & ~x555 & ~x558 & ~x563 & ~x564 & ~x581 & ~x586 & ~x593 & ~x609 & ~x621 & ~x648 & ~x678 & ~x679 & ~x692 & ~x696 & ~x704 & ~x707 & ~x710 & ~x713 & ~x717 & ~x724 & ~x725 & ~x726 & ~x727 & ~x739 & ~x742 & ~x745 & ~x746 & ~x748 & ~x755 & ~x758 & ~x759 & ~x767 & ~x776 & ~x777 & ~x779 & ~x781 & ~x783;
assign c81 =  x658 & ~x17 & ~x18 & ~x36 & ~x39 & ~x58 & ~x67 & ~x72 & ~x74 & ~x77 & ~x94 & ~x98 & ~x99 & ~x111 & ~x137 & ~x142 & ~x170 & ~x196 & ~x200 & ~x225 & ~x341 & ~x365 & ~x394 & ~x418 & ~x421 & ~x473 & ~x477 & ~x481 & ~x482 & ~x503 & ~x506 & ~x511 & ~x513 & ~x514 & ~x515 & ~x516 & ~x545 & ~x560 & ~x589 & ~x614 & ~x618 & ~x666 & ~x671 & ~x673 & ~x707 & ~x725 & ~x729 & ~x734 & ~x741 & ~x751 & ~x755 & ~x759 & ~x760 & ~x775 & ~x780;
assign c83 =  x294 & ~x73 & ~x216 & ~x271 & ~x335 & ~x360 & ~x386 & ~x579 & ~x580 & ~x625 & ~x654 & ~x736 & ~x771;
assign c85 = ~x0 & ~x3 & ~x8 & ~x10 & ~x18 & ~x21 & ~x23 & ~x25 & ~x30 & ~x31 & ~x35 & ~x43 & ~x46 & ~x48 & ~x64 & ~x65 & ~x66 & ~x72 & ~x75 & ~x76 & ~x79 & ~x83 & ~x93 & ~x104 & ~x105 & ~x109 & ~x110 & ~x112 & ~x120 & ~x122 & ~x123 & ~x140 & ~x142 & ~x143 & ~x155 & ~x196 & ~x200 & ~x225 & ~x251 & ~x253 & ~x279 & ~x280 & ~x282 & ~x334 & ~x339 & ~x363 & ~x392 & ~x394 & ~x421 & ~x423 & ~x424 & ~x445 & ~x447 & ~x452 & ~x475 & ~x477 & ~x530 & ~x533 & ~x535 & ~x537 & ~x540 & ~x556 & ~x560 & ~x565 & ~x566 & ~x568 & ~x569 & ~x584 & ~x585 & ~x596 & ~x603 & ~x605 & ~x606 & ~x612 & ~x614 & ~x615 & ~x617 & ~x619 & ~x623 & ~x631 & ~x632 & ~x633 & ~x634 & ~x643 & ~x645 & ~x649 & ~x659 & ~x661 & ~x662 & ~x668 & ~x669 & ~x671 & ~x675 & ~x677 & ~x690 & ~x695 & ~x696 & ~x699 & ~x715 & ~x724 & ~x727 & ~x744 & ~x746 & ~x748 & ~x751 & ~x753 & ~x757 & ~x762 & ~x767 & ~x770 & ~x771;
assign c87 =  x543 &  x544 &  x570 & ~x15 & ~x19 & ~x83 & ~x116 & ~x248 & ~x257 & ~x285 & ~x312 & ~x343 & ~x505 & ~x506 & ~x530 & ~x646 & ~x655 & ~x657 & ~x658 & ~x683 & ~x687 & ~x691 & ~x709 & ~x729 & ~x740 & ~x754 & ~x772 & ~x775 & ~x783;
assign c89 =  x483 & ~x27 & ~x44 & ~x47 & ~x50 & ~x57 & ~x112 & ~x138 & ~x378 & ~x379 & ~x447 & ~x502 & ~x503 & ~x614 & ~x710 & ~x750 & ~x775 & ~x783;
assign c811 = ~x7 & ~x11 & ~x13 & ~x14 & ~x19 & ~x26 & ~x30 & ~x31 & ~x37 & ~x44 & ~x47 & ~x48 & ~x51 & ~x58 & ~x80 & ~x86 & ~x89 & ~x108 & ~x110 & ~x111 & ~x140 & ~x167 & ~x193 & ~x197 & ~x220 & ~x221 & ~x224 & ~x225 & ~x229 & ~x248 & ~x249 & ~x250 & ~x264 & ~x265 & ~x266 & ~x277 & ~x278 & ~x284 & ~x291 & ~x292 & ~x293 & ~x311 & ~x319 & ~x320 & ~x334 & ~x335 & ~x340 & ~x346 & ~x362 & ~x363 & ~x364 & ~x368 & ~x374 & ~x448 & ~x450 & ~x502 & ~x530 & ~x531 & ~x532 & ~x589 & ~x615 & ~x643 & ~x660 & ~x662 & ~x671 & ~x684 & ~x688 & ~x690 & ~x696 & ~x697 & ~x698 & ~x703 & ~x704 & ~x705 & ~x710 & ~x712 & ~x717 & ~x718 & ~x721 & ~x724 & ~x727 & ~x732 & ~x735 & ~x738 & ~x740 & ~x747 & ~x756 & ~x758 & ~x760 & ~x761 & ~x762 & ~x768 & ~x782;
assign c813 = ~x2 & ~x3 & ~x4 & ~x5 & ~x6 & ~x11 & ~x12 & ~x16 & ~x19 & ~x21 & ~x24 & ~x25 & ~x28 & ~x32 & ~x36 & ~x38 & ~x40 & ~x41 & ~x42 & ~x44 & ~x45 & ~x49 & ~x56 & ~x60 & ~x62 & ~x63 & ~x66 & ~x68 & ~x69 & ~x75 & ~x88 & ~x90 & ~x91 & ~x104 & ~x105 & ~x106 & ~x109 & ~x110 & ~x111 & ~x113 & ~x134 & ~x135 & ~x137 & ~x141 & ~x143 & ~x163 & ~x166 & ~x167 & ~x192 & ~x195 & ~x196 & ~x199 & ~x201 & ~x219 & ~x220 & ~x226 & ~x229 & ~x248 & ~x253 & ~x275 & ~x277 & ~x294 & ~x304 & ~x306 & ~x339 & ~x340 & ~x349 & ~x350 & ~x361 & ~x366 & ~x368 & ~x369 & ~x370 & ~x376 & ~x388 & ~x390 & ~x392 & ~x393 & ~x403 & ~x451 & ~x474 & ~x477 & ~x480 & ~x506 & ~x507 & ~x559 & ~x584 & ~x588 & ~x590 & ~x618 & ~x642 & ~x643 & ~x649 & ~x670 & ~x671 & ~x674 & ~x676 & ~x696 & ~x699 & ~x700 & ~x701 & ~x715 & ~x726 & ~x727 & ~x732 & ~x733 & ~x741 & ~x744 & ~x746 & ~x751 & ~x753 & ~x755 & ~x756 & ~x757 & ~x759 & ~x763 & ~x764 & ~x766 & ~x767 & ~x773 & ~x776 & ~x779 & ~x780 & ~x782;
assign c815 = ~x7 & ~x20 & ~x39 & ~x41 & ~x63 & ~x65 & ~x76 & ~x90 & ~x115 & ~x167 & ~x195 & ~x199 & ~x221 & ~x251 & ~x252 & ~x429 & ~x433 & ~x434 & ~x447 & ~x458 & ~x459 & ~x486 & ~x487 & ~x488 & ~x501 & ~x504 & ~x530 & ~x558 & ~x587 & ~x589 & ~x614 & ~x643 & ~x644 & ~x647 & ~x698 & ~x699 & ~x709 & ~x732 & ~x749 & ~x756;
assign c817 =  x408 &  x436 & ~x1 & ~x15 & ~x23 & ~x29 & ~x35 & ~x37 & ~x53 & ~x55 & ~x56 & ~x62 & ~x63 & ~x65 & ~x75 & ~x88 & ~x95 & ~x109 & ~x110 & ~x138 & ~x142 & ~x162 & ~x170 & ~x190 & ~x192 & ~x195 & ~x227 & ~x249 & ~x251 & ~x254 & ~x276 & ~x303 & ~x306 & ~x307 & ~x309 & ~x322 & ~x330 & ~x331 & ~x335 & ~x340 & ~x349 & ~x361 & ~x448 & ~x474 & ~x478 & ~x533 & ~x659 & ~x672 & ~x687 & ~x698 & ~x727 & ~x751 & ~x762 & ~x768 & ~x769 & ~x774 & ~x780 & ~x782;
assign c819 =  x162;
assign c821 =  x517 & ~x4 & ~x9 & ~x12 & ~x25 & ~x35 & ~x39 & ~x48 & ~x50 & ~x64 & ~x65 & ~x82 & ~x83 & ~x97 & ~x99 & ~x106 & ~x108 & ~x132 & ~x164 & ~x168 & ~x189 & ~x220 & ~x281 & ~x285 & ~x291 & ~x318 & ~x330 & ~x344 & ~x366 & ~x395 & ~x396 & ~x412 & ~x419 & ~x424 & ~x450 & ~x498 & ~x505 & ~x506 & ~x511 & ~x586 & ~x587 & ~x613 & ~x614 & ~x645 & ~x667 & ~x671 & ~x694 & ~x697 & ~x698 & ~x699 & ~x701 & ~x713 & ~x715 & ~x730 & ~x731 & ~x748 & ~x752;
assign c823 =  x584;
assign c825 = ~x33 & ~x53 & ~x74 & ~x115 & ~x119 & ~x135 & ~x185 & ~x211 & ~x214 & ~x378 & ~x390 & ~x500 & ~x529 & ~x593 & ~x615 & ~x647 & ~x728 & ~x729;
assign c827 = ~x3 & ~x14 & ~x15 & ~x42 & ~x46 & ~x52 & ~x60 & ~x65 & ~x85 & ~x87 & ~x88 & ~x98 & ~x110 & ~x113 & ~x118 & ~x124 & ~x140 & ~x141 & ~x143 & ~x168 & ~x225 & ~x253 & ~x280 & ~x307 & ~x334 & ~x339 & ~x364 & ~x390 & ~x406 & ~x407 & ~x408 & ~x436 & ~x445 & ~x447 & ~x462 & ~x489 & ~x490 & ~x502 & ~x504 & ~x534 & ~x559 & ~x563 & ~x586 & ~x590 & ~x612 & ~x642 & ~x670 & ~x705 & ~x726 & ~x727 & ~x729 & ~x731 & ~x733 & ~x741 & ~x748 & ~x749 & ~x763 & ~x764 & ~x782;
assign c829 =  x653 & ~x5 & ~x43 & ~x82 & ~x83 & ~x96 & ~x103 & ~x279 & ~x364 & ~x416 & ~x455 & ~x482 & ~x485 & ~x515 & ~x639 & ~x754 & ~x763;
assign c831 = ~x11 & ~x16 & ~x17 & ~x19 & ~x26 & ~x30 & ~x46 & ~x47 & ~x48 & ~x49 & ~x52 & ~x57 & ~x69 & ~x74 & ~x84 & ~x103 & ~x110 & ~x114 & ~x115 & ~x135 & ~x140 & ~x142 & ~x169 & ~x170 & ~x225 & ~x250 & ~x251 & ~x252 & ~x264 & ~x265 & ~x266 & ~x275 & ~x276 & ~x277 & ~x280 & ~x282 & ~x285 & ~x287 & ~x290 & ~x291 & ~x292 & ~x293 & ~x305 & ~x308 & ~x317 & ~x319 & ~x320 & ~x338 & ~x344 & ~x345 & ~x346 & ~x363 & ~x369 & ~x389 & ~x392 & ~x394 & ~x398 & ~x417 & ~x419 & ~x420 & ~x422 & ~x449 & ~x450 & ~x614 & ~x616 & ~x618 & ~x620 & ~x646 & ~x647 & ~x666 & ~x673 & ~x691 & ~x693 & ~x699 & ~x705 & ~x719 & ~x721 & ~x722 & ~x725 & ~x733 & ~x744 & ~x751 & ~x752 & ~x758 & ~x759 & ~x761 & ~x769 & ~x773 & ~x776 & ~x777 & ~x783;
assign c833 = ~x0 & ~x1 & ~x2 & ~x8 & ~x9 & ~x17 & ~x20 & ~x22 & ~x32 & ~x33 & ~x38 & ~x47 & ~x50 & ~x57 & ~x60 & ~x61 & ~x64 & ~x65 & ~x68 & ~x76 & ~x79 & ~x80 & ~x88 & ~x89 & ~x104 & ~x106 & ~x107 & ~x115 & ~x116 & ~x117 & ~x134 & ~x135 & ~x138 & ~x141 & ~x143 & ~x163 & ~x168 & ~x190 & ~x192 & ~x196 & ~x197 & ~x198 & ~x219 & ~x222 & ~x227 & ~x248 & ~x249 & ~x253 & ~x278 & ~x281 & ~x307 & ~x311 & ~x333 & ~x335 & ~x350 & ~x362 & ~x364 & ~x366 & ~x377 & ~x394 & ~x417 & ~x418 & ~x420 & ~x432 & ~x445 & ~x450 & ~x451 & ~x474 & ~x502 & ~x503 & ~x504 & ~x531 & ~x536 & ~x557 & ~x558 & ~x561 & ~x585 & ~x589 & ~x591 & ~x613 & ~x615 & ~x641 & ~x671 & ~x672 & ~x673 & ~x692 & ~x693 & ~x695 & ~x697 & ~x700 & ~x701 & ~x710 & ~x713 & ~x723 & ~x724 & ~x730 & ~x731 & ~x733 & ~x739 & ~x740 & ~x748 & ~x752 & ~x756 & ~x761 & ~x766 & ~x767 & ~x768 & ~x772 & ~x774 & ~x776 & ~x777 & ~x781;
assign c835 =  x374 &  x375 &  x429 &  x430 &  x457 & ~x4 & ~x8 & ~x11 & ~x17 & ~x18 & ~x25 & ~x29 & ~x32 & ~x39 & ~x41 & ~x44 & ~x45 & ~x46 & ~x49 & ~x50 & ~x56 & ~x61 & ~x64 & ~x69 & ~x74 & ~x75 & ~x83 & ~x87 & ~x91 & ~x92 & ~x97 & ~x111 & ~x112 & ~x114 & ~x122 & ~x140 & ~x143 & ~x145 & ~x148 & ~x168 & ~x169 & ~x171 & ~x176 & ~x177 & ~x179 & ~x196 & ~x200 & ~x203 & ~x204 & ~x229 & ~x231 & ~x232 & ~x233 & ~x251 & ~x252 & ~x253 & ~x259 & ~x277 & ~x278 & ~x281 & ~x286 & ~x308 & ~x310 & ~x312 & ~x314 & ~x332 & ~x340 & ~x341 & ~x343 & ~x360 & ~x361 & ~x362 & ~x370 & ~x388 & ~x389 & ~x390 & ~x392 & ~x418 & ~x420 & ~x424 & ~x449 & ~x451 & ~x452 & ~x473 & ~x501 & ~x502 & ~x504 & ~x505 & ~x506 & ~x507 & ~x529 & ~x530 & ~x532 & ~x533 & ~x534 & ~x535 & ~x563 & ~x608 & ~x613 & ~x616 & ~x620 & ~x621 & ~x637 & ~x639 & ~x641 & ~x649 & ~x650 & ~x663 & ~x665 & ~x666 & ~x667 & ~x669 & ~x673 & ~x688 & ~x689 & ~x693 & ~x696 & ~x697 & ~x706 & ~x709 & ~x715 & ~x716 & ~x719 & ~x721 & ~x726 & ~x736 & ~x737 & ~x738 & ~x742 & ~x749 & ~x750 & ~x752 & ~x756 & ~x758 & ~x760 & ~x761 & ~x762 & ~x763 & ~x765 & ~x771 & ~x775 & ~x778 & ~x780 & ~x783;
assign c837 =  x566 &  x569 & ~x6 & ~x38 & ~x40 & ~x50 & ~x58 & ~x71 & ~x78 & ~x81 & ~x86 & ~x91 & ~x114 & ~x118 & ~x168 & ~x222 & ~x248 & ~x283 & ~x303 & ~x306 & ~x310 & ~x332 & ~x339 & ~x390 & ~x446 & ~x471 & ~x500 & ~x531 & ~x534 & ~x559 & ~x589 & ~x616 & ~x672 & ~x679 & ~x696 & ~x707 & ~x718 & ~x719 & ~x724 & ~x731 & ~x732 & ~x734 & ~x736 & ~x737 & ~x754 & ~x767;
assign c839 =  x146;
assign c841 = ~x4 & ~x7 & ~x10 & ~x14 & ~x20 & ~x25 & ~x26 & ~x31 & ~x37 & ~x41 & ~x42 & ~x45 & ~x48 & ~x63 & ~x69 & ~x70 & ~x71 & ~x80 & ~x87 & ~x90 & ~x94 & ~x95 & ~x98 & ~x105 & ~x107 & ~x110 & ~x111 & ~x113 & ~x114 & ~x134 & ~x135 & ~x141 & ~x145 & ~x166 & ~x169 & ~x170 & ~x195 & ~x196 & ~x198 & ~x225 & ~x226 & ~x254 & ~x280 & ~x310 & ~x311 & ~x313 & ~x315 & ~x333 & ~x338 & ~x339 & ~x340 & ~x342 & ~x363 & ~x366 & ~x368 & ~x370 & ~x392 & ~x394 & ~x397 & ~x399 & ~x417 & ~x420 & ~x425 & ~x427 & ~x455 & ~x456 & ~x480 & ~x485 & ~x486 & ~x504 & ~x515 & ~x516 & ~x532 & ~x534 & ~x615 & ~x643 & ~x645 & ~x693 & ~x694 & ~x696 & ~x715 & ~x720 & ~x722 & ~x726 & ~x728 & ~x729 & ~x748 & ~x767 & ~x776 & ~x777;
assign c843 = ~x0 & ~x4 & ~x9 & ~x11 & ~x17 & ~x22 & ~x42 & ~x44 & ~x45 & ~x51 & ~x55 & ~x56 & ~x61 & ~x62 & ~x64 & ~x65 & ~x68 & ~x81 & ~x109 & ~x114 & ~x117 & ~x133 & ~x137 & ~x142 & ~x174 & ~x196 & ~x198 & ~x225 & ~x227 & ~x229 & ~x248 & ~x254 & ~x255 & ~x256 & ~x279 & ~x312 & ~x313 & ~x336 & ~x366 & ~x389 & ~x391 & ~x394 & ~x445 & ~x447 & ~x477 & ~x530 & ~x531 & ~x533 & ~x535 & ~x558 & ~x564 & ~x565 & ~x581 & ~x586 & ~x589 & ~x590 & ~x595 & ~x596 & ~x617 & ~x630 & ~x632 & ~x638 & ~x639 & ~x641 & ~x643 & ~x649 & ~x660 & ~x661 & ~x667 & ~x668 & ~x670 & ~x676 & ~x687 & ~x688 & ~x695 & ~x696 & ~x701 & ~x705 & ~x718 & ~x719 & ~x731 & ~x738 & ~x743 & ~x746 & ~x758 & ~x763 & ~x765 & ~x769 & ~x772 & ~x782;
assign c845 =  x578 & ~x301 & ~x330 & ~x616 & ~x652 & ~x656 & ~x659 & ~x660 & ~x683 & ~x687;
assign c847 =  x268 & ~x12 & ~x20 & ~x66 & ~x87 & ~x138 & ~x154 & ~x183 & ~x203 & ~x210 & ~x231 & ~x308 & ~x329 & ~x331 & ~x333 & ~x342 & ~x359 & ~x422 & ~x641 & ~x696 & ~x699 & ~x708 & ~x753;
assign c849 = ~x3 & ~x4 & ~x10 & ~x12 & ~x14 & ~x16 & ~x26 & ~x33 & ~x47 & ~x61 & ~x63 & ~x72 & ~x75 & ~x79 & ~x87 & ~x96 & ~x100 & ~x102 & ~x108 & ~x121 & ~x125 & ~x127 & ~x157 & ~x165 & ~x170 & ~x174 & ~x181 & ~x195 & ~x250 & ~x251 & ~x253 & ~x306 & ~x333 & ~x358 & ~x359 & ~x360 & ~x364 & ~x365 & ~x387 & ~x388 & ~x390 & ~x393 & ~x479 & ~x532 & ~x533 & ~x601 & ~x602 & ~x629 & ~x643 & ~x656 & ~x657 & ~x667 & ~x676 & ~x683 & ~x684 & ~x711 & ~x723 & ~x727 & ~x740 & ~x754 & ~x755 & ~x757 & ~x758 & ~x761 & ~x763 & ~x771;
assign c851 =  x599 &  x626 & ~x2 & ~x15 & ~x18 & ~x20 & ~x23 & ~x25 & ~x26 & ~x28 & ~x34 & ~x40 & ~x42 & ~x44 & ~x50 & ~x52 & ~x60 & ~x65 & ~x75 & ~x83 & ~x90 & ~x93 & ~x99 & ~x107 & ~x112 & ~x113 & ~x116 & ~x143 & ~x144 & ~x164 & ~x171 & ~x251 & ~x252 & ~x253 & ~x334 & ~x336 & ~x339 & ~x362 & ~x363 & ~x365 & ~x367 & ~x368 & ~x389 & ~x394 & ~x395 & ~x419 & ~x449 & ~x450 & ~x452 & ~x457 & ~x475 & ~x487 & ~x500 & ~x502 & ~x506 & ~x528 & ~x533 & ~x555 & ~x557 & ~x584 & ~x585 & ~x589 & ~x616 & ~x648 & ~x676 & ~x692 & ~x701 & ~x713 & ~x714 & ~x720 & ~x723 & ~x746 & ~x748 & ~x752 & ~x754 & ~x755 & ~x757 & ~x758 & ~x759 & ~x761 & ~x765 & ~x769 & ~x776 & ~x778 & ~x779 & ~x780;
assign c853 = ~x1 & ~x7 & ~x17 & ~x20 & ~x25 & ~x26 & ~x35 & ~x40 & ~x44 & ~x47 & ~x49 & ~x50 & ~x51 & ~x59 & ~x62 & ~x67 & ~x90 & ~x94 & ~x112 & ~x117 & ~x118 & ~x144 & ~x145 & ~x150 & ~x154 & ~x200 & ~x225 & ~x253 & ~x275 & ~x280 & ~x282 & ~x336 & ~x390 & ~x423 & ~x445 & ~x448 & ~x473 & ~x477 & ~x499 & ~x502 & ~x503 & ~x505 & ~x506 & ~x530 & ~x533 & ~x558 & ~x562 & ~x601 & ~x610 & ~x612 & ~x628 & ~x642 & ~x644 & ~x655 & ~x684 & ~x695 & ~x723 & ~x736 & ~x738 & ~x751 & ~x753 & ~x767 & ~x768 & ~x771 & ~x772 & ~x777;
assign c855 = ~x0 & ~x1 & ~x13 & ~x15 & ~x25 & ~x27 & ~x30 & ~x33 & ~x43 & ~x46 & ~x56 & ~x61 & ~x84 & ~x87 & ~x89 & ~x90 & ~x102 & ~x104 & ~x105 & ~x112 & ~x119 & ~x129 & ~x133 & ~x163 & ~x165 & ~x166 & ~x168 & ~x169 & ~x172 & ~x201 & ~x222 & ~x248 & ~x257 & ~x278 & ~x279 & ~x336 & ~x394 & ~x395 & ~x419 & ~x473 & ~x480 & ~x507 & ~x527 & ~x532 & ~x536 & ~x557 & ~x563 & ~x564 & ~x565 & ~x566 & ~x568 & ~x571 & ~x578 & ~x580 & ~x592 & ~x597 & ~x598 & ~x620 & ~x621 & ~x636 & ~x637 & ~x642 & ~x667 & ~x707 & ~x719 & ~x728 & ~x731 & ~x734 & ~x736 & ~x741 & ~x757 & ~x765 & ~x767 & ~x771 & ~x778 & ~x779 & ~x781 & ~x783;
assign c857 =  x125 & ~x349;
assign c859 = ~x18 & ~x22 & ~x25 & ~x26 & ~x27 & ~x30 & ~x37 & ~x42 & ~x45 & ~x50 & ~x63 & ~x64 & ~x65 & ~x71 & ~x75 & ~x77 & ~x79 & ~x80 & ~x84 & ~x91 & ~x142 & ~x194 & ~x195 & ~x196 & ~x230 & ~x278 & ~x307 & ~x310 & ~x339 & ~x379 & ~x392 & ~x406 & ~x407 & ~x408 & ~x436 & ~x437 & ~x451 & ~x474 & ~x504 & ~x530 & ~x533 & ~x560 & ~x561 & ~x562 & ~x642 & ~x646 & ~x673 & ~x676 & ~x688 & ~x703 & ~x714 & ~x720 & ~x723 & ~x728 & ~x729 & ~x743 & ~x746 & ~x750 & ~x755 & ~x779;
assign c861 =  x596 & ~x0 & ~x4 & ~x5 & ~x7 & ~x8 & ~x9 & ~x17 & ~x26 & ~x28 & ~x30 & ~x34 & ~x36 & ~x43 & ~x44 & ~x46 & ~x48 & ~x50 & ~x61 & ~x63 & ~x66 & ~x67 & ~x73 & ~x88 & ~x92 & ~x99 & ~x103 & ~x106 & ~x107 & ~x110 & ~x114 & ~x170 & ~x171 & ~x196 & ~x198 & ~x199 & ~x223 & ~x228 & ~x253 & ~x255 & ~x279 & ~x307 & ~x308 & ~x309 & ~x337 & ~x362 & ~x390 & ~x393 & ~x395 & ~x396 & ~x416 & ~x420 & ~x421 & ~x422 & ~x445 & ~x452 & ~x456 & ~x473 & ~x476 & ~x485 & ~x488 & ~x530 & ~x531 & ~x556 & ~x560 & ~x561 & ~x613 & ~x646 & ~x667 & ~x668 & ~x674 & ~x675 & ~x694 & ~x701 & ~x702 & ~x715 & ~x717 & ~x734 & ~x737 & ~x740 & ~x741 & ~x747 & ~x751 & ~x754 & ~x755 & ~x757 & ~x760 & ~x770 & ~x778 & ~x783;
assign c863 = ~x33 & ~x90 & ~x99 & ~x111 & ~x116 & ~x139 & ~x169 & ~x199 & ~x253 & ~x259 & ~x263 & ~x276 & ~x279 & ~x286 & ~x289 & ~x290 & ~x298 & ~x299 & ~x300 & ~x307 & ~x310 & ~x314 & ~x328 & ~x330 & ~x331 & ~x340 & ~x343 & ~x344 & ~x356 & ~x364 & ~x387 & ~x395 & ~x416 & ~x417 & ~x424 & ~x447 & ~x477 & ~x481 & ~x504 & ~x507 & ~x557 & ~x591 & ~x617 & ~x641 & ~x675 & ~x701 & ~x726 & ~x737 & ~x741 & ~x745 & ~x748 & ~x751 & ~x773;
assign c865 = ~x9 & ~x10 & ~x12 & ~x13 & ~x25 & ~x37 & ~x38 & ~x41 & ~x44 & ~x50 & ~x58 & ~x60 & ~x62 & ~x64 & ~x71 & ~x72 & ~x86 & ~x88 & ~x91 & ~x99 & ~x104 & ~x107 & ~x116 & ~x121 & ~x130 & ~x131 & ~x138 & ~x151 & ~x154 & ~x158 & ~x197 & ~x224 & ~x247 & ~x303 & ~x304 & ~x337 & ~x363 & ~x365 & ~x366 & ~x447 & ~x450 & ~x501 & ~x532 & ~x534 & ~x560 & ~x563 & ~x572 & ~x586 & ~x587 & ~x598 & ~x599 & ~x618 & ~x619 & ~x626 & ~x639 & ~x647 & ~x649 & ~x654 & ~x668 & ~x677 & ~x681 & ~x682 & ~x724 & ~x752 & ~x759 & ~x762 & ~x773 & ~x776;
assign c867 = ~x3 & ~x5 & ~x8 & ~x13 & ~x29 & ~x35 & ~x37 & ~x46 & ~x48 & ~x53 & ~x55 & ~x60 & ~x66 & ~x68 & ~x69 & ~x76 & ~x80 & ~x83 & ~x94 & ~x95 & ~x109 & ~x119 & ~x121 & ~x138 & ~x142 & ~x144 & ~x145 & ~x146 & ~x149 & ~x169 & ~x197 & ~x224 & ~x226 & ~x251 & ~x281 & ~x287 & ~x302 & ~x303 & ~x306 & ~x323 & ~x324 & ~x325 & ~x327 & ~x328 & ~x329 & ~x330 & ~x337 & ~x338 & ~x352 & ~x355 & ~x356 & ~x358 & ~x359 & ~x360 & ~x363 & ~x364 & ~x385 & ~x386 & ~x390 & ~x397 & ~x419 & ~x423 & ~x425 & ~x450 & ~x451 & ~x452 & ~x472 & ~x473 & ~x474 & ~x499 & ~x507 & ~x531 & ~x534 & ~x562 & ~x564 & ~x583 & ~x585 & ~x586 & ~x615 & ~x616 & ~x636 & ~x637 & ~x640 & ~x643 & ~x647 & ~x663 & ~x665 & ~x668 & ~x671 & ~x672 & ~x675 & ~x676 & ~x679 & ~x692 & ~x695 & ~x696 & ~x698 & ~x699 & ~x705 & ~x722 & ~x726 & ~x728 & ~x730 & ~x731 & ~x732 & ~x737 & ~x740 & ~x750 & ~x755 & ~x756 & ~x761 & ~x764 & ~x765 & ~x768 & ~x772 & ~x773 & ~x780 & ~x781;
assign c869 =  x547 & ~x14 & ~x40 & ~x106 & ~x112 & ~x114 & ~x166 & ~x194 & ~x335 & ~x390 & ~x392 & ~x419 & ~x422 & ~x445 & ~x477 & ~x508 & ~x556 & ~x558 & ~x571 & ~x607 & ~x624 & ~x627 & ~x644 & ~x652 & ~x654 & ~x733 & ~x734 & ~x746;
assign c871 = ~x27 & ~x28 & ~x112 & ~x135 & ~x140 & ~x141 & ~x142 & ~x162 & ~x175 & ~x193 & ~x200 & ~x224 & ~x248 & ~x250 & ~x274 & ~x284 & ~x294 & ~x312 & ~x322 & ~x323 & ~x333 & ~x337 & ~x447 & ~x471 & ~x656 & ~x658 & ~x659 & ~x673 & ~x689 & ~x699 & ~x724 & ~x734 & ~x736 & ~x768 & ~x771;
assign c873 = ~x34 & ~x37 & ~x57 & ~x71 & ~x78 & ~x86 & ~x93 & ~x113 & ~x117 & ~x143 & ~x156 & ~x200 & ~x226 & ~x252 & ~x255 & ~x277 & ~x283 & ~x312 & ~x335 & ~x340 & ~x349 & ~x361 & ~x363 & ~x391 & ~x396 & ~x446 & ~x449 & ~x476 & ~x478 & ~x555 & ~x588 & ~x589 & ~x596 & ~x597 & ~x598 & ~x611 & ~x624 & ~x625 & ~x639 & ~x648 & ~x650 & ~x660 & ~x661 & ~x667 & ~x671 & ~x672 & ~x673 & ~x679 & ~x717 & ~x724 & ~x730 & ~x733 & ~x744 & ~x746 & ~x760 & ~x763 & ~x768 & ~x773;
assign c875 = ~x2 & ~x5 & ~x10 & ~x14 & ~x16 & ~x20 & ~x21 & ~x25 & ~x29 & ~x31 & ~x32 & ~x34 & ~x40 & ~x44 & ~x46 & ~x47 & ~x49 & ~x60 & ~x62 & ~x78 & ~x108 & ~x111 & ~x112 & ~x135 & ~x142 & ~x144 & ~x199 & ~x228 & ~x250 & ~x255 & ~x282 & ~x307 & ~x309 & ~x337 & ~x351 & ~x364 & ~x365 & ~x380 & ~x395 & ~x417 & ~x421 & ~x422 & ~x443 & ~x446 & ~x451 & ~x480 & ~x488 & ~x517 & ~x534 & ~x535 & ~x559 & ~x584 & ~x588 & ~x612 & ~x615 & ~x670 & ~x677 & ~x689 & ~x707 & ~x719 & ~x726 & ~x730 & ~x733 & ~x734 & ~x746 & ~x759 & ~x766 & ~x782;
assign c877 = ~x4 & ~x7 & ~x8 & ~x9 & ~x10 & ~x13 & ~x15 & ~x22 & ~x25 & ~x32 & ~x38 & ~x54 & ~x55 & ~x56 & ~x60 & ~x65 & ~x67 & ~x75 & ~x76 & ~x79 & ~x81 & ~x84 & ~x85 & ~x88 & ~x89 & ~x90 & ~x92 & ~x110 & ~x114 & ~x116 & ~x117 & ~x138 & ~x141 & ~x143 & ~x173 & ~x194 & ~x199 & ~x223 & ~x252 & ~x253 & ~x254 & ~x265 & ~x275 & ~x280 & ~x292 & ~x303 & ~x305 & ~x310 & ~x311 & ~x317 & ~x318 & ~x319 & ~x337 & ~x338 & ~x340 & ~x343 & ~x345 & ~x357 & ~x363 & ~x364 & ~x366 & ~x386 & ~x390 & ~x392 & ~x395 & ~x399 & ~x413 & ~x415 & ~x417 & ~x418 & ~x442 & ~x446 & ~x448 & ~x476 & ~x477 & ~x479 & ~x506 & ~x534 & ~x558 & ~x560 & ~x585 & ~x586 & ~x589 & ~x641 & ~x647 & ~x681 & ~x682 & ~x684 & ~x685 & ~x686 & ~x687 & ~x688 & ~x702 & ~x704 & ~x710 & ~x711 & ~x712 & ~x713 & ~x724 & ~x726 & ~x728 & ~x733 & ~x743 & ~x745 & ~x746 & ~x749 & ~x753 & ~x754 & ~x756 & ~x758 & ~x765 & ~x766 & ~x773 & ~x781 & ~x782;
assign c879 =  x426 & ~x12 & ~x14 & ~x15 & ~x18 & ~x32 & ~x35 & ~x36 & ~x77 & ~x81 & ~x82 & ~x87 & ~x110 & ~x119 & ~x131 & ~x144 & ~x224 & ~x279 & ~x282 & ~x283 & ~x284 & ~x419 & ~x420 & ~x446 & ~x589 & ~x614 & ~x638 & ~x703 & ~x730 & ~x737 & ~x749 & ~x761;
assign c881 =  x118;
assign c883 = ~x0 & ~x2 & ~x5 & ~x6 & ~x7 & ~x9 & ~x10 & ~x11 & ~x16 & ~x18 & ~x22 & ~x23 & ~x26 & ~x29 & ~x31 & ~x38 & ~x41 & ~x47 & ~x50 & ~x51 & ~x54 & ~x56 & ~x57 & ~x59 & ~x61 & ~x63 & ~x68 & ~x71 & ~x82 & ~x85 & ~x91 & ~x93 & ~x95 & ~x97 & ~x99 & ~x104 & ~x106 & ~x107 & ~x112 & ~x115 & ~x118 & ~x136 & ~x137 & ~x139 & ~x165 & ~x166 & ~x170 & ~x171 & ~x196 & ~x197 & ~x199 & ~x225 & ~x252 & ~x254 & ~x255 & ~x276 & ~x279 & ~x280 & ~x303 & ~x304 & ~x306 & ~x307 & ~x308 & ~x330 & ~x332 & ~x340 & ~x359 & ~x361 & ~x362 & ~x365 & ~x366 & ~x367 & ~x368 & ~x391 & ~x395 & ~x416 & ~x417 & ~x418 & ~x419 & ~x423 & ~x452 & ~x473 & ~x476 & ~x478 & ~x479 & ~x504 & ~x505 & ~x511 & ~x513 & ~x515 & ~x530 & ~x534 & ~x537 & ~x538 & ~x542 & ~x544 & ~x545 & ~x546 & ~x558 & ~x560 & ~x562 & ~x563 & ~x564 & ~x565 & ~x584 & ~x589 & ~x613 & ~x614 & ~x640 & ~x644 & ~x672 & ~x674 & ~x694 & ~x696 & ~x698 & ~x703 & ~x722 & ~x728 & ~x729 & ~x733 & ~x737 & ~x739 & ~x741 & ~x748 & ~x760 & ~x763 & ~x764 & ~x766 & ~x770 & ~x773 & ~x774 & ~x775 & ~x776 & ~x777 & ~x778 & ~x779 & ~x781 & ~x783;
assign c885 =  x209 &  x212 & ~x34 & ~x35 & ~x37 & ~x42 & ~x82 & ~x94 & ~x111 & ~x120 & ~x137 & ~x141 & ~x169 & ~x224 & ~x248 & ~x432 & ~x433 & ~x458 & ~x474 & ~x475 & ~x477 & ~x500 & ~x506 & ~x561 & ~x615 & ~x617 & ~x676 & ~x702 & ~x704 & ~x723 & ~x760 & ~x766 & ~x779 & ~x783;
assign c887 =  x466 &  x548 & ~x0 & ~x16 & ~x18 & ~x35 & ~x37 & ~x79 & ~x85 & ~x93 & ~x222 & ~x250 & ~x332 & ~x333 & ~x416 & ~x461 & ~x504 & ~x533 & ~x555 & ~x610 & ~x617 & ~x637 & ~x645 & ~x664 & ~x668 & ~x671 & ~x696 & ~x722 & ~x759 & ~x782;
assign c889 =  x465 &  x492 &  x518 &  x519 &  x520 &  x546 & ~x56 & ~x80 & ~x87 & ~x111 & ~x114 & ~x143 & ~x224 & ~x251 & ~x281 & ~x288 & ~x289 & ~x306 & ~x315 & ~x332 & ~x341 & ~x342 & ~x343 & ~x419 & ~x473 & ~x478 & ~x663 & ~x670 & ~x685 & ~x686 & ~x687 & ~x692 & ~x698 & ~x703 & ~x730 & ~x742 & ~x747 & ~x760;
assign c891 = ~x0 & ~x2 & ~x4 & ~x6 & ~x7 & ~x8 & ~x9 & ~x12 & ~x15 & ~x18 & ~x19 & ~x21 & ~x29 & ~x31 & ~x37 & ~x38 & ~x40 & ~x43 & ~x45 & ~x50 & ~x54 & ~x56 & ~x58 & ~x67 & ~x72 & ~x78 & ~x82 & ~x83 & ~x90 & ~x92 & ~x95 & ~x102 & ~x103 & ~x104 & ~x112 & ~x118 & ~x119 & ~x134 & ~x135 & ~x136 & ~x139 & ~x166 & ~x168 & ~x171 & ~x193 & ~x194 & ~x196 & ~x198 & ~x199 & ~x221 & ~x226 & ~x279 & ~x280 & ~x336 & ~x363 & ~x364 & ~x366 & ~x377 & ~x378 & ~x392 & ~x402 & ~x403 & ~x405 & ~x420 & ~x422 & ~x430 & ~x448 & ~x475 & ~x476 & ~x478 & ~x503 & ~x505 & ~x507 & ~x535 & ~x561 & ~x589 & ~x590 & ~x648 & ~x696 & ~x718 & ~x723 & ~x724 & ~x728 & ~x730 & ~x734 & ~x746 & ~x748 & ~x752 & ~x754 & ~x755 & ~x759 & ~x766 & ~x771 & ~x772 & ~x777;
assign c893 = ~x1 & ~x4 & ~x7 & ~x23 & ~x30 & ~x34 & ~x35 & ~x38 & ~x42 & ~x49 & ~x51 & ~x54 & ~x59 & ~x63 & ~x65 & ~x66 & ~x91 & ~x92 & ~x106 & ~x141 & ~x149 & ~x167 & ~x170 & ~x204 & ~x224 & ~x226 & ~x228 & ~x231 & ~x254 & ~x257 & ~x279 & ~x283 & ~x312 & ~x314 & ~x330 & ~x340 & ~x358 & ~x360 & ~x362 & ~x389 & ~x391 & ~x419 & ~x421 & ~x445 & ~x472 & ~x473 & ~x478 & ~x504 & ~x506 & ~x532 & ~x589 & ~x590 & ~x613 & ~x615 & ~x625 & ~x630 & ~x646 & ~x652 & ~x653 & ~x658 & ~x668 & ~x680 & ~x684 & ~x686 & ~x694 & ~x700 & ~x707 & ~x708 & ~x709 & ~x721 & ~x722 & ~x728 & ~x729 & ~x731 & ~x735 & ~x737 & ~x756 & ~x760 & ~x762 & ~x768 & ~x769 & ~x772 & ~x782;
assign c895 = ~x4 & ~x13 & ~x26 & ~x34 & ~x40 & ~x44 & ~x47 & ~x58 & ~x64 & ~x78 & ~x82 & ~x87 & ~x145 & ~x169 & ~x221 & ~x226 & ~x249 & ~x250 & ~x260 & ~x261 & ~x277 & ~x283 & ~x312 & ~x316 & ~x326 & ~x331 & ~x337 & ~x343 & ~x356 & ~x361 & ~x362 & ~x369 & ~x385 & ~x449 & ~x475 & ~x479 & ~x480 & ~x508 & ~x509 & ~x536 & ~x559 & ~x587 & ~x614 & ~x654 & ~x656 & ~x663 & ~x669 & ~x671 & ~x686 & ~x713 & ~x727 & ~x735 & ~x747 & ~x753 & ~x760 & ~x765 & ~x779;
assign c897 =  x376 & ~x17 & ~x62 & ~x67 & ~x80 & ~x289 & ~x334 & ~x343 & ~x360 & ~x474 & ~x478 & ~x483 & ~x485 & ~x515 & ~x752 & ~x760 & ~x765 & ~x777;
assign c899 =  x441 & ~x51 & ~x82 & ~x141 & ~x284 & ~x361 & ~x562 & ~x594 & ~x670 & ~x704 & ~x738;
assign c8101 =  x434 &  x463 &  x491 &  x518 & ~x26 & ~x46 & ~x51 & ~x57 & ~x61 & ~x75 & ~x81 & ~x89 & ~x94 & ~x110 & ~x129 & ~x159 & ~x201 & ~x332 & ~x363 & ~x395 & ~x424 & ~x474 & ~x533 & ~x535 & ~x537 & ~x540 & ~x542 & ~x551 & ~x570 & ~x578 & ~x634 & ~x663 & ~x693 & ~x723;
assign c8103 = ~x0 & ~x4 & ~x14 & ~x15 & ~x18 & ~x21 & ~x23 & ~x24 & ~x28 & ~x29 & ~x34 & ~x35 & ~x37 & ~x38 & ~x40 & ~x44 & ~x49 & ~x54 & ~x57 & ~x64 & ~x66 & ~x70 & ~x77 & ~x80 & ~x81 & ~x82 & ~x85 & ~x89 & ~x94 & ~x111 & ~x112 & ~x122 & ~x135 & ~x142 & ~x169 & ~x192 & ~x194 & ~x196 & ~x197 & ~x201 & ~x222 & ~x223 & ~x224 & ~x249 & ~x276 & ~x278 & ~x281 & ~x282 & ~x304 & ~x322 & ~x340 & ~x348 & ~x349 & ~x365 & ~x367 & ~x369 & ~x375 & ~x376 & ~x394 & ~x402 & ~x403 & ~x420 & ~x450 & ~x529 & ~x532 & ~x534 & ~x590 & ~x616 & ~x645 & ~x668 & ~x669 & ~x672 & ~x674 & ~x686 & ~x689 & ~x690 & ~x721 & ~x728 & ~x729 & ~x730 & ~x731 & ~x732 & ~x742 & ~x747 & ~x748 & ~x749 & ~x751 & ~x753 & ~x754 & ~x756 & ~x759 & ~x764 & ~x766 & ~x770 & ~x771 & ~x776;
assign c8105 =  x649;
assign c8107 =  x409 &  x436 &  x437 & ~x14 & ~x22 & ~x25 & ~x38 & ~x41 & ~x43 & ~x46 & ~x50 & ~x51 & ~x52 & ~x71 & ~x72 & ~x73 & ~x76 & ~x80 & ~x89 & ~x90 & ~x101 & ~x103 & ~x109 & ~x115 & ~x117 & ~x120 & ~x121 & ~x128 & ~x129 & ~x130 & ~x131 & ~x132 & ~x138 & ~x140 & ~x141 & ~x144 & ~x145 & ~x153 & ~x156 & ~x161 & ~x163 & ~x166 & ~x194 & ~x197 & ~x278 & ~x279 & ~x307 & ~x309 & ~x335 & ~x360 & ~x364 & ~x387 & ~x393 & ~x416 & ~x422 & ~x423 & ~x448 & ~x475 & ~x477 & ~x500 & ~x506 & ~x510 & ~x529 & ~x531 & ~x540 & ~x558 & ~x564 & ~x568 & ~x583 & ~x588 & ~x589 & ~x590 & ~x609 & ~x612 & ~x613 & ~x616 & ~x620 & ~x621 & ~x635 & ~x644 & ~x674 & ~x723 & ~x733 & ~x756 & ~x758 & ~x762 & ~x766 & ~x772 & ~x774 & ~x781 & ~x783;
assign c8109 =  x469 &  x523 &  x524 & ~x19 & ~x30 & ~x71 & ~x134 & ~x162 & ~x166 & ~x225 & ~x364 & ~x480 & ~x733 & ~x758;
assign c8111 =  x577 &  x578 &  x603 & ~x10 & ~x44 & ~x56 & ~x96 & ~x104 & ~x113 & ~x195 & ~x196 & ~x317 & ~x330 & ~x343 & ~x362 & ~x370 & ~x371 & ~x397 & ~x477 & ~x493 & ~x502 & ~x503 & ~x586 & ~x612 & ~x614 & ~x617 & ~x640 & ~x674 & ~x689 & ~x733 & ~x767 & ~x780;
assign c8113 = ~x12 & ~x15 & ~x16 & ~x37 & ~x43 & ~x53 & ~x55 & ~x63 & ~x65 & ~x75 & ~x78 & ~x89 & ~x90 & ~x122 & ~x123 & ~x124 & ~x126 & ~x140 & ~x151 & ~x156 & ~x157 & ~x169 & ~x175 & ~x282 & ~x306 & ~x307 & ~x335 & ~x365 & ~x390 & ~x500 & ~x513 & ~x514 & ~x516 & ~x559 & ~x587 & ~x589 & ~x665 & ~x667 & ~x668 & ~x688 & ~x701 & ~x718 & ~x724 & ~x725 & ~x760 & ~x779 & ~x780 & ~x781;
assign c8115 = ~x5 & ~x14 & ~x16 & ~x18 & ~x27 & ~x32 & ~x38 & ~x46 & ~x48 & ~x49 & ~x52 & ~x54 & ~x56 & ~x59 & ~x60 & ~x62 & ~x65 & ~x78 & ~x103 & ~x110 & ~x116 & ~x118 & ~x123 & ~x155 & ~x156 & ~x166 & ~x168 & ~x193 & ~x194 & ~x196 & ~x200 & ~x252 & ~x254 & ~x279 & ~x280 & ~x281 & ~x284 & ~x309 & ~x332 & ~x395 & ~x449 & ~x501 & ~x529 & ~x532 & ~x536 & ~x537 & ~x538 & ~x559 & ~x564 & ~x567 & ~x575 & ~x577 & ~x586 & ~x590 & ~x621 & ~x630 & ~x631 & ~x642 & ~x645 & ~x646 & ~x647 & ~x648 & ~x660 & ~x661 & ~x687 & ~x696 & ~x697 & ~x699 & ~x724 & ~x725 & ~x729 & ~x742 & ~x745 & ~x746 & ~x751 & ~x754 & ~x756 & ~x761 & ~x765 & ~x767 & ~x768 & ~x770 & ~x773 & ~x777 & ~x778 & ~x782;
assign c8117 =  x543 & ~x449 & ~x533 & ~x656 & ~x658 & ~x659 & ~x682 & ~x688;
assign c8119 =  x175 & ~x291 & ~x318;
assign c8121 = ~x7 & ~x15 & ~x25 & ~x42 & ~x43 & ~x46 & ~x50 & ~x57 & ~x61 & ~x66 & ~x93 & ~x102 & ~x109 & ~x138 & ~x198 & ~x222 & ~x225 & ~x248 & ~x251 & ~x252 & ~x276 & ~x281 & ~x282 & ~x304 & ~x306 & ~x332 & ~x336 & ~x358 & ~x365 & ~x394 & ~x395 & ~x396 & ~x422 & ~x424 & ~x447 & ~x474 & ~x475 & ~x479 & ~x482 & ~x485 & ~x486 & ~x488 & ~x490 & ~x506 & ~x514 & ~x517 & ~x529 & ~x587 & ~x642 & ~x667 & ~x669 & ~x672 & ~x674 & ~x695 & ~x699 & ~x700 & ~x719 & ~x725 & ~x726 & ~x730 & ~x734 & ~x743 & ~x748 & ~x754 & ~x765 & ~x776;
assign c8123 =  x574 & ~x4 & ~x13 & ~x15 & ~x20 & ~x28 & ~x33 & ~x42 & ~x46 & ~x57 & ~x61 & ~x66 & ~x74 & ~x82 & ~x88 & ~x105 & ~x130 & ~x131 & ~x140 & ~x142 & ~x157 & ~x165 & ~x166 & ~x187 & ~x251 & ~x283 & ~x306 & ~x308 & ~x361 & ~x368 & ~x390 & ~x420 & ~x421 & ~x475 & ~x476 & ~x530 & ~x531 & ~x590 & ~x608 & ~x615 & ~x617 & ~x620 & ~x623 & ~x626 & ~x653 & ~x664 & ~x665 & ~x673 & ~x676 & ~x677 & ~x680 & ~x690 & ~x692 & ~x694 & ~x695 & ~x727 & ~x746 & ~x751 & ~x752 & ~x762 & ~x765 & ~x772 & ~x777 & ~x779;
assign c8125 =  x241 &  x296 &  x323 &  x351 &  x352 &  x379 &  x380 &  x406 & ~x5 & ~x11 & ~x24 & ~x38 & ~x42 & ~x44 & ~x56 & ~x59 & ~x87 & ~x94 & ~x168 & ~x199 & ~x225 & ~x247 & ~x251 & ~x252 & ~x333 & ~x335 & ~x362 & ~x391 & ~x397 & ~x454 & ~x471 & ~x476 & ~x480 & ~x484 & ~x494 & ~x506 & ~x509 & ~x521 & ~x526 & ~x537 & ~x558 & ~x614 & ~x618 & ~x641 & ~x695 & ~x702 & ~x705 & ~x724 & ~x725 & ~x739 & ~x751 & ~x757 & ~x772 & ~x775;
assign c8127 = ~x3 & ~x15 & ~x44 & ~x48 & ~x70 & ~x80 & ~x86 & ~x88 & ~x99 & ~x102 & ~x120 & ~x127 & ~x130 & ~x136 & ~x164 & ~x191 & ~x282 & ~x340 & ~x388 & ~x395 & ~x418 & ~x419 & ~x506 & ~x563 & ~x571 & ~x579 & ~x584 & ~x588 & ~x596 & ~x598 & ~x610 & ~x615 & ~x617 & ~x622 & ~x623 & ~x626 & ~x644 & ~x653 & ~x665 & ~x669 & ~x701 & ~x705 & ~x747 & ~x752 & ~x776 & ~x779;
assign c8129 =  x353 &  x381 & ~x17 & ~x24 & ~x50 & ~x72 & ~x105 & ~x106 & ~x116 & ~x183 & ~x197 & ~x220 & ~x275 & ~x334 & ~x363 & ~x449 & ~x554 & ~x557 & ~x560 & ~x561 & ~x618 & ~x639 & ~x648 & ~x661 & ~x674 & ~x676 & ~x689 & ~x701 & ~x757 & ~x760 & ~x767 & ~x770 & ~x775 & ~x782;
assign c8131 = ~x1 & ~x2 & ~x11 & ~x19 & ~x26 & ~x45 & ~x50 & ~x56 & ~x69 & ~x110 & ~x118 & ~x122 & ~x123 & ~x132 & ~x145 & ~x151 & ~x157 & ~x158 & ~x165 & ~x173 & ~x174 & ~x179 & ~x193 & ~x254 & ~x279 & ~x308 & ~x311 & ~x339 & ~x449 & ~x458 & ~x459 & ~x480 & ~x527 & ~x533 & ~x549 & ~x591 & ~x594 & ~x615 & ~x636 & ~x637 & ~x664 & ~x697 & ~x744 & ~x745 & ~x747 & ~x748 & ~x749 & ~x771 & ~x774 & ~x776;
assign c8133 = ~x7 & ~x18 & ~x20 & ~x72 & ~x114 & ~x153 & ~x166 & ~x168 & ~x282 & ~x312 & ~x333 & ~x394 & ~x419 & ~x446 & ~x561 & ~x566 & ~x594 & ~x601 & ~x602 & ~x630 & ~x632 & ~x640 & ~x645 & ~x657 & ~x686 & ~x689 & ~x697 & ~x739 & ~x756 & ~x763;
assign c8135 =  x466 & ~x5 & ~x6 & ~x7 & ~x8 & ~x12 & ~x15 & ~x17 & ~x25 & ~x28 & ~x29 & ~x31 & ~x36 & ~x50 & ~x60 & ~x67 & ~x68 & ~x71 & ~x72 & ~x90 & ~x91 & ~x113 & ~x117 & ~x136 & ~x137 & ~x139 & ~x142 & ~x143 & ~x144 & ~x162 & ~x166 & ~x172 & ~x191 & ~x195 & ~x202 & ~x222 & ~x223 & ~x228 & ~x230 & ~x250 & ~x255 & ~x280 & ~x281 & ~x283 & ~x302 & ~x306 & ~x312 & ~x322 & ~x323 & ~x330 & ~x332 & ~x334 & ~x336 & ~x337 & ~x338 & ~x358 & ~x365 & ~x366 & ~x392 & ~x393 & ~x416 & ~x417 & ~x421 & ~x447 & ~x450 & ~x474 & ~x475 & ~x500 & ~x501 & ~x507 & ~x531 & ~x533 & ~x535 & ~x559 & ~x561 & ~x563 & ~x564 & ~x585 & ~x614 & ~x618 & ~x619 & ~x639 & ~x644 & ~x645 & ~x666 & ~x669 & ~x674 & ~x677 & ~x680 & ~x693 & ~x706 & ~x722 & ~x723 & ~x724 & ~x725 & ~x727 & ~x729 & ~x730 & ~x738 & ~x739 & ~x747 & ~x763 & ~x769 & ~x779 & ~x782;
assign c8137 =  x710 & ~x513 & ~x542;
assign c8139 =  x210 &  x552 & ~x18 & ~x33 & ~x46 & ~x62 & ~x64 & ~x76 & ~x105 & ~x131 & ~x168 & ~x199 & ~x432 & ~x462 & ~x473 & ~x588 & ~x590 & ~x642 & ~x728 & ~x760;
assign c8141 = ~x2 & ~x4 & ~x6 & ~x7 & ~x10 & ~x12 & ~x13 & ~x14 & ~x15 & ~x17 & ~x20 & ~x22 & ~x23 & ~x24 & ~x28 & ~x32 & ~x36 & ~x45 & ~x46 & ~x55 & ~x56 & ~x57 & ~x58 & ~x63 & ~x78 & ~x79 & ~x80 & ~x85 & ~x87 & ~x88 & ~x107 & ~x114 & ~x133 & ~x135 & ~x141 & ~x142 & ~x144 & ~x145 & ~x162 & ~x165 & ~x168 & ~x171 & ~x172 & ~x173 & ~x194 & ~x195 & ~x196 & ~x199 & ~x200 & ~x201 & ~x219 & ~x225 & ~x226 & ~x227 & ~x245 & ~x246 & ~x249 & ~x252 & ~x253 & ~x255 & ~x273 & ~x274 & ~x275 & ~x278 & ~x280 & ~x281 & ~x283 & ~x284 & ~x301 & ~x302 & ~x306 & ~x329 & ~x331 & ~x335 & ~x336 & ~x340 & ~x367 & ~x391 & ~x392 & ~x394 & ~x397 & ~x420 & ~x421 & ~x423 & ~x424 & ~x446 & ~x447 & ~x448 & ~x449 & ~x451 & ~x476 & ~x478 & ~x479 & ~x503 & ~x504 & ~x506 & ~x508 & ~x531 & ~x558 & ~x562 & ~x587 & ~x588 & ~x590 & ~x615 & ~x618 & ~x620 & ~x631 & ~x632 & ~x644 & ~x645 & ~x646 & ~x648 & ~x657 & ~x658 & ~x659 & ~x660 & ~x662 & ~x669 & ~x671 & ~x672 & ~x673 & ~x685 & ~x686 & ~x688 & ~x689 & ~x690 & ~x692 & ~x700 & ~x701 & ~x705 & ~x706 & ~x714 & ~x717 & ~x718 & ~x719 & ~x728 & ~x729 & ~x733 & ~x735 & ~x736 & ~x737 & ~x739 & ~x742 & ~x743 & ~x753 & ~x754 & ~x764 & ~x765 & ~x766 & ~x769 & ~x775 & ~x776 & ~x778 & ~x780 & ~x781;
assign c8143 = ~x1 & ~x2 & ~x12 & ~x17 & ~x18 & ~x23 & ~x26 & ~x36 & ~x40 & ~x41 & ~x42 & ~x43 & ~x44 & ~x46 & ~x47 & ~x51 & ~x52 & ~x55 & ~x61 & ~x63 & ~x65 & ~x68 & ~x75 & ~x77 & ~x86 & ~x89 & ~x92 & ~x95 & ~x105 & ~x106 & ~x110 & ~x119 & ~x134 & ~x138 & ~x143 & ~x145 & ~x161 & ~x168 & ~x198 & ~x224 & ~x251 & ~x252 & ~x257 & ~x259 & ~x281 & ~x287 & ~x310 & ~x334 & ~x341 & ~x364 & ~x368 & ~x387 & ~x393 & ~x395 & ~x420 & ~x421 & ~x442 & ~x444 & ~x448 & ~x455 & ~x474 & ~x476 & ~x485 & ~x486 & ~x488 & ~x499 & ~x504 & ~x527 & ~x533 & ~x534 & ~x562 & ~x563 & ~x564 & ~x585 & ~x586 & ~x588 & ~x616 & ~x617 & ~x619 & ~x638 & ~x644 & ~x645 & ~x647 & ~x662 & ~x664 & ~x668 & ~x673 & ~x687 & ~x688 & ~x690 & ~x691 & ~x693 & ~x696 & ~x700 & ~x719 & ~x730 & ~x732 & ~x733 & ~x735 & ~x740 & ~x741 & ~x744 & ~x755 & ~x763 & ~x779;
assign c8145 = ~x14 & ~x15 & ~x24 & ~x31 & ~x36 & ~x41 & ~x47 & ~x54 & ~x56 & ~x69 & ~x70 & ~x109 & ~x115 & ~x143 & ~x167 & ~x199 & ~x224 & ~x227 & ~x248 & ~x249 & ~x265 & ~x277 & ~x281 & ~x293 & ~x301 & ~x312 & ~x320 & ~x336 & ~x347 & ~x361 & ~x375 & ~x390 & ~x392 & ~x400 & ~x401 & ~x402 & ~x421 & ~x424 & ~x446 & ~x452 & ~x500 & ~x506 & ~x557 & ~x561 & ~x585 & ~x587 & ~x647 & ~x671 & ~x699 & ~x718 & ~x736 & ~x739 & ~x742 & ~x745 & ~x746 & ~x750 & ~x752 & ~x759 & ~x764 & ~x768 & ~x769 & ~x770 & ~x776;
assign c8147 =  x521 & ~x0 & ~x16 & ~x21 & ~x25 & ~x43 & ~x50 & ~x57 & ~x58 & ~x61 & ~x66 & ~x85 & ~x106 & ~x107 & ~x137 & ~x199 & ~x202 & ~x225 & ~x230 & ~x232 & ~x251 & ~x252 & ~x253 & ~x260 & ~x278 & ~x304 & ~x337 & ~x368 & ~x379 & ~x391 & ~x445 & ~x533 & ~x591 & ~x634 & ~x635 & ~x640 & ~x641 & ~x642 & ~x663 & ~x708 & ~x716 & ~x724 & ~x727 & ~x732 & ~x741 & ~x749 & ~x751 & ~x753 & ~x759 & ~x763 & ~x777;
assign c8149 =  x494 &  x521 &  x576 & ~x25 & ~x41 & ~x48 & ~x52 & ~x56 & ~x70 & ~x86 & ~x134 & ~x135 & ~x137 & ~x141 & ~x142 & ~x166 & ~x172 & ~x336 & ~x351 & ~x388 & ~x416 & ~x445 & ~x447 & ~x478 & ~x557 & ~x613 & ~x619 & ~x645 & ~x646 & ~x667 & ~x732 & ~x779 & ~x782;
assign c8151 =  x522 &  x524 &  x548 & ~x2 & ~x19 & ~x43 & ~x54 & ~x58 & ~x90 & ~x136 & ~x140 & ~x164 & ~x220 & ~x226 & ~x227 & ~x252 & ~x254 & ~x280 & ~x283 & ~x311 & ~x391 & ~x476 & ~x477 & ~x478 & ~x504 & ~x591 & ~x635 & ~x636 & ~x643 & ~x662 & ~x663 & ~x696 & ~x720 & ~x749 & ~x761 & ~x763 & ~x769 & ~x771 & ~x779;
assign c8153 =  x354 &  x438 &  x493 &  x520 & ~x4 & ~x16 & ~x25 & ~x32 & ~x34 & ~x58 & ~x61 & ~x70 & ~x82 & ~x84 & ~x107 & ~x109 & ~x124 & ~x141 & ~x145 & ~x172 & ~x222 & ~x223 & ~x246 & ~x276 & ~x307 & ~x366 & ~x395 & ~x450 & ~x561 & ~x582 & ~x587 & ~x589 & ~x615 & ~x616 & ~x620 & ~x665 & ~x674 & ~x676 & ~x738 & ~x748 & ~x754 & ~x755 & ~x759 & ~x765 & ~x771 & ~x781;
assign c8155 = ~x0 & ~x2 & ~x5 & ~x8 & ~x9 & ~x17 & ~x22 & ~x23 & ~x27 & ~x34 & ~x47 & ~x51 & ~x53 & ~x55 & ~x62 & ~x64 & ~x67 & ~x68 & ~x69 & ~x70 & ~x73 & ~x75 & ~x82 & ~x84 & ~x87 & ~x92 & ~x93 & ~x97 & ~x100 & ~x101 & ~x102 & ~x106 & ~x109 & ~x111 & ~x121 & ~x138 & ~x169 & ~x195 & ~x196 & ~x222 & ~x224 & ~x226 & ~x249 & ~x253 & ~x276 & ~x277 & ~x281 & ~x303 & ~x304 & ~x305 & ~x306 & ~x310 & ~x333 & ~x337 & ~x359 & ~x363 & ~x386 & ~x390 & ~x414 & ~x418 & ~x445 & ~x448 & ~x450 & ~x474 & ~x476 & ~x478 & ~x481 & ~x482 & ~x483 & ~x501 & ~x512 & ~x531 & ~x532 & ~x533 & ~x541 & ~x542 & ~x543 & ~x544 & ~x546 & ~x555 & ~x557 & ~x561 & ~x583 & ~x589 & ~x613 & ~x614 & ~x615 & ~x616 & ~x642 & ~x669 & ~x675 & ~x696 & ~x701 & ~x703 & ~x708 & ~x723 & ~x724 & ~x727 & ~x730 & ~x733 & ~x737 & ~x740 & ~x741 & ~x758 & ~x776 & ~x779 & ~x780 & ~x783;
assign c8157 =  x266 & ~x142 & ~x149 & ~x157 & ~x206 & ~x456 & ~x514 & ~x542 & ~x671 & ~x695 & ~x699 & ~x759;
assign c8159 =  x466 &  x494 &  x548 & ~x0 & ~x1 & ~x18 & ~x21 & ~x26 & ~x27 & ~x31 & ~x41 & ~x42 & ~x45 & ~x51 & ~x52 & ~x54 & ~x55 & ~x60 & ~x64 & ~x66 & ~x67 & ~x72 & ~x73 & ~x74 & ~x75 & ~x76 & ~x78 & ~x79 & ~x80 & ~x81 & ~x82 & ~x84 & ~x85 & ~x90 & ~x91 & ~x92 & ~x115 & ~x135 & ~x142 & ~x144 & ~x145 & ~x147 & ~x162 & ~x169 & ~x192 & ~x196 & ~x197 & ~x199 & ~x220 & ~x222 & ~x223 & ~x224 & ~x228 & ~x229 & ~x248 & ~x277 & ~x303 & ~x307 & ~x308 & ~x312 & ~x363 & ~x364 & ~x365 & ~x388 & ~x389 & ~x390 & ~x423 & ~x446 & ~x473 & ~x475 & ~x478 & ~x480 & ~x503 & ~x528 & ~x534 & ~x554 & ~x560 & ~x561 & ~x581 & ~x585 & ~x586 & ~x593 & ~x594 & ~x609 & ~x610 & ~x638 & ~x639 & ~x640 & ~x665 & ~x672 & ~x676 & ~x677 & ~x680 & ~x696 & ~x700 & ~x704 & ~x705 & ~x707 & ~x709 & ~x722 & ~x723 & ~x726 & ~x728 & ~x729 & ~x731 & ~x742 & ~x743 & ~x749 & ~x750 & ~x751 & ~x754 & ~x759 & ~x760 & ~x763 & ~x765;
assign c8161 =  x569 &  x600 & ~x13 & ~x14 & ~x16 & ~x21 & ~x22 & ~x27 & ~x31 & ~x41 & ~x42 & ~x47 & ~x52 & ~x69 & ~x82 & ~x83 & ~x84 & ~x112 & ~x139 & ~x142 & ~x167 & ~x169 & ~x194 & ~x199 & ~x201 & ~x225 & ~x230 & ~x231 & ~x280 & ~x283 & ~x284 & ~x285 & ~x302 & ~x307 & ~x311 & ~x334 & ~x339 & ~x340 & ~x359 & ~x361 & ~x364 & ~x392 & ~x394 & ~x395 & ~x423 & ~x449 & ~x452 & ~x487 & ~x528 & ~x530 & ~x533 & ~x534 & ~x560 & ~x585 & ~x588 & ~x610 & ~x639 & ~x640 & ~x646 & ~x671 & ~x694 & ~x720 & ~x721 & ~x729 & ~x737 & ~x749 & ~x756 & ~x761 & ~x765 & ~x772 & ~x780;
assign c8163 =  x382 &  x410 &  x465 & ~x5 & ~x6 & ~x8 & ~x9 & ~x10 & ~x18 & ~x21 & ~x25 & ~x31 & ~x38 & ~x54 & ~x89 & ~x93 & ~x125 & ~x140 & ~x142 & ~x152 & ~x170 & ~x194 & ~x196 & ~x197 & ~x305 & ~x333 & ~x336 & ~x359 & ~x416 & ~x447 & ~x474 & ~x556 & ~x557 & ~x568 & ~x592 & ~x610 & ~x613 & ~x616 & ~x638 & ~x639 & ~x672 & ~x688 & ~x716 & ~x723 & ~x725 & ~x732 & ~x734 & ~x745 & ~x746 & ~x754 & ~x769 & ~x776;
assign c8165 =  x319 & ~x4 & ~x10 & ~x11 & ~x20 & ~x29 & ~x30 & ~x31 & ~x34 & ~x35 & ~x36 & ~x43 & ~x44 & ~x45 & ~x48 & ~x51 & ~x53 & ~x55 & ~x69 & ~x79 & ~x85 & ~x86 & ~x106 & ~x109 & ~x112 & ~x115 & ~x118 & ~x134 & ~x137 & ~x140 & ~x146 & ~x166 & ~x170 & ~x171 & ~x195 & ~x198 & ~x225 & ~x226 & ~x256 & ~x259 & ~x365 & ~x392 & ~x393 & ~x395 & ~x418 & ~x423 & ~x433 & ~x434 & ~x446 & ~x447 & ~x448 & ~x460 & ~x462 & ~x475 & ~x477 & ~x479 & ~x505 & ~x528 & ~x530 & ~x531 & ~x559 & ~x563 & ~x584 & ~x586 & ~x610 & ~x620 & ~x640 & ~x645 & ~x647 & ~x668 & ~x673 & ~x677 & ~x706 & ~x719 & ~x722 & ~x733 & ~x744 & ~x745 & ~x748 & ~x749 & ~x751 & ~x758 & ~x763 & ~x764 & ~x765 & ~x771 & ~x776;
assign c8167 =  x501;
assign c8169 =  x429 & ~x2 & ~x5 & ~x8 & ~x12 & ~x19 & ~x23 & ~x25 & ~x28 & ~x30 & ~x32 & ~x42 & ~x45 & ~x49 & ~x59 & ~x76 & ~x83 & ~x109 & ~x110 & ~x131 & ~x141 & ~x156 & ~x157 & ~x197 & ~x198 & ~x226 & ~x278 & ~x280 & ~x284 & ~x304 & ~x306 & ~x333 & ~x336 & ~x337 & ~x363 & ~x365 & ~x368 & ~x389 & ~x394 & ~x419 & ~x447 & ~x448 & ~x477 & ~x480 & ~x503 & ~x508 & ~x532 & ~x535 & ~x556 & ~x560 & ~x562 & ~x584 & ~x588 & ~x589 & ~x590 & ~x591 & ~x594 & ~x597 & ~x614 & ~x617 & ~x621 & ~x623 & ~x625 & ~x638 & ~x641 & ~x642 & ~x645 & ~x646 & ~x674 & ~x696 & ~x702 & ~x705 & ~x724 & ~x726 & ~x727 & ~x730 & ~x753 & ~x758 & ~x760 & ~x762 & ~x770 & ~x772 & ~x775 & ~x776 & ~x778 & ~x779 & ~x783;
assign c8171 = ~x1 & ~x3 & ~x4 & ~x5 & ~x6 & ~x8 & ~x10 & ~x11 & ~x13 & ~x14 & ~x15 & ~x16 & ~x18 & ~x20 & ~x21 & ~x27 & ~x29 & ~x30 & ~x31 & ~x32 & ~x34 & ~x36 & ~x37 & ~x38 & ~x44 & ~x46 & ~x51 & ~x54 & ~x55 & ~x57 & ~x58 & ~x64 & ~x66 & ~x76 & ~x78 & ~x79 & ~x80 & ~x82 & ~x83 & ~x86 & ~x87 & ~x89 & ~x90 & ~x91 & ~x92 & ~x94 & ~x107 & ~x110 & ~x116 & ~x118 & ~x140 & ~x142 & ~x144 & ~x145 & ~x165 & ~x166 & ~x168 & ~x169 & ~x191 & ~x192 & ~x194 & ~x198 & ~x199 & ~x222 & ~x251 & ~x252 & ~x254 & ~x275 & ~x277 & ~x282 & ~x283 & ~x284 & ~x303 & ~x305 & ~x308 & ~x310 & ~x331 & ~x332 & ~x336 & ~x339 & ~x360 & ~x364 & ~x388 & ~x389 & ~x390 & ~x391 & ~x394 & ~x417 & ~x420 & ~x447 & ~x448 & ~x472 & ~x474 & ~x502 & ~x505 & ~x506 & ~x530 & ~x531 & ~x533 & ~x534 & ~x558 & ~x561 & ~x587 & ~x588 & ~x589 & ~x613 & ~x615 & ~x616 & ~x617 & ~x618 & ~x629 & ~x630 & ~x631 & ~x632 & ~x633 & ~x643 & ~x657 & ~x658 & ~x660 & ~x661 & ~x672 & ~x673 & ~x674 & ~x687 & ~x688 & ~x689 & ~x690 & ~x691 & ~x705 & ~x715 & ~x716 & ~x727 & ~x730 & ~x734 & ~x737 & ~x738 & ~x742 & ~x744 & ~x748 & ~x749 & ~x751 & ~x754 & ~x755 & ~x758 & ~x759 & ~x761 & ~x763 & ~x768 & ~x772 & ~x773 & ~x774 & ~x779 & ~x782 & ~x783;
assign c8173 = ~x2 & ~x3 & ~x9 & ~x11 & ~x18 & ~x24 & ~x25 & ~x27 & ~x28 & ~x31 & ~x39 & ~x46 & ~x49 & ~x51 & ~x57 & ~x58 & ~x62 & ~x63 & ~x66 & ~x70 & ~x71 & ~x75 & ~x83 & ~x91 & ~x96 & ~x97 & ~x99 & ~x107 & ~x108 & ~x116 & ~x118 & ~x139 & ~x166 & ~x170 & ~x224 & ~x249 & ~x253 & ~x277 & ~x279 & ~x283 & ~x312 & ~x362 & ~x365 & ~x386 & ~x387 & ~x414 & ~x416 & ~x422 & ~x423 & ~x424 & ~x449 & ~x451 & ~x474 & ~x476 & ~x478 & ~x483 & ~x488 & ~x489 & ~x509 & ~x510 & ~x512 & ~x513 & ~x515 & ~x516 & ~x529 & ~x535 & ~x557 & ~x561 & ~x563 & ~x565 & ~x582 & ~x586 & ~x614 & ~x616 & ~x617 & ~x636 & ~x645 & ~x665 & ~x667 & ~x669 & ~x692 & ~x694 & ~x695 & ~x698 & ~x726 & ~x755 & ~x760 & ~x762 & ~x766 & ~x768 & ~x773;
assign c8175 =  x544 & ~x9 & ~x12 & ~x21 & ~x23 & ~x32 & ~x38 & ~x40 & ~x51 & ~x58 & ~x59 & ~x79 & ~x81 & ~x86 & ~x92 & ~x108 & ~x111 & ~x117 & ~x142 & ~x164 & ~x196 & ~x228 & ~x252 & ~x276 & ~x280 & ~x281 & ~x304 & ~x310 & ~x314 & ~x322 & ~x331 & ~x332 & ~x340 & ~x367 & ~x392 & ~x393 & ~x478 & ~x532 & ~x613 & ~x615 & ~x617 & ~x640 & ~x656 & ~x660 & ~x675 & ~x684 & ~x685 & ~x686 & ~x690 & ~x692 & ~x694 & ~x696 & ~x700 & ~x713 & ~x715 & ~x724 & ~x728 & ~x731 & ~x744 & ~x746 & ~x754 & ~x756 & ~x758 & ~x761 & ~x774 & ~x777 & ~x778 & ~x780 & ~x783;
assign c8177 = ~x0 & ~x3 & ~x4 & ~x11 & ~x12 & ~x16 & ~x18 & ~x21 & ~x24 & ~x29 & ~x30 & ~x38 & ~x39 & ~x41 & ~x51 & ~x53 & ~x54 & ~x55 & ~x57 & ~x58 & ~x62 & ~x69 & ~x79 & ~x82 & ~x83 & ~x89 & ~x95 & ~x97 & ~x112 & ~x139 & ~x142 & ~x145 & ~x170 & ~x254 & ~x255 & ~x284 & ~x305 & ~x309 & ~x350 & ~x351 & ~x353 & ~x354 & ~x361 & ~x367 & ~x378 & ~x379 & ~x380 & ~x381 & ~x382 & ~x383 & ~x392 & ~x394 & ~x410 & ~x419 & ~x449 & ~x474 & ~x502 & ~x503 & ~x584 & ~x591 & ~x620 & ~x640 & ~x645 & ~x668 & ~x670 & ~x671 & ~x672 & ~x677 & ~x694 & ~x698 & ~x701 & ~x703 & ~x705 & ~x706 & ~x730 & ~x732 & ~x735 & ~x736 & ~x738 & ~x742 & ~x752 & ~x754 & ~x755 & ~x756 & ~x757 & ~x774 & ~x778 & ~x780 & ~x782;
assign c8179 =  x430 &  x486 & ~x2 & ~x10 & ~x32 & ~x36 & ~x37 & ~x42 & ~x88 & ~x114 & ~x143 & ~x146 & ~x164 & ~x169 & ~x216 & ~x243 & ~x247 & ~x251 & ~x257 & ~x276 & ~x278 & ~x315 & ~x342 & ~x360 & ~x361 & ~x389 & ~x448 & ~x476 & ~x478 & ~x502 & ~x505 & ~x535 & ~x558 & ~x561 & ~x614 & ~x623 & ~x635 & ~x645 & ~x648 & ~x653 & ~x662 & ~x668 & ~x683 & ~x690 & ~x694 & ~x696 & ~x698 & ~x718 & ~x722 & ~x727 & ~x735 & ~x753 & ~x757 & ~x760 & ~x766 & ~x770 & ~x771 & ~x783;
assign c8181 =  x443;
assign c8183 =  x508;
assign c8185 =  x412 &  x467 &  x522 & ~x11 & ~x48 & ~x109 & ~x117 & ~x134 & ~x143 & ~x144 & ~x170 & ~x195 & ~x275 & ~x335 & ~x390 & ~x448 & ~x528 & ~x530 & ~x588 & ~x646 & ~x707 & ~x736 & ~x740 & ~x750 & ~x757 & ~x781;
assign c8187 =  x439 & ~x6 & ~x18 & ~x23 & ~x26 & ~x34 & ~x35 & ~x39 & ~x64 & ~x79 & ~x80 & ~x81 & ~x91 & ~x116 & ~x120 & ~x124 & ~x126 & ~x145 & ~x171 & ~x172 & ~x194 & ~x249 & ~x366 & ~x386 & ~x390 & ~x392 & ~x394 & ~x414 & ~x415 & ~x473 & ~x559 & ~x608 & ~x618 & ~x647 & ~x652 & ~x675 & ~x680 & ~x681 & ~x682 & ~x704 & ~x720 & ~x726 & ~x730 & ~x733 & ~x735 & ~x737 & ~x750 & ~x756 & ~x760 & ~x766 & ~x776 & ~x783;
assign c8189 =  x442 &  x469 & ~x446 & ~x500;
assign c8191 = ~x9 & ~x14 & ~x26 & ~x29 & ~x35 & ~x62 & ~x68 & ~x70 & ~x78 & ~x82 & ~x92 & ~x95 & ~x223 & ~x307 & ~x339 & ~x394 & ~x403 & ~x404 & ~x417 & ~x421 & ~x434 & ~x515 & ~x516 & ~x645 & ~x668 & ~x724 & ~x730 & ~x731;
assign c8193 = ~x6 & ~x7 & ~x12 & ~x16 & ~x17 & ~x19 & ~x22 & ~x37 & ~x41 & ~x42 & ~x43 & ~x50 & ~x51 & ~x56 & ~x58 & ~x59 & ~x62 & ~x66 & ~x72 & ~x78 & ~x80 & ~x84 & ~x89 & ~x93 & ~x95 & ~x96 & ~x100 & ~x102 & ~x103 & ~x110 & ~x114 & ~x115 & ~x120 & ~x121 & ~x125 & ~x126 & ~x129 & ~x134 & ~x141 & ~x143 & ~x150 & ~x154 & ~x158 & ~x182 & ~x223 & ~x252 & ~x254 & ~x279 & ~x312 & ~x334 & ~x360 & ~x365 & ~x387 & ~x393 & ~x394 & ~x419 & ~x447 & ~x476 & ~x500 & ~x503 & ~x505 & ~x534 & ~x535 & ~x536 & ~x537 & ~x541 & ~x542 & ~x543 & ~x558 & ~x562 & ~x566 & ~x567 & ~x613 & ~x618 & ~x668 & ~x671 & ~x698 & ~x700 & ~x702 & ~x703 & ~x726 & ~x730 & ~x733 & ~x750 & ~x754 & ~x763 & ~x772 & ~x773 & ~x775 & ~x778 & ~x781;
assign c8195 =  x435 & ~x9 & ~x15 & ~x17 & ~x25 & ~x78 & ~x113 & ~x122 & ~x131 & ~x136 & ~x142 & ~x157 & ~x171 & ~x200 & ~x252 & ~x254 & ~x304 & ~x369 & ~x445 & ~x477 & ~x504 & ~x565 & ~x590 & ~x591 & ~x594 & ~x597 & ~x604 & ~x613 & ~x620 & ~x623 & ~x632 & ~x633 & ~x690 & ~x699 & ~x718 & ~x730 & ~x759 & ~x772 & ~x779 & ~x780;
assign c8197 = ~x0 & ~x9 & ~x13 & ~x16 & ~x18 & ~x20 & ~x21 & ~x32 & ~x38 & ~x42 & ~x44 & ~x47 & ~x49 & ~x61 & ~x65 & ~x75 & ~x83 & ~x98 & ~x116 & ~x143 & ~x200 & ~x225 & ~x251 & ~x252 & ~x306 & ~x364 & ~x418 & ~x452 & ~x473 & ~x478 & ~x484 & ~x486 & ~x502 & ~x516 & ~x532 & ~x534 & ~x542 & ~x544 & ~x545 & ~x563 & ~x589 & ~x610 & ~x615 & ~x619 & ~x640 & ~x645 & ~x667 & ~x669 & ~x672 & ~x674 & ~x691 & ~x695 & ~x702 & ~x717 & ~x726 & ~x734 & ~x738 & ~x742 & ~x760 & ~x763 & ~x765;
assign c8199 = ~x0 & ~x5 & ~x10 & ~x11 & ~x13 & ~x14 & ~x17 & ~x18 & ~x24 & ~x27 & ~x32 & ~x44 & ~x47 & ~x49 & ~x53 & ~x56 & ~x67 & ~x68 & ~x69 & ~x75 & ~x76 & ~x80 & ~x82 & ~x84 & ~x89 & ~x95 & ~x102 & ~x104 & ~x108 & ~x109 & ~x112 & ~x117 & ~x119 & ~x135 & ~x138 & ~x142 & ~x146 & ~x224 & ~x226 & ~x249 & ~x250 & ~x251 & ~x252 & ~x278 & ~x295 & ~x303 & ~x304 & ~x306 & ~x320 & ~x321 & ~x322 & ~x333 & ~x337 & ~x338 & ~x346 & ~x347 & ~x359 & ~x362 & ~x364 & ~x374 & ~x389 & ~x392 & ~x393 & ~x401 & ~x427 & ~x428 & ~x445 & ~x446 & ~x448 & ~x503 & ~x506 & ~x642 & ~x643 & ~x644 & ~x646 & ~x667 & ~x672 & ~x699 & ~x703 & ~x720 & ~x727 & ~x730 & ~x733 & ~x734 & ~x744 & ~x746 & ~x747 & ~x749 & ~x754 & ~x758 & ~x759 & ~x761 & ~x764 & ~x765 & ~x769 & ~x777 & ~x778 & ~x781;
assign c8201 = ~x66 & ~x110 & ~x111 & ~x197 & ~x253 & ~x280 & ~x353 & ~x447 & ~x459 & ~x461 & ~x488 & ~x490 & ~x502 & ~x585 & ~x618 & ~x667 & ~x719 & ~x735 & ~x742;
assign c8203 =  x238 & ~x22 & ~x25 & ~x28 & ~x43 & ~x54 & ~x58 & ~x59 & ~x61 & ~x77 & ~x143 & ~x226 & ~x243 & ~x247 & ~x251 & ~x255 & ~x279 & ~x302 & ~x317 & ~x335 & ~x343 & ~x384 & ~x385 & ~x413 & ~x415 & ~x422 & ~x446 & ~x477 & ~x482 & ~x500 & ~x595 & ~x645 & ~x671 & ~x677 & ~x678 & ~x681 & ~x694 & ~x696 & ~x707 & ~x716 & ~x729 & ~x746 & ~x750 & ~x770 & ~x783;
assign c8205 =  x625 & ~x2 & ~x18 & ~x27 & ~x63 & ~x87 & ~x98 & ~x106 & ~x139 & ~x196 & ~x199 & ~x225 & ~x257 & ~x310 & ~x334 & ~x388 & ~x421 & ~x424 & ~x447 & ~x481 & ~x482 & ~x483 & ~x509 & ~x510 & ~x511 & ~x512 & ~x514 & ~x533 & ~x541 & ~x559 & ~x613 & ~x670 & ~x699 & ~x711 & ~x756 & ~x758;
assign c8207 = ~x6 & ~x8 & ~x15 & ~x19 & ~x20 & ~x22 & ~x26 & ~x28 & ~x30 & ~x31 & ~x32 & ~x37 & ~x38 & ~x43 & ~x47 & ~x55 & ~x56 & ~x58 & ~x71 & ~x72 & ~x76 & ~x80 & ~x84 & ~x87 & ~x97 & ~x109 & ~x111 & ~x140 & ~x141 & ~x167 & ~x225 & ~x254 & ~x283 & ~x311 & ~x330 & ~x363 & ~x367 & ~x393 & ~x395 & ~x458 & ~x459 & ~x460 & ~x461 & ~x473 & ~x483 & ~x488 & ~x489 & ~x490 & ~x517 & ~x518 & ~x529 & ~x533 & ~x559 & ~x561 & ~x562 & ~x588 & ~x612 & ~x615 & ~x666 & ~x692 & ~x696 & ~x702 & ~x716 & ~x717 & ~x718 & ~x721 & ~x725 & ~x736 & ~x740 & ~x745 & ~x753 & ~x757 & ~x772 & ~x775;
assign c8209 = ~x0 & ~x3 & ~x6 & ~x7 & ~x8 & ~x11 & ~x13 & ~x16 & ~x17 & ~x18 & ~x20 & ~x21 & ~x22 & ~x24 & ~x25 & ~x28 & ~x30 & ~x31 & ~x32 & ~x35 & ~x38 & ~x44 & ~x45 & ~x48 & ~x54 & ~x57 & ~x58 & ~x61 & ~x77 & ~x78 & ~x81 & ~x83 & ~x85 & ~x105 & ~x111 & ~x114 & ~x116 & ~x133 & ~x138 & ~x139 & ~x140 & ~x141 & ~x142 & ~x163 & ~x168 & ~x195 & ~x220 & ~x221 & ~x222 & ~x225 & ~x228 & ~x248 & ~x252 & ~x255 & ~x275 & ~x276 & ~x280 & ~x281 & ~x284 & ~x304 & ~x307 & ~x310 & ~x332 & ~x333 & ~x334 & ~x335 & ~x338 & ~x339 & ~x340 & ~x362 & ~x364 & ~x365 & ~x419 & ~x420 & ~x422 & ~x446 & ~x477 & ~x505 & ~x531 & ~x614 & ~x615 & ~x616 & ~x620 & ~x624 & ~x625 & ~x626 & ~x641 & ~x642 & ~x643 & ~x646 & ~x652 & ~x653 & ~x654 & ~x655 & ~x656 & ~x657 & ~x658 & ~x660 & ~x661 & ~x668 & ~x670 & ~x672 & ~x673 & ~x679 & ~x680 & ~x682 & ~x685 & ~x688 & ~x689 & ~x700 & ~x701 & ~x703 & ~x704 & ~x708 & ~x719 & ~x728 & ~x732 & ~x738 & ~x742 & ~x744 & ~x747 & ~x749 & ~x751 & ~x752 & ~x755 & ~x762 & ~x763 & ~x764 & ~x765 & ~x769 & ~x772 & ~x773 & ~x775 & ~x776 & ~x777 & ~x778 & ~x780 & ~x782 & ~x783;
assign c8211 =  x407 &  x518 & ~x3 & ~x7 & ~x10 & ~x12 & ~x17 & ~x19 & ~x20 & ~x23 & ~x24 & ~x34 & ~x36 & ~x38 & ~x39 & ~x40 & ~x52 & ~x53 & ~x62 & ~x67 & ~x74 & ~x85 & ~x86 & ~x87 & ~x92 & ~x94 & ~x120 & ~x132 & ~x134 & ~x138 & ~x142 & ~x146 & ~x148 & ~x159 & ~x165 & ~x167 & ~x168 & ~x174 & ~x196 & ~x200 & ~x222 & ~x225 & ~x226 & ~x304 & ~x305 & ~x308 & ~x333 & ~x366 & ~x388 & ~x419 & ~x421 & ~x442 & ~x451 & ~x475 & ~x476 & ~x508 & ~x510 & ~x529 & ~x530 & ~x539 & ~x541 & ~x562 & ~x567 & ~x577 & ~x588 & ~x594 & ~x606 & ~x614 & ~x615 & ~x616 & ~x623 & ~x635 & ~x638 & ~x643 & ~x671 & ~x674 & ~x702 & ~x703 & ~x720 & ~x722 & ~x727 & ~x730 & ~x733 & ~x737 & ~x745 & ~x748 & ~x751 & ~x762 & ~x763;
assign c8213 = ~x0 & ~x17 & ~x24 & ~x25 & ~x32 & ~x50 & ~x59 & ~x83 & ~x85 & ~x91 & ~x110 & ~x115 & ~x161 & ~x173 & ~x217 & ~x225 & ~x251 & ~x252 & ~x254 & ~x261 & ~x269 & ~x270 & ~x280 & ~x298 & ~x304 & ~x313 & ~x315 & ~x328 & ~x337 & ~x338 & ~x340 & ~x358 & ~x361 & ~x370 & ~x371 & ~x396 & ~x419 & ~x420 & ~x425 & ~x611 & ~x614 & ~x644 & ~x663 & ~x676 & ~x682 & ~x686 & ~x690 & ~x691 & ~x704 & ~x710 & ~x712 & ~x724 & ~x750 & ~x761 & ~x763 & ~x764 & ~x782;
assign c8215 = ~x5 & ~x9 & ~x18 & ~x52 & ~x75 & ~x80 & ~x110 & ~x197 & ~x302 & ~x332 & ~x336 & ~x363 & ~x392 & ~x393 & ~x415 & ~x445 & ~x476 & ~x483 & ~x511 & ~x512 & ~x513 & ~x514 & ~x515 & ~x517 & ~x532 & ~x561 & ~x584 & ~x617 & ~x647 & ~x702 & ~x704 & ~x733 & ~x766 & ~x768 & ~x781;
assign c8217 = ~x22 & ~x26 & ~x29 & ~x39 & ~x50 & ~x89 & ~x106 & ~x114 & ~x119 & ~x138 & ~x173 & ~x254 & ~x282 & ~x309 & ~x337 & ~x348 & ~x349 & ~x350 & ~x377 & ~x394 & ~x404 & ~x431 & ~x458 & ~x475 & ~x507 & ~x532 & ~x588 & ~x673 & ~x751 & ~x756 & ~x764 & ~x773;
assign c8219 = ~x7 & ~x17 & ~x22 & ~x25 & ~x27 & ~x30 & ~x50 & ~x65 & ~x66 & ~x71 & ~x76 & ~x80 & ~x86 & ~x92 & ~x98 & ~x102 & ~x104 & ~x108 & ~x110 & ~x114 & ~x117 & ~x118 & ~x119 & ~x126 & ~x132 & ~x140 & ~x146 & ~x167 & ~x196 & ~x198 & ~x202 & ~x225 & ~x227 & ~x230 & ~x251 & ~x256 & ~x258 & ~x283 & ~x335 & ~x336 & ~x363 & ~x364 & ~x387 & ~x392 & ~x415 & ~x420 & ~x421 & ~x422 & ~x448 & ~x451 & ~x452 & ~x470 & ~x472 & ~x479 & ~x507 & ~x510 & ~x511 & ~x513 & ~x514 & ~x515 & ~x516 & ~x530 & ~x532 & ~x544 & ~x552 & ~x553 & ~x557 & ~x559 & ~x562 & ~x581 & ~x585 & ~x590 & ~x611 & ~x635 & ~x639 & ~x640 & ~x641 & ~x647 & ~x669 & ~x674 & ~x694 & ~x699 & ~x703 & ~x719 & ~x722 & ~x734 & ~x773 & ~x774 & ~x776 & ~x780 & ~x781;
assign c8221 = ~x16 & ~x57 & ~x241 & ~x249 & ~x270 & ~x271 & ~x277 & ~x301 & ~x477 & ~x585 & ~x595 & ~x658 & ~x685 & ~x696;
assign c8223 =  x632 & ~x5 & ~x6 & ~x14 & ~x19 & ~x21 & ~x26 & ~x28 & ~x31 & ~x33 & ~x38 & ~x40 & ~x44 & ~x46 & ~x47 & ~x61 & ~x62 & ~x71 & ~x73 & ~x76 & ~x79 & ~x81 & ~x83 & ~x91 & ~x103 & ~x107 & ~x109 & ~x111 & ~x116 & ~x118 & ~x168 & ~x194 & ~x195 & ~x224 & ~x225 & ~x252 & ~x277 & ~x280 & ~x283 & ~x304 & ~x331 & ~x336 & ~x361 & ~x362 & ~x365 & ~x366 & ~x367 & ~x389 & ~x391 & ~x425 & ~x449 & ~x450 & ~x454 & ~x455 & ~x476 & ~x478 & ~x485 & ~x515 & ~x516 & ~x518 & ~x529 & ~x531 & ~x556 & ~x584 & ~x588 & ~x618 & ~x647 & ~x677 & ~x678 & ~x696 & ~x697 & ~x699 & ~x718 & ~x735 & ~x741 & ~x748 & ~x751 & ~x753 & ~x754 & ~x756 & ~x762 & ~x765 & ~x770 & ~x778 & ~x779;
assign c8225 =  x398 &  x399 &  x426 & ~x418 & ~x449 & ~x751 & ~x780;
assign c8227 =  x493 & ~x9 & ~x43 & ~x46 & ~x47 & ~x59 & ~x63 & ~x79 & ~x87 & ~x90 & ~x91 & ~x109 & ~x141 & ~x143 & ~x166 & ~x253 & ~x256 & ~x277 & ~x323 & ~x324 & ~x329 & ~x340 & ~x352 & ~x386 & ~x389 & ~x394 & ~x420 & ~x421 & ~x442 & ~x446 & ~x477 & ~x588 & ~x616 & ~x670 & ~x690 & ~x691 & ~x692 & ~x699 & ~x703 & ~x724 & ~x726 & ~x733 & ~x743;
assign c8229 = ~x2 & ~x11 & ~x25 & ~x26 & ~x27 & ~x36 & ~x38 & ~x40 & ~x49 & ~x54 & ~x63 & ~x64 & ~x65 & ~x70 & ~x72 & ~x79 & ~x85 & ~x94 & ~x101 & ~x110 & ~x168 & ~x171 & ~x173 & ~x251 & ~x255 & ~x310 & ~x311 & ~x331 & ~x334 & ~x337 & ~x341 & ~x369 & ~x390 & ~x391 & ~x393 & ~x397 & ~x419 & ~x424 & ~x442 & ~x443 & ~x446 & ~x447 & ~x470 & ~x483 & ~x484 & ~x486 & ~x500 & ~x502 & ~x503 & ~x506 & ~x508 & ~x516 & ~x528 & ~x545 & ~x557 & ~x583 & ~x611 & ~x615 & ~x642 & ~x666 & ~x699 & ~x703 & ~x704 & ~x708 & ~x721 & ~x727 & ~x733 & ~x738 & ~x754 & ~x755 & ~x756 & ~x758 & ~x760 & ~x766 & ~x767 & ~x770 & ~x771 & ~x774 & ~x776 & ~x778;
assign c8231 = ~x3 & ~x13 & ~x14 & ~x25 & ~x26 & ~x27 & ~x28 & ~x31 & ~x38 & ~x39 & ~x42 & ~x46 & ~x53 & ~x55 & ~x59 & ~x65 & ~x67 & ~x70 & ~x73 & ~x75 & ~x77 & ~x80 & ~x84 & ~x85 & ~x98 & ~x101 & ~x105 & ~x106 & ~x107 & ~x109 & ~x120 & ~x121 & ~x124 & ~x126 & ~x132 & ~x138 & ~x146 & ~x150 & ~x151 & ~x174 & ~x194 & ~x195 & ~x197 & ~x201 & ~x225 & ~x227 & ~x252 & ~x303 & ~x306 & ~x331 & ~x366 & ~x388 & ~x395 & ~x417 & ~x422 & ~x423 & ~x450 & ~x451 & ~x473 & ~x503 & ~x505 & ~x506 & ~x535 & ~x558 & ~x560 & ~x572 & ~x583 & ~x595 & ~x597 & ~x599 & ~x617 & ~x619 & ~x622 & ~x624 & ~x640 & ~x643 & ~x646 & ~x647 & ~x666 & ~x668 & ~x670 & ~x674 & ~x675 & ~x676 & ~x677 & ~x678 & ~x694 & ~x696 & ~x697 & ~x699 & ~x706 & ~x723 & ~x725 & ~x730 & ~x731 & ~x733 & ~x737 & ~x754 & ~x756 & ~x757 & ~x762 & ~x766 & ~x770 & ~x771 & ~x777;
assign c8233 =  x291 &  x346 &  x374 &  x402 & ~x11 & ~x23 & ~x24 & ~x39 & ~x40 & ~x45 & ~x46 & ~x49 & ~x54 & ~x61 & ~x75 & ~x86 & ~x99 & ~x103 & ~x112 & ~x113 & ~x115 & ~x116 & ~x120 & ~x121 & ~x129 & ~x143 & ~x171 & ~x252 & ~x254 & ~x284 & ~x302 & ~x307 & ~x312 & ~x313 & ~x361 & ~x392 & ~x448 & ~x453 & ~x473 & ~x504 & ~x541 & ~x559 & ~x563 & ~x582 & ~x586 & ~x612 & ~x614 & ~x621 & ~x638 & ~x640 & ~x672 & ~x674 & ~x692 & ~x693 & ~x702 & ~x705 & ~x729 & ~x779;
assign c8235 =  x296 &  x324 &  x489 & ~x100 & ~x143 & ~x274 & ~x275 & ~x317 & ~x318 & ~x319 & ~x320 & ~x419 & ~x421 & ~x507 & ~x589 & ~x735;
assign c8237 = ~x0 & ~x5 & ~x6 & ~x10 & ~x11 & ~x12 & ~x17 & ~x19 & ~x25 & ~x28 & ~x29 & ~x30 & ~x33 & ~x35 & ~x39 & ~x44 & ~x45 & ~x46 & ~x49 & ~x50 & ~x52 & ~x53 & ~x54 & ~x58 & ~x63 & ~x65 & ~x67 & ~x71 & ~x73 & ~x75 & ~x76 & ~x78 & ~x83 & ~x86 & ~x91 & ~x104 & ~x105 & ~x107 & ~x108 & ~x109 & ~x110 & ~x116 & ~x119 & ~x136 & ~x142 & ~x164 & ~x165 & ~x166 & ~x173 & ~x196 & ~x197 & ~x220 & ~x222 & ~x225 & ~x253 & ~x266 & ~x276 & ~x277 & ~x279 & ~x280 & ~x292 & ~x293 & ~x303 & ~x305 & ~x309 & ~x311 & ~x316 & ~x320 & ~x321 & ~x331 & ~x332 & ~x334 & ~x335 & ~x336 & ~x338 & ~x339 & ~x345 & ~x347 & ~x348 & ~x360 & ~x364 & ~x368 & ~x369 & ~x372 & ~x374 & ~x390 & ~x393 & ~x396 & ~x398 & ~x400 & ~x416 & ~x417 & ~x418 & ~x422 & ~x423 & ~x443 & ~x444 & ~x445 & ~x446 & ~x448 & ~x449 & ~x450 & ~x451 & ~x473 & ~x474 & ~x476 & ~x501 & ~x503 & ~x530 & ~x532 & ~x533 & ~x535 & ~x557 & ~x560 & ~x587 & ~x589 & ~x614 & ~x616 & ~x617 & ~x642 & ~x644 & ~x645 & ~x646 & ~x670 & ~x671 & ~x674 & ~x694 & ~x704 & ~x706 & ~x715 & ~x718 & ~x722 & ~x723 & ~x731 & ~x733 & ~x734 & ~x736 & ~x737 & ~x738 & ~x741 & ~x744 & ~x746 & ~x748 & ~x753 & ~x757 & ~x761 & ~x764 & ~x766 & ~x777 & ~x778 & ~x781 & ~x782;
assign c8239 =  x523 &  x550 & ~x2 & ~x7 & ~x8 & ~x196 & ~x201 & ~x279 & ~x392 & ~x407 & ~x417 & ~x613 & ~x641 & ~x741 & ~x750 & ~x752;
assign c8241 = ~x2 & ~x17 & ~x18 & ~x20 & ~x30 & ~x31 & ~x54 & ~x57 & ~x66 & ~x71 & ~x72 & ~x77 & ~x78 & ~x96 & ~x103 & ~x116 & ~x134 & ~x164 & ~x165 & ~x194 & ~x200 & ~x201 & ~x219 & ~x227 & ~x236 & ~x246 & ~x248 & ~x252 & ~x260 & ~x264 & ~x275 & ~x290 & ~x291 & ~x300 & ~x304 & ~x306 & ~x309 & ~x310 & ~x311 & ~x313 & ~x317 & ~x329 & ~x335 & ~x341 & ~x343 & ~x345 & ~x358 & ~x369 & ~x371 & ~x397 & ~x398 & ~x419 & ~x422 & ~x426 & ~x444 & ~x450 & ~x456 & ~x470 & ~x474 & ~x504 & ~x507 & ~x529 & ~x584 & ~x590 & ~x642 & ~x645 & ~x647 & ~x670 & ~x675 & ~x694 & ~x702 & ~x703 & ~x711 & ~x715 & ~x720 & ~x723 & ~x724 & ~x725 & ~x734 & ~x735 & ~x742 & ~x749 & ~x751 & ~x762 & ~x773 & ~x780;
assign c8243 =  x270 & ~x10 & ~x13 & ~x17 & ~x20 & ~x21 & ~x26 & ~x31 & ~x35 & ~x50 & ~x59 & ~x80 & ~x94 & ~x102 & ~x113 & ~x120 & ~x124 & ~x139 & ~x141 & ~x145 & ~x165 & ~x169 & ~x180 & ~x181 & ~x182 & ~x183 & ~x209 & ~x227 & ~x252 & ~x253 & ~x332 & ~x335 & ~x362 & ~x366 & ~x390 & ~x422 & ~x507 & ~x535 & ~x556 & ~x557 & ~x635 & ~x641 & ~x645 & ~x671 & ~x676 & ~x697 & ~x700 & ~x719 & ~x765 & ~x776;
assign c8245 = ~x0 & ~x4 & ~x6 & ~x8 & ~x13 & ~x26 & ~x28 & ~x31 & ~x35 & ~x43 & ~x44 & ~x46 & ~x48 & ~x49 & ~x50 & ~x57 & ~x60 & ~x62 & ~x75 & ~x76 & ~x77 & ~x79 & ~x83 & ~x87 & ~x92 & ~x93 & ~x108 & ~x110 & ~x116 & ~x118 & ~x119 & ~x124 & ~x137 & ~x143 & ~x144 & ~x146 & ~x153 & ~x169 & ~x170 & ~x182 & ~x193 & ~x195 & ~x197 & ~x220 & ~x222 & ~x248 & ~x277 & ~x280 & ~x282 & ~x303 & ~x305 & ~x306 & ~x307 & ~x309 & ~x332 & ~x336 & ~x389 & ~x390 & ~x392 & ~x447 & ~x451 & ~x474 & ~x475 & ~x476 & ~x477 & ~x502 & ~x533 & ~x534 & ~x557 & ~x563 & ~x588 & ~x593 & ~x602 & ~x612 & ~x617 & ~x630 & ~x631 & ~x641 & ~x643 & ~x645 & ~x648 & ~x649 & ~x658 & ~x659 & ~x669 & ~x687 & ~x714 & ~x724 & ~x728 & ~x729 & ~x730 & ~x749 & ~x754 & ~x755 & ~x767 & ~x782 & ~x783;
assign c8247 =  x372 &  x427 &  x455 & ~x6 & ~x12 & ~x25 & ~x26 & ~x35 & ~x37 & ~x39 & ~x41 & ~x48 & ~x50 & ~x52 & ~x66 & ~x67 & ~x80 & ~x90 & ~x109 & ~x111 & ~x115 & ~x116 & ~x119 & ~x127 & ~x138 & ~x140 & ~x141 & ~x227 & ~x392 & ~x477 & ~x504 & ~x507 & ~x530 & ~x536 & ~x564 & ~x592 & ~x673 & ~x676 & ~x701 & ~x702 & ~x730 & ~x732 & ~x735 & ~x740 & ~x755 & ~x768 & ~x778 & ~x781;
assign c8249 =  x580 & ~x191 & ~x195 & ~x197 & ~x291 & ~x343 & ~x615 & ~x779;
assign c8251 =  x322 &  x517 &  x545 & ~x7 & ~x26 & ~x160 & ~x187 & ~x199 & ~x303 & ~x317 & ~x345 & ~x371;
assign c8253 =  x542 & ~x1 & ~x3 & ~x16 & ~x20 & ~x53 & ~x170 & ~x223 & ~x224 & ~x250 & ~x251 & ~x258 & ~x313 & ~x314 & ~x338 & ~x342 & ~x358 & ~x361 & ~x362 & ~x447 & ~x452 & ~x560 & ~x587 & ~x616 & ~x627 & ~x655 & ~x658 & ~x660 & ~x671 & ~x682 & ~x684 & ~x686 & ~x687 & ~x691 & ~x692 & ~x702 & ~x725 & ~x738 & ~x748 & ~x751;
assign c8255 =  x148;
assign c8257 =  x268 & ~x64 & ~x109 & ~x135 & ~x191 & ~x219 & ~x245 & ~x246 & ~x247 & ~x273 & ~x292 & ~x342 & ~x347 & ~x355 & ~x373 & ~x383 & ~x397 & ~x401 & ~x503 & ~x677 & ~x695 & ~x700;
assign c8259 = ~x10 & ~x13 & ~x17 & ~x19 & ~x23 & ~x31 & ~x39 & ~x41 & ~x59 & ~x65 & ~x66 & ~x69 & ~x88 & ~x92 & ~x100 & ~x194 & ~x227 & ~x237 & ~x247 & ~x252 & ~x255 & ~x256 & ~x263 & ~x264 & ~x277 & ~x278 & ~x282 & ~x290 & ~x291 & ~x292 & ~x306 & ~x312 & ~x314 & ~x315 & ~x318 & ~x330 & ~x335 & ~x340 & ~x345 & ~x358 & ~x364 & ~x368 & ~x369 & ~x370 & ~x371 & ~x372 & ~x386 & ~x396 & ~x422 & ~x428 & ~x443 & ~x444 & ~x448 & ~x471 & ~x474 & ~x500 & ~x501 & ~x505 & ~x644 & ~x674 & ~x677 & ~x712 & ~x716 & ~x719 & ~x728 & ~x739 & ~x743 & ~x745 & ~x747 & ~x760 & ~x762 & ~x765 & ~x766 & ~x775;
assign c8261 =  x441 & ~x377;
assign c8263 =  x296 & ~x29 & ~x45 & ~x111 & ~x181 & ~x208 & ~x236 & ~x307 & ~x341 & ~x444 & ~x604 & ~x632 & ~x647 & ~x660 & ~x689 & ~x702 & ~x715;
assign c8265 = ~x0 & ~x8 & ~x10 & ~x15 & ~x16 & ~x20 & ~x34 & ~x44 & ~x51 & ~x61 & ~x69 & ~x71 & ~x73 & ~x74 & ~x77 & ~x87 & ~x90 & ~x94 & ~x95 & ~x100 & ~x117 & ~x137 & ~x140 & ~x199 & ~x223 & ~x248 & ~x251 & ~x277 & ~x281 & ~x305 & ~x334 & ~x362 & ~x367 & ~x415 & ~x416 & ~x418 & ~x420 & ~x444 & ~x447 & ~x455 & ~x473 & ~x474 & ~x475 & ~x483 & ~x484 & ~x501 & ~x513 & ~x514 & ~x515 & ~x517 & ~x543 & ~x544 & ~x546 & ~x558 & ~x585 & ~x590 & ~x611 & ~x613 & ~x616 & ~x638 & ~x642 & ~x645 & ~x646 & ~x647 & ~x649 & ~x669 & ~x670 & ~x671 & ~x673 & ~x676 & ~x701 & ~x702 & ~x725 & ~x730 & ~x733 & ~x734 & ~x735 & ~x740 & ~x753 & ~x756;
assign c8267 =  x656 & ~x10 & ~x17 & ~x19 & ~x21 & ~x26 & ~x30 & ~x39 & ~x48 & ~x54 & ~x55 & ~x64 & ~x68 & ~x74 & ~x75 & ~x77 & ~x84 & ~x93 & ~x94 & ~x95 & ~x108 & ~x140 & ~x170 & ~x196 & ~x198 & ~x252 & ~x386 & ~x388 & ~x390 & ~x392 & ~x397 & ~x421 & ~x485 & ~x500 & ~x501 & ~x514 & ~x515 & ~x544 & ~x563 & ~x564 & ~x566 & ~x587 & ~x643 & ~x674 & ~x697 & ~x699 & ~x720 & ~x721 & ~x724 & ~x746 & ~x751 & ~x766 & ~x773 & ~x776 & ~x782;
assign c8269 = ~x3 & ~x11 & ~x13 & ~x14 & ~x18 & ~x22 & ~x24 & ~x25 & ~x29 & ~x30 & ~x32 & ~x42 & ~x48 & ~x49 & ~x50 & ~x56 & ~x58 & ~x75 & ~x76 & ~x88 & ~x90 & ~x105 & ~x106 & ~x108 & ~x115 & ~x116 & ~x133 & ~x136 & ~x137 & ~x140 & ~x141 & ~x143 & ~x171 & ~x195 & ~x221 & ~x224 & ~x226 & ~x250 & ~x280 & ~x310 & ~x312 & ~x336 & ~x338 & ~x363 & ~x382 & ~x390 & ~x393 & ~x395 & ~x409 & ~x418 & ~x420 & ~x422 & ~x436 & ~x437 & ~x445 & ~x448 & ~x450 & ~x451 & ~x463 & ~x464 & ~x465 & ~x480 & ~x491 & ~x493 & ~x503 & ~x519 & ~x530 & ~x534 & ~x536 & ~x564 & ~x588 & ~x613 & ~x616 & ~x646 & ~x671 & ~x675 & ~x687 & ~x691 & ~x692 & ~x696 & ~x699 & ~x705 & ~x706 & ~x707 & ~x710 & ~x714 & ~x717 & ~x718 & ~x719 & ~x723 & ~x735 & ~x737 & ~x753 & ~x754 & ~x757 & ~x758 & ~x760 & ~x761 & ~x764 & ~x765 & ~x768 & ~x771 & ~x775 & ~x778 & ~x779 & ~x780 & ~x783;
assign c8271 =  x572 &  x573 & ~x0 & ~x1 & ~x7 & ~x9 & ~x11 & ~x19 & ~x29 & ~x30 & ~x36 & ~x42 & ~x45 & ~x52 & ~x57 & ~x68 & ~x76 & ~x77 & ~x78 & ~x81 & ~x82 & ~x88 & ~x92 & ~x94 & ~x107 & ~x112 & ~x117 & ~x167 & ~x188 & ~x189 & ~x199 & ~x216 & ~x226 & ~x248 & ~x288 & ~x299 & ~x300 & ~x306 & ~x311 & ~x313 & ~x330 & ~x336 & ~x338 & ~x343 & ~x358 & ~x390 & ~x415 & ~x416 & ~x505 & ~x507 & ~x508 & ~x510 & ~x529 & ~x535 & ~x558 & ~x559 & ~x587 & ~x592 & ~x594 & ~x614 & ~x615 & ~x645 & ~x646 & ~x662 & ~x686 & ~x703 & ~x716 & ~x722 & ~x723 & ~x725 & ~x732 & ~x737 & ~x747 & ~x768 & ~x769 & ~x783;
assign c8273 =  x739;
assign c8275 =  x297 &  x299 & ~x12 & ~x19 & ~x75 & ~x76 & ~x483 & ~x513 & ~x514 & ~x635 & ~x661 & ~x720;
assign c8277 = ~x0 & ~x2 & ~x3 & ~x6 & ~x7 & ~x8 & ~x9 & ~x10 & ~x15 & ~x16 & ~x20 & ~x21 & ~x23 & ~x25 & ~x26 & ~x27 & ~x31 & ~x37 & ~x43 & ~x45 & ~x46 & ~x51 & ~x54 & ~x56 & ~x57 & ~x59 & ~x60 & ~x61 & ~x63 & ~x64 & ~x67 & ~x75 & ~x78 & ~x83 & ~x84 & ~x88 & ~x97 & ~x100 & ~x103 & ~x107 & ~x110 & ~x111 & ~x113 & ~x131 & ~x132 & ~x137 & ~x138 & ~x139 & ~x144 & ~x166 & ~x167 & ~x168 & ~x169 & ~x171 & ~x172 & ~x193 & ~x197 & ~x222 & ~x224 & ~x247 & ~x248 & ~x250 & ~x253 & ~x275 & ~x276 & ~x303 & ~x305 & ~x309 & ~x310 & ~x321 & ~x336 & ~x337 & ~x339 & ~x347 & ~x348 & ~x362 & ~x364 & ~x365 & ~x366 & ~x373 & ~x374 & ~x375 & ~x392 & ~x395 & ~x398 & ~x400 & ~x401 & ~x402 & ~x403 & ~x419 & ~x420 & ~x445 & ~x446 & ~x451 & ~x473 & ~x476 & ~x479 & ~x502 & ~x504 & ~x505 & ~x530 & ~x560 & ~x561 & ~x586 & ~x589 & ~x618 & ~x641 & ~x645 & ~x646 & ~x671 & ~x696 & ~x697 & ~x700 & ~x718 & ~x719 & ~x721 & ~x722 & ~x728 & ~x731 & ~x739 & ~x745 & ~x749 & ~x757 & ~x759 & ~x760 & ~x762 & ~x763 & ~x768 & ~x774 & ~x778 & ~x779 & ~x781 & ~x782 & ~x783;
assign c8279 =  x679 &  x706;
assign c8281 =  x654 & ~x2 & ~x3 & ~x4 & ~x5 & ~x14 & ~x16 & ~x20 & ~x23 & ~x35 & ~x41 & ~x48 & ~x61 & ~x64 & ~x65 & ~x71 & ~x75 & ~x77 & ~x81 & ~x83 & ~x85 & ~x89 & ~x101 & ~x104 & ~x106 & ~x108 & ~x109 & ~x118 & ~x144 & ~x220 & ~x222 & ~x226 & ~x254 & ~x255 & ~x280 & ~x281 & ~x308 & ~x334 & ~x336 & ~x361 & ~x389 & ~x391 & ~x393 & ~x422 & ~x423 & ~x424 & ~x447 & ~x455 & ~x474 & ~x476 & ~x485 & ~x505 & ~x515 & ~x516 & ~x560 & ~x589 & ~x643 & ~x668 & ~x702 & ~x703 & ~x712 & ~x714 & ~x728 & ~x731 & ~x734 & ~x740 & ~x745 & ~x750 & ~x751 & ~x753 & ~x755 & ~x757 & ~x762 & ~x769 & ~x780;
assign c8283 =  x455 & ~x0 & ~x3 & ~x18 & ~x30 & ~x41 & ~x47 & ~x48 & ~x61 & ~x66 & ~x67 & ~x114 & ~x118 & ~x165 & ~x166 & ~x167 & ~x197 & ~x253 & ~x281 & ~x304 & ~x305 & ~x333 & ~x335 & ~x363 & ~x394 & ~x417 & ~x477 & ~x530 & ~x532 & ~x562 & ~x590 & ~x616 & ~x617 & ~x643 & ~x654 & ~x655 & ~x668 & ~x681 & ~x683 & ~x697 & ~x698 & ~x700 & ~x702 & ~x706 & ~x712 & ~x726 & ~x737 & ~x740 & ~x741 & ~x742 & ~x747 & ~x751 & ~x761 & ~x768 & ~x772 & ~x777;
assign c8285 =  x483 & ~x379 & ~x669 & ~x779;
assign c8287 =  x439 &  x493 &  x521 & ~x0 & ~x7 & ~x9 & ~x11 & ~x12 & ~x17 & ~x18 & ~x20 & ~x21 & ~x23 & ~x28 & ~x30 & ~x36 & ~x37 & ~x39 & ~x45 & ~x51 & ~x54 & ~x56 & ~x63 & ~x65 & ~x69 & ~x73 & ~x77 & ~x81 & ~x82 & ~x83 & ~x86 & ~x92 & ~x108 & ~x111 & ~x113 & ~x114 & ~x118 & ~x121 & ~x139 & ~x140 & ~x145 & ~x147 & ~x165 & ~x167 & ~x191 & ~x192 & ~x194 & ~x197 & ~x199 & ~x200 & ~x224 & ~x226 & ~x227 & ~x255 & ~x277 & ~x279 & ~x281 & ~x284 & ~x304 & ~x305 & ~x309 & ~x335 & ~x336 & ~x360 & ~x361 & ~x362 & ~x364 & ~x366 & ~x389 & ~x392 & ~x421 & ~x422 & ~x446 & ~x448 & ~x449 & ~x451 & ~x479 & ~x528 & ~x529 & ~x533 & ~x534 & ~x535 & ~x560 & ~x588 & ~x589 & ~x592 & ~x608 & ~x618 & ~x620 & ~x637 & ~x639 & ~x640 & ~x642 & ~x645 & ~x662 & ~x664 & ~x668 & ~x672 & ~x678 & ~x691 & ~x692 & ~x694 & ~x695 & ~x701 & ~x705 & ~x719 & ~x722 & ~x727 & ~x732 & ~x734 & ~x737 & ~x744 & ~x751 & ~x754 & ~x760 & ~x763 & ~x764 & ~x768 & ~x771 & ~x774 & ~x777 & ~x778 & ~x780 & ~x781 & ~x783;
assign c8289 =  x441 &  x496 &  x523 & ~x2 & ~x18 & ~x27 & ~x32 & ~x33 & ~x52 & ~x58 & ~x82 & ~x89 & ~x107 & ~x114 & ~x162 & ~x249 & ~x279 & ~x365 & ~x448 & ~x473 & ~x475 & ~x504 & ~x506 & ~x532 & ~x559 & ~x617 & ~x620 & ~x639 & ~x647 & ~x670 & ~x671 & ~x723 & ~x726 & ~x741 & ~x744 & ~x754 & ~x755 & ~x758;
assign c8291 = ~x4 & ~x18 & ~x23 & ~x24 & ~x26 & ~x27 & ~x30 & ~x61 & ~x70 & ~x71 & ~x74 & ~x92 & ~x96 & ~x98 & ~x100 & ~x118 & ~x121 & ~x141 & ~x142 & ~x164 & ~x194 & ~x223 & ~x248 & ~x277 & ~x281 & ~x282 & ~x306 & ~x307 & ~x331 & ~x363 & ~x370 & ~x387 & ~x393 & ~x398 & ~x446 & ~x475 & ~x477 & ~x502 & ~x510 & ~x511 & ~x537 & ~x539 & ~x540 & ~x541 & ~x543 & ~x560 & ~x562 & ~x571 & ~x572 & ~x573 & ~x595 & ~x612 & ~x613 & ~x615 & ~x644 & ~x665 & ~x668 & ~x673 & ~x675 & ~x704 & ~x706 & ~x724 & ~x727 & ~x729 & ~x733 & ~x750 & ~x751 & ~x752 & ~x783;
assign c8293 =  x320 &  x375 &  x492 & ~x0 & ~x4 & ~x17 & ~x27 & ~x36 & ~x38 & ~x39 & ~x44 & ~x52 & ~x59 & ~x70 & ~x83 & ~x91 & ~x98 & ~x108 & ~x111 & ~x141 & ~x178 & ~x197 & ~x200 & ~x206 & ~x225 & ~x228 & ~x252 & ~x256 & ~x257 & ~x258 & ~x259 & ~x260 & ~x284 & ~x285 & ~x308 & ~x309 & ~x311 & ~x313 & ~x339 & ~x340 & ~x363 & ~x364 & ~x365 & ~x367 & ~x389 & ~x391 & ~x393 & ~x447 & ~x478 & ~x501 & ~x504 & ~x506 & ~x589 & ~x590 & ~x612 & ~x639 & ~x640 & ~x666 & ~x673 & ~x675 & ~x676 & ~x686 & ~x694 & ~x697 & ~x701 & ~x702 & ~x705 & ~x714 & ~x717 & ~x727 & ~x728 & ~x749 & ~x751 & ~x759 & ~x763 & ~x765 & ~x766 & ~x767 & ~x769 & ~x773 & ~x778 & ~x782;
assign c8295 = ~x11 & ~x14 & ~x17 & ~x33 & ~x41 & ~x54 & ~x56 & ~x72 & ~x75 & ~x85 & ~x87 & ~x88 & ~x92 & ~x113 & ~x137 & ~x140 & ~x170 & ~x195 & ~x200 & ~x216 & ~x220 & ~x244 & ~x248 & ~x262 & ~x263 & ~x271 & ~x272 & ~x277 & ~x278 & ~x284 & ~x301 & ~x304 & ~x317 & ~x327 & ~x334 & ~x336 & ~x337 & ~x341 & ~x345 & ~x362 & ~x369 & ~x370 & ~x388 & ~x389 & ~x417 & ~x446 & ~x448 & ~x450 & ~x453 & ~x478 & ~x505 & ~x537 & ~x559 & ~x561 & ~x563 & ~x592 & ~x593 & ~x618 & ~x623 & ~x638 & ~x639 & ~x641 & ~x643 & ~x645 & ~x652 & ~x670 & ~x679 & ~x696 & ~x698 & ~x699 & ~x700 & ~x704 & ~x705 & ~x709 & ~x713 & ~x722 & ~x726 & ~x730 & ~x732 & ~x735 & ~x748 & ~x749 & ~x767 & ~x769 & ~x777;
assign c8297 =  x162 & ~x325;
assign c8299 =  x178 &  x182 & ~x0 & ~x2 & ~x9 & ~x10 & ~x12 & ~x13 & ~x17 & ~x19 & ~x20 & ~x25 & ~x27 & ~x30 & ~x35 & ~x43 & ~x45 & ~x54 & ~x56 & ~x63 & ~x70 & ~x73 & ~x76 & ~x80 & ~x81 & ~x87 & ~x92 & ~x98 & ~x101 & ~x109 & ~x113 & ~x115 & ~x133 & ~x136 & ~x138 & ~x139 & ~x144 & ~x163 & ~x164 & ~x191 & ~x192 & ~x193 & ~x219 & ~x226 & ~x227 & ~x251 & ~x253 & ~x276 & ~x282 & ~x292 & ~x308 & ~x313 & ~x315 & ~x316 & ~x317 & ~x318 & ~x330 & ~x338 & ~x340 & ~x342 & ~x343 & ~x344 & ~x358 & ~x362 & ~x368 & ~x369 & ~x371 & ~x386 & ~x389 & ~x390 & ~x397 & ~x417 & ~x421 & ~x422 & ~x424 & ~x446 & ~x448 & ~x449 & ~x450 & ~x451 & ~x476 & ~x477 & ~x505 & ~x506 & ~x507 & ~x530 & ~x558 & ~x589 & ~x613 & ~x614 & ~x618 & ~x645 & ~x692 & ~x695 & ~x697 & ~x699 & ~x701 & ~x706 & ~x720 & ~x726 & ~x727 & ~x728 & ~x733 & ~x738 & ~x742 & ~x744 & ~x747 & ~x750 & ~x755 & ~x759 & ~x760 & ~x764 & ~x765 & ~x772 & ~x782;
assign c90 =  x206 &  x693;
assign c92 =  x350 &  x408 & ~x19 & ~x21 & ~x52 & ~x158 & ~x160 & ~x166 & ~x179 & ~x206 & ~x221 & ~x280 & ~x387 & ~x468 & ~x522 & ~x550 & ~x555 & ~x579 & ~x611 & ~x632;
assign c94 =  x170;
assign c96 =  x206 & ~x2 & ~x5 & ~x6 & ~x13 & ~x15 & ~x19 & ~x21 & ~x23 & ~x29 & ~x32 & ~x33 & ~x35 & ~x38 & ~x41 & ~x43 & ~x45 & ~x46 & ~x51 & ~x55 & ~x56 & ~x60 & ~x61 & ~x69 & ~x70 & ~x72 & ~x75 & ~x78 & ~x81 & ~x83 & ~x84 & ~x85 & ~x89 & ~x92 & ~x95 & ~x102 & ~x113 & ~x115 & ~x117 & ~x118 & ~x121 & ~x129 & ~x130 & ~x131 & ~x136 & ~x144 & ~x147 & ~x148 & ~x158 & ~x159 & ~x161 & ~x162 & ~x168 & ~x170 & ~x172 & ~x173 & ~x174 & ~x188 & ~x189 & ~x192 & ~x194 & ~x196 & ~x197 & ~x199 & ~x215 & ~x218 & ~x219 & ~x221 & ~x224 & ~x246 & ~x248 & ~x255 & ~x256 & ~x264 & ~x274 & ~x275 & ~x282 & ~x283 & ~x284 & ~x291 & ~x293 & ~x303 & ~x304 & ~x310 & ~x331 & ~x333 & ~x334 & ~x335 & ~x336 & ~x338 & ~x361 & ~x386 & ~x390 & ~x391 & ~x417 & ~x443 & ~x450 & ~x451 & ~x462 & ~x471 & ~x476 & ~x477 & ~x488 & ~x498 & ~x499 & ~x502 & ~x505 & ~x509 & ~x526 & ~x527 & ~x529 & ~x556 & ~x558 & ~x561 & ~x565 & ~x566 & ~x584 & ~x585 & ~x587 & ~x589 & ~x590 & ~x594 & ~x624 & ~x644 & ~x648 & ~x652 & ~x669 & ~x672 & ~x674 & ~x675 & ~x679 & ~x680 & ~x681 & ~x697 & ~x706 & ~x708 & ~x723 & ~x725 & ~x732 & ~x735 & ~x742 & ~x744 & ~x745 & ~x746 & ~x752 & ~x754 & ~x756 & ~x759 & ~x760 & ~x761 & ~x763 & ~x765 & ~x767 & ~x768 & ~x772 & ~x778 & ~x781 & ~x783;
assign c98 =  x208 & ~x0 & ~x5 & ~x8 & ~x15 & ~x16 & ~x19 & ~x24 & ~x28 & ~x36 & ~x40 & ~x41 & ~x43 & ~x48 & ~x50 & ~x54 & ~x56 & ~x63 & ~x65 & ~x71 & ~x76 & ~x78 & ~x79 & ~x83 & ~x85 & ~x87 & ~x89 & ~x91 & ~x92 & ~x95 & ~x96 & ~x104 & ~x106 & ~x108 & ~x112 & ~x113 & ~x118 & ~x119 & ~x120 & ~x121 & ~x122 & ~x131 & ~x132 & ~x138 & ~x139 & ~x140 & ~x143 & ~x146 & ~x159 & ~x160 & ~x163 & ~x167 & ~x169 & ~x173 & ~x187 & ~x188 & ~x189 & ~x195 & ~x196 & ~x199 & ~x200 & ~x217 & ~x219 & ~x222 & ~x223 & ~x224 & ~x227 & ~x252 & ~x255 & ~x273 & ~x278 & ~x279 & ~x281 & ~x309 & ~x311 & ~x320 & ~x331 & ~x335 & ~x336 & ~x337 & ~x338 & ~x357 & ~x361 & ~x363 & ~x365 & ~x366 & ~x387 & ~x395 & ~x396 & ~x413 & ~x414 & ~x417 & ~x420 & ~x421 & ~x445 & ~x446 & ~x448 & ~x451 & ~x476 & ~x478 & ~x479 & ~x501 & ~x502 & ~x503 & ~x528 & ~x529 & ~x533 & ~x534 & ~x554 & ~x555 & ~x557 & ~x560 & ~x563 & ~x565 & ~x573 & ~x581 & ~x586 & ~x588 & ~x589 & ~x592 & ~x593 & ~x594 & ~x598 & ~x599 & ~x600 & ~x611 & ~x619 & ~x623 & ~x639 & ~x641 & ~x642 & ~x644 & ~x645 & ~x647 & ~x649 & ~x666 & ~x670 & ~x673 & ~x674 & ~x676 & ~x679 & ~x682 & ~x695 & ~x702 & ~x709 & ~x710 & ~x712 & ~x713 & ~x714 & ~x725 & ~x726 & ~x729 & ~x730 & ~x731 & ~x732 & ~x737 & ~x738 & ~x740 & ~x744 & ~x756 & ~x758 & ~x759 & ~x760 & ~x761 & ~x763 & ~x766 & ~x767 & ~x769 & ~x771 & ~x773 & ~x779 & ~x783;
assign c910 =  x216 &  x406;
assign c912 =  x751;
assign c914 =  x666 &  x695;
assign c916 = ~x1 & ~x6 & ~x10 & ~x15 & ~x16 & ~x19 & ~x20 & ~x21 & ~x22 & ~x23 & ~x25 & ~x26 & ~x27 & ~x28 & ~x29 & ~x32 & ~x34 & ~x35 & ~x41 & ~x43 & ~x45 & ~x46 & ~x48 & ~x49 & ~x51 & ~x53 & ~x54 & ~x56 & ~x58 & ~x60 & ~x64 & ~x66 & ~x70 & ~x71 & ~x75 & ~x86 & ~x87 & ~x89 & ~x90 & ~x91 & ~x92 & ~x95 & ~x97 & ~x99 & ~x101 & ~x102 & ~x103 & ~x105 & ~x113 & ~x114 & ~x115 & ~x118 & ~x122 & ~x123 & ~x124 & ~x128 & ~x132 & ~x133 & ~x134 & ~x136 & ~x137 & ~x138 & ~x139 & ~x140 & ~x141 & ~x147 & ~x148 & ~x151 & ~x152 & ~x153 & ~x154 & ~x155 & ~x156 & ~x158 & ~x162 & ~x163 & ~x164 & ~x168 & ~x173 & ~x176 & ~x178 & ~x179 & ~x191 & ~x193 & ~x194 & ~x195 & ~x197 & ~x202 & ~x204 & ~x205 & ~x206 & ~x221 & ~x225 & ~x226 & ~x229 & ~x230 & ~x232 & ~x233 & ~x249 & ~x250 & ~x252 & ~x255 & ~x259 & ~x275 & ~x281 & ~x283 & ~x284 & ~x285 & ~x304 & ~x308 & ~x310 & ~x311 & ~x312 & ~x313 & ~x332 & ~x341 & ~x342 & ~x343 & ~x361 & ~x362 & ~x365 & ~x369 & ~x390 & ~x393 & ~x398 & ~x412 & ~x415 & ~x420 & ~x421 & ~x422 & ~x424 & ~x426 & ~x427 & ~x440 & ~x443 & ~x444 & ~x445 & ~x450 & ~x451 & ~x453 & ~x454 & ~x467 & ~x469 & ~x472 & ~x473 & ~x477 & ~x479 & ~x481 & ~x495 & ~x498 & ~x501 & ~x504 & ~x509 & ~x510 & ~x511 & ~x523 & ~x524 & ~x525 & ~x527 & ~x529 & ~x530 & ~x532 & ~x534 & ~x535 & ~x552 & ~x555 & ~x557 & ~x558 & ~x559 & ~x561 & ~x562 & ~x563 & ~x564 & ~x566 & ~x568 & ~x570 & ~x581 & ~x584 & ~x585 & ~x590 & ~x591 & ~x592 & ~x596 & ~x597 & ~x598 & ~x607 & ~x608 & ~x610 & ~x612 & ~x616 & ~x624 & ~x626 & ~x634 & ~x635 & ~x643 & ~x645 & ~x646 & ~x649 & ~x650 & ~x651 & ~x653 & ~x662 & ~x663 & ~x665 & ~x666 & ~x667 & ~x673 & ~x677 & ~x678 & ~x680 & ~x683 & ~x691 & ~x693 & ~x694 & ~x695 & ~x696 & ~x701 & ~x704 & ~x706 & ~x707 & ~x719 & ~x720 & ~x722 & ~x728 & ~x735 & ~x738 & ~x746 & ~x748 & ~x749 & ~x750 & ~x751 & ~x756 & ~x759 & ~x761 & ~x763 & ~x764 & ~x765 & ~x767 & ~x768 & ~x769 & ~x770 & ~x772 & ~x775 & ~x778 & ~x780 & ~x781 & ~x783;
assign c918 =  x380 & ~x0 & ~x8 & ~x10 & ~x11 & ~x13 & ~x15 & ~x16 & ~x17 & ~x19 & ~x21 & ~x22 & ~x24 & ~x25 & ~x26 & ~x30 & ~x32 & ~x36 & ~x41 & ~x43 & ~x45 & ~x47 & ~x49 & ~x53 & ~x57 & ~x59 & ~x60 & ~x61 & ~x64 & ~x65 & ~x67 & ~x69 & ~x70 & ~x71 & ~x72 & ~x76 & ~x85 & ~x89 & ~x90 & ~x91 & ~x94 & ~x98 & ~x100 & ~x104 & ~x107 & ~x108 & ~x109 & ~x115 & ~x120 & ~x124 & ~x128 & ~x131 & ~x133 & ~x136 & ~x144 & ~x145 & ~x150 & ~x159 & ~x160 & ~x163 & ~x165 & ~x167 & ~x172 & ~x186 & ~x195 & ~x200 & ~x217 & ~x221 & ~x225 & ~x226 & ~x229 & ~x230 & ~x231 & ~x243 & ~x247 & ~x249 & ~x256 & ~x258 & ~x272 & ~x274 & ~x280 & ~x284 & ~x285 & ~x303 & ~x307 & ~x308 & ~x309 & ~x310 & ~x314 & ~x328 & ~x330 & ~x334 & ~x336 & ~x337 & ~x355 & ~x358 & ~x359 & ~x362 & ~x370 & ~x387 & ~x388 & ~x389 & ~x411 & ~x415 & ~x416 & ~x421 & ~x423 & ~x424 & ~x426 & ~x427 & ~x441 & ~x443 & ~x450 & ~x452 & ~x453 & ~x454 & ~x455 & ~x469 & ~x478 & ~x496 & ~x501 & ~x503 & ~x512 & ~x518 & ~x532 & ~x535 & ~x536 & ~x537 & ~x545 & ~x552 & ~x555 & ~x557 & ~x558 & ~x563 & ~x564 & ~x565 & ~x571 & ~x585 & ~x592 & ~x612 & ~x615 & ~x639 & ~x640 & ~x645 & ~x650 & ~x651 & ~x667 & ~x668 & ~x675 & ~x678 & ~x680 & ~x693 & ~x698 & ~x702 & ~x704 & ~x706 & ~x711 & ~x713 & ~x721 & ~x723 & ~x727 & ~x730 & ~x731 & ~x732 & ~x733 & ~x755 & ~x756 & ~x758 & ~x761 & ~x763 & ~x764 & ~x769 & ~x770 & ~x775;
assign c920 =  x640;
assign c922 =  x280;
assign c924 =  x379 & ~x0 & ~x12 & ~x22 & ~x27 & ~x38 & ~x39 & ~x40 & ~x41 & ~x46 & ~x52 & ~x53 & ~x81 & ~x82 & ~x96 & ~x98 & ~x106 & ~x111 & ~x113 & ~x115 & ~x118 & ~x122 & ~x123 & ~x129 & ~x131 & ~x132 & ~x136 & ~x142 & ~x144 & ~x159 & ~x163 & ~x166 & ~x170 & ~x188 & ~x190 & ~x191 & ~x199 & ~x203 & ~x254 & ~x276 & ~x279 & ~x281 & ~x284 & ~x287 & ~x295 & ~x308 & ~x358 & ~x360 & ~x392 & ~x396 & ~x397 & ~x412 & ~x418 & ~x445 & ~x446 & ~x449 & ~x454 & ~x478 & ~x481 & ~x488 & ~x510 & ~x511 & ~x528 & ~x541 & ~x542 & ~x553 & ~x565 & ~x581 & ~x634 & ~x639 & ~x641 & ~x647 & ~x648 & ~x664 & ~x671 & ~x673 & ~x674 & ~x676 & ~x697 & ~x706 & ~x729 & ~x732 & ~x737 & ~x746 & ~x752 & ~x758 & ~x765 & ~x769;
assign c926 =  x214 &  x405 & ~x36 & ~x39 & ~x52 & ~x72 & ~x76 & ~x90 & ~x95 & ~x107 & ~x109 & ~x131 & ~x142 & ~x151 & ~x165 & ~x179 & ~x180 & ~x228 & ~x259 & ~x306 & ~x314 & ~x362 & ~x390 & ~x443 & ~x472 & ~x481 & ~x495 & ~x510 & ~x536 & ~x549 & ~x550 & ~x584 & ~x592 & ~x595 & ~x604 & ~x606 & ~x611 & ~x614 & ~x620 & ~x630 & ~x636 & ~x673 & ~x676 & ~x685 & ~x748 & ~x758 & ~x759 & ~x778;
assign c928 =  x319 & ~x2 & ~x6 & ~x7 & ~x10 & ~x21 & ~x25 & ~x27 & ~x32 & ~x35 & ~x41 & ~x47 & ~x61 & ~x63 & ~x77 & ~x79 & ~x81 & ~x91 & ~x100 & ~x107 & ~x109 & ~x110 & ~x111 & ~x132 & ~x135 & ~x136 & ~x138 & ~x147 & ~x162 & ~x164 & ~x179 & ~x180 & ~x203 & ~x205 & ~x219 & ~x229 & ~x234 & ~x255 & ~x257 & ~x262 & ~x310 & ~x312 & ~x332 & ~x337 & ~x362 & ~x363 & ~x364 & ~x370 & ~x387 & ~x414 & ~x419 & ~x444 & ~x450 & ~x467 & ~x499 & ~x501 & ~x503 & ~x504 & ~x508 & ~x533 & ~x534 & ~x538 & ~x553 & ~x554 & ~x556 & ~x558 & ~x563 & ~x564 & ~x576 & ~x577 & ~x578 & ~x591 & ~x594 & ~x595 & ~x609 & ~x610 & ~x615 & ~x618 & ~x621 & ~x643 & ~x647 & ~x668 & ~x670 & ~x675 & ~x677 & ~x688 & ~x701 & ~x722 & ~x732 & ~x736 & ~x743 & ~x744 & ~x748 & ~x751 & ~x753 & ~x759 & ~x765 & ~x766 & ~x775 & ~x777 & ~x779 & ~x781 & ~x783;
assign c930 =  x207 &  x692;
assign c932 =  x723;
assign c934 =  x460 & ~x5 & ~x19 & ~x58 & ~x73 & ~x78 & ~x88 & ~x95 & ~x126 & ~x136 & ~x149 & ~x152 & ~x169 & ~x192 & ~x196 & ~x197 & ~x204 & ~x255 & ~x284 & ~x360 & ~x366 & ~x377 & ~x404 & ~x418 & ~x421 & ~x443 & ~x446 & ~x451 & ~x469 & ~x480 & ~x525 & ~x532 & ~x537 & ~x541 & ~x542 & ~x543 & ~x555 & ~x563 & ~x570 & ~x578 & ~x583 & ~x587 & ~x620 & ~x622 & ~x640 & ~x644 & ~x651 & ~x692 & ~x703 & ~x725 & ~x726 & ~x779 & ~x781;
assign c936 =  x211 & ~x0 & ~x13 & ~x17 & ~x24 & ~x25 & ~x38 & ~x40 & ~x46 & ~x50 & ~x60 & ~x61 & ~x71 & ~x75 & ~x78 & ~x79 & ~x81 & ~x87 & ~x89 & ~x90 & ~x93 & ~x96 & ~x102 & ~x111 & ~x113 & ~x114 & ~x128 & ~x130 & ~x132 & ~x134 & ~x144 & ~x152 & ~x154 & ~x156 & ~x161 & ~x162 & ~x163 & ~x164 & ~x165 & ~x168 & ~x202 & ~x204 & ~x206 & ~x231 & ~x244 & ~x245 & ~x246 & ~x247 & ~x249 & ~x250 & ~x255 & ~x274 & ~x275 & ~x285 & ~x331 & ~x332 & ~x335 & ~x337 & ~x340 & ~x341 & ~x359 & ~x364 & ~x365 & ~x369 & ~x385 & ~x387 & ~x390 & ~x391 & ~x393 & ~x412 & ~x415 & ~x443 & ~x446 & ~x454 & ~x472 & ~x474 & ~x475 & ~x481 & ~x482 & ~x500 & ~x501 & ~x502 & ~x503 & ~x508 & ~x525 & ~x557 & ~x558 & ~x568 & ~x569 & ~x582 & ~x589 & ~x591 & ~x600 & ~x615 & ~x617 & ~x618 & ~x621 & ~x623 & ~x636 & ~x637 & ~x638 & ~x642 & ~x643 & ~x645 & ~x646 & ~x648 & ~x649 & ~x654 & ~x655 & ~x666 & ~x670 & ~x682 & ~x683 & ~x695 & ~x712 & ~x722 & ~x725 & ~x731 & ~x732 & ~x734 & ~x735 & ~x744 & ~x749 & ~x756 & ~x762 & ~x763 & ~x765 & ~x777 & ~x780;
assign c938 =  x722;
assign c940 =  x240 &  x410 &  x457 & ~x9 & ~x14 & ~x71 & ~x78 & ~x90 & ~x124 & ~x155 & ~x180 & ~x222 & ~x232 & ~x279 & ~x309 & ~x366 & ~x392 & ~x419 & ~x422 & ~x469 & ~x504 & ~x538 & ~x539 & ~x562 & ~x597 & ~x612 & ~x622 & ~x676 & ~x677 & ~x692 & ~x774;
assign c942 =  x209 &  x211 &  x344 &  x355 & ~x7 & ~x32 & ~x34 & ~x38 & ~x50 & ~x80 & ~x93 & ~x110 & ~x115 & ~x125 & ~x131 & ~x161 & ~x170 & ~x230 & ~x331 & ~x337 & ~x339 & ~x392 & ~x393 & ~x448 & ~x478 & ~x501 & ~x554 & ~x561 & ~x582 & ~x587 & ~x599 & ~x611 & ~x613 & ~x649 & ~x650 & ~x671 & ~x698 & ~x730 & ~x746 & ~x759 & ~x768 & ~x770;
assign c944 =  x721;
assign c946 =  x342 & ~x36 & ~x185 & ~x229 & ~x248 & ~x275 & ~x347 & ~x443 & ~x528 & ~x571 & ~x600 & ~x631;
assign c948 =  x208 &  x404 & ~x6 & ~x7 & ~x11 & ~x12 & ~x15 & ~x17 & ~x18 & ~x23 & ~x25 & ~x31 & ~x32 & ~x33 & ~x36 & ~x37 & ~x38 & ~x39 & ~x40 & ~x41 & ~x43 & ~x50 & ~x53 & ~x57 & ~x59 & ~x60 & ~x63 & ~x64 & ~x65 & ~x70 & ~x74 & ~x77 & ~x81 & ~x83 & ~x86 & ~x93 & ~x95 & ~x98 & ~x99 & ~x100 & ~x105 & ~x109 & ~x110 & ~x111 & ~x114 & ~x115 & ~x118 & ~x119 & ~x121 & ~x132 & ~x134 & ~x136 & ~x137 & ~x143 & ~x146 & ~x163 & ~x167 & ~x169 & ~x171 & ~x172 & ~x174 & ~x192 & ~x193 & ~x196 & ~x197 & ~x201 & ~x220 & ~x222 & ~x223 & ~x224 & ~x248 & ~x276 & ~x280 & ~x281 & ~x282 & ~x283 & ~x284 & ~x305 & ~x306 & ~x311 & ~x332 & ~x334 & ~x337 & ~x340 & ~x387 & ~x389 & ~x390 & ~x396 & ~x397 & ~x423 & ~x442 & ~x443 & ~x444 & ~x445 & ~x446 & ~x448 & ~x453 & ~x455 & ~x456 & ~x457 & ~x458 & ~x459 & ~x460 & ~x461 & ~x471 & ~x474 & ~x479 & ~x480 & ~x483 & ~x487 & ~x488 & ~x489 & ~x497 & ~x500 & ~x505 & ~x506 & ~x508 & ~x526 & ~x532 & ~x536 & ~x558 & ~x562 & ~x582 & ~x584 & ~x585 & ~x588 & ~x589 & ~x592 & ~x611 & ~x617 & ~x618 & ~x621 & ~x638 & ~x641 & ~x642 & ~x645 & ~x647 & ~x669 & ~x675 & ~x677 & ~x704 & ~x705 & ~x720 & ~x726 & ~x728 & ~x729 & ~x732 & ~x744 & ~x747 & ~x749 & ~x753 & ~x755 & ~x761 & ~x767 & ~x769 & ~x782 & ~x783;
assign c950 =  x211 &  x382 &  x433 &  x465 & ~x1 & ~x7 & ~x10 & ~x12 & ~x16 & ~x17 & ~x24 & ~x25 & ~x27 & ~x29 & ~x30 & ~x34 & ~x39 & ~x45 & ~x47 & ~x55 & ~x56 & ~x71 & ~x77 & ~x90 & ~x91 & ~x96 & ~x101 & ~x104 & ~x107 & ~x115 & ~x117 & ~x119 & ~x134 & ~x138 & ~x139 & ~x143 & ~x145 & ~x148 & ~x149 & ~x161 & ~x167 & ~x170 & ~x173 & ~x174 & ~x196 & ~x201 & ~x202 & ~x226 & ~x227 & ~x254 & ~x255 & ~x256 & ~x277 & ~x280 & ~x281 & ~x307 & ~x311 & ~x334 & ~x340 & ~x360 & ~x366 & ~x393 & ~x394 & ~x444 & ~x451 & ~x535 & ~x543 & ~x567 & ~x587 & ~x588 & ~x591 & ~x618 & ~x619 & ~x645 & ~x649 & ~x650 & ~x666 & ~x690 & ~x699 & ~x700 & ~x701 & ~x705 & ~x724 & ~x728 & ~x730 & ~x732 & ~x743 & ~x750 & ~x759 & ~x762 & ~x765 & ~x769 & ~x771 & ~x781;
assign c952 =  x350 &  x351 &  x352 & ~x5 & ~x15 & ~x23 & ~x24 & ~x33 & ~x36 & ~x41 & ~x61 & ~x64 & ~x66 & ~x70 & ~x77 & ~x94 & ~x95 & ~x96 & ~x99 & ~x100 & ~x101 & ~x105 & ~x115 & ~x121 & ~x123 & ~x128 & ~x130 & ~x138 & ~x150 & ~x151 & ~x152 & ~x161 & ~x162 & ~x166 & ~x172 & ~x178 & ~x196 & ~x204 & ~x257 & ~x258 & ~x278 & ~x281 & ~x284 & ~x305 & ~x309 & ~x311 & ~x332 & ~x390 & ~x395 & ~x400 & ~x416 & ~x418 & ~x420 & ~x421 & ~x423 & ~x450 & ~x452 & ~x456 & ~x457 & ~x459 & ~x476 & ~x479 & ~x483 & ~x484 & ~x487 & ~x495 & ~x503 & ~x504 & ~x507 & ~x508 & ~x511 & ~x512 & ~x513 & ~x523 & ~x532 & ~x538 & ~x555 & ~x566 & ~x579 & ~x581 & ~x585 & ~x590 & ~x594 & ~x595 & ~x623 & ~x636 & ~x669 & ~x674 & ~x703 & ~x724 & ~x733 & ~x743 & ~x747 & ~x749 & ~x754 & ~x755 & ~x761 & ~x777 & ~x780;
assign c954 = ~x0 & ~x2 & ~x4 & ~x9 & ~x14 & ~x18 & ~x26 & ~x29 & ~x31 & ~x36 & ~x37 & ~x39 & ~x45 & ~x46 & ~x73 & ~x76 & ~x80 & ~x81 & ~x83 & ~x85 & ~x88 & ~x95 & ~x98 & ~x102 & ~x103 & ~x109 & ~x110 & ~x112 & ~x122 & ~x124 & ~x126 & ~x127 & ~x133 & ~x139 & ~x144 & ~x150 & ~x160 & ~x162 & ~x167 & ~x170 & ~x175 & ~x187 & ~x188 & ~x191 & ~x203 & ~x213 & ~x219 & ~x221 & ~x223 & ~x228 & ~x230 & ~x248 & ~x274 & ~x282 & ~x292 & ~x303 & ~x305 & ~x307 & ~x310 & ~x336 & ~x337 & ~x361 & ~x364 & ~x367 & ~x390 & ~x392 & ~x443 & ~x446 & ~x447 & ~x448 & ~x454 & ~x472 & ~x483 & ~x499 & ~x529 & ~x535 & ~x536 & ~x538 & ~x539 & ~x554 & ~x561 & ~x569 & ~x574 & ~x592 & ~x593 & ~x596 & ~x599 & ~x601 & ~x612 & ~x614 & ~x622 & ~x624 & ~x626 & ~x627 & ~x642 & ~x647 & ~x648 & ~x654 & ~x667 & ~x671 & ~x675 & ~x682 & ~x695 & ~x699 & ~x700 & ~x701 & ~x704 & ~x705 & ~x706 & ~x709 & ~x710 & ~x722 & ~x727 & ~x729 & ~x733 & ~x735 & ~x751 & ~x752 & ~x756 & ~x761 & ~x762 & ~x769 & ~x775 & ~x778 & ~x779 & ~x781;
assign c956 =  x279;
assign c958 =  x208 &  x235 & ~x15 & ~x17 & ~x22 & ~x26 & ~x33 & ~x37 & ~x39 & ~x40 & ~x47 & ~x50 & ~x57 & ~x61 & ~x64 & ~x69 & ~x76 & ~x78 & ~x86 & ~x87 & ~x96 & ~x97 & ~x105 & ~x108 & ~x113 & ~x124 & ~x125 & ~x134 & ~x175 & ~x176 & ~x177 & ~x189 & ~x192 & ~x200 & ~x201 & ~x203 & ~x218 & ~x222 & ~x228 & ~x251 & ~x253 & ~x281 & ~x304 & ~x311 & ~x319 & ~x333 & ~x335 & ~x337 & ~x361 & ~x388 & ~x389 & ~x390 & ~x392 & ~x419 & ~x471 & ~x473 & ~x474 & ~x478 & ~x499 & ~x500 & ~x507 & ~x528 & ~x533 & ~x534 & ~x583 & ~x601 & ~x610 & ~x611 & ~x614 & ~x618 & ~x620 & ~x623 & ~x624 & ~x641 & ~x648 & ~x649 & ~x655 & ~x669 & ~x677 & ~x680 & ~x681 & ~x709 & ~x710 & ~x711 & ~x712 & ~x721 & ~x731 & ~x739 & ~x743 & ~x752 & ~x758 & ~x761 & ~x763 & ~x767 & ~x771 & ~x775 & ~x776 & ~x779 & ~x781 & ~x782;
assign c960 =  x475;
assign c962 =  x291 &  x346 &  x379 & ~x6 & ~x8 & ~x15 & ~x35 & ~x41 & ~x42 & ~x43 & ~x46 & ~x47 & ~x53 & ~x76 & ~x89 & ~x91 & ~x95 & ~x97 & ~x112 & ~x113 & ~x116 & ~x120 & ~x126 & ~x129 & ~x130 & ~x132 & ~x134 & ~x150 & ~x152 & ~x160 & ~x164 & ~x166 & ~x171 & ~x174 & ~x175 & ~x176 & ~x178 & ~x188 & ~x194 & ~x216 & ~x217 & ~x221 & ~x222 & ~x223 & ~x224 & ~x225 & ~x226 & ~x228 & ~x230 & ~x248 & ~x255 & ~x261 & ~x273 & ~x274 & ~x276 & ~x281 & ~x282 & ~x307 & ~x314 & ~x315 & ~x333 & ~x336 & ~x342 & ~x360 & ~x362 & ~x364 & ~x367 & ~x386 & ~x388 & ~x390 & ~x395 & ~x414 & ~x415 & ~x423 & ~x424 & ~x426 & ~x427 & ~x445 & ~x452 & ~x467 & ~x479 & ~x480 & ~x500 & ~x502 & ~x506 & ~x507 & ~x510 & ~x535 & ~x539 & ~x618 & ~x619 & ~x621 & ~x638 & ~x644 & ~x669 & ~x670 & ~x672 & ~x693 & ~x695 & ~x696 & ~x700 & ~x728 & ~x757 & ~x773 & ~x781 & ~x782 & ~x783;
assign c964 =  x327 &  x354 &  x433 &  x437 & ~x6 & ~x55 & ~x59 & ~x133 & ~x148 & ~x163 & ~x192 & ~x202 & ~x203 & ~x221 & ~x223 & ~x254 & ~x389 & ~x396 & ~x444 & ~x472 & ~x567 & ~x604 & ~x645 & ~x670 & ~x697 & ~x714 & ~x741 & ~x754 & ~x766 & ~x771;
assign c966 =  x182 &  x183 & ~x2 & ~x10 & ~x11 & ~x17 & ~x20 & ~x21 & ~x24 & ~x31 & ~x32 & ~x44 & ~x47 & ~x49 & ~x52 & ~x60 & ~x66 & ~x67 & ~x74 & ~x75 & ~x77 & ~x79 & ~x82 & ~x85 & ~x89 & ~x95 & ~x96 & ~x98 & ~x100 & ~x102 & ~x105 & ~x112 & ~x122 & ~x132 & ~x134 & ~x138 & ~x145 & ~x148 & ~x149 & ~x159 & ~x161 & ~x171 & ~x176 & ~x197 & ~x203 & ~x222 & ~x223 & ~x229 & ~x230 & ~x247 & ~x248 & ~x250 & ~x255 & ~x256 & ~x275 & ~x276 & ~x279 & ~x285 & ~x303 & ~x310 & ~x331 & ~x333 & ~x336 & ~x339 & ~x349 & ~x361 & ~x365 & ~x387 & ~x391 & ~x415 & ~x416 & ~x420 & ~x443 & ~x451 & ~x476 & ~x478 & ~x498 & ~x500 & ~x502 & ~x524 & ~x525 & ~x533 & ~x537 & ~x553 & ~x557 & ~x564 & ~x569 & ~x595 & ~x596 & ~x599 & ~x610 & ~x611 & ~x618 & ~x620 & ~x623 & ~x639 & ~x648 & ~x669 & ~x670 & ~x671 & ~x672 & ~x676 & ~x678 & ~x680 & ~x681 & ~x698 & ~x699 & ~x700 & ~x704 & ~x707 & ~x723 & ~x724 & ~x729 & ~x730 & ~x731 & ~x737 & ~x744 & ~x746 & ~x749 & ~x750 & ~x752 & ~x757 & ~x766 & ~x774 & ~x782;
assign c968 =  x238 &  x290 &  x438 &  x458 & ~x0 & ~x2 & ~x4 & ~x7 & ~x10 & ~x17 & ~x19 & ~x36 & ~x61 & ~x63 & ~x93 & ~x104 & ~x105 & ~x107 & ~x109 & ~x110 & ~x115 & ~x120 & ~x125 & ~x126 & ~x172 & ~x196 & ~x204 & ~x224 & ~x230 & ~x249 & ~x309 & ~x310 & ~x332 & ~x360 & ~x392 & ~x417 & ~x423 & ~x445 & ~x446 & ~x447 & ~x476 & ~x502 & ~x532 & ~x561 & ~x565 & ~x566 & ~x569 & ~x587 & ~x592 & ~x598 & ~x619 & ~x622 & ~x623 & ~x647 & ~x649 & ~x667 & ~x669 & ~x701 & ~x704 & ~x705 & ~x706 & ~x723 & ~x726 & ~x753 & ~x756 & ~x759 & ~x763 & ~x766 & ~x775 & ~x782 & ~x783;
assign c970 =  x35;
assign c972 =  x211 &  x352 &  x379 & ~x1 & ~x4 & ~x19 & ~x24 & ~x25 & ~x33 & ~x38 & ~x41 & ~x45 & ~x47 & ~x50 & ~x53 & ~x54 & ~x60 & ~x76 & ~x78 & ~x92 & ~x99 & ~x119 & ~x123 & ~x124 & ~x129 & ~x145 & ~x152 & ~x154 & ~x167 & ~x172 & ~x175 & ~x177 & ~x189 & ~x191 & ~x250 & ~x274 & ~x275 & ~x277 & ~x278 & ~x308 & ~x311 & ~x312 & ~x313 & ~x385 & ~x388 & ~x394 & ~x413 & ~x416 & ~x417 & ~x420 & ~x423 & ~x442 & ~x448 & ~x450 & ~x470 & ~x471 & ~x473 & ~x481 & ~x496 & ~x498 & ~x500 & ~x506 & ~x507 & ~x509 & ~x516 & ~x528 & ~x532 & ~x533 & ~x543 & ~x557 & ~x565 & ~x567 & ~x584 & ~x586 & ~x592 & ~x596 & ~x639 & ~x644 & ~x648 & ~x650 & ~x664 & ~x666 & ~x674 & ~x690 & ~x691 & ~x706 & ~x733 & ~x734 & ~x735 & ~x739 & ~x753 & ~x758 & ~x763 & ~x764 & ~x765 & ~x766 & ~x768 & ~x779;
assign c974 =  x214 & ~x30 & ~x32 & ~x34 & ~x41 & ~x50 & ~x65 & ~x67 & ~x68 & ~x69 & ~x78 & ~x92 & ~x101 & ~x107 & ~x108 & ~x131 & ~x132 & ~x143 & ~x147 & ~x153 & ~x165 & ~x176 & ~x178 & ~x201 & ~x205 & ~x221 & ~x230 & ~x234 & ~x250 & ~x253 & ~x332 & ~x333 & ~x369 & ~x388 & ~x397 & ~x415 & ~x417 & ~x419 & ~x422 & ~x424 & ~x450 & ~x470 & ~x476 & ~x477 & ~x522 & ~x526 & ~x530 & ~x535 & ~x550 & ~x568 & ~x576 & ~x604 & ~x605 & ~x608 & ~x630 & ~x631 & ~x632 & ~x639 & ~x657 & ~x658 & ~x659 & ~x685 & ~x687 & ~x689 & ~x703 & ~x712 & ~x718 & ~x724 & ~x725 & ~x730 & ~x731 & ~x745 & ~x761 & ~x765 & ~x779;
assign c976 =  x214 &  x328 &  x383 &  x411 & ~x14 & ~x19 & ~x24 & ~x28 & ~x36 & ~x40 & ~x57 & ~x72 & ~x81 & ~x95 & ~x131 & ~x132 & ~x135 & ~x147 & ~x149 & ~x162 & ~x163 & ~x168 & ~x195 & ~x251 & ~x255 & ~x276 & ~x278 & ~x283 & ~x333 & ~x476 & ~x500 & ~x564 & ~x618 & ~x688 & ~x697 & ~x704 & ~x740 & ~x741 & ~x742 & ~x753 & ~x754 & ~x763 & ~x779 & ~x781;
assign c978 = ~x1 & ~x3 & ~x5 & ~x6 & ~x7 & ~x8 & ~x12 & ~x14 & ~x22 & ~x23 & ~x27 & ~x28 & ~x30 & ~x31 & ~x34 & ~x35 & ~x36 & ~x38 & ~x41 & ~x42 & ~x43 & ~x51 & ~x53 & ~x54 & ~x55 & ~x62 & ~x64 & ~x65 & ~x66 & ~x67 & ~x71 & ~x75 & ~x80 & ~x84 & ~x87 & ~x89 & ~x95 & ~x104 & ~x106 & ~x111 & ~x119 & ~x120 & ~x124 & ~x126 & ~x127 & ~x130 & ~x132 & ~x133 & ~x141 & ~x143 & ~x145 & ~x147 & ~x149 & ~x159 & ~x163 & ~x166 & ~x167 & ~x169 & ~x171 & ~x186 & ~x190 & ~x199 & ~x202 & ~x215 & ~x219 & ~x220 & ~x226 & ~x228 & ~x229 & ~x246 & ~x247 & ~x252 & ~x256 & ~x258 & ~x273 & ~x274 & ~x275 & ~x283 & ~x303 & ~x307 & ~x308 & ~x310 & ~x314 & ~x329 & ~x332 & ~x339 & ~x340 & ~x342 & ~x343 & ~x359 & ~x360 & ~x361 & ~x365 & ~x372 & ~x385 & ~x388 & ~x391 & ~x392 & ~x397 & ~x398 & ~x413 & ~x415 & ~x417 & ~x418 & ~x420 & ~x421 & ~x424 & ~x425 & ~x426 & ~x428 & ~x441 & ~x442 & ~x452 & ~x456 & ~x469 & ~x470 & ~x471 & ~x476 & ~x479 & ~x480 & ~x485 & ~x501 & ~x505 & ~x506 & ~x507 & ~x510 & ~x517 & ~x522 & ~x524 & ~x527 & ~x530 & ~x532 & ~x533 & ~x534 & ~x540 & ~x543 & ~x550 & ~x557 & ~x559 & ~x561 & ~x562 & ~x563 & ~x565 & ~x566 & ~x581 & ~x588 & ~x590 & ~x595 & ~x596 & ~x606 & ~x609 & ~x610 & ~x613 & ~x614 & ~x617 & ~x618 & ~x622 & ~x625 & ~x637 & ~x643 & ~x647 & ~x648 & ~x650 & ~x651 & ~x663 & ~x666 & ~x669 & ~x671 & ~x672 & ~x691 & ~x699 & ~x702 & ~x703 & ~x707 & ~x722 & ~x724 & ~x725 & ~x727 & ~x728 & ~x730 & ~x735 & ~x737 & ~x739 & ~x744 & ~x745 & ~x749 & ~x750 & ~x755 & ~x756 & ~x757 & ~x759 & ~x762 & ~x775 & ~x782;
assign c980 =  x197;
assign c982 =  x265 &  x266 &  x316 &  x460 & ~x154 & ~x201 & ~x570;
assign c984 =  x668;
assign c986 =  x236 & ~x0 & ~x2 & ~x8 & ~x12 & ~x19 & ~x32 & ~x33 & ~x36 & ~x41 & ~x47 & ~x50 & ~x53 & ~x55 & ~x65 & ~x66 & ~x73 & ~x78 & ~x88 & ~x91 & ~x93 & ~x99 & ~x100 & ~x113 & ~x116 & ~x117 & ~x120 & ~x121 & ~x129 & ~x132 & ~x136 & ~x142 & ~x144 & ~x149 & ~x150 & ~x160 & ~x161 & ~x164 & ~x167 & ~x174 & ~x177 & ~x188 & ~x198 & ~x199 & ~x205 & ~x217 & ~x218 & ~x219 & ~x224 & ~x225 & ~x248 & ~x251 & ~x253 & ~x255 & ~x273 & ~x278 & ~x285 & ~x286 & ~x287 & ~x308 & ~x313 & ~x333 & ~x337 & ~x358 & ~x362 & ~x364 & ~x397 & ~x416 & ~x417 & ~x420 & ~x426 & ~x443 & ~x445 & ~x451 & ~x453 & ~x471 & ~x472 & ~x483 & ~x496 & ~x499 & ~x507 & ~x513 & ~x515 & ~x517 & ~x523 & ~x532 & ~x533 & ~x537 & ~x538 & ~x541 & ~x543 & ~x552 & ~x553 & ~x555 & ~x559 & ~x562 & ~x563 & ~x568 & ~x569 & ~x571 & ~x579 & ~x582 & ~x583 & ~x586 & ~x609 & ~x610 & ~x611 & ~x613 & ~x638 & ~x639 & ~x643 & ~x644 & ~x645 & ~x647 & ~x648 & ~x649 & ~x664 & ~x667 & ~x668 & ~x670 & ~x673 & ~x674 & ~x678 & ~x695 & ~x708 & ~x718 & ~x719 & ~x722 & ~x725 & ~x730 & ~x756 & ~x758 & ~x760 & ~x761 & ~x764;
assign c988 =  x340;
assign c990 = ~x0 & ~x12 & ~x19 & ~x20 & ~x24 & ~x27 & ~x35 & ~x38 & ~x40 & ~x42 & ~x46 & ~x48 & ~x50 & ~x55 & ~x64 & ~x67 & ~x70 & ~x76 & ~x93 & ~x95 & ~x98 & ~x116 & ~x139 & ~x141 & ~x142 & ~x148 & ~x151 & ~x152 & ~x155 & ~x160 & ~x164 & ~x178 & ~x179 & ~x194 & ~x203 & ~x206 & ~x216 & ~x218 & ~x228 & ~x232 & ~x233 & ~x247 & ~x248 & ~x250 & ~x253 & ~x257 & ~x258 & ~x273 & ~x275 & ~x277 & ~x304 & ~x309 & ~x330 & ~x338 & ~x356 & ~x358 & ~x364 & ~x383 & ~x385 & ~x393 & ~x395 & ~x418 & ~x425 & ~x427 & ~x438 & ~x444 & ~x453 & ~x478 & ~x483 & ~x484 & ~x497 & ~x502 & ~x509 & ~x528 & ~x531 & ~x540 & ~x544 & ~x557 & ~x561 & ~x565 & ~x568 & ~x585 & ~x593 & ~x607 & ~x613 & ~x614 & ~x616 & ~x618 & ~x621 & ~x636 & ~x642 & ~x669 & ~x670 & ~x677 & ~x695 & ~x699 & ~x703 & ~x710 & ~x732 & ~x738 & ~x748 & ~x751 & ~x755 & ~x756 & ~x763 & ~x781;
assign c992 =  x182 &  x183 &  x184 &  x409 &  x436 &  x464 & ~x2 & ~x11 & ~x14 & ~x15 & ~x17 & ~x25 & ~x34 & ~x36 & ~x41 & ~x43 & ~x45 & ~x49 & ~x54 & ~x55 & ~x57 & ~x59 & ~x67 & ~x68 & ~x76 & ~x79 & ~x81 & ~x84 & ~x86 & ~x96 & ~x102 & ~x110 & ~x111 & ~x112 & ~x118 & ~x121 & ~x132 & ~x135 & ~x136 & ~x137 & ~x142 & ~x148 & ~x149 & ~x160 & ~x161 & ~x162 & ~x163 & ~x175 & ~x176 & ~x192 & ~x194 & ~x197 & ~x199 & ~x201 & ~x202 & ~x203 & ~x204 & ~x219 & ~x223 & ~x224 & ~x227 & ~x230 & ~x231 & ~x248 & ~x252 & ~x253 & ~x256 & ~x266 & ~x274 & ~x275 & ~x276 & ~x279 & ~x280 & ~x282 & ~x307 & ~x310 & ~x311 & ~x313 & ~x330 & ~x334 & ~x336 & ~x338 & ~x339 & ~x358 & ~x366 & ~x369 & ~x389 & ~x393 & ~x397 & ~x415 & ~x416 & ~x418 & ~x419 & ~x420 & ~x426 & ~x440 & ~x441 & ~x444 & ~x445 & ~x447 & ~x454 & ~x468 & ~x470 & ~x474 & ~x479 & ~x480 & ~x481 & ~x482 & ~x495 & ~x499 & ~x505 & ~x509 & ~x525 & ~x530 & ~x534 & ~x536 & ~x537 & ~x538 & ~x540 & ~x552 & ~x555 & ~x556 & ~x559 & ~x565 & ~x567 & ~x568 & ~x579 & ~x585 & ~x589 & ~x594 & ~x595 & ~x608 & ~x610 & ~x613 & ~x614 & ~x616 & ~x618 & ~x619 & ~x620 & ~x621 & ~x622 & ~x638 & ~x639 & ~x640 & ~x641 & ~x642 & ~x643 & ~x647 & ~x649 & ~x663 & ~x664 & ~x668 & ~x672 & ~x692 & ~x694 & ~x695 & ~x699 & ~x700 & ~x707 & ~x717 & ~x720 & ~x724 & ~x731 & ~x734 & ~x736 & ~x742 & ~x746 & ~x747 & ~x750 & ~x751 & ~x761 & ~x764 & ~x765 & ~x766 & ~x767 & ~x770 & ~x772 & ~x780;
assign c994 =  x749;
assign c996 =  x378 & ~x1 & ~x2 & ~x3 & ~x6 & ~x15 & ~x20 & ~x22 & ~x24 & ~x25 & ~x26 & ~x28 & ~x31 & ~x36 & ~x39 & ~x43 & ~x46 & ~x47 & ~x49 & ~x58 & ~x59 & ~x64 & ~x68 & ~x73 & ~x76 & ~x77 & ~x79 & ~x80 & ~x81 & ~x94 & ~x97 & ~x98 & ~x106 & ~x107 & ~x109 & ~x112 & ~x117 & ~x118 & ~x125 & ~x130 & ~x131 & ~x135 & ~x136 & ~x141 & ~x147 & ~x150 & ~x152 & ~x163 & ~x165 & ~x176 & ~x177 & ~x178 & ~x192 & ~x193 & ~x200 & ~x204 & ~x205 & ~x224 & ~x225 & ~x228 & ~x230 & ~x249 & ~x254 & ~x255 & ~x257 & ~x258 & ~x279 & ~x282 & ~x284 & ~x285 & ~x306 & ~x312 & ~x335 & ~x393 & ~x415 & ~x416 & ~x419 & ~x421 & ~x424 & ~x427 & ~x446 & ~x448 & ~x451 & ~x453 & ~x455 & ~x456 & ~x457 & ~x466 & ~x477 & ~x478 & ~x483 & ~x487 & ~x494 & ~x512 & ~x513 & ~x514 & ~x521 & ~x529 & ~x537 & ~x538 & ~x540 & ~x541 & ~x548 & ~x549 & ~x551 & ~x556 & ~x557 & ~x558 & ~x559 & ~x562 & ~x576 & ~x579 & ~x585 & ~x586 & ~x587 & ~x588 & ~x592 & ~x605 & ~x608 & ~x610 & ~x615 & ~x632 & ~x633 & ~x643 & ~x647 & ~x661 & ~x666 & ~x668 & ~x691 & ~x694 & ~x699 & ~x716 & ~x719 & ~x721 & ~x725 & ~x747 & ~x753 & ~x757 & ~x758 & ~x760 & ~x761 & ~x762 & ~x769 & ~x773 & ~x777 & ~x783;
assign c998 =  x89;
assign c9100 =  x324 &  x378 & ~x2 & ~x4 & ~x7 & ~x11 & ~x13 & ~x14 & ~x15 & ~x23 & ~x26 & ~x29 & ~x30 & ~x40 & ~x52 & ~x53 & ~x57 & ~x58 & ~x65 & ~x66 & ~x67 & ~x71 & ~x74 & ~x77 & ~x78 & ~x85 & ~x89 & ~x96 & ~x97 & ~x109 & ~x113 & ~x114 & ~x115 & ~x116 & ~x118 & ~x123 & ~x133 & ~x134 & ~x137 & ~x139 & ~x141 & ~x142 & ~x145 & ~x146 & ~x148 & ~x154 & ~x155 & ~x158 & ~x160 & ~x161 & ~x167 & ~x168 & ~x170 & ~x172 & ~x173 & ~x174 & ~x186 & ~x193 & ~x194 & ~x195 & ~x218 & ~x220 & ~x224 & ~x226 & ~x245 & ~x254 & ~x256 & ~x257 & ~x274 & ~x275 & ~x276 & ~x281 & ~x284 & ~x285 & ~x304 & ~x307 & ~x311 & ~x312 & ~x330 & ~x340 & ~x361 & ~x389 & ~x391 & ~x419 & ~x420 & ~x423 & ~x424 & ~x440 & ~x447 & ~x450 & ~x474 & ~x478 & ~x481 & ~x489 & ~x502 & ~x507 & ~x508 & ~x509 & ~x510 & ~x511 & ~x512 & ~x517 & ~x529 & ~x530 & ~x531 & ~x536 & ~x544 & ~x555 & ~x559 & ~x561 & ~x562 & ~x563 & ~x570 & ~x582 & ~x584 & ~x586 & ~x588 & ~x592 & ~x593 & ~x596 & ~x615 & ~x617 & ~x623 & ~x624 & ~x638 & ~x639 & ~x642 & ~x644 & ~x647 & ~x651 & ~x670 & ~x676 & ~x678 & ~x694 & ~x695 & ~x696 & ~x706 & ~x726 & ~x727 & ~x728 & ~x729 & ~x735 & ~x739 & ~x756 & ~x760 & ~x765 & ~x768 & ~x780;
assign c9102 =  x238 & ~x0 & ~x15 & ~x28 & ~x37 & ~x53 & ~x63 & ~x66 & ~x68 & ~x70 & ~x74 & ~x75 & ~x80 & ~x84 & ~x94 & ~x102 & ~x114 & ~x119 & ~x127 & ~x130 & ~x133 & ~x139 & ~x147 & ~x152 & ~x154 & ~x162 & ~x168 & ~x170 & ~x180 & ~x203 & ~x206 & ~x207 & ~x224 & ~x233 & ~x254 & ~x259 & ~x275 & ~x279 & ~x287 & ~x305 & ~x307 & ~x331 & ~x335 & ~x339 & ~x365 & ~x370 & ~x424 & ~x449 & ~x451 & ~x455 & ~x499 & ~x507 & ~x508 & ~x509 & ~x525 & ~x528 & ~x556 & ~x566 & ~x571 & ~x579 & ~x580 & ~x586 & ~x590 & ~x597 & ~x605 & ~x607 & ~x609 & ~x617 & ~x622 & ~x624 & ~x635 & ~x643 & ~x645 & ~x648 & ~x651 & ~x694 & ~x699 & ~x705 & ~x719 & ~x728 & ~x730 & ~x731 & ~x736 & ~x745 & ~x748 & ~x750 & ~x751 & ~x753 & ~x759 & ~x773;
assign c9104 =  x238 &  x240 &  x290 &  x372 &  x432 & ~x46 & ~x59 & ~x68 & ~x74 & ~x82 & ~x89 & ~x93 & ~x94 & ~x99 & ~x118 & ~x125 & ~x128 & ~x143 & ~x145 & ~x154 & ~x162 & ~x226 & ~x255 & ~x393 & ~x473 & ~x502 & ~x568 & ~x593 & ~x611 & ~x639 & ~x645 & ~x649 & ~x650 & ~x692 & ~x704 & ~x727 & ~x728 & ~x730 & ~x764 & ~x765;
assign c9106 =  x209 &  x236 & ~x1 & ~x12 & ~x14 & ~x20 & ~x21 & ~x22 & ~x26 & ~x36 & ~x51 & ~x52 & ~x65 & ~x70 & ~x79 & ~x107 & ~x115 & ~x129 & ~x138 & ~x139 & ~x142 & ~x144 & ~x145 & ~x147 & ~x150 & ~x153 & ~x161 & ~x164 & ~x172 & ~x173 & ~x179 & ~x191 & ~x193 & ~x195 & ~x198 & ~x200 & ~x206 & ~x215 & ~x217 & ~x221 & ~x224 & ~x227 & ~x230 & ~x232 & ~x244 & ~x254 & ~x259 & ~x283 & ~x302 & ~x307 & ~x308 & ~x314 & ~x330 & ~x334 & ~x339 & ~x358 & ~x361 & ~x364 & ~x370 & ~x390 & ~x391 & ~x395 & ~x396 & ~x411 & ~x413 & ~x417 & ~x421 & ~x422 & ~x425 & ~x442 & ~x444 & ~x466 & ~x471 & ~x477 & ~x481 & ~x494 & ~x522 & ~x523 & ~x527 & ~x540 & ~x554 & ~x563 & ~x566 & ~x583 & ~x584 & ~x585 & ~x587 & ~x588 & ~x589 & ~x590 & ~x591 & ~x607 & ~x619 & ~x622 & ~x635 & ~x636 & ~x641 & ~x645 & ~x649 & ~x651 & ~x667 & ~x668 & ~x679 & ~x691 & ~x695 & ~x696 & ~x700 & ~x701 & ~x702 & ~x705 & ~x719 & ~x732 & ~x738 & ~x749 & ~x755 & ~x765 & ~x766 & ~x775 & ~x777;
assign c9108 =  x53;
assign c9110 =  x178 &  x259 &  x429 & ~x318;
assign c9112 =  x213 &  x409 &  x436 & ~x2 & ~x14 & ~x16 & ~x18 & ~x46 & ~x48 & ~x64 & ~x77 & ~x91 & ~x97 & ~x104 & ~x106 & ~x122 & ~x141 & ~x142 & ~x147 & ~x148 & ~x152 & ~x171 & ~x201 & ~x208 & ~x229 & ~x234 & ~x282 & ~x305 & ~x340 & ~x419 & ~x444 & ~x448 & ~x476 & ~x478 & ~x496 & ~x501 & ~x508 & ~x523 & ~x531 & ~x550 & ~x555 & ~x556 & ~x565 & ~x579 & ~x583 & ~x587 & ~x632 & ~x635 & ~x637 & ~x720 & ~x721 & ~x738 & ~x740 & ~x752 & ~x777 & ~x780;
assign c9114 = ~x12 & ~x13 & ~x45 & ~x54 & ~x62 & ~x74 & ~x95 & ~x103 & ~x108 & ~x112 & ~x116 & ~x119 & ~x126 & ~x127 & ~x132 & ~x146 & ~x147 & ~x162 & ~x168 & ~x190 & ~x199 & ~x223 & ~x224 & ~x225 & ~x227 & ~x310 & ~x321 & ~x333 & ~x337 & ~x346 & ~x373 & ~x387 & ~x403 & ~x416 & ~x478 & ~x503 & ~x533 & ~x562 & ~x575 & ~x594 & ~x601 & ~x602 & ~x630 & ~x651 & ~x654 & ~x655 & ~x656 & ~x671 & ~x672 & ~x682 & ~x683 & ~x685 & ~x705 & ~x707 & ~x709 & ~x712 & ~x714 & ~x724 & ~x728 & ~x741 & ~x750 & ~x760 & ~x769 & ~x781;
assign c9116 =  x1;
assign c9118 =  x667;
assign c9120 =  x740;
assign c9124 =  x241 &  x355 &  x428 & ~x154 & ~x232 & ~x257 & ~x509 & ~x594 & ~x595 & ~x606;
assign c9126 =  x280;
assign c9128 =  x504;
assign c9130 =  x407 & ~x7 & ~x12 & ~x15 & ~x32 & ~x37 & ~x53 & ~x58 & ~x74 & ~x88 & ~x89 & ~x108 & ~x114 & ~x117 & ~x120 & ~x125 & ~x134 & ~x150 & ~x170 & ~x172 & ~x173 & ~x174 & ~x178 & ~x221 & ~x223 & ~x231 & ~x249 & ~x281 & ~x282 & ~x284 & ~x288 & ~x334 & ~x340 & ~x343 & ~x359 & ~x361 & ~x390 & ~x399 & ~x411 & ~x422 & ~x424 & ~x440 & ~x451 & ~x453 & ~x465 & ~x469 & ~x474 & ~x475 & ~x495 & ~x527 & ~x529 & ~x532 & ~x536 & ~x539 & ~x541 & ~x557 & ~x558 & ~x561 & ~x562 & ~x565 & ~x567 & ~x575 & ~x577 & ~x578 & ~x580 & ~x584 & ~x586 & ~x605 & ~x608 & ~x616 & ~x632 & ~x637 & ~x666 & ~x674 & ~x677 & ~x694 & ~x705 & ~x722 & ~x726 & ~x743 & ~x745 & ~x749 & ~x758 & ~x769 & ~x770 & ~x779 & ~x781 & ~x782 & ~x783;
assign c9132 =  x206 &  x207 &  x353 &  x409 & ~x0 & ~x2 & ~x7 & ~x10 & ~x12 & ~x13 & ~x35 & ~x40 & ~x42 & ~x44 & ~x48 & ~x52 & ~x55 & ~x58 & ~x63 & ~x66 & ~x67 & ~x72 & ~x88 & ~x98 & ~x114 & ~x115 & ~x120 & ~x128 & ~x129 & ~x132 & ~x134 & ~x137 & ~x138 & ~x143 & ~x146 & ~x157 & ~x158 & ~x160 & ~x161 & ~x162 & ~x168 & ~x173 & ~x186 & ~x188 & ~x191 & ~x194 & ~x195 & ~x200 & ~x216 & ~x217 & ~x218 & ~x222 & ~x224 & ~x244 & ~x247 & ~x252 & ~x256 & ~x284 & ~x307 & ~x308 & ~x310 & ~x359 & ~x366 & ~x367 & ~x390 & ~x392 & ~x393 & ~x413 & ~x416 & ~x419 & ~x446 & ~x448 & ~x470 & ~x471 & ~x473 & ~x480 & ~x500 & ~x511 & ~x513 & ~x528 & ~x529 & ~x534 & ~x542 & ~x545 & ~x546 & ~x555 & ~x556 & ~x559 & ~x561 & ~x562 & ~x592 & ~x612 & ~x619 & ~x642 & ~x646 & ~x648 & ~x672 & ~x673 & ~x677 & ~x678 & ~x696 & ~x703 & ~x706 & ~x709 & ~x712 & ~x723 & ~x727 & ~x730 & ~x733 & ~x737 & ~x750 & ~x754 & ~x756 & ~x763 & ~x770 & ~x777;
assign c9134 =  x185 & ~x18 & ~x42 & ~x48 & ~x100 & ~x179 & ~x233 & ~x254 & ~x341 & ~x343 & ~x367 & ~x398 & ~x444 & ~x468 & ~x541 & ~x578 & ~x581 & ~x603 & ~x615 & ~x667 & ~x761;
assign c9136 =  x209 &  x210 & ~x3 & ~x9 & ~x13 & ~x14 & ~x16 & ~x20 & ~x21 & ~x24 & ~x25 & ~x29 & ~x33 & ~x35 & ~x40 & ~x41 & ~x42 & ~x44 & ~x45 & ~x46 & ~x48 & ~x50 & ~x51 & ~x52 & ~x58 & ~x61 & ~x69 & ~x75 & ~x76 & ~x77 & ~x78 & ~x80 & ~x84 & ~x87 & ~x89 & ~x95 & ~x98 & ~x99 & ~x103 & ~x106 & ~x110 & ~x111 & ~x114 & ~x121 & ~x122 & ~x124 & ~x129 & ~x130 & ~x132 & ~x133 & ~x134 & ~x142 & ~x143 & ~x144 & ~x146 & ~x148 & ~x157 & ~x158 & ~x164 & ~x165 & ~x170 & ~x172 & ~x173 & ~x174 & ~x175 & ~x186 & ~x188 & ~x189 & ~x190 & ~x191 & ~x196 & ~x197 & ~x200 & ~x202 & ~x215 & ~x217 & ~x218 & ~x226 & ~x247 & ~x248 & ~x249 & ~x257 & ~x265 & ~x274 & ~x275 & ~x277 & ~x278 & ~x279 & ~x282 & ~x283 & ~x284 & ~x303 & ~x304 & ~x309 & ~x332 & ~x336 & ~x337 & ~x339 & ~x360 & ~x361 & ~x364 & ~x365 & ~x366 & ~x416 & ~x418 & ~x424 & ~x441 & ~x443 & ~x452 & ~x453 & ~x469 & ~x471 & ~x475 & ~x476 & ~x480 & ~x482 & ~x498 & ~x502 & ~x505 & ~x507 & ~x508 & ~x509 & ~x510 & ~x526 & ~x531 & ~x532 & ~x533 & ~x538 & ~x545 & ~x554 & ~x557 & ~x561 & ~x563 & ~x582 & ~x583 & ~x592 & ~x594 & ~x595 & ~x609 & ~x611 & ~x612 & ~x613 & ~x615 & ~x619 & ~x637 & ~x638 & ~x639 & ~x640 & ~x645 & ~x648 & ~x649 & ~x650 & ~x651 & ~x652 & ~x667 & ~x670 & ~x672 & ~x673 & ~x675 & ~x679 & ~x700 & ~x705 & ~x712 & ~x722 & ~x725 & ~x727 & ~x730 & ~x731 & ~x734 & ~x735 & ~x737 & ~x738 & ~x747 & ~x756 & ~x760 & ~x763 & ~x765 & ~x766 & ~x768 & ~x771 & ~x772 & ~x773 & ~x774 & ~x779;
assign c9138 =  x708;
assign c9140 =  x211 &  x343 &  x411 & ~x1 & ~x2 & ~x4 & ~x5 & ~x6 & ~x7 & ~x9 & ~x11 & ~x12 & ~x14 & ~x15 & ~x16 & ~x18 & ~x21 & ~x22 & ~x23 & ~x28 & ~x33 & ~x37 & ~x39 & ~x43 & ~x44 & ~x45 & ~x50 & ~x53 & ~x54 & ~x62 & ~x63 & ~x64 & ~x66 & ~x68 & ~x72 & ~x73 & ~x74 & ~x75 & ~x76 & ~x79 & ~x81 & ~x83 & ~x88 & ~x90 & ~x92 & ~x98 & ~x99 & ~x102 & ~x106 & ~x107 & ~x110 & ~x111 & ~x113 & ~x114 & ~x117 & ~x118 & ~x119 & ~x122 & ~x123 & ~x124 & ~x128 & ~x130 & ~x131 & ~x133 & ~x141 & ~x142 & ~x144 & ~x149 & ~x150 & ~x164 & ~x167 & ~x174 & ~x176 & ~x177 & ~x192 & ~x193 & ~x197 & ~x198 & ~x201 & ~x202 & ~x204 & ~x221 & ~x222 & ~x248 & ~x249 & ~x250 & ~x255 & ~x257 & ~x278 & ~x282 & ~x283 & ~x284 & ~x305 & ~x333 & ~x337 & ~x340 & ~x361 & ~x362 & ~x364 & ~x367 & ~x368 & ~x388 & ~x389 & ~x393 & ~x394 & ~x417 & ~x444 & ~x472 & ~x473 & ~x475 & ~x476 & ~x477 & ~x498 & ~x499 & ~x503 & ~x505 & ~x506 & ~x527 & ~x528 & ~x532 & ~x533 & ~x534 & ~x555 & ~x558 & ~x560 & ~x563 & ~x564 & ~x582 & ~x587 & ~x590 & ~x591 & ~x593 & ~x597 & ~x610 & ~x611 & ~x616 & ~x620 & ~x621 & ~x623 & ~x624 & ~x625 & ~x637 & ~x639 & ~x640 & ~x643 & ~x645 & ~x646 & ~x647 & ~x648 & ~x649 & ~x651 & ~x652 & ~x668 & ~x671 & ~x672 & ~x674 & ~x677 & ~x678 & ~x679 & ~x680 & ~x694 & ~x698 & ~x704 & ~x721 & ~x724 & ~x725 & ~x730 & ~x732 & ~x735 & ~x747 & ~x749 & ~x755 & ~x762 & ~x763 & ~x765 & ~x767 & ~x769 & ~x770 & ~x771;
assign c9142 =  x484 &  x515 & ~x4 & ~x101 & ~x104 & ~x148 & ~x202 & ~x229 & ~x404 & ~x415 & ~x470 & ~x535 & ~x568 & ~x598 & ~x626 & ~x652;
assign c9144 =  x368;
assign c9146 =  x184 &  x437 & ~x0 & ~x5 & ~x12 & ~x16 & ~x21 & ~x24 & ~x25 & ~x33 & ~x35 & ~x41 & ~x42 & ~x44 & ~x45 & ~x46 & ~x49 & ~x60 & ~x66 & ~x73 & ~x85 & ~x87 & ~x91 & ~x97 & ~x99 & ~x104 & ~x105 & ~x106 & ~x110 & ~x123 & ~x133 & ~x134 & ~x136 & ~x137 & ~x151 & ~x165 & ~x171 & ~x175 & ~x177 & ~x192 & ~x196 & ~x198 & ~x201 & ~x222 & ~x224 & ~x268 & ~x275 & ~x280 & ~x294 & ~x295 & ~x313 & ~x335 & ~x359 & ~x364 & ~x365 & ~x393 & ~x396 & ~x414 & ~x419 & ~x424 & ~x449 & ~x470 & ~x471 & ~x474 & ~x480 & ~x504 & ~x507 & ~x532 & ~x558 & ~x561 & ~x565 & ~x578 & ~x579 & ~x580 & ~x585 & ~x591 & ~x594 & ~x597 & ~x609 & ~x616 & ~x635 & ~x636 & ~x637 & ~x650 & ~x674 & ~x692 & ~x723 & ~x726 & ~x737 & ~x740 & ~x743 & ~x748 & ~x757 & ~x758 & ~x759 & ~x761 & ~x783;
assign c9148 =  x55;
assign c9150 =  x212 & ~x10 & ~x29 & ~x38 & ~x64 & ~x113 & ~x142 & ~x151 & ~x176 & ~x199 & ~x204 & ~x205 & ~x219 & ~x220 & ~x229 & ~x253 & ~x255 & ~x295 & ~x339 & ~x340 & ~x359 & ~x440 & ~x478 & ~x501 & ~x507 & ~x555 & ~x561 & ~x562 & ~x570 & ~x578 & ~x598 & ~x615 & ~x623 & ~x645 & ~x661 & ~x676 & ~x690 & ~x691 & ~x709 & ~x751;
assign c9152 =  x31;
assign c9154 =  x210 &  x211 &  x435 &  x487 & ~x25 & ~x33 & ~x49 & ~x57 & ~x88 & ~x117 & ~x131 & ~x166 & ~x178 & ~x191 & ~x197 & ~x202 & ~x231 & ~x259 & ~x306 & ~x365 & ~x404 & ~x414 & ~x469 & ~x508 & ~x533 & ~x583 & ~x598 & ~x616 & ~x698 & ~x729 & ~x781;
assign c9156 =  x186 &  x187 &  x264 &  x400 & ~x205 & ~x229;
assign c9158 =  x379 &  x380 & ~x2 & ~x7 & ~x8 & ~x9 & ~x11 & ~x19 & ~x22 & ~x23 & ~x30 & ~x31 & ~x32 & ~x42 & ~x51 & ~x61 & ~x68 & ~x75 & ~x77 & ~x91 & ~x92 & ~x102 & ~x104 & ~x107 & ~x108 & ~x112 & ~x115 & ~x116 & ~x123 & ~x125 & ~x127 & ~x129 & ~x130 & ~x131 & ~x133 & ~x140 & ~x143 & ~x144 & ~x148 & ~x153 & ~x154 & ~x155 & ~x156 & ~x157 & ~x158 & ~x166 & ~x172 & ~x178 & ~x180 & ~x192 & ~x196 & ~x204 & ~x205 & ~x206 & ~x221 & ~x223 & ~x230 & ~x232 & ~x249 & ~x252 & ~x253 & ~x257 & ~x260 & ~x279 & ~x286 & ~x311 & ~x333 & ~x339 & ~x340 & ~x357 & ~x362 & ~x365 & ~x367 & ~x384 & ~x385 & ~x388 & ~x395 & ~x412 & ~x416 & ~x421 & ~x442 & ~x445 & ~x448 & ~x450 & ~x472 & ~x473 & ~x474 & ~x475 & ~x497 & ~x501 & ~x502 & ~x504 & ~x509 & ~x532 & ~x551 & ~x553 & ~x555 & ~x556 & ~x564 & ~x566 & ~x595 & ~x615 & ~x617 & ~x620 & ~x622 & ~x658 & ~x676 & ~x694 & ~x697 & ~x698 & ~x721 & ~x723 & ~x725 & ~x727 & ~x728 & ~x729 & ~x741 & ~x751 & ~x755 & ~x757 & ~x758 & ~x759 & ~x765 & ~x775;
assign c9160 =  x239 &  x317 &  x345 &  x401 &  x431 & ~x1 & ~x8 & ~x18 & ~x22 & ~x26 & ~x28 & ~x58 & ~x73 & ~x88 & ~x99 & ~x100 & ~x108 & ~x112 & ~x121 & ~x123 & ~x132 & ~x135 & ~x143 & ~x174 & ~x175 & ~x200 & ~x219 & ~x229 & ~x248 & ~x275 & ~x313 & ~x391 & ~x392 & ~x419 & ~x422 & ~x424 & ~x454 & ~x477 & ~x483 & ~x501 & ~x531 & ~x538 & ~x570 & ~x625 & ~x644 & ~x671 & ~x674 & ~x677 & ~x691 & ~x700 & ~x724 & ~x726 & ~x732 & ~x751 & ~x754 & ~x763 & ~x776;
assign c9162 =  x400 &  x428 &  x437 & ~x4 & ~x10 & ~x12 & ~x16 & ~x21 & ~x26 & ~x28 & ~x32 & ~x38 & ~x51 & ~x57 & ~x59 & ~x60 & ~x67 & ~x75 & ~x79 & ~x82 & ~x86 & ~x92 & ~x99 & ~x103 & ~x116 & ~x117 & ~x118 & ~x125 & ~x128 & ~x129 & ~x132 & ~x135 & ~x137 & ~x175 & ~x177 & ~x195 & ~x196 & ~x220 & ~x226 & ~x227 & ~x228 & ~x229 & ~x230 & ~x231 & ~x252 & ~x254 & ~x258 & ~x276 & ~x304 & ~x308 & ~x310 & ~x333 & ~x337 & ~x348 & ~x359 & ~x361 & ~x362 & ~x364 & ~x365 & ~x375 & ~x377 & ~x392 & ~x396 & ~x403 & ~x415 & ~x417 & ~x422 & ~x441 & ~x442 & ~x443 & ~x447 & ~x453 & ~x498 & ~x500 & ~x505 & ~x527 & ~x529 & ~x532 & ~x533 & ~x534 & ~x537 & ~x553 & ~x556 & ~x561 & ~x564 & ~x585 & ~x587 & ~x588 & ~x594 & ~x595 & ~x614 & ~x616 & ~x619 & ~x623 & ~x642 & ~x646 & ~x673 & ~x674 & ~x675 & ~x698 & ~x700 & ~x725 & ~x749 & ~x753 & ~x754 & ~x755 & ~x756 & ~x758 & ~x759 & ~x767 & ~x768 & ~x770 & ~x776 & ~x778 & ~x779 & ~x781;
assign c9164 =  x746;
assign c9166 =  x385 &  x396 &  x413;
assign c9168 =  x212 &  x355 &  x383 & ~x7 & ~x8 & ~x10 & ~x11 & ~x20 & ~x23 & ~x27 & ~x32 & ~x43 & ~x67 & ~x68 & ~x70 & ~x78 & ~x85 & ~x90 & ~x95 & ~x99 & ~x101 & ~x109 & ~x113 & ~x117 & ~x123 & ~x126 & ~x136 & ~x137 & ~x151 & ~x164 & ~x166 & ~x167 & ~x192 & ~x195 & ~x198 & ~x200 & ~x226 & ~x227 & ~x231 & ~x232 & ~x233 & ~x251 & ~x257 & ~x281 & ~x285 & ~x286 & ~x309 & ~x366 & ~x367 & ~x390 & ~x392 & ~x395 & ~x414 & ~x417 & ~x421 & ~x441 & ~x449 & ~x469 & ~x471 & ~x502 & ~x526 & ~x529 & ~x558 & ~x581 & ~x635 & ~x662 & ~x663 & ~x675 & ~x691 & ~x699 & ~x731 & ~x732 & ~x739 & ~x743 & ~x751 & ~x755 & ~x757 & ~x758 & ~x777 & ~x779;
assign c9170 =  x183 &  x184 &  x291 &  x382 &  x465 & ~x5 & ~x7 & ~x9 & ~x16 & ~x21 & ~x26 & ~x29 & ~x30 & ~x34 & ~x35 & ~x37 & ~x39 & ~x42 & ~x44 & ~x48 & ~x49 & ~x57 & ~x60 & ~x63 & ~x64 & ~x65 & ~x68 & ~x69 & ~x76 & ~x81 & ~x90 & ~x93 & ~x97 & ~x98 & ~x99 & ~x100 & ~x103 & ~x104 & ~x106 & ~x107 & ~x111 & ~x112 & ~x115 & ~x116 & ~x120 & ~x121 & ~x125 & ~x127 & ~x130 & ~x132 & ~x141 & ~x144 & ~x148 & ~x161 & ~x166 & ~x172 & ~x173 & ~x174 & ~x175 & ~x191 & ~x195 & ~x196 & ~x205 & ~x220 & ~x223 & ~x227 & ~x247 & ~x255 & ~x279 & ~x280 & ~x281 & ~x283 & ~x284 & ~x286 & ~x314 & ~x331 & ~x333 & ~x334 & ~x338 & ~x340 & ~x341 & ~x363 & ~x366 & ~x368 & ~x388 & ~x395 & ~x425 & ~x450 & ~x453 & ~x470 & ~x473 & ~x523 & ~x524 & ~x531 & ~x534 & ~x536 & ~x554 & ~x556 & ~x586 & ~x591 & ~x592 & ~x606 & ~x610 & ~x620 & ~x637 & ~x664 & ~x676 & ~x691 & ~x693 & ~x698 & ~x721 & ~x729 & ~x734 & ~x740 & ~x741 & ~x746 & ~x752 & ~x759 & ~x775 & ~x780 & ~x781;
assign c9172 =  x211 &  x212 &  x356 &  x411 & ~x4 & ~x18 & ~x24 & ~x29 & ~x32 & ~x47 & ~x48 & ~x49 & ~x54 & ~x59 & ~x60 & ~x61 & ~x62 & ~x75 & ~x79 & ~x90 & ~x92 & ~x94 & ~x104 & ~x106 & ~x107 & ~x117 & ~x121 & ~x124 & ~x165 & ~x166 & ~x177 & ~x192 & ~x193 & ~x201 & ~x202 & ~x220 & ~x229 & ~x249 & ~x253 & ~x281 & ~x306 & ~x310 & ~x312 & ~x323 & ~x338 & ~x339 & ~x366 & ~x389 & ~x390 & ~x423 & ~x445 & ~x476 & ~x477 & ~x499 & ~x500 & ~x501 & ~x502 & ~x508 & ~x531 & ~x532 & ~x560 & ~x568 & ~x582 & ~x609 & ~x617 & ~x618 & ~x637 & ~x642 & ~x646 & ~x672 & ~x695 & ~x720 & ~x723 & ~x727 & ~x729 & ~x736 & ~x742 & ~x751 & ~x752 & ~x757 & ~x758 & ~x760 & ~x761 & ~x769 & ~x774 & ~x777;
assign c9174 =  x235 &  x261 &  x344 & ~x15 & ~x40 & ~x44 & ~x61 & ~x71 & ~x74 & ~x76 & ~x78 & ~x80 & ~x92 & ~x116 & ~x124 & ~x131 & ~x140 & ~x148 & ~x150 & ~x186 & ~x191 & ~x192 & ~x215 & ~x257 & ~x305 & ~x368 & ~x386 & ~x398 & ~x417 & ~x426 & ~x453 & ~x473 & ~x476 & ~x478 & ~x529 & ~x533 & ~x534 & ~x535 & ~x568 & ~x572 & ~x594 & ~x614 & ~x623 & ~x624 & ~x654 & ~x674 & ~x698 & ~x722 & ~x738 & ~x756 & ~x764 & ~x778;
assign c9176 =  x211 &  x237 & ~x1 & ~x4 & ~x6 & ~x7 & ~x14 & ~x26 & ~x30 & ~x49 & ~x53 & ~x55 & ~x59 & ~x64 & ~x66 & ~x75 & ~x84 & ~x85 & ~x95 & ~x97 & ~x103 & ~x108 & ~x111 & ~x117 & ~x122 & ~x124 & ~x132 & ~x143 & ~x152 & ~x155 & ~x164 & ~x172 & ~x173 & ~x174 & ~x175 & ~x180 & ~x193 & ~x226 & ~x234 & ~x247 & ~x249 & ~x250 & ~x254 & ~x257 & ~x258 & ~x261 & ~x284 & ~x288 & ~x312 & ~x331 & ~x336 & ~x340 & ~x358 & ~x388 & ~x395 & ~x397 & ~x414 & ~x426 & ~x448 & ~x452 & ~x478 & ~x480 & ~x497 & ~x501 & ~x502 & ~x538 & ~x552 & ~x562 & ~x593 & ~x607 & ~x613 & ~x626 & ~x634 & ~x637 & ~x664 & ~x665 & ~x666 & ~x671 & ~x678 & ~x695 & ~x707 & ~x709 & ~x719 & ~x733 & ~x736 & ~x737 & ~x738 & ~x751 & ~x753 & ~x761 & ~x777;
assign c9178 =  x212 &  x380 &  x463 & ~x4 & ~x5 & ~x6 & ~x7 & ~x8 & ~x9 & ~x10 & ~x11 & ~x21 & ~x24 & ~x31 & ~x34 & ~x37 & ~x46 & ~x48 & ~x51 & ~x56 & ~x66 & ~x68 & ~x72 & ~x75 & ~x80 & ~x84 & ~x88 & ~x89 & ~x95 & ~x102 & ~x104 & ~x105 & ~x109 & ~x110 & ~x116 & ~x119 & ~x124 & ~x128 & ~x135 & ~x136 & ~x139 & ~x146 & ~x147 & ~x165 & ~x172 & ~x175 & ~x178 & ~x180 & ~x194 & ~x195 & ~x205 & ~x228 & ~x229 & ~x231 & ~x233 & ~x250 & ~x252 & ~x255 & ~x256 & ~x261 & ~x277 & ~x286 & ~x312 & ~x337 & ~x341 & ~x343 & ~x344 & ~x360 & ~x363 & ~x364 & ~x368 & ~x370 & ~x397 & ~x413 & ~x417 & ~x423 & ~x439 & ~x440 & ~x445 & ~x446 & ~x449 & ~x453 & ~x455 & ~x467 & ~x468 & ~x473 & ~x474 & ~x478 & ~x479 & ~x499 & ~x521 & ~x522 & ~x524 & ~x530 & ~x537 & ~x551 & ~x553 & ~x556 & ~x557 & ~x558 & ~x562 & ~x563 & ~x564 & ~x578 & ~x588 & ~x589 & ~x595 & ~x606 & ~x613 & ~x616 & ~x638 & ~x643 & ~x647 & ~x659 & ~x664 & ~x666 & ~x669 & ~x694 & ~x699 & ~x700 & ~x703 & ~x715 & ~x717 & ~x720 & ~x726 & ~x729 & ~x735 & ~x744 & ~x750 & ~x751 & ~x764 & ~x770 & ~x773 & ~x774 & ~x775 & ~x779 & ~x783;
assign c9180 =  x181 &  x182 &  x409 &  x437 & ~x9 & ~x34 & ~x42 & ~x57 & ~x58 & ~x84 & ~x125 & ~x130 & ~x139 & ~x143 & ~x169 & ~x172 & ~x174 & ~x176 & ~x200 & ~x218 & ~x222 & ~x255 & ~x256 & ~x259 & ~x275 & ~x292 & ~x312 & ~x360 & ~x394 & ~x443 & ~x471 & ~x530 & ~x535 & ~x552 & ~x580 & ~x608 & ~x613 & ~x623 & ~x637 & ~x665 & ~x677 & ~x733 & ~x743 & ~x748 & ~x774 & ~x777;
assign c9182 =  x380 &  x717 & ~x229 & ~x657;
assign c9184 =  x213 &  x382 & ~x68 & ~x104 & ~x111 & ~x180 & ~x196 & ~x231 & ~x232 & ~x296 & ~x442 & ~x444 & ~x541 & ~x550 & ~x605 & ~x745 & ~x782;
assign c9186 =  x209 &  x210 &  x373 & ~x24 & ~x27 & ~x28 & ~x30 & ~x54 & ~x57 & ~x61 & ~x71 & ~x75 & ~x92 & ~x99 & ~x101 & ~x106 & ~x113 & ~x117 & ~x122 & ~x125 & ~x129 & ~x137 & ~x142 & ~x143 & ~x147 & ~x160 & ~x171 & ~x187 & ~x224 & ~x228 & ~x230 & ~x292 & ~x320 & ~x334 & ~x337 & ~x338 & ~x366 & ~x392 & ~x395 & ~x396 & ~x417 & ~x420 & ~x426 & ~x427 & ~x448 & ~x452 & ~x475 & ~x480 & ~x483 & ~x499 & ~x502 & ~x507 & ~x509 & ~x511 & ~x514 & ~x539 & ~x559 & ~x566 & ~x583 & ~x588 & ~x608 & ~x664 & ~x671 & ~x676 & ~x677 & ~x696 & ~x700 & ~x721 & ~x730 & ~x732 & ~x749 & ~x750 & ~x767 & ~x770 & ~x772;
assign c9188 =  x210 & ~x12 & ~x24 & ~x142 & ~x159 & ~x199 & ~x202 & ~x244 & ~x276 & ~x304 & ~x315 & ~x356 & ~x411 & ~x412 & ~x451 & ~x466 & ~x482 & ~x493 & ~x550 & ~x570 & ~x576 & ~x621 & ~x633 & ~x659 & ~x706;
assign c9190 =  x208 &  x401 & ~x15 & ~x34 & ~x35 & ~x40 & ~x49 & ~x62 & ~x75 & ~x82 & ~x83 & ~x85 & ~x96 & ~x99 & ~x115 & ~x128 & ~x132 & ~x135 & ~x140 & ~x141 & ~x147 & ~x160 & ~x163 & ~x170 & ~x172 & ~x188 & ~x191 & ~x219 & ~x228 & ~x246 & ~x248 & ~x274 & ~x319 & ~x320 & ~x348 & ~x366 & ~x422 & ~x443 & ~x478 & ~x538 & ~x541 & ~x543 & ~x544 & ~x589 & ~x613 & ~x616 & ~x667 & ~x674 & ~x680 & ~x696 & ~x697 & ~x698 & ~x727 & ~x743 & ~x757 & ~x766 & ~x768 & ~x779;
assign c9192 =  x239 &  x355 &  x398 &  x459 & ~x82 & ~x89 & ~x155 & ~x156 & ~x278 & ~x282 & ~x389 & ~x423 & ~x504 & ~x535 & ~x566 & ~x568 & ~x701 & ~x727;
assign c9194 =  x370 & ~x158 & ~x188 & ~x218 & ~x319 & ~x372 & ~x374 & ~x600 & ~x602 & ~x655 & ~x656 & ~x683;
assign c9196 =  x206 &  x352 &  x662 & ~x185 & ~x256 & ~x715;
assign c9198 =  x214 &  x265 &  x456 & ~x26 & ~x109 & ~x110 & ~x115 & ~x164 & ~x205 & ~x207 & ~x252 & ~x259 & ~x390 & ~x415 & ~x422 & ~x470 & ~x507 & ~x566 & ~x617 & ~x662 & ~x724 & ~x766;
assign c9200 =  x692 &  x720;
assign c9202 =  x240 &  x403 & ~x65 & ~x178 & ~x206 & ~x231 & ~x232 & ~x548 & ~x549 & ~x568 & ~x644 & ~x687;
assign c9204 =  x210 &  x326 &  x354 &  x378 &  x409 & ~x8 & ~x29 & ~x111 & ~x145 & ~x150 & ~x191 & ~x202 & ~x224 & ~x248 & ~x393 & ~x418 & ~x419 & ~x482 & ~x513 & ~x523 & ~x535 & ~x542 & ~x589 & ~x596 & ~x622 & ~x671 & ~x704 & ~x718 & ~x723 & ~x732 & ~x761;
assign c9206 =  x240 &  x381 &  x406 &  x409 &  x437 & ~x17 & ~x18 & ~x29 & ~x33 & ~x50 & ~x81 & ~x84 & ~x91 & ~x94 & ~x102 & ~x117 & ~x140 & ~x153 & ~x166 & ~x177 & ~x193 & ~x203 & ~x205 & ~x221 & ~x224 & ~x259 & ~x277 & ~x394 & ~x418 & ~x502 & ~x505 & ~x525 & ~x561 & ~x570 & ~x594 & ~x652 & ~x702 & ~x703 & ~x725 & ~x731 & ~x756;
assign c9208 =  x211 &  x215 &  x409 &  x437 &  x464 &  x492 & ~x4 & ~x16 & ~x20 & ~x21 & ~x22 & ~x23 & ~x24 & ~x25 & ~x30 & ~x31 & ~x33 & ~x35 & ~x41 & ~x44 & ~x50 & ~x53 & ~x54 & ~x64 & ~x71 & ~x73 & ~x79 & ~x84 & ~x90 & ~x97 & ~x98 & ~x99 & ~x104 & ~x106 & ~x118 & ~x127 & ~x128 & ~x142 & ~x143 & ~x150 & ~x162 & ~x163 & ~x168 & ~x195 & ~x201 & ~x223 & ~x224 & ~x228 & ~x229 & ~x249 & ~x250 & ~x257 & ~x282 & ~x309 & ~x311 & ~x332 & ~x333 & ~x340 & ~x397 & ~x424 & ~x443 & ~x444 & ~x445 & ~x446 & ~x448 & ~x449 & ~x472 & ~x475 & ~x501 & ~x502 & ~x506 & ~x523 & ~x524 & ~x525 & ~x526 & ~x532 & ~x533 & ~x534 & ~x561 & ~x563 & ~x566 & ~x583 & ~x587 & ~x588 & ~x593 & ~x596 & ~x619 & ~x623 & ~x634 & ~x636 & ~x641 & ~x667 & ~x672 & ~x698 & ~x703 & ~x704 & ~x723 & ~x735 & ~x739 & ~x740 & ~x741 & ~x743 & ~x751 & ~x754 & ~x755 & ~x757 & ~x761 & ~x764 & ~x771 & ~x773 & ~x774 & ~x776 & ~x777;
assign c9210 =  x705;
assign c9212 =  x720;
assign c9214 =  x694;
assign c9216 =  x405 & ~x11 & ~x15 & ~x24 & ~x27 & ~x31 & ~x33 & ~x35 & ~x38 & ~x39 & ~x44 & ~x52 & ~x53 & ~x54 & ~x56 & ~x62 & ~x63 & ~x69 & ~x70 & ~x84 & ~x88 & ~x94 & ~x96 & ~x97 & ~x101 & ~x108 & ~x112 & ~x116 & ~x122 & ~x133 & ~x141 & ~x147 & ~x149 & ~x158 & ~x159 & ~x161 & ~x166 & ~x169 & ~x177 & ~x188 & ~x191 & ~x192 & ~x194 & ~x220 & ~x224 & ~x225 & ~x250 & ~x253 & ~x255 & ~x280 & ~x283 & ~x307 & ~x311 & ~x335 & ~x364 & ~x366 & ~x388 & ~x390 & ~x418 & ~x427 & ~x449 & ~x450 & ~x452 & ~x453 & ~x460 & ~x461 & ~x482 & ~x484 & ~x502 & ~x508 & ~x511 & ~x513 & ~x515 & ~x516 & ~x524 & ~x535 & ~x539 & ~x553 & ~x555 & ~x565 & ~x566 & ~x579 & ~x580 & ~x586 & ~x587 & ~x606 & ~x607 & ~x614 & ~x620 & ~x621 & ~x623 & ~x641 & ~x643 & ~x651 & ~x663 & ~x664 & ~x670 & ~x672 & ~x676 & ~x678 & ~x691 & ~x700 & ~x703 & ~x706 & ~x729 & ~x731 & ~x734 & ~x746 & ~x747 & ~x748 & ~x755 & ~x756 & ~x757 & ~x764 & ~x767 & ~x769 & ~x771 & ~x772 & ~x777 & ~x780 & ~x781 & ~x783;
assign c9218 =  x210 &  x409 & ~x0 & ~x3 & ~x10 & ~x12 & ~x17 & ~x18 & ~x19 & ~x26 & ~x31 & ~x34 & ~x35 & ~x36 & ~x37 & ~x38 & ~x39 & ~x47 & ~x48 & ~x49 & ~x50 & ~x51 & ~x56 & ~x58 & ~x64 & ~x69 & ~x70 & ~x75 & ~x76 & ~x80 & ~x82 & ~x83 & ~x84 & ~x86 & ~x88 & ~x89 & ~x90 & ~x91 & ~x92 & ~x103 & ~x111 & ~x113 & ~x114 & ~x115 & ~x116 & ~x118 & ~x120 & ~x123 & ~x124 & ~x125 & ~x127 & ~x129 & ~x133 & ~x135 & ~x138 & ~x140 & ~x141 & ~x144 & ~x148 & ~x162 & ~x169 & ~x172 & ~x174 & ~x191 & ~x198 & ~x201 & ~x203 & ~x219 & ~x225 & ~x230 & ~x246 & ~x249 & ~x251 & ~x252 & ~x253 & ~x254 & ~x255 & ~x257 & ~x281 & ~x282 & ~x306 & ~x307 & ~x320 & ~x330 & ~x331 & ~x339 & ~x364 & ~x365 & ~x367 & ~x386 & ~x388 & ~x389 & ~x390 & ~x393 & ~x394 & ~x397 & ~x413 & ~x414 & ~x416 & ~x420 & ~x424 & ~x441 & ~x442 & ~x445 & ~x447 & ~x451 & ~x469 & ~x472 & ~x498 & ~x508 & ~x525 & ~x529 & ~x533 & ~x537 & ~x553 & ~x554 & ~x563 & ~x564 & ~x583 & ~x585 & ~x592 & ~x609 & ~x618 & ~x620 & ~x622 & ~x624 & ~x628 & ~x629 & ~x642 & ~x646 & ~x648 & ~x665 & ~x669 & ~x673 & ~x674 & ~x680 & ~x695 & ~x697 & ~x699 & ~x704 & ~x705 & ~x710 & ~x711 & ~x722 & ~x723 & ~x724 & ~x726 & ~x729 & ~x735 & ~x738 & ~x752 & ~x753 & ~x759 & ~x769 & ~x772 & ~x775 & ~x777 & ~x778;
assign c9220 =  x723;
assign c9222 =  x0;
assign c9224 =  x7;
assign c9226 =  x323 & ~x10 & ~x18 & ~x24 & ~x34 & ~x42 & ~x55 & ~x57 & ~x61 & ~x62 & ~x63 & ~x64 & ~x66 & ~x67 & ~x68 & ~x69 & ~x73 & ~x74 & ~x77 & ~x78 & ~x82 & ~x83 & ~x84 & ~x87 & ~x88 & ~x91 & ~x93 & ~x94 & ~x99 & ~x105 & ~x107 & ~x110 & ~x117 & ~x120 & ~x121 & ~x123 & ~x124 & ~x128 & ~x129 & ~x136 & ~x138 & ~x140 & ~x141 & ~x144 & ~x146 & ~x147 & ~x149 & ~x158 & ~x162 & ~x163 & ~x164 & ~x167 & ~x169 & ~x171 & ~x176 & ~x187 & ~x190 & ~x192 & ~x195 & ~x199 & ~x200 & ~x218 & ~x219 & ~x222 & ~x223 & ~x224 & ~x229 & ~x231 & ~x245 & ~x246 & ~x250 & ~x252 & ~x255 & ~x273 & ~x277 & ~x278 & ~x281 & ~x284 & ~x285 & ~x286 & ~x302 & ~x304 & ~x305 & ~x308 & ~x312 & ~x331 & ~x332 & ~x334 & ~x335 & ~x341 & ~x357 & ~x358 & ~x359 & ~x362 & ~x364 & ~x366 & ~x369 & ~x384 & ~x388 & ~x389 & ~x390 & ~x395 & ~x396 & ~x397 & ~x398 & ~x413 & ~x414 & ~x418 & ~x420 & ~x423 & ~x440 & ~x445 & ~x449 & ~x450 & ~x461 & ~x468 & ~x469 & ~x474 & ~x476 & ~x477 & ~x478 & ~x481 & ~x482 & ~x488 & ~x495 & ~x496 & ~x499 & ~x500 & ~x502 & ~x504 & ~x508 & ~x516 & ~x522 & ~x524 & ~x525 & ~x530 & ~x532 & ~x533 & ~x534 & ~x535 & ~x540 & ~x543 & ~x560 & ~x565 & ~x584 & ~x586 & ~x588 & ~x591 & ~x610 & ~x617 & ~x635 & ~x639 & ~x642 & ~x648 & ~x651 & ~x662 & ~x664 & ~x666 & ~x670 & ~x675 & ~x677 & ~x678 & ~x691 & ~x698 & ~x699 & ~x702 & ~x703 & ~x708 & ~x718 & ~x721 & ~x727 & ~x731 & ~x732 & ~x734 & ~x746 & ~x750 & ~x752 & ~x753 & ~x754 & ~x761 & ~x764 & ~x767 & ~x769 & ~x778;
assign c9228 =  x207 &  x411 &  x523 & ~x39 & ~x159 & ~x188 & ~x245 & ~x443 & ~x572 & ~x600 & ~x649;
assign c9230 =  x397 & ~x2 & ~x126 & ~x161 & ~x229 & ~x346 & ~x373 & ~x443;
assign c9232 =  x209 &  x372 &  x429 & ~x31 & ~x45 & ~x58 & ~x62 & ~x71 & ~x75 & ~x82 & ~x91 & ~x121 & ~x124 & ~x130 & ~x141 & ~x163 & ~x174 & ~x189 & ~x220 & ~x224 & ~x226 & ~x246 & ~x276 & ~x305 & ~x365 & ~x395 & ~x454 & ~x455 & ~x534 & ~x541 & ~x553 & ~x560 & ~x571 & ~x590 & ~x596 & ~x639 & ~x672 & ~x676 & ~x704 & ~x735 & ~x749 & ~x778;
assign c9234 =  x210 &  x212 & ~x4 & ~x26 & ~x31 & ~x35 & ~x40 & ~x52 & ~x53 & ~x58 & ~x69 & ~x72 & ~x79 & ~x88 & ~x94 & ~x97 & ~x107 & ~x108 & ~x110 & ~x115 & ~x137 & ~x140 & ~x152 & ~x164 & ~x177 & ~x178 & ~x218 & ~x225 & ~x229 & ~x246 & ~x252 & ~x257 & ~x267 & ~x280 & ~x294 & ~x303 & ~x307 & ~x309 & ~x310 & ~x312 & ~x334 & ~x340 & ~x341 & ~x359 & ~x419 & ~x447 & ~x474 & ~x477 & ~x480 & ~x502 & ~x527 & ~x529 & ~x537 & ~x538 & ~x552 & ~x564 & ~x565 & ~x584 & ~x586 & ~x592 & ~x598 & ~x607 & ~x609 & ~x613 & ~x616 & ~x644 & ~x649 & ~x663 & ~x666 & ~x671 & ~x672 & ~x724 & ~x726 & ~x728 & ~x731 & ~x744 & ~x748 & ~x751 & ~x753 & ~x763 & ~x768 & ~x777 & ~x780;
assign c9236 =  x182 &  x241 & ~x526 & ~x556 & ~x625 & ~x629 & ~x685 & ~x707 & ~x775;
assign c9238 =  x212 &  x404 & ~x3 & ~x6 & ~x14 & ~x15 & ~x35 & ~x53 & ~x71 & ~x94 & ~x95 & ~x101 & ~x106 & ~x107 & ~x118 & ~x124 & ~x135 & ~x138 & ~x154 & ~x155 & ~x156 & ~x179 & ~x180 & ~x191 & ~x192 & ~x198 & ~x199 & ~x204 & ~x227 & ~x229 & ~x231 & ~x396 & ~x419 & ~x453 & ~x454 & ~x499 & ~x514 & ~x538 & ~x539 & ~x540 & ~x552 & ~x555 & ~x566 & ~x567 & ~x579 & ~x594 & ~x604 & ~x616 & ~x631 & ~x632 & ~x648 & ~x664 & ~x726 & ~x762 & ~x775 & ~x780;
assign c9240 =  x184 & ~x6 & ~x7 & ~x16 & ~x19 & ~x20 & ~x23 & ~x33 & ~x45 & ~x50 & ~x52 & ~x60 & ~x61 & ~x62 & ~x72 & ~x86 & ~x87 & ~x90 & ~x97 & ~x102 & ~x103 & ~x105 & ~x107 & ~x112 & ~x113 & ~x114 & ~x117 & ~x125 & ~x126 & ~x127 & ~x128 & ~x138 & ~x140 & ~x143 & ~x148 & ~x150 & ~x164 & ~x166 & ~x173 & ~x176 & ~x193 & ~x194 & ~x202 & ~x220 & ~x221 & ~x231 & ~x247 & ~x251 & ~x253 & ~x256 & ~x284 & ~x296 & ~x305 & ~x338 & ~x349 & ~x362 & ~x365 & ~x366 & ~x377 & ~x387 & ~x394 & ~x415 & ~x417 & ~x419 & ~x422 & ~x444 & ~x446 & ~x473 & ~x500 & ~x508 & ~x528 & ~x531 & ~x534 & ~x556 & ~x557 & ~x558 & ~x559 & ~x583 & ~x596 & ~x599 & ~x613 & ~x614 & ~x615 & ~x620 & ~x622 & ~x623 & ~x624 & ~x626 & ~x638 & ~x640 & ~x648 & ~x653 & ~x671 & ~x672 & ~x681 & ~x695 & ~x705 & ~x706 & ~x709 & ~x710 & ~x711 & ~x723 & ~x731 & ~x733 & ~x734 & ~x739 & ~x749 & ~x758 & ~x762 & ~x767 & ~x768 & ~x773 & ~x774 & ~x777 & ~x781;
assign c9242 =  x380 & ~x1 & ~x4 & ~x8 & ~x10 & ~x11 & ~x12 & ~x14 & ~x15 & ~x21 & ~x22 & ~x23 & ~x26 & ~x29 & ~x30 & ~x32 & ~x34 & ~x36 & ~x37 & ~x40 & ~x43 & ~x44 & ~x45 & ~x47 & ~x50 & ~x51 & ~x54 & ~x55 & ~x58 & ~x63 & ~x73 & ~x78 & ~x86 & ~x87 & ~x89 & ~x93 & ~x94 & ~x97 & ~x100 & ~x103 & ~x104 & ~x105 & ~x108 & ~x110 & ~x111 & ~x114 & ~x118 & ~x122 & ~x125 & ~x127 & ~x128 & ~x133 & ~x143 & ~x158 & ~x159 & ~x161 & ~x163 & ~x165 & ~x167 & ~x168 & ~x169 & ~x171 & ~x173 & ~x174 & ~x175 & ~x176 & ~x184 & ~x186 & ~x188 & ~x189 & ~x190 & ~x195 & ~x197 & ~x199 & ~x200 & ~x202 & ~x217 & ~x222 & ~x227 & ~x229 & ~x242 & ~x243 & ~x245 & ~x246 & ~x247 & ~x249 & ~x252 & ~x255 & ~x256 & ~x258 & ~x271 & ~x272 & ~x273 & ~x278 & ~x280 & ~x284 & ~x285 & ~x300 & ~x305 & ~x306 & ~x311 & ~x331 & ~x333 & ~x336 & ~x337 & ~x340 & ~x355 & ~x356 & ~x357 & ~x361 & ~x364 & ~x367 & ~x383 & ~x384 & ~x385 & ~x390 & ~x393 & ~x394 & ~x396 & ~x397 & ~x412 & ~x414 & ~x417 & ~x419 & ~x423 & ~x424 & ~x425 & ~x440 & ~x444 & ~x451 & ~x452 & ~x453 & ~x455 & ~x468 & ~x469 & ~x471 & ~x472 & ~x473 & ~x474 & ~x477 & ~x483 & ~x484 & ~x497 & ~x502 & ~x504 & ~x505 & ~x509 & ~x512 & ~x525 & ~x528 & ~x532 & ~x533 & ~x535 & ~x538 & ~x553 & ~x555 & ~x559 & ~x560 & ~x565 & ~x566 & ~x567 & ~x568 & ~x583 & ~x584 & ~x588 & ~x589 & ~x595 & ~x610 & ~x611 & ~x612 & ~x614 & ~x617 & ~x618 & ~x619 & ~x622 & ~x638 & ~x641 & ~x642 & ~x643 & ~x651 & ~x667 & ~x669 & ~x672 & ~x674 & ~x676 & ~x677 & ~x679 & ~x680 & ~x694 & ~x701 & ~x702 & ~x705 & ~x709 & ~x738 & ~x748 & ~x749 & ~x758 & ~x762 & ~x773 & ~x774 & ~x775 & ~x781;
assign c9244 =  x209 &  x315 &  x342 &  x370 & ~x18 & ~x30 & ~x46 & ~x47 & ~x52 & ~x77 & ~x96 & ~x97 & ~x124 & ~x127 & ~x141 & ~x159 & ~x173 & ~x189 & ~x199 & ~x217 & ~x319 & ~x363 & ~x444 & ~x500 & ~x559 & ~x561 & ~x570 & ~x591 & ~x594 & ~x651 & ~x673 & ~x674 & ~x678 & ~x750 & ~x773 & ~x777 & ~x779 & ~x782;
assign c9246 =  x210 &  x290 &  x407 &  x434 & ~x2 & ~x11 & ~x15 & ~x19 & ~x21 & ~x28 & ~x37 & ~x42 & ~x44 & ~x46 & ~x52 & ~x57 & ~x59 & ~x60 & ~x64 & ~x74 & ~x78 & ~x84 & ~x87 & ~x93 & ~x98 & ~x109 & ~x112 & ~x113 & ~x115 & ~x117 & ~x118 & ~x128 & ~x130 & ~x133 & ~x135 & ~x140 & ~x141 & ~x142 & ~x145 & ~x159 & ~x160 & ~x161 & ~x167 & ~x171 & ~x174 & ~x187 & ~x194 & ~x195 & ~x196 & ~x197 & ~x198 & ~x199 & ~x203 & ~x205 & ~x218 & ~x219 & ~x221 & ~x222 & ~x223 & ~x232 & ~x246 & ~x249 & ~x250 & ~x257 & ~x258 & ~x278 & ~x279 & ~x282 & ~x304 & ~x306 & ~x307 & ~x308 & ~x310 & ~x312 & ~x336 & ~x338 & ~x359 & ~x360 & ~x365 & ~x387 & ~x388 & ~x415 & ~x426 & ~x447 & ~x454 & ~x471 & ~x472 & ~x475 & ~x478 & ~x481 & ~x503 & ~x510 & ~x516 & ~x532 & ~x537 & ~x544 & ~x557 & ~x558 & ~x566 & ~x581 & ~x582 & ~x583 & ~x586 & ~x587 & ~x592 & ~x613 & ~x616 & ~x624 & ~x635 & ~x644 & ~x645 & ~x647 & ~x650 & ~x666 & ~x667 & ~x676 & ~x693 & ~x694 & ~x697 & ~x698 & ~x702 & ~x706 & ~x723 & ~x748 & ~x753 & ~x754 & ~x755 & ~x759 & ~x760 & ~x761 & ~x768 & ~x769 & ~x776 & ~x777 & ~x778 & ~x782 & ~x783;
assign c9248 =  x455 & ~x18 & ~x130 & ~x191 & ~x229 & ~x334 & ~x374 & ~x376 & ~x422 & ~x602 & ~x629 & ~x630;
assign c9250 =  x208 &  x209 &  x409 &  x465 & ~x31 & ~x36 & ~x45 & ~x62 & ~x63 & ~x67 & ~x68 & ~x95 & ~x106 & ~x112 & ~x114 & ~x115 & ~x117 & ~x120 & ~x128 & ~x142 & ~x145 & ~x150 & ~x152 & ~x162 & ~x187 & ~x194 & ~x197 & ~x205 & ~x216 & ~x227 & ~x230 & ~x231 & ~x246 & ~x251 & ~x253 & ~x257 & ~x308 & ~x333 & ~x340 & ~x358 & ~x361 & ~x365 & ~x368 & ~x369 & ~x390 & ~x440 & ~x443 & ~x447 & ~x448 & ~x473 & ~x475 & ~x498 & ~x501 & ~x504 & ~x525 & ~x538 & ~x552 & ~x565 & ~x572 & ~x612 & ~x615 & ~x616 & ~x648 & ~x674 & ~x694 & ~x735 & ~x756 & ~x757 & ~x766 & ~x773 & ~x778;
assign c9252 =  x211 &  x263 &  x466 & ~x8 & ~x12 & ~x18 & ~x35 & ~x41 & ~x42 & ~x52 & ~x54 & ~x57 & ~x61 & ~x68 & ~x84 & ~x89 & ~x96 & ~x100 & ~x105 & ~x107 & ~x108 & ~x112 & ~x115 & ~x134 & ~x139 & ~x141 & ~x167 & ~x168 & ~x173 & ~x193 & ~x196 & ~x224 & ~x230 & ~x255 & ~x285 & ~x308 & ~x334 & ~x359 & ~x414 & ~x442 & ~x446 & ~x450 & ~x471 & ~x479 & ~x500 & ~x528 & ~x532 & ~x555 & ~x564 & ~x566 & ~x596 & ~x609 & ~x616 & ~x623 & ~x637 & ~x643 & ~x646 & ~x649 & ~x666 & ~x672 & ~x682 & ~x710 & ~x711 & ~x721 & ~x725 & ~x738 & ~x747 & ~x750 & ~x752 & ~x768 & ~x771 & ~x779 & ~x780;
assign c9254 =  x240 &  x266 & ~x1 & ~x6 & ~x7 & ~x16 & ~x25 & ~x30 & ~x32 & ~x38 & ~x45 & ~x48 & ~x52 & ~x57 & ~x71 & ~x75 & ~x84 & ~x92 & ~x100 & ~x101 & ~x109 & ~x114 & ~x117 & ~x134 & ~x149 & ~x154 & ~x156 & ~x160 & ~x183 & ~x194 & ~x201 & ~x206 & ~x209 & ~x228 & ~x230 & ~x231 & ~x253 & ~x262 & ~x279 & ~x343 & ~x392 & ~x414 & ~x443 & ~x447 & ~x468 & ~x480 & ~x496 & ~x501 & ~x524 & ~x529 & ~x532 & ~x537 & ~x550 & ~x554 & ~x605 & ~x618 & ~x644 & ~x665 & ~x701 & ~x702 & ~x731;
assign c9256 =  x209 &  x353 & ~x10 & ~x15 & ~x21 & ~x22 & ~x25 & ~x32 & ~x41 & ~x43 & ~x48 & ~x49 & ~x50 & ~x57 & ~x59 & ~x61 & ~x64 & ~x69 & ~x71 & ~x72 & ~x74 & ~x82 & ~x84 & ~x85 & ~x86 & ~x88 & ~x89 & ~x91 & ~x94 & ~x95 & ~x100 & ~x101 & ~x102 & ~x104 & ~x112 & ~x114 & ~x115 & ~x121 & ~x124 & ~x131 & ~x132 & ~x136 & ~x137 & ~x142 & ~x147 & ~x152 & ~x160 & ~x162 & ~x167 & ~x169 & ~x172 & ~x175 & ~x186 & ~x187 & ~x188 & ~x191 & ~x192 & ~x197 & ~x198 & ~x204 & ~x223 & ~x225 & ~x226 & ~x227 & ~x229 & ~x231 & ~x245 & ~x246 & ~x254 & ~x255 & ~x258 & ~x273 & ~x274 & ~x277 & ~x281 & ~x302 & ~x304 & ~x308 & ~x309 & ~x313 & ~x332 & ~x334 & ~x338 & ~x339 & ~x361 & ~x366 & ~x368 & ~x415 & ~x416 & ~x419 & ~x423 & ~x443 & ~x445 & ~x446 & ~x448 & ~x449 & ~x450 & ~x453 & ~x455 & ~x469 & ~x474 & ~x476 & ~x480 & ~x482 & ~x500 & ~x503 & ~x505 & ~x508 & ~x524 & ~x526 & ~x534 & ~x536 & ~x539 & ~x540 & ~x554 & ~x556 & ~x557 & ~x559 & ~x560 & ~x565 & ~x566 & ~x581 & ~x582 & ~x587 & ~x588 & ~x590 & ~x592 & ~x594 & ~x595 & ~x597 & ~x598 & ~x599 & ~x608 & ~x613 & ~x618 & ~x619 & ~x620 & ~x624 & ~x637 & ~x641 & ~x646 & ~x650 & ~x651 & ~x668 & ~x669 & ~x671 & ~x672 & ~x692 & ~x693 & ~x694 & ~x697 & ~x698 & ~x700 & ~x707 & ~x722 & ~x723 & ~x728 & ~x747 & ~x749 & ~x752 & ~x755 & ~x756 & ~x757 & ~x767 & ~x769 & ~x770 & ~x772 & ~x776 & ~x778 & ~x780 & ~x781 & ~x783;
assign c9258 =  x144;
assign c9260 =  x238 &  x404 & ~x3 & ~x5 & ~x6 & ~x15 & ~x41 & ~x43 & ~x66 & ~x83 & ~x85 & ~x87 & ~x90 & ~x95 & ~x98 & ~x119 & ~x121 & ~x124 & ~x127 & ~x129 & ~x130 & ~x134 & ~x148 & ~x149 & ~x152 & ~x153 & ~x155 & ~x156 & ~x158 & ~x159 & ~x161 & ~x169 & ~x173 & ~x174 & ~x178 & ~x202 & ~x203 & ~x204 & ~x221 & ~x250 & ~x255 & ~x279 & ~x280 & ~x285 & ~x307 & ~x312 & ~x364 & ~x388 & ~x419 & ~x443 & ~x444 & ~x457 & ~x472 & ~x502 & ~x504 & ~x508 & ~x511 & ~x527 & ~x535 & ~x540 & ~x567 & ~x595 & ~x605 & ~x612 & ~x616 & ~x632 & ~x637 & ~x663 & ~x671 & ~x673 & ~x677 & ~x678 & ~x697 & ~x704 & ~x705 & ~x723 & ~x731 & ~x748 & ~x750 & ~x751 & ~x763 & ~x764 & ~x769;
assign c9262 =  x89;
assign c9264 =  x180 &  x181 &  x234 &  x410 &  x493 & ~x6 & ~x12 & ~x13 & ~x17 & ~x18 & ~x23 & ~x25 & ~x27 & ~x28 & ~x29 & ~x36 & ~x37 & ~x38 & ~x40 & ~x52 & ~x54 & ~x56 & ~x63 & ~x69 & ~x70 & ~x76 & ~x83 & ~x84 & ~x87 & ~x89 & ~x91 & ~x94 & ~x96 & ~x99 & ~x101 & ~x104 & ~x107 & ~x108 & ~x111 & ~x114 & ~x116 & ~x117 & ~x119 & ~x121 & ~x134 & ~x138 & ~x147 & ~x160 & ~x171 & ~x172 & ~x174 & ~x175 & ~x176 & ~x195 & ~x196 & ~x203 & ~x225 & ~x231 & ~x250 & ~x251 & ~x254 & ~x256 & ~x265 & ~x275 & ~x278 & ~x303 & ~x305 & ~x307 & ~x308 & ~x309 & ~x310 & ~x312 & ~x313 & ~x333 & ~x335 & ~x337 & ~x340 & ~x361 & ~x362 & ~x363 & ~x365 & ~x367 & ~x368 & ~x369 & ~x387 & ~x388 & ~x393 & ~x397 & ~x416 & ~x421 & ~x422 & ~x423 & ~x442 & ~x443 & ~x447 & ~x451 & ~x470 & ~x471 & ~x472 & ~x476 & ~x477 & ~x481 & ~x497 & ~x498 & ~x500 & ~x504 & ~x505 & ~x506 & ~x507 & ~x533 & ~x534 & ~x536 & ~x542 & ~x558 & ~x560 & ~x561 & ~x582 & ~x591 & ~x611 & ~x612 & ~x616 & ~x618 & ~x619 & ~x640 & ~x642 & ~x667 & ~x668 & ~x671 & ~x672 & ~x673 & ~x695 & ~x696 & ~x697 & ~x698 & ~x702 & ~x721 & ~x723 & ~x724 & ~x733 & ~x735 & ~x737 & ~x738 & ~x739 & ~x743 & ~x745 & ~x746 & ~x751 & ~x752 & ~x753 & ~x758 & ~x760 & ~x768 & ~x769 & ~x770 & ~x773 & ~x776 & ~x779 & ~x781 & ~x783;
assign c9266 =  x214 &  x238 & ~x0 & ~x9 & ~x15 & ~x17 & ~x18 & ~x22 & ~x26 & ~x27 & ~x36 & ~x39 & ~x40 & ~x41 & ~x42 & ~x50 & ~x52 & ~x59 & ~x62 & ~x66 & ~x87 & ~x89 & ~x96 & ~x97 & ~x100 & ~x101 & ~x102 & ~x106 & ~x114 & ~x115 & ~x128 & ~x129 & ~x131 & ~x144 & ~x149 & ~x152 & ~x154 & ~x155 & ~x157 & ~x162 & ~x168 & ~x169 & ~x173 & ~x175 & ~x180 & ~x191 & ~x203 & ~x207 & ~x208 & ~x222 & ~x223 & ~x226 & ~x228 & ~x280 & ~x282 & ~x284 & ~x335 & ~x337 & ~x366 & ~x368 & ~x390 & ~x392 & ~x393 & ~x415 & ~x424 & ~x442 & ~x444 & ~x446 & ~x450 & ~x467 & ~x470 & ~x471 & ~x475 & ~x479 & ~x500 & ~x502 & ~x503 & ~x522 & ~x535 & ~x537 & ~x538 & ~x554 & ~x556 & ~x562 & ~x567 & ~x578 & ~x590 & ~x605 & ~x608 & ~x610 & ~x612 & ~x614 & ~x615 & ~x618 & ~x620 & ~x637 & ~x664 & ~x665 & ~x670 & ~x673 & ~x689 & ~x692 & ~x693 & ~x699 & ~x702 & ~x717 & ~x723 & ~x751 & ~x754 & ~x755 & ~x758 & ~x762 & ~x763 & ~x764 & ~x776 & ~x778;
assign c9268 =  x183 &  x380 &  x408 & ~x4 & ~x5 & ~x6 & ~x13 & ~x20 & ~x23 & ~x25 & ~x29 & ~x33 & ~x36 & ~x39 & ~x43 & ~x44 & ~x46 & ~x47 & ~x50 & ~x55 & ~x58 & ~x65 & ~x70 & ~x73 & ~x75 & ~x76 & ~x77 & ~x89 & ~x90 & ~x92 & ~x94 & ~x96 & ~x100 & ~x103 & ~x105 & ~x109 & ~x112 & ~x113 & ~x116 & ~x117 & ~x120 & ~x124 & ~x125 & ~x126 & ~x128 & ~x131 & ~x133 & ~x137 & ~x143 & ~x144 & ~x145 & ~x146 & ~x147 & ~x148 & ~x151 & ~x161 & ~x163 & ~x164 & ~x165 & ~x168 & ~x169 & ~x171 & ~x175 & ~x189 & ~x195 & ~x198 & ~x202 & ~x206 & ~x217 & ~x222 & ~x223 & ~x224 & ~x225 & ~x226 & ~x229 & ~x231 & ~x233 & ~x244 & ~x245 & ~x248 & ~x249 & ~x251 & ~x252 & ~x254 & ~x257 & ~x272 & ~x276 & ~x277 & ~x282 & ~x283 & ~x284 & ~x302 & ~x307 & ~x310 & ~x311 & ~x313 & ~x314 & ~x329 & ~x333 & ~x334 & ~x335 & ~x336 & ~x338 & ~x339 & ~x344 & ~x357 & ~x359 & ~x363 & ~x366 & ~x367 & ~x369 & ~x371 & ~x384 & ~x387 & ~x389 & ~x393 & ~x399 & ~x400 & ~x412 & ~x415 & ~x416 & ~x420 & ~x424 & ~x426 & ~x428 & ~x441 & ~x442 & ~x444 & ~x445 & ~x450 & ~x451 & ~x453 & ~x457 & ~x467 & ~x480 & ~x483 & ~x498 & ~x501 & ~x502 & ~x508 & ~x509 & ~x510 & ~x524 & ~x527 & ~x532 & ~x533 & ~x534 & ~x535 & ~x536 & ~x537 & ~x538 & ~x539 & ~x541 & ~x556 & ~x559 & ~x560 & ~x563 & ~x565 & ~x569 & ~x580 & ~x583 & ~x585 & ~x586 & ~x587 & ~x591 & ~x594 & ~x608 & ~x609 & ~x615 & ~x616 & ~x622 & ~x623 & ~x639 & ~x641 & ~x642 & ~x643 & ~x645 & ~x648 & ~x650 & ~x666 & ~x667 & ~x668 & ~x670 & ~x692 & ~x693 & ~x694 & ~x696 & ~x698 & ~x702 & ~x705 & ~x720 & ~x721 & ~x722 & ~x723 & ~x724 & ~x725 & ~x728 & ~x730 & ~x731 & ~x733 & ~x736 & ~x742 & ~x749 & ~x755 & ~x756 & ~x762 & ~x764 & ~x765 & ~x769 & ~x770 & ~x771 & ~x772 & ~x775 & ~x777 & ~x782;
assign c9270 =  x171;
assign c9272 =  x669;
assign c9274 =  x209 & ~x1 & ~x2 & ~x4 & ~x5 & ~x6 & ~x7 & ~x8 & ~x9 & ~x10 & ~x11 & ~x12 & ~x13 & ~x15 & ~x16 & ~x17 & ~x18 & ~x19 & ~x20 & ~x21 & ~x22 & ~x23 & ~x25 & ~x26 & ~x27 & ~x28 & ~x30 & ~x31 & ~x32 & ~x34 & ~x35 & ~x36 & ~x37 & ~x38 & ~x39 & ~x40 & ~x41 & ~x42 & ~x44 & ~x45 & ~x46 & ~x47 & ~x48 & ~x49 & ~x50 & ~x51 & ~x52 & ~x53 & ~x54 & ~x55 & ~x57 & ~x58 & ~x59 & ~x60 & ~x61 & ~x62 & ~x64 & ~x65 & ~x66 & ~x67 & ~x69 & ~x70 & ~x71 & ~x72 & ~x73 & ~x75 & ~x76 & ~x77 & ~x78 & ~x79 & ~x80 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x86 & ~x87 & ~x88 & ~x89 & ~x90 & ~x91 & ~x92 & ~x93 & ~x94 & ~x95 & ~x96 & ~x97 & ~x98 & ~x99 & ~x100 & ~x101 & ~x102 & ~x103 & ~x104 & ~x105 & ~x106 & ~x107 & ~x109 & ~x110 & ~x111 & ~x112 & ~x113 & ~x115 & ~x116 & ~x117 & ~x118 & ~x120 & ~x121 & ~x122 & ~x123 & ~x124 & ~x125 & ~x126 & ~x127 & ~x129 & ~x130 & ~x131 & ~x132 & ~x133 & ~x134 & ~x135 & ~x136 & ~x137 & ~x138 & ~x139 & ~x140 & ~x141 & ~x142 & ~x143 & ~x144 & ~x145 & ~x146 & ~x147 & ~x148 & ~x150 & ~x157 & ~x158 & ~x159 & ~x160 & ~x162 & ~x163 & ~x164 & ~x165 & ~x166 & ~x167 & ~x168 & ~x169 & ~x170 & ~x171 & ~x172 & ~x173 & ~x174 & ~x175 & ~x186 & ~x187 & ~x188 & ~x189 & ~x191 & ~x192 & ~x195 & ~x198 & ~x199 & ~x200 & ~x202 & ~x215 & ~x216 & ~x217 & ~x219 & ~x220 & ~x221 & ~x223 & ~x224 & ~x226 & ~x227 & ~x228 & ~x229 & ~x243 & ~x244 & ~x245 & ~x246 & ~x248 & ~x249 & ~x250 & ~x251 & ~x252 & ~x253 & ~x254 & ~x255 & ~x256 & ~x257 & ~x272 & ~x273 & ~x274 & ~x275 & ~x276 & ~x278 & ~x279 & ~x280 & ~x281 & ~x282 & ~x283 & ~x302 & ~x303 & ~x304 & ~x305 & ~x306 & ~x308 & ~x310 & ~x311 & ~x312 & ~x313 & ~x330 & ~x331 & ~x332 & ~x333 & ~x334 & ~x335 & ~x336 & ~x337 & ~x338 & ~x339 & ~x340 & ~x341 & ~x342 & ~x357 & ~x358 & ~x359 & ~x360 & ~x361 & ~x362 & ~x363 & ~x364 & ~x365 & ~x366 & ~x367 & ~x368 & ~x369 & ~x370 & ~x387 & ~x388 & ~x389 & ~x391 & ~x392 & ~x396 & ~x397 & ~x413 & ~x414 & ~x415 & ~x416 & ~x417 & ~x420 & ~x421 & ~x422 & ~x423 & ~x424 & ~x425 & ~x426 & ~x427 & ~x442 & ~x443 & ~x444 & ~x445 & ~x446 & ~x447 & ~x449 & ~x450 & ~x451 & ~x454 & ~x469 & ~x470 & ~x471 & ~x473 & ~x475 & ~x476 & ~x477 & ~x478 & ~x481 & ~x482 & ~x483 & ~x484 & ~x485 & ~x497 & ~x498 & ~x499 & ~x500 & ~x501 & ~x502 & ~x503 & ~x504 & ~x505 & ~x506 & ~x507 & ~x508 & ~x509 & ~x510 & ~x511 & ~x512 & ~x513 & ~x514 & ~x515 & ~x516 & ~x517 & ~x524 & ~x525 & ~x527 & ~x528 & ~x530 & ~x531 & ~x532 & ~x533 & ~x534 & ~x535 & ~x536 & ~x537 & ~x539 & ~x540 & ~x542 & ~x543 & ~x553 & ~x554 & ~x555 & ~x556 & ~x558 & ~x559 & ~x560 & ~x562 & ~x563 & ~x564 & ~x565 & ~x568 & ~x571 & ~x581 & ~x582 & ~x583 & ~x584 & ~x585 & ~x586 & ~x587 & ~x588 & ~x589 & ~x590 & ~x591 & ~x592 & ~x593 & ~x594 & ~x595 & ~x610 & ~x611 & ~x613 & ~x614 & ~x615 & ~x617 & ~x618 & ~x619 & ~x620 & ~x622 & ~x623 & ~x624 & ~x625 & ~x637 & ~x638 & ~x639 & ~x640 & ~x642 & ~x643 & ~x644 & ~x646 & ~x647 & ~x648 & ~x649 & ~x650 & ~x651 & ~x652 & ~x667 & ~x668 & ~x669 & ~x671 & ~x672 & ~x673 & ~x674 & ~x675 & ~x676 & ~x677 & ~x678 & ~x680 & ~x692 & ~x694 & ~x695 & ~x696 & ~x697 & ~x698 & ~x699 & ~x702 & ~x703 & ~x704 & ~x705 & ~x706 & ~x708 & ~x721 & ~x722 & ~x724 & ~x726 & ~x727 & ~x728 & ~x733 & ~x734 & ~x736 & ~x737 & ~x738 & ~x739 & ~x741 & ~x751 & ~x752 & ~x753 & ~x754 & ~x755 & ~x756 & ~x757 & ~x759 & ~x760 & ~x761 & ~x762 & ~x763 & ~x764 & ~x765 & ~x768 & ~x770 & ~x771 & ~x772 & ~x773 & ~x774 & ~x775 & ~x776 & ~x778 & ~x779 & ~x780 & ~x781 & ~x782 & ~x783;
assign c9276 =  x584;
assign c9278 =  x732;
assign c9280 =  x238 &  x433 &  x436 & ~x6 & ~x12 & ~x26 & ~x28 & ~x30 & ~x39 & ~x40 & ~x54 & ~x56 & ~x61 & ~x74 & ~x87 & ~x101 & ~x114 & ~x128 & ~x139 & ~x142 & ~x144 & ~x181 & ~x198 & ~x205 & ~x226 & ~x310 & ~x312 & ~x333 & ~x337 & ~x362 & ~x363 & ~x370 & ~x390 & ~x481 & ~x534 & ~x541 & ~x551 & ~x552 & ~x554 & ~x565 & ~x566 & ~x567 & ~x592 & ~x619 & ~x633 & ~x648 & ~x728 & ~x734 & ~x750 & ~x752 & ~x775 & ~x780;
assign c9282 = ~x15 & ~x45 & ~x48 & ~x57 & ~x79 & ~x158 & ~x175 & ~x185 & ~x201 & ~x215 & ~x246 & ~x255 & ~x309 & ~x310 & ~x347 & ~x415 & ~x447 & ~x528 & ~x548 & ~x603 & ~x625 & ~x632 & ~x652 & ~x653 & ~x670 & ~x671 & ~x680 & ~x763;
assign c9284 =  x488 & ~x0 & ~x1 & ~x21 & ~x25 & ~x27 & ~x29 & ~x40 & ~x48 & ~x60 & ~x66 & ~x74 & ~x77 & ~x96 & ~x116 & ~x126 & ~x127 & ~x139 & ~x140 & ~x143 & ~x144 & ~x147 & ~x163 & ~x166 & ~x171 & ~x174 & ~x189 & ~x193 & ~x229 & ~x252 & ~x254 & ~x332 & ~x361 & ~x362 & ~x393 & ~x403 & ~x443 & ~x451 & ~x479 & ~x528 & ~x530 & ~x546 & ~x558 & ~x563 & ~x594 & ~x600 & ~x601 & ~x616 & ~x653 & ~x676 & ~x680 & ~x682 & ~x711 & ~x713 & ~x736 & ~x764 & ~x781 & ~x782;
assign c9286 =  x239 &  x356 &  x412 & ~x7 & ~x13 & ~x18 & ~x33 & ~x58 & ~x61 & ~x71 & ~x84 & ~x105 & ~x123 & ~x130 & ~x149 & ~x162 & ~x173 & ~x192 & ~x201 & ~x228 & ~x256 & ~x283 & ~x295 & ~x389 & ~x582;
assign c9288 =  x207 &  x690 & ~x185 & ~x213;
assign c9290 =  x208 &  x342 & ~x2 & ~x4 & ~x28 & ~x34 & ~x44 & ~x46 & ~x47 & ~x52 & ~x56 & ~x58 & ~x64 & ~x81 & ~x83 & ~x88 & ~x95 & ~x99 & ~x101 & ~x103 & ~x105 & ~x111 & ~x115 & ~x117 & ~x125 & ~x134 & ~x135 & ~x139 & ~x164 & ~x172 & ~x192 & ~x198 & ~x219 & ~x226 & ~x227 & ~x248 & ~x249 & ~x256 & ~x278 & ~x279 & ~x292 & ~x304 & ~x305 & ~x306 & ~x319 & ~x333 & ~x345 & ~x347 & ~x348 & ~x361 & ~x362 & ~x394 & ~x421 & ~x444 & ~x472 & ~x499 & ~x505 & ~x532 & ~x535 & ~x556 & ~x558 & ~x560 & ~x563 & ~x564 & ~x587 & ~x591 & ~x625 & ~x648 & ~x649 & ~x679 & ~x701 & ~x708 & ~x728 & ~x733 & ~x747 & ~x757 & ~x762 & ~x763 & ~x764 & ~x767 & ~x769 & ~x770 & ~x775 & ~x783;
assign c9292 =  x584;
assign c9294 =  x728;
assign c9296 =  x346 &  x376 & ~x2 & ~x3 & ~x4 & ~x6 & ~x14 & ~x37 & ~x43 & ~x50 & ~x54 & ~x64 & ~x75 & ~x80 & ~x81 & ~x82 & ~x84 & ~x85 & ~x90 & ~x94 & ~x96 & ~x98 & ~x109 & ~x110 & ~x111 & ~x126 & ~x129 & ~x135 & ~x142 & ~x143 & ~x160 & ~x161 & ~x174 & ~x189 & ~x190 & ~x192 & ~x199 & ~x201 & ~x224 & ~x231 & ~x279 & ~x334 & ~x339 & ~x359 & ~x387 & ~x393 & ~x398 & ~x424 & ~x444 & ~x445 & ~x457 & ~x472 & ~x500 & ~x505 & ~x529 & ~x541 & ~x556 & ~x559 & ~x568 & ~x569 & ~x579 & ~x587 & ~x590 & ~x592 & ~x605 & ~x608 & ~x610 & ~x620 & ~x646 & ~x671 & ~x720 & ~x727 & ~x747 & ~x752 & ~x765 & ~x772;
assign c9298 =  x239 &  x406 &  x431 & ~x17 & ~x19 & ~x36 & ~x82 & ~x89 & ~x112 & ~x125 & ~x144 & ~x149 & ~x155 & ~x156 & ~x157 & ~x162 & ~x164 & ~x165 & ~x180 & ~x195 & ~x225 & ~x249 & ~x257 & ~x334 & ~x478 & ~x507 & ~x514 & ~x528 & ~x541 & ~x542 & ~x568 & ~x592 & ~x595 & ~x616 & ~x691 & ~x693 & ~x755 & ~x759 & ~x762;
assign c91 =  x433 &  x461 & ~x3 & ~x6 & ~x12 & ~x13 & ~x14 & ~x16 & ~x21 & ~x22 & ~x32 & ~x38 & ~x39 & ~x40 & ~x42 & ~x48 & ~x53 & ~x54 & ~x57 & ~x58 & ~x59 & ~x60 & ~x62 & ~x68 & ~x71 & ~x72 & ~x80 & ~x82 & ~x105 & ~x107 & ~x108 & ~x109 & ~x111 & ~x112 & ~x119 & ~x121 & ~x125 & ~x136 & ~x141 & ~x144 & ~x145 & ~x148 & ~x164 & ~x168 & ~x169 & ~x171 & ~x199 & ~x222 & ~x223 & ~x225 & ~x229 & ~x250 & ~x251 & ~x252 & ~x253 & ~x255 & ~x265 & ~x284 & ~x306 & ~x309 & ~x310 & ~x312 & ~x334 & ~x335 & ~x359 & ~x362 & ~x365 & ~x369 & ~x391 & ~x392 & ~x397 & ~x415 & ~x418 & ~x447 & ~x448 & ~x452 & ~x472 & ~x473 & ~x476 & ~x477 & ~x500 & ~x501 & ~x506 & ~x509 & ~x525 & ~x526 & ~x528 & ~x531 & ~x533 & ~x534 & ~x537 & ~x556 & ~x559 & ~x560 & ~x561 & ~x585 & ~x586 & ~x591 & ~x593 & ~x611 & ~x613 & ~x623 & ~x638 & ~x639 & ~x640 & ~x645 & ~x646 & ~x647 & ~x649 & ~x666 & ~x675 & ~x679 & ~x693 & ~x694 & ~x695 & ~x700 & ~x703 & ~x706 & ~x707 & ~x708 & ~x709 & ~x719 & ~x721 & ~x723 & ~x726 & ~x728 & ~x730 & ~x731 & ~x737 & ~x739 & ~x750 & ~x753 & ~x754 & ~x755 & ~x757 & ~x759 & ~x760 & ~x761 & ~x764 & ~x772 & ~x780 & ~x782;
assign c93 =  x443;
assign c95 =  x271 & ~x8 & ~x38 & ~x74 & ~x83 & ~x106 & ~x156 & ~x183 & ~x184 & ~x199 & ~x211 & ~x212 & ~x239 & ~x240 & ~x337 & ~x423 & ~x499 & ~x652 & ~x679 & ~x680 & ~x709 & ~x760 & ~x767 & ~x775;
assign c97 =  x602 & ~x4 & ~x12 & ~x13 & ~x14 & ~x18 & ~x23 & ~x28 & ~x31 & ~x36 & ~x43 & ~x47 & ~x54 & ~x57 & ~x60 & ~x63 & ~x75 & ~x76 & ~x77 & ~x85 & ~x88 & ~x112 & ~x115 & ~x122 & ~x132 & ~x141 & ~x145 & ~x160 & ~x162 & ~x197 & ~x198 & ~x308 & ~x311 & ~x338 & ~x349 & ~x377 & ~x378 & ~x393 & ~x405 & ~x418 & ~x419 & ~x420 & ~x421 & ~x432 & ~x433 & ~x447 & ~x473 & ~x478 & ~x488 & ~x507 & ~x533 & ~x558 & ~x587 & ~x588 & ~x590 & ~x609 & ~x613 & ~x618 & ~x620 & ~x637 & ~x639 & ~x640 & ~x667 & ~x669 & ~x679 & ~x691 & ~x719 & ~x725 & ~x727 & ~x728 & ~x730 & ~x734 & ~x747 & ~x754 & ~x756 & ~x769 & ~x782;
assign c99 =  x542 &  x570 & ~x2 & ~x3 & ~x7 & ~x10 & ~x14 & ~x15 & ~x16 & ~x29 & ~x34 & ~x35 & ~x37 & ~x50 & ~x52 & ~x54 & ~x59 & ~x61 & ~x62 & ~x67 & ~x72 & ~x77 & ~x80 & ~x86 & ~x88 & ~x93 & ~x95 & ~x108 & ~x109 & ~x113 & ~x114 & ~x116 & ~x132 & ~x139 & ~x141 & ~x144 & ~x147 & ~x149 & ~x162 & ~x164 & ~x166 & ~x170 & ~x171 & ~x172 & ~x190 & ~x194 & ~x196 & ~x201 & ~x223 & ~x250 & ~x252 & ~x280 & ~x283 & ~x285 & ~x307 & ~x308 & ~x309 & ~x310 & ~x336 & ~x337 & ~x338 & ~x363 & ~x365 & ~x366 & ~x418 & ~x419 & ~x446 & ~x450 & ~x477 & ~x501 & ~x502 & ~x503 & ~x530 & ~x531 & ~x532 & ~x533 & ~x534 & ~x560 & ~x562 & ~x587 & ~x589 & ~x591 & ~x592 & ~x615 & ~x618 & ~x620 & ~x648 & ~x650 & ~x662 & ~x664 & ~x674 & ~x676 & ~x678 & ~x679 & ~x692 & ~x694 & ~x702 & ~x705 & ~x706 & ~x716 & ~x717 & ~x723 & ~x726 & ~x727 & ~x732 & ~x736 & ~x740 & ~x741 & ~x744 & ~x745 & ~x750 & ~x752 & ~x759 & ~x760 & ~x762 & ~x763 & ~x767 & ~x770 & ~x772 & ~x774 & ~x777 & ~x778 & ~x781 & ~x782 & ~x783;
assign c911 =  x321 &  x348 &  x375 &  x601 & ~x419 & ~x423 & ~x504 & ~x674 & ~x687 & ~x717 & ~x737 & ~x740 & ~x751 & ~x758;
assign c913 = ~x4 & ~x5 & ~x10 & ~x24 & ~x35 & ~x36 & ~x37 & ~x38 & ~x41 & ~x51 & ~x61 & ~x79 & ~x81 & ~x85 & ~x91 & ~x104 & ~x115 & ~x142 & ~x143 & ~x156 & ~x182 & ~x192 & ~x227 & ~x254 & ~x278 & ~x281 & ~x307 & ~x310 & ~x334 & ~x376 & ~x377 & ~x404 & ~x414 & ~x415 & ~x416 & ~x433 & ~x460 & ~x500 & ~x514 & ~x526 & ~x528 & ~x530 & ~x539 & ~x557 & ~x561 & ~x564 & ~x568 & ~x618 & ~x620 & ~x646 & ~x648 & ~x664 & ~x667 & ~x669 & ~x692 & ~x723 & ~x730 & ~x731 & ~x733 & ~x748 & ~x753 & ~x759 & ~x766 & ~x783;
assign c915 = ~x46 & ~x97 & ~x194 & ~x287 & ~x291 & ~x292 & ~x315 & ~x317 & ~x342 & ~x424 & ~x674 & ~x705;
assign c917 =  x485 &  x568;
assign c919 = ~x0 & ~x1 & ~x3 & ~x5 & ~x10 & ~x28 & ~x35 & ~x37 & ~x41 & ~x55 & ~x65 & ~x66 & ~x71 & ~x77 & ~x82 & ~x83 & ~x107 & ~x114 & ~x116 & ~x135 & ~x136 & ~x142 & ~x143 & ~x151 & ~x174 & ~x179 & ~x187 & ~x207 & ~x224 & ~x235 & ~x254 & ~x276 & ~x305 & ~x307 & ~x336 & ~x361 & ~x362 & ~x363 & ~x389 & ~x392 & ~x424 & ~x443 & ~x445 & ~x446 & ~x452 & ~x475 & ~x500 & ~x502 & ~x503 & ~x504 & ~x507 & ~x532 & ~x534 & ~x560 & ~x561 & ~x585 & ~x587 & ~x593 & ~x595 & ~x611 & ~x615 & ~x617 & ~x620 & ~x622 & ~x624 & ~x639 & ~x645 & ~x667 & ~x670 & ~x674 & ~x677 & ~x680 & ~x700 & ~x703 & ~x709 & ~x711 & ~x713 & ~x714 & ~x715 & ~x716 & ~x717 & ~x720 & ~x721 & ~x724 & ~x734 & ~x740 & ~x741 & ~x742 & ~x743 & ~x745 & ~x752 & ~x758 & ~x759 & ~x761 & ~x768 & ~x782;
assign c921 =  x125;
assign c923 = ~x1 & ~x11 & ~x16 & ~x32 & ~x42 & ~x49 & ~x74 & ~x103 & ~x106 & ~x133 & ~x149 & ~x154 & ~x165 & ~x184 & ~x185 & ~x222 & ~x226 & ~x227 & ~x240 & ~x252 & ~x254 & ~x282 & ~x283 & ~x421 & ~x423 & ~x424 & ~x449 & ~x504 & ~x558 & ~x588 & ~x619 & ~x633 & ~x649 & ~x671 & ~x698 & ~x702 & ~x724 & ~x728 & ~x733 & ~x743 & ~x746 & ~x749 & ~x750 & ~x761 & ~x763 & ~x769 & ~x774 & ~x782;
assign c925 = ~x1 & ~x6 & ~x15 & ~x21 & ~x25 & ~x37 & ~x38 & ~x52 & ~x57 & ~x59 & ~x77 & ~x81 & ~x85 & ~x90 & ~x99 & ~x107 & ~x113 & ~x118 & ~x140 & ~x141 & ~x169 & ~x191 & ~x219 & ~x252 & ~x283 & ~x292 & ~x331 & ~x333 & ~x334 & ~x335 & ~x340 & ~x345 & ~x361 & ~x370 & ~x371 & ~x420 & ~x421 & ~x504 & ~x530 & ~x559 & ~x560 & ~x643 & ~x697 & ~x700 & ~x737 & ~x744 & ~x746 & ~x769 & ~x774;
assign c927 =  x434 & ~x0 & ~x9 & ~x29 & ~x37 & ~x39 & ~x42 & ~x44 & ~x57 & ~x59 & ~x60 & ~x66 & ~x69 & ~x70 & ~x72 & ~x80 & ~x86 & ~x94 & ~x109 & ~x114 & ~x116 & ~x124 & ~x137 & ~x142 & ~x151 & ~x167 & ~x168 & ~x171 & ~x175 & ~x195 & ~x221 & ~x250 & ~x255 & ~x256 & ~x284 & ~x301 & ~x305 & ~x306 & ~x311 & ~x331 & ~x332 & ~x337 & ~x354 & ~x357 & ~x358 & ~x362 & ~x364 & ~x365 & ~x366 & ~x388 & ~x390 & ~x391 & ~x416 & ~x421 & ~x444 & ~x450 & ~x451 & ~x454 & ~x473 & ~x475 & ~x504 & ~x533 & ~x558 & ~x590 & ~x592 & ~x611 & ~x614 & ~x641 & ~x665 & ~x667 & ~x675 & ~x676 & ~x680 & ~x681 & ~x682 & ~x700 & ~x716 & ~x717 & ~x718 & ~x725 & ~x733 & ~x735 & ~x736 & ~x740 & ~x741 & ~x742 & ~x743 & ~x748 & ~x751 & ~x752 & ~x756 & ~x763 & ~x779 & ~x780 & ~x782;
assign c929 =  x305;
assign c931 =  x497 & ~x11 & ~x17 & ~x20 & ~x34 & ~x54 & ~x57 & ~x84 & ~x89 & ~x114 & ~x116 & ~x136 & ~x143 & ~x198 & ~x220 & ~x313 & ~x422 & ~x505 & ~x531 & ~x584 & ~x611 & ~x615 & ~x643 & ~x666 & ~x693 & ~x696 & ~x712 & ~x713 & ~x714 & ~x720 & ~x721 & ~x730 & ~x733 & ~x743 & ~x748 & ~x750 & ~x756 & ~x765 & ~x773;
assign c933 = ~x9 & ~x32 & ~x66 & ~x76 & ~x77 & ~x95 & ~x96 & ~x117 & ~x148 & ~x251 & ~x256 & ~x277 & ~x291 & ~x306 & ~x310 & ~x312 & ~x316 & ~x317 & ~x319 & ~x342 & ~x367 & ~x419 & ~x444 & ~x505 & ~x555 & ~x558 & ~x695 & ~x722 & ~x726 & ~x753 & ~x758 & ~x764 & ~x765;
assign c935 = ~x2 & ~x17 & ~x23 & ~x31 & ~x34 & ~x39 & ~x43 & ~x60 & ~x63 & ~x78 & ~x80 & ~x83 & ~x85 & ~x89 & ~x90 & ~x101 & ~x106 & ~x108 & ~x109 & ~x133 & ~x136 & ~x137 & ~x179 & ~x180 & ~x194 & ~x198 & ~x209 & ~x237 & ~x266 & ~x335 & ~x337 & ~x364 & ~x417 & ~x447 & ~x474 & ~x504 & ~x506 & ~x528 & ~x530 & ~x533 & ~x536 & ~x559 & ~x595 & ~x597 & ~x644 & ~x653 & ~x679 & ~x682 & ~x699 & ~x701 & ~x704 & ~x707 & ~x708 & ~x710 & ~x724 & ~x729 & ~x734 & ~x737 & ~x738 & ~x740 & ~x752 & ~x759 & ~x763 & ~x776 & ~x782 & ~x783;
assign c937 = ~x0 & ~x5 & ~x10 & ~x11 & ~x13 & ~x16 & ~x21 & ~x24 & ~x58 & ~x61 & ~x64 & ~x83 & ~x89 & ~x97 & ~x109 & ~x110 & ~x111 & ~x148 & ~x200 & ~x228 & ~x326 & ~x337 & ~x338 & ~x352 & ~x382 & ~x411 & ~x449 & ~x472 & ~x483 & ~x620 & ~x639 & ~x642 & ~x648 & ~x735 & ~x744;
assign c939 = ~x352 & ~x353 & ~x382 & ~x384 & ~x426;
assign c941 = ~x6 & ~x14 & ~x16 & ~x39 & ~x40 & ~x43 & ~x50 & ~x57 & ~x64 & ~x69 & ~x73 & ~x74 & ~x75 & ~x78 & ~x80 & ~x85 & ~x95 & ~x99 & ~x102 & ~x105 & ~x116 & ~x136 & ~x138 & ~x140 & ~x142 & ~x157 & ~x164 & ~x165 & ~x176 & ~x185 & ~x195 & ~x199 & ~x213 & ~x223 & ~x224 & ~x251 & ~x257 & ~x258 & ~x259 & ~x281 & ~x282 & ~x284 & ~x285 & ~x296 & ~x306 & ~x308 & ~x312 & ~x323 & ~x361 & ~x417 & ~x449 & ~x451 & ~x471 & ~x478 & ~x480 & ~x504 & ~x508 & ~x529 & ~x530 & ~x531 & ~x536 & ~x557 & ~x558 & ~x587 & ~x591 & ~x611 & ~x612 & ~x616 & ~x617 & ~x639 & ~x642 & ~x643 & ~x646 & ~x650 & ~x664 & ~x673 & ~x679 & ~x691 & ~x692 & ~x698 & ~x700 & ~x701 & ~x706 & ~x718 & ~x720 & ~x721 & ~x735 & ~x737 & ~x738 & ~x740 & ~x742 & ~x743 & ~x746 & ~x751 & ~x753 & ~x756 & ~x769 & ~x770 & ~x771 & ~x773 & ~x779 & ~x783;
assign c943 =  x128;
assign c945 =  x269 & ~x1 & ~x10 & ~x13 & ~x22 & ~x23 & ~x26 & ~x27 & ~x31 & ~x35 & ~x40 & ~x41 & ~x42 & ~x44 & ~x58 & ~x60 & ~x62 & ~x67 & ~x78 & ~x81 & ~x83 & ~x92 & ~x101 & ~x113 & ~x119 & ~x120 & ~x121 & ~x123 & ~x125 & ~x130 & ~x132 & ~x138 & ~x139 & ~x143 & ~x146 & ~x148 & ~x155 & ~x157 & ~x165 & ~x170 & ~x172 & ~x191 & ~x222 & ~x250 & ~x279 & ~x282 & ~x306 & ~x332 & ~x333 & ~x349 & ~x350 & ~x360 & ~x365 & ~x367 & ~x377 & ~x387 & ~x392 & ~x414 & ~x417 & ~x419 & ~x421 & ~x425 & ~x432 & ~x443 & ~x450 & ~x459 & ~x460 & ~x468 & ~x471 & ~x475 & ~x486 & ~x501 & ~x502 & ~x529 & ~x533 & ~x534 & ~x536 & ~x555 & ~x560 & ~x567 & ~x568 & ~x581 & ~x586 & ~x587 & ~x588 & ~x593 & ~x595 & ~x608 & ~x611 & ~x618 & ~x620 & ~x636 & ~x641 & ~x646 & ~x664 & ~x701 & ~x703 & ~x721 & ~x725 & ~x728 & ~x757 & ~x761 & ~x773 & ~x781 & ~x783;
assign c947 =  x304;
assign c949 =  x220;
assign c951 =  x579 & ~x268 & ~x358;
assign c953 =  x264 & ~x1 & ~x7 & ~x10 & ~x14 & ~x17 & ~x20 & ~x23 & ~x28 & ~x35 & ~x37 & ~x45 & ~x52 & ~x54 & ~x59 & ~x73 & ~x82 & ~x89 & ~x91 & ~x93 & ~x95 & ~x96 & ~x97 & ~x98 & ~x104 & ~x117 & ~x120 & ~x137 & ~x141 & ~x145 & ~x146 & ~x150 & ~x151 & ~x165 & ~x169 & ~x170 & ~x175 & ~x191 & ~x192 & ~x193 & ~x278 & ~x334 & ~x336 & ~x337 & ~x361 & ~x376 & ~x405 & ~x415 & ~x419 & ~x421 & ~x423 & ~x433 & ~x455 & ~x475 & ~x476 & ~x478 & ~x479 & ~x484 & ~x502 & ~x504 & ~x505 & ~x510 & ~x512 & ~x514 & ~x530 & ~x540 & ~x555 & ~x563 & ~x567 & ~x581 & ~x586 & ~x587 & ~x591 & ~x594 & ~x615 & ~x618 & ~x619 & ~x643 & ~x648 & ~x649 & ~x670 & ~x674 & ~x675 & ~x700 & ~x701 & ~x703 & ~x704 & ~x726 & ~x748 & ~x751 & ~x752 & ~x755 & ~x761 & ~x765 & ~x766;
assign c955 = ~x12 & ~x14 & ~x79 & ~x84 & ~x114 & ~x134 & ~x151 & ~x180 & ~x196 & ~x209 & ~x403 & ~x432 & ~x446 & ~x451 & ~x460 & ~x484 & ~x486 & ~x487 & ~x504 & ~x506 & ~x534 & ~x560 & ~x584 & ~x645 & ~x695 & ~x728 & ~x762;
assign c957 = ~x12 & ~x18 & ~x19 & ~x54 & ~x78 & ~x86 & ~x89 & ~x117 & ~x120 & ~x134 & ~x155 & ~x165 & ~x168 & ~x173 & ~x179 & ~x191 & ~x220 & ~x334 & ~x336 & ~x349 & ~x375 & ~x391 & ~x402 & ~x403 & ~x404 & ~x419 & ~x430 & ~x457 & ~x458 & ~x475 & ~x500 & ~x506 & ~x564 & ~x586 & ~x588 & ~x593 & ~x614 & ~x666 & ~x698 & ~x700 & ~x726 & ~x727 & ~x779;
assign c959 =  x572 & ~x0 & ~x4 & ~x17 & ~x26 & ~x31 & ~x37 & ~x38 & ~x52 & ~x54 & ~x58 & ~x71 & ~x81 & ~x89 & ~x93 & ~x106 & ~x133 & ~x136 & ~x139 & ~x167 & ~x187 & ~x223 & ~x224 & ~x281 & ~x312 & ~x365 & ~x366 & ~x368 & ~x394 & ~x396 & ~x425 & ~x447 & ~x501 & ~x534 & ~x559 & ~x584 & ~x612 & ~x614 & ~x647 & ~x676 & ~x678 & ~x681 & ~x682 & ~x683 & ~x699 & ~x702 & ~x704 & ~x708 & ~x718 & ~x720 & ~x722 & ~x726 & ~x737 & ~x740 & ~x746 & ~x747 & ~x760 & ~x769 & ~x779;
assign c961 =  x241 &  x462 & ~x13 & ~x17 & ~x39 & ~x50 & ~x63 & ~x88 & ~x338 & ~x368 & ~x369 & ~x399 & ~x401 & ~x428 & ~x452 & ~x472 & ~x478 & ~x482 & ~x502 & ~x530 & ~x533 & ~x645 & ~x674 & ~x698 & ~x719 & ~x727;
assign c963 =  x630 & ~x94 & ~x111 & ~x121 & ~x325 & ~x326 & ~x336 & ~x366 & ~x370 & ~x452 & ~x505 & ~x669 & ~x700 & ~x713 & ~x714 & ~x780;
assign c965 =  x189 & ~x356;
assign c967 =  x231 &  x236 & ~x429 & ~x445 & ~x458;
assign c969 =  x577 &  x602 & ~x9 & ~x14 & ~x80 & ~x89 & ~x139 & ~x172 & ~x222 & ~x355 & ~x392 & ~x531 & ~x713 & ~x755 & ~x771;
assign c971 =  x517 &  x572 & ~x59 & ~x69 & ~x89 & ~x93 & ~x150 & ~x228 & ~x333 & ~x350 & ~x378 & ~x391 & ~x425 & ~x453 & ~x454 & ~x457 & ~x481 & ~x503 & ~x508 & ~x511 & ~x531 & ~x588 & ~x622 & ~x745 & ~x759 & ~x760;
assign c973 =  x594;
assign c975 =  x220;
assign c977 =  x571 &  x599 & ~x1 & ~x4 & ~x9 & ~x14 & ~x15 & ~x17 & ~x19 & ~x20 & ~x24 & ~x30 & ~x32 & ~x38 & ~x39 & ~x48 & ~x57 & ~x62 & ~x64 & ~x72 & ~x73 & ~x74 & ~x75 & ~x88 & ~x91 & ~x92 & ~x94 & ~x98 & ~x110 & ~x115 & ~x117 & ~x120 & ~x121 & ~x125 & ~x135 & ~x136 & ~x144 & ~x170 & ~x171 & ~x174 & ~x176 & ~x194 & ~x195 & ~x224 & ~x228 & ~x250 & ~x253 & ~x279 & ~x280 & ~x282 & ~x306 & ~x308 & ~x310 & ~x311 & ~x340 & ~x359 & ~x361 & ~x362 & ~x363 & ~x365 & ~x391 & ~x395 & ~x416 & ~x417 & ~x419 & ~x444 & ~x446 & ~x453 & ~x475 & ~x478 & ~x482 & ~x506 & ~x507 & ~x529 & ~x531 & ~x560 & ~x561 & ~x562 & ~x585 & ~x590 & ~x612 & ~x615 & ~x619 & ~x622 & ~x624 & ~x642 & ~x650 & ~x653 & ~x677 & ~x693 & ~x698 & ~x710 & ~x733 & ~x740 & ~x744 & ~x745 & ~x747 & ~x752 & ~x754 & ~x757 & ~x763 & ~x765 & ~x766 & ~x768 & ~x769 & ~x775;
assign c979 = ~x0 & ~x8 & ~x13 & ~x14 & ~x15 & ~x20 & ~x22 & ~x26 & ~x40 & ~x53 & ~x55 & ~x59 & ~x68 & ~x73 & ~x74 & ~x75 & ~x77 & ~x83 & ~x100 & ~x103 & ~x104 & ~x116 & ~x139 & ~x143 & ~x200 & ~x254 & ~x334 & ~x336 & ~x362 & ~x393 & ~x409 & ~x411 & ~x418 & ~x422 & ~x477 & ~x501 & ~x505 & ~x530 & ~x531 & ~x533 & ~x556 & ~x558 & ~x620 & ~x647 & ~x675 & ~x702 & ~x718 & ~x722 & ~x736 & ~x738 & ~x742 & ~x744 & ~x767 & ~x780 & ~x783;
assign c981 =  x185 &  x405 & ~x1 & ~x5 & ~x22 & ~x28 & ~x30 & ~x36 & ~x41 & ~x42 & ~x47 & ~x53 & ~x59 & ~x64 & ~x79 & ~x80 & ~x85 & ~x88 & ~x97 & ~x124 & ~x137 & ~x139 & ~x140 & ~x165 & ~x167 & ~x193 & ~x197 & ~x225 & ~x303 & ~x307 & ~x311 & ~x332 & ~x333 & ~x334 & ~x359 & ~x384 & ~x388 & ~x413 & ~x417 & ~x423 & ~x448 & ~x450 & ~x451 & ~x474 & ~x478 & ~x501 & ~x507 & ~x508 & ~x529 & ~x531 & ~x562 & ~x617 & ~x618 & ~x641 & ~x696 & ~x706 & ~x707 & ~x709 & ~x719 & ~x720 & ~x721 & ~x724 & ~x725 & ~x733 & ~x737 & ~x772 & ~x780;
assign c983 =  x549 & ~x12 & ~x30 & ~x60 & ~x224 & ~x278 & ~x280 & ~x341 & ~x369 & ~x370 & ~x391 & ~x395 & ~x409 & ~x500 & ~x531 & ~x589 & ~x638 & ~x664 & ~x675 & ~x692 & ~x708 & ~x709 & ~x716 & ~x719 & ~x738 & ~x752;
assign c985 = ~x0 & ~x4 & ~x5 & ~x14 & ~x16 & ~x24 & ~x26 & ~x38 & ~x42 & ~x43 & ~x47 & ~x57 & ~x58 & ~x62 & ~x70 & ~x73 & ~x77 & ~x79 & ~x85 & ~x89 & ~x90 & ~x93 & ~x98 & ~x105 & ~x112 & ~x115 & ~x119 & ~x132 & ~x140 & ~x147 & ~x153 & ~x167 & ~x171 & ~x182 & ~x201 & ~x210 & ~x229 & ~x238 & ~x251 & ~x255 & ~x258 & ~x266 & ~x280 & ~x306 & ~x309 & ~x363 & ~x365 & ~x366 & ~x367 & ~x393 & ~x445 & ~x447 & ~x499 & ~x502 & ~x506 & ~x527 & ~x532 & ~x533 & ~x534 & ~x536 & ~x538 & ~x555 & ~x561 & ~x570 & ~x584 & ~x587 & ~x591 & ~x597 & ~x598 & ~x616 & ~x618 & ~x620 & ~x640 & ~x644 & ~x646 & ~x650 & ~x654 & ~x674 & ~x675 & ~x678 & ~x680 & ~x699 & ~x727 & ~x732 & ~x734 & ~x737 & ~x741 & ~x742 & ~x744 & ~x745 & ~x746 & ~x758 & ~x762 & ~x764 & ~x772 & ~x773 & ~x774 & ~x780;
assign c987 =  x247;
assign c989 =  x513 &  x540 & ~x397 & ~x399;
assign c991 =  x655 &  x660 & ~x296 & ~x386 & ~x477;
assign c993 =  x235 & ~x26 & ~x40 & ~x45 & ~x104 & ~x106 & ~x113 & ~x141 & ~x143 & ~x165 & ~x168 & ~x193 & ~x226 & ~x310 & ~x349 & ~x361 & ~x374 & ~x428 & ~x454 & ~x472 & ~x534 & ~x667 & ~x674 & ~x699 & ~x724;
assign c995 =  x160;
assign c997 =  x158 & ~x329 & ~x544 & ~x572;
assign c999 =  x291 & ~x4 & ~x23 & ~x24 & ~x26 & ~x28 & ~x36 & ~x54 & ~x56 & ~x62 & ~x64 & ~x78 & ~x92 & ~x95 & ~x111 & ~x119 & ~x129 & ~x130 & ~x134 & ~x158 & ~x169 & ~x174 & ~x184 & ~x185 & ~x196 & ~x212 & ~x221 & ~x279 & ~x351 & ~x365 & ~x378 & ~x396 & ~x419 & ~x447 & ~x450 & ~x504 & ~x565 & ~x590 & ~x592 & ~x610 & ~x615 & ~x617 & ~x621 & ~x676 & ~x677 & ~x693 & ~x694 & ~x700 & ~x704 & ~x705 & ~x707 & ~x721 & ~x742 & ~x748 & ~x768;
assign c9101 = ~x0 & ~x8 & ~x10 & ~x13 & ~x16 & ~x18 & ~x23 & ~x24 & ~x25 & ~x27 & ~x29 & ~x36 & ~x38 & ~x39 & ~x40 & ~x41 & ~x42 & ~x43 & ~x49 & ~x52 & ~x54 & ~x60 & ~x61 & ~x66 & ~x72 & ~x79 & ~x80 & ~x82 & ~x86 & ~x87 & ~x94 & ~x102 & ~x106 & ~x108 & ~x109 & ~x113 & ~x116 & ~x128 & ~x136 & ~x141 & ~x152 & ~x154 & ~x163 & ~x167 & ~x168 & ~x169 & ~x181 & ~x182 & ~x194 & ~x196 & ~x197 & ~x198 & ~x209 & ~x210 & ~x237 & ~x238 & ~x250 & ~x251 & ~x252 & ~x253 & ~x266 & ~x278 & ~x280 & ~x281 & ~x306 & ~x307 & ~x338 & ~x363 & ~x364 & ~x420 & ~x421 & ~x422 & ~x450 & ~x474 & ~x476 & ~x503 & ~x504 & ~x506 & ~x527 & ~x528 & ~x558 & ~x561 & ~x562 & ~x584 & ~x588 & ~x593 & ~x594 & ~x596 & ~x612 & ~x617 & ~x619 & ~x622 & ~x624 & ~x640 & ~x643 & ~x644 & ~x645 & ~x649 & ~x671 & ~x676 & ~x679 & ~x680 & ~x682 & ~x700 & ~x703 & ~x704 & ~x705 & ~x706 & ~x708 & ~x719 & ~x728 & ~x736 & ~x751 & ~x754 & ~x755 & ~x756 & ~x757 & ~x762 & ~x763 & ~x764 & ~x766 & ~x774 & ~x777 & ~x778 & ~x782 & ~x783;
assign c9103 =  x98;
assign c9105 =  x581;
assign c9107 =  x460 &  x542 & ~x4 & ~x5 & ~x9 & ~x10 & ~x19 & ~x25 & ~x26 & ~x32 & ~x37 & ~x60 & ~x108 & ~x136 & ~x145 & ~x165 & ~x282 & ~x335 & ~x397 & ~x417 & ~x422 & ~x423 & ~x445 & ~x451 & ~x482 & ~x535 & ~x563 & ~x650 & ~x672 & ~x676 & ~x678 & ~x706 & ~x740 & ~x749 & ~x751 & ~x760 & ~x763 & ~x783;
assign c9109 =  x133;
assign c9111 =  x459 & ~x1 & ~x3 & ~x17 & ~x18 & ~x20 & ~x22 & ~x23 & ~x25 & ~x27 & ~x30 & ~x31 & ~x32 & ~x34 & ~x35 & ~x40 & ~x41 & ~x43 & ~x51 & ~x55 & ~x57 & ~x59 & ~x65 & ~x67 & ~x69 & ~x71 & ~x75 & ~x82 & ~x85 & ~x90 & ~x91 & ~x95 & ~x96 & ~x103 & ~x136 & ~x137 & ~x139 & ~x140 & ~x141 & ~x144 & ~x171 & ~x197 & ~x198 & ~x201 & ~x224 & ~x227 & ~x229 & ~x251 & ~x256 & ~x281 & ~x282 & ~x338 & ~x341 & ~x358 & ~x365 & ~x390 & ~x392 & ~x393 & ~x394 & ~x395 & ~x397 & ~x399 & ~x416 & ~x417 & ~x418 & ~x421 & ~x423 & ~x425 & ~x426 & ~x446 & ~x448 & ~x451 & ~x471 & ~x475 & ~x478 & ~x479 & ~x499 & ~x503 & ~x506 & ~x507 & ~x530 & ~x533 & ~x559 & ~x560 & ~x562 & ~x587 & ~x589 & ~x616 & ~x619 & ~x640 & ~x645 & ~x646 & ~x665 & ~x669 & ~x671 & ~x672 & ~x677 & ~x678 & ~x692 & ~x696 & ~x700 & ~x703 & ~x704 & ~x705 & ~x707 & ~x708 & ~x709 & ~x712 & ~x713 & ~x714 & ~x715 & ~x716 & ~x717 & ~x726 & ~x727 & ~x732 & ~x734 & ~x736 & ~x737 & ~x741 & ~x745 & ~x747 & ~x755 & ~x757 & ~x758 & ~x760 & ~x762 & ~x764 & ~x765 & ~x767 & ~x773 & ~x774 & ~x776 & ~x777 & ~x780 & ~x781;
assign c9113 = ~x8 & ~x17 & ~x21 & ~x29 & ~x30 & ~x35 & ~x37 & ~x39 & ~x40 & ~x41 & ~x42 & ~x47 & ~x48 & ~x49 & ~x50 & ~x53 & ~x55 & ~x57 & ~x61 & ~x63 & ~x79 & ~x113 & ~x142 & ~x172 & ~x186 & ~x197 & ~x200 & ~x202 & ~x229 & ~x232 & ~x241 & ~x253 & ~x258 & ~x259 & ~x261 & ~x278 & ~x280 & ~x283 & ~x419 & ~x448 & ~x450 & ~x451 & ~x476 & ~x480 & ~x503 & ~x527 & ~x529 & ~x532 & ~x533 & ~x560 & ~x564 & ~x586 & ~x588 & ~x613 & ~x615 & ~x617 & ~x639 & ~x643 & ~x648 & ~x668 & ~x670 & ~x672 & ~x673 & ~x689 & ~x693 & ~x694 & ~x700 & ~x703 & ~x705 & ~x713 & ~x714 & ~x716 & ~x719 & ~x720 & ~x721 & ~x723 & ~x724 & ~x727 & ~x731 & ~x734 & ~x739 & ~x740 & ~x742 & ~x745 & ~x747 & ~x751 & ~x753 & ~x757 & ~x761 & ~x775 & ~x778;
assign c9115 = ~x4 & ~x9 & ~x10 & ~x13 & ~x14 & ~x15 & ~x22 & ~x23 & ~x24 & ~x28 & ~x31 & ~x35 & ~x37 & ~x38 & ~x41 & ~x42 & ~x44 & ~x51 & ~x53 & ~x62 & ~x63 & ~x65 & ~x66 & ~x67 & ~x70 & ~x74 & ~x79 & ~x88 & ~x89 & ~x96 & ~x97 & ~x98 & ~x100 & ~x102 & ~x104 & ~x107 & ~x108 & ~x120 & ~x131 & ~x132 & ~x133 & ~x135 & ~x136 & ~x139 & ~x140 & ~x141 & ~x143 & ~x145 & ~x154 & ~x155 & ~x162 & ~x166 & ~x171 & ~x172 & ~x182 & ~x194 & ~x197 & ~x198 & ~x210 & ~x218 & ~x221 & ~x223 & ~x225 & ~x228 & ~x238 & ~x249 & ~x251 & ~x266 & ~x277 & ~x279 & ~x282 & ~x304 & ~x305 & ~x307 & ~x308 & ~x309 & ~x310 & ~x334 & ~x361 & ~x363 & ~x365 & ~x366 & ~x390 & ~x392 & ~x393 & ~x418 & ~x420 & ~x421 & ~x446 & ~x473 & ~x475 & ~x501 & ~x502 & ~x526 & ~x529 & ~x557 & ~x562 & ~x582 & ~x584 & ~x586 & ~x590 & ~x591 & ~x595 & ~x616 & ~x617 & ~x618 & ~x622 & ~x624 & ~x638 & ~x639 & ~x641 & ~x642 & ~x643 & ~x649 & ~x652 & ~x664 & ~x665 & ~x667 & ~x669 & ~x670 & ~x675 & ~x676 & ~x680 & ~x696 & ~x697 & ~x701 & ~x702 & ~x706 & ~x707 & ~x708 & ~x723 & ~x727 & ~x732 & ~x734 & ~x735 & ~x738 & ~x740 & ~x742 & ~x743 & ~x744 & ~x745 & ~x746 & ~x747 & ~x748 & ~x749 & ~x750 & ~x755 & ~x759 & ~x760 & ~x766 & ~x769 & ~x780 & ~x781 & ~x782;
assign c9117 =  x177 & ~x131 & ~x287 & ~x369 & ~x395;
assign c9119 =  x264 &  x266 & ~x0 & ~x1 & ~x8 & ~x21 & ~x25 & ~x36 & ~x43 & ~x46 & ~x49 & ~x53 & ~x60 & ~x63 & ~x67 & ~x71 & ~x75 & ~x88 & ~x89 & ~x95 & ~x130 & ~x140 & ~x161 & ~x163 & ~x166 & ~x168 & ~x170 & ~x176 & ~x177 & ~x199 & ~x249 & ~x276 & ~x304 & ~x307 & ~x309 & ~x361 & ~x375 & ~x376 & ~x389 & ~x402 & ~x418 & ~x421 & ~x443 & ~x447 & ~x448 & ~x450 & ~x457 & ~x479 & ~x481 & ~x482 & ~x486 & ~x534 & ~x537 & ~x558 & ~x566 & ~x568 & ~x582 & ~x585 & ~x593 & ~x615 & ~x616 & ~x621 & ~x647 & ~x669 & ~x670 & ~x675 & ~x676 & ~x693 & ~x702 & ~x703 & ~x749 & ~x755 & ~x762 & ~x765;
assign c9121 = ~x7 & ~x8 & ~x11 & ~x27 & ~x43 & ~x51 & ~x52 & ~x73 & ~x76 & ~x88 & ~x95 & ~x102 & ~x115 & ~x144 & ~x165 & ~x324 & ~x337 & ~x365 & ~x389 & ~x420 & ~x421 & ~x446 & ~x463 & ~x464 & ~x474 & ~x475 & ~x493 & ~x504 & ~x532 & ~x563 & ~x585 & ~x589 & ~x612 & ~x613 & ~x645 & ~x702 & ~x721 & ~x747 & ~x749 & ~x766 & ~x769 & ~x780;
assign c9123 =  x581 & ~x353 & ~x380;
assign c9125 =  x516 &  x629 &  x658 & ~x39 & ~x89 & ~x111 & ~x125 & ~x255 & ~x334 & ~x392 & ~x484 & ~x531 & ~x614 & ~x699 & ~x756;
assign c9127 =  x432 &  x433 &  x487 & ~x12 & ~x51 & ~x77 & ~x83 & ~x279 & ~x341 & ~x371 & ~x372 & ~x394 & ~x443 & ~x475 & ~x768;
assign c9129 = ~x6 & ~x10 & ~x12 & ~x13 & ~x21 & ~x23 & ~x32 & ~x42 & ~x43 & ~x46 & ~x75 & ~x78 & ~x82 & ~x84 & ~x85 & ~x89 & ~x92 & ~x105 & ~x108 & ~x112 & ~x114 & ~x130 & ~x137 & ~x138 & ~x142 & ~x143 & ~x157 & ~x167 & ~x172 & ~x185 & ~x196 & ~x201 & ~x212 & ~x213 & ~x222 & ~x224 & ~x240 & ~x241 & ~x268 & ~x278 & ~x295 & ~x296 & ~x304 & ~x308 & ~x335 & ~x339 & ~x361 & ~x366 & ~x367 & ~x420 & ~x422 & ~x423 & ~x449 & ~x474 & ~x475 & ~x476 & ~x478 & ~x479 & ~x501 & ~x503 & ~x533 & ~x535 & ~x562 & ~x563 & ~x564 & ~x583 & ~x584 & ~x585 & ~x595 & ~x610 & ~x621 & ~x638 & ~x639 & ~x644 & ~x646 & ~x648 & ~x650 & ~x666 & ~x667 & ~x675 & ~x689 & ~x690 & ~x691 & ~x693 & ~x694 & ~x698 & ~x699 & ~x703 & ~x705 & ~x727 & ~x730 & ~x734 & ~x737 & ~x738 & ~x741 & ~x742 & ~x746 & ~x754 & ~x756 & ~x757 & ~x769 & ~x772 & ~x776;
assign c9131 =  x405 &  x406 & ~x6 & ~x7 & ~x16 & ~x18 & ~x19 & ~x21 & ~x22 & ~x24 & ~x25 & ~x29 & ~x31 & ~x32 & ~x33 & ~x37 & ~x40 & ~x41 & ~x57 & ~x59 & ~x65 & ~x67 & ~x77 & ~x82 & ~x86 & ~x87 & ~x93 & ~x95 & ~x97 & ~x99 & ~x103 & ~x108 & ~x110 & ~x111 & ~x113 & ~x122 & ~x130 & ~x134 & ~x137 & ~x140 & ~x144 & ~x145 & ~x147 & ~x163 & ~x194 & ~x195 & ~x197 & ~x199 & ~x223 & ~x227 & ~x277 & ~x278 & ~x282 & ~x311 & ~x315 & ~x326 & ~x332 & ~x337 & ~x339 & ~x341 & ~x417 & ~x444 & ~x450 & ~x475 & ~x478 & ~x503 & ~x506 & ~x533 & ~x536 & ~x558 & ~x562 & ~x584 & ~x586 & ~x589 & ~x611 & ~x612 & ~x616 & ~x640 & ~x644 & ~x671 & ~x672 & ~x674 & ~x677 & ~x678 & ~x691 & ~x692 & ~x694 & ~x698 & ~x702 & ~x707 & ~x718 & ~x727 & ~x730 & ~x731 & ~x732 & ~x737 & ~x742 & ~x743 & ~x745 & ~x751 & ~x754 & ~x756 & ~x761 & ~x762 & ~x763 & ~x764 & ~x774 & ~x775 & ~x777;
assign c9133 =  x178 &  x462 & ~x399;
assign c9135 =  x347 & ~x354 & ~x517;
assign c9137 =  x461 &  x630 & ~x34 & ~x59 & ~x80 & ~x110 & ~x119 & ~x120 & ~x222 & ~x332 & ~x383 & ~x410 & ~x411 & ~x412 & ~x418 & ~x423 & ~x477 & ~x507 & ~x556 & ~x584 & ~x671 & ~x729 & ~x739 & ~x763 & ~x773;
assign c9141 =  x163;
assign c9143 = ~x2 & ~x68 & ~x306 & ~x317 & ~x320 & ~x346 & ~x371 & ~x385 & ~x398 & ~x624 & ~x737 & ~x749 & ~x750;
assign c9145 = ~x0 & ~x10 & ~x11 & ~x15 & ~x16 & ~x27 & ~x38 & ~x45 & ~x46 & ~x49 & ~x50 & ~x51 & ~x53 & ~x57 & ~x59 & ~x63 & ~x66 & ~x75 & ~x79 & ~x81 & ~x83 & ~x84 & ~x87 & ~x97 & ~x99 & ~x100 & ~x102 & ~x108 & ~x112 & ~x113 & ~x120 & ~x131 & ~x132 & ~x138 & ~x139 & ~x140 & ~x141 & ~x142 & ~x143 & ~x146 & ~x159 & ~x161 & ~x167 & ~x192 & ~x193 & ~x194 & ~x196 & ~x198 & ~x200 & ~x221 & ~x225 & ~x251 & ~x253 & ~x255 & ~x278 & ~x279 & ~x280 & ~x283 & ~x304 & ~x307 & ~x308 & ~x310 & ~x311 & ~x322 & ~x333 & ~x337 & ~x339 & ~x350 & ~x351 & ~x362 & ~x378 & ~x389 & ~x391 & ~x393 & ~x395 & ~x405 & ~x416 & ~x418 & ~x419 & ~x421 & ~x423 & ~x432 & ~x444 & ~x449 & ~x450 & ~x460 & ~x473 & ~x474 & ~x476 & ~x478 & ~x480 & ~x501 & ~x503 & ~x505 & ~x507 & ~x515 & ~x527 & ~x528 & ~x529 & ~x531 & ~x534 & ~x543 & ~x554 & ~x560 & ~x561 & ~x564 & ~x584 & ~x588 & ~x591 & ~x612 & ~x613 & ~x619 & ~x620 & ~x621 & ~x622 & ~x637 & ~x640 & ~x645 & ~x648 & ~x665 & ~x668 & ~x669 & ~x673 & ~x674 & ~x677 & ~x694 & ~x697 & ~x700 & ~x703 & ~x706 & ~x722 & ~x726 & ~x730 & ~x749 & ~x750 & ~x753 & ~x755 & ~x756 & ~x761 & ~x763 & ~x780 & ~x782;
assign c9147 =  x326 & ~x5 & ~x10 & ~x20 & ~x22 & ~x31 & ~x41 & ~x49 & ~x50 & ~x60 & ~x61 & ~x68 & ~x89 & ~x109 & ~x144 & ~x150 & ~x158 & ~x164 & ~x195 & ~x251 & ~x252 & ~x310 & ~x349 & ~x350 & ~x362 & ~x363 & ~x364 & ~x377 & ~x394 & ~x404 & ~x405 & ~x417 & ~x420 & ~x432 & ~x442 & ~x445 & ~x451 & ~x459 & ~x475 & ~x482 & ~x483 & ~x509 & ~x514 & ~x527 & ~x529 & ~x536 & ~x556 & ~x558 & ~x609 & ~x610 & ~x644 & ~x649 & ~x693 & ~x722 & ~x730 & ~x732 & ~x752 & ~x759 & ~x775 & ~x776 & ~x782;
assign c9149 =  x658 & ~x7 & ~x32 & ~x224 & ~x325 & ~x326 & ~x341 & ~x464 & ~x771;
assign c9151 =  x293 & ~x16 & ~x22 & ~x23 & ~x29 & ~x49 & ~x64 & ~x70 & ~x73 & ~x81 & ~x82 & ~x89 & ~x98 & ~x105 & ~x117 & ~x121 & ~x132 & ~x177 & ~x308 & ~x336 & ~x380 & ~x459 & ~x460 & ~x475 & ~x486 & ~x487 & ~x529 & ~x559 & ~x562 & ~x585 & ~x670 & ~x695 & ~x733 & ~x755 & ~x764;
assign c9153 =  x191;
assign c9155 =  x300 & ~x37 & ~x378 & ~x428 & ~x440 & ~x455 & ~x510 & ~x559;
assign c9157 = ~x80 & ~x81 & ~x88 & ~x119 & ~x120 & ~x141 & ~x148 & ~x167 & ~x194 & ~x228 & ~x249 & ~x306 & ~x309 & ~x321 & ~x338 & ~x377 & ~x403 & ~x425 & ~x426 & ~x430 & ~x452 & ~x456 & ~x472 & ~x562 & ~x621 & ~x696 & ~x702 & ~x770 & ~x779 & ~x780;
assign c9159 =  x348 &  x632 & ~x1 & ~x80 & ~x619 & ~x693 & ~x743 & ~x766 & ~x783;
assign c9161 =  x494 & ~x0 & ~x5 & ~x10 & ~x50 & ~x55 & ~x82 & ~x86 & ~x97 & ~x106 & ~x167 & ~x249 & ~x329 & ~x330 & ~x336 & ~x355 & ~x356 & ~x363 & ~x392 & ~x393 & ~x473 & ~x553 & ~x638 & ~x639 & ~x668 & ~x692 & ~x704 & ~x717 & ~x720 & ~x732 & ~x735 & ~x736 & ~x746 & ~x757 & ~x774;
assign c9163 =  x538;
assign c9165 = ~x42 & ~x74 & ~x137 & ~x252 & ~x320 & ~x334 & ~x340 & ~x344 & ~x345 & ~x364 & ~x369 & ~x398 & ~x421 & ~x423 & ~x448 & ~x476 & ~x560 & ~x690 & ~x704 & ~x725 & ~x765 & ~x781;
assign c9167 =  x241 &  x269 & ~x1 & ~x2 & ~x7 & ~x25 & ~x26 & ~x29 & ~x30 & ~x34 & ~x40 & ~x45 & ~x49 & ~x52 & ~x59 & ~x60 & ~x74 & ~x76 & ~x77 & ~x79 & ~x87 & ~x97 & ~x98 & ~x99 & ~x102 & ~x104 & ~x139 & ~x141 & ~x145 & ~x155 & ~x169 & ~x172 & ~x191 & ~x194 & ~x211 & ~x217 & ~x224 & ~x227 & ~x273 & ~x303 & ~x391 & ~x421 & ~x423 & ~x451 & ~x475 & ~x478 & ~x503 & ~x527 & ~x533 & ~x555 & ~x558 & ~x560 & ~x565 & ~x585 & ~x589 & ~x594 & ~x595 & ~x610 & ~x611 & ~x614 & ~x639 & ~x646 & ~x668 & ~x697 & ~x702 & ~x706 & ~x709 & ~x719 & ~x723 & ~x726 & ~x730 & ~x734 & ~x736 & ~x738 & ~x741 & ~x743 & ~x747 & ~x752 & ~x754 & ~x757 & ~x767 & ~x772 & ~x775 & ~x776 & ~x782;
assign c9169 =  x239 &  x263 &  x264 &  x265 & ~x12 & ~x21 & ~x67 & ~x101 & ~x118 & ~x252 & ~x255 & ~x335 & ~x392 & ~x451 & ~x497 & ~x588 & ~x665 & ~x667 & ~x696 & ~x698 & ~x701 & ~x716 & ~x742 & ~x743 & ~x753 & ~x763 & ~x775 & ~x776 & ~x778;
assign c9171 =  x539 & ~x204 & ~x662 & ~x688 & ~x689;
assign c9173 =  x484 &  x512 &  x626;
assign c9175 =  x176 & ~x44 & ~x116 & ~x313;
assign c9177 =  x218 & ~x410;
assign c9179 =  x572 & ~x8 & ~x23 & ~x27 & ~x38 & ~x46 & ~x55 & ~x58 & ~x79 & ~x82 & ~x84 & ~x88 & ~x105 & ~x107 & ~x109 & ~x113 & ~x115 & ~x129 & ~x134 & ~x137 & ~x140 & ~x165 & ~x166 & ~x168 & ~x176 & ~x226 & ~x280 & ~x285 & ~x312 & ~x313 & ~x340 & ~x392 & ~x419 & ~x421 & ~x474 & ~x502 & ~x505 & ~x530 & ~x531 & ~x532 & ~x614 & ~x616 & ~x618 & ~x635 & ~x639 & ~x648 & ~x649 & ~x663 & ~x664 & ~x665 & ~x668 & ~x678 & ~x680 & ~x689 & ~x691 & ~x692 & ~x696 & ~x700 & ~x711 & ~x716 & ~x731 & ~x737 & ~x750 & ~x758 & ~x766 & ~x774 & ~x775;
assign c9181 =  x527;
assign c9183 =  x566 & ~x605;
assign c9185 =  x189 & ~x383;
assign c9187 =  x430 & ~x35 & ~x55 & ~x118 & ~x136 & ~x137 & ~x163 & ~x170 & ~x171 & ~x174 & ~x303 & ~x359 & ~x368 & ~x476 & ~x501 & ~x504 & ~x534 & ~x544 & ~x558 & ~x593 & ~x610 & ~x619 & ~x700 & ~x713 & ~x716 & ~x718 & ~x719 & ~x723 & ~x771;
assign c9189 = ~x54 & ~x94 & ~x99 & ~x105 & ~x110 & ~x118 & ~x144 & ~x149 & ~x170 & ~x178 & ~x351 & ~x403 & ~x427 & ~x429 & ~x430 & ~x483 & ~x512 & ~x533 & ~x555 & ~x563 & ~x583 & ~x609 & ~x611 & ~x640 & ~x666 & ~x775 & ~x780;
assign c9191 =  x201;
assign c9193 =  x569 & ~x408 & ~x720;
assign c9195 =  x129;
assign c9197 =  x159 & ~x317;
assign c9199 = ~x12 & ~x14 & ~x23 & ~x25 & ~x26 & ~x38 & ~x42 & ~x43 & ~x44 & ~x46 & ~x50 & ~x54 & ~x58 & ~x62 & ~x65 & ~x66 & ~x70 & ~x72 & ~x73 & ~x77 & ~x82 & ~x83 & ~x99 & ~x101 & ~x109 & ~x110 & ~x117 & ~x122 & ~x125 & ~x128 & ~x131 & ~x134 & ~x137 & ~x138 & ~x139 & ~x141 & ~x150 & ~x162 & ~x164 & ~x166 & ~x170 & ~x174 & ~x180 & ~x190 & ~x191 & ~x192 & ~x193 & ~x201 & ~x225 & ~x306 & ~x308 & ~x331 & ~x333 & ~x334 & ~x359 & ~x361 & ~x364 & ~x376 & ~x378 & ~x387 & ~x406 & ~x422 & ~x447 & ~x448 & ~x449 & ~x451 & ~x473 & ~x474 & ~x479 & ~x486 & ~x487 & ~x502 & ~x516 & ~x528 & ~x542 & ~x543 & ~x553 & ~x554 & ~x555 & ~x561 & ~x566 & ~x581 & ~x584 & ~x585 & ~x594 & ~x609 & ~x612 & ~x620 & ~x625 & ~x626 & ~x637 & ~x638 & ~x639 & ~x646 & ~x653 & ~x664 & ~x667 & ~x677 & ~x682 & ~x693 & ~x699 & ~x705 & ~x708 & ~x720 & ~x722 & ~x723 & ~x724 & ~x736 & ~x749 & ~x750 & ~x756 & ~x757 & ~x759 & ~x762 & ~x771 & ~x776 & ~x779 & ~x782;
assign c9201 =  x149;
assign c9203 = ~x5 & ~x7 & ~x8 & ~x12 & ~x26 & ~x41 & ~x55 & ~x62 & ~x65 & ~x67 & ~x68 & ~x69 & ~x71 & ~x77 & ~x80 & ~x91 & ~x100 & ~x105 & ~x106 & ~x111 & ~x118 & ~x127 & ~x135 & ~x144 & ~x155 & ~x156 & ~x199 & ~x251 & ~x253 & ~x276 & ~x305 & ~x308 & ~x338 & ~x361 & ~x367 & ~x377 & ~x378 & ~x396 & ~x404 & ~x405 & ~x416 & ~x421 & ~x431 & ~x432 & ~x450 & ~x460 & ~x485 & ~x487 & ~x501 & ~x512 & ~x558 & ~x567 & ~x595 & ~x614 & ~x640 & ~x671 & ~x672 & ~x676 & ~x678 & ~x696 & ~x697 & ~x698 & ~x719 & ~x727 & ~x749 & ~x752 & ~x778;
assign c9205 =  x228;
assign c9207 = ~x0 & ~x8 & ~x16 & ~x18 & ~x24 & ~x25 & ~x26 & ~x28 & ~x33 & ~x37 & ~x40 & ~x43 & ~x44 & ~x46 & ~x48 & ~x57 & ~x59 & ~x62 & ~x66 & ~x79 & ~x89 & ~x90 & ~x93 & ~x94 & ~x96 & ~x103 & ~x112 & ~x113 & ~x116 & ~x137 & ~x138 & ~x139 & ~x145 & ~x154 & ~x155 & ~x156 & ~x167 & ~x173 & ~x183 & ~x184 & ~x193 & ~x195 & ~x198 & ~x210 & ~x212 & ~x223 & ~x239 & ~x254 & ~x266 & ~x277 & ~x278 & ~x279 & ~x305 & ~x333 & ~x337 & ~x361 & ~x365 & ~x390 & ~x392 & ~x394 & ~x395 & ~x417 & ~x445 & ~x448 & ~x478 & ~x499 & ~x509 & ~x527 & ~x529 & ~x537 & ~x555 & ~x556 & ~x557 & ~x559 & ~x563 & ~x565 & ~x583 & ~x584 & ~x589 & ~x615 & ~x617 & ~x619 & ~x620 & ~x622 & ~x639 & ~x641 & ~x644 & ~x645 & ~x667 & ~x674 & ~x675 & ~x679 & ~x693 & ~x696 & ~x705 & ~x720 & ~x722 & ~x724 & ~x725 & ~x730 & ~x731 & ~x743 & ~x747 & ~x753 & ~x760 & ~x761 & ~x762 & ~x769 & ~x776;
assign c9209 =  x433 & ~x25 & ~x35 & ~x75 & ~x92 & ~x164 & ~x217 & ~x299 & ~x326 & ~x339 & ~x354 & ~x363 & ~x423 & ~x451 & ~x475 & ~x506 & ~x565 & ~x618 & ~x691 & ~x705 & ~x711 & ~x713 & ~x718 & ~x720 & ~x735 & ~x737 & ~x743 & ~x749 & ~x760 & ~x773;
assign c9211 =  x272 &  x299 & ~x2 & ~x7 & ~x8 & ~x10 & ~x11 & ~x12 & ~x13 & ~x16 & ~x17 & ~x22 & ~x28 & ~x30 & ~x39 & ~x41 & ~x42 & ~x43 & ~x49 & ~x50 & ~x70 & ~x74 & ~x77 & ~x78 & ~x88 & ~x90 & ~x103 & ~x107 & ~x108 & ~x116 & ~x117 & ~x125 & ~x127 & ~x129 & ~x136 & ~x137 & ~x138 & ~x145 & ~x157 & ~x167 & ~x185 & ~x186 & ~x213 & ~x221 & ~x222 & ~x226 & ~x251 & ~x336 & ~x338 & ~x359 & ~x360 & ~x366 & ~x389 & ~x447 & ~x478 & ~x503 & ~x530 & ~x536 & ~x555 & ~x560 & ~x612 & ~x618 & ~x619 & ~x650 & ~x666 & ~x668 & ~x671 & ~x673 & ~x696 & ~x703 & ~x706 & ~x719 & ~x726 & ~x731 & ~x742 & ~x747 & ~x757 & ~x767 & ~x776 & ~x777 & ~x781;
assign c9213 =  x162;
assign c9215 =  x467 & ~x1 & ~x3 & ~x6 & ~x10 & ~x12 & ~x15 & ~x19 & ~x20 & ~x29 & ~x38 & ~x44 & ~x70 & ~x80 & ~x82 & ~x83 & ~x88 & ~x89 & ~x99 & ~x108 & ~x111 & ~x113 & ~x115 & ~x119 & ~x144 & ~x166 & ~x169 & ~x196 & ~x223 & ~x224 & ~x247 & ~x249 & ~x250 & ~x281 & ~x288 & ~x310 & ~x312 & ~x342 & ~x363 & ~x364 & ~x419 & ~x448 & ~x476 & ~x505 & ~x532 & ~x562 & ~x563 & ~x612 & ~x616 & ~x640 & ~x643 & ~x647 & ~x665 & ~x668 & ~x670 & ~x674 & ~x678 & ~x691 & ~x692 & ~x693 & ~x695 & ~x697 & ~x698 & ~x700 & ~x702 & ~x711 & ~x728 & ~x730 & ~x734 & ~x739 & ~x743 & ~x746 & ~x747 & ~x757 & ~x760 & ~x763 & ~x769;
assign c9217 =  x218 &  x245 & ~x24 & ~x385 & ~x386 & ~x512;
assign c9219 = ~x3 & ~x4 & ~x5 & ~x9 & ~x16 & ~x19 & ~x23 & ~x26 & ~x29 & ~x32 & ~x35 & ~x38 & ~x39 & ~x44 & ~x47 & ~x53 & ~x55 & ~x58 & ~x62 & ~x64 & ~x67 & ~x70 & ~x73 & ~x77 & ~x78 & ~x82 & ~x83 & ~x86 & ~x95 & ~x97 & ~x104 & ~x106 & ~x108 & ~x109 & ~x111 & ~x115 & ~x121 & ~x136 & ~x139 & ~x143 & ~x153 & ~x154 & ~x156 & ~x167 & ~x168 & ~x170 & ~x171 & ~x182 & ~x183 & ~x195 & ~x197 & ~x198 & ~x200 & ~x210 & ~x211 & ~x224 & ~x225 & ~x238 & ~x239 & ~x250 & ~x252 & ~x254 & ~x266 & ~x267 & ~x281 & ~x294 & ~x295 & ~x308 & ~x309 & ~x310 & ~x335 & ~x336 & ~x338 & ~x363 & ~x392 & ~x421 & ~x422 & ~x447 & ~x478 & ~x501 & ~x503 & ~x505 & ~x506 & ~x531 & ~x532 & ~x533 & ~x557 & ~x561 & ~x562 & ~x565 & ~x582 & ~x583 & ~x584 & ~x585 & ~x586 & ~x587 & ~x594 & ~x597 & ~x611 & ~x613 & ~x614 & ~x616 & ~x618 & ~x622 & ~x623 & ~x639 & ~x640 & ~x641 & ~x644 & ~x645 & ~x650 & ~x670 & ~x676 & ~x682 & ~x696 & ~x700 & ~x701 & ~x702 & ~x706 & ~x709 & ~x721 & ~x723 & ~x727 & ~x731 & ~x732 & ~x734 & ~x737 & ~x740 & ~x743 & ~x746 & ~x747 & ~x748 & ~x750 & ~x751 & ~x756 & ~x761 & ~x762 & ~x767 & ~x775 & ~x776 & ~x783;
assign c9221 = ~x24 & ~x48 & ~x72 & ~x73 & ~x86 & ~x120 & ~x122 & ~x198 & ~x280 & ~x309 & ~x321 & ~x335 & ~x347 & ~x348 & ~x360 & ~x402 & ~x443 & ~x444 & ~x456 & ~x476 & ~x483 & ~x502 & ~x535 & ~x558 & ~x588 & ~x704 & ~x728 & ~x730 & ~x734;
assign c9223 =  x498 & ~x396 & ~x769;
assign c9225 =  x240 & ~x6 & ~x16 & ~x77 & ~x141 & ~x306 & ~x322 & ~x350 & ~x368 & ~x374 & ~x399 & ~x425 & ~x528 & ~x588 & ~x730;
assign c9227 =  x500;
assign c9229 =  x434 & ~x0 & ~x7 & ~x23 & ~x25 & ~x65 & ~x82 & ~x91 & ~x92 & ~x109 & ~x111 & ~x133 & ~x141 & ~x164 & ~x192 & ~x224 & ~x254 & ~x284 & ~x344 & ~x346 & ~x347 & ~x365 & ~x367 & ~x530 & ~x642 & ~x673 & ~x697 & ~x701 & ~x704 & ~x722 & ~x741 & ~x756 & ~x772;
assign c9231 =  x159 &  x657;
assign c9233 =  x209 & ~x14 & ~x36 & ~x41 & ~x48 & ~x58 & ~x65 & ~x66 & ~x80 & ~x86 & ~x92 & ~x93 & ~x109 & ~x117 & ~x138 & ~x139 & ~x142 & ~x166 & ~x168 & ~x195 & ~x199 & ~x201 & ~x202 & ~x258 & ~x286 & ~x288 & ~x290 & ~x316 & ~x331 & ~x333 & ~x340 & ~x342 & ~x362 & ~x368 & ~x390 & ~x415 & ~x420 & ~x474 & ~x526 & ~x532 & ~x533 & ~x585 & ~x587 & ~x588 & ~x612 & ~x614 & ~x640 & ~x668 & ~x675 & ~x703 & ~x713 & ~x714 & ~x729 & ~x734 & ~x740 & ~x745 & ~x752 & ~x758 & ~x761 & ~x764 & ~x775;
assign c9235 =  x432 & ~x0 & ~x7 & ~x12 & ~x13 & ~x31 & ~x35 & ~x44 & ~x45 & ~x51 & ~x61 & ~x65 & ~x67 & ~x76 & ~x80 & ~x91 & ~x93 & ~x97 & ~x100 & ~x103 & ~x108 & ~x110 & ~x128 & ~x150 & ~x164 & ~x171 & ~x174 & ~x196 & ~x198 & ~x200 & ~x252 & ~x254 & ~x255 & ~x256 & ~x306 & ~x312 & ~x332 & ~x341 & ~x343 & ~x361 & ~x363 & ~x370 & ~x371 & ~x373 & ~x387 & ~x389 & ~x397 & ~x420 & ~x421 & ~x448 & ~x470 & ~x474 & ~x475 & ~x476 & ~x501 & ~x503 & ~x504 & ~x557 & ~x561 & ~x592 & ~x637 & ~x639 & ~x643 & ~x649 & ~x666 & ~x668 & ~x672 & ~x696 & ~x698 & ~x700 & ~x702 & ~x717 & ~x718 & ~x721 & ~x725 & ~x734 & ~x744 & ~x753 & ~x754 & ~x761 & ~x763 & ~x771 & ~x776 & ~x777 & ~x782;
assign c9237 = ~x20 & ~x26 & ~x41 & ~x42 & ~x72 & ~x74 & ~x79 & ~x82 & ~x84 & ~x96 & ~x104 & ~x108 & ~x292 & ~x310 & ~x311 & ~x318 & ~x333 & ~x334 & ~x342 & ~x344 & ~x360 & ~x369 & ~x396 & ~x450 & ~x721 & ~x722 & ~x729 & ~x742 & ~x748 & ~x749 & ~x773 & ~x776;
assign c9239 =  x214 &  x376 &  x402 & ~x12 & ~x17 & ~x36 & ~x49 & ~x73 & ~x107 & ~x138 & ~x145 & ~x277 & ~x356 & ~x369 & ~x388 & ~x418 & ~x448 & ~x535 & ~x612 & ~x743 & ~x752 & ~x756 & ~x760 & ~x767 & ~x778 & ~x780;
assign c9241 = ~x7 & ~x10 & ~x23 & ~x32 & ~x39 & ~x42 & ~x47 & ~x49 & ~x53 & ~x54 & ~x55 & ~x57 & ~x59 & ~x63 & ~x64 & ~x74 & ~x75 & ~x76 & ~x78 & ~x89 & ~x96 & ~x100 & ~x101 & ~x106 & ~x110 & ~x117 & ~x119 & ~x132 & ~x137 & ~x142 & ~x143 & ~x170 & ~x171 & ~x198 & ~x227 & ~x253 & ~x279 & ~x282 & ~x284 & ~x307 & ~x313 & ~x315 & ~x320 & ~x342 & ~x343 & ~x345 & ~x363 & ~x395 & ~x422 & ~x450 & ~x499 & ~x505 & ~x508 & ~x531 & ~x533 & ~x559 & ~x561 & ~x562 & ~x586 & ~x587 & ~x589 & ~x614 & ~x615 & ~x616 & ~x643 & ~x670 & ~x691 & ~x698 & ~x704 & ~x719 & ~x728 & ~x732 & ~x733 & ~x737 & ~x753 & ~x766 & ~x769 & ~x774 & ~x775;
assign c9243 =  x156 & ~x234 & ~x235 & ~x340 & ~x684;
assign c9245 =  x543 &  x598 &  x599 & ~x2 & ~x3 & ~x10 & ~x12 & ~x14 & ~x19 & ~x20 & ~x22 & ~x23 & ~x28 & ~x32 & ~x39 & ~x45 & ~x50 & ~x54 & ~x56 & ~x57 & ~x60 & ~x61 & ~x62 & ~x64 & ~x70 & ~x71 & ~x74 & ~x76 & ~x81 & ~x89 & ~x92 & ~x106 & ~x114 & ~x116 & ~x119 & ~x121 & ~x139 & ~x141 & ~x142 & ~x167 & ~x171 & ~x173 & ~x193 & ~x198 & ~x200 & ~x224 & ~x227 & ~x228 & ~x251 & ~x252 & ~x253 & ~x280 & ~x281 & ~x283 & ~x340 & ~x361 & ~x362 & ~x366 & ~x367 & ~x391 & ~x395 & ~x451 & ~x473 & ~x474 & ~x500 & ~x558 & ~x586 & ~x587 & ~x589 & ~x613 & ~x614 & ~x615 & ~x644 & ~x650 & ~x668 & ~x669 & ~x671 & ~x673 & ~x678 & ~x679 & ~x680 & ~x692 & ~x693 & ~x696 & ~x697 & ~x703 & ~x705 & ~x707 & ~x708 & ~x717 & ~x720 & ~x722 & ~x728 & ~x735 & ~x746 & ~x750 & ~x753 & ~x754 & ~x760 & ~x764 & ~x767;
assign c9247 =  x131;
assign c9249 = ~x0 & ~x3 & ~x14 & ~x25 & ~x38 & ~x50 & ~x56 & ~x57 & ~x58 & ~x59 & ~x62 & ~x63 & ~x77 & ~x82 & ~x83 & ~x87 & ~x114 & ~x140 & ~x141 & ~x168 & ~x169 & ~x173 & ~x176 & ~x184 & ~x185 & ~x202 & ~x222 & ~x226 & ~x232 & ~x240 & ~x251 & ~x254 & ~x283 & ~x314 & ~x323 & ~x334 & ~x338 & ~x361 & ~x388 & ~x389 & ~x390 & ~x393 & ~x417 & ~x421 & ~x449 & ~x450 & ~x474 & ~x476 & ~x498 & ~x500 & ~x505 & ~x508 & ~x526 & ~x530 & ~x557 & ~x558 & ~x559 & ~x565 & ~x567 & ~x581 & ~x593 & ~x616 & ~x618 & ~x621 & ~x651 & ~x666 & ~x669 & ~x675 & ~x693 & ~x695 & ~x698 & ~x700 & ~x702 & ~x708 & ~x727 & ~x731 & ~x743 & ~x746 & ~x749 & ~x754 & ~x759 & ~x774 & ~x776 & ~x777 & ~x780 & ~x782 & ~x783;
assign c9251 =  x597 & ~x113 & ~x251 & ~x340 & ~x354 & ~x643 & ~x702 & ~x725 & ~x752;
assign c9253 =  x463 & ~x1 & ~x3 & ~x5 & ~x13 & ~x14 & ~x16 & ~x17 & ~x19 & ~x20 & ~x21 & ~x26 & ~x27 & ~x31 & ~x33 & ~x34 & ~x36 & ~x41 & ~x42 & ~x44 & ~x47 & ~x53 & ~x54 & ~x58 & ~x61 & ~x69 & ~x72 & ~x75 & ~x78 & ~x79 & ~x80 & ~x86 & ~x88 & ~x92 & ~x101 & ~x108 & ~x110 & ~x111 & ~x112 & ~x133 & ~x136 & ~x139 & ~x140 & ~x142 & ~x144 & ~x147 & ~x167 & ~x169 & ~x183 & ~x196 & ~x199 & ~x211 & ~x222 & ~x227 & ~x252 & ~x267 & ~x279 & ~x280 & ~x284 & ~x295 & ~x306 & ~x311 & ~x335 & ~x337 & ~x361 & ~x366 & ~x367 & ~x389 & ~x390 & ~x395 & ~x418 & ~x421 & ~x423 & ~x445 & ~x450 & ~x476 & ~x480 & ~x502 & ~x503 & ~x504 & ~x509 & ~x538 & ~x560 & ~x565 & ~x584 & ~x586 & ~x587 & ~x588 & ~x589 & ~x622 & ~x643 & ~x645 & ~x647 & ~x650 & ~x651 & ~x668 & ~x671 & ~x676 & ~x694 & ~x696 & ~x706 & ~x718 & ~x720 & ~x721 & ~x725 & ~x726 & ~x727 & ~x728 & ~x730 & ~x731 & ~x732 & ~x734 & ~x736 & ~x739 & ~x741 & ~x742 & ~x750 & ~x753 & ~x754 & ~x755 & ~x763 & ~x764 & ~x766 & ~x769 & ~x770 & ~x771 & ~x775 & ~x776 & ~x777 & ~x779 & ~x783;
assign c9255 =  x473;
assign c9257 = ~x0 & ~x2 & ~x4 & ~x17 & ~x33 & ~x36 & ~x40 & ~x54 & ~x78 & ~x79 & ~x81 & ~x87 & ~x96 & ~x109 & ~x118 & ~x134 & ~x136 & ~x137 & ~x163 & ~x167 & ~x191 & ~x195 & ~x250 & ~x253 & ~x280 & ~x307 & ~x311 & ~x376 & ~x392 & ~x403 & ~x404 & ~x430 & ~x452 & ~x458 & ~x459 & ~x502 & ~x514 & ~x530 & ~x541 & ~x582 & ~x589 & ~x616 & ~x643 & ~x647 & ~x718 & ~x728 & ~x767 & ~x775 & ~x778;
assign c9259 = ~x24 & ~x51 & ~x55 & ~x57 & ~x91 & ~x101 & ~x116 & ~x194 & ~x199 & ~x222 & ~x225 & ~x302 & ~x364 & ~x375 & ~x394 & ~x402 & ~x429 & ~x447 & ~x451 & ~x458 & ~x478 & ~x484 & ~x485 & ~x486 & ~x540 & ~x591 & ~x610 & ~x613 & ~x615 & ~x616 & ~x618 & ~x701 & ~x721 & ~x728 & ~x756 & ~x780;
assign c9261 =  x472;
assign c9263 =  x660 & ~x31 & ~x34 & ~x39 & ~x67 & ~x81 & ~x90 & ~x95 & ~x107 & ~x109 & ~x112 & ~x116 & ~x150 & ~x154 & ~x181 & ~x209 & ~x309 & ~x417 & ~x421 & ~x451 & ~x477 & ~x510 & ~x539 & ~x542 & ~x557 & ~x567 & ~x583 & ~x584 & ~x600 & ~x701 & ~x721 & ~x732 & ~x745;
assign c9265 =  x99;
assign c9267 =  x175;
assign c9269 = ~x0 & ~x1 & ~x2 & ~x4 & ~x10 & ~x12 & ~x13 & ~x14 & ~x17 & ~x22 & ~x23 & ~x24 & ~x28 & ~x35 & ~x41 & ~x45 & ~x47 & ~x48 & ~x49 & ~x50 & ~x52 & ~x53 & ~x59 & ~x61 & ~x62 & ~x63 & ~x64 & ~x65 & ~x66 & ~x67 & ~x69 & ~x70 & ~x76 & ~x78 & ~x83 & ~x84 & ~x85 & ~x88 & ~x90 & ~x94 & ~x97 & ~x102 & ~x103 & ~x104 & ~x105 & ~x107 & ~x110 & ~x111 & ~x113 & ~x115 & ~x116 & ~x117 & ~x120 & ~x126 & ~x133 & ~x137 & ~x138 & ~x139 & ~x140 & ~x141 & ~x144 & ~x148 & ~x154 & ~x166 & ~x167 & ~x168 & ~x171 & ~x172 & ~x182 & ~x192 & ~x194 & ~x195 & ~x196 & ~x198 & ~x199 & ~x200 & ~x210 & ~x222 & ~x225 & ~x226 & ~x238 & ~x254 & ~x255 & ~x256 & ~x266 & ~x277 & ~x278 & ~x281 & ~x282 & ~x283 & ~x284 & ~x294 & ~x305 & ~x307 & ~x309 & ~x311 & ~x321 & ~x336 & ~x337 & ~x339 & ~x364 & ~x365 & ~x389 & ~x390 & ~x391 & ~x394 & ~x416 & ~x417 & ~x418 & ~x423 & ~x445 & ~x447 & ~x449 & ~x450 & ~x452 & ~x474 & ~x475 & ~x479 & ~x499 & ~x500 & ~x501 & ~x506 & ~x508 & ~x527 & ~x528 & ~x533 & ~x534 & ~x537 & ~x538 & ~x556 & ~x558 & ~x559 & ~x560 & ~x563 & ~x564 & ~x566 & ~x568 & ~x569 & ~x582 & ~x586 & ~x587 & ~x590 & ~x593 & ~x594 & ~x611 & ~x615 & ~x617 & ~x618 & ~x620 & ~x621 & ~x639 & ~x641 & ~x648 & ~x666 & ~x667 & ~x669 & ~x671 & ~x672 & ~x673 & ~x675 & ~x676 & ~x678 & ~x679 & ~x694 & ~x695 & ~x699 & ~x700 & ~x702 & ~x705 & ~x706 & ~x707 & ~x709 & ~x722 & ~x724 & ~x725 & ~x726 & ~x730 & ~x732 & ~x733 & ~x735 & ~x736 & ~x740 & ~x742 & ~x744 & ~x745 & ~x747 & ~x748 & ~x750 & ~x753 & ~x755 & ~x756 & ~x763 & ~x764 & ~x766 & ~x767 & ~x768 & ~x770 & ~x773 & ~x776 & ~x778 & ~x780 & ~x782 & ~x783;
assign c9271 =  x578 & ~x84 & ~x93 & ~x100 & ~x101 & ~x122 & ~x126 & ~x196 & ~x333 & ~x341 & ~x344 & ~x363 & ~x366 & ~x369 & ~x370 & ~x371 & ~x399 & ~x504 & ~x530 & ~x557 & ~x560 & ~x561 & ~x641 & ~x671 & ~x674 & ~x729 & ~x730 & ~x766 & ~x773;
assign c9273 = ~x4 & ~x8 & ~x9 & ~x12 & ~x13 & ~x14 & ~x16 & ~x17 & ~x18 & ~x19 & ~x21 & ~x22 & ~x31 & ~x32 & ~x34 & ~x35 & ~x42 & ~x49 & ~x52 & ~x54 & ~x55 & ~x56 & ~x57 & ~x60 & ~x62 & ~x65 & ~x71 & ~x73 & ~x74 & ~x75 & ~x78 & ~x79 & ~x80 & ~x81 & ~x83 & ~x87 & ~x89 & ~x91 & ~x99 & ~x100 & ~x101 & ~x105 & ~x106 & ~x107 & ~x112 & ~x113 & ~x114 & ~x115 & ~x119 & ~x136 & ~x137 & ~x139 & ~x144 & ~x153 & ~x164 & ~x165 & ~x166 & ~x168 & ~x181 & ~x193 & ~x194 & ~x197 & ~x209 & ~x224 & ~x236 & ~x237 & ~x251 & ~x255 & ~x266 & ~x276 & ~x278 & ~x279 & ~x281 & ~x283 & ~x292 & ~x304 & ~x308 & ~x309 & ~x333 & ~x337 & ~x361 & ~x362 & ~x363 & ~x365 & ~x366 & ~x392 & ~x393 & ~x417 & ~x420 & ~x422 & ~x446 & ~x450 & ~x473 & ~x476 & ~x477 & ~x499 & ~x500 & ~x501 & ~x502 & ~x503 & ~x507 & ~x530 & ~x532 & ~x534 & ~x536 & ~x555 & ~x559 & ~x561 & ~x562 & ~x563 & ~x567 & ~x586 & ~x587 & ~x588 & ~x590 & ~x595 & ~x611 & ~x615 & ~x642 & ~x646 & ~x648 & ~x652 & ~x654 & ~x668 & ~x669 & ~x676 & ~x677 & ~x678 & ~x679 & ~x680 & ~x681 & ~x698 & ~x702 & ~x704 & ~x705 & ~x707 & ~x708 & ~x709 & ~x710 & ~x724 & ~x726 & ~x727 & ~x730 & ~x736 & ~x738 & ~x739 & ~x746 & ~x749 & ~x752 & ~x754 & ~x759 & ~x763 & ~x770 & ~x771 & ~x772 & ~x773 & ~x778 & ~x779 & ~x780 & ~x783;
assign c9275 =  x264 &  x318 & ~x12 & ~x13 & ~x28 & ~x39 & ~x47 & ~x50 & ~x51 & ~x53 & ~x58 & ~x68 & ~x85 & ~x86 & ~x91 & ~x96 & ~x97 & ~x100 & ~x114 & ~x123 & ~x133 & ~x137 & ~x149 & ~x173 & ~x196 & ~x197 & ~x224 & ~x252 & ~x256 & ~x259 & ~x312 & ~x336 & ~x360 & ~x368 & ~x378 & ~x379 & ~x445 & ~x479 & ~x488 & ~x505 & ~x515 & ~x542 & ~x587 & ~x588 & ~x636 & ~x639 & ~x691 & ~x694 & ~x705 & ~x706 & ~x720 & ~x724 & ~x728 & ~x769 & ~x775;
assign c9277 =  x404 &  x486 & ~x398;
assign c9279 =  x163;
assign c9281 = ~x1 & ~x3 & ~x7 & ~x10 & ~x12 & ~x19 & ~x23 & ~x26 & ~x27 & ~x29 & ~x30 & ~x39 & ~x40 & ~x41 & ~x42 & ~x45 & ~x55 & ~x57 & ~x59 & ~x61 & ~x62 & ~x76 & ~x77 & ~x79 & ~x81 & ~x83 & ~x85 & ~x105 & ~x106 & ~x109 & ~x110 & ~x113 & ~x117 & ~x119 & ~x120 & ~x134 & ~x136 & ~x140 & ~x145 & ~x156 & ~x173 & ~x176 & ~x184 & ~x191 & ~x193 & ~x195 & ~x199 & ~x200 & ~x201 & ~x211 & ~x220 & ~x223 & ~x227 & ~x228 & ~x229 & ~x230 & ~x239 & ~x250 & ~x252 & ~x253 & ~x257 & ~x277 & ~x279 & ~x281 & ~x311 & ~x312 & ~x334 & ~x335 & ~x336 & ~x340 & ~x362 & ~x364 & ~x365 & ~x417 & ~x419 & ~x420 & ~x421 & ~x446 & ~x449 & ~x473 & ~x474 & ~x476 & ~x477 & ~x502 & ~x504 & ~x505 & ~x506 & ~x554 & ~x557 & ~x560 & ~x561 & ~x562 & ~x563 & ~x565 & ~x566 & ~x592 & ~x593 & ~x610 & ~x611 & ~x614 & ~x616 & ~x640 & ~x642 & ~x646 & ~x648 & ~x650 & ~x669 & ~x672 & ~x678 & ~x679 & ~x680 & ~x690 & ~x694 & ~x696 & ~x706 & ~x707 & ~x717 & ~x719 & ~x721 & ~x723 & ~x724 & ~x729 & ~x732 & ~x737 & ~x742 & ~x743 & ~x745 & ~x746 & ~x752 & ~x753 & ~x756 & ~x760 & ~x761 & ~x763 & ~x766 & ~x767 & ~x768 & ~x770 & ~x783;
assign c9283 =  x468 &  x469 & ~x85 & ~x285 & ~x312 & ~x313 & ~x341 & ~x368 & ~x396;
assign c9285 =  x471;
assign c9287 =  x154 & ~x108 & ~x316 & ~x324;
assign c9289 =  x256;
assign c9291 = ~x0 & ~x1 & ~x2 & ~x3 & ~x4 & ~x6 & ~x7 & ~x10 & ~x12 & ~x13 & ~x14 & ~x16 & ~x17 & ~x18 & ~x19 & ~x20 & ~x21 & ~x22 & ~x24 & ~x28 & ~x29 & ~x31 & ~x32 & ~x34 & ~x36 & ~x37 & ~x39 & ~x41 & ~x42 & ~x45 & ~x46 & ~x47 & ~x51 & ~x52 & ~x54 & ~x55 & ~x59 & ~x60 & ~x61 & ~x62 & ~x64 & ~x65 & ~x66 & ~x70 & ~x71 & ~x77 & ~x79 & ~x80 & ~x82 & ~x84 & ~x85 & ~x88 & ~x89 & ~x91 & ~x93 & ~x94 & ~x95 & ~x97 & ~x98 & ~x99 & ~x102 & ~x103 & ~x105 & ~x107 & ~x108 & ~x110 & ~x112 & ~x115 & ~x116 & ~x117 & ~x118 & ~x119 & ~x121 & ~x122 & ~x124 & ~x125 & ~x126 & ~x133 & ~x134 & ~x137 & ~x138 & ~x139 & ~x140 & ~x142 & ~x143 & ~x144 & ~x153 & ~x162 & ~x164 & ~x167 & ~x170 & ~x171 & ~x181 & ~x182 & ~x192 & ~x193 & ~x194 & ~x196 & ~x198 & ~x209 & ~x210 & ~x223 & ~x224 & ~x226 & ~x238 & ~x249 & ~x253 & ~x277 & ~x278 & ~x280 & ~x307 & ~x308 & ~x332 & ~x333 & ~x336 & ~x337 & ~x360 & ~x361 & ~x362 & ~x363 & ~x366 & ~x390 & ~x391 & ~x392 & ~x393 & ~x416 & ~x418 & ~x420 & ~x421 & ~x446 & ~x447 & ~x449 & ~x451 & ~x475 & ~x478 & ~x479 & ~x503 & ~x504 & ~x505 & ~x507 & ~x526 & ~x529 & ~x530 & ~x531 & ~x532 & ~x533 & ~x557 & ~x559 & ~x562 & ~x566 & ~x567 & ~x568 & ~x582 & ~x583 & ~x584 & ~x585 & ~x586 & ~x590 & ~x591 & ~x592 & ~x593 & ~x594 & ~x598 & ~x611 & ~x613 & ~x615 & ~x616 & ~x617 & ~x618 & ~x621 & ~x624 & ~x638 & ~x639 & ~x641 & ~x643 & ~x646 & ~x647 & ~x648 & ~x653 & ~x654 & ~x666 & ~x669 & ~x672 & ~x673 & ~x674 & ~x679 & ~x680 & ~x681 & ~x682 & ~x695 & ~x696 & ~x697 & ~x698 & ~x699 & ~x703 & ~x704 & ~x705 & ~x707 & ~x708 & ~x710 & ~x711 & ~x721 & ~x722 & ~x724 & ~x725 & ~x726 & ~x727 & ~x728 & ~x731 & ~x732 & ~x733 & ~x734 & ~x735 & ~x736 & ~x737 & ~x738 & ~x740 & ~x743 & ~x744 & ~x746 & ~x749 & ~x750 & ~x751 & ~x752 & ~x753 & ~x758 & ~x759 & ~x763 & ~x765 & ~x766 & ~x768 & ~x772 & ~x775 & ~x778 & ~x780 & ~x782 & ~x783;
assign c9293 = ~x10 & ~x28 & ~x102 & ~x143 & ~x159 & ~x171 & ~x186 & ~x213 & ~x280 & ~x282 & ~x363 & ~x366 & ~x393 & ~x639 & ~x662 & ~x663 & ~x676 & ~x689 & ~x692 & ~x713 & ~x715 & ~x716 & ~x718 & ~x719 & ~x720 & ~x731 & ~x733 & ~x746 & ~x767 & ~x783;
assign c9295 =  x238 &  x623;
assign c9297 =  x240 & ~x8 & ~x10 & ~x41 & ~x44 & ~x69 & ~x75 & ~x80 & ~x85 & ~x96 & ~x114 & ~x126 & ~x136 & ~x220 & ~x281 & ~x336 & ~x349 & ~x364 & ~x376 & ~x387 & ~x443 & ~x446 & ~x458 & ~x459 & ~x474 & ~x486 & ~x504 & ~x513 & ~x533 & ~x540 & ~x559 & ~x560 & ~x567 & ~x585 & ~x586 & ~x615 & ~x634 & ~x665 & ~x746;
assign c9299 =  x201;

endmodule