module tm( x0,x1,x2,x3,x4,x5,x6,x7,x8,x9,x10,x11,x12,x13,x14,x15,x16,x17,x18,x19,x20,x21,x22,x23,x24,x25,x26,x27,x28,x29,x30,x31,x32,x33,x34,x35,x36,x37,x38,x39,x40,x41,x42,x43,x44,x45,x46,x47,x48,x49,x50,x51,x52,x53,x54,x55,x56,x57,x58,x59,x60,x61,x62,x63,x64,x65,x66,x67,x68,x69,x70,x71,x72,x73,x74,x75,x76,x77,x78,x79,x80,x81,x82,x83,x84,x85,x86,x87,x88,x89,x90,x91,x92,x93,x94,x95,x96,x97,x98,x99,x100,x101,x102,x103,x104,x105,x106,x107,x108,x109,x110,x111,x112,x113,x114,x115,x116,x117,x118,x119,x120,x121,x122,x123,x124,x125,x126,x127,x128,x129,x130,x131,x132,x133,x134,x135,x136,x137,x138,x139,x140,x141,x142,x143,x144,x145,x146,x147,x148,x149,x150,x151,x152,x153,x154,x155,x156,x157,x158,x159,x160,x161,x162,x163,x164,x165,x166,x167,x168,x169,x170,x171,x172,x173,x174,x175,x176,x177,x178,x179,x180,x181,x182,x183,x184,x185,x186,x187,x188,x189,x190,x191,x192,x193,x194,x195,x196,x197,x198,x199,x200,x201,x202,x203,x204,x205,x206,x207,x208,x209,x210,x211,x212,x213,x214,x215,x216,x217,x218,x219,x220,x221,x222,x223,x224,x225,x226,x227,x228,x229,x230,x231,x232,x233,x234,x235,x236,x237,x238,x239,x240,x241,x242,x243,x244,x245,x246,x247,x248,x249,x250,x251,x252,x253,x254,x255,x256,x257,x258,x259,x260,x261,x262,x263,x264,x265,x266,x267,x268,x269,x270,x271,x272,x273,x274,x275,x276,x277,x278,x279,x280,x281,x282,x283,x284,x285,x286,x287,x288,x289,x290,x291,x292,x293,x294,x295,x296,x297,x298,x299,x300,x301,x302,x303,x304,x305,x306,x307,x308,x309,x310,x311,x312,x313,x314,x315,x316,x317,x318,x319,x320,x321,x322,x323,c1119,c0367,c0364,c0576,c0245,c0110,c1262,c024,c082,c0522,c0171,c033,c1362,c1380,c0270,c0170,c0357,c1269,c1288,c1415,c0555,c150,c1519,c0174,c1551,c1186,c053,c0517,c0309,c1185,c0429,c0135,c1478,c059,c017,c122,c177,c0331,c0472,c0286,c1175,c1483,c1333,c0375,c1254,c1503,c1530,c0141,c0218,c0302,c0189,c1147,c083,c0225,c0253,c1253,c1369,c0548,c0124,c0579,c1258,c1316,c181,c041,c1531,c1237,c1304,c1444,c1202,c1492,c145,c1421,c0336,c0116,c0500,c0459,c1354,c015,c16,c1217,c1430,c036,c034,c0285,c0105,c167,c1145,c1522,c1475,c1401,c1577,c0129,c0453,c1130,c0136,c1146,c0502,c0437,c1441,c1571,c0268,c0172,c1236,c1222,c0339,c1457,c116,c09,c089,c0516,c0133,c0251,c0407,c0585,c0209,c1218,c0413,c1498,c1140,c1112,c114,c0187,c049,c1157,c0523,c1301,c1411,c1451,c0321,c1550,c039,c0456,c08,c1377,c1311,c120,c1173,c1489,c026,c1124,c1233,c0195,c0373,c1244,c1460,c0448,c1267,c043,c1342,c1201,c1447,c0589,c0599,c173,c0197,c1139,c154,c1248,c0164,c0263,c1108,c0181,c1540,c1213,c0127,c1151,c0451,c1331,c0363,c1115,c0418,c04,c1232,c1306,c0568,c0536,c099,c0301,c0157,c149,c1183,c0120,c175,c0125,c1129,c1259,c1315,c0445,c1382,c0307,c1454,c1558,c0319,c0360,c0385,c0206,c0355,c0239,c1449,c174,c080,c023,c0554,c0395,c1167,c1160,c0188,c016,c0406,c0203,c0365,c10,c1466,c1590,c1163,c1501,c1404,c0320,c0490,c0542,c0119,c1172,c1400,c0370,c1107,c0228,c0257,c1545,c1357,c18,c0540,c1325,c0326,c1599,c0570,c169,c1219,c1341,c0444,c0290,c0313,c1413,c1491,c1588,c1543,c1414,c0574,c0178,c1479,c0508,c1536,c0100,c0481,c0550,c1136,c0298,c0381,c1358,c1456,c1572,c1121,c1347,c0467,c144,c075,c151,c0167,c1264,c021,c0386,c1225,c0246,c0211,c192,c0292,c0122,c0549,c1106,c1320,c1505,c0306,c0108,c1509,c0162,c186,c1526,c1191,c0510,c191,c1435,c1585,c0297,c0371,c0495,c0432,c0260,c1582,c1469,c1474,c1595,c110,c061,c0295,c0252,c1100,c182,c143,c1229,c00,c040,c0543,c1434,c0457,c1378,c0323,c0196,c160,c1274,c0224,c1228,c1396,c0345,c1127,c1207,c1339,c1312,c1143,c0349,c1329,c1493,c1559,c1512,c132,c0494,c1391,c1496,c1534,c0256,c176,c1374,c090,c1334,c0521,c1544,c1486,c1256,c165,c0352,c0596,c1179,c0236,c136,c030,c1481,c0440,c0318,c0397,c1587,c0426,c0208,c0534,c1349,c0222,c0462,c0411,c071,c1162,c0186,c0595,c1508,c1363,c0308,c1480,c032,c171,c0466,c1497,c1570,c078,c0243,c1517,c0294,c0498,c0571,c1223,c1557,c085,c1181,c1532,c1116,c0553,c0535,c194,c0584,c1278,c0427,c1174,c0344,c0422,c0564,c1390,c1323,c0315,c076,c0160,c0410,c1405,c1542,c0400,c1277,c0376,c1446,c0131,c1573,c0281,c1275,c0346,c1148,c1307,c068,c0289,c1261,c1149,c1279,c1273,c1134,c1182,c195,c062,c0291,c1464,c1507,c196,c1500,c0166,c1180,c1578,c1389,c1513,c0458,c1346,c0204,c1352,c155,c1548,c1376,c1224,c0202,c0470,c0279,c0305,c1592,c0223,c0322,c1247,c0399,c0401,c1554,c19,c074,c1563,c0396,c152,c1165,c0531,c0175,c1520,c0539,c1345,c1424,c1516,c11,c0591,c1206,c1271,c127,c1196,c193,c1159,c0350,c1427,c096,c0450,c0198,c0551,c1423,c0541,c079,c1227,c0177,c0303,c0325,c1298,c1221,c0532,c1490,c0390,c0137,c0168,c1178,c1539,c12,c140,c0377,c0192,c0237,c0485,c0509,c1210,c0342,c058,c06,c0561,c1338,c0388,c095,c0484,c0329,c0361,c0241,c1212,c1443,c0158,c0161,c0391,c1327,c0526,c0275,c0507,c0402,c1366,c0389,c1399,c1524,c1132,c1569,c0491,c1128,c092,c1120,c1281,c0496,c047,c0358,c1117,c1194,c0238,c0151,c0431,c0276,c088,c1296,c112,c1310,c1420,c1515,c1368,c0577,c0580,c1523,c0111,c1152,c087,c1158,c0578,c1321,c1251,c1371,c1238,c011,c057,c129,c1453,c1239,c1195,c0269,c1156,c1459,c1302,c0559,c0583,c01,c1260,c0128,c0199,c1169,c184,c0497,c0152,c0335,c1437,c1439,c1408,c0538,c0235,c159,c0274,c156,c162,c1266,c1205,c1249,c1211,c0465,c1485,c0146,c1407,c0156,c0537,c124,c073,c1370,c1596,c1294,c1289,c0392,c1387,c0316,c0101,c0525,c0492,c0159,c1436,c137,c1226,c0452,c0562,c0259,c1470,c146,c1549,c025,c1560,c0103,c0219,c142,c178,c1409,c1445,c199,c0288,c1504,c1553,c1214,c1208,c1154,c0374,c0176,c0366,c1330,c0304,c158,c180,c197,c1137,c1197,c0117,c1383,c0519,c1252,c0415,c031,c1384,c1353,c0480,c1133,c1309,c1326,c0372,c0277,c0436,c0511,c0566,c0588,c0227,c1565,c1395,c0130,c0378,c0271,c1332,c0347,c1461,c1537,c1473,c0150,c0126,c0382,c1209,c045,c0191,c0293,c0340,c1308,c0132,c0441,c1581,c0478,c0107,c1412,c1193,c0205,c1280,c0143,c0311,c0487,c1388,c0231,c1283,c027,c1385,c0499,c1416,c1463,c1255,c0512,c0518,c0102,c0545,c0479,c163,c0461,c0575,c1476,c0240,c1367,c0327,c0513,c0483,c1243,c010,c0248,c0501,c1580,c051,c17,c0332,c054,c0182,c0183,c0351,c1350,c1552,c1402,c0121,c118,c0393,c056,c1290,c1458,c0149,c0317,c0387,c0438,c0212,c1240,c1518,c1365,c164,c1155,c0560,c0547,c0190,c0338,c1564,c119,c1297,c0282,c0454,c060,c0563,c0384,c1286,c187,c0598,c1114,c1591,c1340,c1336,c1131,c1246,c1272,c1419,c130,c1198,c1538,c0463,c02,c0250,c0412,c0213,c1142,c1438,c1440,c0486,c0417,c1230,c1190,c135,c1429,c190,c0520,c1200,c0439,c0420,c1356,c1494,c1176,c0200,c1514,c018,c1562,c0469,c052,c1101,c1450,c0104,c046,c086,c0179,c0379,c1527,c1584,c1428,c1344,c1245,c1511,c042,c069,c1343,c0194,c1287,c1295,c0214,c1487,c064,c05,c0324,c0592,c0201,c198,c1468,c0398,c0220,c0524,c1521,c0383,c1216,c022,c0138,c0359,c0428,c0300,c1372,c0255,c189,c0266,c0247,c1510,c157,c1586,c0460,c14,c0242,c1150,c1184,c1337,c1319,c077,c1547,c13,c0442,c0414,c0165,c0114,c126,c0249,c0433,c029,c0435,c148,c1561,c128,c1103,c0416,c15,c028,c1533,c1102,c0506,c1471,c0408,c1242,c1386,c0343,c170,c0264,c0155,c1276,c093,c1525,c0528,c1110,c1318,c1528,c0299,c117,c1433,c0226,c1314,c1364,c0505,c0262,c1220,c1392,c0185,c1125,c0362,c1231,c1442,c0173,c0341,c0482,c0233,c1348,c1235,c037,c1135,c1317,c1541,c0380,c0404,c0546,c0567,c0169,c1282,c1452,c0443,c121,c1360,c161,c0283,c1546,c1141,c0493,c038,c0594,c0409,c0284,c067,c0145,c168,c0215,c1418,c1355,c1373,c1597,c1576,c133,c1484,c1455,c0232,c0229,c0134,c0477,c188,c0514,c055,c050,c013,c0423,c1432,c1482,c1189,c1361,c1324,c1393,c1292,c0348,c0476,c1203,c0515,c0421,c0434,c1328,c0504,c0184,c1506,c125,c172,c1535,c153,c0582,c0312,c0527,c1187,c0586,c1168,c183,c1574,c138,c1556,c0244,c019,c1126,c0328,c1394,c139,c0280,c1566,c0314,c0569,c0272,c0261,c0217,c1417,c0587,c0153,c0430,c0207,c1123,c0147,c1403,c0337,c07,c0265,c070,c1177,c094,c091,c0113,c1166,c1313,c1579,c072,c1598,c0109,c0258,c1583,c1322,c0180,c0356,c0488,c1170,c0163,c1488,c0419,c0193,c1144,c1299,c1351,c1192,c0449,c1268,c1397,c0572,c0230,c1467,c1118,c0597,c048,c1188,c0446,c1594,c0533,c1161,c098,c0573,c1381,c0334,c0210,c0254,c1379,c0425,c1293,c147,c179,c1215,c044,c1426,c1270,c1359,c014,c1431,c1265,c065,c0140,c166,c0593,c1502,c1472,c1122,c1263,c1241,c1465,c1567,c084,c0115,c1234,c1422,c0148,c0455,c1398,c185,c1555,c1593,c1199,c0544,c063,c0474,c0330,c123,c1109,c1171,c0556,c0581,c1425,c035,c1568,c0473,c1499,c1529,c0475,c0565,c1575,c1300,c131,c1495,c1305,c0530,c0468,c0552,c0369,c0278,c0216,c081,c134,c1285,c111,c0558,c1250,c0106,c0296,c0112,c012,c0234,c0424,c03,c0123,c0267,c0273,c020,c0403,c0405,c0142,c0489,c1138,c0503,c1164,c1375,c097,c0144,c0333,c0354,c0529,c1462,c0139,c0310,c1335,c1204,c0368,c1589,c0353,c1113,c1406,c0471,c1257,c1448,c0154,c0394,c1104,c0447,c0557,c0287,c1284,c1410,c1303,c0118,c1105,c1477,c1291,c141,c0590,c0221,c1153,c066,c113,c0464,c1111,c115 );

input x0;
input x1;
input x2;
input x3;
input x4;
input x5;
input x6;
input x7;
input x8;
input x9;
input x10;
input x11;
input x12;
input x13;
input x14;
input x15;
input x16;
input x17;
input x18;
input x19;
input x20;
input x21;
input x22;
input x23;
input x24;
input x25;
input x26;
input x27;
input x28;
input x29;
input x30;
input x31;
input x32;
input x33;
input x34;
input x35;
input x36;
input x37;
input x38;
input x39;
input x40;
input x41;
input x42;
input x43;
input x44;
input x45;
input x46;
input x47;
input x48;
input x49;
input x50;
input x51;
input x52;
input x53;
input x54;
input x55;
input x56;
input x57;
input x58;
input x59;
input x60;
input x61;
input x62;
input x63;
input x64;
input x65;
input x66;
input x67;
input x68;
input x69;
input x70;
input x71;
input x72;
input x73;
input x74;
input x75;
input x76;
input x77;
input x78;
input x79;
input x80;
input x81;
input x82;
input x83;
input x84;
input x85;
input x86;
input x87;
input x88;
input x89;
input x90;
input x91;
input x92;
input x93;
input x94;
input x95;
input x96;
input x97;
input x98;
input x99;
input x100;
input x101;
input x102;
input x103;
input x104;
input x105;
input x106;
input x107;
input x108;
input x109;
input x110;
input x111;
input x112;
input x113;
input x114;
input x115;
input x116;
input x117;
input x118;
input x119;
input x120;
input x121;
input x122;
input x123;
input x124;
input x125;
input x126;
input x127;
input x128;
input x129;
input x130;
input x131;
input x132;
input x133;
input x134;
input x135;
input x136;
input x137;
input x138;
input x139;
input x140;
input x141;
input x142;
input x143;
input x144;
input x145;
input x146;
input x147;
input x148;
input x149;
input x150;
input x151;
input x152;
input x153;
input x154;
input x155;
input x156;
input x157;
input x158;
input x159;
input x160;
input x161;
input x162;
input x163;
input x164;
input x165;
input x166;
input x167;
input x168;
input x169;
input x170;
input x171;
input x172;
input x173;
input x174;
input x175;
input x176;
input x177;
input x178;
input x179;
input x180;
input x181;
input x182;
input x183;
input x184;
input x185;
input x186;
input x187;
input x188;
input x189;
input x190;
input x191;
input x192;
input x193;
input x194;
input x195;
input x196;
input x197;
input x198;
input x199;
input x200;
input x201;
input x202;
input x203;
input x204;
input x205;
input x206;
input x207;
input x208;
input x209;
input x210;
input x211;
input x212;
input x213;
input x214;
input x215;
input x216;
input x217;
input x218;
input x219;
input x220;
input x221;
input x222;
input x223;
input x224;
input x225;
input x226;
input x227;
input x228;
input x229;
input x230;
input x231;
input x232;
input x233;
input x234;
input x235;
input x236;
input x237;
input x238;
input x239;
input x240;
input x241;
input x242;
input x243;
input x244;
input x245;
input x246;
input x247;
input x248;
input x249;
input x250;
input x251;
input x252;
input x253;
input x254;
input x255;
input x256;
input x257;
input x258;
input x259;
input x260;
input x261;
input x262;
input x263;
input x264;
input x265;
input x266;
input x267;
input x268;
input x269;
input x270;
input x271;
input x272;
input x273;
input x274;
input x275;
input x276;
input x277;
input x278;
input x279;
input x280;
input x281;
input x282;
input x283;
input x284;
input x285;
input x286;
input x287;
input x288;
input x289;
input x290;
input x291;
input x292;
input x293;
input x294;
input x295;
input x296;
input x297;
input x298;
input x299;
input x300;
input x301;
input x302;
input x303;
input x304;
input x305;
input x306;
input x307;
input x308;
input x309;
input x310;
input x311;
input x312;
input x313;
input x314;
input x315;
input x316;
input x317;
input x318;
input x319;
input x320;
input x321;
input x322;
input x323;
output c1119;
output c0367;
output c0364;
output c0576;
output c0245;
output c0110;
output c1262;
output c024;
output c082;
output c0522;
output c0171;
output c033;
output c1362;
output c1380;
output c0270;
output c0170;
output c0357;
output c1269;
output c1288;
output c1415;
output c0555;
output c150;
output c1519;
output c0174;
output c1551;
output c1186;
output c053;
output c0517;
output c0309;
output c1185;
output c0429;
output c0135;
output c1478;
output c059;
output c017;
output c122;
output c177;
output c0331;
output c0472;
output c0286;
output c1175;
output c1483;
output c1333;
output c0375;
output c1254;
output c1503;
output c1530;
output c0141;
output c0218;
output c0302;
output c0189;
output c1147;
output c083;
output c0225;
output c0253;
output c1253;
output c1369;
output c0548;
output c0124;
output c0579;
output c1258;
output c1316;
output c181;
output c041;
output c1531;
output c1237;
output c1304;
output c1444;
output c1202;
output c1492;
output c145;
output c1421;
output c0336;
output c0116;
output c0500;
output c0459;
output c1354;
output c015;
output c16;
output c1217;
output c1430;
output c036;
output c034;
output c0285;
output c0105;
output c167;
output c1145;
output c1522;
output c1475;
output c1401;
output c1577;
output c0129;
output c0453;
output c1130;
output c0136;
output c1146;
output c0502;
output c0437;
output c1441;
output c1571;
output c0268;
output c0172;
output c1236;
output c1222;
output c0339;
output c1457;
output c116;
output c09;
output c089;
output c0516;
output c0133;
output c0251;
output c0407;
output c0585;
output c0209;
output c1218;
output c0413;
output c1498;
output c1140;
output c1112;
output c114;
output c0187;
output c049;
output c1157;
output c0523;
output c1301;
output c1411;
output c1451;
output c0321;
output c1550;
output c039;
output c0456;
output c08;
output c1377;
output c1311;
output c120;
output c1173;
output c1489;
output c026;
output c1124;
output c1233;
output c0195;
output c0373;
output c1244;
output c1460;
output c0448;
output c1267;
output c043;
output c1342;
output c1201;
output c1447;
output c0589;
output c0599;
output c173;
output c0197;
output c1139;
output c154;
output c1248;
output c0164;
output c0263;
output c1108;
output c0181;
output c1540;
output c1213;
output c0127;
output c1151;
output c0451;
output c1331;
output c0363;
output c1115;
output c0418;
output c04;
output c1232;
output c1306;
output c0568;
output c0536;
output c099;
output c0301;
output c0157;
output c149;
output c1183;
output c0120;
output c175;
output c0125;
output c1129;
output c1259;
output c1315;
output c0445;
output c1382;
output c0307;
output c1454;
output c1558;
output c0319;
output c0360;
output c0385;
output c0206;
output c0355;
output c0239;
output c1449;
output c174;
output c080;
output c023;
output c0554;
output c0395;
output c1167;
output c1160;
output c0188;
output c016;
output c0406;
output c0203;
output c0365;
output c10;
output c1466;
output c1590;
output c1163;
output c1501;
output c1404;
output c0320;
output c0490;
output c0542;
output c0119;
output c1172;
output c1400;
output c0370;
output c1107;
output c0228;
output c0257;
output c1545;
output c1357;
output c18;
output c0540;
output c1325;
output c0326;
output c1599;
output c0570;
output c169;
output c1219;
output c1341;
output c0444;
output c0290;
output c0313;
output c1413;
output c1491;
output c1588;
output c1543;
output c1414;
output c0574;
output c0178;
output c1479;
output c0508;
output c1536;
output c0100;
output c0481;
output c0550;
output c1136;
output c0298;
output c0381;
output c1358;
output c1456;
output c1572;
output c1121;
output c1347;
output c0467;
output c144;
output c075;
output c151;
output c0167;
output c1264;
output c021;
output c0386;
output c1225;
output c0246;
output c0211;
output c192;
output c0292;
output c0122;
output c0549;
output c1106;
output c1320;
output c1505;
output c0306;
output c0108;
output c1509;
output c0162;
output c186;
output c1526;
output c1191;
output c0510;
output c191;
output c1435;
output c1585;
output c0297;
output c0371;
output c0495;
output c0432;
output c0260;
output c1582;
output c1469;
output c1474;
output c1595;
output c110;
output c061;
output c0295;
output c0252;
output c1100;
output c182;
output c143;
output c1229;
output c00;
output c040;
output c0543;
output c1434;
output c0457;
output c1378;
output c0323;
output c0196;
output c160;
output c1274;
output c0224;
output c1228;
output c1396;
output c0345;
output c1127;
output c1207;
output c1339;
output c1312;
output c1143;
output c0349;
output c1329;
output c1493;
output c1559;
output c1512;
output c132;
output c0494;
output c1391;
output c1496;
output c1534;
output c0256;
output c176;
output c1374;
output c090;
output c1334;
output c0521;
output c1544;
output c1486;
output c1256;
output c165;
output c0352;
output c0596;
output c1179;
output c0236;
output c136;
output c030;
output c1481;
output c0440;
output c0318;
output c0397;
output c1587;
output c0426;
output c0208;
output c0534;
output c1349;
output c0222;
output c0462;
output c0411;
output c071;
output c1162;
output c0186;
output c0595;
output c1508;
output c1363;
output c0308;
output c1480;
output c032;
output c171;
output c0466;
output c1497;
output c1570;
output c078;
output c0243;
output c1517;
output c0294;
output c0498;
output c0571;
output c1223;
output c1557;
output c085;
output c1181;
output c1532;
output c1116;
output c0553;
output c0535;
output c194;
output c0584;
output c1278;
output c0427;
output c1174;
output c0344;
output c0422;
output c0564;
output c1390;
output c1323;
output c0315;
output c076;
output c0160;
output c0410;
output c1405;
output c1542;
output c0400;
output c1277;
output c0376;
output c1446;
output c0131;
output c1573;
output c0281;
output c1275;
output c0346;
output c1148;
output c1307;
output c068;
output c0289;
output c1261;
output c1149;
output c1279;
output c1273;
output c1134;
output c1182;
output c195;
output c062;
output c0291;
output c1464;
output c1507;
output c196;
output c1500;
output c0166;
output c1180;
output c1578;
output c1389;
output c1513;
output c0458;
output c1346;
output c0204;
output c1352;
output c155;
output c1548;
output c1376;
output c1224;
output c0202;
output c0470;
output c0279;
output c0305;
output c1592;
output c0223;
output c0322;
output c1247;
output c0399;
output c0401;
output c1554;
output c19;
output c074;
output c1563;
output c0396;
output c152;
output c1165;
output c0531;
output c0175;
output c1520;
output c0539;
output c1345;
output c1424;
output c1516;
output c11;
output c0591;
output c1206;
output c1271;
output c127;
output c1196;
output c193;
output c1159;
output c0350;
output c1427;
output c096;
output c0450;
output c0198;
output c0551;
output c1423;
output c0541;
output c079;
output c1227;
output c0177;
output c0303;
output c0325;
output c1298;
output c1221;
output c0532;
output c1490;
output c0390;
output c0137;
output c0168;
output c1178;
output c1539;
output c12;
output c140;
output c0377;
output c0192;
output c0237;
output c0485;
output c0509;
output c1210;
output c0342;
output c058;
output c06;
output c0561;
output c1338;
output c0388;
output c095;
output c0484;
output c0329;
output c0361;
output c0241;
output c1212;
output c1443;
output c0158;
output c0161;
output c0391;
output c1327;
output c0526;
output c0275;
output c0507;
output c0402;
output c1366;
output c0389;
output c1399;
output c1524;
output c1132;
output c1569;
output c0491;
output c1128;
output c092;
output c1120;
output c1281;
output c0496;
output c047;
output c0358;
output c1117;
output c1194;
output c0238;
output c0151;
output c0431;
output c0276;
output c088;
output c1296;
output c112;
output c1310;
output c1420;
output c1515;
output c1368;
output c0577;
output c0580;
output c1523;
output c0111;
output c1152;
output c087;
output c1158;
output c0578;
output c1321;
output c1251;
output c1371;
output c1238;
output c011;
output c057;
output c129;
output c1453;
output c1239;
output c1195;
output c0269;
output c1156;
output c1459;
output c1302;
output c0559;
output c0583;
output c01;
output c1260;
output c0128;
output c0199;
output c1169;
output c184;
output c0497;
output c0152;
output c0335;
output c1437;
output c1439;
output c1408;
output c0538;
output c0235;
output c159;
output c0274;
output c156;
output c162;
output c1266;
output c1205;
output c1249;
output c1211;
output c0465;
output c1485;
output c0146;
output c1407;
output c0156;
output c0537;
output c124;
output c073;
output c1370;
output c1596;
output c1294;
output c1289;
output c0392;
output c1387;
output c0316;
output c0101;
output c0525;
output c0492;
output c0159;
output c1436;
output c137;
output c1226;
output c0452;
output c0562;
output c0259;
output c1470;
output c146;
output c1549;
output c025;
output c1560;
output c0103;
output c0219;
output c142;
output c178;
output c1409;
output c1445;
output c199;
output c0288;
output c1504;
output c1553;
output c1214;
output c1208;
output c1154;
output c0374;
output c0176;
output c0366;
output c1330;
output c0304;
output c158;
output c180;
output c197;
output c1137;
output c1197;
output c0117;
output c1383;
output c0519;
output c1252;
output c0415;
output c031;
output c1384;
output c1353;
output c0480;
output c1133;
output c1309;
output c1326;
output c0372;
output c0277;
output c0436;
output c0511;
output c0566;
output c0588;
output c0227;
output c1565;
output c1395;
output c0130;
output c0378;
output c0271;
output c1332;
output c0347;
output c1461;
output c1537;
output c1473;
output c0150;
output c0126;
output c0382;
output c1209;
output c045;
output c0191;
output c0293;
output c0340;
output c1308;
output c0132;
output c0441;
output c1581;
output c0478;
output c0107;
output c1412;
output c1193;
output c0205;
output c1280;
output c0143;
output c0311;
output c0487;
output c1388;
output c0231;
output c1283;
output c027;
output c1385;
output c0499;
output c1416;
output c1463;
output c1255;
output c0512;
output c0518;
output c0102;
output c0545;
output c0479;
output c163;
output c0461;
output c0575;
output c1476;
output c0240;
output c1367;
output c0327;
output c0513;
output c0483;
output c1243;
output c010;
output c0248;
output c0501;
output c1580;
output c051;
output c17;
output c0332;
output c054;
output c0182;
output c0183;
output c0351;
output c1350;
output c1552;
output c1402;
output c0121;
output c118;
output c0393;
output c056;
output c1290;
output c1458;
output c0149;
output c0317;
output c0387;
output c0438;
output c0212;
output c1240;
output c1518;
output c1365;
output c164;
output c1155;
output c0560;
output c0547;
output c0190;
output c0338;
output c1564;
output c119;
output c1297;
output c0282;
output c0454;
output c060;
output c0563;
output c0384;
output c1286;
output c187;
output c0598;
output c1114;
output c1591;
output c1340;
output c1336;
output c1131;
output c1246;
output c1272;
output c1419;
output c130;
output c1198;
output c1538;
output c0463;
output c02;
output c0250;
output c0412;
output c0213;
output c1142;
output c1438;
output c1440;
output c0486;
output c0417;
output c1230;
output c1190;
output c135;
output c1429;
output c190;
output c0520;
output c1200;
output c0439;
output c0420;
output c1356;
output c1494;
output c1176;
output c0200;
output c1514;
output c018;
output c1562;
output c0469;
output c052;
output c1101;
output c1450;
output c0104;
output c046;
output c086;
output c0179;
output c0379;
output c1527;
output c1584;
output c1428;
output c1344;
output c1245;
output c1511;
output c042;
output c069;
output c1343;
output c0194;
output c1287;
output c1295;
output c0214;
output c1487;
output c064;
output c05;
output c0324;
output c0592;
output c0201;
output c198;
output c1468;
output c0398;
output c0220;
output c0524;
output c1521;
output c0383;
output c1216;
output c022;
output c0138;
output c0359;
output c0428;
output c0300;
output c1372;
output c0255;
output c189;
output c0266;
output c0247;
output c1510;
output c157;
output c1586;
output c0460;
output c14;
output c0242;
output c1150;
output c1184;
output c1337;
output c1319;
output c077;
output c1547;
output c13;
output c0442;
output c0414;
output c0165;
output c0114;
output c126;
output c0249;
output c0433;
output c029;
output c0435;
output c148;
output c1561;
output c128;
output c1103;
output c0416;
output c15;
output c028;
output c1533;
output c1102;
output c0506;
output c1471;
output c0408;
output c1242;
output c1386;
output c0343;
output c170;
output c0264;
output c0155;
output c1276;
output c093;
output c1525;
output c0528;
output c1110;
output c1318;
output c1528;
output c0299;
output c117;
output c1433;
output c0226;
output c1314;
output c1364;
output c0505;
output c0262;
output c1220;
output c1392;
output c0185;
output c1125;
output c0362;
output c1231;
output c1442;
output c0173;
output c0341;
output c0482;
output c0233;
output c1348;
output c1235;
output c037;
output c1135;
output c1317;
output c1541;
output c0380;
output c0404;
output c0546;
output c0567;
output c0169;
output c1282;
output c1452;
output c0443;
output c121;
output c1360;
output c161;
output c0283;
output c1546;
output c1141;
output c0493;
output c038;
output c0594;
output c0409;
output c0284;
output c067;
output c0145;
output c168;
output c0215;
output c1418;
output c1355;
output c1373;
output c1597;
output c1576;
output c133;
output c1484;
output c1455;
output c0232;
output c0229;
output c0134;
output c0477;
output c188;
output c0514;
output c055;
output c050;
output c013;
output c0423;
output c1432;
output c1482;
output c1189;
output c1361;
output c1324;
output c1393;
output c1292;
output c0348;
output c0476;
output c1203;
output c0515;
output c0421;
output c0434;
output c1328;
output c0504;
output c0184;
output c1506;
output c125;
output c172;
output c1535;
output c153;
output c0582;
output c0312;
output c0527;
output c1187;
output c0586;
output c1168;
output c183;
output c1574;
output c138;
output c1556;
output c0244;
output c019;
output c1126;
output c0328;
output c1394;
output c139;
output c0280;
output c1566;
output c0314;
output c0569;
output c0272;
output c0261;
output c0217;
output c1417;
output c0587;
output c0153;
output c0430;
output c0207;
output c1123;
output c0147;
output c1403;
output c0337;
output c07;
output c0265;
output c070;
output c1177;
output c094;
output c091;
output c0113;
output c1166;
output c1313;
output c1579;
output c072;
output c1598;
output c0109;
output c0258;
output c1583;
output c1322;
output c0180;
output c0356;
output c0488;
output c1170;
output c0163;
output c1488;
output c0419;
output c0193;
output c1144;
output c1299;
output c1351;
output c1192;
output c0449;
output c1268;
output c1397;
output c0572;
output c0230;
output c1467;
output c1118;
output c0597;
output c048;
output c1188;
output c0446;
output c1594;
output c0533;
output c1161;
output c098;
output c0573;
output c1381;
output c0334;
output c0210;
output c0254;
output c1379;
output c0425;
output c1293;
output c147;
output c179;
output c1215;
output c044;
output c1426;
output c1270;
output c1359;
output c014;
output c1431;
output c1265;
output c065;
output c0140;
output c166;
output c0593;
output c1502;
output c1472;
output c1122;
output c1263;
output c1241;
output c1465;
output c1567;
output c084;
output c0115;
output c1234;
output c1422;
output c0148;
output c0455;
output c1398;
output c185;
output c1555;
output c1593;
output c1199;
output c0544;
output c063;
output c0474;
output c0330;
output c123;
output c1109;
output c1171;
output c0556;
output c0581;
output c1425;
output c035;
output c1568;
output c0473;
output c1499;
output c1529;
output c0475;
output c0565;
output c1575;
output c1300;
output c131;
output c1495;
output c1305;
output c0530;
output c0468;
output c0552;
output c0369;
output c0278;
output c0216;
output c081;
output c134;
output c1285;
output c111;
output c0558;
output c1250;
output c0106;
output c0296;
output c0112;
output c012;
output c0234;
output c0424;
output c03;
output c0123;
output c0267;
output c0273;
output c020;
output c0403;
output c0405;
output c0142;
output c0489;
output c1138;
output c0503;
output c1164;
output c1375;
output c097;
output c0144;
output c0333;
output c0354;
output c0529;
output c1462;
output c0139;
output c0310;
output c1335;
output c1204;
output c0368;
output c1589;
output c0353;
output c1113;
output c1406;
output c0471;
output c1257;
output c1448;
output c0154;
output c0394;
output c1104;
output c0447;
output c0557;
output c0287;
output c1284;
output c1410;
output c1303;
output c0118;
output c1105;
output c1477;
output c1291;
output c141;
output c0590;
output c0221;
output c1153;
output c066;
output c113;
output c0464;
output c1111;
output c115;

assign c00 =  x40 &  x290 & ~x145;
assign c02 = ~x157 & ~x160 & ~x287 & ~x309 & ~x321;
assign c04 =  x107 & ~x71 & ~x257 & ~x278;
assign c06 =  x131 &  x294 &  x310 &  x321;
assign c08 =  x206 &  x287 & ~x2 & ~x309;
assign c010 =  x51 &  x276 &  x308 & ~x217;
assign c012 =  x20 &  x213 & ~x163 & ~x264;
assign c014 =  x6 &  x58 &  x193 &  x202 & ~x318;
assign c016 =  x270 & ~x33 & ~x106 & ~x134;
assign c018 =  x203 &  x226 & ~x102 & ~x197;
assign c020 =  x24 & ~x84 & ~x138 & ~x174 & ~x270;
assign c022 =  x103 &  x105 & ~x21;
assign c024 =  x268 &  x288 &  x294 & ~x115;
assign c026 =  x15 &  x47 &  x74 &  x249 & ~x320;
assign c028 =  x49 &  x132 &  x158;
assign c030 =  x235 &  x258 & ~x32 & ~x157 & ~x319;
assign c032 =  x97 &  x123 &  x262 &  x285 & ~x21 & ~x111;
assign c034 =  x303 & ~x291 & ~x318 & ~x322;
assign c036 =  x16 & ~x32 & ~x195;
assign c038 =  x93 &  x187 & ~x100 & ~x105;
assign c040 =  x96 &  x193 & ~x264;
assign c042 =  x272 & ~x127 & ~x144 & ~x275;
assign c044 =  x60 &  x96 &  x283 & ~x107;
assign c046 =  x103 &  x132 &  x133 &  x312 &  x323;
assign c048 =  x24 &  x56 & ~x189 & ~x244;
assign c050 =  x16 &  x25 &  x97 & ~x289;
assign c052 =  x209 &  x268 &  x281 & ~x149 & ~x291;
assign c054 =  x101 &  x205 & ~x282;
assign c056 = ~x83 & ~x191 & ~x197 & ~x224;
assign c058 = ~x9 & ~x14 & ~x96 & ~x202 & ~x294;
assign c060 =  x14 &  x71 &  x96 &  x123 &  x155;
assign c062 =  x111 &  x143 & ~x154 & ~x159;
assign c064 =  x49 &  x90 &  x105 & ~x140;
assign c066 =  x104 &  x275 & ~x103;
assign c068 =  x38 & ~x100 & ~x291;
assign c070 =  x205 & ~x134 & ~x267 & ~x315;
assign c072 =  x166 &  x301 &  x312 &  x316 & ~x212;
assign c074 =  x150 & ~x228 & ~x264;
assign c076 =  x24 &  x77 & ~x129;
assign c078 =  x91 &  x208 & ~x133 & ~x157 & ~x296;
assign c080 =  x18 &  x24 & ~x95 & ~x255;
assign c082 =  x160 &  x273 & ~x284 & ~x289;
assign c084 =  x289 & ~x259 & ~x290;
assign c086 =  x206 &  x312 & ~x127;
assign c088 =  x20 & ~x174 & ~x216;
assign c090 = ~x191 & ~x218 & ~x269 & ~x283 & ~x294 & ~x320;
assign c092 =  x101 &  x303 &  x306 & ~x156 & ~x291;
assign c094 =  x76 &  x202 &  x312;
assign c096 = ~x2 & ~x65 & ~x107 & ~x192 & ~x223;
assign c098 =  x87 &  x101 &  x128 &  x232 &  x260 &  x263;
assign c0100 =  x173 &  x268 &  x311;
assign c0102 =  x121 &  x269 &  x293 & ~x271;
assign c0104 = ~x295 & ~x320 & ~x323;
assign c0106 =  x43 & ~x23 & ~x123 & ~x262;
assign c0108 =  x68 &  x73 & ~x101;
assign c0110 =  x110 &  x285 & ~x282;
assign c0112 =  x155 & ~x39 & ~x275;
assign c0114 =  x31 &  x290 & ~x43 & ~x59;
assign c0116 =  x114 &  x154 & ~x39 & ~x111 & ~x138;
assign c0118 =  x96 &  x258 &  x290 & ~x7 & ~x111;
assign c0120 = ~x263 & ~x269;
assign c0122 =  x199 & ~x228 & ~x236 & ~x237 & ~x286 & ~x317;
assign c0124 =  x239 &  x267 & ~x241 & ~x291;
assign c0126 =  x212 &  x226 & ~x116;
assign c0128 =  x279 &  x315 & ~x280;
assign c0130 =  x186 & ~x273 & ~x313;
assign c0132 =  x16 & ~x63 & ~x105 & ~x106;
assign c0134 =  x25 & ~x100 & ~x103 & ~x104;
assign c0136 = ~x143 & ~x160 & ~x321 & ~x323;
assign c0138 =  x10 &  x96 &  x131 &  x323 & ~x250;
assign c0140 = ~x120 & ~x149 & ~x152 & ~x184 & ~x287;
assign c0142 =  x157 &  x267 &  x269 &  x312;
assign c0144 =  x18 &  x105 &  x106 & ~x129 & ~x277;
assign c0146 =  x103 &  x132 &  x316 & ~x7;
assign c0148 =  x258 &  x266 & ~x144 & ~x300;
assign c0150 =  x100 &  x128 &  x132 & ~x120 & ~x255;
assign c0152 =  x191 &  x289 & ~x295;
assign c0154 =  x97 &  x137 &  x160 &  x268 &  x294 & ~x118;
assign c0156 =  x117 &  x234 &  x302 & ~x201;
assign c0158 = ~x10 & ~x19 & ~x37 & ~x105 & ~x186 & ~x212;
assign c0160 =  x19 & ~x254 & ~x316;
assign c0162 =  x123 & ~x68 & ~x212;
assign c0164 =  x76 &  x133 &  x215 &  x294 &  x321;
assign c0166 =  x40 &  x94 & ~x208;
assign c0168 =  x87 &  x101 &  x123 &  x213 & ~x295;
assign c0170 =  x101 &  x175 & ~x48;
assign c0172 =  x24 &  x41 &  x253 & ~x130;
assign c0174 =  x105 & ~x295 & ~x323;
assign c0176 = ~x9 & ~x150 & ~x193 & ~x319;
assign c0178 =  x80 &  x313 &  x317;
assign c0180 =  x24 &  x103 &  x168 &  x312;
assign c0182 =  x159 &  x267 & ~x55 & ~x302;
assign c0184 =  x133 &  x269 & ~x221;
assign c0186 =  x193 &  x213 &  x316 & ~x251;
assign c0188 =  x203 &  x298 & ~x237 & ~x322;
assign c0190 =  x159 &  x316 & ~x244;
assign c0192 =  x105 &  x267 & ~x129 & ~x286;
assign c0194 =  x92 &  x155 & ~x53 & ~x99 & ~x130;
assign c0196 =  x24 &  x96 &  x263 &  x305;
assign c0198 =  x46 & ~x34 & ~x58 & ~x305;
assign c0200 =  x4 &  x148 &  x197 &  x315 & ~x225;
assign c0202 =  x67 &  x127 &  x177 & ~x286;
assign c0204 =  x129 & ~x46 & ~x105;
assign c0206 =  x16 &  x21 & ~x283 & ~x306;
assign c0208 =  x88 & ~x100 & ~x106;
assign c0210 =  x102 &  x316 & ~x262;
assign c0212 =  x16 &  x178 & ~x104 & ~x105 & ~x107;
assign c0214 =  x289 & ~x290 & ~x319 & ~x322;
assign c0216 =  x79 & ~x229 & ~x288;
assign c0218 =  x115 &  x282 &  x295 & ~x267;
assign c0220 = ~x107 & ~x159 & ~x218 & ~x268 & ~x293 & ~x319;
assign c0222 =  x43 &  x297 & ~x223;
assign c0224 = ~x162 & ~x234 & ~x296;
assign c0226 =  x245 & ~x131 & ~x208;
assign c0228 =  x96 &  x134 &  x233 &  x310;
assign c0230 =  x21 &  x94 &  x128 & ~x107;
assign c0232 =  x109 &  x258 & ~x165;
assign c0234 =  x101 &  x310 &  x316;
assign c0236 =  x226 &  x257 & ~x304;
assign c0238 =  x84 &  x291 & ~x27 & ~x197;
assign c0240 =  x105 &  x159 &  x310 & ~x194;
assign c0242 =  x172 & ~x156 & ~x255 & ~x264 & ~x317;
assign c0244 =  x271 & ~x197 & ~x259 & ~x266;
assign c0246 =  x16 &  x151 &  x250 &  x259 & ~x36 & ~x127 & ~x257;
assign c0248 =  x96 &  x161 & ~x23 & ~x178;
assign c0250 =  x315 & ~x84 & ~x190;
assign c0252 =  x49 &  x70 &  x102 & ~x73 & ~x118;
assign c0254 = ~x76 & ~x105 & ~x117 & ~x153;
assign c0256 =  x123 &  x150 &  x312 & ~x84;
assign c0258 =  x48 &  x318 & ~x5 & ~x40;
assign c0260 =  x106 &  x294 & ~x117 & ~x120 & ~x140;
assign c0262 =  x263 & ~x181 & ~x212 & ~x217;
assign c0264 =  x11 & ~x256 & ~x278 & ~x279 & ~x284;
assign c0266 =  x128 &  x248 &  x316 & ~x198;
assign c0268 =  x158 &  x159 &  x161 &  x267 &  x287 & ~x280;
assign c0270 = ~x152 & ~x265 & ~x316;
assign c0272 = ~x241 & ~x263 & ~x296;
assign c0274 = ~x39 & ~x138 & ~x273 & ~x291;
assign c0276 =  x105 &  x292 &  x296 &  x316;
assign c0278 =  x55;
assign c0280 = ~x101 & ~x125 & ~x134 & ~x151;
assign c0282 =  x163 & ~x295 & ~x318 & ~x322;
assign c0284 =  x56 &  x213 &  x227 & ~x153;
assign c0286 =  x70 &  x178 &  x320 & ~x39 & ~x111;
assign c0288 =  x58 &  x121 &  x266 & ~x174;
assign c0290 =  x191 &  x289 &  x302;
assign c0292 = ~x213 & ~x247 & ~x310;
assign c0294 =  x101 &  x133 &  x269;
assign c0296 =  x87 &  x148 &  x204 &  x231 &  x316;
assign c0298 = ~x175 & ~x305;
assign c0300 =  x87 &  x96 &  x101 &  x128 & ~x48;
assign c0302 =  x26 &  x95 &  x162 & ~x75;
assign c0304 =  x97 &  x112 &  x193 &  x295;
assign c0306 =  x102 &  x222 &  x311 & ~x319;
assign c0308 =  x96 &  x268 & ~x255 & ~x271;
assign c0310 =  x33 &  x87 &  x123 &  x307 & ~x66;
assign c0312 =  x195 &  x289 & ~x201 & ~x237 & ~x295;
assign c0314 = ~x6 & ~x109 & ~x219 & ~x274;
assign c0316 =  x180 & ~x56 & ~x101 & ~x323;
assign c0318 =  x207 &  x258 & ~x129;
assign c0320 =  x80 &  x101 &  x215 &  x287 &  x312;
assign c0322 =  x155 &  x215 &  x290 &  x308 & ~x275;
assign c0324 =  x142 & ~x0 & ~x51 & ~x240;
assign c0326 = ~x126 & ~x129 & ~x157 & ~x252 & ~x256;
assign c0328 =  x122 &  x303 & ~x291 & ~x318;
assign c0330 =  x148 &  x285 & ~x111;
assign c0332 = ~x0 & ~x137 & ~x191 & ~x201;
assign c0334 =  x258 &  x312 & ~x120 & ~x145 & ~x250;
assign c0336 =  x20 &  x42 &  x47 &  x87 &  x142 & ~x217;
assign c0338 = ~x27 & ~x65 & ~x173 & ~x200 & ~x238 & ~x267 & ~x294;
assign c0340 = ~x63 & ~x162 & ~x208;
assign c0342 =  x160 & ~x64 & ~x111;
assign c0344 =  x104 & ~x94 & ~x167 & ~x264;
assign c0346 =  x53 &  x90 &  x206 &  x213;
assign c0348 =  x182 & ~x144 & ~x153 & ~x185;
assign c0350 =  x133 & ~x241 & ~x300;
assign c0352 = ~x105 & ~x186 & ~x288;
assign c0354 =  x132 &  x308 &  x319 & ~x34;
assign c0356 =  x44 & ~x101 & ~x102 & ~x103 & ~x294;
assign c0358 =  x307 & ~x248 & ~x275;
assign c0360 =  x20 &  x24 &  x119 &  x209 &  x258;
assign c0362 =  x42 &  x96 &  x117 &  x240 &  x269;
assign c0364 =  x290 & ~x154 & ~x262;
assign c0366 =  x114 &  x211 & ~x250;
assign c0368 = ~x6 & ~x37 & ~x157 & ~x220;
assign c0370 =  x178 &  x243 & ~x192 & ~x301;
assign c0372 =  x265 & ~x93 & ~x275 & ~x302;
assign c0374 =  x62 &  x76 & ~x273;
assign c0376 =  x40 &  x49 &  x51 &  x312 & ~x199;
assign c0378 =  x21 &  x79 & ~x169;
assign c0380 =  x256 &  x260 & ~x43;
assign c0382 =  x32 & ~x202 & ~x253 & ~x265;
assign c0384 =  x181 & ~x24 & ~x28 & ~x274;
assign c0386 =  x158 &  x208 & ~x130;
assign c0388 = ~x115 & ~x120 & ~x135 & ~x207;
assign c0390 =  x33 &  x134 &  x154 &  x265 &  x289;
assign c0392 =  x27 &  x96 &  x106 &  x123 & ~x115;
assign c0394 = ~x0 & ~x9 & ~x195 & ~x220 & ~x238;
assign c0396 =  x102 &  x121 &  x168 &  x316 & ~x271;
assign c0398 = ~x89 & ~x259 & ~x314 & ~x322;
assign c0400 =  x12 &  x16 & ~x6 & ~x121;
assign c0402 =  x160 &  x236 & ~x117 & ~x123;
assign c0404 =  x101 &  x258 & ~x2;
assign c0406 =  x77 &  x284 & ~x241 & ~x286 & ~x290;
assign c0408 =  x26 &  x240 &  x321 & ~x68 & ~x248;
assign c0410 = ~x0 & ~x24 & ~x268 & ~x269;
assign c0412 = ~x129 & ~x241 & ~x317 & ~x318 & ~x321;
assign c0414 =  x285 & ~x248 & ~x280;
assign c0416 =  x12 &  x273 & ~x87 & ~x193;
assign c0418 =  x128 &  x150 & ~x86 & ~x120;
assign c0420 =  x67 &  x121 &  x238;
assign c0422 =  x42 &  x123 &  x268 &  x293;
assign c0424 =  x110 &  x132 & ~x255 & ~x256;
assign c0426 =  x118 & ~x124 & ~x312;
assign c0428 = ~x95 & ~x158 & ~x261 & ~x262;
assign c0430 =  x159 &  x263 &  x321 & ~x302;
assign c0432 =  x24 &  x87 &  x102 &  x175 & ~x136;
assign c0434 =  x182 & ~x223;
assign c0436 =  x102 &  x150 &  x292;
assign c0438 =  x294 & ~x100 & ~x131 & ~x248;
assign c0440 =  x183 & ~x55 & ~x227 & ~x254 & ~x301;
assign c0442 = ~x197 & ~x216 & ~x233 & ~x242 & ~x269;
assign c0444 =  x56 &  x200 & ~x77 & ~x248;
assign c0446 =  x33 &  x103 &  x133 & ~x226;
assign c0448 =  x312 & ~x113 & ~x203 & ~x253;
assign c0450 =  x202 &  x236 & ~x298;
assign c0452 =  x106 &  x132 &  x150 & ~x250 & ~x275;
assign c0454 = ~x217 & ~x266 & ~x284 & ~x307;
assign c0456 =  x68 & ~x295 & ~x296;
assign c0458 =  x19 &  x25 &  x230 & ~x1 & ~x313;
assign c0460 = ~x130 & ~x148 & ~x152 & ~x242 & ~x256 & ~x265;
assign c0462 =  x38 &  x259 & ~x198;
assign c0464 =  x203 & ~x10 & ~x133 & ~x222 & ~x301 & ~x311;
assign c0466 =  x101 &  x102 &  x316 & ~x84;
assign c0468 =  x158 &  x168 & ~x48;
assign c0470 =  x30 & ~x96 & ~x150 & ~x274;
assign c0472 = ~x71 & ~x148 & ~x188 & ~x269 & ~x283;
assign c0474 = ~x18 & ~x131 & ~x154 & ~x262;
assign c0476 = ~x4 & ~x206 & ~x306;
assign c0478 =  x22 &  x150 & ~x216;
assign c0480 =  x321 & ~x48 & ~x194;
assign c0482 =  x123 &  x134 &  x240 &  x276;
assign c0484 =  x60 &  x76 &  x196 &  x310;
assign c0486 = ~x5 & ~x32 & ~x201 & ~x306;
assign c0488 =  x230 & ~x148 & ~x184 & ~x306;
assign c0490 =  x133 &  x268 &  x323 & ~x286;
assign c0492 =  x128 & ~x100 & ~x318;
assign c0494 = ~x57 & ~x223 & ~x259 & ~x274;
assign c0496 = ~x0 & ~x169 & ~x192 & ~x219;
assign c0498 =  x35 &  x97 &  x316 & ~x262;
assign c0500 =  x312 &  x316 & ~x91 & ~x118 & ~x253;
assign c0502 =  x24 &  x33 &  x152;
assign c0504 =  x65 & ~x50 & ~x318;
assign c0506 =  x259 & ~x127 & ~x145 & ~x243;
assign c0508 =  x96 &  x101 &  x128 &  x148;
assign c0510 =  x79 & ~x99 & ~x105 & ~x126 & ~x132 & ~x268;
assign c0512 =  x128 &  x193 &  x293;
assign c0514 =  x40 &  x107 &  x316;
assign c0516 =  x71 &  x148 &  x152 & ~x221;
assign c0518 =  x5 &  x25 & ~x230 & ~x280;
assign c0520 =  x76 &  x97 & ~x73 & ~x271;
assign c0522 =  x240 &  x263 &  x290 & ~x10;
assign c0524 =  x22 &  x96 &  x101 & ~x183 & ~x246;
assign c0526 =  x312 & ~x160 & ~x265 & ~x268;
assign c0528 = ~x68 & ~x111 & ~x255;
assign c0530 = ~x160 & ~x241 & ~x300 & ~x319;
assign c0532 =  x214 & ~x105 & ~x107 & ~x288;
assign c0534 =  x264 & ~x96 & ~x99 & ~x106 & ~x127;
assign c0536 =  x206 &  x240 & ~x39;
assign c0538 = ~x113 & ~x201 & ~x217 & ~x248;
assign c0540 = ~x45;
assign c0542 =  x105 &  x132 & ~x21 & ~x124 & ~x286;
assign c0544 =  x164 &  x230 &  x240;
assign c0546 =  x22 &  x24 & ~x271;
assign c0548 = ~x269 & ~x285;
assign c0550 =  x196 &  x269 &  x312 & ~x275;
assign c0552 =  x11 &  x209 & ~x162 & ~x296;
assign c0554 =  x161 &  x265 & ~x1;
assign c0556 =  x128 &  x191 & ~x291;
assign c0558 =  x27 &  x139 & ~x149;
assign c0560 =  x25 &  x70 &  x129 &  x178 & ~x32;
assign c0562 = ~x1 & ~x152 & ~x163 & ~x259 & ~x263;
assign c0564 =  x97 & ~x54 & ~x288 & ~x289;
assign c0566 = ~x36 & ~x95 & ~x104 & ~x105 & ~x127;
assign c0568 =  x132 & ~x152 & ~x228;
assign c0570 = ~x17 & ~x219 & ~x245 & ~x298;
assign c0572 = ~x61 & ~x65 & ~x162 & ~x223;
assign c0574 =  x258 &  x290 &  x317 & ~x138 & ~x271;
assign c0576 =  x6 &  x157 &  x215 &  x247;
assign c0578 = ~x86 & ~x113 & ~x131 & ~x261 & ~x279;
assign c0580 =  x177 &  x231 & ~x237;
assign c0582 =  x67 &  x150 &  x186 &  x258 &  x285;
assign c0584 = ~x8 & ~x86 & ~x155 & ~x265;
assign c0586 =  x192 &  x219 &  x294 & ~x280 & ~x309;
assign c0588 =  x11 &  x25 &  x52 &  x65 &  x259 & ~x19 & ~x153;
assign c0590 =  x195 &  x219 &  x315;
assign c0592 =  x208 & ~x128 & ~x151 & ~x319;
assign c0594 =  x120 & ~x28 & ~x78 & ~x162 & ~x228;
assign c0596 =  x306 & ~x179 & ~x319 & ~x322;
assign c0598 = ~x1 & ~x30 & ~x56 & ~x106 & ~x188 & ~x192;
assign c01 =  x85 &  x239 &  x288;
assign c03 =  x28 &  x139 & ~x33;
assign c05 =  x279 & ~x96 & ~x285;
assign c07 =  x219 &  x229 &  x239 &  x301 & ~x110;
assign c09 = ~x90 & ~x192 & ~x239 & ~x274;
assign c011 =  x165 &  x318 & ~x198;
assign c013 =  x279 & ~x238 & ~x239 & ~x323;
assign c015 =  x60 &  x168 & ~x92 & ~x186;
assign c017 =  x212 &  x285 & ~x21 & ~x209;
assign c019 =  x55 &  x190 &  x219 & ~x49 & ~x184 & ~x256;
assign c021 =  x3 &  x174 & ~x69 & ~x141;
assign c023 =  x228 &  x233 & ~x173;
assign c025 = ~x17 & ~x54 & ~x231;
assign c027 =  x98 &  x173 & ~x209 & ~x303;
assign c029 =  x26 &  x156 &  x240 &  x291;
assign c031 =  x45 &  x109 & ~x141 & ~x142;
assign c033 =  x11 &  x289 & ~x98;
assign c035 =  x59 & ~x35 & ~x89;
assign c037 = ~x90 & ~x94 & ~x103 & ~x225 & ~x297;
assign c039 =  x319 & ~x24 & ~x135;
assign c041 =  x55 &  x190 &  x218 &  x219 &  x322 & ~x40;
assign c043 =  x291 & ~x286;
assign c045 = ~x212 & ~x224 & ~x238 & ~x239 & ~x297;
assign c047 =  x125 &  x301 & ~x42;
assign c049 =  x192 & ~x69 & ~x315 & ~x320;
assign c051 =  x125 & ~x69 & ~x70 & ~x114 & ~x177;
assign c053 =  x68 &  x271 &  x295 &  x297;
assign c055 =  x116 &  x179 &  x250 & ~x11;
assign c057 =  x70 & ~x13 & ~x209;
assign c059 =  x33 &  x42 &  x115 & ~x245;
assign c061 = ~x46 & ~x91 & ~x159 & ~x253;
assign c063 =  x18 &  x38 & ~x69 & ~x195;
assign c065 =  x9 &  x17 & ~x222;
assign c067 =  x127 &  x128 &  x263 &  x289 & ~x240;
assign c069 =  x54 &  x322 & ~x315;
assign c071 =  x100 &  x119 &  x228 & ~x169;
assign c073 =  x210 &  x211 &  x282 &  x292;
assign c075 =  x207 &  x279 & ~x5 & ~x315;
assign c077 =  x72 &  x207 &  x253 &  x279 & ~x241 & ~x260;
assign c079 =  x174 &  x176 & ~x157;
assign c081 =  x49 &  x291 & ~x17 & ~x53;
assign c083 =  x25 &  x258 & ~x152 & ~x229;
assign c085 = ~x31 & ~x54 & ~x89 & ~x96 & ~x174 & ~x189;
assign c087 =  x252 & ~x69 & ~x184;
assign c089 =  x127 &  x206 & ~x247;
assign c091 =  x53 &  x108 &  x251 & ~x61;
assign c093 = ~x240 & ~x241 & ~x303 & ~x304;
assign c095 =  x122 &  x174 &  x189;
assign c097 = ~x149 & ~x231 & ~x238 & ~x239 & ~x303 & ~x310;
assign c099 =  x99 &  x288 & ~x84 & ~x171;
assign c0101 =  x147 & ~x26 & ~x89 & ~x98 & ~x261;
assign c0103 = ~x182 & ~x209 & ~x225 & ~x255;
assign c0105 =  x14 &  x45 &  x46 &  x180 &  x267;
assign c0107 =  x178 & ~x200 & ~x201 & ~x244 & ~x245;
assign c0109 =  x45 &  x125 &  x180 &  x199 &  x271 & ~x205;
assign c0111 =  x69 &  x115 & ~x20 & ~x71;
assign c0113 =  x99 &  x301 & ~x49 & ~x241;
assign c0115 =  x72 &  x207 &  x279 & ~x44 & ~x142;
assign c0117 =  x27 &  x302 &  x315;
assign c0119 = ~x17 & ~x26 & ~x89 & ~x98 & ~x190 & ~x289;
assign c0121 =  x83 & ~x80 & ~x220;
assign c0123 =  x99 & ~x171;
assign c0125 =  x85 &  x107 &  x227;
assign c0127 =  x140 &  x239 &  x311 & ~x173;
assign c0129 =  x27 & ~x142 & ~x177 & ~x214;
assign c0131 =  x144 &  x161 &  x207 & ~x242;
assign c0133 =  x34 &  x304 &  x309 & ~x207;
assign c0135 =  x48 &  x88 &  x183 &  x255 &  x292;
assign c0137 = ~x97 & ~x250 & ~x285;
assign c0139 =  x76 &  x147 &  x210 &  x211 &  x318;
assign c0141 =  x206 & ~x52 & ~x251;
assign c0143 =  x43 &  x153 & ~x173 & ~x190;
assign c0145 =  x26 &  x98 &  x237 & ~x35;
assign c0147 =  x137 &  x279 & ~x128 & ~x238;
assign c0149 =  x13 &  x84 &  x93 & ~x80 & ~x152;
assign c0151 =  x9 &  x17 &  x89 & ~x22 & ~x180;
assign c0153 =  x54 &  x166 & ~x98;
assign c0155 =  x2 &  x3 &  x12 & ~x245 & ~x278;
assign c0157 = ~x87 & ~x88 & ~x308;
assign c0159 =  x210 & ~x303 & ~x322;
assign c0161 =  x184 &  x248 & ~x74 & ~x208;
assign c0163 =  x144 &  x161 &  x279 & ~x10 & ~x173;
assign c0165 =  x44 &  x48 &  x183 &  x205 &  x277 & ~x64;
assign c0167 =  x219 &  x220 &  x238 &  x318;
assign c0169 =  x147 &  x219 & ~x89;
assign c0171 = ~x50 & ~x70 & ~x76;
assign c0173 =  x202 &  x219 & ~x195;
assign c0175 =  x56 &  x278 & ~x231;
assign c0177 =  x5 & ~x67 & ~x198 & ~x200;
assign c0179 =  x291 &  x305 & ~x90 & ~x144;
assign c0181 =  x127 &  x155 &  x235 & ~x116 & ~x251;
assign c0183 =  x21 &  x93 & ~x53 & ~x78 & ~x188;
assign c0185 =  x236 &  x253 & ~x18;
assign c0187 =  x9 &  x26 &  x29 &  x174;
assign c0189 =  x48 &  x251 & ~x18;
assign c0191 =  x256 & ~x23 & ~x26 & ~x95 & ~x102;
assign c0193 =  x34 &  x35 &  x169 & ~x290;
assign c0195 =  x22 & ~x15 & ~x321;
assign c0197 =  x3 &  x242 &  x314 & ~x76;
assign c0199 =  x121 & ~x52 & ~x138 & ~x217;
assign c0201 =  x5 &  x314 & ~x189 & ~x312;
assign c0203 =  x189 & ~x2 & ~x177 & ~x186;
assign c0205 =  x86 &  x119 &  x253 & ~x242;
assign c0207 =  x250 & ~x26 & ~x210 & ~x274;
assign c0209 =  x15 &  x87 &  x88 &  x96 & ~x180;
assign c0211 =  x32 &  x167 &  x176 & ~x10 & ~x11 & ~x56 & ~x191;
assign c0213 =  x43 &  x245 & ~x127;
assign c0215 =  x277 &  x280 &  x281 & ~x176;
assign c0217 =  x79 &  x126 &  x186 &  x250;
assign c0219 =  x6 &  x89 &  x99 & ~x71;
assign c0221 =  x39 &  x85 & ~x42;
assign c0223 =  x192 & ~x42 & ~x88;
assign c0225 =  x70 &  x210 &  x282 & ~x56;
assign c0227 = ~x72 & ~x105 & ~x132 & ~x299 & ~x321;
assign c0229 =  x55 &  x57 &  x139;
assign c0231 =  x124 &  x142 &  x153;
assign c0233 =  x12 & ~x136 & ~x270;
assign c0235 =  x95 &  x102 &  x225 &  x302;
assign c0237 = ~x228 & ~x238 & ~x239 & ~x297;
assign c0239 =  x220 &  x229 &  x230 &  x238 &  x301 &  x302;
assign c0241 =  x72 &  x144 &  x279 & ~x158 & ~x229 & ~x239 & ~x311;
assign c0243 =  x91 &  x109 &  x283;
assign c0245 = ~x16 & ~x114 & ~x295;
assign c0247 =  x26 &  x30 & ~x251;
assign c0249 =  x109 &  x135 &  x136 &  x282 & ~x50;
assign c0251 =  x284 & ~x71 & ~x175 & ~x248;
assign c0253 =  x26 &  x99 & ~x208 & ~x281;
assign c0255 =  x46 &  x109 & ~x44 & ~x179 & ~x250;
assign c0257 =  x201 & ~x49 & ~x72 & ~x199;
assign c0259 =  x39 &  x311 &  x319;
assign c0261 =  x223 & ~x56 & ~x172 & ~x200;
assign c0263 =  x169 &  x256 & ~x156;
assign c0265 =  x210 &  x246 &  x273 & ~x171;
assign c0267 =  x24 &  x279 & ~x13 & ~x85 & ~x290;
assign c0269 =  x5 &  x48 &  x49 &  x121 & ~x87;
assign c0271 =  x95 &  x180 &  x268 & ~x237;
assign c0273 =  x85 &  x194 &  x201 & ~x50 & ~x213;
assign c0275 =  x59 &  x140 &  x212;
assign c0277 =  x202 &  x210 &  x211 &  x273 & ~x69;
assign c0279 = ~x105 & ~x141 & ~x321;
assign c0281 =  x122 & ~x233 & ~x234;
assign c0283 =  x124 & ~x256 & ~x306 & ~x314;
assign c0285 =  x113 & ~x84 & ~x200 & ~x299;
assign c0287 =  x205 & ~x26 & ~x216 & ~x225;
assign c0289 =  x6 &  x48 &  x111 &  x207;
assign c0291 =  x206 &  x253 &  x279 & ~x12;
assign c0293 =  x1 &  x142 &  x253 &  x277;
assign c0295 =  x121 &  x256 & ~x5 & ~x294;
assign c0297 =  x99 & ~x175 & ~x184 & ~x246 & ~x247;
assign c0299 =  x23 &  x86 &  x306 & ~x256;
assign c0301 =  x109 &  x155 & ~x250;
assign c0303 =  x0 &  x8 &  x58 &  x176;
assign c0305 =  x48 & ~x63 & ~x71;
assign c0307 =  x3 &  x4 &  x12 &  x39 &  x40 &  x112;
assign c0309 =  x37 &  x149 & ~x184 & ~x249;
assign c0311 = ~x75 & ~x213 & ~x288;
assign c0313 =  x129 &  x263 & ~x256;
assign c0315 =  x0 &  x8 & ~x62 & ~x168;
assign c0317 =  x53 &  x93 &  x125 & ~x141;
assign c0319 =  x1 &  x207 &  x226 &  x279;
assign c0321 =  x249 & ~x26 & ~x53 & ~x162 & ~x179;
assign c0323 =  x205 & ~x50 & ~x270;
assign c0325 =  x47 &  x207 &  x226 &  x254;
assign c0327 =  x4 &  x5 &  x13 &  x39 &  x246;
assign c0329 =  x55 &  x190 &  x230 &  x239 &  x318;
assign c0331 =  x130 &  x150 &  x212 & ~x166;
assign c0333 =  x42 &  x86 &  x114 & ~x37 & ~x109 & ~x246;
assign c0335 =  x131 & ~x216 & ~x224 & ~x225;
assign c0337 =  x115 &  x132 &  x251 & ~x98;
assign c0339 =  x145 &  x213 &  x289 &  x290 & ~x179;
assign c0341 =  x136 &  x168 &  x198 &  x243;
assign c0343 =  x27 &  x37 &  x171 &  x192;
assign c0345 =  x212 & ~x74 & ~x92 & ~x145 & ~x280;
assign c0347 = ~x0 & ~x26 & ~x52 & ~x192 & ~x227 & ~x309;
assign c0349 =  x141 &  x144 &  x219;
assign c0351 =  x33 &  x170 &  x215;
assign c0353 = ~x16 & ~x182 & ~x254 & ~x280;
assign c0355 =  x14 &  x177 & ~x38 & ~x182 & ~x272;
assign c0357 =  x1 &  x90 &  x134 & ~x154;
assign c0359 =  x167 &  x321 & ~x22 & ~x94;
assign c0361 =  x265 & ~x137 & ~x209 & ~x223;
assign c0363 =  x139 &  x275 & ~x242;
assign c0365 =  x35 &  x113 &  x129 &  x170 & ~x300;
assign c0367 = ~x51 & ~x56 & ~x57 & ~x226;
assign c0369 =  x229 & ~x105 & ~x299;
assign c0371 =  x31 &  x277 & ~x26;
assign c0373 =  x57 &  x248 & ~x179 & ~x237;
assign c0375 =  x153 &  x217 &  x289 & ~x61;
assign c0377 =  x108 &  x135 &  x252 & ~x155;
assign c0379 =  x124 &  x187 &  x218 & ~x197;
assign c0381 =  x141 & ~x36 & ~x179 & ~x318;
assign c0383 =  x91 &  x128 & ~x85 & ~x98;
assign c0385 =  x100 & ~x23 & ~x177;
assign c0387 =  x112 &  x113 &  x175 &  x176 & ~x221;
assign c0389 =  x268 &  x269 & ~x155 & ~x316;
assign c0391 =  x69 &  x203 &  x223 & ~x179;
assign c0393 =  x1 &  x30 &  x165 &  x237;
assign c0395 =  x88 &  x91 &  x138 & ~x22 & ~x94;
assign c0397 =  x30 &  x194 &  x221 & ~x148;
assign c0399 =  x286 & ~x21 & ~x209 & ~x280;
assign c0401 =  x88 &  x92 &  x137 &  x218;
assign c0403 =  x70 & ~x3 & ~x12 & ~x13 & ~x21;
assign c0405 =  x0 &  x2 &  x9 &  x228;
assign c0407 =  x68 &  x144 &  x207 &  x264 &  x279;
assign c0409 =  x111 &  x112 &  x257 & ~x15;
assign c0411 =  x134 & ~x30 & ~x51 & ~x214 & ~x241;
assign c0413 = ~x22 & ~x84 & ~x93 & ~x180 & ~x315;
assign c0415 =  x134 &  x189 & ~x154;
assign c0417 =  x39 &  x40 &  x112 &  x174 &  x242;
assign c0419 =  x201 & ~x20 & ~x152;
assign c0421 =  x28 &  x163 &  x192 & ~x61 & ~x168;
assign c0423 =  x45 &  x125 &  x171 &  x199;
assign c0425 =  x54 &  x190 &  x219 & ~x168;
assign c0427 =  x45 &  x53 &  x125 & ~x71;
assign c0429 =  x79 &  x151 &  x228 &  x288;
assign c0431 =  x128 &  x154 &  x289 & ~x105 & ~x231 & ~x303;
assign c0433 =  x70 &  x318 & ~x23 & ~x144;
assign c0435 =  x114 &  x127 &  x264 & ~x110 & ~x245;
assign c0437 =  x234 &  x306 & ~x37 & ~x171 & ~x213;
assign c0439 =  x46 & ~x40 & ~x61 & ~x62 & ~x112;
assign c0441 =  x141 & ~x23 & ~x26 & ~x98;
assign c0443 =  x275 &  x290 &  x291 & ~x71;
assign c0445 =  x142 &  x205 & ~x165 & ~x173 & ~x267;
assign c0447 =  x1 &  x158 & ~x303;
assign c0449 =  x68 &  x279 & ~x111 & ~x112;
assign c0451 =  x310 &  x319 & ~x42 & ~x135;
assign c0453 =  x167 & ~x51 & ~x124 & ~x284;
assign c0455 =  x85 &  x108 &  x136 & ~x156;
assign c0457 =  x14 &  x50 &  x86 &  x94 & ~x200;
assign c0459 =  x29 &  x164 &  x278;
assign c0461 =  x78 &  x232 &  x234 &  x306;
assign c0463 =  x251 & ~x23 & ~x102 & ~x225;
assign c0465 =  x29 &  x126 &  x157 &  x158 &  x173;
assign c0467 =  x283 & ~x14 & ~x93 & ~x279;
assign c0469 =  x82 &  x293 & ~x179;
assign c0471 =  x14 &  x81 &  x99;
assign c0473 =  x8 &  x27 & ~x245;
assign c0475 =  x55 &  x192 &  x219 & ~x0;
assign c0477 =  x35 &  x54 &  x62 &  x197 &  x265;
assign c0479 =  x118 &  x253 &  x281 & ~x213 & ~x241 & ~x285;
assign c0481 =  x48 &  x154 & ~x50;
assign c0483 =  x5 &  x90 &  x219;
assign c0485 =  x192 &  x219 & ~x5 & ~x6;
assign c0487 =  x95 &  x233 &  x306 & ~x11;
assign c0489 =  x250 &  x261 & ~x238;
assign c0491 =  x53 &  x77 &  x89 &  x149 &  x284;
assign c0493 =  x182 & ~x17 & ~x26 & ~x102 & ~x103;
assign c0495 =  x271 &  x301 &  x310 &  x318;
assign c0497 =  x55 &  x163 &  x164 &  x275 & ~x180 & ~x252;
assign c0499 =  x39 &  x41 &  x151 &  x174;
assign c0501 =  x70 &  x205 &  x206 & ~x38 & ~x307;
assign c0503 =  x224 &  x225 &  x305 & ~x42 & ~x177;
assign c0505 = ~x163 & ~x171 & ~x194 & ~x306;
assign c0507 =  x2 &  x28 &  x122 &  x190 &  x218 & ~x176;
assign c0509 =  x129 &  x298 & ~x175;
assign c0511 =  x93 &  x186 &  x263 &  x288;
assign c0513 =  x75 &  x138 &  x270 & ~x44;
assign c0515 =  x14 &  x90 &  x99 &  x216 &  x297;
assign c0517 =  x11 &  x30 &  x165 &  x272 & ~x69;
assign c0519 =  x167 & ~x29 & ~x231 & ~x241;
assign c0521 =  x99 &  x279 & ~x319;
assign c0523 =  x36 & ~x65 & ~x200 & ~x246;
assign c0525 =  x94 &  x270 & ~x39 & ~x238;
assign c0527 =  x174 &  x204 &  x246 & ~x254;
assign c0529 =  x179 & ~x297 & ~x299;
assign c0531 =  x23 &  x94 &  x223 &  x288;
assign c0533 =  x218 & ~x115 & ~x127 & ~x128;
assign c0535 =  x5 &  x48 &  x120 &  x319;
assign c0537 =  x53 &  x81 &  x116 & ~x13;
assign c0539 =  x210 &  x274 & ~x145 & ~x207;
assign c0541 =  x8 &  x171 & ~x51;
assign c0543 =  x0 &  x293 & ~x19;
assign c0545 =  x14 &  x21 &  x120 &  x145 &  x208;
assign c0547 =  x3 &  x34 &  x35 &  x232;
assign c0549 =  x41 &  x61 &  x167 & ~x69;
assign c0551 =  x48 &  x112 &  x120 &  x129 &  x183 &  x256;
assign c0553 =  x0 &  x89 & ~x303;
assign c0555 =  x32 &  x124 &  x136 &  x271 & ~x164;
assign c0557 = ~x188 & ~x196 & ~x221 & ~x260;
assign c0559 =  x36 &  x108 & ~x47 & ~x73 & ~x182 & ~x209;
assign c0561 =  x49 &  x205 &  x318;
assign c0563 =  x77 &  x149 & ~x67 & ~x139;
assign c0565 =  x50 &  x248 & ~x39 & ~x53 & ~x259;
assign c0567 =  x49 &  x122 &  x315 & ~x26 & ~x97;
assign c0569 =  x77 &  x122 &  x149 &  x212 &  x290 & ~x245;
assign c0571 = ~x26 & ~x90 & ~x98 & ~x229 & ~x235 & ~x297;
assign c0573 =  x205 &  x210 & ~x302;
assign c0575 =  x82 & ~x139 & ~x186 & ~x274;
assign c0577 =  x75 &  x132 &  x210 &  x282 & ~x22;
assign c0579 =  x146 &  x198 &  x224 &  x270 &  x271 &  x281;
assign c0581 =  x60 &  x305 & ~x186 & ~x258 & ~x322;
assign c0583 =  x230 &  x261 &  x300 &  x311;
assign c0585 =  x232 & ~x227 & ~x299;
assign c0587 =  x34 &  x89 &  x99 &  x246;
assign c0589 =  x13 &  x48 &  x120 &  x319;
assign c0591 =  x82 & ~x79 & ~x305;
assign c0593 =  x26 &  x198 &  x264;
assign c0595 =  x117 &  x164 & ~x214;
assign c0597 =  x224 &  x233 & ~x29 & ~x56 & ~x162;
assign c0599 = ~x72 & ~x207 & ~x249;
assign c10 =  x250 &  x262 & ~x69;
assign c12 =  x69 &  x234 & ~x112;
assign c14 =  x130 & ~x31 & ~x209;
assign c16 =  x141 &  x264 & ~x238 & ~x295;
assign c18 =  x168 & ~x116 & ~x216;
assign c110 =  x306 & ~x213 & ~x261;
assign c112 =  x31 &  x64 &  x135 &  x189 &  x270;
assign c114 =  x93 &  x126 &  x127 &  x129;
assign c116 = ~x75 & ~x76 & ~x225 & ~x234;
assign c118 = ~x22 & ~x72 & ~x224 & ~x234 & ~x297;
assign c120 =  x205 & ~x17 & ~x26 & ~x98 & ~x226;
assign c122 = ~x17 & ~x24 & ~x96 & ~x105 & ~x320;
assign c124 =  x234 &  x291 & ~x112;
assign c126 =  x253 & ~x43 & ~x116 & ~x178 & ~x282;
assign c128 =  x164 &  x218 &  x219 & ~x60 & ~x195 & ~x196;
assign c130 =  x53 &  x125 &  x151 &  x291;
assign c132 =  x0 &  x176 & ~x148;
assign c134 =  x148 &  x210 &  x283 & ~x252;
assign c136 =  x237 &  x300 &  x301 &  x304;
assign c138 =  x234 &  x235 & ~x116 & ~x173;
assign c140 =  x55 &  x77 &  x149 &  x318;
assign c142 =  x146 & ~x180 & ~x186;
assign c144 =  x127 & ~x18 & ~x301;
assign c146 =  x41 & ~x100 & ~x127 & ~x128 & ~x155 & ~x290;
assign c148 =  x275 & ~x26 & ~x74 & ~x319;
assign c150 =  x238 &  x310 &  x318;
assign c152 =  x53 &  x125 &  x134 & ~x104;
assign c154 =  x212 &  x292 & ~x47 & ~x74 & ~x254;
assign c156 =  x41 & ~x83 & ~x110 & ~x231;
assign c158 =  x217 &  x219 &  x220 &  x302;
assign c160 =  x165 &  x316 &  x318;
assign c162 =  x183 & ~x45 & ~x117 & ~x180 & ~x252 & ~x310;
assign c164 =  x34 & ~x171 & ~x175;
assign c166 =  x86 &  x176 &  x223 & ~x56;
assign c168 =  x13 & ~x15 & ~x226;
assign c170 =  x3 &  x4 &  x21 &  x48 &  x232;
assign c172 =  x146 &  x281 & ~x23 & ~x61 & ~x168;
assign c174 =  x74 &  x85 & ~x185 & ~x191;
assign c176 =  x112 &  x175 &  x198 & ~x74;
assign c178 =  x223 & ~x241;
assign c180 =  x14 &  x78 &  x154 &  x241;
assign c182 =  x111 &  x169 & ~x270;
assign c184 =  x158 &  x284 &  x293 &  x313 & ~x112;
assign c186 =  x12 &  x187 &  x288 &  x290;
assign c188 =  x8 &  x16 &  x126 &  x153;
assign c190 =  x279 & ~x254 & ~x283;
assign c192 =  x127 &  x128 &  x156 &  x262 &  x263 &  x264 &  x291;
assign c194 =  x1 &  x127 &  x153 &  x154 &  x289;
assign c196 =  x78 &  x115 &  x165 &  x250;
assign c198 = ~x89 & ~x98 & ~x102 & ~x110;
assign c1100 =  x95 & ~x141 & ~x214;
assign c1102 =  x77 &  x149 &  x212 &  x224 &  x284;
assign c1104 =  x194 & ~x55 & ~x93 & ~x133;
assign c1106 =  x194 &  x268 &  x295 &  x322;
assign c1108 =  x77 & ~x114 & ~x214;
assign c1110 =  x252 & ~x141 & ~x237 & ~x276;
assign c1112 =  x270 &  x321 & ~x200 & ~x274;
assign c1114 =  x119 &  x127 &  x254 &  x280 & ~x188;
assign c1116 =  x75 &  x147 & ~x63 & ~x190;
assign c1118 =  x229 & ~x110 & ~x236 & ~x245;
assign c1120 =  x89 &  x99 &  x107 &  x296;
assign c1122 =  x60 &  x63 & ~x93;
assign c1124 =  x42 & ~x0 & ~x131 & ~x171;
assign c1126 =  x288 &  x323 & ~x133 & ~x160;
assign c1128 =  x118 &  x198 &  x207 &  x279 & ~x133;
assign c1130 =  x100 &  x217 &  x259;
assign c1132 =  x100 &  x201 &  x273 & ~x49 & ~x121;
assign c1134 =  x34 &  x203 &  x304 & ~x90;
assign c1136 =  x252 &  x253 & ~x213 & ~x286;
assign c1138 =  x15 &  x69 &  x144 &  x279 & ~x128;
assign c1140 =  x183 & ~x24 & ~x222;
assign c1142 = ~x4 & ~x12 & ~x13 & ~x21 & ~x36 & ~x84;
assign c1144 =  x86 & ~x20 & ~x303;
assign c1146 =  x10 &  x279 & ~x238;
assign c1148 =  x69 &  x223 & ~x31 & ~x162;
assign c1150 =  x270 &  x271 & ~x44 & ~x205;
assign c1152 =  x216 &  x292 &  x302;
assign c1154 =  x242 &  x304 & ~x58 & ~x192;
assign c1156 =  x217 &  x288 & ~x46;
assign c1158 =  x18 &  x86 & ~x31;
assign c1160 =  x138 &  x149 &  x212 &  x275;
assign c1162 =  x263 & ~x135 & ~x231;
assign c1164 =  x81 & ~x20 & ~x252;
assign c1166 =  x205 &  x242 &  x314 & ~x18 & ~x298;
assign c1168 =  x93 &  x134 &  x281;
assign c1170 = ~x18 & ~x47 & ~x91 & ~x284;
assign c1172 =  x129 & ~x142 & ~x179;
assign c1174 =  x0 &  x174 &  x319 & ~x306;
assign c1176 =  x57 &  x65 &  x300 & ~x167;
assign c1178 = ~x96 & ~x114 & ~x222;
assign c1180 = ~x5 & ~x13 & ~x21 & ~x225;
assign c1182 =  x110 &  x111 & ~x46 & ~x302;
assign c1184 = ~x203 & ~x204 & ~x290;
assign c1186 =  x45 &  x243 &  x256 & ~x128;
assign c1188 =  x99 &  x194 &  x288;
assign c1190 =  x129 &  x284 & ~x178 & ~x251;
assign c1192 =  x166 &  x167 & ~x128 & ~x154;
assign c1194 =  x89 &  x98 &  x99 & ~x242;
assign c1196 =  x10 &  x255 & ~x65;
assign c1198 =  x142 &  x143 &  x220 & ~x60;
assign c1200 =  x41 & ~x38 & ~x92 & ~x298;
assign c1202 =  x70 &  x251 &  x313;
assign c1204 =  x14 &  x86 & ~x112 & ~x175 & ~x256;
assign c1206 =  x129 &  x155 &  x212 &  x263;
assign c1208 = ~x67 & ~x96 & ~x178;
assign c1210 =  x26 &  x28 &  x81 &  x164 &  x228;
assign c1212 =  x18 &  x89 & ~x171 & ~x177;
assign c1214 =  x312 & ~x182 & ~x254 & ~x290 & ~x307;
assign c1216 =  x274 & ~x234 & ~x296;
assign c1218 =  x244 &  x252 &  x273 & ~x127;
assign c1220 =  x69 & ~x0 & ~x32 & ~x44 & ~x179;
assign c1222 =  x301 &  x302 &  x310 & ~x20 & ~x92;
assign c1224 =  x142 &  x277 & ~x18 & ~x235;
assign c1226 =  x82 &  x94 & ~x215;
assign c1228 =  x113 &  x270 & ~x153;
assign c1230 =  x100 &  x117 &  x179 & ~x289;
assign c1232 =  x219 &  x318 & ~x61;
assign c1234 =  x219 & ~x212 & ~x264;
assign c1236 =  x194 &  x224 &  x234;
assign c1238 =  x55 &  x291 & ~x71;
assign c1240 =  x153 &  x217 &  x220 &  x288;
assign c1242 =  x27 &  x45 &  x108 & ~x61;
assign c1244 =  x36 &  x273 & ~x76 & ~x147;
assign c1246 =  x3 &  x27 &  x319;
assign c1248 =  x90 & ~x78 & ~x106;
assign c1250 =  x0 &  x192 &  x261 & ~x61;
assign c1252 = ~x234 & ~x238 & ~x288 & ~x297 & ~x306 & ~x315;
assign c1254 =  x266 & ~x29 & ~x173 & ~x217;
assign c1256 =  x10 &  x75 &  x210;
assign c1258 =  x4 & ~x144 & ~x194;
assign c1260 =  x201 & ~x78 & ~x146 & ~x276;
assign c1262 =  x256 &  x307 & ~x58;
assign c1264 =  x69 &  x144 &  x207 & ~x17 & ~x89;
assign c1266 =  x75 &  x283 & ~x267;
assign c1268 =  x219 & ~x98 & ~x169;
assign c1270 =  x223 &  x224 &  x234 & ~x173;
assign c1272 =  x79 &  x210 &  x218 &  x282;
assign c1274 =  x160 &  x189 &  x190 &  x270;
assign c1276 =  x149 &  x237 &  x238 &  x309;
assign c1278 =  x122 &  x140 &  x232 & ~x188;
assign c1280 =  x14 &  x302 &  x318;
assign c1282 =  x4 &  x33 &  x83 &  x174;
assign c1284 =  x70 & ~x37 & ~x66 & ~x201 & ~x272;
assign c1286 =  x53 &  x153 & ~x257;
assign c1288 =  x0 &  x89 &  x165 &  x315;
assign c1290 =  x32 &  x59 &  x68 &  x167 &  x274 &  x282;
assign c1292 =  x89 &  x100 & ~x13;
assign c1294 =  x105 &  x219 &  x230 &  x258;
assign c1296 =  x219 &  x220 &  x228 &  x301 & ~x168 & ~x195;
assign c1298 =  x305 & ~x96 & ~x281;
assign c1300 =  x139 & ~x22 & ~x93 & ~x179;
assign c1302 = ~x98 & ~x125 & ~x232;
assign c1304 =  x52 &  x194 &  x221 &  x288;
assign c1306 =  x121 &  x241 & ~x139 & ~x225;
assign c1308 =  x229 &  x273 &  x300 & ~x216;
assign c1310 =  x140 &  x222 &  x236 & ~x214;
assign c1312 =  x182 & ~x27 & ~x31 & ~x162 & ~x266;
assign c1314 =  x276 &  x313 & ~x26 & ~x173 & ~x216;
assign c1316 =  x116 &  x125 & ~x42 & ~x177;
assign c1318 =  x121 &  x218 & ~x26;
assign c1320 =  x10 &  x219 &  x228 & ~x49;
assign c1322 =  x210 &  x234 &  x282 & ~x257;
assign c1324 =  x200 &  x310 & ~x47 & ~x120 & ~x156;
assign c1326 =  x61 &  x71 &  x176 & ~x83;
assign c1328 =  x64 &  x125 &  x251 & ~x13;
assign c1330 =  x168 & ~x234 & ~x235;
assign c1332 =  x309 & ~x25 & ~x51 & ~x258;
assign c1334 =  x37 &  x244 &  x283 & ~x74 & ~x207;
assign c1336 =  x35 &  x62 &  x108;
assign c1338 =  x29 &  x69 & ~x180 & ~x252;
assign c1340 = ~x53 & ~x92 & ~x117 & ~x254;
assign c1342 =  x142 &  x143 & ~x59 & ~x98;
assign c1344 =  x95 &  x207 &  x296 & ~x35;
assign c1346 =  x19 &  x55 &  x82 &  x301;
assign c1348 =  x300 &  x311 &  x318 &  x319;
assign c1350 =  x1 &  x26 &  x89 &  x99;
assign c1352 =  x31 & ~x17 & ~x98 & ~x99;
assign c1354 =  x0 &  x8 & ~x234 & ~x303;
assign c1356 =  x220 &  x264 & ~x195;
assign c1358 =  x66 &  x138 &  x286 & ~x16;
assign c1360 =  x170 & ~x135 & ~x270;
assign c1362 =  x207 &  x208 & ~x44 & ~x169;
assign c1364 =  x139 & ~x213;
assign c1366 = ~x97 & ~x183 & ~x240 & ~x303;
assign c1368 =  x53 &  x288 & ~x168;
assign c1370 =  x21 &  x85 &  x111 & ~x58;
assign c1372 =  x108 &  x109 &  x243 & ~x184 & ~x185;
assign c1374 =  x44 &  x169 &  x179 & ~x95;
assign c1376 =  x13 &  x84 &  x85 &  x93 &  x253 & ~x152;
assign c1378 =  x39 &  x126 &  x237;
assign c1380 =  x55 &  x189 &  x198 &  x317;
assign c1382 =  x161 &  x288 & ~x160;
assign c1384 =  x112 &  x113 &  x176 &  x248 & ~x276;
assign c1386 =  x22 &  x94 & ~x25 & ~x242;
assign c1388 =  x1 &  x18 &  x86 &  x95;
assign c1390 =  x34 &  x35 &  x233 & ~x269;
assign c1392 = ~x31 & ~x35 & ~x55 & ~x148;
assign c1394 =  x99 &  x207 & ~x3 & ~x238;
assign c1396 =  x6 &  x34 &  x127 &  x128 &  x155 &  x262;
assign c1398 =  x70 &  x167 &  x178 &  x250 & ~x64 & ~x172;
assign c1400 =  x29 &  x210 & ~x278;
assign c1402 =  x34 &  x93 &  x169 & ~x67 & ~x202;
assign c1404 =  x157 &  x173 & ~x101;
assign c1406 =  x85 & ~x24 & ~x114;
assign c1408 =  x260 & ~x19 & ~x47 & ~x235;
assign c1410 =  x223 &  x235 & ~x112;
assign c1412 =  x120 &  x147 & ~x118 & ~x285;
assign c1414 =  x269 &  x270 & ~x205;
assign c1416 =  x64 &  x77 &  x125;
assign c1418 =  x72 &  x207 & ~x238 & ~x301 & ~x319;
assign c1420 =  x174 & ~x130 & ~x203 & ~x240;
assign c1422 =  x75 &  x234 &  x306 & ~x303;
assign c1424 = ~x98 & ~x192 & ~x202 & ~x216 & ~x229;
assign c1426 = ~x98 & ~x225 & ~x258;
assign c1428 =  x27 & ~x114 & ~x176 & ~x187;
assign c1430 =  x60 & ~x35 & ~x36 & ~x238;
assign c1432 =  x194 &  x223 &  x225 &  x297;
assign c1434 =  x138 &  x143 &  x220 &  x278;
assign c1436 =  x0 &  x48 & ~x103;
assign c1438 =  x38 &  x81 & ~x177 & ~x204;
assign c1440 =  x131 &  x279 &  x312 &  x320;
assign c1442 =  x212 &  x238 & ~x80;
assign c1444 =  x63 & ~x51 & ~x123 & ~x263;
assign c1446 =  x118 & ~x96 & ~x240 & ~x312;
assign c1448 =  x156 &  x297 &  x302;
assign c1450 =  x68 &  x252 & ~x38 & ~x137;
assign c1452 =  x85 &  x146 & ~x123 & ~x229;
assign c1454 =  x100 &  x207 &  x249 & ~x13;
assign c1456 =  x55 &  x218 &  x304 & ~x187;
assign c1458 =  x62 &  x218 & ~x220;
assign c1460 = ~x52 & ~x185 & ~x285 & ~x290;
assign c1462 =  x314 & ~x230 & ~x316;
assign c1464 =  x182 &  x255 & ~x18 & ~x225;
assign c1466 =  x44 &  x203 & ~x180;
assign c1468 =  x60 & ~x31 & ~x173 & ~x190;
assign c1470 =  x9 &  x201 & ~x63 & ~x270;
assign c1472 =  x66 &  x92 &  x289 &  x307;
assign c1474 =  x70 &  x142 &  x202 & ~x21;
assign c1476 =  x210 &  x304 & ~x194 & ~x216;
assign c1478 =  x85 & ~x69 & ~x70 & ~x204 & ~x205;
assign c1480 =  x69 &  x130 &  x288 & ~x172;
assign c1482 =  x108 &  x192 & ~x242;
assign c1484 =  x4 &  x5 &  x13 & ~x42;
assign c1486 =  x46 &  x119 & ~x98 & ~x315;
assign c1488 =  x0 &  x48 &  x291;
assign c1490 = ~x38 & ~x150 & ~x241 & ~x313;
assign c1492 =  x48 &  x93 & ~x28 & ~x69 & ~x276;
assign c1494 =  x75 & ~x17 & ~x84 & ~x169;
assign c1496 =  x207 & ~x25 & ~x54 & ~x97;
assign c1498 =  x230 & ~x31 & ~x166 & ~x179 & ~x197 & ~x262;
assign c1500 =  x75 &  x223 &  x234 &  x306;
assign c1502 =  x89 & ~x34 & ~x231;
assign c1504 =  x77 &  x212 &  x275 &  x284 & ~x120 & ~x254;
assign c1506 =  x158 &  x201 & ~x68 & ~x204;
assign c1508 =  x31 &  x39 &  x111 &  x313;
assign c1510 =  x232 &  x263 &  x290 & ~x29 & ~x35;
assign c1512 =  x35 &  x96 &  x142;
assign c1514 =  x217 &  x218 &  x219;
assign c1516 =  x41 &  x68 &  x207 &  x270 & ~x179;
assign c1518 =  x81 &  x98 & ~x22 & ~x142;
assign c1520 =  x135 &  x169 & ~x156 & ~x192 & ~x202;
assign c1522 =  x86 &  x206 & ~x240 & ~x312;
assign c1524 =  x146 &  x185 &  x281 & ~x42;
assign c1526 =  x224 &  x234 & ~x163 & ~x303;
assign c1528 =  x34 &  x111 &  x169 &  x237 &  x304;
assign c1530 =  x3 &  x4 &  x304 &  x319;
assign c1532 =  x8 & ~x38 & ~x104;
assign c1534 =  x99 &  x100 &  x217 &  x301;
assign c1536 =  x5 &  x48 &  x183 & ~x260;
assign c1538 =  x36 &  x37 &  x284 & ~x204;
assign c1540 =  x223 &  x226 &  x297 &  x300;
assign c1542 =  x153 &  x187 &  x261 &  x288;
assign c1544 =  x35 &  x115 &  x165 &  x182;
assign c1546 =  x174 & ~x0 & ~x282;
assign c1548 =  x270 &  x279 & ~x283 & ~x310 & ~x319;
assign c1550 =  x2 &  x16 &  x55 &  x127;
assign c1552 =  x81 &  x134 &  x212 & ~x182;
assign c1554 =  x122 &  x279 & ~x75 & ~x173;
assign c1556 =  x81 &  x191 & ~x75 & ~x148;
assign c1558 =  x9 &  x81 &  x89 &  x165 &  x174;
assign c1560 =  x39 &  x111 &  x112 &  x175 &  x184 &  x246 &  x247 & ~x22;
assign c1562 =  x277 &  x318 & ~x95;
assign c1564 =  x37 &  x238 & ~x114 & ~x141 & ~x177;
assign c1566 =  x305 & ~x64 & ~x260 & ~x301;
assign c1568 =  x0 &  x8 &  x244 & ~x262;
assign c1570 =  x84 &  x169 &  x262 & ~x71;
assign c1572 =  x14 &  x194 & ~x131 & ~x247;
assign c1574 =  x104 &  x169 & ~x234 & ~x306;
assign c1576 =  x116 &  x125 & ~x61 & ~x177;
assign c1578 =  x270 & ~x13 & ~x237 & ~x238 & ~x310;
assign c1580 =  x53 &  x108 &  x179 & ~x231;
assign c1582 =  x76 &  x211 &  x302 & ~x314;
assign c1584 =  x117 &  x295 & ~x75;
assign c1586 =  x122 &  x318 & ~x127;
assign c1588 =  x35 & ~x74 & ~x98 & ~x136;
assign c1590 = ~x4 & ~x13 & ~x21 & ~x81 & ~x300;
assign c1592 =  x138 &  x197 &  x274 & ~x177;
assign c1594 =  x30 &  x96 &  x165 &  x312 &  x313;
assign c1596 =  x135 &  x136 &  x199 &  x270 & ~x81 & ~x314;
assign c1598 =  x157 &  x265 &  x283 & ~x312;
assign c11 =  x199 &  x253 & ~x74;
assign c13 =  x20 &  x69 & ~x55 & ~x56 & ~x163 & ~x192 & ~x218 & ~x219;
assign c15 =  x7 &  x289 & ~x155 & ~x318;
assign c17 =  x94 &  x200 &  x303 & ~x226;
assign c19 =  x35 & ~x112 & ~x127;
assign c111 =  x87 &  x303 &  x307 & ~x295 & ~x322;
assign c113 = ~x33 & ~x55 & ~x101 & ~x310 & ~x319;
assign c115 =  x124 &  x264 & ~x18 & ~x19;
assign c117 =  x67 &  x96 &  x175 &  x294 & ~x84;
assign c119 =  x92 &  x150 & ~x37;
assign c121 =  x169 &  x312 &  x316;
assign c123 =  x102 &  x302 & ~x147;
assign c125 =  x65 &  x294 & ~x237;
assign c127 =  x236 & ~x154 & ~x212 & ~x252;
assign c129 =  x155 &  x247 &  x263 &  x312 &  x323;
assign c131 =  x317 & ~x32;
assign c133 =  x181 &  x212 & ~x130 & ~x134 & ~x259 & ~x265 & ~x269;
assign c135 = ~x65 & ~x78 & ~x81 & ~x159 & ~x228 & ~x267;
assign c137 =  x21 & ~x104 & ~x105 & ~x127;
assign c139 =  x229 &  x246 &  x298;
assign c141 =  x122 &  x150 & ~x156;
assign c143 =  x24 &  x123 &  x150 &  x213 &  x240 & ~x48;
assign c145 =  x93 &  x151 & ~x126 & ~x131;
assign c147 = ~x93 & ~x111 & ~x291;
assign c149 =  x105 &  x134 &  x213 & ~x120;
assign c151 =  x88 & ~x96 & ~x258 & ~x288;
assign c153 =  x304 & ~x77 & ~x127;
assign c155 =  x13 &  x312 &  x316 & ~x181;
assign c157 =  x77 & ~x5 & ~x70 & ~x129 & ~x269;
assign c159 = ~x128 & ~x227 & ~x268 & ~x305;
assign c161 =  x150 &  x209 &  x258 & ~x120;
assign c163 =  x137 &  x196 & ~x10;
assign c165 =  x14 &  x127 &  x241 & ~x82;
assign c167 =  x156 & ~x41 & ~x283;
assign c169 =  x33 & ~x99 & ~x255;
assign c171 =  x84 & ~x1 & ~x27 & ~x98 & ~x101;
assign c173 =  x83 &  x211 &  x312;
assign c175 =  x11 &  x173 &  x209 & ~x118 & ~x313;
assign c177 =  x168 &  x242 & ~x94 & ~x286;
assign c179 =  x182 & ~x154 & ~x186 & ~x283;
assign c181 =  x310 &  x315 & ~x199 & ~x208;
assign c183 = ~x60 & ~x167 & ~x266;
assign c185 =  x144 & ~x58 & ~x201 & ~x312;
assign c187 =  x103 &  x132 &  x155 & ~x275;
assign c189 =  x209 &  x259 &  x321;
assign c191 =  x50 &  x96 &  x186 & ~x84;
assign c193 =  x78 & ~x68 & ~x114;
assign c195 =  x203 & ~x129 & ~x235 & ~x263;
assign c197 =  x101 &  x161 &  x184 &  x269;
assign c199 =  x180 &  x189 &  x307 & ~x174;
assign c1101 =  x51 &  x77 &  x96 &  x123 &  x229 & ~x264;
assign c1103 =  x157 &  x161 &  x263 &  x305 &  x312;
assign c1105 =  x275 & ~x129 & ~x318;
assign c1107 =  x96 &  x132 &  x133 &  x137 &  x245 & ~x255;
assign c1109 = ~x233 & ~x257 & ~x289 & ~x303;
assign c1111 =  x112 &  x119 & ~x250;
assign c1113 =  x297 & ~x97 & ~x201 & ~x219;
assign c1115 = ~x101 & ~x124 & ~x134 & ~x259;
assign c1117 =  x127 & ~x2 & ~x8 & ~x65 & ~x163 & ~x173;
assign c1119 =  x87 &  x106 &  x154 & ~x59;
assign c1121 = ~x77 & ~x82 & ~x118 & ~x208 & ~x284;
assign c1123 =  x96 &  x99 &  x289;
assign c1125 =  x159 &  x267 & ~x151 & ~x322;
assign c1127 =  x24 &  x132 &  x242 & ~x264;
assign c1129 =  x51 &  x186 &  x242 &  x314 & ~x48;
assign c1131 =  x105 & ~x44 & ~x236 & ~x286;
assign c1133 =  x28 &  x105 & ~x147 & ~x250 & ~x313;
assign c1135 =  x51 &  x80 &  x209 &  x277 & ~x217;
assign c1137 =  x80 &  x87 &  x117 &  x128;
assign c1139 =  x102 &  x123 &  x175 &  x310;
assign c1141 =  x174 & ~x5 & ~x128 & ~x211 & ~x288;
assign c1143 =  x43 &  x214 & ~x117 & ~x134 & ~x154 & ~x266;
assign c1145 =  x289 & ~x273 & ~x277 & ~x322;
assign c1147 =  x16 &  x120 &  x187 & ~x104;
assign c1149 = ~x76 & ~x158 & ~x257 & ~x261 & ~x292;
assign c1151 =  x235 &  x249 & ~x295 & ~x319 & ~x320 & ~x322;
assign c1153 =  x187 & ~x127 & ~x132;
assign c1155 =  x154 &  x303 & ~x291 & ~x319;
assign c1157 =  x76 &  x133 &  x211 &  x294 &  x295 & ~x122;
assign c1159 =  x38 &  x239 & ~x300;
assign c1161 =  x230 & ~x99 & ~x322;
assign c1163 =  x178 & ~x0 & ~x1 & ~x162 & ~x193;
assign c1165 =  x96 & ~x264 & ~x281;
assign c1167 = ~x121 & ~x157 & ~x296 & ~x316;
assign c1169 = ~x161 & ~x192 & ~x314 & ~x316;
assign c1171 =  x263 &  x272 & ~x262;
assign c1173 =  x230 &  x284 & ~x1 & ~x313;
assign c1175 =  x140 & ~x33 & ~x114;
assign c1177 =  x212 &  x218 &  x222 &  x307 & ~x277;
assign c1179 =  x267 & ~x86 & ~x116 & ~x277;
assign c1181 =  x281 & ~x248 & ~x279 & ~x284;
assign c1183 =  x47 &  x173 &  x239 & ~x255;
assign c1185 =  x123 &  x312 & ~x226 & ~x246 & ~x271 & ~x298;
assign c1187 =  x76 &  x102 &  x133 &  x168 &  x310;
assign c1189 = ~x1 & ~x58 & ~x196 & ~x285;
assign c1191 =  x67 &  x132 &  x209 &  x238;
assign c1193 = ~x5 & ~x41 & ~x265 & ~x316;
assign c1195 =  x203 & ~x193 & ~x228 & ~x263;
assign c1197 =  x240 & ~x46 & ~x248 & ~x284;
assign c1199 =  x63 & ~x22 & ~x289;
assign c1201 =  x204 & ~x1 & ~x295 & ~x300 & ~x321;
assign c1203 =  x79 &  x315 &  x321;
assign c1205 =  x246 & ~x162 & ~x197 & ~x269;
assign c1207 =  x15 &  x125 &  x236 & ~x271;
assign c1209 =  x222 & ~x291 & ~x321 & ~x322;
assign c1211 =  x24 &  x262 &  x323 & ~x34;
assign c1213 =  x99 &  x285 & ~x298;
assign c1215 =  x218 &  x295 & ~x276 & ~x284;
assign c1217 =  x133 &  x267 & ~x16 & ~x203;
assign c1219 = ~x125 & ~x153 & ~x224 & ~x256 & ~x284;
assign c1221 =  x51 &  x78 &  x186 &  x240 &  x308;
assign c1223 =  x133 &  x292 &  x316 & ~x250;
assign c1225 =  x35 &  x67 & ~x212;
assign c1227 =  x259 & ~x91 & ~x261 & ~x274;
assign c1229 =  x33 & ~x154 & ~x212 & ~x266;
assign c1231 = ~x33 & ~x192 & ~x197;
assign c1233 =  x90 &  x316 & ~x216;
assign c1235 =  x258 &  x268 &  x293 & ~x120;
assign c1237 =  x80 &  x238 & ~x2;
assign c1239 =  x58 &  x168 &  x213 &  x223;
assign c1241 =  x24 &  x85 &  x202 &  x317 & ~x174;
assign c1243 =  x84 &  x151 & ~x154 & ~x280 & ~x289;
assign c1245 = ~x4 & ~x24 & ~x130 & ~x161;
assign c1247 =  x149 &  x275 & ~x155 & ~x211;
assign c1249 =  x71 &  x105 &  x215 &  x242;
assign c1251 =  x236 &  x272 & ~x132;
assign c1253 =  x4 &  x148 &  x285;
assign c1255 =  x102 &  x128 & ~x145 & ~x253;
assign c1257 =  x69 &  x83 &  x93 &  x276;
assign c1259 =  x96 &  x123 &  x240 & ~x115 & ~x142;
assign c1261 =  x6 & ~x99 & ~x104;
assign c1263 =  x121 &  x267 &  x268 &  x312;
assign c1265 = ~x145 & ~x257 & ~x294;
assign c1267 =  x199 & ~x211 & ~x229 & ~x312;
assign c1269 =  x121 &  x155 & ~x156;
assign c1271 =  x47 &  x187 &  x241 & ~x310;
assign c1273 = ~x201 & ~x286 & ~x318;
assign c1275 =  x25 &  x160 &  x200 & ~x100;
assign c1277 =  x213 &  x265 &  x276 &  x312 &  x316;
assign c1279 =  x154 &  x222 &  x266 & ~x291 & ~x318;
assign c1281 =  x16 &  x214 &  x270 & ~x105;
assign c1283 =  x137 &  x151 & ~x104 & ~x139;
assign c1285 =  x101 &  x123 & ~x243 & ~x273;
assign c1287 =  x213 &  x303 & ~x34 & ~x189;
assign c1289 =  x96 &  x316 & ~x115;
assign c1291 =  x133 &  x137 & ~x3 & ~x228;
assign c1293 =  x272 & ~x49 & ~x144 & ~x153 & ~x154 & ~x184 & ~x265;
assign c1295 = ~x188 & ~x263 & ~x315;
assign c1297 =  x148 &  x168 &  x197 &  x316;
assign c1299 =  x142 &  x241 & ~x27 & ~x134 & ~x192;
assign c1301 =  x164 &  x209 &  x315 & ~x255;
assign c1303 =  x105 &  x107 &  x132 & ~x124;
assign c1305 = ~x131 & ~x219 & ~x260 & ~x264 & ~x265;
assign c1307 =  x96 &  x128 &  x213 & ~x129;
assign c1309 = ~x76 & ~x160 & ~x161 & ~x274 & ~x288;
assign c1311 =  x182 & ~x203 & ~x255;
assign c1313 =  x4 &  x25 &  x294 & ~x113;
assign c1315 =  x42 &  x129 &  x168 &  x207 &  x263;
assign c1317 = ~x126 & ~x157;
assign c1319 =  x96 &  x193 &  x312;
assign c1321 =  x265 & ~x120 & ~x205;
assign c1323 =  x101 &  x161 &  x206 &  x287 &  x296;
assign c1325 =  x87 &  x148 &  x269 &  x306;
assign c1327 =  x105 &  x168 & ~x255 & ~x308;
assign c1329 =  x210 &  x322 & ~x262 & ~x280 & ~x306;
assign c1331 =  x307 &  x311 & ~x156;
assign c1333 =  x92 & ~x82 & ~x111 & ~x174;
assign c1335 =  x71 &  x96 &  x128 &  x254;
assign c1337 =  x204 & ~x217 & ~x292;
assign c1339 =  x41 &  x82 &  x195 & ~x291;
assign c1341 =  x289 & ~x99 & ~x156 & ~x291;
assign c1343 =  x106 &  x110 & ~x75;
assign c1345 =  x27 &  x133 & ~x34;
assign c1347 =  x103 &  x105 &  x197 &  x321;
assign c1349 =  x88 &  x277 & ~x0 & ~x207 & ~x216;
assign c1351 =  x231 & ~x49 & ~x80 & ~x287;
assign c1353 =  x203 & ~x0 & ~x57 & ~x300 & ~x319 & ~x320;
assign c1355 =  x150 &  x312 & ~x122;
assign c1357 =  x128 &  x141 & ~x99 & ~x246 & ~x264;
assign c1359 =  x101 &  x317 & ~x116;
assign c1361 =  x175 &  x323 & ~x221;
assign c1363 = ~x159 & ~x238 & ~x268;
assign c1365 =  x136 & ~x129 & ~x151 & ~x152 & ~x264 & ~x282;
assign c1367 = ~x5 & ~x15 & ~x28 & ~x86 & ~x272;
assign c1369 =  x20 &  x213 & ~x208;
assign c1371 =  x184 &  x290 & ~x141 & ~x248;
assign c1373 =  x31 &  x94 & ~x105;
assign c1375 =  x95 & ~x105 & ~x173 & ~x268 & ~x311 & ~x320;
assign c1377 =  x15 &  x87 &  x307 & ~x99 & ~x320;
assign c1379 =  x102 &  x168 &  x197 &  x283 &  x323;
assign c1381 =  x22 &  x103 &  x168 &  x215 &  x316;
assign c1383 =  x155 &  x300 & ~x131;
assign c1385 =  x132 &  x311 & ~x160;
assign c1387 =  x138 &  x312 & ~x86;
assign c1389 =  x103 &  x105 &  x157 & ~x217;
assign c1391 = ~x1 & ~x33 & ~x60 & ~x128;
assign c1393 = ~x128 & ~x134 & ~x159 & ~x294 & ~x315;
assign c1395 =  x56 &  x263 &  x312 & ~x305;
assign c1397 =  x19 &  x50 &  x105 &  x127;
assign c1399 = ~x57 & ~x137 & ~x264 & ~x319;
assign c1401 =  x250 &  x300 & ~x99;
assign c1403 = ~x100 & ~x118 & ~x154;
assign c1405 =  x71 & ~x168 & ~x219;
assign c1407 = ~x19 & ~x91 & ~x105 & ~x107 & ~x258;
assign c1409 =  x136 & ~x134 & ~x148 & ~x281 & ~x287;
assign c1411 =  x240 & ~x12 & ~x34 & ~x99;
assign c1413 =  x255 & ~x60 & ~x192;
assign c1415 =  x24 &  x223 & ~x138 & ~x183;
assign c1417 =  x199 & ~x120 & ~x264;
assign c1419 =  x101 &  x153 &  x317 & ~x3;
assign c1421 =  x52 &  x93 & ~x105;
assign c1423 = ~x121 & ~x148 & ~x257 & ~x288 & ~x297;
assign c1425 =  x71 &  x98 &  x188 & ~x172;
assign c1427 =  x276 & ~x244 & ~x270 & ~x297;
assign c1429 =  x96 &  x101 & ~x201;
assign c1431 =  x156 &  x291 & ~x99 & ~x132;
assign c1433 =  x80 &  x159 & ~x255;
assign c1435 =  x316 & ~x280 & ~x302;
assign c1437 =  x270 & ~x268 & ~x310 & ~x316;
assign c1439 =  x152 &  x316 &  x321;
assign c1441 =  x92 &  x150 &  x207 &  x281;
assign c1443 =  x149 & ~x241 & ~x292 & ~x322;
assign c1445 =  x50 &  x255 & ~x28 & ~x299 & ~x319;
assign c1447 =  x15 &  x33 &  x184 &  x186;
assign c1449 =  x16 &  x151 & ~x96 & ~x104;
assign c1451 =  x6 &  x11 &  x272 & ~x140;
assign c1453 =  x58 &  x166 &  x294 & ~x145;
assign c1455 =  x102 &  x240 &  x316 &  x321;
assign c1457 =  x24 &  x92 &  x123 & ~x57;
assign c1459 =  x151 &  x214 &  x232 &  x295 & ~x280;
assign c1461 =  x132 &  x266;
assign c1463 =  x49 &  x159 & ~x253;
assign c1465 =  x184 & ~x7 & ~x43 & ~x217;
assign c1467 =  x213 &  x236 & ~x304;
assign c1469 =  x240 &  x258 &  x294 & ~x282;
assign c1471 =  x117 &  x268 &  x294 & ~x250;
assign c1473 =  x42 &  x92 &  x141 &  x304 & ~x198;
assign c1475 =  x157 &  x233 &  x317;
assign c1477 =  x236 &  x260 &  x299;
assign c1479 =  x17 &  x21 &  x236;
assign c1481 =  x103 &  x240 & ~x120 & ~x203;
assign c1483 =  x166 &  x312 &  x315 & ~x280;
assign c1485 =  x123 &  x126 &  x134 &  x265 & ~x21;
assign c1487 =  x140 & ~x155 & ~x308 & ~x317 & ~x322 & ~x323;
assign c1489 =  x227 & ~x100 & ~x105;
assign c1491 =  x82 & ~x49 & ~x53 & ~x71 & ~x99;
assign c1493 =  x175 &  x312 &  x317 & ~x282;
assign c1495 =  x77 &  x137 & ~x264 & ~x317;
assign c1497 =  x17 &  x299 &  x308 & ~x63 & ~x318;
assign c1499 =  x94 &  x128 &  x148 &  x252 &  x308;
assign c1501 =  x15 &  x262 & ~x148 & ~x291 & ~x322;
assign c1503 =  x321 &  x323 & ~x122;
assign c1505 =  x74 &  x308 & ~x149 & ~x257;
assign c1507 =  x74 &  x146 & ~x153 & ~x271 & ~x319;
assign c1509 =  x50 & ~x192 & ~x293 & ~x320;
assign c1511 =  x11 & ~x39 & ~x67 & ~x123;
assign c1513 =  x185 & ~x166 & ~x265;
assign c1515 =  x266 & ~x125 & ~x290 & ~x321;
assign c1517 =  x97 &  x159 &  x184;
assign c1519 =  x150 &  x266 &  x316 &  x323;
assign c1521 =  x5 &  x33 &  x168 &  x316 & ~x298;
assign c1523 =  x171 &  x308 &  x321 & ~x115;
assign c1525 =  x87 &  x105 &  x310;
assign c1527 =  x96 &  x157 &  x266 &  x269;
assign c1529 =  x60 &  x101 &  x269 &  x293;
assign c1531 = ~x102 & ~x124 & ~x128 & ~x133 & ~x134 & ~x159 & ~x269;
assign c1533 =  x5 &  x97 & ~x145;
assign c1535 =  x242 &  x312 & ~x216 & ~x218 & ~x298;
assign c1537 =  x192 &  x198 & ~x140;
assign c1539 =  x241 & ~x64 & ~x133 & ~x136 & ~x180;
assign c1541 = ~x54 & ~x117 & ~x131 & ~x279;
assign c1543 =  x52 &  x58 &  x200;
assign c1545 =  x142 & ~x99 & ~x104 & ~x132;
assign c1547 =  x298 & ~x146 & ~x209;
assign c1549 =  x226 & ~x146 & ~x295 & ~x323;
assign c1551 =  x193 &  x206 & ~x23 & ~x41;
assign c1553 =  x111 & ~x1 & ~x6 & ~x319;
assign c1555 = ~x67 & ~x106 & ~x154;
assign c1557 =  x24 &  x96 &  x101 &  x267 & ~x255;
assign c1559 =  x178 & ~x192 & ~x242 & ~x321;
assign c1561 =  x256 &  x312 & ~x136;
assign c1563 =  x143 & ~x90 & ~x105 & ~x163;
assign c1565 =  x92 &  x128 & ~x225;
assign c1567 =  x258 & ~x228;
assign c1569 =  x60 &  x242 &  x308;
assign c1571 =  x221 & ~x277 & ~x319 & ~x323;
assign c1573 =  x24 &  x197 &  x262 &  x313 & ~x226;
assign c1575 =  x97 &  x124 &  x137 & ~x112;
assign c1577 =  x0 & ~x120;
assign c1579 =  x67 &  x143 &  x157 &  x184 & ~x280;
assign c1581 =  x94 &  x117 &  x133 &  x161 &  x175;
assign c1583 =  x19 & ~x120 & ~x125 & ~x255;
assign c1585 =  x101 &  x121 &  x292 &  x321 & ~x217;
assign c1587 =  x200 & ~x306;
assign c1589 =  x101 &  x150 & ~x183;
assign c1591 =  x77 & ~x232 & ~x291;
assign c1593 =  x20 &  x123 & ~x68 & ~x264;
assign c1595 =  x123 &  x184 &  x256 &  x312;
assign c1597 =  x297 & ~x2 & ~x103 & ~x269;
assign c1599 = ~x18 & ~x105 & ~x131 & ~x154 & ~x265;

endmodule