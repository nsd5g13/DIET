module tm( x0,x1,x2,x3,x4,x5,x6,x7,x8,x9,x10,x11,x12,x13,x14,x15,x16,x17,x18,x19,x20,x21,x22,x23,x24,x25,x26,x27,x28,x29,x30,x31,x32,x33,x34,x35,x36,x37,x38,x39,x40,x41,x42,x43,x44,x45,x46,x47,x48,x49,x50,x51,x52,x53,x54,x55,x56,x57,x58,x59,x60,x61,x62,x63,x64,x65,x66,x67,x68,x69,x70,x71,x72,x73,x74,x75,x76,x77,x78,x79,x80,x81,x82,x83,x84,x85,x86,x87,x88,x89,x90,x91,x92,x93,x94,x95,x96,x97,x98,x99,x100,x101,x102,x103,x104,x105,x106,x107,x108,x109,x110,x111,x112,x113,x114,x115,x116,x117,x118,x119,x120,x121,x122,x123,x124,x125,x126,x127,x128,x129,x130,x131,x132,x133,x134,x135,x136,x137,x138,x139,x140,x141,x142,x143,x144,x145,x146,x147,x148,x149,x150,x151,x152,x153,x154,x155,x156,x157,x158,x159,x160,x161,x162,x163,x164,x165,x166,x167,x168,x169,x170,x171,x172,x173,x174,x175,x176,x177,x178,x179,x180,x181,x182,x183,x184,x185,x186,x187,x188,x189,x190,x191,x192,x193,x194,x195,x196,x197,x198,x199,x200,x201,x202,x203,x204,x205,x206,x207,x208,x209,x210,x211,x212,x213,x214,x215,x216,x217,x218,x219,x220,x221,x222,x223,x224,x225,x226,x227,x228,x229,x230,x231,x232,x233,x234,x235,x236,x237,x238,x239,x240,x241,x242,x243,x244,x245,x246,x247,x248,x249,x250,x251,x252,x253,x254,x255,x256,x257,x258,x259,x260,x261,x262,x263,x264,x265,x266,x267,x268,x269,x270,x271,x272,x273,x274,x275,x276,x277,x278,x279,x280,x281,x282,x283,x284,x285,x286,x287,x288,x289,x290,x291,x292,x293,x294,x295,x296,x297,x298,x299,x300,x301,x302,x303,x304,x305,x306,x307,x308,x309,x310,x311,x312,x313,x314,x315,x316,x317,x318,x319,x320,x321,x322,x323,x324,x325,x326,x327,x328,x329,x330,x331,x332,x333,x334,x335,x336,x337,x338,x339,x340,x341,x342,x343,x344,x345,x346,x347,x348,x349,x350,x351,x352,x353,x354,x355,x356,x357,x358,x359,x360,x361,x362,x363,x364,x365,x366,x367,x368,x369,x370,x371,x372,x373,x374,x375,x376,x377,x378,x379,x380,x381,x382,x383,x384,x385,x386,x387,x388,x389,x390,x391,x392,x393,x394,x395,x396,x397,x398,x399,x400,x401,x402,x403,x404,x405,x406,x407,x408,x409,x410,x411,x412,x413,x414,x415,x416,x417,x418,x419,x420,x421,x422,x423,x424,x425,x426,x427,x428,x429,x430,x431,x432,x433,x434,x435,x436,x437,x438,x439,x440,x441,x442,x443,x444,x445,x446,x447,x448,x449,x450,x451,x452,x453,x454,x455,x456,x457,x458,x459,x460,x461,x462,x463,x464,x465,x466,x467,x468,x469,x470,x471,x472,x473,x474,x475,x476,x477,x478,x479,x480,x481,x482,x483,x484,x485,x486,x487,x488,x489,x490,x491,x492,x493,x494,x495,x496,x497,x498,x499,x500,x501,x502,x503,x504,x505,x506,x507,x508,x509,x510,x511,x512,x513,x514,x515,x516,x517,x518,x519,x520,x521,x522,x523,x524,x525,x526,x527,x528,x529,x530,x531,x532,x533,x534,x535,x536,x537,x538,x539,x540,x541,x542,x543,x544,x545,x546,x547,x548,x549,x550,x551,x552,x553,x554,x555,x556,x557,x558,x559,x560,x561,x562,x563,x564,x565,x566,x567,x568,x569,x570,x571,x572,x573,x574,x575,x576,x577,x578,x579,x580,x581,x582,x583,x584,x585,x586,x587,x588,x589,x590,x591,x592,x593,x594,x595,x596,x597,x598,x599,x600,x601,x602,x603,x604,x605,x606,x607,x608,x609,x610,x611,x612,x613,x614,x615,x616,x617,x618,x619,x620,x621,x622,x623,x624,x625,x626,x627,x628,x629,x630,x631,x632,x633,x634,x635,x636,x637,x638,x639,x640,x641,x642,x643,x644,x645,x646,x647,x648,x649,x650,x651,x652,x653,x654,x655,x656,x657,x658,x659,x660,x661,x662,x663,x664,x665,x666,x667,x668,x669,x670,x671,x672,x673,x674,x675,x676,x677,x678,x679,x680,x681,x682,x683,x684,x685,x686,x687,x688,x689,x690,x691,x692,x693,x694,x695,x696,x697,x698,x699,x700,x701,x702,x703,x704,x705,x706,x707,x708,x709,x710,x711,x712,x713,x714,x715,x716,x717,x718,x719,x720,x721,x722,x723,x724,x725,x726,x727,x728,x729,x730,x731,x732,x733,x734,x735,x736,x737,x738,x739,x740,x741,x742,x743,x744,x745,x746,x747,x748,x749,x750,x751,x752,x753,x754,x755,x756,x757,x758,x759,x760,x761,x762,x763,x764,x765,x766,x767,x768,x769,x770,x771,x772,x773,x774,x775,x776,x777,x778,x779,x780,x781,x782,x783,x784,x785,x786,x787,x788,x789,x790,x791,x792,x793,x794,x795,x796,x797,x798,x799,x800,x801,x802,x803,x804,x805,x806,x807,x808,x809,x810,x811,x812,x813,x814,x815,x816,x817,x818,x819,x820,x821,x822,x823,x824,x825,x826,x827,x828,x829,x830,x831,x832,x833,x834,x835,x836,x837,x838,x839,x840,x841,x842,x843,x844,x845,x846,x847,x848,x849,x850,x851,x852,x853,x854,x855,x856,x857,x858,x859,x860,x861,x862,x863,x864,x865,x866,x867,x868,x869,x870,x871,x872,x873,x874,x875,x876,x877,x878,x879,x880,x881,x882,x883,x884,x885,x886,x887,x888,x889,x890,x891,x892,x893,x894,x895,x896,x897,x898,x899,x900,x901,x902,x903,x904,x905,x906,x907,x908,x909,x910,x911,x912,x913,x914,x915,x916,x917,x918,x919,x920,x921,x922,x923,x924,x925,x926,x927,x928,x929,x930,x931,x932,x933,x934,x935,x936,x937,x938,x939,x940,x941,x942,x943,x944,x945,x946,x947,x948,x949,x950,x951,x952,x953,x954,x955,x956,x957,x958,x959,x960,x961,x962,x963,x964,x965,x966,x967,x968,x969,x970,x971,x972,x973,x974,x975,x976,x977,x978,x979,x980,x981,x982,x983,x984,x985,x986,x987,x988,x989,x990,x991,x992,x993,x994,x995,x996,x997,x998,x999,x1000,x1001,x1002,x1003,x1004,x1005,x1006,x1007,x1008,x1009,x1010,x1011,x1012,x1013,x1014,x1015,x1016,x1017,x1018,x1019,x1020,x1021,x1022,x1023,x1024,x1025,x1026,x1027,x1028,x1029,x1030,x1031,x1032,x1033,x1034,x1035,x1036,x1037,x1038,x1039,x1040,x1041,x1042,x1043,x1044,x1045,x1046,x1047,x1048,x1049,x1050,x1051,x1052,x1053,x1054,x1055,x1056,x1057,x1058,x1059,x1060,x1061,x1062,x1063,x1064,x1065,x1066,x1067,x1068,x1069,x1070,x1071,x1072,x1073,x1074,x1075,x1076,x1077,x1078,x1079,x1080,x1081,x1082,x1083,x1084,x1085,x1086,x1087,x1088,x1089,x1090,x1091,x1092,x1093,x1094,x1095,x1096,x1097,x1098,x1099,x1100,x1101,x1102,x1103,x1104,x1105,x1106,x1107,x1108,x1109,x1110,x1111,x1112,x1113,x1114,x1115,x1116,x1117,x1118,x1119,x1120,x1121,x1122,x1123,x1124,x1125,x1126,x1127,x1128,x1129,x1130,c4223,c036,c259,c5176,c6274,c7287,c2295,c732,c7122,c6221,c524,c121,c3237,c1212,c6217,c6159,c6190,c6143,c3223,c3110,c3293,c3236,c568,c3221,c2118,c06,c2270,c334,c261,c183,c7160,c6230,c6175,c1155,c4294,c5168,c4253,c3143,c1226,c5228,c1175,c451,c579,c236,c7289,c1194,c6151,c562,c6145,c6268,c493,c2228,c3204,c748,c4229,c515,c725,c3139,c7123,c4231,c219,c7267,c292,c65,c1235,c3252,c46,c1243,c651,c643,c354,c391,c6192,c3227,c7234,c1197,c31,c4145,c2182,c5130,c20,c5182,c434,c3288,c4122,c689,c636,c38,c6176,c1169,c2112,c1192,c048,c3172,c57,c5274,c5265,c0198,c1151,c1150,c362,c7210,c342,c7180,c211,c1129,c273,c454,c7219,c0207,c3286,c435,c4111,c1154,c2271,c2251,c1128,c5122,c547,c2272,c2107,c4207,c715,c6164,c234,c3262,c4230,c728,c4152,c046,c14,c3180,c347,c2204,c291,c4161,c7213,c6216,c343,c1220,c1113,c2256,c1149,c1255,c340,c1259,c766,c0267,c1114,c527,c060,c156,c3299,c3280,c1180,c4283,c45,c330,c1284,c043,c724,c0182,c2131,c621,c5102,c413,c0295,c0249,c0287,c7217,c358,c685,c3199,c4244,c541,c5224,c74,c2254,c28,c4267,c742,c693,c3174,c798,c1118,c282,c658,c173,c2114,c1158,c1279,c093,c09,c191,c2296,c3222,c367,c5250,c224,c3168,c4259,c611,c091,c37,c7169,c041,c087,c614,c673,c1181,c2242,c5157,c3135,c596,c0129,c1252,c3107,c5292,c4139,c0128,c6113,c0167,c366,c115,c491,c126,c084,c016,c7233,c1270,c755,c4212,c1146,c2117,c3260,c460,c086,c1251,c761,c7268,c6207,c2142,c3212,c1139,c7155,c7145,c3244,c6122,c269,c610,c7256,c0245,c539,c0166,c736,c5222,c258,c3178,c7105,c0291,c2249,c6119,c6285,c4171,c4128,c5237,c0140,c373,c2132,c6165,c034,c1272,c230,c625,c0272,c6102,c6129,c387,c238,c3238,c3219,c3185,c0105,c6171,c180,c3287,c7247,c3165,c0268,c08,c2241,c7276,c6189,c3157,c511,c299,c556,c7258,c25,c07,c780,c3251,c2115,c0229,c7154,c2105,c627,c52,c757,c4188,c395,c7202,c586,c426,c0168,c5143,c7159,c1227,c361,c1229,c0223,c6117,c5106,c370,c6225,c075,c6224,c247,c3106,c4125,c1201,c744,c239,c5132,c061,c64,c2195,c331,c1241,c0113,c228,c381,c7198,c2169,c4189,c711,c768,c735,c733,c4241,c05,c1120,c6266,c30,c1132,c3208,c7193,c5271,c067,c758,c140,c3184,c223,c3283,c545,c297,c1157,c4184,c16,c5159,c1167,c3217,c6148,c3131,c0282,c3101,c044,c333,c3183,c058,c4187,c6173,c443,c2176,c339,c4272,c0145,c2202,c1224,c3133,c6283,c740,c7115,c59,c216,c0114,c2172,c2200,c438,c4146,c4239,c195,c2261,c6211,c0241,c4154,c4247,c5218,c459,c4287,c324,c773,c0220,c6105,c722,c452,c6229,c525,c4180,c0102,c376,c6142,c0211,c6179,c10,c0205,c2144,c4248,c543,c519,c335,c1287,c1119,c5287,c0165,c1292,c3259,c792,c1190,c7146,c7241,c3104,c1123,c235,c187,c233,c5110,c5154,c531,c6130,c6238,c6128,c229,c36,c348,c731,c4198,c271,c3194,c3250,c430,c7152,c559,c6218,c1230,c63,c5111,c769,c799,c01,c7149,c2275,c752,c389,c7111,c420,c015,c251,c2273,c4130,c791,c578,c7244,c172,c013,c4269,c589,c380,c0219,c1237,c2122,c517,c222,c497,c244,c7295,c7165,c2247,c053,c7163,c011,c5249,c622,c2159,c4124,c4101,c631,c1168,c499,c7172,c145,c4140,c1256,c4222,c364,c17,c7191,c3277,c794,c3254,c5108,c1248,c5262,c7230,c660,c5298,c0226,c2227,c6166,c316,c3121,c2234,c727,c2133,c0225,c1278,c558,c552,c5170,c116,c3214,c4160,c2152,c3140,c49,c020,c494,c6125,c7109,c617,c7255,c0202,c337,c6153,c582,c71,c112,c6296,c55,c7288,c496,c1176,c7179,c4276,c274,c2179,c7299,c0298,c0164,c5236,c669,c2281,c135,c4183,c3270,c667,c5116,c18,c3122,c3176,c117,c7224,c0254,c5136,c4127,c2192,c686,c154,c7117,c0273,c398,c2146,c1193,c6249,c0175,c597,c577,c1156,c6144,c6279,c7157,c0159,c2217,c5261,c536,c226,c6198,c1208,c3102,c3203,c394,c764,c1174,c5276,c215,c7283,c4118,c2189,c0119,c696,c6136,c77,c2214,c2259,c593,c240,c464,c444,c6127,c7185,c6202,c3173,c1210,c2237,c485,c5266,c1105,c2130,c648,c6290,c796,c1211,c7278,c5134,c119,c0177,c5121,c467,c045,c7134,c159,c4255,c3189,c13,c5181,c070,c083,c0253,c4273,c4245,c4205,c2160,c6186,c7296,c139,c0185,c5260,c4115,c2292,c4268,c6108,c4119,c7226,c7206,c3170,c638,c388,c6265,c7168,c4210,c128,c137,c7297,c166,c072,c3228,c0151,c698,c0265,c138,c2139,c0237,c6258,c056,c789,c7221,c0111,c0277,c6185,c5221,c3215,c3220,c5296,c294,c0172,c410,c377,c415,c0122,c637,c3161,c4256,c1126,c160,c1280,c7102,c39,c2119,c1276,c095,c2252,c3231,c047,c1178,c1117,c3258,c3150,c0250,c0127,c136,c583,c3278,c04,c2231,c5238,c7238,c5171,c6293,c0150,c4217,c288,c7199,c1133,c462,c5187,c263,c7266,c2149,c6152,c793,c3247,c7107,c078,c421,c784,c633,c476,c4208,c7232,c7120,c6204,c385,c6182,c349,c129,c141,c4275,c245,c19,c153,c2226,c6246,c0153,c3242,c040,c3253,c22,c528,c6226,c2137,c487,c599,c2167,c5280,c0269,c6231,c1161,c50,c360,c3144,c017,c668,c619,c418,c481,c4165,c3290,c0137,c0108,c114,c4144,c6257,c6219,c72,c032,c0278,c6169,c7161,c4129,c2175,c7133,c296,c7194,c537,c063,c6112,c2294,c1218,c019,c5259,c4258,c049,c7162,c3226,c255,c346,c2253,c2267,c2246,c0124,c4131,c7187,c429,c155,c1131,c374,c2243,c2255,c0209,c58,c6104,c783,c386,c1148,c6247,c7188,c7269,c1253,c530,c2290,c1205,c5207,c2165,c4143,c6264,c0144,c6299,c3274,c1294,c774,c2224,c2180,c629,c4233,c4176,c1203,c7239,c442,c1187,c4249,c523,c592,c664,c5196,c0138,c0215,c7174,c5144,c518,c495,c2282,c2109,c1107,c351,c6100,c2138,c5160,c029,c0125,c220,c3147,c4148,c461,c130,c6157,c1185,c4279,c7127,c094,c4116,c5210,c0297,c7261,c591,c7119,c5138,c2245,c7290,c074,c7147,c4297,c721,c5215,c146,c6263,c2170,c1234,c218,c4274,c3148,c133,c0244,c6103,c1247,c7197,c3191,c148,c051,c3273,c0169,c2197,c3196,c6292,c6245,c2262,c620,c1225,c1166,c039,c4179,c672,c720,c2264,c4224,c532,c439,c131,c2126,c2268,c0294,c73,c692,c2235,c7139,c165,c2106,c0188,c2229,c110,c486,c474,c7257,c7121,c0240,c3190,c32,c6286,c174,c5120,c2277,c1274,c6297,c1290,c375,c7189,c569,c699,c557,c4290,c2129,c7207,c5251,c0246,c134,c6281,c7177,c2174,c397,c5139,c7216,c2293,c513,c2258,c5284,c5267,c3298,c3100,c4270,c1196,c4175,c428,c6294,c763,c3153,c281,c795,c1182,c6270,c69,c62,c797,c2248,c3292,c080,c0197,c3234,c4200,c1165,c2154,c535,c6201,c7277,c7282,c449,c089,c5185,c5186,c0196,c5203,c5257,c7274,c2164,c3145,c650,c1124,c3279,c34,c6250,c225,c563,c5225,c4246,c2121,c5165,c6200,c7280,c0262,c653,c623,c0115,c2212,c055,c6170,c4214,c5279,c5193,c5232,c7271,c7141,c4254,c5105,c0275,c332,c1122,c5202,c7132,c5149,c3243,c2211,c1141,c0109,c284,c2265,c0280,c5263,c6256,c0149,c0195,c5169,c5178,c5208,c188,c0285,c0116,c2153,c5180,c2143,c1296,c190,c5252,c5288,c2110,c27,c670,c6140,c785,c53,c5270,c5275,c5283,c012,c498,c1268,c7273,c6213,c417,c3188,c4138,c6203,c489,c5201,c6121,c7170,c5184,c1159,c383,c3197,c3108,c7279,c6237,c4238,c5214,c695,c2209,c540,c2171,c1202,c3235,c5268,c176,c1153,c4102,c688,c2299,c1223,c1102,c6120,c782,c170,c393,c483,c7292,c5239,c729,c5285,c3245,c250,c70,c6168,c412,c7135,c3138,c448,c6239,c1145,c5217,c3115,c4163,c1217,c161,c1179,c6187,c4134,c6195,c042,c6260,c7130,c2113,c5254,c7281,c550,c030,c754,c2238,c588,c6163,c778,c416,c0251,c432,c210,c0271,c575,c1222,c475,c2222,c321,c5189,c29,c3136,c3255,c4192,c7298,c6253,c1143,c7228,c3213,c5241,c6199,c6244,c4213,c1104,c546,c0157,c2260,c7144,c4281,c5195,c7240,c635,c2280,c3141,c3256,c4227,c3120,c565,c697,c5167,c062,c4169,c746,c252,c1171,c1195,c4237,c2279,c7200,c1233,c5290,c5204,c5226,c7246,c0184,c0118,c520,c7104,c2166,c1281,c6271,c02,c123,c2285,c2297,c7209,c2184,c639,c0224,c587,c5192,c2136,c1127,c4215,c5246,c776,c3128,c7136,c2155,c4177,c4156,c4167,c712,c3186,c427,c6240,c456,c314,c1232,c0112,c573,c6251,c0187,c265,c311,c2128,c379,c3294,c327,c6232,c4186,c064,c477,c7229,c2188,c0243,c2123,c4150,c1213,c414,c618,c0228,c4206,c6156,c382,c6254,c7176,c4137,c2135,c4257,c7138,c0186,c553,c1136,c694,c4288,c4159,c647,c6298,c2150,c0216,c0106,c192,c661,c167,c6233,c510,c318,c290,c7190,c5247,c4166,c2177,c079,c671,c4242,c7103,c5103,c4295,c2116,c6126,c750,c642,c248,c2147,c268,c359,c576,c5163,c4196,c4221,c458,c7285,c471,c232,c4293,c5293,c3285,c1130,c4181,c4142,c7291,c4266,c026,c242,c3296,c378,c169,c4172,c4278,c1228,c280,c3109,c3132,c6272,c162,c7203,c3123,c071,c488,c3114,c0270,c1289,c734,c221,c4298,c3232,c312,c2210,c2266,c1231,c6131,c4232,c3265,c3224,c7126,c3207,c2289,c0206,c1221,c7215,c295,c788,c1188,c512,c615,c6158,c7231,c2225,c352,c1109,c6178,c1101,c6269,c021,c7259,c612,c6223,c3162,c6278,c1298,c4263,c5199,c0201,c189,c730,c326,c317,c2199,c0258,c2168,c4225,c1291,c0173,c1263,c3111,c0141,c613,c027,c2274,c469,c5240,c150,c538,c7286,c2286,c7183,c5198,c0264,c7118,c771,c6288,c7129,c2104,c099,c2257,c3264,c7275,c2162,c594,c4164,c54,c344,c645,c665,c1200,c433,c3239,c5151,c760,c0135,c315,c7237,c470,c0193,c1238,c6191,c7181,c262,c1286,c0217,c595,c3156,c7214,c4228,c2127,c6261,c185,c254,c683,c0248,c025,c177,c5146,c097,c5125,c7164,c7114,c4178,c1283,c0163,c777,c7227,c4282,c7128,c678,c5200,c3182,c7218,c5118,c164,c186,c5156,c4240,c33,c472,c6295,c6101,c122,c6115,c7220,c4286,c659,c2151,c2218,c5291,c4277,c0279,c5223,c492,c6255,c463,c6174,c677,c7245,c3158,c329,c2156,c544,c7251,c270,c1273,c5227,c7125,c264,c1257,c0231,c212,c285,c522,c7250,c152,c466,c142,c2206,c5256,c3218,c0233,c6114,c717,c0132,c6222,c6181,c6193,c473,c253,c666,c4123,c199,c42,c431,c3275,c4147,c266,c2148,c634,c5115,c5161,c5183,c3261,c446,c0218,c1198,c057,c120,c1277,c2158,c1254,c0227,c5155,c3202,c1269,c5114,c2120,c616,c480,c751,c5128,c0208,c6227,c3152,c6277,c6141,c7264,c163,c368,c0221,c6262,c0286,c786,c7153,c175,c4201,c4105,c213,c5277,c1103,c350,c2185,c1135,c775,c0255,c4104,c7112,c1116,c7222,c3198,c0257,c6154,c490,c082,c3263,c5175,c5101,c090,c2239,c0276,c2276,c7196,c5206,c6106,c1138,c023,c0232,c256,c3151,c014,c3103,c3230,c1170,c2232,c7260,c035,c1293,c5295,c5142,c4170,c5243,c5177,c5233,c3205,c356,c3126,c7236,c4168,c4121,c2198,c2134,c118,c0117,c4284,c0110,c4292,c5123,c5153,c0296,c719,c6177,c548,c5299,c5145,c293,c0101,c1189,c1282,c3257,c4199,c0107,c7272,c3209,c4218,c4203,c1297,c392,c2250,c038,c2220,c4110,c4193,c79,c15,c319,c0142,c4264,c0242,c037,c2230,c4252,c0100,c726,c184,c4173,c6282,c716,c6111,c43,c4195,c2205,c033,c4296,c0180,c0103,c031,c298,c5190,c3267,c365,c424,c384,c3266,c2125,c3175,c5230,c6243,c3179,c691,c390,c6196,c7108,c5133,c5137,c2288,c5219,c762,c7212,c178,c0214,c632,c1160,c6167,c179,c534,c5135,c0123,c555,c5117,c147,c2244,c6150,c790,c7171,c0247,c440,c2194,c5281,c714,c363,c0147,c4133,c3268,c1246,c5119,c572,c143,c40,c4243,c3159,c6228,c1216,c749,c3113,c0288,c743,c3124,c024,c6110,c125,c5179,c7116,c287,c5245,c574,c2141,c2183,c0261,c5297,c0156,c567,c1264,c0133,c0210,c23,c7110,c484,c7182,c4220,c6214,c628,c4155,c151,c468,c0281,c0139,c441,c24,c5131,c144,c772,c1260,c56,c4113,c1236,c5209,c3164,c1295,c3246,c447,c7284,c4235,c7151,c2216,c2223,c2284,c2157,c7253,c0200,c2193,c3160,c5166,c0176,c4158,c6291,c521,c5191,c6135,c5152,c310,c3166,c479,c6160,c6116,c3241,c584,c1242,c3210,c4162,c6284,c4109,c5212,c3192,c2173,c0120,c4174,c2196,c371,c0238,c5188,c5205,c2186,c66,c4285,c3193,c756,c241,c425,c78,c2102,c739,c6259,c3289,c0259,c7167,c7294,c214,c0178,c4141,c0121,c6133,c052,c0204,c6220,c5269,c2291,c5216,c7166,c7223,c372,c7186,c5150,c4153,c453,c4261,c7270,c0174,c2208,c077,c069,c1110,c3169,c6180,c322,c345,c277,c6212,c590,c7265,c4236,c3125,c6194,c5289,c4209,c0152,c0148,c652,c747,c5172,c0235,c2145,c3167,c581,c6172,c3134,c3142,c2207,c4100,c0283,c3195,c1240,c1258,c4132,c0256,c2201,c237,c1207,c181,c243,c4216,c1266,c2181,c3248,c570,c5235,c7175,c423,c437,c1267,c158,c7225,c5158,c323,c1245,c276,c529,c3282,c6236,c246,c2263,c564,c687,c640,c336,c3118,c3225,c4191,c4106,c092,c0234,c4114,c081,c193,c1288,c113,c0289,c3201,c0260,c6134,c0130,c6162,c6188,c1164,c00,c1214,c624,c6209,c1108,c0155,c0299,c3249,c2108,c6276,c765,c283,c7173,c1261,c5147,c1206,c4149,c0192,c1299,c560,c066,c1209,c2111,c5282,c0213,c580,c436,c6183,c679,c2203,c085,c111,c5258,c630,c2298,c4103,c7124,c566,c6248,c1147,c60,c194,c551,c5129,c585,c1191,c289,c6289,c4299,c3211,c1112,c4234,c4190,c010,c561,c6161,c132,c171,c0158,c48,c5211,c738,c278,c1204,c684,c0230,c1106,c3146,c6287,c018,c355,c227,c5294,c279,c51,c149,c1100,c1177,c76,c4262,c272,c0274,c182,c656,c4211,c61,c7184,c124,c4108,c5272,c5278,c2103,c0162,c674,c157,c3187,c770,c2140,c5174,c325,c655,c4151,c068,c571,c6215,c198,c21,c680,c0212,c710,c2215,c6107,c682,c0181,c7192,c0203,c663,c6273,c0179,c2161,c3149,c2283,c7293,c6210,c6118,c088,c5124,c028,c450,c059,c3181,c7243,c7106,c7142,c7195,c0190,c7254,c4251,c1219,c4226,c787,c1137,c6235,c5104,c073,c2269,c1239,c767,c0292,c3127,c6280,c723,c197,c759,c6123,c3155,c641,c0160,c1275,c2219,c4120,c050,c0236,c3171,c196,c7208,c0134,c1186,c0136,c3163,c2278,c0126,c6139,c3117,c4126,c5141,c4280,c4265,c5248,c3233,c6252,c6234,c3112,c2191,c4135,c1250,c3137,c2213,c741,c5231,c7178,c12,c5197,c353,c7100,c6197,c0171,c7143,c526,c399,c0194,c516,c781,c022,c4289,c7248,c737,c455,c2178,c076,c338,c7137,c369,c1121,c0183,c396,c1244,c4204,c6147,c549,c7204,c1134,c5244,c3177,c1152,c1249,c260,c411,c5112,c2124,c0239,c6275,c0154,c1183,c1262,c67,c646,c422,c626,c0263,c554,c0104,c0199,c168,c7205,c249,c065,c41,c2240,c257,c5253,c7211,c745,c3105,c0252,c4117,c096,c7235,c6109,c313,c5107,c6184,c44,c6149,c644,c7113,c3216,c217,c4202,c5234,c7140,c1184,c7263,c482,c5220,c5113,c2236,c7156,c098,c2101,c4107,c5140,c127,c3276,c5162,c4197,c1142,c35,c6132,c328,c3206,c5242,c0146,c1140,c1162,c7249,c657,c1265,c26,c598,c5164,c662,c690,c2233,c4219,c0161,c7262,c5229,c1199,c7158,c2221,c3295,c1285,c341,c6138,c4260,c478,c0189,c6267,c0222,c1172,c3200,c2287,c6208,c1144,c675,c6124,c5100,c75,c1215,c654,c3284,c676,c7252,c5264,c0293,c3281,c5126,c4182,c275,c0143,c5194,c357,c3119,c1163,c2187,c4271,c4136,c47,c5273,c718,c5255,c7150,c1111,c7242,c457,c514,c753,c11,c649,c6205,c267,c7101,c465,c1125,c2190,c3229,c4112,c6155,c286,c4194,c779,c3271,c3130,c6206,c6241,c7201,c7148,c5148,c6242,c713,c4291,c5173,c3240,c445,c0284,c1271,c4185,c320,c3154,c3291,c2163,c533,c5127,c68,c3297,c7131,c1173,c681,c542,c5286,c3272,c5109,c1115,c6137,c054,c0131,c3116,c0266,c0170,c3269,c2100,c0290,c0191,c4250,c3129,c419,c6146,c4157,c231,c03,c5213 );

input x0;
input x1;
input x2;
input x3;
input x4;
input x5;
input x6;
input x7;
input x8;
input x9;
input x10;
input x11;
input x12;
input x13;
input x14;
input x15;
input x16;
input x17;
input x18;
input x19;
input x20;
input x21;
input x22;
input x23;
input x24;
input x25;
input x26;
input x27;
input x28;
input x29;
input x30;
input x31;
input x32;
input x33;
input x34;
input x35;
input x36;
input x37;
input x38;
input x39;
input x40;
input x41;
input x42;
input x43;
input x44;
input x45;
input x46;
input x47;
input x48;
input x49;
input x50;
input x51;
input x52;
input x53;
input x54;
input x55;
input x56;
input x57;
input x58;
input x59;
input x60;
input x61;
input x62;
input x63;
input x64;
input x65;
input x66;
input x67;
input x68;
input x69;
input x70;
input x71;
input x72;
input x73;
input x74;
input x75;
input x76;
input x77;
input x78;
input x79;
input x80;
input x81;
input x82;
input x83;
input x84;
input x85;
input x86;
input x87;
input x88;
input x89;
input x90;
input x91;
input x92;
input x93;
input x94;
input x95;
input x96;
input x97;
input x98;
input x99;
input x100;
input x101;
input x102;
input x103;
input x104;
input x105;
input x106;
input x107;
input x108;
input x109;
input x110;
input x111;
input x112;
input x113;
input x114;
input x115;
input x116;
input x117;
input x118;
input x119;
input x120;
input x121;
input x122;
input x123;
input x124;
input x125;
input x126;
input x127;
input x128;
input x129;
input x130;
input x131;
input x132;
input x133;
input x134;
input x135;
input x136;
input x137;
input x138;
input x139;
input x140;
input x141;
input x142;
input x143;
input x144;
input x145;
input x146;
input x147;
input x148;
input x149;
input x150;
input x151;
input x152;
input x153;
input x154;
input x155;
input x156;
input x157;
input x158;
input x159;
input x160;
input x161;
input x162;
input x163;
input x164;
input x165;
input x166;
input x167;
input x168;
input x169;
input x170;
input x171;
input x172;
input x173;
input x174;
input x175;
input x176;
input x177;
input x178;
input x179;
input x180;
input x181;
input x182;
input x183;
input x184;
input x185;
input x186;
input x187;
input x188;
input x189;
input x190;
input x191;
input x192;
input x193;
input x194;
input x195;
input x196;
input x197;
input x198;
input x199;
input x200;
input x201;
input x202;
input x203;
input x204;
input x205;
input x206;
input x207;
input x208;
input x209;
input x210;
input x211;
input x212;
input x213;
input x214;
input x215;
input x216;
input x217;
input x218;
input x219;
input x220;
input x221;
input x222;
input x223;
input x224;
input x225;
input x226;
input x227;
input x228;
input x229;
input x230;
input x231;
input x232;
input x233;
input x234;
input x235;
input x236;
input x237;
input x238;
input x239;
input x240;
input x241;
input x242;
input x243;
input x244;
input x245;
input x246;
input x247;
input x248;
input x249;
input x250;
input x251;
input x252;
input x253;
input x254;
input x255;
input x256;
input x257;
input x258;
input x259;
input x260;
input x261;
input x262;
input x263;
input x264;
input x265;
input x266;
input x267;
input x268;
input x269;
input x270;
input x271;
input x272;
input x273;
input x274;
input x275;
input x276;
input x277;
input x278;
input x279;
input x280;
input x281;
input x282;
input x283;
input x284;
input x285;
input x286;
input x287;
input x288;
input x289;
input x290;
input x291;
input x292;
input x293;
input x294;
input x295;
input x296;
input x297;
input x298;
input x299;
input x300;
input x301;
input x302;
input x303;
input x304;
input x305;
input x306;
input x307;
input x308;
input x309;
input x310;
input x311;
input x312;
input x313;
input x314;
input x315;
input x316;
input x317;
input x318;
input x319;
input x320;
input x321;
input x322;
input x323;
input x324;
input x325;
input x326;
input x327;
input x328;
input x329;
input x330;
input x331;
input x332;
input x333;
input x334;
input x335;
input x336;
input x337;
input x338;
input x339;
input x340;
input x341;
input x342;
input x343;
input x344;
input x345;
input x346;
input x347;
input x348;
input x349;
input x350;
input x351;
input x352;
input x353;
input x354;
input x355;
input x356;
input x357;
input x358;
input x359;
input x360;
input x361;
input x362;
input x363;
input x364;
input x365;
input x366;
input x367;
input x368;
input x369;
input x370;
input x371;
input x372;
input x373;
input x374;
input x375;
input x376;
input x377;
input x378;
input x379;
input x380;
input x381;
input x382;
input x383;
input x384;
input x385;
input x386;
input x387;
input x388;
input x389;
input x390;
input x391;
input x392;
input x393;
input x394;
input x395;
input x396;
input x397;
input x398;
input x399;
input x400;
input x401;
input x402;
input x403;
input x404;
input x405;
input x406;
input x407;
input x408;
input x409;
input x410;
input x411;
input x412;
input x413;
input x414;
input x415;
input x416;
input x417;
input x418;
input x419;
input x420;
input x421;
input x422;
input x423;
input x424;
input x425;
input x426;
input x427;
input x428;
input x429;
input x430;
input x431;
input x432;
input x433;
input x434;
input x435;
input x436;
input x437;
input x438;
input x439;
input x440;
input x441;
input x442;
input x443;
input x444;
input x445;
input x446;
input x447;
input x448;
input x449;
input x450;
input x451;
input x452;
input x453;
input x454;
input x455;
input x456;
input x457;
input x458;
input x459;
input x460;
input x461;
input x462;
input x463;
input x464;
input x465;
input x466;
input x467;
input x468;
input x469;
input x470;
input x471;
input x472;
input x473;
input x474;
input x475;
input x476;
input x477;
input x478;
input x479;
input x480;
input x481;
input x482;
input x483;
input x484;
input x485;
input x486;
input x487;
input x488;
input x489;
input x490;
input x491;
input x492;
input x493;
input x494;
input x495;
input x496;
input x497;
input x498;
input x499;
input x500;
input x501;
input x502;
input x503;
input x504;
input x505;
input x506;
input x507;
input x508;
input x509;
input x510;
input x511;
input x512;
input x513;
input x514;
input x515;
input x516;
input x517;
input x518;
input x519;
input x520;
input x521;
input x522;
input x523;
input x524;
input x525;
input x526;
input x527;
input x528;
input x529;
input x530;
input x531;
input x532;
input x533;
input x534;
input x535;
input x536;
input x537;
input x538;
input x539;
input x540;
input x541;
input x542;
input x543;
input x544;
input x545;
input x546;
input x547;
input x548;
input x549;
input x550;
input x551;
input x552;
input x553;
input x554;
input x555;
input x556;
input x557;
input x558;
input x559;
input x560;
input x561;
input x562;
input x563;
input x564;
input x565;
input x566;
input x567;
input x568;
input x569;
input x570;
input x571;
input x572;
input x573;
input x574;
input x575;
input x576;
input x577;
input x578;
input x579;
input x580;
input x581;
input x582;
input x583;
input x584;
input x585;
input x586;
input x587;
input x588;
input x589;
input x590;
input x591;
input x592;
input x593;
input x594;
input x595;
input x596;
input x597;
input x598;
input x599;
input x600;
input x601;
input x602;
input x603;
input x604;
input x605;
input x606;
input x607;
input x608;
input x609;
input x610;
input x611;
input x612;
input x613;
input x614;
input x615;
input x616;
input x617;
input x618;
input x619;
input x620;
input x621;
input x622;
input x623;
input x624;
input x625;
input x626;
input x627;
input x628;
input x629;
input x630;
input x631;
input x632;
input x633;
input x634;
input x635;
input x636;
input x637;
input x638;
input x639;
input x640;
input x641;
input x642;
input x643;
input x644;
input x645;
input x646;
input x647;
input x648;
input x649;
input x650;
input x651;
input x652;
input x653;
input x654;
input x655;
input x656;
input x657;
input x658;
input x659;
input x660;
input x661;
input x662;
input x663;
input x664;
input x665;
input x666;
input x667;
input x668;
input x669;
input x670;
input x671;
input x672;
input x673;
input x674;
input x675;
input x676;
input x677;
input x678;
input x679;
input x680;
input x681;
input x682;
input x683;
input x684;
input x685;
input x686;
input x687;
input x688;
input x689;
input x690;
input x691;
input x692;
input x693;
input x694;
input x695;
input x696;
input x697;
input x698;
input x699;
input x700;
input x701;
input x702;
input x703;
input x704;
input x705;
input x706;
input x707;
input x708;
input x709;
input x710;
input x711;
input x712;
input x713;
input x714;
input x715;
input x716;
input x717;
input x718;
input x719;
input x720;
input x721;
input x722;
input x723;
input x724;
input x725;
input x726;
input x727;
input x728;
input x729;
input x730;
input x731;
input x732;
input x733;
input x734;
input x735;
input x736;
input x737;
input x738;
input x739;
input x740;
input x741;
input x742;
input x743;
input x744;
input x745;
input x746;
input x747;
input x748;
input x749;
input x750;
input x751;
input x752;
input x753;
input x754;
input x755;
input x756;
input x757;
input x758;
input x759;
input x760;
input x761;
input x762;
input x763;
input x764;
input x765;
input x766;
input x767;
input x768;
input x769;
input x770;
input x771;
input x772;
input x773;
input x774;
input x775;
input x776;
input x777;
input x778;
input x779;
input x780;
input x781;
input x782;
input x783;
input x784;
input x785;
input x786;
input x787;
input x788;
input x789;
input x790;
input x791;
input x792;
input x793;
input x794;
input x795;
input x796;
input x797;
input x798;
input x799;
input x800;
input x801;
input x802;
input x803;
input x804;
input x805;
input x806;
input x807;
input x808;
input x809;
input x810;
input x811;
input x812;
input x813;
input x814;
input x815;
input x816;
input x817;
input x818;
input x819;
input x820;
input x821;
input x822;
input x823;
input x824;
input x825;
input x826;
input x827;
input x828;
input x829;
input x830;
input x831;
input x832;
input x833;
input x834;
input x835;
input x836;
input x837;
input x838;
input x839;
input x840;
input x841;
input x842;
input x843;
input x844;
input x845;
input x846;
input x847;
input x848;
input x849;
input x850;
input x851;
input x852;
input x853;
input x854;
input x855;
input x856;
input x857;
input x858;
input x859;
input x860;
input x861;
input x862;
input x863;
input x864;
input x865;
input x866;
input x867;
input x868;
input x869;
input x870;
input x871;
input x872;
input x873;
input x874;
input x875;
input x876;
input x877;
input x878;
input x879;
input x880;
input x881;
input x882;
input x883;
input x884;
input x885;
input x886;
input x887;
input x888;
input x889;
input x890;
input x891;
input x892;
input x893;
input x894;
input x895;
input x896;
input x897;
input x898;
input x899;
input x900;
input x901;
input x902;
input x903;
input x904;
input x905;
input x906;
input x907;
input x908;
input x909;
input x910;
input x911;
input x912;
input x913;
input x914;
input x915;
input x916;
input x917;
input x918;
input x919;
input x920;
input x921;
input x922;
input x923;
input x924;
input x925;
input x926;
input x927;
input x928;
input x929;
input x930;
input x931;
input x932;
input x933;
input x934;
input x935;
input x936;
input x937;
input x938;
input x939;
input x940;
input x941;
input x942;
input x943;
input x944;
input x945;
input x946;
input x947;
input x948;
input x949;
input x950;
input x951;
input x952;
input x953;
input x954;
input x955;
input x956;
input x957;
input x958;
input x959;
input x960;
input x961;
input x962;
input x963;
input x964;
input x965;
input x966;
input x967;
input x968;
input x969;
input x970;
input x971;
input x972;
input x973;
input x974;
input x975;
input x976;
input x977;
input x978;
input x979;
input x980;
input x981;
input x982;
input x983;
input x984;
input x985;
input x986;
input x987;
input x988;
input x989;
input x990;
input x991;
input x992;
input x993;
input x994;
input x995;
input x996;
input x997;
input x998;
input x999;
input x1000;
input x1001;
input x1002;
input x1003;
input x1004;
input x1005;
input x1006;
input x1007;
input x1008;
input x1009;
input x1010;
input x1011;
input x1012;
input x1013;
input x1014;
input x1015;
input x1016;
input x1017;
input x1018;
input x1019;
input x1020;
input x1021;
input x1022;
input x1023;
input x1024;
input x1025;
input x1026;
input x1027;
input x1028;
input x1029;
input x1030;
input x1031;
input x1032;
input x1033;
input x1034;
input x1035;
input x1036;
input x1037;
input x1038;
input x1039;
input x1040;
input x1041;
input x1042;
input x1043;
input x1044;
input x1045;
input x1046;
input x1047;
input x1048;
input x1049;
input x1050;
input x1051;
input x1052;
input x1053;
input x1054;
input x1055;
input x1056;
input x1057;
input x1058;
input x1059;
input x1060;
input x1061;
input x1062;
input x1063;
input x1064;
input x1065;
input x1066;
input x1067;
input x1068;
input x1069;
input x1070;
input x1071;
input x1072;
input x1073;
input x1074;
input x1075;
input x1076;
input x1077;
input x1078;
input x1079;
input x1080;
input x1081;
input x1082;
input x1083;
input x1084;
input x1085;
input x1086;
input x1087;
input x1088;
input x1089;
input x1090;
input x1091;
input x1092;
input x1093;
input x1094;
input x1095;
input x1096;
input x1097;
input x1098;
input x1099;
input x1100;
input x1101;
input x1102;
input x1103;
input x1104;
input x1105;
input x1106;
input x1107;
input x1108;
input x1109;
input x1110;
input x1111;
input x1112;
input x1113;
input x1114;
input x1115;
input x1116;
input x1117;
input x1118;
input x1119;
input x1120;
input x1121;
input x1122;
input x1123;
input x1124;
input x1125;
input x1126;
input x1127;
input x1128;
input x1129;
input x1130;
output c4223;
output c036;
output c259;
output c5176;
output c6274;
output c7287;
output c2295;
output c732;
output c7122;
output c6221;
output c524;
output c121;
output c3237;
output c1212;
output c6217;
output c6159;
output c6190;
output c6143;
output c3223;
output c3110;
output c3293;
output c3236;
output c568;
output c3221;
output c2118;
output c06;
output c2270;
output c334;
output c261;
output c183;
output c7160;
output c6230;
output c6175;
output c1155;
output c4294;
output c5168;
output c4253;
output c3143;
output c1226;
output c5228;
output c1175;
output c451;
output c579;
output c236;
output c7289;
output c1194;
output c6151;
output c562;
output c6145;
output c6268;
output c493;
output c2228;
output c3204;
output c748;
output c4229;
output c515;
output c725;
output c3139;
output c7123;
output c4231;
output c219;
output c7267;
output c292;
output c65;
output c1235;
output c3252;
output c46;
output c1243;
output c651;
output c643;
output c354;
output c391;
output c6192;
output c3227;
output c7234;
output c1197;
output c31;
output c4145;
output c2182;
output c5130;
output c20;
output c5182;
output c434;
output c3288;
output c4122;
output c689;
output c636;
output c38;
output c6176;
output c1169;
output c2112;
output c1192;
output c048;
output c3172;
output c57;
output c5274;
output c5265;
output c0198;
output c1151;
output c1150;
output c362;
output c7210;
output c342;
output c7180;
output c211;
output c1129;
output c273;
output c454;
output c7219;
output c0207;
output c3286;
output c435;
output c4111;
output c1154;
output c2271;
output c2251;
output c1128;
output c5122;
output c547;
output c2272;
output c2107;
output c4207;
output c715;
output c6164;
output c234;
output c3262;
output c4230;
output c728;
output c4152;
output c046;
output c14;
output c3180;
output c347;
output c2204;
output c291;
output c4161;
output c7213;
output c6216;
output c343;
output c1220;
output c1113;
output c2256;
output c1149;
output c1255;
output c340;
output c1259;
output c766;
output c0267;
output c1114;
output c527;
output c060;
output c156;
output c3299;
output c3280;
output c1180;
output c4283;
output c45;
output c330;
output c1284;
output c043;
output c724;
output c0182;
output c2131;
output c621;
output c5102;
output c413;
output c0295;
output c0249;
output c0287;
output c7217;
output c358;
output c685;
output c3199;
output c4244;
output c541;
output c5224;
output c74;
output c2254;
output c28;
output c4267;
output c742;
output c693;
output c3174;
output c798;
output c1118;
output c282;
output c658;
output c173;
output c2114;
output c1158;
output c1279;
output c093;
output c09;
output c191;
output c2296;
output c3222;
output c367;
output c5250;
output c224;
output c3168;
output c4259;
output c611;
output c091;
output c37;
output c7169;
output c041;
output c087;
output c614;
output c673;
output c1181;
output c2242;
output c5157;
output c3135;
output c596;
output c0129;
output c1252;
output c3107;
output c5292;
output c4139;
output c0128;
output c6113;
output c0167;
output c366;
output c115;
output c491;
output c126;
output c084;
output c016;
output c7233;
output c1270;
output c755;
output c4212;
output c1146;
output c2117;
output c3260;
output c460;
output c086;
output c1251;
output c761;
output c7268;
output c6207;
output c2142;
output c3212;
output c1139;
output c7155;
output c7145;
output c3244;
output c6122;
output c269;
output c610;
output c7256;
output c0245;
output c539;
output c0166;
output c736;
output c5222;
output c258;
output c3178;
output c7105;
output c0291;
output c2249;
output c6119;
output c6285;
output c4171;
output c4128;
output c5237;
output c0140;
output c373;
output c2132;
output c6165;
output c034;
output c1272;
output c230;
output c625;
output c0272;
output c6102;
output c6129;
output c387;
output c238;
output c3238;
output c3219;
output c3185;
output c0105;
output c6171;
output c180;
output c3287;
output c7247;
output c3165;
output c0268;
output c08;
output c2241;
output c7276;
output c6189;
output c3157;
output c511;
output c299;
output c556;
output c7258;
output c25;
output c07;
output c780;
output c3251;
output c2115;
output c0229;
output c7154;
output c2105;
output c627;
output c52;
output c757;
output c4188;
output c395;
output c7202;
output c586;
output c426;
output c0168;
output c5143;
output c7159;
output c1227;
output c361;
output c1229;
output c0223;
output c6117;
output c5106;
output c370;
output c6225;
output c075;
output c6224;
output c247;
output c3106;
output c4125;
output c1201;
output c744;
output c239;
output c5132;
output c061;
output c64;
output c2195;
output c331;
output c1241;
output c0113;
output c228;
output c381;
output c7198;
output c2169;
output c4189;
output c711;
output c768;
output c735;
output c733;
output c4241;
output c05;
output c1120;
output c6266;
output c30;
output c1132;
output c3208;
output c7193;
output c5271;
output c067;
output c758;
output c140;
output c3184;
output c223;
output c3283;
output c545;
output c297;
output c1157;
output c4184;
output c16;
output c5159;
output c1167;
output c3217;
output c6148;
output c3131;
output c0282;
output c3101;
output c044;
output c333;
output c3183;
output c058;
output c4187;
output c6173;
output c443;
output c2176;
output c339;
output c4272;
output c0145;
output c2202;
output c1224;
output c3133;
output c6283;
output c740;
output c7115;
output c59;
output c216;
output c0114;
output c2172;
output c2200;
output c438;
output c4146;
output c4239;
output c195;
output c2261;
output c6211;
output c0241;
output c4154;
output c4247;
output c5218;
output c459;
output c4287;
output c324;
output c773;
output c0220;
output c6105;
output c722;
output c452;
output c6229;
output c525;
output c4180;
output c0102;
output c376;
output c6142;
output c0211;
output c6179;
output c10;
output c0205;
output c2144;
output c4248;
output c543;
output c519;
output c335;
output c1287;
output c1119;
output c5287;
output c0165;
output c1292;
output c3259;
output c792;
output c1190;
output c7146;
output c7241;
output c3104;
output c1123;
output c235;
output c187;
output c233;
output c5110;
output c5154;
output c531;
output c6130;
output c6238;
output c6128;
output c229;
output c36;
output c348;
output c731;
output c4198;
output c271;
output c3194;
output c3250;
output c430;
output c7152;
output c559;
output c6218;
output c1230;
output c63;
output c5111;
output c769;
output c799;
output c01;
output c7149;
output c2275;
output c752;
output c389;
output c7111;
output c420;
output c015;
output c251;
output c2273;
output c4130;
output c791;
output c578;
output c7244;
output c172;
output c013;
output c4269;
output c589;
output c380;
output c0219;
output c1237;
output c2122;
output c517;
output c222;
output c497;
output c244;
output c7295;
output c7165;
output c2247;
output c053;
output c7163;
output c011;
output c5249;
output c622;
output c2159;
output c4124;
output c4101;
output c631;
output c1168;
output c499;
output c7172;
output c145;
output c4140;
output c1256;
output c4222;
output c364;
output c17;
output c7191;
output c3277;
output c794;
output c3254;
output c5108;
output c1248;
output c5262;
output c7230;
output c660;
output c5298;
output c0226;
output c2227;
output c6166;
output c316;
output c3121;
output c2234;
output c727;
output c2133;
output c0225;
output c1278;
output c558;
output c552;
output c5170;
output c116;
output c3214;
output c4160;
output c2152;
output c3140;
output c49;
output c020;
output c494;
output c6125;
output c7109;
output c617;
output c7255;
output c0202;
output c337;
output c6153;
output c582;
output c71;
output c112;
output c6296;
output c55;
output c7288;
output c496;
output c1176;
output c7179;
output c4276;
output c274;
output c2179;
output c7299;
output c0298;
output c0164;
output c5236;
output c669;
output c2281;
output c135;
output c4183;
output c3270;
output c667;
output c5116;
output c18;
output c3122;
output c3176;
output c117;
output c7224;
output c0254;
output c5136;
output c4127;
output c2192;
output c686;
output c154;
output c7117;
output c0273;
output c398;
output c2146;
output c1193;
output c6249;
output c0175;
output c597;
output c577;
output c1156;
output c6144;
output c6279;
output c7157;
output c0159;
output c2217;
output c5261;
output c536;
output c226;
output c6198;
output c1208;
output c3102;
output c3203;
output c394;
output c764;
output c1174;
output c5276;
output c215;
output c7283;
output c4118;
output c2189;
output c0119;
output c696;
output c6136;
output c77;
output c2214;
output c2259;
output c593;
output c240;
output c464;
output c444;
output c6127;
output c7185;
output c6202;
output c3173;
output c1210;
output c2237;
output c485;
output c5266;
output c1105;
output c2130;
output c648;
output c6290;
output c796;
output c1211;
output c7278;
output c5134;
output c119;
output c0177;
output c5121;
output c467;
output c045;
output c7134;
output c159;
output c4255;
output c3189;
output c13;
output c5181;
output c070;
output c083;
output c0253;
output c4273;
output c4245;
output c4205;
output c2160;
output c6186;
output c7296;
output c139;
output c0185;
output c5260;
output c4115;
output c2292;
output c4268;
output c6108;
output c4119;
output c7226;
output c7206;
output c3170;
output c638;
output c388;
output c6265;
output c7168;
output c4210;
output c128;
output c137;
output c7297;
output c166;
output c072;
output c3228;
output c0151;
output c698;
output c0265;
output c138;
output c2139;
output c0237;
output c6258;
output c056;
output c789;
output c7221;
output c0111;
output c0277;
output c6185;
output c5221;
output c3215;
output c3220;
output c5296;
output c294;
output c0172;
output c410;
output c377;
output c415;
output c0122;
output c637;
output c3161;
output c4256;
output c1126;
output c160;
output c1280;
output c7102;
output c39;
output c2119;
output c1276;
output c095;
output c2252;
output c3231;
output c047;
output c1178;
output c1117;
output c3258;
output c3150;
output c0250;
output c0127;
output c136;
output c583;
output c3278;
output c04;
output c2231;
output c5238;
output c7238;
output c5171;
output c6293;
output c0150;
output c4217;
output c288;
output c7199;
output c1133;
output c462;
output c5187;
output c263;
output c7266;
output c2149;
output c6152;
output c793;
output c3247;
output c7107;
output c078;
output c421;
output c784;
output c633;
output c476;
output c4208;
output c7232;
output c7120;
output c6204;
output c385;
output c6182;
output c349;
output c129;
output c141;
output c4275;
output c245;
output c19;
output c153;
output c2226;
output c6246;
output c0153;
output c3242;
output c040;
output c3253;
output c22;
output c528;
output c6226;
output c2137;
output c487;
output c599;
output c2167;
output c5280;
output c0269;
output c6231;
output c1161;
output c50;
output c360;
output c3144;
output c017;
output c668;
output c619;
output c418;
output c481;
output c4165;
output c3290;
output c0137;
output c0108;
output c114;
output c4144;
output c6257;
output c6219;
output c72;
output c032;
output c0278;
output c6169;
output c7161;
output c4129;
output c2175;
output c7133;
output c296;
output c7194;
output c537;
output c063;
output c6112;
output c2294;
output c1218;
output c019;
output c5259;
output c4258;
output c049;
output c7162;
output c3226;
output c255;
output c346;
output c2253;
output c2267;
output c2246;
output c0124;
output c4131;
output c7187;
output c429;
output c155;
output c1131;
output c374;
output c2243;
output c2255;
output c0209;
output c58;
output c6104;
output c783;
output c386;
output c1148;
output c6247;
output c7188;
output c7269;
output c1253;
output c530;
output c2290;
output c1205;
output c5207;
output c2165;
output c4143;
output c6264;
output c0144;
output c6299;
output c3274;
output c1294;
output c774;
output c2224;
output c2180;
output c629;
output c4233;
output c4176;
output c1203;
output c7239;
output c442;
output c1187;
output c4249;
output c523;
output c592;
output c664;
output c5196;
output c0138;
output c0215;
output c7174;
output c5144;
output c518;
output c495;
output c2282;
output c2109;
output c1107;
output c351;
output c6100;
output c2138;
output c5160;
output c029;
output c0125;
output c220;
output c3147;
output c4148;
output c461;
output c130;
output c6157;
output c1185;
output c4279;
output c7127;
output c094;
output c4116;
output c5210;
output c0297;
output c7261;
output c591;
output c7119;
output c5138;
output c2245;
output c7290;
output c074;
output c7147;
output c4297;
output c721;
output c5215;
output c146;
output c6263;
output c2170;
output c1234;
output c218;
output c4274;
output c3148;
output c133;
output c0244;
output c6103;
output c1247;
output c7197;
output c3191;
output c148;
output c051;
output c3273;
output c0169;
output c2197;
output c3196;
output c6292;
output c6245;
output c2262;
output c620;
output c1225;
output c1166;
output c039;
output c4179;
output c672;
output c720;
output c2264;
output c4224;
output c532;
output c439;
output c131;
output c2126;
output c2268;
output c0294;
output c73;
output c692;
output c2235;
output c7139;
output c165;
output c2106;
output c0188;
output c2229;
output c110;
output c486;
output c474;
output c7257;
output c7121;
output c0240;
output c3190;
output c32;
output c6286;
output c174;
output c5120;
output c2277;
output c1274;
output c6297;
output c1290;
output c375;
output c7189;
output c569;
output c699;
output c557;
output c4290;
output c2129;
output c7207;
output c5251;
output c0246;
output c134;
output c6281;
output c7177;
output c2174;
output c397;
output c5139;
output c7216;
output c2293;
output c513;
output c2258;
output c5284;
output c5267;
output c3298;
output c3100;
output c4270;
output c1196;
output c4175;
output c428;
output c6294;
output c763;
output c3153;
output c281;
output c795;
output c1182;
output c6270;
output c69;
output c62;
output c797;
output c2248;
output c3292;
output c080;
output c0197;
output c3234;
output c4200;
output c1165;
output c2154;
output c535;
output c6201;
output c7277;
output c7282;
output c449;
output c089;
output c5185;
output c5186;
output c0196;
output c5203;
output c5257;
output c7274;
output c2164;
output c3145;
output c650;
output c1124;
output c3279;
output c34;
output c6250;
output c225;
output c563;
output c5225;
output c4246;
output c2121;
output c5165;
output c6200;
output c7280;
output c0262;
output c653;
output c623;
output c0115;
output c2212;
output c055;
output c6170;
output c4214;
output c5279;
output c5193;
output c5232;
output c7271;
output c7141;
output c4254;
output c5105;
output c0275;
output c332;
output c1122;
output c5202;
output c7132;
output c5149;
output c3243;
output c2211;
output c1141;
output c0109;
output c284;
output c2265;
output c0280;
output c5263;
output c6256;
output c0149;
output c0195;
output c5169;
output c5178;
output c5208;
output c188;
output c0285;
output c0116;
output c2153;
output c5180;
output c2143;
output c1296;
output c190;
output c5252;
output c5288;
output c2110;
output c27;
output c670;
output c6140;
output c785;
output c53;
output c5270;
output c5275;
output c5283;
output c012;
output c498;
output c1268;
output c7273;
output c6213;
output c417;
output c3188;
output c4138;
output c6203;
output c489;
output c5201;
output c6121;
output c7170;
output c5184;
output c1159;
output c383;
output c3197;
output c3108;
output c7279;
output c6237;
output c4238;
output c5214;
output c695;
output c2209;
output c540;
output c2171;
output c1202;
output c3235;
output c5268;
output c176;
output c1153;
output c4102;
output c688;
output c2299;
output c1223;
output c1102;
output c6120;
output c782;
output c170;
output c393;
output c483;
output c7292;
output c5239;
output c729;
output c5285;
output c3245;
output c250;
output c70;
output c6168;
output c412;
output c7135;
output c3138;
output c448;
output c6239;
output c1145;
output c5217;
output c3115;
output c4163;
output c1217;
output c161;
output c1179;
output c6187;
output c4134;
output c6195;
output c042;
output c6260;
output c7130;
output c2113;
output c5254;
output c7281;
output c550;
output c030;
output c754;
output c2238;
output c588;
output c6163;
output c778;
output c416;
output c0251;
output c432;
output c210;
output c0271;
output c575;
output c1222;
output c475;
output c2222;
output c321;
output c5189;
output c29;
output c3136;
output c3255;
output c4192;
output c7298;
output c6253;
output c1143;
output c7228;
output c3213;
output c5241;
output c6199;
output c6244;
output c4213;
output c1104;
output c546;
output c0157;
output c2260;
output c7144;
output c4281;
output c5195;
output c7240;
output c635;
output c2280;
output c3141;
output c3256;
output c4227;
output c3120;
output c565;
output c697;
output c5167;
output c062;
output c4169;
output c746;
output c252;
output c1171;
output c1195;
output c4237;
output c2279;
output c7200;
output c1233;
output c5290;
output c5204;
output c5226;
output c7246;
output c0184;
output c0118;
output c520;
output c7104;
output c2166;
output c1281;
output c6271;
output c02;
output c123;
output c2285;
output c2297;
output c7209;
output c2184;
output c639;
output c0224;
output c587;
output c5192;
output c2136;
output c1127;
output c4215;
output c5246;
output c776;
output c3128;
output c7136;
output c2155;
output c4177;
output c4156;
output c4167;
output c712;
output c3186;
output c427;
output c6240;
output c456;
output c314;
output c1232;
output c0112;
output c573;
output c6251;
output c0187;
output c265;
output c311;
output c2128;
output c379;
output c3294;
output c327;
output c6232;
output c4186;
output c064;
output c477;
output c7229;
output c2188;
output c0243;
output c2123;
output c4150;
output c1213;
output c414;
output c618;
output c0228;
output c4206;
output c6156;
output c382;
output c6254;
output c7176;
output c4137;
output c2135;
output c4257;
output c7138;
output c0186;
output c553;
output c1136;
output c694;
output c4288;
output c4159;
output c647;
output c6298;
output c2150;
output c0216;
output c0106;
output c192;
output c661;
output c167;
output c6233;
output c510;
output c318;
output c290;
output c7190;
output c5247;
output c4166;
output c2177;
output c079;
output c671;
output c4242;
output c7103;
output c5103;
output c4295;
output c2116;
output c6126;
output c750;
output c642;
output c248;
output c2147;
output c268;
output c359;
output c576;
output c5163;
output c4196;
output c4221;
output c458;
output c7285;
output c471;
output c232;
output c4293;
output c5293;
output c3285;
output c1130;
output c4181;
output c4142;
output c7291;
output c4266;
output c026;
output c242;
output c3296;
output c378;
output c169;
output c4172;
output c4278;
output c1228;
output c280;
output c3109;
output c3132;
output c6272;
output c162;
output c7203;
output c3123;
output c071;
output c488;
output c3114;
output c0270;
output c1289;
output c734;
output c221;
output c4298;
output c3232;
output c312;
output c2210;
output c2266;
output c1231;
output c6131;
output c4232;
output c3265;
output c3224;
output c7126;
output c3207;
output c2289;
output c0206;
output c1221;
output c7215;
output c295;
output c788;
output c1188;
output c512;
output c615;
output c6158;
output c7231;
output c2225;
output c352;
output c1109;
output c6178;
output c1101;
output c6269;
output c021;
output c7259;
output c612;
output c6223;
output c3162;
output c6278;
output c1298;
output c4263;
output c5199;
output c0201;
output c189;
output c730;
output c326;
output c317;
output c2199;
output c0258;
output c2168;
output c4225;
output c1291;
output c0173;
output c1263;
output c3111;
output c0141;
output c613;
output c027;
output c2274;
output c469;
output c5240;
output c150;
output c538;
output c7286;
output c2286;
output c7183;
output c5198;
output c0264;
output c7118;
output c771;
output c6288;
output c7129;
output c2104;
output c099;
output c2257;
output c3264;
output c7275;
output c2162;
output c594;
output c4164;
output c54;
output c344;
output c645;
output c665;
output c1200;
output c433;
output c3239;
output c5151;
output c760;
output c0135;
output c315;
output c7237;
output c470;
output c0193;
output c1238;
output c6191;
output c7181;
output c262;
output c1286;
output c0217;
output c595;
output c3156;
output c7214;
output c4228;
output c2127;
output c6261;
output c185;
output c254;
output c683;
output c0248;
output c025;
output c177;
output c5146;
output c097;
output c5125;
output c7164;
output c7114;
output c4178;
output c1283;
output c0163;
output c777;
output c7227;
output c4282;
output c7128;
output c678;
output c5200;
output c3182;
output c7218;
output c5118;
output c164;
output c186;
output c5156;
output c4240;
output c33;
output c472;
output c6295;
output c6101;
output c122;
output c6115;
output c7220;
output c4286;
output c659;
output c2151;
output c2218;
output c5291;
output c4277;
output c0279;
output c5223;
output c492;
output c6255;
output c463;
output c6174;
output c677;
output c7245;
output c3158;
output c329;
output c2156;
output c544;
output c7251;
output c270;
output c1273;
output c5227;
output c7125;
output c264;
output c1257;
output c0231;
output c212;
output c285;
output c522;
output c7250;
output c152;
output c466;
output c142;
output c2206;
output c5256;
output c3218;
output c0233;
output c6114;
output c717;
output c0132;
output c6222;
output c6181;
output c6193;
output c473;
output c253;
output c666;
output c4123;
output c199;
output c42;
output c431;
output c3275;
output c4147;
output c266;
output c2148;
output c634;
output c5115;
output c5161;
output c5183;
output c3261;
output c446;
output c0218;
output c1198;
output c057;
output c120;
output c1277;
output c2158;
output c1254;
output c0227;
output c5155;
output c3202;
output c1269;
output c5114;
output c2120;
output c616;
output c480;
output c751;
output c5128;
output c0208;
output c6227;
output c3152;
output c6277;
output c6141;
output c7264;
output c163;
output c368;
output c0221;
output c6262;
output c0286;
output c786;
output c7153;
output c175;
output c4201;
output c4105;
output c213;
output c5277;
output c1103;
output c350;
output c2185;
output c1135;
output c775;
output c0255;
output c4104;
output c7112;
output c1116;
output c7222;
output c3198;
output c0257;
output c6154;
output c490;
output c082;
output c3263;
output c5175;
output c5101;
output c090;
output c2239;
output c0276;
output c2276;
output c7196;
output c5206;
output c6106;
output c1138;
output c023;
output c0232;
output c256;
output c3151;
output c014;
output c3103;
output c3230;
output c1170;
output c2232;
output c7260;
output c035;
output c1293;
output c5295;
output c5142;
output c4170;
output c5243;
output c5177;
output c5233;
output c3205;
output c356;
output c3126;
output c7236;
output c4168;
output c4121;
output c2198;
output c2134;
output c118;
output c0117;
output c4284;
output c0110;
output c4292;
output c5123;
output c5153;
output c0296;
output c719;
output c6177;
output c548;
output c5299;
output c5145;
output c293;
output c0101;
output c1189;
output c1282;
output c3257;
output c4199;
output c0107;
output c7272;
output c3209;
output c4218;
output c4203;
output c1297;
output c392;
output c2250;
output c038;
output c2220;
output c4110;
output c4193;
output c79;
output c15;
output c319;
output c0142;
output c4264;
output c0242;
output c037;
output c2230;
output c4252;
output c0100;
output c726;
output c184;
output c4173;
output c6282;
output c716;
output c6111;
output c43;
output c4195;
output c2205;
output c033;
output c4296;
output c0180;
output c0103;
output c031;
output c298;
output c5190;
output c3267;
output c365;
output c424;
output c384;
output c3266;
output c2125;
output c3175;
output c5230;
output c6243;
output c3179;
output c691;
output c390;
output c6196;
output c7108;
output c5133;
output c5137;
output c2288;
output c5219;
output c762;
output c7212;
output c178;
output c0214;
output c632;
output c1160;
output c6167;
output c179;
output c534;
output c5135;
output c0123;
output c555;
output c5117;
output c147;
output c2244;
output c6150;
output c790;
output c7171;
output c0247;
output c440;
output c2194;
output c5281;
output c714;
output c363;
output c0147;
output c4133;
output c3268;
output c1246;
output c5119;
output c572;
output c143;
output c40;
output c4243;
output c3159;
output c6228;
output c1216;
output c749;
output c3113;
output c0288;
output c743;
output c3124;
output c024;
output c6110;
output c125;
output c5179;
output c7116;
output c287;
output c5245;
output c574;
output c2141;
output c2183;
output c0261;
output c5297;
output c0156;
output c567;
output c1264;
output c0133;
output c0210;
output c23;
output c7110;
output c484;
output c7182;
output c4220;
output c6214;
output c628;
output c4155;
output c151;
output c468;
output c0281;
output c0139;
output c441;
output c24;
output c5131;
output c144;
output c772;
output c1260;
output c56;
output c4113;
output c1236;
output c5209;
output c3164;
output c1295;
output c3246;
output c447;
output c7284;
output c4235;
output c7151;
output c2216;
output c2223;
output c2284;
output c2157;
output c7253;
output c0200;
output c2193;
output c3160;
output c5166;
output c0176;
output c4158;
output c6291;
output c521;
output c5191;
output c6135;
output c5152;
output c310;
output c3166;
output c479;
output c6160;
output c6116;
output c3241;
output c584;
output c1242;
output c3210;
output c4162;
output c6284;
output c4109;
output c5212;
output c3192;
output c2173;
output c0120;
output c4174;
output c2196;
output c371;
output c0238;
output c5188;
output c5205;
output c2186;
output c66;
output c4285;
output c3193;
output c756;
output c241;
output c425;
output c78;
output c2102;
output c739;
output c6259;
output c3289;
output c0259;
output c7167;
output c7294;
output c214;
output c0178;
output c4141;
output c0121;
output c6133;
output c052;
output c0204;
output c6220;
output c5269;
output c2291;
output c5216;
output c7166;
output c7223;
output c372;
output c7186;
output c5150;
output c4153;
output c453;
output c4261;
output c7270;
output c0174;
output c2208;
output c077;
output c069;
output c1110;
output c3169;
output c6180;
output c322;
output c345;
output c277;
output c6212;
output c590;
output c7265;
output c4236;
output c3125;
output c6194;
output c5289;
output c4209;
output c0152;
output c0148;
output c652;
output c747;
output c5172;
output c0235;
output c2145;
output c3167;
output c581;
output c6172;
output c3134;
output c3142;
output c2207;
output c4100;
output c0283;
output c3195;
output c1240;
output c1258;
output c4132;
output c0256;
output c2201;
output c237;
output c1207;
output c181;
output c243;
output c4216;
output c1266;
output c2181;
output c3248;
output c570;
output c5235;
output c7175;
output c423;
output c437;
output c1267;
output c158;
output c7225;
output c5158;
output c323;
output c1245;
output c276;
output c529;
output c3282;
output c6236;
output c246;
output c2263;
output c564;
output c687;
output c640;
output c336;
output c3118;
output c3225;
output c4191;
output c4106;
output c092;
output c0234;
output c4114;
output c081;
output c193;
output c1288;
output c113;
output c0289;
output c3201;
output c0260;
output c6134;
output c0130;
output c6162;
output c6188;
output c1164;
output c00;
output c1214;
output c624;
output c6209;
output c1108;
output c0155;
output c0299;
output c3249;
output c2108;
output c6276;
output c765;
output c283;
output c7173;
output c1261;
output c5147;
output c1206;
output c4149;
output c0192;
output c1299;
output c560;
output c066;
output c1209;
output c2111;
output c5282;
output c0213;
output c580;
output c436;
output c6183;
output c679;
output c2203;
output c085;
output c111;
output c5258;
output c630;
output c2298;
output c4103;
output c7124;
output c566;
output c6248;
output c1147;
output c60;
output c194;
output c551;
output c5129;
output c585;
output c1191;
output c289;
output c6289;
output c4299;
output c3211;
output c1112;
output c4234;
output c4190;
output c010;
output c561;
output c6161;
output c132;
output c171;
output c0158;
output c48;
output c5211;
output c738;
output c278;
output c1204;
output c684;
output c0230;
output c1106;
output c3146;
output c6287;
output c018;
output c355;
output c227;
output c5294;
output c279;
output c51;
output c149;
output c1100;
output c1177;
output c76;
output c4262;
output c272;
output c0274;
output c182;
output c656;
output c4211;
output c61;
output c7184;
output c124;
output c4108;
output c5272;
output c5278;
output c2103;
output c0162;
output c674;
output c157;
output c3187;
output c770;
output c2140;
output c5174;
output c325;
output c655;
output c4151;
output c068;
output c571;
output c6215;
output c198;
output c21;
output c680;
output c0212;
output c710;
output c2215;
output c6107;
output c682;
output c0181;
output c7192;
output c0203;
output c663;
output c6273;
output c0179;
output c2161;
output c3149;
output c2283;
output c7293;
output c6210;
output c6118;
output c088;
output c5124;
output c028;
output c450;
output c059;
output c3181;
output c7243;
output c7106;
output c7142;
output c7195;
output c0190;
output c7254;
output c4251;
output c1219;
output c4226;
output c787;
output c1137;
output c6235;
output c5104;
output c073;
output c2269;
output c1239;
output c767;
output c0292;
output c3127;
output c6280;
output c723;
output c197;
output c759;
output c6123;
output c3155;
output c641;
output c0160;
output c1275;
output c2219;
output c4120;
output c050;
output c0236;
output c3171;
output c196;
output c7208;
output c0134;
output c1186;
output c0136;
output c3163;
output c2278;
output c0126;
output c6139;
output c3117;
output c4126;
output c5141;
output c4280;
output c4265;
output c5248;
output c3233;
output c6252;
output c6234;
output c3112;
output c2191;
output c4135;
output c1250;
output c3137;
output c2213;
output c741;
output c5231;
output c7178;
output c12;
output c5197;
output c353;
output c7100;
output c6197;
output c0171;
output c7143;
output c526;
output c399;
output c0194;
output c516;
output c781;
output c022;
output c4289;
output c7248;
output c737;
output c455;
output c2178;
output c076;
output c338;
output c7137;
output c369;
output c1121;
output c0183;
output c396;
output c1244;
output c4204;
output c6147;
output c549;
output c7204;
output c1134;
output c5244;
output c3177;
output c1152;
output c1249;
output c260;
output c411;
output c5112;
output c2124;
output c0239;
output c6275;
output c0154;
output c1183;
output c1262;
output c67;
output c646;
output c422;
output c626;
output c0263;
output c554;
output c0104;
output c0199;
output c168;
output c7205;
output c249;
output c065;
output c41;
output c2240;
output c257;
output c5253;
output c7211;
output c745;
output c3105;
output c0252;
output c4117;
output c096;
output c7235;
output c6109;
output c313;
output c5107;
output c6184;
output c44;
output c6149;
output c644;
output c7113;
output c3216;
output c217;
output c4202;
output c5234;
output c7140;
output c1184;
output c7263;
output c482;
output c5220;
output c5113;
output c2236;
output c7156;
output c098;
output c2101;
output c4107;
output c5140;
output c127;
output c3276;
output c5162;
output c4197;
output c1142;
output c35;
output c6132;
output c328;
output c3206;
output c5242;
output c0146;
output c1140;
output c1162;
output c7249;
output c657;
output c1265;
output c26;
output c598;
output c5164;
output c662;
output c690;
output c2233;
output c4219;
output c0161;
output c7262;
output c5229;
output c1199;
output c7158;
output c2221;
output c3295;
output c1285;
output c341;
output c6138;
output c4260;
output c478;
output c0189;
output c6267;
output c0222;
output c1172;
output c3200;
output c2287;
output c6208;
output c1144;
output c675;
output c6124;
output c5100;
output c75;
output c1215;
output c654;
output c3284;
output c676;
output c7252;
output c5264;
output c0293;
output c3281;
output c5126;
output c4182;
output c275;
output c0143;
output c5194;
output c357;
output c3119;
output c1163;
output c2187;
output c4271;
output c4136;
output c47;
output c5273;
output c718;
output c5255;
output c7150;
output c1111;
output c7242;
output c457;
output c514;
output c753;
output c11;
output c649;
output c6205;
output c267;
output c7101;
output c465;
output c1125;
output c2190;
output c3229;
output c4112;
output c6155;
output c286;
output c4194;
output c779;
output c3271;
output c3130;
output c6206;
output c6241;
output c7201;
output c7148;
output c5148;
output c6242;
output c713;
output c4291;
output c5173;
output c3240;
output c445;
output c0284;
output c1271;
output c4185;
output c320;
output c3154;
output c3291;
output c2163;
output c533;
output c5127;
output c68;
output c3297;
output c7131;
output c1173;
output c681;
output c542;
output c5286;
output c3272;
output c5109;
output c1115;
output c6137;
output c054;
output c0131;
output c3116;
output c0266;
output c0170;
output c3269;
output c2100;
output c0290;
output c0191;
output c4250;
output c3129;
output c419;
output c6146;
output c4157;
output c231;
output c03;
output c5213;

assign c00 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x74 &  x77 &  x80 &  x82 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x121 &  x122 &  x125 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x157 &  x158 &  x160 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x195 &  x196 &  x199 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x234 &  x235 &  x236 &  x238 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x274 &  x275 &  x277 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x314 &  x317 &  x320 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x355 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x391 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x433 &  x434 &  x437 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x472 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x497 &  x500 &  x503 &  x506 &  x509 &  x511 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x550 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x628 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x821 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x980 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130 & ~x180 & ~x279 & ~x585 & ~x624 & ~x663 & ~x741 & ~x780 & ~x819;
assign c02 =  x8 &  x11 &  x20 &  x26 &  x29 &  x41 &  x47 &  x50 &  x53 &  x62 &  x68 &  x71 &  x74 &  x80 &  x86 &  x95 &  x104 &  x113 &  x125 &  x128 &  x131 &  x134 &  x140 &  x146 &  x152 &  x155 &  x161 &  x164 &  x173 &  x176 &  x179 &  x181 &  x182 &  x185 &  x197 &  x200 &  x203 &  x206 &  x209 &  x218 &  x220 &  x221 &  x224 &  x230 &  x233 &  x236 &  x241 &  x242 &  x245 &  x247 &  x254 &  x257 &  x260 &  x263 &  x269 &  x272 &  x275 &  x278 &  x281 &  x287 &  x296 &  x299 &  x314 &  x320 &  x323 &  x326 &  x331 &  x332 &  x335 &  x338 &  x350 &  x353 &  x359 &  x362 &  x368 &  x374 &  x383 &  x386 &  x389 &  x395 &  x398 &  x407 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x443 &  x446 &  x455 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x491 &  x500 &  x503 &  x515 &  x518 &  x524 &  x527 &  x533 &  x539 &  x548 &  x551 &  x554 &  x557 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x587 &  x590 &  x596 &  x608 &  x611 &  x617 &  x620 &  x623 &  x626 &  x635 &  x647 &  x650 &  x653 &  x656 &  x662 &  x668 &  x671 &  x677 &  x686 &  x692 &  x695 &  x701 &  x703 &  x704 &  x710 &  x713 &  x719 &  x722 &  x725 &  x731 &  x737 &  x742 &  x743 &  x746 &  x755 &  x758 &  x764 &  x776 &  x779 &  x781 &  x782 &  x788 &  x791 &  x794 &  x803 &  x809 &  x812 &  x815 &  x818 &  x821 &  x830 &  x833 &  x839 &  x842 &  x845 &  x848 &  x857 &  x860 &  x866 &  x869 &  x881 &  x887 &  x898 &  x899 &  x901 &  x902 &  x908 &  x914 &  x917 &  x920 &  x923 &  x940 &  x941 &  x947 &  x959 &  x962 &  x968 &  x971 &  x976 &  x979 &  x980 &  x983 &  x998 &  x1001 &  x1004 &  x1007 &  x1018 &  x1031 &  x1034 &  x1040 &  x1043 &  x1049 &  x1052 &  x1054 &  x1055 &  x1061 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x273 & ~x312 & ~x432 & ~x471 & ~x510 & ~x867;
assign c04 =  x2 &  x5 &  x8 &  x11 &  x23 &  x26 &  x29 &  x38 &  x47 &  x50 &  x53 &  x56 &  x62 &  x65 &  x74 &  x77 &  x83 &  x92 &  x98 &  x101 &  x104 &  x113 &  x122 &  x125 &  x128 &  x134 &  x137 &  x140 &  x146 &  x149 &  x151 &  x155 &  x158 &  x161 &  x182 &  x185 &  x188 &  x203 &  x209 &  x215 &  x218 &  x224 &  x230 &  x233 &  x236 &  x242 &  x247 &  x251 &  x254 &  x269 &  x272 &  x278 &  x286 &  x287 &  x296 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x325 &  x326 &  x338 &  x341 &  x344 &  x350 &  x353 &  x359 &  x362 &  x364 &  x365 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x404 &  x407 &  x410 &  x413 &  x419 &  x425 &  x428 &  x431 &  x440 &  x443 &  x446 &  x449 &  x452 &  x461 &  x464 &  x467 &  x473 &  x476 &  x482 &  x488 &  x491 &  x500 &  x503 &  x512 &  x521 &  x524 &  x530 &  x533 &  x539 &  x554 &  x566 &  x578 &  x580 &  x584 &  x587 &  x590 &  x593 &  x599 &  x602 &  x608 &  x611 &  x617 &  x620 &  x623 &  x629 &  x632 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x671 &  x674 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x701 &  x704 &  x706 &  x710 &  x713 &  x722 &  x725 &  x728 &  x731 &  x737 &  x740 &  x745 &  x746 &  x749 &  x758 &  x761 &  x764 &  x776 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x806 &  x809 &  x812 &  x815 &  x821 &  x827 &  x830 &  x833 &  x839 &  x842 &  x845 &  x848 &  x850 &  x854 &  x857 &  x863 &  x869 &  x875 &  x880 &  x881 &  x884 &  x887 &  x893 &  x899 &  x902 &  x905 &  x908 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x949 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x977 &  x983 &  x989 &  x992 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1033 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 &  x1130;
assign c06 =  x2 &  x5 &  x11 &  x17 &  x20 &  x23 &  x26 &  x29 &  x35 &  x38 &  x47 &  x50 &  x56 &  x59 &  x62 &  x65 &  x74 &  x77 &  x80 &  x83 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x149 &  x152 &  x155 &  x158 &  x167 &  x170 &  x173 &  x176 &  x182 &  x185 &  x194 &  x196 &  x197 &  x200 &  x209 &  x215 &  x221 &  x230 &  x233 &  x234 &  x235 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x263 &  x272 &  x274 &  x275 &  x277 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x308 &  x313 &  x314 &  x316 &  x317 &  x320 &  x326 &  x332 &  x338 &  x341 &  x350 &  x352 &  x353 &  x355 &  x356 &  x359 &  x368 &  x371 &  x374 &  x380 &  x383 &  x386 &  x389 &  x391 &  x392 &  x398 &  x407 &  x410 &  x416 &  x419 &  x425 &  x433 &  x434 &  x437 &  x440 &  x443 &  x446 &  x461 &  x467 &  x470 &  x471 &  x472 &  x476 &  x479 &  x485 &  x488 &  x494 &  x497 &  x500 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x545 &  x550 &  x569 &  x572 &  x578 &  x587 &  x589 &  x596 &  x605 &  x608 &  x611 &  x614 &  x617 &  x623 &  x626 &  x632 &  x638 &  x641 &  x647 &  x650 &  x653 &  x659 &  x665 &  x668 &  x671 &  x677 &  x686 &  x698 &  x701 &  x704 &  x713 &  x719 &  x722 &  x728 &  x731 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x767 &  x770 &  x785 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x815 &  x818 &  x821 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x851 &  x860 &  x863 &  x869 &  x872 &  x875 &  x881 &  x887 &  x890 &  x893 &  x896 &  x899 &  x905 &  x908 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x935 &  x938 &  x950 &  x953 &  x959 &  x962 &  x968 &  x974 &  x977 &  x986 &  x992 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1019 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1058 &  x1061 &  x1073 &  x1085 &  x1088 &  x1097 &  x1109 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x201 & ~x219 & ~x240 & ~x297 & ~x318 & ~x702 & ~x741;
assign c08 =  x8 &  x17 &  x23 &  x68 &  x77 &  x83 &  x89 &  x101 &  x107 &  x113 &  x119 &  x143 &  x146 &  x152 &  x155 &  x173 &  x179 &  x185 &  x191 &  x197 &  x227 &  x242 &  x248 &  x263 &  x281 &  x299 &  x302 &  x308 &  x320 &  x326 &  x329 &  x341 &  x344 &  x377 &  x407 &  x431 &  x434 &  x449 &  x452 &  x455 &  x464 &  x479 &  x491 &  x505 &  x509 &  x512 &  x527 &  x539 &  x542 &  x545 &  x566 &  x617 &  x629 &  x658 &  x680 &  x704 &  x710 &  x737 &  x752 &  x754 &  x758 &  x767 &  x770 &  x773 &  x779 &  x785 &  x791 &  x809 &  x814 &  x818 &  x821 &  x827 &  x836 &  x845 &  x848 &  x852 &  x853 &  x857 &  x887 &  x901 &  x914 &  x917 &  x941 &  x953 &  x962 &  x965 &  x976 &  x980 &  x986 &  x995 &  x1015 &  x1019 &  x1022 &  x1025 &  x1031 &  x1037 &  x1048 &  x1054 &  x1058 &  x1061 &  x1082 &  x1096 &  x1100 &  x1121 &  x1126;
assign c010 =  x14 &  x23 &  x26 &  x29 &  x35 &  x53 &  x65 &  x71 &  x83 &  x104 &  x107 &  x119 &  x130 &  x140 &  x143 &  x152 &  x158 &  x167 &  x169 &  x191 &  x203 &  x212 &  x230 &  x245 &  x251 &  x266 &  x269 &  x293 &  x299 &  x305 &  x320 &  x325 &  x356 &  x362 &  x374 &  x386 &  x389 &  x395 &  x401 &  x410 &  x422 &  x428 &  x437 &  x452 &  x467 &  x470 &  x479 &  x482 &  x485 &  x581 &  x587 &  x589 &  x608 &  x644 &  x653 &  x659 &  x662 &  x677 &  x680 &  x683 &  x686 &  x698 &  x704 &  x713 &  x719 &  x722 &  x731 &  x740 &  x749 &  x764 &  x767 &  x791 &  x797 &  x815 &  x818 &  x821 &  x827 &  x830 &  x845 &  x848 &  x854 &  x857 &  x863 &  x866 &  x878 &  x881 &  x910 &  x935 &  x938 &  x944 &  x947 &  x965 &  x977 &  x986 &  x989 &  x992 &  x998 &  x1010 &  x1013 &  x1031 &  x1055 &  x1058 &  x1067 &  x1072 &  x1085 &  x1094 &  x1103 &  x1109 &  x1124 &  x1127 &  x1130 & ~x138 & ~x453 & ~x846 & ~x1092;
assign c012 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x44 &  x47 &  x50 &  x53 &  x62 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x104 &  x110 &  x116 &  x122 &  x125 &  x131 &  x134 &  x137 &  x143 &  x149 &  x155 &  x158 &  x161 &  x164 &  x167 &  x176 &  x182 &  x185 &  x191 &  x194 &  x197 &  x200 &  x203 &  x209 &  x215 &  x218 &  x221 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x257 &  x260 &  x263 &  x266 &  x275 &  x278 &  x281 &  x284 &  x287 &  x293 &  x302 &  x308 &  x311 &  x320 &  x323 &  x329 &  x338 &  x341 &  x344 &  x347 &  x350 &  x356 &  x359 &  x371 &  x380 &  x386 &  x389 &  x392 &  x395 &  x401 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x434 &  x437 &  x443 &  x446 &  x449 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x479 &  x482 &  x485 &  x488 &  x500 &  x503 &  x512 &  x518 &  x524 &  x533 &  x536 &  x539 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x587 &  x593 &  x596 &  x602 &  x608 &  x611 &  x620 &  x625 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x663 &  x664 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x692 &  x695 &  x698 &  x703 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x731 &  x734 &  x737 &  x740 &  x741 &  x742 &  x743 &  x746 &  x749 &  x752 &  x758 &  x761 &  x764 &  x767 &  x770 &  x776 &  x780 &  x781 &  x782 &  x785 &  x788 &  x791 &  x794 &  x800 &  x806 &  x809 &  x812 &  x815 &  x820 &  x821 &  x827 &  x830 &  x833 &  x839 &  x845 &  x851 &  x854 &  x858 &  x859 &  x860 &  x866 &  x869 &  x872 &  x881 &  x890 &  x893 &  x896 &  x897 &  x901 &  x905 &  x914 &  x920 &  x929 &  x932 &  x935 &  x940 &  x944 &  x947 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x976 &  x979 &  x980 &  x989 &  x995 &  x1001 &  x1007 &  x1015 &  x1016 &  x1018 &  x1019 &  x1022 &  x1031 &  x1034 &  x1049 &  x1052 &  x1054 &  x1058 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x234 & ~x273 & ~x312 & ~x351 & ~x393 & ~x432 & ~x708 & ~x747 & ~x786;
assign c014 =  x2 &  x11 &  x14 &  x17 &  x20 &  x23 &  x32 &  x41 &  x53 &  x62 &  x65 &  x68 &  x71 &  x77 &  x83 &  x92 &  x95 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x134 &  x137 &  x140 &  x143 &  x146 &  x152 &  x155 &  x158 &  x161 &  x167 &  x173 &  x176 &  x179 &  x182 &  x191 &  x197 &  x200 &  x203 &  x206 &  x209 &  x218 &  x221 &  x230 &  x233 &  x236 &  x242 &  x245 &  x257 &  x266 &  x269 &  x272 &  x278 &  x281 &  x287 &  x293 &  x299 &  x308 &  x311 &  x314 &  x317 &  x323 &  x326 &  x332 &  x335 &  x341 &  x344 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x380 &  x383 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x413 &  x419 &  x422 &  x431 &  x433 &  x434 &  x437 &  x440 &  x446 &  x449 &  x458 &  x461 &  x464 &  x472 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x510 &  x512 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x548 &  x550 &  x554 &  x563 &  x566 &  x569 &  x572 &  x575 &  x581 &  x584 &  x588 &  x590 &  x593 &  x596 &  x599 &  x605 &  x608 &  x611 &  x614 &  x628 &  x629 &  x632 &  x635 &  x638 &  x641 &  x647 &  x650 &  x659 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x695 &  x698 &  x704 &  x707 &  x710 &  x716 &  x722 &  x727 &  x731 &  x734 &  x737 &  x749 &  x755 &  x758 &  x766 &  x770 &  x773 &  x779 &  x782 &  x794 &  x797 &  x803 &  x809 &  x812 &  x818 &  x824 &  x827 &  x830 &  x833 &  x842 &  x845 &  x848 &  x851 &  x869 &  x887 &  x890 &  x902 &  x910 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x941 &  x947 &  x949 &  x950 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x988 &  x989 &  x992 &  x995 &  x998 &  x1007 &  x1010 &  x1022 &  x1025 &  x1027 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1103 &  x1105 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x483 & ~x522 & ~x561 & ~x600 & ~x819 & ~x897 & ~x1041 & ~x1053 & ~x1092 & ~x1125;
assign c016 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x323 &  x326 &  x332 &  x335 &  x338 &  x344 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x386 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x430 &  x431 &  x434 &  x437 &  x440 &  x443 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x468 &  x469 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x494 &  x497 &  x500 &  x503 &  x506 &  x507 &  x508 &  x509 &  x515 &  x518 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x546 &  x547 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x625 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x703 &  x706 &  x707 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x742 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x781 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x820 &  x821 &  x823 &  x824 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x851 &  x854 &  x857 &  x859 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x898 &  x899 &  x901 &  x902 &  x905 &  x908 &  x911 &  x914 &  x920 &  x923 &  x926 &  x929 &  x935 &  x938 &  x940 &  x941 &  x944 &  x947 &  x950 &  x953 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x976 &  x977 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1057 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 & ~x474 & ~x513 & ~x552 & ~x675;
assign c018 =  x17 &  x26 &  x35 &  x38 &  x44 &  x50 &  x53 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x89 &  x92 &  x104 &  x128 &  x131 &  x134 &  x149 &  x158 &  x161 &  x164 &  x167 &  x170 &  x194 &  x197 &  x203 &  x212 &  x221 &  x227 &  x239 &  x245 &  x248 &  x251 &  x254 &  x274 &  x284 &  x290 &  x293 &  x299 &  x302 &  x305 &  x314 &  x317 &  x320 &  x323 &  x335 &  x344 &  x347 &  x352 &  x353 &  x362 &  x365 &  x371 &  x374 &  x383 &  x386 &  x392 &  x394 &  x395 &  x398 &  x404 &  x407 &  x419 &  x428 &  x431 &  x433 &  x434 &  x446 &  x461 &  x464 &  x467 &  x472 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x511 &  x512 &  x515 &  x530 &  x533 &  x539 &  x545 &  x550 &  x551 &  x554 &  x569 &  x575 &  x581 &  x593 &  x596 &  x605 &  x623 &  x629 &  x641 &  x644 &  x650 &  x653 &  x662 &  x665 &  x671 &  x683 &  x686 &  x689 &  x716 &  x740 &  x743 &  x751 &  x752 &  x755 &  x761 &  x767 &  x770 &  x773 &  x779 &  x782 &  x791 &  x797 &  x800 &  x811 &  x818 &  x824 &  x827 &  x830 &  x836 &  x838 &  x842 &  x845 &  x851 &  x854 &  x860 &  x869 &  x872 &  x887 &  x893 &  x905 &  x908 &  x914 &  x916 &  x920 &  x923 &  x932 &  x950 &  x955 &  x956 &  x962 &  x967 &  x974 &  x983 &  x986 &  x989 &  x1001 &  x1016 &  x1019 &  x1031 &  x1043 &  x1049 &  x1061 &  x1064 &  x1079 &  x1085 &  x1094 &  x1097 &  x1106 &  x1109 &  x1118 &  x1124 &  x1127 & ~x135 & ~x141 & ~x585;
assign c020 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x274 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x312 &  x313 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x351 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x390 &  x391 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x429 &  x431 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x469 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x508 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x547 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x575 &  x578 &  x581 &  x584 &  x586 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x611 &  x614 &  x617 &  x620 &  x623 &  x625 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x667 &  x668 &  x671 &  x674 &  x677 &  x680 &  x686 &  x692 &  x695 &  x698 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x812 &  x815 &  x818 &  x821 &  x827 &  x830 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130 & ~x318 & ~x357 & ~x358 & ~x396 & ~x435 & ~x474 & ~x558;
assign c022 =  x2 &  x8 &  x14 &  x17 &  x20 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x59 &  x65 &  x68 &  x92 &  x95 &  x98 &  x101 &  x113 &  x116 &  x119 &  x134 &  x137 &  x149 &  x155 &  x158 &  x161 &  x167 &  x176 &  x179 &  x182 &  x185 &  x191 &  x194 &  x197 &  x200 &  x202 &  x203 &  x209 &  x212 &  x221 &  x227 &  x239 &  x241 &  x245 &  x251 &  x260 &  x266 &  x278 &  x281 &  x293 &  x296 &  x299 &  x311 &  x314 &  x317 &  x329 &  x344 &  x350 &  x356 &  x359 &  x362 &  x365 &  x371 &  x377 &  x380 &  x386 &  x389 &  x392 &  x398 &  x404 &  x410 &  x413 &  x416 &  x425 &  x431 &  x434 &  x437 &  x445 &  x446 &  x449 &  x455 &  x461 &  x464 &  x470 &  x479 &  x481 &  x488 &  x494 &  x506 &  x509 &  x512 &  x515 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x551 &  x557 &  x587 &  x593 &  x596 &  x602 &  x605 &  x608 &  x614 &  x617 &  x635 &  x644 &  x647 &  x650 &  x653 &  x659 &  x664 &  x665 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x692 &  x701 &  x703 &  x707 &  x710 &  x713 &  x719 &  x722 &  x731 &  x734 &  x737 &  x740 &  x742 &  x746 &  x749 &  x758 &  x761 &  x764 &  x770 &  x781 &  x785 &  x788 &  x791 &  x797 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x820 &  x821 &  x823 &  x824 &  x833 &  x836 &  x842 &  x845 &  x851 &  x854 &  x857 &  x859 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x898 &  x899 &  x902 &  x911 &  x914 &  x920 &  x926 &  x929 &  x935 &  x938 &  x944 &  x947 &  x950 &  x953 &  x956 &  x962 &  x968 &  x971 &  x974 &  x976 &  x992 &  x995 &  x1004 &  x1015 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1057 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1106 &  x1118 & ~x432 & ~x510 & ~x630 & ~x648 & ~x669 & ~x708 & ~x747 & ~x786;
assign c024 =  x8 &  x11 &  x14 &  x17 &  x23 &  x26 &  x29 &  x32 &  x35 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x92 &  x98 &  x101 &  x104 &  x107 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x140 &  x143 &  x146 &  x149 &  x158 &  x161 &  x167 &  x170 &  x173 &  x176 &  x179 &  x188 &  x194 &  x197 &  x203 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x308 &  x314 &  x317 &  x320 &  x323 &  x325 &  x326 &  x329 &  x335 &  x338 &  x341 &  x347 &  x350 &  x356 &  x359 &  x362 &  x368 &  x383 &  x389 &  x392 &  x398 &  x401 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x431 &  x434 &  x437 &  x440 &  x452 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x509 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x563 &  x566 &  x569 &  x572 &  x575 &  x581 &  x584 &  x587 &  x590 &  x593 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x625 &  x632 &  x635 &  x638 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x671 &  x674 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x703 &  x707 &  x710 &  x716 &  x719 &  x722 &  x725 &  x731 &  x734 &  x737 &  x742 &  x743 &  x746 &  x749 &  x752 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x788 &  x791 &  x794 &  x803 &  x806 &  x809 &  x812 &  x815 &  x820 &  x821 &  x824 &  x830 &  x833 &  x839 &  x842 &  x845 &  x851 &  x854 &  x857 &  x859 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x890 &  x893 &  x898 &  x899 &  x902 &  x905 &  x908 &  x914 &  x917 &  x923 &  x929 &  x932 &  x935 &  x937 &  x938 &  x940 &  x941 &  x944 &  x950 &  x953 &  x956 &  x962 &  x971 &  x974 &  x976 &  x977 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1013 &  x1022 &  x1025 &  x1028 &  x1037 &  x1043 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 & ~x237 & ~x393 & ~x432 & ~x471 & ~x549 & ~x669 & ~x709 & ~x747 & ~x786 & ~x795 & ~x825 & ~x834 & ~x903;
assign c026 =  x2 &  x5 &  x11 &  x14 &  x17 &  x26 &  x29 &  x35 &  x40 &  x47 &  x53 &  x59 &  x62 &  x68 &  x74 &  x77 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x110 &  x113 &  x119 &  x122 &  x125 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x164 &  x167 &  x170 &  x176 &  x182 &  x188 &  x191 &  x203 &  x206 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x236 &  x239 &  x245 &  x248 &  x260 &  x262 &  x269 &  x272 &  x275 &  x278 &  x284 &  x287 &  x290 &  x293 &  x296 &  x301 &  x302 &  x308 &  x314 &  x323 &  x326 &  x332 &  x335 &  x341 &  x347 &  x350 &  x356 &  x359 &  x362 &  x365 &  x368 &  x377 &  x392 &  x397 &  x406 &  x410 &  x413 &  x416 &  x418 &  x419 &  x428 &  x437 &  x443 &  x445 &  x452 &  x458 &  x461 &  x464 &  x470 &  x473 &  x479 &  x484 &  x485 &  x488 &  x496 &  x500 &  x512 &  x518 &  x520 &  x521 &  x524 &  x527 &  x533 &  x542 &  x545 &  x548 &  x554 &  x557 &  x563 &  x569 &  x575 &  x578 &  x584 &  x590 &  x593 &  x596 &  x599 &  x605 &  x608 &  x617 &  x620 &  x626 &  x629 &  x635 &  x647 &  x650 &  x656 &  x662 &  x664 &  x665 &  x671 &  x674 &  x677 &  x680 &  x686 &  x689 &  x695 &  x698 &  x701 &  x703 &  x713 &  x716 &  x719 &  x722 &  x728 &  x737 &  x740 &  x742 &  x743 &  x746 &  x761 &  x764 &  x770 &  x779 &  x782 &  x785 &  x788 &  x797 &  x800 &  x803 &  x809 &  x812 &  x818 &  x820 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x845 &  x848 &  x851 &  x854 &  x869 &  x878 &  x896 &  x905 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x936 &  x938 &  x941 &  x944 &  x950 &  x953 &  x956 &  x974 &  x975 &  x976 &  x980 &  x983 &  x986 &  x989 &  x1001 &  x1004 &  x1010 &  x1014 &  x1016 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1054 &  x1061 &  x1064 &  x1070 &  x1073 &  x1079 &  x1082 &  x1088 &  x1091 &  x1097 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x432 & ~x510 & ~x708;
assign c028 =  x2 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x62 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x143 &  x152 &  x161 &  x167 &  x173 &  x176 &  x179 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x227 &  x233 &  x235 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x274 &  x275 &  x281 &  x287 &  x290 &  x293 &  x296 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x368 &  x371 &  x377 &  x383 &  x386 &  x389 &  x391 &  x392 &  x394 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x430 &  x431 &  x433 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x455 &  x458 &  x461 &  x464 &  x470 &  x472 &  x473 &  x476 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x506 &  x509 &  x511 &  x512 &  x515 &  x521 &  x530 &  x536 &  x539 &  x545 &  x548 &  x550 &  x551 &  x554 &  x560 &  x569 &  x572 &  x575 &  x584 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x680 &  x683 &  x686 &  x688 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x830 &  x833 &  x836 &  x839 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x977 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1055 &  x1058 &  x1061 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1121 &  x1127 &  x1130 & ~x201 & ~x219 & ~x240 & ~x258 & ~x259 & ~x279 & ~x297 & ~x318 & ~x438 & ~x477 & ~x516;
assign c030 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x23 &  x26 &  x32 &  x35 &  x38 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x68 &  x77 &  x83 &  x86 &  x89 &  x95 &  x101 &  x104 &  x110 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x137 &  x140 &  x146 &  x149 &  x155 &  x158 &  x161 &  x164 &  x170 &  x173 &  x176 &  x182 &  x185 &  x188 &  x191 &  x197 &  x200 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x320 &  x323 &  x326 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x362 &  x365 &  x377 &  x380 &  x383 &  x389 &  x392 &  x401 &  x404 &  x407 &  x410 &  x413 &  x419 &  x422 &  x425 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x461 &  x467 &  x470 &  x473 &  x476 &  x479 &  x491 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x550 &  x551 &  x554 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x589 &  x599 &  x602 &  x605 &  x611 &  x614 &  x620 &  x623 &  x625 &  x626 &  x628 &  x629 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x659 &  x662 &  x664 &  x665 &  x667 &  x668 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x703 &  x704 &  x705 &  x706 &  x713 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x744 &  x746 &  x752 &  x755 &  x758 &  x770 &  x773 &  x776 &  x782 &  x783 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x809 &  x815 &  x818 &  x821 &  x823 &  x824 &  x827 &  x833 &  x836 &  x839 &  x842 &  x845 &  x851 &  x854 &  x862 &  x866 &  x875 &  x878 &  x881 &  x884 &  x890 &  x893 &  x896 &  x899 &  x901 &  x902 &  x908 &  x914 &  x917 &  x932 &  x935 &  x940 &  x944 &  x947 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1039 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1078 &  x1079 &  x1082 &  x1085 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1130 & ~x495 & ~x1041 & ~x1080;
assign c032 =  x2 &  x5 &  x7 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x32 &  x35 &  x41 &  x44 &  x47 &  x53 &  x59 &  x62 &  x65 &  x85 &  x86 &  x89 &  x92 &  x95 &  x101 &  x107 &  x110 &  x113 &  x125 &  x134 &  x140 &  x146 &  x149 &  x155 &  x158 &  x167 &  x169 &  x182 &  x191 &  x194 &  x197 &  x200 &  x202 &  x203 &  x206 &  x208 &  x215 &  x218 &  x221 &  x224 &  x227 &  x232 &  x241 &  x245 &  x247 &  x248 &  x251 &  x254 &  x257 &  x259 &  x260 &  x266 &  x269 &  x272 &  x284 &  x287 &  x293 &  x296 &  x298 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x329 &  x332 &  x335 &  x347 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x395 &  x404 &  x407 &  x413 &  x416 &  x425 &  x431 &  x434 &  x437 &  x440 &  x461 &  x467 &  x470 &  x473 &  x479 &  x488 &  x494 &  x497 &  x500 &  x506 &  x509 &  x512 &  x515 &  x521 &  x524 &  x527 &  x536 &  x539 &  x542 &  x545 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x587 &  x593 &  x596 &  x599 &  x602 &  x608 &  x611 &  x617 &  x623 &  x626 &  x632 &  x635 &  x638 &  x641 &  x647 &  x650 &  x656 &  x662 &  x664 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x704 &  x707 &  x710 &  x713 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x742 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x779 &  x781 &  x782 &  x785 &  x791 &  x794 &  x797 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x830 &  x836 &  x839 &  x842 &  x848 &  x857 &  x860 &  x862 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x893 &  x898 &  x902 &  x905 &  x908 &  x911 &  x920 &  x923 &  x926 &  x935 &  x937 &  x938 &  x940 &  x941 &  x947 &  x950 &  x953 &  x956 &  x959 &  x968 &  x971 &  x979 &  x980 &  x983 &  x989 &  x992 &  x998 &  x1001 &  x1007 &  x1013 &  x1018 &  x1019 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1115 &  x1121 &  x1127 &  x1130 & ~x78 & ~x117 & ~x156 & ~x195 & ~x234 & ~x237 & ~x276 & ~x315 & ~x354 & ~x393;
assign c034 =  x5 &  x8 &  x11 &  x14 &  x17 &  x29 &  x38 &  x44 &  x47 &  x50 &  x53 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x95 &  x98 &  x101 &  x107 &  x110 &  x113 &  x119 &  x122 &  x125 &  x128 &  x131 &  x143 &  x149 &  x158 &  x161 &  x167 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x209 &  x212 &  x215 &  x221 &  x224 &  x230 &  x233 &  x236 &  x245 &  x248 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x284 &  x296 &  x299 &  x302 &  x305 &  x314 &  x320 &  x323 &  x326 &  x338 &  x344 &  x347 &  x350 &  x353 &  x356 &  x362 &  x365 &  x368 &  x371 &  x377 &  x380 &  x386 &  x395 &  x401 &  x404 &  x407 &  x413 &  x416 &  x419 &  x428 &  x437 &  x440 &  x446 &  x449 &  x458 &  x461 &  x467 &  x470 &  x473 &  x485 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x518 &  x521 &  x524 &  x533 &  x536 &  x539 &  x542 &  x548 &  x551 &  x554 &  x557 &  x560 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x589 &  x590 &  x593 &  x596 &  x599 &  x602 &  x608 &  x611 &  x617 &  x620 &  x623 &  x628 &  x641 &  x644 &  x653 &  x656 &  x659 &  x662 &  x665 &  x667 &  x671 &  x677 &  x680 &  x683 &  x686 &  x689 &  x695 &  x701 &  x704 &  x705 &  x706 &  x707 &  x710 &  x713 &  x716 &  x722 &  x725 &  x731 &  x733 &  x734 &  x737 &  x743 &  x744 &  x745 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x772 &  x782 &  x783 &  x784 &  x785 &  x788 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x811 &  x815 &  x821 &  x823 &  x824 &  x827 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x849 &  x851 &  x854 &  x862 &  x863 &  x866 &  x872 &  x878 &  x881 &  x884 &  x889 &  x890 &  x893 &  x896 &  x899 &  x901 &  x905 &  x911 &  x914 &  x917 &  x920 &  x929 &  x932 &  x935 &  x938 &  x940 &  x941 &  x950 &  x962 &  x968 &  x971 &  x974 &  x977 &  x979 &  x980 &  x986 &  x992 &  x998 &  x1001 &  x1004 &  x1007 &  x1025 &  x1028 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130;
assign c036 =  x8 &  x17 &  x20 &  x23 &  x26 &  x32 &  x35 &  x38 &  x41 &  x44 &  x53 &  x56 &  x59 &  x62 &  x65 &  x74 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x164 &  x167 &  x176 &  x179 &  x182 &  x185 &  x188 &  x194 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x247 &  x248 &  x254 &  x257 &  x260 &  x263 &  x266 &  x272 &  x278 &  x281 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x323 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x389 &  x392 &  x398 &  x404 &  x413 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x491 &  x500 &  x503 &  x509 &  x511 &  x512 &  x515 &  x518 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x550 &  x554 &  x557 &  x560 &  x566 &  x569 &  x572 &  x575 &  x581 &  x584 &  x587 &  x589 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x627 &  x628 &  x632 &  x641 &  x644 &  x647 &  x650 &  x653 &  x659 &  x662 &  x665 &  x666 &  x667 &  x668 &  x671 &  x677 &  x680 &  x683 &  x689 &  x692 &  x695 &  x701 &  x704 &  x705 &  x706 &  x707 &  x710 &  x716 &  x719 &  x722 &  x725 &  x728 &  x734 &  x737 &  x743 &  x744 &  x745 &  x746 &  x749 &  x752 &  x758 &  x761 &  x764 &  x773 &  x776 &  x779 &  x782 &  x783 &  x784 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x890 &  x896 &  x899 &  x901 &  x902 &  x905 &  x908 &  x911 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1058 &  x1060 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1088 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x0 & ~x156 & ~x195 & ~x495 & ~x534;
assign c038 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x312 &  x313 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x380 &  x383 &  x386 &  x389 &  x391 &  x394 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x430 &  x431 &  x433 &  x434 &  x437 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x469 &  x470 &  x472 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x508 &  x511 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x550 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x628 &  x629 &  x632 &  x635 &  x638 &  x644 &  x647 &  x653 &  x656 &  x662 &  x665 &  x667 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x695 &  x701 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x812 &  x815 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x877 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x905 &  x908 &  x914 &  x916 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x336 & ~x375 & ~x522 & ~x561 & ~x702 & ~x741 & ~x780 & ~x819 & ~x858;
assign c040 =  x5 &  x8 &  x14 &  x17 &  x20 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x143 &  x149 &  x152 &  x155 &  x161 &  x170 &  x173 &  x176 &  x182 &  x185 &  x188 &  x191 &  x197 &  x209 &  x212 &  x221 &  x224 &  x227 &  x230 &  x233 &  x235 &  x245 &  x251 &  x254 &  x257 &  x260 &  x263 &  x269 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x317 &  x320 &  x323 &  x329 &  x335 &  x338 &  x341 &  x347 &  x350 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x391 &  x392 &  x394 &  x395 &  x398 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x430 &  x431 &  x434 &  x437 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x472 &  x473 &  x476 &  x485 &  x494 &  x500 &  x503 &  x506 &  x509 &  x511 &  x512 &  x515 &  x521 &  x527 &  x539 &  x545 &  x550 &  x557 &  x560 &  x563 &  x566 &  x569 &  x575 &  x578 &  x581 &  x587 &  x590 &  x593 &  x596 &  x602 &  x604 &  x617 &  x620 &  x623 &  x629 &  x632 &  x635 &  x638 &  x641 &  x642 &  x644 &  x647 &  x650 &  x653 &  x656 &  x662 &  x665 &  x668 &  x671 &  x674 &  x680 &  x682 &  x683 &  x686 &  x689 &  x698 &  x701 &  x707 &  x710 &  x713 &  x716 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x743 &  x746 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x815 &  x818 &  x821 &  x824 &  x827 &  x833 &  x836 &  x839 &  x842 &  x845 &  x851 &  x854 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x905 &  x908 &  x914 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x950 &  x953 &  x959 &  x962 &  x965 &  x968 &  x974 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1067 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x258 & ~x780 & ~x819 & ~x858;
assign c042 =  x5 &  x8 &  x11 &  x17 &  x26 &  x29 &  x32 &  x38 &  x44 &  x47 &  x53 &  x56 &  x68 &  x71 &  x74 &  x77 &  x83 &  x86 &  x89 &  x101 &  x104 &  x107 &  x119 &  x122 &  x131 &  x134 &  x137 &  x152 &  x155 &  x164 &  x167 &  x173 &  x176 &  x182 &  x187 &  x188 &  x197 &  x200 &  x206 &  x209 &  x212 &  x218 &  x230 &  x233 &  x236 &  x245 &  x248 &  x254 &  x260 &  x263 &  x265 &  x271 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x296 &  x299 &  x305 &  x308 &  x311 &  x317 &  x320 &  x323 &  x326 &  x332 &  x338 &  x341 &  x347 &  x350 &  x353 &  x356 &  x365 &  x371 &  x377 &  x380 &  x386 &  x389 &  x398 &  x404 &  x407 &  x413 &  x416 &  x419 &  x422 &  x431 &  x443 &  x446 &  x455 &  x461 &  x464 &  x467 &  x476 &  x479 &  x488 &  x491 &  x497 &  x509 &  x512 &  x521 &  x524 &  x533 &  x539 &  x542 &  x545 &  x572 &  x581 &  x584 &  x587 &  x590 &  x593 &  x605 &  x608 &  x617 &  x623 &  x626 &  x635 &  x638 &  x641 &  x647 &  x665 &  x668 &  x671 &  x674 &  x680 &  x686 &  x692 &  x698 &  x710 &  x716 &  x722 &  x731 &  x734 &  x740 &  x745 &  x746 &  x749 &  x752 &  x761 &  x770 &  x784 &  x785 &  x788 &  x794 &  x800 &  x803 &  x809 &  x812 &  x815 &  x821 &  x824 &  x839 &  x848 &  x861 &  x862 &  x866 &  x869 &  x881 &  x896 &  x900 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x940 &  x941 &  x950 &  x953 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x977 &  x979 &  x980 &  x989 &  x995 &  x998 &  x1001 &  x1010 &  x1013 &  x1016 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1049 &  x1055 &  x1058 &  x1064 &  x1076 &  x1079 &  x1082 &  x1085 &  x1094 &  x1100 &  x1106 &  x1109 &  x1112 &  x1114 &  x1115 &  x1118 &  x1127 & ~x789 & ~x828 & ~x906;
assign c044 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x124 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x325 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x364 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x704 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x916 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x955 &  x959 &  x962 &  x965 &  x968 &  x974 &  x977 &  x983 &  x986 &  x989 &  x992 &  x994 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1072 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1111 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x174 & ~x252 & ~x330;
assign c046 =  x5 &  x8 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x89 &  x92 &  x95 &  x98 &  x101 &  x107 &  x110 &  x113 &  x116 &  x122 &  x125 &  x131 &  x134 &  x137 &  x140 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x173 &  x179 &  x182 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x266 &  x269 &  x272 &  x275 &  x281 &  x284 &  x290 &  x293 &  x299 &  x305 &  x308 &  x314 &  x317 &  x323 &  x326 &  x329 &  x332 &  x335 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x437 &  x440 &  x443 &  x446 &  x452 &  x455 &  x458 &  x464 &  x467 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x625 &  x626 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x703 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x742 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x781 &  x785 &  x788 &  x791 &  x794 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x820 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x851 &  x854 &  x859 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x893 &  x896 &  x898 &  x899 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x935 &  x938 &  x940 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x976 &  x977 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1015 &  x1016 &  x1018 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1054 &  x1055 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 & ~x276 & ~x354 & ~x393 & ~x432 & ~x471 & ~x510 & ~x549 & ~x630 & ~x669 & ~x670 & ~x708 & ~x747 & ~x748 & ~x786 & ~x787 & ~x831 & ~x864 & ~x870;
assign c048 =  x2 &  x5 &  x8 &  x11 &  x23 &  x26 &  x35 &  x38 &  x44 &  x62 &  x65 &  x89 &  x92 &  x95 &  x98 &  x107 &  x110 &  x125 &  x128 &  x131 &  x140 &  x149 &  x155 &  x158 &  x161 &  x173 &  x179 &  x185 &  x188 &  x194 &  x209 &  x215 &  x221 &  x224 &  x230 &  x233 &  x235 &  x239 &  x248 &  x251 &  x254 &  x257 &  x273 &  x281 &  x284 &  x287 &  x290 &  x293 &  x311 &  x314 &  x317 &  x320 &  x335 &  x347 &  x352 &  x359 &  x374 &  x377 &  x386 &  x398 &  x401 &  x410 &  x413 &  x419 &  x434 &  x440 &  x443 &  x446 &  x461 &  x467 &  x470 &  x482 &  x485 &  x512 &  x515 &  x518 &  x521 &  x527 &  x530 &  x536 &  x542 &  x548 &  x551 &  x557 &  x560 &  x569 &  x572 &  x578 &  x587 &  x593 &  x602 &  x611 &  x614 &  x620 &  x623 &  x626 &  x632 &  x635 &  x637 &  x638 &  x644 &  x650 &  x653 &  x668 &  x674 &  x676 &  x686 &  x695 &  x698 &  x707 &  x710 &  x719 &  x722 &  x737 &  x755 &  x764 &  x767 &  x770 &  x773 &  x776 &  x794 &  x806 &  x812 &  x824 &  x827 &  x833 &  x839 &  x854 &  x863 &  x878 &  x881 &  x884 &  x893 &  x896 &  x905 &  x908 &  x914 &  x920 &  x932 &  x941 &  x965 &  x968 &  x974 &  x980 &  x983 &  x986 &  x992 &  x1001 &  x1010 &  x1013 &  x1025 &  x1028 &  x1034 &  x1040 &  x1043 &  x1049 &  x1052 &  x1061 &  x1064 &  x1073 &  x1079 &  x1088 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1130 & ~x123 & ~x162 & ~x201 & ~x213 & ~x321 & ~x360 & ~x399 & ~x705 & ~x1056;
assign c050 =  x8 &  x11 &  x20 &  x35 &  x38 &  x44 &  x47 &  x56 &  x59 &  x68 &  x71 &  x74 &  x89 &  x92 &  x98 &  x104 &  x110 &  x116 &  x119 &  x128 &  x131 &  x140 &  x143 &  x149 &  x152 &  x155 &  x167 &  x170 &  x173 &  x176 &  x179 &  x185 &  x194 &  x197 &  x206 &  x218 &  x224 &  x227 &  x230 &  x236 &  x254 &  x260 &  x266 &  x278 &  x281 &  x287 &  x293 &  x296 &  x311 &  x317 &  x323 &  x329 &  x332 &  x335 &  x338 &  x344 &  x350 &  x356 &  x362 &  x368 &  x380 &  x383 &  x389 &  x392 &  x395 &  x410 &  x419 &  x422 &  x428 &  x431 &  x433 &  x437 &  x446 &  x452 &  x461 &  x467 &  x472 &  x473 &  x476 &  x479 &  x488 &  x491 &  x500 &  x510 &  x511 &  x521 &  x530 &  x533 &  x549 &  x550 &  x551 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x587 &  x588 &  x596 &  x599 &  x605 &  x608 &  x611 &  x620 &  x628 &  x632 &  x641 &  x656 &  x659 &  x662 &  x665 &  x667 &  x671 &  x677 &  x689 &  x701 &  x706 &  x716 &  x725 &  x728 &  x737 &  x740 &  x745 &  x749 &  x752 &  x758 &  x761 &  x764 &  x770 &  x784 &  x785 &  x788 &  x800 &  x803 &  x812 &  x823 &  x827 &  x842 &  x857 &  x863 &  x872 &  x878 &  x883 &  x899 &  x905 &  x911 &  x914 &  x917 &  x929 &  x938 &  x950 &  x953 &  x956 &  x962 &  x965 &  x971 &  x974 &  x980 &  x989 &  x1004 &  x1013 &  x1022 &  x1025 &  x1031 &  x1037 &  x1040 &  x1043 &  x1055 &  x1061 &  x1064 &  x1076 &  x1079 &  x1094 &  x1103 &  x1109 &  x1112 &  x1115 &  x1121 &  x1127 &  x1130 & ~x0 & ~x222 & ~x261 & ~x300 & ~x741 & ~x780 & ~x1014;
assign c052 =  x2 &  x8 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x89 &  x92 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x122 &  x131 &  x134 &  x140 &  x146 &  x149 &  x155 &  x158 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x200 &  x203 &  x206 &  x212 &  x215 &  x218 &  x224 &  x233 &  x236 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x272 &  x278 &  x281 &  x284 &  x286 &  x287 &  x293 &  x296 &  x305 &  x311 &  x314 &  x317 &  x323 &  x325 &  x326 &  x329 &  x335 &  x341 &  x344 &  x347 &  x350 &  x353 &  x359 &  x362 &  x365 &  x374 &  x383 &  x386 &  x392 &  x407 &  x410 &  x416 &  x419 &  x422 &  x428 &  x434 &  x440 &  x443 &  x446 &  x449 &  x452 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x491 &  x494 &  x497 &  x506 &  x512 &  x515 &  x518 &  x521 &  x527 &  x530 &  x536 &  x539 &  x542 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x580 &  x581 &  x584 &  x590 &  x593 &  x596 &  x599 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x638 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x743 &  x746 &  x752 &  x755 &  x758 &  x761 &  x770 &  x782 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x842 &  x845 &  x848 &  x854 &  x856 &  x857 &  x860 &  x863 &  x866 &  x872 &  x875 &  x881 &  x884 &  x887 &  x893 &  x896 &  x899 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x941 &  x944 &  x947 &  x953 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x983 &  x986 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 & ~x81 & ~x120 & ~x159 & ~x243 & ~x276 & ~x315 & ~x354 & ~x393 & ~x432 & ~x630 & ~x747;
assign c054 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x104 &  x107 &  x110 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x391 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x429 &  x430 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x468 &  x469 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x508 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x547 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x625 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x703 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x733 &  x734 &  x737 &  x740 &  x742 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x955 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x994 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x474;
assign c056 =  x2 &  x5 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x163 &  x164 &  x167 &  x170 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x236 &  x239 &  x242 &  x245 &  x247 &  x248 &  x251 &  x254 &  x257 &  x266 &  x269 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x389 &  x392 &  x395 &  x401 &  x404 &  x407 &  x410 &  x413 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x545 &  x548 &  x550 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x587 &  x596 &  x599 &  x602 &  x605 &  x611 &  x617 &  x620 &  x623 &  x626 &  x627 &  x628 &  x632 &  x635 &  x638 &  x644 &  x647 &  x650 &  x653 &  x659 &  x662 &  x665 &  x666 &  x667 &  x668 &  x671 &  x674 &  x680 &  x683 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x705 &  x706 &  x707 &  x710 &  x713 &  x716 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x744 &  x745 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x803 &  x806 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x830 &  x839 &  x842 &  x848 &  x851 &  x854 &  x857 &  x860 &  x866 &  x869 &  x872 &  x875 &  x878 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x941 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1033 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1072 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1127 & ~x0 & ~x39 & ~x78 & ~x117 & ~x339 & ~x378 & ~x417 & ~x1014 & ~x1053 & ~x1092;
assign c058 =  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x80 &  x86 &  x89 &  x91 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x164 &  x167 &  x169 &  x170 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x667 &  x668 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x706 &  x707 &  x710 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x920 &  x922 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x949 &  x950 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x980 &  x982 &  x983 &  x986 &  x988 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1027 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1066 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1105 &  x1106 &  x1109 &  x1111 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x39 & ~x78 & ~x117 & ~x300 & ~x339 & ~x378 & ~x1014 & ~x1053 & ~x1092;
assign c060 =  x2 &  x5 &  x14 &  x17 &  x23 &  x26 &  x32 &  x41 &  x53 &  x56 &  x59 &  x62 &  x68 &  x77 &  x80 &  x92 &  x95 &  x101 &  x107 &  x110 &  x113 &  x116 &  x119 &  x125 &  x137 &  x143 &  x146 &  x155 &  x158 &  x167 &  x173 &  x182 &  x191 &  x194 &  x200 &  x209 &  x218 &  x221 &  x227 &  x230 &  x236 &  x242 &  x254 &  x260 &  x266 &  x269 &  x272 &  x311 &  x314 &  x320 &  x332 &  x338 &  x341 &  x344 &  x347 &  x362 &  x365 &  x368 &  x374 &  x380 &  x392 &  x395 &  x398 &  x404 &  x407 &  x419 &  x431 &  x434 &  x437 &  x440 &  x449 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x494 &  x497 &  x506 &  x509 &  x515 &  x533 &  x539 &  x563 &  x581 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x628 &  x635 &  x638 &  x647 &  x662 &  x667 &  x671 &  x692 &  x695 &  x704 &  x707 &  x713 &  x716 &  x725 &  x728 &  x731 &  x740 &  x746 &  x752 &  x755 &  x758 &  x764 &  x806 &  x812 &  x815 &  x833 &  x836 &  x845 &  x857 &  x860 &  x872 &  x878 &  x881 &  x884 &  x890 &  x893 &  x902 &  x908 &  x911 &  x926 &  x938 &  x944 &  x950 &  x953 &  x956 &  x968 &  x971 &  x980 &  x986 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1031 &  x1033 &  x1034 &  x1037 &  x1049 &  x1055 &  x1058 &  x1067 &  x1072 &  x1073 &  x1076 &  x1088 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1124 & ~x369 & ~x396 & ~x696 & ~x702 & ~x735 & ~x741 & ~x774 & ~x1041 & ~x1080;
assign c062 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x122 &  x125 &  x128 &  x134 &  x137 &  x140 &  x146 &  x149 &  x152 &  x155 &  x158 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x230 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x323 &  x326 &  x329 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x359 &  x362 &  x365 &  x374 &  x377 &  x380 &  x386 &  x389 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x430 &  x434 &  x437 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x467 &  x468 &  x469 &  x470 &  x479 &  x482 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x507 &  x508 &  x509 &  x511 &  x512 &  x515 &  x518 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x547 &  x548 &  x550 &  x551 &  x554 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x589 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x625 &  x626 &  x628 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x659 &  x664 &  x665 &  x667 &  x668 &  x671 &  x674 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x703 &  x704 &  x706 &  x707 &  x710 &  x719 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x742 &  x743 &  x745 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x809 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x836 &  x839 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x871 &  x872 &  x875 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x910 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x940 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1124 &  x1127 &  x1130 & ~x474 & ~x513 & ~x552 & ~x597;
assign c064 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x32 &  x38 &  x47 &  x50 &  x56 &  x59 &  x65 &  x68 &  x71 &  x80 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x113 &  x116 &  x122 &  x128 &  x131 &  x134 &  x137 &  x143 &  x146 &  x173 &  x185 &  x191 &  x196 &  x200 &  x203 &  x206 &  x215 &  x221 &  x224 &  x230 &  x233 &  x235 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x257 &  x260 &  x263 &  x269 &  x272 &  x273 &  x274 &  x275 &  x277 &  x281 &  x284 &  x287 &  x293 &  x296 &  x299 &  x305 &  x311 &  x313 &  x316 &  x317 &  x326 &  x329 &  x332 &  x338 &  x347 &  x350 &  x353 &  x354 &  x356 &  x359 &  x362 &  x365 &  x371 &  x377 &  x386 &  x401 &  x404 &  x410 &  x422 &  x425 &  x433 &  x440 &  x449 &  x455 &  x464 &  x467 &  x470 &  x471 &  x472 &  x476 &  x494 &  x497 &  x500 &  x503 &  x509 &  x510 &  x512 &  x524 &  x527 &  x533 &  x536 &  x539 &  x542 &  x545 &  x550 &  x554 &  x557 &  x569 &  x572 &  x581 &  x584 &  x587 &  x589 &  x590 &  x596 &  x602 &  x608 &  x614 &  x620 &  x623 &  x626 &  x628 &  x629 &  x632 &  x635 &  x638 &  x641 &  x647 &  x653 &  x656 &  x665 &  x668 &  x677 &  x680 &  x683 &  x686 &  x689 &  x695 &  x710 &  x713 &  x728 &  x734 &  x740 &  x749 &  x764 &  x770 &  x791 &  x794 &  x797 &  x803 &  x806 &  x812 &  x815 &  x818 &  x821 &  x824 &  x830 &  x839 &  x845 &  x848 &  x851 &  x854 &  x866 &  x872 &  x875 &  x881 &  x887 &  x893 &  x899 &  x905 &  x917 &  x923 &  x926 &  x929 &  x932 &  x938 &  x941 &  x944 &  x947 &  x950 &  x956 &  x962 &  x965 &  x968 &  x974 &  x977 &  x980 &  x986 &  x989 &  x992 &  x998 &  x1001 &  x1007 &  x1010 &  x1019 &  x1022 &  x1025 &  x1031 &  x1040 &  x1043 &  x1049 &  x1058 &  x1061 &  x1067 &  x1082 &  x1085 &  x1091 &  x1100 &  x1106 &  x1109 &  x1118 &  x1121 &  x1124 &  x1130 & ~x201 & ~x240 & ~x702 & ~x741 & ~x780 & ~x819;
assign c066 =  x5 &  x14 &  x17 &  x20 &  x26 &  x29 &  x35 &  x44 &  x62 &  x68 &  x71 &  x74 &  x77 &  x86 &  x89 &  x92 &  x95 &  x101 &  x104 &  x110 &  x119 &  x122 &  x131 &  x134 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x164 &  x173 &  x176 &  x179 &  x191 &  x197 &  x200 &  x203 &  x209 &  x212 &  x215 &  x221 &  x230 &  x232 &  x242 &  x248 &  x251 &  x257 &  x260 &  x266 &  x269 &  x272 &  x275 &  x281 &  x284 &  x290 &  x296 &  x299 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x386 &  x389 &  x392 &  x395 &  x398 &  x404 &  x407 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x437 &  x440 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x481 &  x482 &  x485 &  x488 &  x494 &  x500 &  x506 &  x512 &  x517 &  x518 &  x524 &  x527 &  x530 &  x533 &  x536 &  x542 &  x551 &  x554 &  x556 &  x557 &  x563 &  x569 &  x575 &  x578 &  x580 &  x581 &  x584 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x611 &  x614 &  x623 &  x629 &  x632 &  x635 &  x647 &  x650 &  x653 &  x662 &  x665 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x695 &  x698 &  x701 &  x703 &  x707 &  x716 &  x728 &  x731 &  x734 &  x737 &  x743 &  x746 &  x752 &  x761 &  x764 &  x776 &  x779 &  x781 &  x782 &  x788 &  x800 &  x806 &  x809 &  x815 &  x818 &  x830 &  x833 &  x839 &  x842 &  x845 &  x854 &  x857 &  x860 &  x866 &  x869 &  x872 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x905 &  x911 &  x914 &  x917 &  x920 &  x923 &  x938 &  x940 &  x941 &  x944 &  x947 &  x950 &  x956 &  x959 &  x965 &  x968 &  x971 &  x979 &  x980 &  x986 &  x989 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1067 &  x1070 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x432 & ~x531 & ~x606;
assign c068 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x65 &  x68 &  x74 &  x80 &  x86 &  x107 &  x119 &  x122 &  x128 &  x137 &  x146 &  x149 &  x155 &  x161 &  x164 &  x169 &  x170 &  x179 &  x197 &  x212 &  x227 &  x230 &  x233 &  x236 &  x245 &  x251 &  x263 &  x284 &  x290 &  x302 &  x314 &  x320 &  x344 &  x347 &  x350 &  x353 &  x359 &  x362 &  x368 &  x371 &  x392 &  x395 &  x398 &  x407 &  x413 &  x425 &  x428 &  x433 &  x434 &  x446 &  x449 &  x455 &  x458 &  x470 &  x472 &  x473 &  x476 &  x479 &  x482 &  x488 &  x494 &  x506 &  x509 &  x512 &  x518 &  x530 &  x542 &  x548 &  x550 &  x578 &  x584 &  x587 &  x590 &  x593 &  x617 &  x632 &  x641 &  x650 &  x665 &  x667 &  x674 &  x677 &  x686 &  x689 &  x698 &  x706 &  x725 &  x728 &  x740 &  x746 &  x749 &  x758 &  x761 &  x767 &  x773 &  x782 &  x785 &  x806 &  x809 &  x821 &  x824 &  x827 &  x833 &  x836 &  x839 &  x842 &  x843 &  x848 &  x851 &  x872 &  x883 &  x884 &  x887 &  x899 &  x902 &  x908 &  x910 &  x911 &  x914 &  x920 &  x926 &  x935 &  x938 &  x941 &  x950 &  x953 &  x956 &  x959 &  x962 &  x974 &  x977 &  x986 &  x989 &  x995 &  x998 &  x1000 &  x1004 &  x1019 &  x1022 &  x1037 &  x1043 &  x1058 &  x1067 &  x1073 &  x1079 &  x1085 &  x1097 &  x1106 &  x1121 &  x1127 &  x1130 & ~x39 & ~x261 & ~x300;
assign c070 =  x5 &  x8 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x77 &  x80 &  x83 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x116 &  x125 &  x128 &  x131 &  x137 &  x143 &  x149 &  x155 &  x161 &  x170 &  x173 &  x176 &  x191 &  x194 &  x209 &  x212 &  x215 &  x230 &  x239 &  x242 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x278 &  x284 &  x286 &  x287 &  x290 &  x293 &  x296 &  x302 &  x304 &  x305 &  x311 &  x320 &  x326 &  x332 &  x335 &  x341 &  x343 &  x344 &  x347 &  x350 &  x353 &  x356 &  x371 &  x377 &  x383 &  x386 &  x392 &  x395 &  x397 &  x401 &  x404 &  x416 &  x419 &  x422 &  x428 &  x434 &  x440 &  x455 &  x467 &  x482 &  x491 &  x494 &  x503 &  x506 &  x509 &  x515 &  x518 &  x524 &  x527 &  x536 &  x539 &  x545 &  x548 &  x554 &  x557 &  x560 &  x572 &  x584 &  x590 &  x605 &  x623 &  x625 &  x626 &  x629 &  x635 &  x638 &  x641 &  x647 &  x656 &  x664 &  x665 &  x677 &  x686 &  x689 &  x692 &  x701 &  x704 &  x707 &  x710 &  x716 &  x725 &  x731 &  x743 &  x746 &  x755 &  x767 &  x770 &  x779 &  x782 &  x785 &  x791 &  x794 &  x797 &  x803 &  x809 &  x812 &  x821 &  x824 &  x827 &  x836 &  x842 &  x854 &  x857 &  x860 &  x862 &  x869 &  x872 &  x878 &  x884 &  x896 &  x899 &  x901 &  x905 &  x908 &  x917 &  x938 &  x940 &  x941 &  x947 &  x950 &  x953 &  x962 &  x965 &  x978 &  x983 &  x986 &  x1001 &  x1007 &  x1010 &  x1018 &  x1022 &  x1025 &  x1031 &  x1040 &  x1043 &  x1046 &  x1052 &  x1058 &  x1061 &  x1073 &  x1085 &  x1091 &  x1097 &  x1100 &  x1103 &  x1112 &  x1130 & ~x234 & ~x273 & ~x393 & ~x432 & ~x573;
assign c072 =  x2 &  x5 &  x8 &  x11 &  x14 &  x32 &  x41 &  x47 &  x50 &  x56 &  x62 &  x77 &  x89 &  x95 &  x110 &  x119 &  x122 &  x131 &  x143 &  x149 &  x152 &  x158 &  x167 &  x170 &  x176 &  x179 &  x182 &  x188 &  x197 &  x215 &  x224 &  x227 &  x233 &  x236 &  x242 &  x251 &  x260 &  x266 &  x269 &  x290 &  x305 &  x308 &  x314 &  x320 &  x323 &  x329 &  x332 &  x335 &  x338 &  x353 &  x356 &  x359 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x386 &  x401 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x434 &  x437 &  x440 &  x443 &  x449 &  x455 &  x467 &  x485 &  x488 &  x494 &  x497 &  x509 &  x512 &  x515 &  x524 &  x530 &  x536 &  x548 &  x551 &  x554 &  x557 &  x560 &  x569 &  x581 &  x587 &  x599 &  x605 &  x617 &  x629 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x659 &  x676 &  x683 &  x686 &  x689 &  x692 &  x698 &  x704 &  x713 &  x716 &  x725 &  x728 &  x731 &  x737 &  x743 &  x746 &  x749 &  x757 &  x758 &  x773 &  x776 &  x779 &  x797 &  x800 &  x803 &  x809 &  x821 &  x824 &  x827 &  x836 &  x839 &  x854 &  x860 &  x863 &  x866 &  x872 &  x875 &  x878 &  x893 &  x899 &  x905 &  x917 &  x926 &  x938 &  x941 &  x944 &  x956 &  x959 &  x962 &  x965 &  x968 &  x977 &  x1010 &  x1013 &  x1019 &  x1022 &  x1031 &  x1040 &  x1052 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1100 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 & ~x201 & ~x213 & ~x219 & ~x240 & ~x279 & ~x357 & ~x402 & ~x480 & ~x867 & ~x984;
assign c074 =  x2 &  x5 &  x11 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x107 &  x113 &  x116 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x317 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x362 &  x365 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x419 &  x422 &  x431 &  x434 &  x437 &  x443 &  x446 &  x449 &  x455 &  x458 &  x461 &  x467 &  x469 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x497 &  x500 &  x506 &  x507 &  x508 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x533 &  x539 &  x542 &  x545 &  x546 &  x547 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x590 &  x593 &  x596 &  x599 &  x605 &  x608 &  x611 &  x617 &  x620 &  x623 &  x625 &  x626 &  x629 &  x632 &  x635 &  x638 &  x647 &  x650 &  x653 &  x656 &  x659 &  x664 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x701 &  x703 &  x704 &  x707 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x737 &  x740 &  x742 &  x743 &  x749 &  x752 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x815 &  x818 &  x820 &  x821 &  x823 &  x824 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x860 &  x862 &  x863 &  x866 &  x869 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x901 &  x902 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x940 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x195 & ~x234 & ~x354 & ~x474 & ~x492 & ~x552 & ~x591;
assign c076 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x508 &  x509 &  x511 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x547 &  x548 &  x550 &  x551 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x625 &  x626 &  x628 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x656 &  x659 &  x662 &  x665 &  x667 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x703 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x731 &  x734 &  x737 &  x740 &  x743 &  x744 &  x745 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x818 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x863 &  x865 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x890 &  x896 &  x899 &  x901 &  x902 &  x905 &  x908 &  x911 &  x914 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x940 &  x941 &  x944 &  x947 &  x949 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130 & ~x513 & ~x552;
assign c078 =  x8 &  x11 &  x35 &  x41 &  x47 &  x65 &  x68 &  x77 &  x80 &  x83 &  x89 &  x95 &  x113 &  x122 &  x128 &  x143 &  x155 &  x158 &  x173 &  x179 &  x182 &  x188 &  x209 &  x218 &  x232 &  x236 &  x239 &  x254 &  x257 &  x265 &  x266 &  x281 &  x290 &  x296 &  x320 &  x323 &  x329 &  x335 &  x338 &  x344 &  x347 &  x353 &  x356 &  x362 &  x365 &  x368 &  x377 &  x392 &  x398 &  x407 &  x422 &  x431 &  x446 &  x449 &  x455 &  x476 &  x481 &  x494 &  x503 &  x530 &  x548 &  x560 &  x562 &  x563 &  x575 &  x578 &  x584 &  x587 &  x635 &  x641 &  x647 &  x650 &  x653 &  x656 &  x665 &  x683 &  x710 &  x716 &  x725 &  x745 &  x749 &  x752 &  x761 &  x767 &  x776 &  x779 &  x809 &  x812 &  x851 &  x878 &  x890 &  x898 &  x900 &  x911 &  x937 &  x950 &  x959 &  x962 &  x974 &  x976 &  x977 &  x979 &  x980 &  x983 &  x986 &  x1013 &  x1018 &  x1031 &  x1040 &  x1046 &  x1049 &  x1056 &  x1082 &  x1091 &  x1124 & ~x306 & ~x312 & ~x423 & ~x462;
assign c080 =  x2 &  x5 &  x11 &  x14 &  x17 &  x20 &  x35 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x68 &  x71 &  x74 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x116 &  x119 &  x122 &  x134 &  x137 &  x140 &  x155 &  x158 &  x161 &  x167 &  x170 &  x173 &  x179 &  x182 &  x185 &  x194 &  x197 &  x203 &  x206 &  x212 &  x221 &  x224 &  x233 &  x239 &  x242 &  x244 &  x245 &  x248 &  x251 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x317 &  x320 &  x323 &  x326 &  x329 &  x341 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x383 &  x386 &  x391 &  x392 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x430 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x469 &  x470 &  x485 &  x491 &  x497 &  x503 &  x506 &  x508 &  x518 &  x524 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x566 &  x569 &  x572 &  x581 &  x587 &  x593 &  x605 &  x608 &  x611 &  x614 &  x616 &  x617 &  x620 &  x623 &  x626 &  x632 &  x635 &  x638 &  x641 &  x644 &  x653 &  x656 &  x659 &  x665 &  x674 &  x677 &  x680 &  x686 &  x692 &  x695 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x746 &  x752 &  x755 &  x764 &  x767 &  x770 &  x773 &  x782 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x815 &  x833 &  x836 &  x842 &  x845 &  x848 &  x851 &  x854 &  x860 &  x863 &  x866 &  x872 &  x875 &  x878 &  x884 &  x887 &  x890 &  x893 &  x902 &  x911 &  x914 &  x920 &  x923 &  x926 &  x929 &  x938 &  x941 &  x949 &  x959 &  x962 &  x965 &  x974 &  x977 &  x980 &  x983 &  x988 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1049 &  x1052 &  x1058 &  x1061 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x6 & ~x45 & ~x855 & ~x1020 & ~x1098;
assign c082 =  x44 &  x50 &  x56 &  x59 &  x68 &  x83 &  x89 &  x95 &  x101 &  x113 &  x119 &  x125 &  x131 &  x143 &  x146 &  x158 &  x167 &  x170 &  x173 &  x179 &  x197 &  x200 &  x212 &  x215 &  x218 &  x227 &  x239 &  x245 &  x248 &  x254 &  x263 &  x275 &  x287 &  x301 &  x302 &  x308 &  x311 &  x314 &  x320 &  x323 &  x338 &  x344 &  x350 &  x365 &  x380 &  x382 &  x401 &  x407 &  x410 &  x422 &  x428 &  x437 &  x449 &  x457 &  x461 &  x464 &  x467 &  x476 &  x482 &  x488 &  x512 &  x518 &  x533 &  x536 &  x545 &  x548 &  x560 &  x566 &  x575 &  x581 &  x584 &  x587 &  x599 &  x602 &  x605 &  x608 &  x617 &  x629 &  x632 &  x638 &  x640 &  x647 &  x656 &  x659 &  x665 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x701 &  x704 &  x713 &  x722 &  x725 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x757 &  x767 &  x770 &  x773 &  x776 &  x782 &  x791 &  x796 &  x803 &  x806 &  x809 &  x812 &  x821 &  x827 &  x830 &  x833 &  x836 &  x848 &  x854 &  x860 &  x863 &  x869 &  x878 &  x884 &  x896 &  x902 &  x911 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x938 &  x944 &  x947 &  x953 &  x956 &  x965 &  x971 &  x974 &  x980 &  x983 &  x986 &  x992 &  x998 &  x1001 &  x1010 &  x1031 &  x1034 &  x1043 &  x1046 &  x1049 &  x1058 &  x1061 &  x1064 &  x1067 &  x1076 &  x1085 &  x1103 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130 & ~x180 & ~x627 & ~x666 & ~x669 & ~x708 & ~x744 & ~x747 & ~x825 & ~x864;
assign c084 =  x2 &  x23 &  x47 &  x59 &  x71 &  x74 &  x89 &  x107 &  x110 &  x113 &  x116 &  x117 &  x121 &  x125 &  x143 &  x152 &  x160 &  x170 &  x188 &  x191 &  x194 &  x197 &  x199 &  x203 &  x212 &  x221 &  x234 &  x235 &  x236 &  x238 &  x239 &  x245 &  x254 &  x266 &  x272 &  x326 &  x329 &  x338 &  x347 &  x350 &  x352 &  x356 &  x362 &  x368 &  x371 &  x374 &  x389 &  x392 &  x394 &  x398 &  x404 &  x422 &  x428 &  x443 &  x446 &  x461 &  x479 &  x482 &  x485 &  x488 &  x491 &  x506 &  x509 &  x518 &  x524 &  x530 &  x536 &  x542 &  x551 &  x578 &  x581 &  x587 &  x590 &  x596 &  x605 &  x614 &  x617 &  x620 &  x623 &  x635 &  x644 &  x659 &  x665 &  x668 &  x677 &  x698 &  x704 &  x710 &  x718 &  x719 &  x722 &  x725 &  x743 &  x749 &  x757 &  x758 &  x760 &  x764 &  x767 &  x776 &  x791 &  x799 &  x806 &  x809 &  x812 &  x818 &  x824 &  x827 &  x830 &  x848 &  x860 &  x872 &  x878 &  x887 &  x893 &  x902 &  x914 &  x926 &  x929 &  x932 &  x938 &  x941 &  x944 &  x956 &  x959 &  x983 &  x998 &  x1001 &  x1004 &  x1019 &  x1028 &  x1031 &  x1034 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1076 &  x1085 &  x1091 &  x1094 &  x1097 &  x1103 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 & ~x220 & ~x375 & ~x819 & ~x858;
assign c086 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x44 &  x47 &  x53 &  x56 &  x59 &  x65 &  x71 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x101 &  x104 &  x107 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x234 &  x235 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x274 &  x275 &  x278 &  x284 &  x287 &  x290 &  x293 &  x299 &  x302 &  x308 &  x311 &  x313 &  x314 &  x316 &  x317 &  x320 &  x323 &  x329 &  x332 &  x338 &  x341 &  x344 &  x350 &  x352 &  x353 &  x355 &  x356 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x391 &  x392 &  x394 &  x395 &  x398 &  x404 &  x407 &  x410 &  x413 &  x419 &  x422 &  x425 &  x431 &  x433 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x458 &  x461 &  x470 &  x472 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x509 &  x511 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x605 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x716 &  x719 &  x722 &  x725 &  x728 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x799 &  x803 &  x806 &  x812 &  x815 &  x818 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x902 &  x905 &  x908 &  x911 &  x914 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 & ~x213 & ~x219 & ~x252 & ~x258 & ~x259 & ~x279 & ~x297 & ~x318 & ~x477 & ~x663 & ~x702 & ~x741 & ~x780 & ~x819 & ~x858;
assign c088 =  x23 &  x38 &  x44 &  x47 &  x53 &  x68 &  x110 &  x155 &  x156 &  x195 &  x199 &  x236 &  x248 &  x277 &  x284 &  x290 &  x356 &  x368 &  x386 &  x391 &  x394 &  x434 &  x472 &  x503 &  x521 &  x569 &  x620 &  x623 &  x656 &  x659 &  x680 &  x681 &  x686 &  x689 &  x709 &  x722 &  x748 &  x760 &  x782 &  x799 &  x821 &  x827 &  x836 &  x893 &  x905 &  x911 &  x923 &  x926 &  x953 &  x980 &  x989 &  x1052 &  x1058 &  x1097 &  x1124 &  x1130 & ~x546 & ~x624 & ~x741;
assign c090 =  x11 &  x14 &  x17 &  x23 &  x26 &  x29 &  x35 &  x44 &  x47 &  x50 &  x56 &  x59 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x107 &  x110 &  x122 &  x134 &  x137 &  x143 &  x158 &  x161 &  x167 &  x173 &  x176 &  x179 &  x191 &  x194 &  x206 &  x209 &  x215 &  x224 &  x227 &  x230 &  x233 &  x236 &  x242 &  x245 &  x251 &  x260 &  x269 &  x275 &  x278 &  x281 &  x287 &  x296 &  x299 &  x305 &  x316 &  x320 &  x323 &  x329 &  x332 &  x335 &  x344 &  x350 &  x353 &  x356 &  x365 &  x368 &  x374 &  x377 &  x389 &  x394 &  x407 &  x410 &  x413 &  x416 &  x425 &  x428 &  x431 &  x437 &  x452 &  x455 &  x461 &  x464 &  x470 &  x473 &  x476 &  x479 &  x494 &  x509 &  x515 &  x521 &  x530 &  x539 &  x545 &  x550 &  x557 &  x560 &  x563 &  x614 &  x617 &  x626 &  x635 &  x638 &  x647 &  x650 &  x653 &  x659 &  x665 &  x674 &  x677 &  x683 &  x689 &  x692 &  x695 &  x698 &  x701 &  x707 &  x719 &  x728 &  x734 &  x737 &  x740 &  x743 &  x746 &  x748 &  x749 &  x752 &  x755 &  x767 &  x770 &  x773 &  x776 &  x782 &  x785 &  x791 &  x818 &  x824 &  x826 &  x827 &  x830 &  x836 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x865 &  x866 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x910 &  x911 &  x914 &  x917 &  x923 &  x935 &  x938 &  x941 &  x947 &  x949 &  x950 &  x953 &  x956 &  x959 &  x965 &  x974 &  x977 &  x980 &  x988 &  x1001 &  x1007 &  x1019 &  x1022 &  x1025 &  x1027 &  x1028 &  x1031 &  x1046 &  x1049 &  x1052 &  x1055 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1094 &  x1097 &  x1103 &  x1106 & ~x99 & ~x702 & ~x735 & ~x774 & ~x963 & ~x1014 & ~x1092;
assign c092 =  x8 &  x17 &  x32 &  x34 &  x35 &  x38 &  x53 &  x56 &  x67 &  x73 &  x74 &  x77 &  x89 &  x106 &  x110 &  x125 &  x128 &  x134 &  x137 &  x140 &  x146 &  x167 &  x182 &  x188 &  x194 &  x212 &  x227 &  x239 &  x242 &  x251 &  x257 &  x263 &  x266 &  x287 &  x290 &  x299 &  x305 &  x311 &  x314 &  x326 &  x329 &  x338 &  x341 &  x347 &  x350 &  x362 &  x365 &  x371 &  x377 &  x383 &  x392 &  x395 &  x404 &  x431 &  x443 &  x449 &  x452 &  x455 &  x461 &  x464 &  x473 &  x482 &  x491 &  x494 &  x497 &  x500 &  x503 &  x512 &  x518 &  x530 &  x533 &  x536 &  x539 &  x542 &  x548 &  x557 &  x563 &  x569 &  x578 &  x584 &  x593 &  x596 &  x605 &  x611 &  x614 &  x617 &  x623 &  x625 &  x635 &  x638 &  x659 &  x662 &  x664 &  x665 &  x667 &  x668 &  x680 &  x683 &  x698 &  x703 &  x713 &  x725 &  x731 &  x737 &  x742 &  x746 &  x761 &  x767 &  x776 &  x806 &  x820 &  x830 &  x839 &  x842 &  x859 &  x862 &  x863 &  x866 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x926 &  x935 &  x941 &  x950 &  x968 &  x1004 &  x1007 &  x1010 &  x1016 &  x1019 &  x1031 &  x1034 &  x1049 &  x1052 &  x1058 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1088 &  x1094 &  x1103 &  x1106 &  x1112 & ~x474 & ~x648 & ~x972;
assign c094 =  x10 &  x56 &  x65 &  x86 &  x95 &  x155 &  x195 &  x235 &  x257 &  x320 &  x326 &  x347 &  x352 &  x365 &  x368 &  x371 &  x394 &  x401 &  x422 &  x446 &  x491 &  x503 &  x526 &  x577 &  x587 &  x590 &  x614 &  x617 &  x626 &  x629 &  x638 &  x642 &  x644 &  x650 &  x659 &  x662 &  x665 &  x689 &  x709 &  x713 &  x716 &  x722 &  x728 &  x740 &  x749 &  x797 &  x803 &  x806 &  x824 &  x839 &  x863 &  x872 &  x908 &  x998 &  x1034 &  x1037 &  x1082 &  x1094 &  x1112;
assign c096 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x212 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x491 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x572 &  x575 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x728 &  x731 &  x734 &  x737 &  x740 &  x742 &  x743 &  x745 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x781 &  x782 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x815 &  x818 &  x820 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x859 &  x860 &  x862 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x898 &  x899 &  x901 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x940 &  x941 &  x944 &  x947 &  x953 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 & ~x150 & ~x177 & ~x189 & ~x306 & ~x345 & ~x378 & ~x567 & ~x606 & ~x645 & ~x648;
assign c098 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x47 &  x50 &  x56 &  x62 &  x65 &  x67 &  x68 &  x71 &  x74 &  x77 &  x80 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x122 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x194 &  x197 &  x200 &  x203 &  x218 &  x221 &  x227 &  x233 &  x239 &  x245 &  x248 &  x251 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x379 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x431 &  x434 &  x436 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x467 &  x470 &  x476 &  x479 &  x482 &  x485 &  x488 &  x497 &  x506 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x545 &  x554 &  x560 &  x562 &  x563 &  x566 &  x569 &  x572 &  x575 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x598 &  x599 &  x601 &  x602 &  x608 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x647 &  x650 &  x656 &  x659 &  x662 &  x668 &  x671 &  x674 &  x680 &  x683 &  x686 &  x689 &  x692 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x740 &  x746 &  x749 &  x752 &  x755 &  x757 &  x758 &  x761 &  x764 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x794 &  x797 &  x806 &  x809 &  x815 &  x818 &  x827 &  x830 &  x833 &  x836 &  x839 &  x845 &  x848 &  x851 &  x857 &  x860 &  x863 &  x869 &  x872 &  x881 &  x887 &  x890 &  x893 &  x899 &  x905 &  x911 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x956 &  x959 &  x962 &  x968 &  x971 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1025 &  x1031 &  x1040 &  x1043 &  x1046 &  x1052 &  x1061 &  x1067 &  x1073 &  x1076 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 & ~x12 & ~x669 & ~x708 & ~x870 & ~x909 & ~x948;
assign c0100 =  x2 &  x5 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x197 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x224 &  x227 &  x239 &  x242 &  x245 &  x247 &  x248 &  x254 &  x257 &  x260 &  x263 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x317 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x362 &  x365 &  x368 &  x371 &  x374 &  x380 &  x383 &  x386 &  x395 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x419 &  x422 &  x428 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x509 &  x512 &  x518 &  x524 &  x527 &  x530 &  x533 &  x536 &  x542 &  x545 &  x548 &  x551 &  x557 &  x560 &  x566 &  x572 &  x575 &  x578 &  x584 &  x586 &  x587 &  x589 &  x593 &  x596 &  x602 &  x608 &  x611 &  x614 &  x617 &  x623 &  x626 &  x628 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x656 &  x662 &  x665 &  x667 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x704 &  x706 &  x707 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x758 &  x760 &  x761 &  x764 &  x767 &  x770 &  x773 &  x779 &  x784 &  x785 &  x788 &  x791 &  x794 &  x798 &  x799 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x836 &  x838 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 & ~x120 & ~x159;
assign c0102 =  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x89 &  x92 &  x95 &  x104 &  x110 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x140 &  x146 &  x149 &  x152 &  x155 &  x158 &  x164 &  x167 &  x173 &  x176 &  x179 &  x182 &  x185 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x281 &  x287 &  x290 &  x293 &  x296 &  x308 &  x311 &  x314 &  x317 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x380 &  x386 &  x392 &  x395 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x431 &  x437 &  x442 &  x443 &  x449 &  x455 &  x461 &  x464 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x506 &  x509 &  x512 &  x518 &  x521 &  x524 &  x530 &  x533 &  x536 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x575 &  x584 &  x593 &  x599 &  x602 &  x605 &  x611 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x668 &  x671 &  x674 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x703 &  x704 &  x707 &  x713 &  x719 &  x722 &  x725 &  x731 &  x734 &  x737 &  x740 &  x742 &  x743 &  x746 &  x752 &  x755 &  x758 &  x761 &  x767 &  x769 &  x770 &  x773 &  x776 &  x779 &  x781 &  x782 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x820 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x847 &  x848 &  x851 &  x854 &  x857 &  x859 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x885 &  x886 &  x887 &  x890 &  x893 &  x896 &  x898 &  x899 &  x901 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x938 &  x940 &  x941 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x979 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1018 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1057 &  x1058 &  x1061 &  x1064 &  x1067 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1096 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1124 &  x1127 &  x1130 & ~x159 & ~x198 & ~x237 & ~x276 & ~x432;
assign c0104 =  x2 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x56 &  x59 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x95 &  x101 &  x104 &  x107 &  x110 &  x113 &  x119 &  x122 &  x125 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x266 &  x269 &  x272 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x298 &  x299 &  x302 &  x305 &  x308 &  x311 &  x317 &  x319 &  x323 &  x326 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x368 &  x374 &  x377 &  x380 &  x386 &  x389 &  x395 &  x398 &  x404 &  x407 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x440 &  x443 &  x445 &  x446 &  x449 &  x452 &  x461 &  x464 &  x467 &  x470 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x503 &  x506 &  x509 &  x512 &  x515 &  x521 &  x524 &  x527 &  x530 &  x539 &  x542 &  x545 &  x551 &  x554 &  x557 &  x563 &  x566 &  x572 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x611 &  x614 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x662 &  x664 &  x665 &  x668 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x703 &  x704 &  x707 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x740 &  x742 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x767 &  x773 &  x776 &  x779 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x803 &  x806 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x836 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x878 &  x881 &  x887 &  x890 &  x893 &  x896 &  x899 &  x901 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x956 &  x959 &  x962 &  x968 &  x971 &  x974 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1019 &  x1022 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x234 & ~x273 & ~x312 & ~x528 & ~x534;
assign c0106 =  x2 &  x5 &  x20 &  x23 &  x26 &  x38 &  x50 &  x53 &  x62 &  x68 &  x77 &  x80 &  x89 &  x92 &  x95 &  x98 &  x101 &  x107 &  x112 &  x116 &  x122 &  x125 &  x134 &  x140 &  x143 &  x146 &  x149 &  x155 &  x158 &  x164 &  x170 &  x178 &  x179 &  x184 &  x188 &  x191 &  x200 &  x217 &  x221 &  x223 &  x227 &  x236 &  x242 &  x245 &  x248 &  x263 &  x269 &  x272 &  x275 &  x278 &  x284 &  x295 &  x301 &  x302 &  x311 &  x314 &  x317 &  x320 &  x326 &  x329 &  x332 &  x338 &  x339 &  x341 &  x347 &  x353 &  x359 &  x362 &  x374 &  x379 &  x386 &  x389 &  x392 &  x400 &  x404 &  x413 &  x416 &  x425 &  x428 &  x439 &  x440 &  x443 &  x452 &  x455 &  x473 &  x476 &  x479 &  x485 &  x497 &  x502 &  x506 &  x515 &  x518 &  x521 &  x523 &  x524 &  x530 &  x533 &  x539 &  x541 &  x542 &  x545 &  x551 &  x557 &  x559 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x593 &  x598 &  x599 &  x602 &  x605 &  x608 &  x614 &  x620 &  x626 &  x632 &  x638 &  x644 &  x647 &  x650 &  x659 &  x671 &  x674 &  x680 &  x686 &  x689 &  x692 &  x695 &  x698 &  x722 &  x725 &  x731 &  x746 &  x752 &  x764 &  x767 &  x770 &  x776 &  x779 &  x791 &  x797 &  x812 &  x818 &  x821 &  x827 &  x830 &  x833 &  x839 &  x845 &  x851 &  x860 &  x863 &  x866 &  x875 &  x878 &  x884 &  x893 &  x899 &  x905 &  x914 &  x917 &  x919 &  x923 &  x929 &  x941 &  x944 &  x950 &  x953 &  x956 &  x958 &  x959 &  x962 &  x971 &  x976 &  x977 &  x980 &  x983 &  x989 &  x998 &  x1010 &  x1013 &  x1016 &  x1022 &  x1031 &  x1037 &  x1040 &  x1043 &  x1055 &  x1058 &  x1061 &  x1070 &  x1076 &  x1091 &  x1100 &  x1115 &  x1118 &  x1124 &  x1127;
assign c0108 =  x53 &  x65 &  x74 &  x86 &  x98 &  x122 &  x134 &  x140 &  x200 &  x203 &  x209 &  x215 &  x221 &  x239 &  x248 &  x284 &  x290 &  x308 &  x329 &  x332 &  x362 &  x365 &  x368 &  x380 &  x395 &  x404 &  x416 &  x470 &  x473 &  x482 &  x488 &  x518 &  x521 &  x539 &  x542 &  x578 &  x587 &  x599 &  x608 &  x647 &  x665 &  x689 &  x701 &  x707 &  x710 &  x728 &  x734 &  x742 &  x746 &  x764 &  x776 &  x779 &  x781 &  x815 &  x830 &  x842 &  x845 &  x854 &  x858 &  x866 &  x869 &  x899 &  x935 &  x936 &  x956 &  x965 &  x968 &  x979 &  x983 &  x1013 &  x1019 &  x1028 &  x1055 &  x1073 &  x1088 &  x1112 & ~x315 & ~x354 & ~x393 & ~x603 & ~x687 & ~x708 & ~x726 & ~x843;
assign c0110 =  x2 &  x5 &  x8 &  x11 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x50 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x113 &  x116 &  x119 &  x122 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x155 &  x158 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x182 &  x185 &  x197 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x220 &  x221 &  x224 &  x227 &  x230 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x259 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x365 &  x368 &  x371 &  x374 &  x389 &  x392 &  x395 &  x398 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x470 &  x473 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x542 &  x545 &  x548 &  x551 &  x554 &  x560 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x590 &  x593 &  x596 &  x599 &  x605 &  x611 &  x617 &  x620 &  x623 &  x625 &  x626 &  x629 &  x632 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x703 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x731 &  x734 &  x737 &  x740 &  x742 &  x746 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x820 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x859 &  x860 &  x862 &  x863 &  x866 &  x869 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x896 &  x898 &  x899 &  x901 &  x902 &  x905 &  x908 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x937 &  x938 &  x941 &  x947 &  x950 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1049 &  x1055 &  x1058 &  x1061 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x234 & ~x273 & ~x393 & ~x489 & ~x513 & ~x552 & ~x630 & ~x631 & ~x669 & ~x708;
assign c0112 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x91 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x236 &  x239 &  x242 &  x245 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x401 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x430 &  x431 &  x434 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x832 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x988 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1027 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x396 & ~x435 & ~x474 & ~x489 & ~x528 & ~x555 & ~x594 & ~x633;
assign c0114 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x32 &  x35 &  x44 &  x50 &  x56 &  x59 &  x65 &  x68 &  x71 &  x74 &  x83 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x167 &  x170 &  x182 &  x188 &  x197 &  x203 &  x212 &  x215 &  x218 &  x221 &  x224 &  x233 &  x235 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x263 &  x266 &  x269 &  x272 &  x273 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x314 &  x316 &  x317 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x355 &  x356 &  x359 &  x362 &  x365 &  x368 &  x374 &  x386 &  x389 &  x391 &  x392 &  x394 &  x395 &  x398 &  x401 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x449 &  x452 &  x455 &  x461 &  x464 &  x470 &  x472 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x503 &  x509 &  x511 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x542 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x575 &  x578 &  x593 &  x599 &  x602 &  x611 &  x614 &  x620 &  x623 &  x632 &  x635 &  x644 &  x650 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x760 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x797 &  x799 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x827 &  x836 &  x839 &  x842 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x881 &  x887 &  x896 &  x902 &  x917 &  x920 &  x926 &  x929 &  x932 &  x938 &  x947 &  x950 &  x959 &  x962 &  x965 &  x968 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1028 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1061 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x213 & ~x219 & ~x258 & ~x585 & ~x663 & ~x741 & ~x780 & ~x819 & ~x822 & ~x858 & ~x900 & ~x939 & ~x1056;
assign c0116 =  x8 &  x11 &  x20 &  x23 &  x26 &  x32 &  x35 &  x47 &  x50 &  x53 &  x56 &  x62 &  x65 &  x71 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x113 &  x117 &  x118 &  x119 &  x122 &  x125 &  x128 &  x137 &  x143 &  x146 &  x152 &  x155 &  x157 &  x158 &  x161 &  x164 &  x170 &  x176 &  x179 &  x182 &  x185 &  x191 &  x196 &  x206 &  x212 &  x215 &  x218 &  x221 &  x233 &  x234 &  x236 &  x248 &  x251 &  x254 &  x257 &  x260 &  x262 &  x269 &  x272 &  x274 &  x278 &  x281 &  x284 &  x293 &  x299 &  x301 &  x302 &  x305 &  x313 &  x314 &  x317 &  x320 &  x326 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x352 &  x359 &  x365 &  x368 &  x374 &  x377 &  x380 &  x386 &  x389 &  x398 &  x401 &  x404 &  x410 &  x413 &  x422 &  x425 &  x428 &  x434 &  x440 &  x446 &  x449 &  x470 &  x473 &  x479 &  x482 &  x485 &  x488 &  x491 &  x500 &  x503 &  x506 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x545 &  x551 &  x557 &  x560 &  x572 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x605 &  x611 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x638 &  x641 &  x644 &  x650 &  x656 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x683 &  x688 &  x692 &  x695 &  x701 &  x716 &  x719 &  x725 &  x727 &  x728 &  x734 &  x737 &  x743 &  x746 &  x752 &  x755 &  x757 &  x758 &  x760 &  x764 &  x766 &  x767 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x794 &  x800 &  x803 &  x806 &  x809 &  x815 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x869 &  x875 &  x877 &  x878 &  x881 &  x896 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x938 &  x941 &  x950 &  x953 &  x956 &  x962 &  x974 &  x980 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1028 &  x1031 &  x1034 &  x1043 &  x1046 &  x1049 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1088 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1130 & ~x123 & ~x282 & ~x861;
assign c0118 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x41 &  x44 &  x47 &  x56 &  x59 &  x62 &  x65 &  x71 &  x74 &  x77 &  x80 &  x83 &  x89 &  x92 &  x95 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x131 &  x134 &  x137 &  x143 &  x146 &  x149 &  x152 &  x155 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x197 &  x200 &  x203 &  x206 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x299 &  x308 &  x311 &  x314 &  x317 &  x320 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x400 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x464 &  x467 &  x469 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x508 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x546 &  x547 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x590 &  x593 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x625 &  x626 &  x632 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x667 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x737 &  x740 &  x742 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x783 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x812 &  x815 &  x818 &  x823 &  x824 &  x827 &  x830 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x857 &  x860 &  x862 &  x863 &  x866 &  x869 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x901 &  x902 &  x908 &  x911 &  x917 &  x920 &  x923 &  x926 &  x929 &  x935 &  x938 &  x940 &  x941 &  x944 &  x950 &  x953 &  x956 &  x959 &  x962 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1130 & ~x492 & ~x531 & ~x570;
assign c0120 =  x2 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x125 &  x131 &  x134 &  x140 &  x149 &  x152 &  x158 &  x161 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x194 &  x197 &  x200 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x239 &  x242 &  x254 &  x257 &  x260 &  x263 &  x266 &  x278 &  x281 &  x284 &  x290 &  x296 &  x299 &  x302 &  x320 &  x323 &  x326 &  x329 &  x335 &  x338 &  x341 &  x350 &  x353 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x380 &  x389 &  x392 &  x395 &  x404 &  x413 &  x431 &  x434 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x467 &  x473 &  x476 &  x479 &  x485 &  x491 &  x503 &  x506 &  x509 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x542 &  x548 &  x554 &  x557 &  x560 &  x566 &  x569 &  x572 &  x575 &  x584 &  x587 &  x590 &  x593 &  x596 &  x602 &  x605 &  x608 &  x620 &  x623 &  x632 &  x635 &  x644 &  x647 &  x653 &  x674 &  x677 &  x680 &  x683 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x710 &  x713 &  x716 &  x719 &  x722 &  x731 &  x734 &  x737 &  x740 &  x758 &  x764 &  x767 &  x770 &  x779 &  x788 &  x797 &  x803 &  x806 &  x812 &  x815 &  x818 &  x824 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x875 &  x878 &  x884 &  x890 &  x893 &  x901 &  x902 &  x908 &  x911 &  x914 &  x917 &  x920 &  x926 &  x935 &  x938 &  x944 &  x947 &  x950 &  x953 &  x959 &  x962 &  x968 &  x971 &  x977 &  x979 &  x980 &  x983 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1055 &  x1057 &  x1058 &  x1061 &  x1064 &  x1067 &  x1076 &  x1079 &  x1082 &  x1085 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x6 & ~x46 & ~x84 & ~x162 & ~x168 & ~x267 & ~x306 & ~x384;
assign c0122 =  x5 &  x11 &  x35 &  x65 &  x104 &  x125 &  x200 &  x206 &  x209 &  x212 &  x248 &  x251 &  x257 &  x260 &  x266 &  x272 &  x278 &  x296 &  x299 &  x302 &  x311 &  x314 &  x338 &  x341 &  x362 &  x368 &  x395 &  x401 &  x404 &  x443 &  x455 &  x482 &  x488 &  x491 &  x500 &  x503 &  x518 &  x521 &  x539 &  x545 &  x547 &  x569 &  x584 &  x596 &  x611 &  x620 &  x644 &  x653 &  x667 &  x677 &  x689 &  x716 &  x725 &  x745 &  x770 &  x782 &  x785 &  x788 &  x809 &  x842 &  x881 &  x884 &  x905 &  x914 &  x917 &  x932 &  x950 &  x953 &  x983 &  x989 &  x1025 &  x1034 &  x1040 &  x1046 &  x1055 &  x1073 &  x1085 &  x1088 &  x1094 &  x1118 &  x1130 & ~x249 & ~x486 & ~x564 & ~x604 & ~x681 & ~x1041 & ~x1080;
assign c0124 =  x8 &  x9 &  x10 &  x14 &  x17 &  x20 &  x23 &  x26 &  x38 &  x44 &  x50 &  x53 &  x59 &  x68 &  x71 &  x82 &  x86 &  x89 &  x98 &  x107 &  x110 &  x113 &  x117 &  x119 &  x125 &  x131 &  x134 &  x137 &  x143 &  x146 &  x149 &  x155 &  x157 &  x160 &  x161 &  x170 &  x179 &  x182 &  x188 &  x191 &  x196 &  x199 &  x203 &  x206 &  x209 &  x215 &  x218 &  x227 &  x230 &  x233 &  x235 &  x236 &  x239 &  x242 &  x248 &  x254 &  x257 &  x260 &  x263 &  x266 &  x272 &  x274 &  x275 &  x277 &  x278 &  x281 &  x293 &  x302 &  x305 &  x316 &  x317 &  x320 &  x338 &  x344 &  x347 &  x353 &  x355 &  x359 &  x362 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x394 &  x395 &  x398 &  x407 &  x410 &  x416 &  x419 &  x433 &  x437 &  x446 &  x452 &  x455 &  x458 &  x460 &  x461 &  x464 &  x467 &  x472 &  x473 &  x476 &  x479 &  x485 &  x488 &  x497 &  x500 &  x503 &  x509 &  x512 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x557 &  x566 &  x569 &  x572 &  x578 &  x581 &  x584 &  x593 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x626 &  x629 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x659 &  x665 &  x674 &  x680 &  x689 &  x692 &  x701 &  x704 &  x710 &  x713 &  x716 &  x719 &  x721 &  x722 &  x725 &  x734 &  x739 &  x740 &  x749 &  x758 &  x760 &  x761 &  x770 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x815 &  x818 &  x827 &  x830 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x872 &  x878 &  x881 &  x884 &  x890 &  x896 &  x899 &  x908 &  x911 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x971 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1058 &  x1061 &  x1073 &  x1076 &  x1088 &  x1103 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 & ~x546 & ~x624 & ~x663 & ~x702 & ~x741 & ~x819 & ~x858;
assign c0126 =  x5 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x56 &  x59 &  x65 &  x74 &  x77 &  x80 &  x89 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x122 &  x125 &  x128 &  x134 &  x137 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x188 &  x191 &  x194 &  x197 &  x203 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x287 &  x296 &  x299 &  x302 &  x305 &  x311 &  x323 &  x326 &  x332 &  x335 &  x338 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x371 &  x377 &  x380 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x437 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x467 &  x469 &  x470 &  x473 &  x482 &  x485 &  x488 &  x491 &  x494 &  x503 &  x506 &  x507 &  x509 &  x512 &  x515 &  x524 &  x530 &  x536 &  x539 &  x542 &  x547 &  x551 &  x557 &  x560 &  x569 &  x572 &  x575 &  x581 &  x584 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x611 &  x617 &  x620 &  x623 &  x625 &  x638 &  x644 &  x650 &  x653 &  x665 &  x674 &  x683 &  x686 &  x689 &  x692 &  x698 &  x701 &  x704 &  x707 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x742 &  x743 &  x749 &  x752 &  x755 &  x764 &  x767 &  x770 &  x773 &  x776 &  x782 &  x785 &  x788 &  x791 &  x797 &  x809 &  x815 &  x818 &  x820 &  x821 &  x824 &  x827 &  x842 &  x848 &  x851 &  x854 &  x857 &  x859 &  x860 &  x863 &  x866 &  x875 &  x878 &  x881 &  x887 &  x898 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x929 &  x932 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x976 &  x977 &  x979 &  x980 &  x986 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1046 &  x1049 &  x1052 &  x1055 &  x1057 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1094 &  x1103 &  x1109 &  x1115 &  x1118 &  x1121 &  x1127 & ~x393 & ~x432 & ~x453 & ~x486 & ~x552 & ~x630 & ~x669;
assign c0128 =  x11 &  x17 &  x20 &  x26 &  x32 &  x35 &  x38 &  x43 &  x47 &  x53 &  x56 &  x62 &  x77 &  x83 &  x86 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x122 &  x125 &  x137 &  x140 &  x143 &  x146 &  x149 &  x155 &  x161 &  x164 &  x176 &  x179 &  x182 &  x185 &  x194 &  x197 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x224 &  x239 &  x248 &  x251 &  x254 &  x260 &  x269 &  x275 &  x278 &  x281 &  x287 &  x290 &  x314 &  x317 &  x320 &  x323 &  x329 &  x338 &  x341 &  x344 &  x356 &  x359 &  x362 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x404 &  x407 &  x419 &  x437 &  x440 &  x452 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x491 &  x503 &  x506 &  x509 &  x512 &  x515 &  x527 &  x530 &  x533 &  x536 &  x548 &  x560 &  x566 &  x569 &  x572 &  x575 &  x584 &  x587 &  x590 &  x599 &  x602 &  x611 &  x617 &  x629 &  x632 &  x647 &  x650 &  x662 &  x664 &  x665 &  x667 &  x674 &  x677 &  x680 &  x686 &  x689 &  x698 &  x701 &  x707 &  x713 &  x716 &  x719 &  x722 &  x731 &  x734 &  x740 &  x742 &  x743 &  x745 &  x746 &  x752 &  x755 &  x761 &  x767 &  x773 &  x776 &  x779 &  x781 &  x788 &  x797 &  x800 &  x803 &  x812 &  x815 &  x818 &  x821 &  x823 &  x827 &  x830 &  x836 &  x839 &  x842 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x893 &  x896 &  x898 &  x902 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x937 &  x941 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x980 &  x986 &  x989 &  x995 &  x1015 &  x1016 &  x1022 &  x1025 &  x1031 &  x1037 &  x1043 &  x1049 &  x1052 &  x1054 &  x1064 &  x1067 &  x1076 &  x1082 &  x1088 &  x1091 &  x1093 &  x1096 &  x1109 &  x1112 &  x1115 &  x1121 & ~x162 & ~x219 & ~x258 & ~x330 & ~x648;
assign c0130 =  x14 &  x17 &  x20 &  x26 &  x50 &  x53 &  x71 &  x77 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x122 &  x128 &  x131 &  x134 &  x143 &  x152 &  x155 &  x158 &  x161 &  x167 &  x179 &  x182 &  x188 &  x197 &  x209 &  x212 &  x215 &  x224 &  x236 &  x242 &  x254 &  x257 &  x266 &  x269 &  x275 &  x284 &  x287 &  x290 &  x293 &  x296 &  x302 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x389 &  x392 &  x395 &  x404 &  x407 &  x410 &  x413 &  x433 &  x434 &  x437 &  x443 &  x452 &  x455 &  x461 &  x464 &  x472 &  x473 &  x479 &  x482 &  x491 &  x500 &  x503 &  x511 &  x515 &  x518 &  x521 &  x527 &  x530 &  x536 &  x539 &  x548 &  x557 &  x560 &  x575 &  x578 &  x584 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x614 &  x626 &  x632 &  x635 &  x641 &  x647 &  x650 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x682 &  x683 &  x692 &  x695 &  x701 &  x707 &  x710 &  x713 &  x716 &  x719 &  x721 &  x730 &  x731 &  x740 &  x743 &  x749 &  x758 &  x760 &  x761 &  x770 &  x773 &  x776 &  x782 &  x788 &  x791 &  x794 &  x797 &  x799 &  x800 &  x806 &  x808 &  x809 &  x812 &  x818 &  x833 &  x838 &  x842 &  x845 &  x847 &  x848 &  x854 &  x856 &  x857 &  x860 &  x869 &  x877 &  x890 &  x893 &  x896 &  x902 &  x905 &  x911 &  x914 &  x917 &  x923 &  x929 &  x932 &  x935 &  x938 &  x941 &  x943 &  x944 &  x950 &  x953 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x986 &  x995 &  x1001 &  x1007 &  x1013 &  x1016 &  x1022 &  x1025 &  x1027 &  x1028 &  x1031 &  x1033 &  x1034 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1061 &  x1066 &  x1073 &  x1076 &  x1079 &  x1085 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1121 &  x1124 & ~x240 & ~x279;
assign c0132 =  x2 &  x8 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x41 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x71 &  x74 &  x77 &  x83 &  x86 &  x95 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x131 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x185 &  x188 &  x194 &  x197 &  x200 &  x203 &  x209 &  x212 &  x218 &  x221 &  x224 &  x227 &  x230 &  x236 &  x239 &  x242 &  x248 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x332 &  x335 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x365 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x488 &  x494 &  x500 &  x503 &  x506 &  x508 &  x521 &  x524 &  x530 &  x533 &  x542 &  x545 &  x547 &  x548 &  x551 &  x560 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x586 &  x587 &  x590 &  x596 &  x599 &  x602 &  x605 &  x611 &  x617 &  x620 &  x625 &  x626 &  x629 &  x632 &  x641 &  x644 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x680 &  x683 &  x686 &  x689 &  x695 &  x698 &  x701 &  x704 &  x707 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x737 &  x740 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x758 &  x764 &  x767 &  x776 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x806 &  x809 &  x812 &  x818 &  x821 &  x824 &  x833 &  x836 &  x839 &  x845 &  x848 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x869 &  x875 &  x878 &  x884 &  x887 &  x890 &  x896 &  x899 &  x901 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x944 &  x947 &  x953 &  x956 &  x959 &  x962 &  x965 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x33 & ~x72 & ~x339 & ~x474 & ~x513 & ~x552 & ~x660 & ~x699 & ~x738 & ~x777;
assign c0134 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x191 &  x194 &  x197 &  x200 &  x203 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x293 &  x296 &  x302 &  x305 &  x308 &  x314 &  x317 &  x320 &  x323 &  x326 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x400 &  x401 &  x404 &  x407 &  x413 &  x416 &  x422 &  x431 &  x434 &  x439 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x470 &  x473 &  x476 &  x479 &  x481 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x506 &  x508 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x546 &  x547 &  x554 &  x557 &  x560 &  x563 &  x566 &  x572 &  x575 &  x578 &  x581 &  x584 &  x585 &  x586 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x624 &  x625 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x742 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x781 &  x782 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x820 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x857 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x898 &  x899 &  x901 &  x902 &  x905 &  x908 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x940 &  x941 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 & ~x525 & ~x564;
assign c0136 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x53 &  x59 &  x68 &  x71 &  x74 &  x80 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x119 &  x122 &  x128 &  x131 &  x137 &  x143 &  x146 &  x152 &  x155 &  x158 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x197 &  x203 &  x206 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x236 &  x239 &  x242 &  x248 &  x251 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x326 &  x329 &  x338 &  x341 &  x344 &  x347 &  x351 &  x352 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x389 &  x390 &  x392 &  x395 &  x398 &  x404 &  x407 &  x410 &  x413 &  x416 &  x425 &  x428 &  x430 &  x431 &  x434 &  x437 &  x443 &  x446 &  x449 &  x452 &  x458 &  x461 &  x469 &  x476 &  x479 &  x482 &  x488 &  x491 &  x494 &  x497 &  x500 &  x508 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x542 &  x545 &  x547 &  x551 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x587 &  x590 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x620 &  x623 &  x626 &  x629 &  x638 &  x641 &  x644 &  x647 &  x650 &  x656 &  x659 &  x662 &  x665 &  x667 &  x668 &  x674 &  x677 &  x680 &  x683 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x706 &  x707 &  x713 &  x716 &  x719 &  x728 &  x734 &  x737 &  x743 &  x746 &  x749 &  x752 &  x758 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x788 &  x791 &  x794 &  x797 &  x806 &  x809 &  x812 &  x815 &  x818 &  x824 &  x827 &  x830 &  x833 &  x839 &  x848 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x887 &  x890 &  x893 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1016 &  x1022 &  x1025 &  x1027 &  x1028 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1061 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1118 &  x1121 &  x1124 & ~x342 & ~x375 & ~x516 & ~x780 & ~x819;
assign c0138 =  x5 &  x8 &  x11 &  x14 &  x17 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x56 &  x59 &  x62 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x167 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x209 &  x215 &  x218 &  x221 &  x227 &  x230 &  x233 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x302 &  x305 &  x308 &  x314 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x341 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x389 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x437 &  x440 &  x446 &  x452 &  x455 &  x458 &  x461 &  x467 &  x470 &  x473 &  x476 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x506 &  x509 &  x515 &  x518 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x589 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x623 &  x626 &  x628 &  x629 &  x635 &  x638 &  x647 &  x650 &  x656 &  x659 &  x662 &  x667 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x731 &  x737 &  x743 &  x745 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x773 &  x779 &  x783 &  x784 &  x785 &  x788 &  x791 &  x794 &  x800 &  x803 &  x806 &  x812 &  x815 &  x821 &  x823 &  x824 &  x836 &  x839 &  x842 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x881 &  x884 &  x893 &  x896 &  x902 &  x905 &  x908 &  x911 &  x916 &  x917 &  x920 &  x926 &  x929 &  x932 &  x938 &  x940 &  x941 &  x944 &  x950 &  x953 &  x955 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x977 &  x983 &  x992 &  x994 &  x1001 &  x1004 &  x1007 &  x1013 &  x1016 &  x1028 &  x1031 &  x1032 &  x1034 &  x1037 &  x1043 &  x1049 &  x1052 &  x1055 &  x1058 &  x1067 &  x1072 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1090 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1124 &  x1127 &  x1130;
assign c0140 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x41 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x92 &  x98 &  x101 &  x104 &  x107 &  x110 &  x116 &  x119 &  x122 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x179 &  x182 &  x188 &  x197 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x251 &  x254 &  x266 &  x269 &  x272 &  x281 &  x284 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x377 &  x380 &  x386 &  x389 &  x391 &  x392 &  x395 &  x398 &  x401 &  x407 &  x413 &  x416 &  x419 &  x425 &  x430 &  x437 &  x440 &  x443 &  x449 &  x452 &  x455 &  x464 &  x467 &  x473 &  x476 &  x479 &  x488 &  x491 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x530 &  x533 &  x536 &  x539 &  x542 &  x548 &  x551 &  x554 &  x557 &  x560 &  x566 &  x569 &  x572 &  x578 &  x581 &  x584 &  x587 &  x593 &  x599 &  x602 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x641 &  x644 &  x647 &  x650 &  x656 &  x659 &  x665 &  x667 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x722 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x745 &  x746 &  x749 &  x752 &  x761 &  x764 &  x767 &  x770 &  x776 &  x779 &  x784 &  x785 &  x788 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x830 &  x833 &  x836 &  x839 &  x845 &  x851 &  x854 &  x857 &  x863 &  x869 &  x872 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x938 &  x944 &  x953 &  x956 &  x959 &  x962 &  x968 &  x971 &  x974 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1049 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x177 & ~x318 & ~x357 & ~x396 & ~x435 & ~x474 & ~x480 & ~x513 & ~x519 & ~x558 & ~x1041 & ~x1080;
assign c0142 =  x2 &  x8 &  x11 &  x14 &  x17 &  x23 &  x26 &  x32 &  x35 &  x41 &  x53 &  x56 &  x62 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x92 &  x95 &  x101 &  x107 &  x110 &  x113 &  x116 &  x119 &  x128 &  x131 &  x134 &  x143 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x170 &  x179 &  x181 &  x182 &  x185 &  x188 &  x191 &  x194 &  x203 &  x206 &  x209 &  x212 &  x218 &  x220 &  x226 &  x230 &  x233 &  x236 &  x242 &  x245 &  x251 &  x254 &  x257 &  x260 &  x263 &  x265 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x298 &  x299 &  x302 &  x305 &  x311 &  x314 &  x320 &  x323 &  x329 &  x332 &  x335 &  x337 &  x338 &  x344 &  x350 &  x359 &  x368 &  x370 &  x371 &  x374 &  x380 &  x383 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x419 &  x422 &  x434 &  x437 &  x446 &  x449 &  x455 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x485 &  x494 &  x497 &  x503 &  x509 &  x512 &  x530 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x566 &  x572 &  x581 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x614 &  x623 &  x629 &  x632 &  x635 &  x638 &  x644 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x677 &  x680 &  x683 &  x689 &  x692 &  x695 &  x698 &  x713 &  x716 &  x719 &  x722 &  x728 &  x734 &  x737 &  x740 &  x742 &  x743 &  x745 &  x746 &  x755 &  x758 &  x764 &  x770 &  x776 &  x779 &  x781 &  x782 &  x784 &  x785 &  x788 &  x791 &  x797 &  x803 &  x818 &  x821 &  x823 &  x830 &  x833 &  x839 &  x851 &  x854 &  x857 &  x859 &  x862 &  x863 &  x866 &  x878 &  x881 &  x890 &  x896 &  x898 &  x899 &  x900 &  x901 &  x902 &  x905 &  x908 &  x911 &  x920 &  x923 &  x929 &  x935 &  x937 &  x939 &  x940 &  x944 &  x947 &  x950 &  x953 &  x956 &  x965 &  x968 &  x971 &  x974 &  x976 &  x978 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1018 &  x1022 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1056 &  x1057 &  x1058 &  x1067 &  x1082 &  x1085 &  x1095 &  x1096 &  x1097 &  x1100 &  x1106 &  x1109 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x273 & ~x312 & ~x351 & ~x471 & ~x510;
assign c0144 =  x16 &  x32 &  x38 &  x41 &  x47 &  x50 &  x55 &  x59 &  x106 &  x113 &  x116 &  x122 &  x125 &  x131 &  x144 &  x155 &  x197 &  x209 &  x212 &  x260 &  x281 &  x289 &  x290 &  x293 &  x296 &  x299 &  x302 &  x320 &  x328 &  x338 &  x344 &  x347 &  x350 &  x353 &  x356 &  x365 &  x371 &  x389 &  x395 &  x413 &  x431 &  x443 &  x488 &  x494 &  x497 &  x512 &  x518 &  x524 &  x527 &  x536 &  x539 &  x542 &  x554 &  x557 &  x562 &  x563 &  x578 &  x593 &  x602 &  x608 &  x626 &  x629 &  x638 &  x640 &  x644 &  x659 &  x662 &  x668 &  x671 &  x692 &  x734 &  x742 &  x752 &  x755 &  x757 &  x758 &  x767 &  x782 &  x785 &  x809 &  x818 &  x824 &  x833 &  x854 &  x859 &  x905 &  x908 &  x914 &  x932 &  x937 &  x944 &  x953 &  x956 &  x962 &  x971 &  x983 &  x986 &  x992 &  x1010 &  x1013 &  x1019 &  x1025 &  x1034 &  x1040 &  x1055 &  x1064 &  x1067 &  x1079 &  x1085 &  x1091 &  x1093 &  x1097 &  x1103 &  x1121 &  x1127 & ~x237 & ~x276 & ~x315 & ~x432 & ~x708 & ~x825 & ~x903;
assign c0146 =  x5 &  x8 &  x17 &  x26 &  x32 &  x35 &  x38 &  x44 &  x47 &  x53 &  x56 &  x59 &  x65 &  x68 &  x74 &  x86 &  x98 &  x104 &  x107 &  x119 &  x125 &  x128 &  x131 &  x134 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x167 &  x170 &  x185 &  x188 &  x200 &  x206 &  x212 &  x215 &  x218 &  x227 &  x230 &  x233 &  x245 &  x248 &  x254 &  x260 &  x269 &  x275 &  x278 &  x281 &  x287 &  x299 &  x302 &  x305 &  x320 &  x326 &  x335 &  x341 &  x353 &  x356 &  x377 &  x383 &  x389 &  x398 &  x401 &  x404 &  x407 &  x413 &  x419 &  x422 &  x425 &  x430 &  x434 &  x437 &  x446 &  x452 &  x458 &  x464 &  x467 &  x470 &  x472 &  x473 &  x476 &  x479 &  x482 &  x485 &  x491 &  x500 &  x503 &  x506 &  x511 &  x524 &  x527 &  x536 &  x539 &  x542 &  x545 &  x548 &  x550 &  x551 &  x557 &  x563 &  x566 &  x569 &  x572 &  x575 &  x584 &  x587 &  x590 &  x593 &  x599 &  x602 &  x614 &  x628 &  x632 &  x635 &  x641 &  x644 &  x650 &  x662 &  x665 &  x668 &  x671 &  x677 &  x683 &  x689 &  x695 &  x701 &  x706 &  x707 &  x710 &  x716 &  x722 &  x743 &  x752 &  x755 &  x761 &  x764 &  x767 &  x770 &  x782 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x824 &  x827 &  x830 &  x833 &  x836 &  x842 &  x845 &  x860 &  x866 &  x869 &  x872 &  x877 &  x878 &  x890 &  x893 &  x896 &  x899 &  x905 &  x908 &  x911 &  x914 &  x923 &  x935 &  x941 &  x950 &  x959 &  x968 &  x974 &  x977 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1010 &  x1016 &  x1019 &  x1025 &  x1034 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1061 &  x1082 &  x1088 &  x1100 &  x1106 &  x1112 &  x1118 &  x1124 &  x1130 & ~x138 & ~x178 & ~x702 & ~x741;
assign c0148 =  x2 &  x8 &  x11 &  x14 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x41 &  x43 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x80 &  x83 &  x89 &  x92 &  x101 &  x104 &  x107 &  x116 &  x119 &  x122 &  x125 &  x137 &  x146 &  x149 &  x155 &  x173 &  x182 &  x194 &  x197 &  x212 &  x218 &  x224 &  x227 &  x230 &  x242 &  x245 &  x251 &  x254 &  x260 &  x263 &  x278 &  x281 &  x284 &  x299 &  x302 &  x308 &  x311 &  x314 &  x317 &  x326 &  x329 &  x338 &  x341 &  x353 &  x355 &  x359 &  x362 &  x365 &  x374 &  x380 &  x383 &  x392 &  x394 &  x395 &  x398 &  x407 &  x410 &  x413 &  x425 &  x428 &  x431 &  x434 &  x440 &  x443 &  x458 &  x470 &  x473 &  x488 &  x500 &  x506 &  x512 &  x518 &  x524 &  x527 &  x548 &  x550 &  x551 &  x554 &  x557 &  x560 &  x563 &  x575 &  x587 &  x589 &  x590 &  x599 &  x605 &  x611 &  x617 &  x623 &  x626 &  x628 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x656 &  x662 &  x671 &  x674 &  x677 &  x683 &  x686 &  x692 &  x701 &  x707 &  x710 &  x713 &  x719 &  x725 &  x731 &  x737 &  x745 &  x748 &  x749 &  x758 &  x761 &  x764 &  x767 &  x773 &  x776 &  x785 &  x787 &  x797 &  x800 &  x803 &  x812 &  x815 &  x818 &  x821 &  x827 &  x830 &  x845 &  x848 &  x851 &  x854 &  x857 &  x866 &  x869 &  x872 &  x878 &  x881 &  x884 &  x887 &  x890 &  x908 &  x914 &  x920 &  x932 &  x935 &  x938 &  x944 &  x953 &  x956 &  x959 &  x965 &  x971 &  x977 &  x980 &  x986 &  x992 &  x995 &  x998 &  x1016 &  x1021 &  x1022 &  x1025 &  x1027 &  x1043 &  x1049 &  x1055 &  x1058 &  x1064 &  x1073 &  x1076 &  x1082 &  x1085 &  x1103 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130 & ~x1122;
assign c0150 =  x5 &  x8 &  x14 &  x20 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x50 &  x53 &  x56 &  x65 &  x68 &  x74 &  x77 &  x80 &  x86 &  x95 &  x98 &  x107 &  x110 &  x119 &  x125 &  x128 &  x131 &  x134 &  x140 &  x146 &  x152 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x182 &  x188 &  x203 &  x206 &  x209 &  x212 &  x233 &  x251 &  x254 &  x263 &  x269 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x302 &  x308 &  x311 &  x317 &  x332 &  x338 &  x344 &  x347 &  x350 &  x353 &  x356 &  x368 &  x371 &  x377 &  x380 &  x392 &  x407 &  x416 &  x419 &  x425 &  x428 &  x434 &  x437 &  x443 &  x449 &  x452 &  x455 &  x461 &  x464 &  x467 &  x481 &  x482 &  x485 &  x494 &  x500 &  x503 &  x506 &  x512 &  x518 &  x521 &  x524 &  x539 &  x542 &  x545 &  x554 &  x560 &  x563 &  x566 &  x569 &  x575 &  x578 &  x581 &  x584 &  x590 &  x596 &  x608 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x641 &  x644 &  x647 &  x653 &  x665 &  x668 &  x671 &  x674 &  x680 &  x683 &  x686 &  x698 &  x710 &  x719 &  x737 &  x740 &  x746 &  x755 &  x758 &  x767 &  x770 &  x773 &  x776 &  x779 &  x788 &  x791 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x842 &  x845 &  x851 &  x854 &  x860 &  x863 &  x878 &  x881 &  x884 &  x887 &  x897 &  x901 &  x905 &  x908 &  x911 &  x917 &  x923 &  x929 &  x932 &  x936 &  x937 &  x938 &  x940 &  x941 &  x956 &  x959 &  x968 &  x971 &  x974 &  x977 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1014 &  x1015 &  x1028 &  x1037 &  x1043 &  x1053 &  x1055 &  x1057 &  x1061 &  x1067 &  x1070 &  x1076 &  x1079 &  x1088 &  x1092 &  x1093 &  x1094 &  x1097 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 & ~x351 & ~x708 & ~x987;
assign c0152 =  x2 &  x11 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x50 &  x59 &  x74 &  x77 &  x80 &  x82 &  x89 &  x104 &  x110 &  x113 &  x119 &  x121 &  x122 &  x125 &  x137 &  x156 &  x158 &  x160 &  x164 &  x170 &  x173 &  x179 &  x182 &  x185 &  x188 &  x194 &  x199 &  x200 &  x203 &  x206 &  x209 &  x221 &  x224 &  x227 &  x230 &  x233 &  x234 &  x238 &  x245 &  x248 &  x254 &  x257 &  x263 &  x266 &  x269 &  x272 &  x274 &  x278 &  x284 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x311 &  x316 &  x320 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x355 &  x371 &  x374 &  x377 &  x383 &  x386 &  x389 &  x398 &  x401 &  x410 &  x413 &  x416 &  x419 &  x428 &  x431 &  x433 &  x440 &  x446 &  x449 &  x455 &  x458 &  x473 &  x476 &  x479 &  x485 &  x488 &  x491 &  x497 &  x500 &  x503 &  x509 &  x512 &  x524 &  x527 &  x545 &  x551 &  x553 &  x554 &  x557 &  x563 &  x566 &  x575 &  x578 &  x581 &  x590 &  x593 &  x596 &  x599 &  x602 &  x604 &  x617 &  x620 &  x626 &  x629 &  x632 &  x638 &  x640 &  x642 &  x644 &  x647 &  x650 &  x653 &  x662 &  x665 &  x668 &  x671 &  x674 &  x689 &  x695 &  x704 &  x716 &  x722 &  x737 &  x740 &  x743 &  x746 &  x755 &  x758 &  x760 &  x764 &  x767 &  x779 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x812 &  x818 &  x821 &  x824 &  x827 &  x833 &  x836 &  x839 &  x845 &  x848 &  x851 &  x854 &  x863 &  x869 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x905 &  x908 &  x914 &  x920 &  x935 &  x941 &  x947 &  x950 &  x953 &  x956 &  x962 &  x968 &  x983 &  x986 &  x989 &  x1022 &  x1025 &  x1028 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1088 &  x1091 &  x1097 &  x1103 &  x1112 &  x1115 &  x1118 &  x1121 &  x1130 & ~x819;
assign c0154 =  x2 &  x17 &  x20 &  x23 &  x29 &  x35 &  x38 &  x41 &  x44 &  x53 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x92 &  x98 &  x101 &  x110 &  x113 &  x116 &  x119 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x152 &  x158 &  x167 &  x170 &  x176 &  x179 &  x185 &  x188 &  x203 &  x206 &  x212 &  x215 &  x218 &  x221 &  x224 &  x236 &  x242 &  x245 &  x248 &  x251 &  x257 &  x260 &  x263 &  x266 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x293 &  x296 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x329 &  x335 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x365 &  x371 &  x374 &  x377 &  x380 &  x383 &  x389 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x449 &  x458 &  x467 &  x476 &  x479 &  x482 &  x485 &  x488 &  x494 &  x497 &  x503 &  x506 &  x508 &  x509 &  x521 &  x527 &  x530 &  x533 &  x542 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x584 &  x586 &  x587 &  x589 &  x593 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x623 &  x626 &  x628 &  x641 &  x647 &  x650 &  x653 &  x655 &  x659 &  x662 &  x665 &  x667 &  x668 &  x680 &  x683 &  x686 &  x692 &  x698 &  x701 &  x707 &  x710 &  x716 &  x719 &  x725 &  x728 &  x734 &  x737 &  x740 &  x745 &  x746 &  x755 &  x758 &  x764 &  x767 &  x770 &  x773 &  x776 &  x782 &  x788 &  x794 &  x797 &  x800 &  x803 &  x806 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x830 &  x833 &  x842 &  x845 &  x848 &  x857 &  x860 &  x862 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x893 &  x896 &  x899 &  x901 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x935 &  x938 &  x940 &  x944 &  x947 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x980 &  x986 &  x989 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1022 &  x1025 &  x1028 &  x1034 &  x1037 &  x1040 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1118 &  x1121 &  x1127 & ~x474 & ~x555 & ~x594 & ~x816;
assign c0156 =  x2 &  x11 &  x29 &  x41 &  x44 &  x50 &  x56 &  x83 &  x92 &  x98 &  x101 &  x104 &  x131 &  x143 &  x149 &  x158 &  x164 &  x176 &  x179 &  x185 &  x188 &  x206 &  x209 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x239 &  x251 &  x257 &  x260 &  x269 &  x272 &  x275 &  x278 &  x284 &  x287 &  x290 &  x296 &  x302 &  x305 &  x308 &  x314 &  x323 &  x335 &  x341 &  x344 &  x353 &  x356 &  x368 &  x377 &  x380 &  x392 &  x395 &  x407 &  x419 &  x422 &  x425 &  x428 &  x434 &  x437 &  x449 &  x461 &  x467 &  x472 &  x476 &  x479 &  x497 &  x503 &  x506 &  x512 &  x530 &  x542 &  x545 &  x551 &  x554 &  x560 &  x566 &  x581 &  x590 &  x602 &  x605 &  x614 &  x617 &  x627 &  x628 &  x629 &  x635 &  x647 &  x650 &  x653 &  x662 &  x665 &  x666 &  x667 &  x668 &  x680 &  x686 &  x692 &  x705 &  x706 &  x710 &  x728 &  x740 &  x743 &  x745 &  x752 &  x755 &  x764 &  x767 &  x782 &  x784 &  x791 &  x800 &  x803 &  x824 &  x827 &  x836 &  x839 &  x848 &  x851 &  x863 &  x869 &  x872 &  x875 &  x881 &  x893 &  x896 &  x899 &  x902 &  x908 &  x917 &  x923 &  x932 &  x938 &  x950 &  x956 &  x962 &  x968 &  x983 &  x988 &  x998 &  x1004 &  x1019 &  x1025 &  x1026 &  x1034 &  x1052 &  x1061 &  x1079 &  x1082 &  x1088 &  x1103 &  x1121 &  x1127 &  x1130;
assign c0158 =  x2 &  x8 &  x11 &  x14 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x50 &  x65 &  x71 &  x74 &  x83 &  x86 &  x98 &  x101 &  x116 &  x117 &  x118 &  x119 &  x137 &  x143 &  x146 &  x155 &  x157 &  x158 &  x160 &  x161 &  x170 &  x173 &  x182 &  x185 &  x191 &  x197 &  x203 &  x206 &  x209 &  x212 &  x215 &  x227 &  x234 &  x235 &  x238 &  x245 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x274 &  x275 &  x278 &  x281 &  x284 &  x293 &  x296 &  x299 &  x305 &  x308 &  x311 &  x313 &  x317 &  x320 &  x323 &  x329 &  x332 &  x335 &  x341 &  x352 &  x359 &  x362 &  x365 &  x371 &  x374 &  x380 &  x383 &  x386 &  x392 &  x394 &  x401 &  x404 &  x407 &  x416 &  x419 &  x425 &  x437 &  x440 &  x455 &  x464 &  x470 &  x472 &  x482 &  x485 &  x488 &  x503 &  x515 &  x533 &  x548 &  x554 &  x557 &  x563 &  x566 &  x578 &  x584 &  x587 &  x590 &  x599 &  x602 &  x604 &  x605 &  x608 &  x620 &  x623 &  x629 &  x635 &  x647 &  x650 &  x656 &  x662 &  x665 &  x668 &  x674 &  x679 &  x682 &  x686 &  x689 &  x692 &  x701 &  x709 &  x710 &  x713 &  x716 &  x718 &  x719 &  x721 &  x725 &  x731 &  x743 &  x748 &  x749 &  x761 &  x764 &  x770 &  x776 &  x779 &  x782 &  x788 &  x791 &  x796 &  x797 &  x799 &  x800 &  x803 &  x809 &  x812 &  x815 &  x821 &  x824 &  x838 &  x839 &  x845 &  x851 &  x854 &  x860 &  x866 &  x875 &  x878 &  x881 &  x884 &  x890 &  x902 &  x904 &  x905 &  x908 &  x914 &  x916 &  x917 &  x920 &  x923 &  x935 &  x938 &  x941 &  x943 &  x950 &  x953 &  x965 &  x968 &  x971 &  x974 &  x983 &  x986 &  x989 &  x998 &  x1004 &  x1007 &  x1019 &  x1040 &  x1046 &  x1055 &  x1058 &  x1067 &  x1073 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1106 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 & ~x939;
assign c0160 =  x2 &  x5 &  x8 &  x14 &  x17 &  x23 &  x29 &  x35 &  x38 &  x41 &  x50 &  x53 &  x68 &  x71 &  x74 &  x77 &  x83 &  x86 &  x89 &  x98 &  x101 &  x104 &  x107 &  x113 &  x116 &  x122 &  x125 &  x131 &  x143 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x176 &  x179 &  x182 &  x185 &  x191 &  x197 &  x200 &  x206 &  x218 &  x227 &  x233 &  x248 &  x251 &  x254 &  x260 &  x263 &  x266 &  x272 &  x275 &  x281 &  x284 &  x290 &  x293 &  x299 &  x305 &  x308 &  x311 &  x320 &  x326 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x356 &  x362 &  x368 &  x374 &  x377 &  x383 &  x389 &  x394 &  x410 &  x413 &  x425 &  x428 &  x430 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x458 &  x461 &  x464 &  x470 &  x472 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x497 &  x500 &  x503 &  x518 &  x527 &  x533 &  x536 &  x542 &  x545 &  x548 &  x550 &  x551 &  x554 &  x560 &  x563 &  x569 &  x575 &  x581 &  x584 &  x590 &  x599 &  x605 &  x614 &  x617 &  x628 &  x632 &  x638 &  x650 &  x653 &  x656 &  x665 &  x667 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x689 &  x692 &  x695 &  x698 &  x701 &  x706 &  x710 &  x713 &  x716 &  x725 &  x728 &  x731 &  x734 &  x737 &  x743 &  x745 &  x749 &  x754 &  x755 &  x761 &  x767 &  x770 &  x773 &  x779 &  x784 &  x785 &  x788 &  x793 &  x797 &  x800 &  x803 &  x806 &  x812 &  x815 &  x818 &  x823 &  x824 &  x827 &  x830 &  x831 &  x833 &  x836 &  x839 &  x842 &  x845 &  x863 &  x866 &  x869 &  x871 &  x872 &  x877 &  x884 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x911 &  x914 &  x916 &  x917 &  x920 &  x923 &  x926 &  x929 &  x935 &  x938 &  x941 &  x947 &  x953 &  x955 &  x962 &  x974 &  x977 &  x983 &  x986 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1031 &  x1034 &  x1037 &  x1043 &  x1064 &  x1067 &  x1070 &  x1072 &  x1076 &  x1079 &  x1082 &  x1088 &  x1094 &  x1100 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1129 & ~x663 & ~x780 & ~x819;
assign c0162 =  x5 &  x8 &  x20 &  x23 &  x26 &  x32 &  x38 &  x41 &  x47 &  x53 &  x59 &  x68 &  x71 &  x74 &  x89 &  x92 &  x95 &  x101 &  x104 &  x107 &  x110 &  x113 &  x125 &  x131 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x161 &  x164 &  x167 &  x170 &  x176 &  x179 &  x182 &  x185 &  x191 &  x194 &  x197 &  x200 &  x209 &  x215 &  x218 &  x224 &  x230 &  x233 &  x239 &  x242 &  x248 &  x251 &  x254 &  x260 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x293 &  x302 &  x305 &  x311 &  x317 &  x320 &  x323 &  x329 &  x332 &  x335 &  x344 &  x350 &  x353 &  x356 &  x368 &  x371 &  x377 &  x380 &  x383 &  x389 &  x395 &  x398 &  x401 &  x404 &  x406 &  x407 &  x410 &  x416 &  x422 &  x425 &  x428 &  x431 &  x449 &  x452 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x488 &  x491 &  x494 &  x500 &  x506 &  x509 &  x518 &  x521 &  x524 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x572 &  x575 &  x578 &  x584 &  x587 &  x590 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x625 &  x626 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x656 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x731 &  x734 &  x737 &  x740 &  x742 &  x743 &  x749 &  x758 &  x761 &  x770 &  x773 &  x779 &  x782 &  x788 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x818 &  x820 &  x821 &  x830 &  x836 &  x842 &  x848 &  x851 &  x854 &  x857 &  x859 &  x860 &  x862 &  x863 &  x866 &  x869 &  x881 &  x884 &  x887 &  x896 &  x898 &  x899 &  x902 &  x908 &  x911 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x937 &  x938 &  x940 &  x941 &  x944 &  x947 &  x950 &  x962 &  x965 &  x968 &  x971 &  x977 &  x979 &  x980 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1018 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1052 &  x1058 &  x1061 &  x1064 &  x1073 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x315 & ~x354 & ~x489 & ~x513 & ~x591 & ~x630 & ~x669 & ~x747 & ~x903;
assign c0164 =  x2 &  x5 &  x8 &  x11 &  x17 &  x23 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x65 &  x68 &  x71 &  x74 &  x77 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x430 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x469 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x511 &  x512 &  x515 &  x518 &  x524 &  x527 &  x533 &  x536 &  x539 &  x545 &  x550 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x589 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130 & ~x69 & ~x186 & ~x852 & ~x855 & ~x891 & ~x930 & ~x969 & ~x1086 & ~x1125;
assign c0166 =  x5 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x35 &  x38 &  x44 &  x53 &  x62 &  x68 &  x74 &  x77 &  x80 &  x86 &  x95 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x122 &  x128 &  x131 &  x134 &  x140 &  x143 &  x155 &  x158 &  x164 &  x170 &  x179 &  x185 &  x188 &  x191 &  x215 &  x218 &  x221 &  x224 &  x230 &  x236 &  x242 &  x248 &  x251 &  x254 &  x263 &  x269 &  x278 &  x281 &  x284 &  x287 &  x293 &  x314 &  x317 &  x323 &  x326 &  x332 &  x344 &  x347 &  x350 &  x356 &  x365 &  x368 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x395 &  x401 &  x404 &  x407 &  x410 &  x416 &  x422 &  x425 &  x434 &  x437 &  x442 &  x443 &  x446 &  x455 &  x467 &  x470 &  x473 &  x485 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x547 &  x551 &  x554 &  x557 &  x560 &  x563 &  x575 &  x581 &  x584 &  x585 &  x587 &  x590 &  x605 &  x608 &  x611 &  x614 &  x620 &  x626 &  x629 &  x632 &  x647 &  x650 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x683 &  x689 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x734 &  x740 &  x743 &  x749 &  x752 &  x758 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x788 &  x803 &  x806 &  x809 &  x818 &  x820 &  x823 &  x842 &  x845 &  x848 &  x854 &  x860 &  x862 &  x863 &  x866 &  x869 &  x875 &  x878 &  x890 &  x893 &  x896 &  x901 &  x902 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x937 &  x938 &  x941 &  x944 &  x947 &  x956 &  x959 &  x962 &  x971 &  x974 &  x976 &  x977 &  x979 &  x989 &  x998 &  x1004 &  x1007 &  x1013 &  x1016 &  x1018 &  x1019 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1052 &  x1055 &  x1064 &  x1067 &  x1070 &  x1073 &  x1085 &  x1088 &  x1094 &  x1097 &  x1103 &  x1106 &  x1115 &  x1124 &  x1127 & ~x525 & ~x564 & ~x603 & ~x630;
assign c0168 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x53 &  x59 &  x65 &  x68 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x113 &  x116 &  x119 &  x122 &  x125 &  x131 &  x134 &  x137 &  x140 &  x146 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x242 &  x245 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x311 &  x313 &  x314 &  x317 &  x320 &  x326 &  x329 &  x335 &  x338 &  x344 &  x347 &  x350 &  x353 &  x356 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x629 &  x635 &  x641 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x707 &  x710 &  x713 &  x716 &  x719 &  x725 &  x728 &  x734 &  x737 &  x743 &  x746 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x772 &  x773 &  x776 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x811 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x950 &  x953 &  x959 &  x965 &  x968 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x994 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1052 &  x1055 &  x1058 &  x1061 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x6 & ~x12 & ~x45 & ~x51 & ~x84 & ~x297 & ~x303 & ~x336 & ~x1059 & ~x1098;
assign c0170 =  x2 &  x23 &  x35 &  x38 &  x47 &  x62 &  x65 &  x74 &  x77 &  x86 &  x89 &  x98 &  x104 &  x110 &  x119 &  x125 &  x131 &  x140 &  x152 &  x158 &  x161 &  x170 &  x176 &  x182 &  x185 &  x188 &  x212 &  x218 &  x227 &  x239 &  x248 &  x260 &  x269 &  x281 &  x284 &  x287 &  x296 &  x299 &  x302 &  x305 &  x308 &  x335 &  x353 &  x359 &  x365 &  x371 &  x392 &  x395 &  x413 &  x425 &  x429 &  x430 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x452 &  x458 &  x469 &  x473 &  x476 &  x482 &  x485 &  x488 &  x494 &  x497 &  x508 &  x511 &  x512 &  x515 &  x545 &  x560 &  x578 &  x587 &  x590 &  x614 &  x617 &  x625 &  x647 &  x653 &  x665 &  x667 &  x668 &  x680 &  x686 &  x689 &  x701 &  x704 &  x705 &  x707 &  x716 &  x719 &  x722 &  x725 &  x742 &  x743 &  x746 &  x764 &  x767 &  x770 &  x784 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x818 &  x821 &  x824 &  x833 &  x845 &  x848 &  x857 &  x863 &  x872 &  x875 &  x878 &  x881 &  x890 &  x902 &  x917 &  x932 &  x938 &  x941 &  x950 &  x953 &  x956 &  x962 &  x986 &  x992 &  x998 &  x1001 &  x1007 &  x1022 &  x1025 &  x1046 &  x1052 &  x1058 &  x1064 &  x1079 &  x1082 &  x1097 &  x1103 &  x1112 &  x1121 &  x1130;
assign c0172 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x469 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x508 &  x509 &  x512 &  x515 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x547 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x625 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x694 &  x695 &  x698 &  x701 &  x703 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x742 &  x743 &  x746 &  x749 &  x752 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x435 & ~x474 & ~x513 & ~x552 & ~x553 & ~x591 & ~x592 & ~x630 & ~x636 & ~x675 & ~x708;
assign c0174 =  x2 &  x5 &  x11 &  x17 &  x20 &  x23 &  x32 &  x41 &  x44 &  x47 &  x53 &  x59 &  x74 &  x77 &  x80 &  x83 &  x92 &  x101 &  x104 &  x107 &  x113 &  x116 &  x119 &  x128 &  x131 &  x134 &  x140 &  x143 &  x146 &  x152 &  x155 &  x161 &  x164 &  x170 &  x173 &  x176 &  x188 &  x191 &  x194 &  x200 &  x203 &  x209 &  x212 &  x215 &  x221 &  x230 &  x233 &  x236 &  x242 &  x245 &  x248 &  x251 &  x260 &  x272 &  x275 &  x278 &  x284 &  x290 &  x308 &  x314 &  x320 &  x323 &  x326 &  x338 &  x341 &  x344 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x380 &  x389 &  x392 &  x398 &  x416 &  x419 &  x425 &  x431 &  x433 &  x434 &  x443 &  x446 &  x455 &  x458 &  x467 &  x485 &  x488 &  x494 &  x497 &  x503 &  x506 &  x509 &  x511 &  x512 &  x515 &  x527 &  x533 &  x536 &  x539 &  x550 &  x557 &  x560 &  x569 &  x572 &  x575 &  x578 &  x581 &  x589 &  x590 &  x593 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x626 &  x628 &  x629 &  x632 &  x635 &  x644 &  x653 &  x656 &  x662 &  x665 &  x666 &  x668 &  x671 &  x677 &  x680 &  x683 &  x692 &  x698 &  x701 &  x705 &  x706 &  x707 &  x713 &  x716 &  x725 &  x728 &  x734 &  x743 &  x745 &  x749 &  x755 &  x758 &  x764 &  x770 &  x779 &  x782 &  x785 &  x797 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x824 &  x830 &  x833 &  x848 &  x850 &  x851 &  x866 &  x872 &  x875 &  x881 &  x883 &  x887 &  x890 &  x893 &  x899 &  x902 &  x908 &  x914 &  x923 &  x926 &  x929 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x962 &  x965 &  x971 &  x977 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1064 &  x1070 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 & ~x306 & ~x600 & ~x663 & ~x702 & ~x819 & ~x858 & ~x936 & ~x975;
assign c0176 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x391 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x429 &  x430 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x469 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x508 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x547 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x625 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x667 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x703 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x742 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x375 & ~x396 & ~x414 & ~x435 & ~x453 & ~x474 & ~x492 & ~x513 & ~x519 & ~x552 & ~x558 & ~x597 & ~x636;
assign c0178 =  x2 &  x5 &  x8 &  x14 &  x17 &  x23 &  x26 &  x29 &  x44 &  x56 &  x59 &  x65 &  x71 &  x74 &  x80 &  x83 &  x86 &  x98 &  x107 &  x110 &  x113 &  x116 &  x122 &  x125 &  x131 &  x140 &  x143 &  x149 &  x152 &  x155 &  x158 &  x161 &  x176 &  x179 &  x182 &  x188 &  x194 &  x200 &  x206 &  x215 &  x221 &  x233 &  x239 &  x251 &  x254 &  x257 &  x275 &  x278 &  x281 &  x284 &  x293 &  x296 &  x305 &  x311 &  x314 &  x317 &  x323 &  x332 &  x335 &  x344 &  x347 &  x350 &  x356 &  x359 &  x362 &  x374 &  x377 &  x380 &  x386 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x428 &  x434 &  x443 &  x446 &  x452 &  x458 &  x464 &  x473 &  x476 &  x479 &  x485 &  x494 &  x506 &  x509 &  x512 &  x515 &  x518 &  x524 &  x533 &  x536 &  x539 &  x548 &  x554 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x596 &  x608 &  x620 &  x623 &  x626 &  x632 &  x635 &  x653 &  x659 &  x662 &  x665 &  x668 &  x677 &  x680 &  x683 &  x689 &  x698 &  x701 &  x704 &  x707 &  x713 &  x716 &  x725 &  x731 &  x737 &  x740 &  x743 &  x746 &  x755 &  x758 &  x761 &  x764 &  x767 &  x779 &  x784 &  x785 &  x794 &  x797 &  x800 &  x806 &  x812 &  x818 &  x820 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x851 &  x854 &  x857 &  x859 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x901 &  x902 &  x908 &  x914 &  x920 &  x926 &  x929 &  x932 &  x935 &  x938 &  x940 &  x944 &  x947 &  x950 &  x953 &  x956 &  x962 &  x965 &  x968 &  x971 &  x976 &  x979 &  x980 &  x986 &  x989 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1018 &  x1022 &  x1025 &  x1037 &  x1043 &  x1046 &  x1052 &  x1058 &  x1067 &  x1070 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1115 &  x1121 &  x1130 & ~x384 & ~x432 & ~x450 & ~x513 & ~x567 & ~x840;
assign c0180 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x227 &  x230 &  x233 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x266 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x437 &  x440 &  x446 &  x452 &  x455 &  x458 &  x461 &  x464 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x503 &  x506 &  x509 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x542 &  x545 &  x548 &  x550 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x627 &  x628 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x667 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x710 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x851 &  x854 &  x857 &  x860 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x902 &  x905 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x977 &  x980 &  x983 &  x986 &  x988 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1019 &  x1025 &  x1027 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1066 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x138 & ~x555 & ~x594 & ~x633 & ~x672 & ~x741 & ~x780 & ~x819 & ~x975 & ~x1014 & ~x1053;
assign c0182 =  x8 &  x11 &  x17 &  x23 &  x26 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x62 &  x68 &  x71 &  x74 &  x77 &  x83 &  x86 &  x89 &  x92 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x124 &  x125 &  x128 &  x131 &  x134 &  x143 &  x158 &  x164 &  x170 &  x173 &  x176 &  x179 &  x185 &  x188 &  x202 &  x203 &  x212 &  x221 &  x230 &  x233 &  x236 &  x241 &  x242 &  x245 &  x251 &  x257 &  x260 &  x263 &  x269 &  x272 &  x278 &  x284 &  x287 &  x299 &  x302 &  x308 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x335 &  x338 &  x350 &  x353 &  x356 &  x362 &  x368 &  x371 &  x380 &  x383 &  x389 &  x392 &  x416 &  x425 &  x428 &  x434 &  x440 &  x443 &  x445 &  x449 &  x452 &  x455 &  x458 &  x470 &  x473 &  x479 &  x491 &  x494 &  x497 &  x503 &  x509 &  x512 &  x527 &  x530 &  x542 &  x554 &  x559 &  x560 &  x563 &  x569 &  x572 &  x575 &  x584 &  x587 &  x596 &  x598 &  x599 &  x602 &  x605 &  x611 &  x614 &  x626 &  x629 &  x632 &  x641 &  x647 &  x656 &  x659 &  x662 &  x664 &  x665 &  x668 &  x671 &  x674 &  x680 &  x683 &  x686 &  x689 &  x695 &  x698 &  x701 &  x703 &  x707 &  x710 &  x716 &  x719 &  x722 &  x725 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x758 &  x761 &  x767 &  x773 &  x776 &  x781 &  x782 &  x785 &  x788 &  x803 &  x815 &  x818 &  x820 &  x821 &  x824 &  x827 &  x830 &  x833 &  x839 &  x845 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x869 &  x878 &  x881 &  x884 &  x887 &  x898 &  x899 &  x901 &  x902 &  x905 &  x908 &  x911 &  x917 &  x920 &  x923 &  x926 &  x935 &  x937 &  x938 &  x940 &  x941 &  x944 &  x947 &  x953 &  x956 &  x959 &  x968 &  x976 &  x980 &  x983 &  x986 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1018 &  x1019 &  x1022 &  x1025 &  x1028 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1061 &  x1064 &  x1070 &  x1073 &  x1085 &  x1091 &  x1094 &  x1096 &  x1106 &  x1124 &  x1127 &  x1130 & ~x432 & ~x471 & ~x687 & ~x726 & ~x765;
assign c0184 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x38 &  x41 &  x44 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x71 &  x74 &  x77 &  x80 &  x83 &  x92 &  x95 &  x101 &  x104 &  x110 &  x113 &  x122 &  x125 &  x128 &  x131 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x182 &  x185 &  x191 &  x194 &  x197 &  x206 &  x209 &  x212 &  x218 &  x221 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x338 &  x341 &  x344 &  x347 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x497 &  x500 &  x503 &  x509 &  x511 &  x512 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x539 &  x545 &  x548 &  x550 &  x551 &  x566 &  x569 &  x572 &  x575 &  x581 &  x584 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x611 &  x614 &  x617 &  x623 &  x632 &  x641 &  x644 &  x647 &  x653 &  x656 &  x659 &  x665 &  x668 &  x671 &  x674 &  x677 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x709 &  x710 &  x713 &  x716 &  x719 &  x722 &  x728 &  x731 &  x734 &  x737 &  x743 &  x746 &  x748 &  x752 &  x755 &  x758 &  x764 &  x767 &  x773 &  x776 &  x779 &  x782 &  x785 &  x797 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x826 &  x827 &  x830 &  x836 &  x839 &  x842 &  x848 &  x857 &  x860 &  x863 &  x866 &  x869 &  x871 &  x875 &  x877 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x905 &  x908 &  x910 &  x914 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x944 &  x947 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x988 &  x992 &  x995 &  x1004 &  x1007 &  x1010 &  x1016 &  x1019 &  x1022 &  x1025 &  x1027 &  x1031 &  x1034 &  x1043 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1066 &  x1067 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1130 & ~x99 & ~x240 & ~x741 & ~x780 & ~x819 & ~x858 & ~x897 & ~x975;
assign c0186 =  x2 &  x11 &  x14 &  x20 &  x26 &  x47 &  x53 &  x59 &  x62 &  x68 &  x83 &  x86 &  x95 &  x101 &  x107 &  x110 &  x113 &  x119 &  x121 &  x122 &  x128 &  x137 &  x140 &  x146 &  x149 &  x156 &  x157 &  x158 &  x160 &  x161 &  x170 &  x191 &  x195 &  x197 &  x203 &  x215 &  x224 &  x227 &  x236 &  x238 &  x254 &  x274 &  x275 &  x278 &  x287 &  x290 &  x293 &  x296 &  x316 &  x317 &  x326 &  x329 &  x335 &  x344 &  x352 &  x355 &  x359 &  x362 &  x365 &  x383 &  x389 &  x392 &  x395 &  x398 &  x407 &  x410 &  x419 &  x422 &  x425 &  x437 &  x443 &  x449 &  x452 &  x476 &  x482 &  x485 &  x488 &  x500 &  x506 &  x515 &  x536 &  x542 &  x545 &  x551 &  x557 &  x572 &  x575 &  x578 &  x587 &  x605 &  x611 &  x620 &  x626 &  x643 &  x644 &  x647 &  x653 &  x656 &  x662 &  x665 &  x677 &  x683 &  x698 &  x704 &  x713 &  x716 &  x719 &  x721 &  x722 &  x731 &  x734 &  x737 &  x740 &  x743 &  x748 &  x749 &  x760 &  x761 &  x770 &  x773 &  x782 &  x791 &  x797 &  x806 &  x812 &  x818 &  x821 &  x830 &  x836 &  x848 &  x851 &  x857 &  x881 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x917 &  x920 &  x926 &  x929 &  x932 &  x938 &  x953 &  x959 &  x989 &  x1007 &  x1016 &  x1025 &  x1031 &  x1040 &  x1043 &  x1046 &  x1052 &  x1058 &  x1073 &  x1079 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 & ~x102 & ~x324 & ~x429 & ~x468 & ~x507 & ~x546 & ~x585 & ~x663 & ~x741 & ~x819;
assign c0188 =  x5 &  x11 &  x14 &  x17 &  x20 &  x26 &  x32 &  x35 &  x38 &  x41 &  x44 &  x50 &  x56 &  x59 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x92 &  x104 &  x110 &  x116 &  x122 &  x125 &  x128 &  x143 &  x152 &  x158 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x185 &  x188 &  x194 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x227 &  x239 &  x242 &  x248 &  x254 &  x257 &  x260 &  x266 &  x269 &  x284 &  x287 &  x293 &  x296 &  x308 &  x311 &  x323 &  x329 &  x335 &  x338 &  x347 &  x353 &  x359 &  x365 &  x368 &  x371 &  x374 &  x383 &  x386 &  x389 &  x392 &  x401 &  x404 &  x410 &  x416 &  x422 &  x425 &  x428 &  x430 &  x431 &  x434 &  x437 &  x440 &  x452 &  x455 &  x458 &  x464 &  x467 &  x468 &  x473 &  x476 &  x479 &  x482 &  x485 &  x491 &  x497 &  x500 &  x509 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x542 &  x545 &  x554 &  x557 &  x563 &  x569 &  x572 &  x586 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x613 &  x620 &  x626 &  x632 &  x647 &  x652 &  x653 &  x659 &  x664 &  x671 &  x674 &  x686 &  x689 &  x692 &  x703 &  x704 &  x707 &  x713 &  x716 &  x728 &  x730 &  x731 &  x737 &  x740 &  x742 &  x746 &  x752 &  x755 &  x761 &  x764 &  x773 &  x781 &  x785 &  x788 &  x791 &  x794 &  x803 &  x806 &  x808 &  x809 &  x812 &  x815 &  x818 &  x820 &  x824 &  x836 &  x848 &  x854 &  x857 &  x859 &  x860 &  x863 &  x866 &  x869 &  x872 &  x878 &  x881 &  x884 &  x887 &  x896 &  x901 &  x902 &  x905 &  x911 &  x914 &  x917 &  x920 &  x929 &  x938 &  x944 &  x947 &  x950 &  x956 &  x959 &  x965 &  x968 &  x974 &  x977 &  x980 &  x983 &  x989 &  x992 &  x1013 &  x1019 &  x1022 &  x1034 &  x1046 &  x1049 &  x1052 &  x1057 &  x1058 &  x1061 &  x1067 &  x1070 &  x1073 &  x1079 &  x1088 &  x1091 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1118 &  x1124 & ~x474 & ~x513 & ~x552 & ~x591;
assign c0190 =  x2 &  x5 &  x8 &  x11 &  x29 &  x32 &  x35 &  x41 &  x44 &  x47 &  x50 &  x56 &  x62 &  x65 &  x68 &  x71 &  x77 &  x80 &  x92 &  x110 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x155 &  x158 &  x164 &  x170 &  x179 &  x191 &  x203 &  x209 &  x212 &  x221 &  x227 &  x230 &  x236 &  x239 &  x254 &  x272 &  x275 &  x281 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x313 &  x320 &  x323 &  x332 &  x350 &  x359 &  x365 &  x371 &  x374 &  x389 &  x392 &  x395 &  x401 &  x404 &  x410 &  x419 &  x425 &  x434 &  x437 &  x440 &  x449 &  x455 &  x461 &  x482 &  x491 &  x494 &  x500 &  x503 &  x509 &  x512 &  x518 &  x521 &  x524 &  x527 &  x539 &  x542 &  x545 &  x548 &  x560 &  x569 &  x575 &  x587 &  x590 &  x602 &  x605 &  x608 &  x611 &  x620 &  x628 &  x629 &  x632 &  x641 &  x647 &  x653 &  x656 &  x662 &  x665 &  x667 &  x668 &  x671 &  x677 &  x683 &  x689 &  x695 &  x704 &  x706 &  x710 &  x716 &  x719 &  x722 &  x731 &  x734 &  x737 &  x745 &  x749 &  x761 &  x764 &  x767 &  x770 &  x776 &  x785 &  x791 &  x794 &  x830 &  x836 &  x839 &  x842 &  x845 &  x851 &  x857 &  x860 &  x866 &  x869 &  x872 &  x875 &  x878 &  x890 &  x896 &  x899 &  x902 &  x908 &  x920 &  x926 &  x932 &  x935 &  x941 &  x944 &  x947 &  x950 &  x962 &  x968 &  x971 &  x974 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1000 &  x1001 &  x1004 &  x1013 &  x1016 &  x1022 &  x1025 &  x1027 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1055 &  x1058 &  x1066 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1103 &  x1106 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x201 & ~x240 & ~x241 & ~x258 & ~x318;
assign c0192 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x35 &  x38 &  x44 &  x47 &  x50 &  x56 &  x62 &  x71 &  x74 &  x77 &  x80 &  x86 &  x92 &  x95 &  x98 &  x101 &  x113 &  x116 &  x119 &  x122 &  x125 &  x131 &  x134 &  x137 &  x143 &  x146 &  x158 &  x167 &  x170 &  x173 &  x176 &  x182 &  x185 &  x194 &  x197 &  x200 &  x203 &  x212 &  x218 &  x221 &  x224 &  x230 &  x233 &  x239 &  x242 &  x251 &  x254 &  x260 &  x263 &  x269 &  x272 &  x275 &  x278 &  x281 &  x287 &  x293 &  x299 &  x302 &  x308 &  x314 &  x320 &  x323 &  x335 &  x341 &  x359 &  x362 &  x368 &  x370 &  x386 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x428 &  x431 &  x434 &  x437 &  x443 &  x445 &  x446 &  x449 &  x452 &  x455 &  x458 &  x467 &  x479 &  x481 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x512 &  x518 &  x521 &  x524 &  x527 &  x536 &  x539 &  x542 &  x548 &  x557 &  x560 &  x566 &  x569 &  x578 &  x581 &  x584 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x611 &  x614 &  x617 &  x620 &  x626 &  x629 &  x638 &  x641 &  x644 &  x650 &  x656 &  x659 &  x662 &  x664 &  x668 &  x671 &  x680 &  x686 &  x689 &  x695 &  x701 &  x703 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x731 &  x734 &  x737 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x781 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x803 &  x806 &  x820 &  x821 &  x824 &  x827 &  x830 &  x836 &  x845 &  x848 &  x851 &  x854 &  x857 &  x859 &  x860 &  x862 &  x863 &  x869 &  x872 &  x875 &  x881 &  x884 &  x890 &  x893 &  x901 &  x902 &  x908 &  x911 &  x914 &  x923 &  x929 &  x932 &  x935 &  x937 &  x938 &  x940 &  x944 &  x947 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x976 &  x977 &  x979 &  x980 &  x986 &  x989 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1018 &  x1022 &  x1031 &  x1037 &  x1040 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1100 &  x1103 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x609 & ~x630 & ~x648 & ~x669 & ~x708 & ~x747 & ~x789 & ~x828;
assign c0194 =  x2 &  x5 &  x29 &  x38 &  x44 &  x53 &  x56 &  x62 &  x65 &  x71 &  x83 &  x89 &  x92 &  x122 &  x131 &  x149 &  x176 &  x194 &  x203 &  x209 &  x212 &  x227 &  x235 &  x245 &  x254 &  x257 &  x263 &  x269 &  x281 &  x299 &  x311 &  x323 &  x329 &  x344 &  x347 &  x356 &  x383 &  x394 &  x419 &  x425 &  x433 &  x446 &  x451 &  x452 &  x458 &  x472 &  x479 &  x482 &  x488 &  x491 &  x497 &  x503 &  x512 &  x518 &  x542 &  x572 &  x590 &  x593 &  x602 &  x620 &  x637 &  x641 &  x668 &  x679 &  x683 &  x686 &  x692 &  x695 &  x698 &  x707 &  x710 &  x715 &  x719 &  x733 &  x737 &  x755 &  x758 &  x767 &  x773 &  x779 &  x785 &  x794 &  x799 &  x800 &  x806 &  x809 &  x812 &  x815 &  x824 &  x836 &  x842 &  x860 &  x875 &  x877 &  x884 &  x889 &  x896 &  x914 &  x920 &  x935 &  x953 &  x974 &  x1004 &  x1022 &  x1025 &  x1031 &  x1037 &  x1046 &  x1073 &  x1076 &  x1079 &  x1082 &  x1088 &  x1115 & ~x984 & ~x1023;
assign c0196 =  x5 &  x8 &  x11 &  x17 &  x32 &  x38 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x80 &  x83 &  x95 &  x98 &  x101 &  x116 &  x119 &  x128 &  x140 &  x149 &  x152 &  x161 &  x176 &  x179 &  x182 &  x185 &  x193 &  x194 &  x200 &  x206 &  x215 &  x218 &  x221 &  x224 &  x230 &  x233 &  x239 &  x254 &  x257 &  x260 &  x287 &  x290 &  x293 &  x296 &  x305 &  x314 &  x320 &  x323 &  x338 &  x344 &  x350 &  x362 &  x365 &  x370 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x401 &  x413 &  x416 &  x419 &  x437 &  x461 &  x464 &  x466 &  x482 &  x485 &  x497 &  x503 &  x506 &  x509 &  x524 &  x530 &  x533 &  x536 &  x548 &  x551 &  x557 &  x572 &  x575 &  x587 &  x608 &  x614 &  x617 &  x632 &  x641 &  x644 &  x650 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x680 &  x689 &  x698 &  x701 &  x707 &  x710 &  x728 &  x734 &  x740 &  x755 &  x770 &  x785 &  x794 &  x809 &  x818 &  x820 &  x830 &  x842 &  x854 &  x866 &  x869 &  x878 &  x899 &  x901 &  x905 &  x917 &  x926 &  x929 &  x938 &  x940 &  x941 &  x947 &  x953 &  x965 &  x968 &  x971 &  x974 &  x979 &  x980 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1015 &  x1016 &  x1025 &  x1040 &  x1046 &  x1049 &  x1052 &  x1057 &  x1064 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1096 &  x1097 &  x1100 &  x1103 &  x1109 &  x1121 &  x1127 & ~x1050 & ~x1129;
assign c0198 =  x5 &  x14 &  x17 &  x23 &  x26 &  x35 &  x41 &  x47 &  x50 &  x62 &  x65 &  x74 &  x83 &  x92 &  x101 &  x113 &  x116 &  x119 &  x131 &  x137 &  x146 &  x149 &  x155 &  x161 &  x164 &  x176 &  x179 &  x185 &  x209 &  x212 &  x215 &  x218 &  x224 &  x230 &  x236 &  x245 &  x260 &  x263 &  x275 &  x287 &  x299 &  x302 &  x308 &  x311 &  x316 &  x317 &  x332 &  x347 &  x352 &  x359 &  x374 &  x377 &  x380 &  x386 &  x389 &  x391 &  x398 &  x404 &  x407 &  x416 &  x422 &  x425 &  x430 &  x431 &  x433 &  x434 &  x443 &  x446 &  x455 &  x476 &  x494 &  x500 &  x511 &  x515 &  x518 &  x530 &  x533 &  x536 &  x538 &  x545 &  x550 &  x557 &  x563 &  x572 &  x578 &  x584 &  x587 &  x596 &  x599 &  x605 &  x617 &  x626 &  x628 &  x632 &  x644 &  x659 &  x662 &  x665 &  x667 &  x671 &  x674 &  x677 &  x680 &  x689 &  x707 &  x710 &  x713 &  x719 &  x722 &  x728 &  x734 &  x746 &  x752 &  x755 &  x761 &  x764 &  x766 &  x767 &  x773 &  x776 &  x779 &  x782 &  x788 &  x794 &  x803 &  x809 &  x815 &  x829 &  x830 &  x833 &  x836 &  x839 &  x845 &  x851 &  x854 &  x857 &  x866 &  x869 &  x872 &  x884 &  x890 &  x899 &  x902 &  x908 &  x920 &  x923 &  x929 &  x932 &  x935 &  x950 &  x953 &  x956 &  x959 &  x962 &  x968 &  x971 &  x974 &  x983 &  x989 &  x992 &  x998 &  x1007 &  x1013 &  x1031 &  x1034 &  x1046 &  x1049 &  x1058 &  x1064 &  x1067 &  x1079 &  x1085 &  x1088 &  x1091 &  x1100 &  x1103 &  x1118 &  x1121 &  x1124 & ~x72;
assign c0200 =  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x92 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x251 &  x260 &  x263 &  x269 &  x272 &  x275 &  x278 &  x284 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x317 &  x320 &  x326 &  x329 &  x332 &  x335 &  x341 &  x344 &  x347 &  x350 &  x353 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x400 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x434 &  x437 &  x439 &  x440 &  x443 &  x446 &  x452 &  x455 &  x458 &  x461 &  x467 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x506 &  x508 &  x509 &  x512 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x542 &  x545 &  x547 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x580 &  x581 &  x584 &  x586 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x626 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x785 &  x791 &  x797 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x851 &  x854 &  x857 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x890 &  x893 &  x896 &  x899 &  x901 &  x902 &  x914 &  x917 &  x920 &  x926 &  x929 &  x932 &  x935 &  x938 &  x940 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x976 &  x977 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x237 & ~x276 & ~x354 & ~x435 & ~x492;
assign c0202 =  x5 &  x14 &  x17 &  x32 &  x38 &  x41 &  x44 &  x56 &  x62 &  x65 &  x74 &  x83 &  x86 &  x89 &  x92 &  x98 &  x101 &  x104 &  x107 &  x113 &  x116 &  x119 &  x134 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x161 &  x164 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x230 &  x236 &  x242 &  x245 &  x251 &  x254 &  x257 &  x263 &  x266 &  x272 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x317 &  x320 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x359 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x395 &  x401 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x443 &  x446 &  x452 &  x455 &  x458 &  x461 &  x464 &  x470 &  x473 &  x476 &  x479 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x506 &  x509 &  x512 &  x515 &  x518 &  x536 &  x542 &  x545 &  x548 &  x551 &  x557 &  x563 &  x566 &  x572 &  x575 &  x578 &  x581 &  x584 &  x590 &  x593 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x664 &  x671 &  x674 &  x677 &  x683 &  x692 &  x701 &  x704 &  x707 &  x710 &  x713 &  x719 &  x722 &  x728 &  x734 &  x740 &  x742 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x779 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x827 &  x830 &  x836 &  x839 &  x842 &  x851 &  x854 &  x857 &  x859 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x893 &  x896 &  x898 &  x911 &  x917 &  x920 &  x923 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x989 &  x992 &  x995 &  x1004 &  x1010 &  x1016 &  x1018 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x120 & ~x159 & ~x198 & ~x201 & ~x237 & ~x315 & ~x318 & ~x432 & ~x471 & ~x648 & ~x669 & ~x747 & ~x867;
assign c0204 =  x2 &  x5 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x53 &  x56 &  x59 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x107 &  x110 &  x113 &  x119 &  x122 &  x125 &  x134 &  x137 &  x146 &  x152 &  x155 &  x158 &  x164 &  x167 &  x173 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x272 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x317 &  x320 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x368 &  x371 &  x374 &  x380 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x410 &  x413 &  x425 &  x428 &  x431 &  x437 &  x440 &  x443 &  x446 &  x452 &  x455 &  x458 &  x464 &  x467 &  x470 &  x473 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x506 &  x512 &  x515 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x547 &  x548 &  x551 &  x554 &  x557 &  x560 &  x566 &  x569 &  x572 &  x575 &  x578 &  x584 &  x587 &  x590 &  x599 &  x602 &  x605 &  x608 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x662 &  x664 &  x665 &  x668 &  x674 &  x680 &  x686 &  x689 &  x692 &  x695 &  x701 &  x703 &  x704 &  x710 &  x713 &  x716 &  x719 &  x722 &  x728 &  x731 &  x742 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x764 &  x767 &  x770 &  x773 &  x781 &  x782 &  x785 &  x788 &  x791 &  x794 &  x803 &  x806 &  x809 &  x818 &  x821 &  x824 &  x827 &  x842 &  x845 &  x848 &  x851 &  x854 &  x859 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x890 &  x893 &  x896 &  x898 &  x899 &  x901 &  x902 &  x905 &  x911 &  x914 &  x920 &  x923 &  x926 &  x929 &  x932 &  x937 &  x938 &  x940 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x968 &  x971 &  x974 &  x976 &  x977 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1049 &  x1052 &  x1058 &  x1064 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x393 & ~x525 & ~x591 & ~x603 & ~x630 & ~x648 & ~x669 & ~x687 & ~x726 & ~x747;
assign c0206 =  x2 &  x8 &  x14 &  x17 &  x23 &  x26 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x56 &  x62 &  x65 &  x68 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x152 &  x155 &  x158 &  x167 &  x170 &  x173 &  x176 &  x179 &  x185 &  x191 &  x194 &  x200 &  x203 &  x206 &  x209 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x248 &  x251 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x314 &  x317 &  x326 &  x329 &  x338 &  x341 &  x344 &  x347 &  x350 &  x356 &  x359 &  x365 &  x368 &  x371 &  x380 &  x383 &  x389 &  x392 &  x395 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x488 &  x491 &  x494 &  x497 &  x503 &  x506 &  x509 &  x512 &  x515 &  x521 &  x530 &  x533 &  x536 &  x542 &  x548 &  x551 &  x554 &  x557 &  x560 &  x566 &  x569 &  x575 &  x578 &  x581 &  x584 &  x586 &  x590 &  x593 &  x596 &  x599 &  x602 &  x608 &  x614 &  x620 &  x623 &  x625 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x698 &  x707 &  x710 &  x713 &  x719 &  x722 &  x725 &  x731 &  x734 &  x740 &  x743 &  x745 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x770 &  x776 &  x779 &  x782 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x818 &  x821 &  x822 &  x823 &  x824 &  x827 &  x830 &  x836 &  x842 &  x848 &  x854 &  x857 &  x860 &  x861 &  x862 &  x866 &  x878 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x900 &  x902 &  x905 &  x911 &  x914 &  x917 &  x920 &  x926 &  x935 &  x938 &  x940 &  x944 &  x947 &  x950 &  x956 &  x962 &  x965 &  x974 &  x977 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1013 &  x1016 &  x1018 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1033 &  x1034 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1067 &  x1070 &  x1072 &  x1073 &  x1082 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1111 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 & ~x489 & ~x756 & ~x795 & ~x834;
assign c0208 =  x2 &  x5 &  x8 &  x20 &  x23 &  x32 &  x35 &  x38 &  x41 &  x47 &  x50 &  x53 &  x59 &  x62 &  x68 &  x71 &  x101 &  x104 &  x110 &  x113 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x146 &  x149 &  x152 &  x167 &  x170 &  x176 &  x182 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x260 &  x263 &  x266 &  x272 &  x281 &  x284 &  x287 &  x293 &  x296 &  x302 &  x305 &  x308 &  x320 &  x323 &  x326 &  x329 &  x335 &  x341 &  x350 &  x374 &  x377 &  x380 &  x383 &  x391 &  x398 &  x410 &  x413 &  x419 &  x422 &  x425 &  x428 &  x431 &  x433 &  x434 &  x437 &  x443 &  x446 &  x455 &  x458 &  x461 &  x467 &  x470 &  x472 &  x473 &  x476 &  x479 &  x482 &  x491 &  x494 &  x497 &  x503 &  x509 &  x515 &  x521 &  x524 &  x530 &  x533 &  x539 &  x545 &  x548 &  x551 &  x557 &  x560 &  x563 &  x572 &  x584 &  x587 &  x590 &  x596 &  x599 &  x605 &  x608 &  x611 &  x614 &  x623 &  x626 &  x628 &  x629 &  x638 &  x641 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x671 &  x674 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x701 &  x706 &  x707 &  x719 &  x722 &  x725 &  x737 &  x743 &  x755 &  x758 &  x761 &  x764 &  x770 &  x773 &  x776 &  x779 &  x782 &  x784 &  x785 &  x787 &  x788 &  x791 &  x794 &  x800 &  x806 &  x815 &  x818 &  x823 &  x824 &  x827 &  x833 &  x836 &  x839 &  x842 &  x845 &  x854 &  x865 &  x866 &  x869 &  x878 &  x881 &  x884 &  x890 &  x896 &  x899 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x935 &  x938 &  x944 &  x956 &  x959 &  x962 &  x965 &  x980 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1010 &  x1016 &  x1019 &  x1022 &  x1031 &  x1034 &  x1043 &  x1052 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1082 &  x1085 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1121 & ~x330 & ~x375 & ~x474 & ~x516 & ~x555;
assign c0210 =  x2 &  x5 &  x11 &  x32 &  x38 &  x59 &  x65 &  x68 &  x74 &  x77 &  x83 &  x86 &  x89 &  x95 &  x98 &  x104 &  x110 &  x113 &  x116 &  x122 &  x125 &  x128 &  x131 &  x143 &  x146 &  x152 &  x161 &  x167 &  x170 &  x179 &  x185 &  x194 &  x200 &  x203 &  x206 &  x215 &  x218 &  x227 &  x236 &  x239 &  x242 &  x248 &  x257 &  x260 &  x263 &  x269 &  x272 &  x275 &  x278 &  x284 &  x287 &  x293 &  x299 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x335 &  x338 &  x341 &  x347 &  x350 &  x356 &  x362 &  x380 &  x383 &  x389 &  x391 &  x395 &  x407 &  x413 &  x419 &  x425 &  x431 &  x434 &  x437 &  x440 &  x446 &  x449 &  x452 &  x455 &  x461 &  x464 &  x470 &  x472 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x509 &  x511 &  x512 &  x521 &  x527 &  x530 &  x533 &  x539 &  x542 &  x548 &  x554 &  x557 &  x560 &  x563 &  x569 &  x572 &  x577 &  x578 &  x581 &  x590 &  x593 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x616 &  x617 &  x623 &  x626 &  x632 &  x638 &  x641 &  x644 &  x647 &  x653 &  x656 &  x662 &  x665 &  x671 &  x677 &  x692 &  x695 &  x698 &  x701 &  x704 &  x713 &  x719 &  x725 &  x731 &  x734 &  x743 &  x746 &  x749 &  x755 &  x761 &  x770 &  x776 &  x779 &  x791 &  x799 &  x803 &  x818 &  x824 &  x827 &  x836 &  x848 &  x854 &  x866 &  x869 &  x872 &  x878 &  x887 &  x896 &  x899 &  x905 &  x908 &  x914 &  x917 &  x920 &  x926 &  x932 &  x938 &  x941 &  x947 &  x950 &  x959 &  x968 &  x971 &  x983 &  x986 &  x989 &  x1001 &  x1019 &  x1022 &  x1025 &  x1031 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1070 &  x1082 &  x1085 &  x1088 &  x1094 &  x1103 &  x1109 &  x1112 &  x1121 &  x1124 &  x1130 & ~x138 & ~x663 & ~x768 & ~x912 & ~x1047;
assign c0212 =  x2 &  x11 &  x14 &  x17 &  x23 &  x29 &  x35 &  x44 &  x47 &  x50 &  x53 &  x65 &  x68 &  x71 &  x74 &  x77 &  x83 &  x89 &  x92 &  x95 &  x98 &  x104 &  x107 &  x110 &  x113 &  x122 &  x125 &  x128 &  x131 &  x137 &  x149 &  x152 &  x164 &  x170 &  x173 &  x176 &  x182 &  x185 &  x188 &  x194 &  x197 &  x203 &  x206 &  x209 &  x212 &  x224 &  x227 &  x233 &  x236 &  x245 &  x248 &  x254 &  x263 &  x266 &  x272 &  x275 &  x278 &  x281 &  x290 &  x298 &  x299 &  x302 &  x317 &  x323 &  x332 &  x338 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x368 &  x370 &  x371 &  x374 &  x377 &  x380 &  x389 &  x392 &  x395 &  x398 &  x407 &  x413 &  x422 &  x425 &  x431 &  x437 &  x443 &  x449 &  x455 &  x458 &  x461 &  x467 &  x470 &  x473 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x509 &  x515 &  x518 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x545 &  x551 &  x554 &  x560 &  x563 &  x569 &  x572 &  x575 &  x581 &  x593 &  x596 &  x599 &  x605 &  x608 &  x617 &  x620 &  x623 &  x626 &  x629 &  x638 &  x641 &  x647 &  x653 &  x659 &  x662 &  x664 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x703 &  x704 &  x707 &  x713 &  x716 &  x719 &  x722 &  x725 &  x731 &  x734 &  x737 &  x740 &  x742 &  x743 &  x752 &  x755 &  x761 &  x767 &  x773 &  x781 &  x788 &  x791 &  x794 &  x803 &  x809 &  x812 &  x818 &  x820 &  x824 &  x833 &  x836 &  x851 &  x857 &  x859 &  x860 &  x862 &  x863 &  x872 &  x875 &  x881 &  x887 &  x893 &  x896 &  x898 &  x899 &  x901 &  x902 &  x905 &  x917 &  x923 &  x926 &  x929 &  x941 &  x944 &  x950 &  x959 &  x962 &  x965 &  x968 &  x971 &  x977 &  x979 &  x986 &  x989 &  x992 &  x998 &  x1004 &  x1007 &  x1010 &  x1013 &  x1015 &  x1017 &  x1018 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1052 &  x1055 &  x1056 &  x1057 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1096 &  x1103 &  x1106 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x273 & ~x312 & ~x351 & ~x669 & ~x723 & ~x747 & ~x762 & ~x786;
assign c0214 =  x2 &  x5 &  x11 &  x17 &  x20 &  x23 &  x29 &  x32 &  x35 &  x41 &  x47 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x98 &  x101 &  x104 &  x110 &  x119 &  x125 &  x128 &  x131 &  x134 &  x140 &  x146 &  x149 &  x152 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x191 &  x194 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x239 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x272 &  x278 &  x281 &  x284 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x317 &  x320 &  x326 &  x329 &  x332 &  x335 &  x341 &  x344 &  x353 &  x356 &  x359 &  x362 &  x365 &  x371 &  x377 &  x383 &  x386 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x416 &  x428 &  x431 &  x434 &  x449 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x482 &  x485 &  x488 &  x491 &  x494 &  x503 &  x506 &  x512 &  x515 &  x518 &  x527 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x550 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x584 &  x587 &  x589 &  x590 &  x596 &  x599 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x628 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x656 &  x659 &  x662 &  x668 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x701 &  x707 &  x710 &  x713 &  x716 &  x719 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x749 &  x752 &  x755 &  x761 &  x764 &  x767 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x845 &  x848 &  x851 &  x854 &  x857 &  x863 &  x866 &  x869 &  x875 &  x878 &  x881 &  x887 &  x890 &  x893 &  x899 &  x902 &  x905 &  x911 &  x916 &  x917 &  x920 &  x926 &  x929 &  x932 &  x938 &  x941 &  x953 &  x954 &  x955 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x986 &  x989 &  x993 &  x994 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1033 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1072 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x6 & ~x138 & ~x177 & ~x1092;
assign c0216 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x26 &  x32 &  x35 &  x38 &  x41 &  x44 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x86 &  x89 &  x95 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x314 &  x317 &  x320 &  x323 &  x329 &  x332 &  x335 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x389 &  x392 &  x394 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x473 &  x476 &  x479 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x589 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x626 &  x628 &  x629 &  x632 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x662 &  x665 &  x668 &  x671 &  x674 &  x680 &  x686 &  x689 &  x695 &  x698 &  x701 &  x707 &  x710 &  x722 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x745 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x773 &  x779 &  x784 &  x788 &  x791 &  x797 &  x803 &  x806 &  x809 &  x811 &  x812 &  x815 &  x818 &  x821 &  x824 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x857 &  x860 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x949 &  x950 &  x953 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x988 &  x989 &  x992 &  x998 &  x1001 &  x1004 &  x1010 &  x1016 &  x1022 &  x1025 &  x1027 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1058 &  x1061 &  x1064 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x27 & ~x93 & ~x555;
assign c0218 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x23 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x101 &  x104 &  x107 &  x110 &  x113 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x170 &  x173 &  x176 &  x179 &  x182 &  x194 &  x197 &  x209 &  x215 &  x221 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x251 &  x254 &  x257 &  x260 &  x266 &  x269 &  x272 &  x274 &  x275 &  x281 &  x284 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x312 &  x314 &  x317 &  x320 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x351 &  x352 &  x353 &  x359 &  x365 &  x368 &  x371 &  x374 &  x380 &  x383 &  x386 &  x391 &  x394 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x430 &  x433 &  x440 &  x443 &  x446 &  x452 &  x455 &  x458 &  x461 &  x469 &  x470 &  x473 &  x476 &  x482 &  x488 &  x491 &  x494 &  x497 &  x500 &  x506 &  x508 &  x509 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x545 &  x547 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x575 &  x578 &  x584 &  x587 &  x593 &  x596 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x625 &  x628 &  x629 &  x632 &  x638 &  x641 &  x644 &  x650 &  x653 &  x656 &  x659 &  x667 &  x668 &  x671 &  x674 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x745 &  x749 &  x752 &  x755 &  x758 &  x764 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x872 &  x875 &  x878 &  x884 &  x887 &  x890 &  x893 &  x902 &  x905 &  x911 &  x914 &  x917 &  x926 &  x929 &  x932 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x977 &  x980 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1036 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1064 &  x1067 &  x1070 &  x1073 &  x1075 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 &  x1130 & ~x396 & ~x435;
assign c0220 =  x11 &  x20 &  x29 &  x38 &  x50 &  x56 &  x65 &  x71 &  x74 &  x77 &  x80 &  x89 &  x92 &  x98 &  x101 &  x107 &  x116 &  x119 &  x131 &  x146 &  x152 &  x170 &  x182 &  x185 &  x191 &  x194 &  x206 &  x209 &  x215 &  x218 &  x221 &  x224 &  x233 &  x236 &  x245 &  x247 &  x248 &  x251 &  x257 &  x260 &  x269 &  x272 &  x275 &  x287 &  x290 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x320 &  x323 &  x329 &  x332 &  x335 &  x347 &  x356 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x404 &  x407 &  x410 &  x419 &  x425 &  x428 &  x434 &  x437 &  x440 &  x458 &  x464 &  x482 &  x485 &  x494 &  x500 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x545 &  x548 &  x551 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x590 &  x599 &  x608 &  x614 &  x620 &  x623 &  x625 &  x626 &  x632 &  x638 &  x641 &  x650 &  x659 &  x664 &  x665 &  x668 &  x671 &  x680 &  x683 &  x692 &  x695 &  x701 &  x703 &  x704 &  x710 &  x713 &  x725 &  x731 &  x734 &  x737 &  x745 &  x755 &  x761 &  x764 &  x770 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x815 &  x820 &  x821 &  x823 &  x824 &  x830 &  x839 &  x842 &  x851 &  x862 &  x863 &  x869 &  x872 &  x884 &  x890 &  x893 &  x898 &  x900 &  x908 &  x917 &  x923 &  x929 &  x932 &  x938 &  x941 &  x944 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x976 &  x978 &  x989 &  x1001 &  x1004 &  x1010 &  x1013 &  x1015 &  x1017 &  x1018 &  x1019 &  x1025 &  x1031 &  x1034 &  x1043 &  x1052 &  x1055 &  x1057 &  x1058 &  x1064 &  x1070 &  x1082 &  x1100 &  x1105 &  x1109 &  x1118 &  x1121 &  x1127 &  x1130 & ~x117 & ~x156 & ~x195 & ~x354 & ~x648;
assign c0222 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x289 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x625 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x703 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x733 &  x734 &  x737 &  x740 &  x742 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x772 &  x773 &  x776 &  x779 &  x781 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x810 &  x811 &  x812 &  x815 &  x818 &  x820 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x850 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x889 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1018 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1096 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130;
assign c0224 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x442 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x625 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x668 &  x671 &  x674 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x703 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x742 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x781 &  x782 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x820 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x859 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x898 &  x899 &  x901 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x940 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1072 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1111 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x354 & ~x393 & ~x432 & ~x591 & ~x630 & ~x669;
assign c0226 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x247 &  x248 &  x254 &  x257 &  x260 &  x263 &  x265 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x296 &  x299 &  x302 &  x304 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x443 &  x446 &  x449 &  x455 &  x458 &  x461 &  x464 &  x470 &  x473 &  x476 &  x479 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x625 &  x626 &  x629 &  x632 &  x638 &  x641 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x698 &  x701 &  x703 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x769 &  x770 &  x773 &  x776 &  x785 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x808 &  x809 &  x812 &  x815 &  x818 &  x821 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x950 &  x953 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1130 & ~x237 & ~x276 & ~x315 & ~x354 & ~x393 & ~x606 & ~x795;
assign c0228 =  x5 &  x14 &  x23 &  x26 &  x32 &  x35 &  x38 &  x56 &  x59 &  x65 &  x68 &  x80 &  x83 &  x89 &  x98 &  x104 &  x110 &  x122 &  x128 &  x137 &  x140 &  x143 &  x146 &  x149 &  x155 &  x164 &  x173 &  x176 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x206 &  x212 &  x221 &  x230 &  x236 &  x245 &  x260 &  x263 &  x269 &  x275 &  x293 &  x305 &  x314 &  x317 &  x323 &  x326 &  x338 &  x344 &  x350 &  x362 &  x365 &  x377 &  x389 &  x392 &  x394 &  x398 &  x404 &  x407 &  x410 &  x419 &  x422 &  x425 &  x437 &  x440 &  x443 &  x449 &  x452 &  x470 &  x476 &  x479 &  x482 &  x491 &  x494 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x527 &  x533 &  x554 &  x560 &  x569 &  x572 &  x578 &  x581 &  x584 &  x587 &  x590 &  x602 &  x605 &  x608 &  x614 &  x617 &  x641 &  x647 &  x650 &  x653 &  x674 &  x677 &  x683 &  x686 &  x695 &  x701 &  x704 &  x710 &  x713 &  x716 &  x722 &  x725 &  x727 &  x734 &  x755 &  x758 &  x761 &  x776 &  x785 &  x788 &  x800 &  x812 &  x815 &  x827 &  x830 &  x832 &  x839 &  x845 &  x851 &  x857 &  x863 &  x869 &  x875 &  x878 &  x884 &  x890 &  x893 &  x902 &  x917 &  x923 &  x935 &  x938 &  x941 &  x950 &  x956 &  x962 &  x965 &  x974 &  x980 &  x986 &  x992 &  x1004 &  x1007 &  x1016 &  x1019 &  x1022 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1064 &  x1076 &  x1079 &  x1082 &  x1088 &  x1094 &  x1100 &  x1103 &  x1106 &  x1115 &  x1121 &  x1124 &  x1130 & ~x516 & ~x555 & ~x582 & ~x852 & ~x885 & ~x924;
assign c0230 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x284 &  x287 &  x290 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x667 &  x668 &  x671 &  x674 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x698 &  x700 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x739 &  x740 &  x743 &  x745 &  x746 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x949 &  x950 &  x953 &  x956 &  x959 &  x962 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x988 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1027 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x198 & ~x237 & ~x276 & ~x315 & ~x354 & ~x393 & ~x570;
assign c0232 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x312 &  x313 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x351 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x390 &  x391 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x430 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x469 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x508 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x547 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x785 &  x788 &  x791 &  x794 &  x797 &  x803 &  x806 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x240 & ~x279 & ~x318 & ~x357 & ~x396 & ~x397 & ~x435 & ~x436 & ~x474 & ~x513 & ~x591 & ~x630 & ~x942 & ~x1020 & ~x1059;
assign c0234 =  x2 &  x5 &  x17 &  x29 &  x32 &  x38 &  x41 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x95 &  x98 &  x104 &  x113 &  x122 &  x128 &  x134 &  x140 &  x146 &  x152 &  x155 &  x161 &  x164 &  x173 &  x176 &  x179 &  x193 &  x197 &  x200 &  x203 &  x206 &  x218 &  x224 &  x227 &  x230 &  x233 &  x245 &  x251 &  x257 &  x263 &  x269 &  x272 &  x275 &  x284 &  x293 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x338 &  x341 &  x344 &  x350 &  x356 &  x362 &  x374 &  x377 &  x380 &  x383 &  x395 &  x398 &  x401 &  x413 &  x422 &  x425 &  x427 &  x428 &  x431 &  x437 &  x440 &  x443 &  x452 &  x458 &  x461 &  x464 &  x473 &  x482 &  x485 &  x488 &  x491 &  x497 &  x509 &  x515 &  x518 &  x521 &  x524 &  x530 &  x533 &  x542 &  x548 &  x551 &  x554 &  x560 &  x563 &  x572 &  x575 &  x581 &  x596 &  x599 &  x611 &  x614 &  x620 &  x626 &  x635 &  x641 &  x650 &  x653 &  x656 &  x662 &  x671 &  x677 &  x680 &  x683 &  x686 &  x692 &  x701 &  x707 &  x710 &  x713 &  x716 &  x719 &  x725 &  x731 &  x734 &  x737 &  x740 &  x758 &  x761 &  x782 &  x791 &  x794 &  x806 &  x809 &  x812 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x848 &  x854 &  x856 &  x866 &  x872 &  x878 &  x881 &  x884 &  x896 &  x899 &  x905 &  x908 &  x911 &  x914 &  x919 &  x920 &  x926 &  x929 &  x938 &  x941 &  x944 &  x947 &  x959 &  x968 &  x980 &  x983 &  x992 &  x1004 &  x1010 &  x1016 &  x1025 &  x1031 &  x1037 &  x1040 &  x1052 &  x1067 &  x1070 &  x1075 &  x1079 &  x1082 &  x1091 &  x1094 &  x1097 &  x1100 &  x1102 &  x1103 &  x1109 &  x1115 &  x1121 & ~x1041;
assign c0236 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x56 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x86 &  x92 &  x95 &  x98 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x156 &  x157 &  x158 &  x167 &  x170 &  x176 &  x179 &  x182 &  x188 &  x195 &  x196 &  x197 &  x206 &  x209 &  x212 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x234 &  x235 &  x236 &  x238 &  x239 &  x242 &  x257 &  x260 &  x263 &  x269 &  x272 &  x273 &  x274 &  x275 &  x284 &  x290 &  x293 &  x296 &  x299 &  x316 &  x320 &  x323 &  x329 &  x338 &  x344 &  x347 &  x352 &  x353 &  x355 &  x356 &  x365 &  x371 &  x374 &  x377 &  x391 &  x392 &  x394 &  x398 &  x401 &  x404 &  x410 &  x416 &  x422 &  x428 &  x431 &  x433 &  x434 &  x446 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x473 &  x476 &  x482 &  x485 &  x494 &  x497 &  x500 &  x509 &  x511 &  x515 &  x518 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x550 &  x551 &  x575 &  x587 &  x593 &  x596 &  x605 &  x608 &  x611 &  x620 &  x626 &  x628 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x674 &  x686 &  x689 &  x695 &  x701 &  x713 &  x716 &  x719 &  x722 &  x731 &  x734 &  x737 &  x746 &  x749 &  x752 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x794 &  x800 &  x803 &  x806 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x842 &  x851 &  x857 &  x860 &  x869 &  x875 &  x878 &  x881 &  x884 &  x890 &  x899 &  x902 &  x908 &  x911 &  x914 &  x917 &  x920 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x959 &  x962 &  x965 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x992 &  x998 &  x1007 &  x1010 &  x1013 &  x1022 &  x1025 &  x1028 &  x1034 &  x1037 &  x1040 &  x1049 &  x1055 &  x1058 &  x1064 &  x1070 &  x1082 &  x1088 &  x1097 &  x1103 &  x1112 &  x1115 &  x1118 &  x1124 &  x1130 & ~x162 & ~x240 & ~x402 & ~x741;
assign c0238 =  x2 &  x5 &  x11 &  x17 &  x20 &  x23 &  x26 &  x32 &  x35 &  x41 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x86 &  x89 &  x92 &  x98 &  x101 &  x104 &  x110 &  x116 &  x122 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x158 &  x161 &  x167 &  x176 &  x179 &  x182 &  x185 &  x194 &  x197 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x257 &  x260 &  x263 &  x272 &  x275 &  x278 &  x281 &  x284 &  x290 &  x299 &  x305 &  x311 &  x314 &  x316 &  x317 &  x320 &  x326 &  x329 &  x332 &  x335 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x355 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x383 &  x389 &  x391 &  x394 &  x395 &  x404 &  x416 &  x419 &  x425 &  x428 &  x431 &  x433 &  x434 &  x440 &  x443 &  x449 &  x461 &  x464 &  x467 &  x472 &  x476 &  x479 &  x482 &  x485 &  x488 &  x494 &  x500 &  x506 &  x511 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x542 &  x545 &  x550 &  x551 &  x554 &  x557 &  x560 &  x566 &  x569 &  x572 &  x575 &  x578 &  x584 &  x587 &  x599 &  x602 &  x605 &  x614 &  x616 &  x617 &  x620 &  x632 &  x635 &  x641 &  x656 &  x668 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x701 &  x704 &  x707 &  x719 &  x722 &  x731 &  x737 &  x740 &  x749 &  x752 &  x758 &  x764 &  x767 &  x770 &  x776 &  x779 &  x785 &  x791 &  x794 &  x797 &  x803 &  x806 &  x811 &  x812 &  x815 &  x821 &  x824 &  x827 &  x830 &  x832 &  x833 &  x836 &  x839 &  x842 &  x845 &  x850 &  x851 &  x854 &  x857 &  x860 &  x866 &  x878 &  x881 &  x883 &  x884 &  x887 &  x890 &  x896 &  x902 &  x905 &  x908 &  x910 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x938 &  x941 &  x944 &  x953 &  x956 &  x965 &  x967 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x994 &  x1004 &  x1006 &  x1016 &  x1019 &  x1022 &  x1028 &  x1031 &  x1033 &  x1034 &  x1037 &  x1040 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 & ~x216 & ~x336 & ~x741 & ~x780 & ~x819;
assign c0240 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x289 &  x290 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x523 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x625 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x703 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x742 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x781 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x820 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x859 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x896 &  x898 &  x899 &  x901 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x937 &  x938 &  x940 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1015 &  x1016 &  x1018 &  x1019 &  x1022 &  x1025 &  x1028 &  x1030 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1054 &  x1055 &  x1057 &  x1058 &  x1061 &  x1064 &  x1067 &  x1068 &  x1069 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1096 &  x1097 &  x1100 &  x1103 &  x1106 &  x1108 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 &  x1130 & ~x753 & ~x792;
assign c0242 =  x5 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x35 &  x38 &  x41 &  x50 &  x53 &  x56 &  x62 &  x65 &  x74 &  x77 &  x83 &  x89 &  x92 &  x98 &  x110 &  x113 &  x116 &  x119 &  x137 &  x140 &  x146 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x230 &  x233 &  x245 &  x248 &  x260 &  x263 &  x266 &  x272 &  x275 &  x278 &  x284 &  x290 &  x293 &  x296 &  x299 &  x302 &  x311 &  x314 &  x320 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x356 &  x359 &  x365 &  x368 &  x374 &  x380 &  x389 &  x395 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x431 &  x434 &  x437 &  x443 &  x449 &  x452 &  x455 &  x461 &  x464 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x551 &  x557 &  x569 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x613 &  x614 &  x620 &  x623 &  x626 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x652 &  x656 &  x662 &  x665 &  x668 &  x671 &  x674 &  x680 &  x683 &  x686 &  x689 &  x690 &  x692 &  x695 &  x701 &  x707 &  x710 &  x712 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x730 &  x731 &  x734 &  x740 &  x743 &  x746 &  x749 &  x761 &  x764 &  x767 &  x769 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x827 &  x830 &  x833 &  x836 &  x839 &  x845 &  x847 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x875 &  x877 &  x881 &  x884 &  x886 &  x887 &  x890 &  x896 &  x902 &  x905 &  x911 &  x914 &  x916 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x941 &  x944 &  x947 &  x950 &  x953 &  x955 &  x965 &  x971 &  x974 &  x977 &  x985 &  x989 &  x991 &  x992 &  x995 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1021 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1060 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130;
assign c0244 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x29 &  x32 &  x35 &  x38 &  x44 &  x47 &  x50 &  x53 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x469 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x812 &  x815 &  x818 &  x821 &  x827 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x435 & ~x474 & ~x489 & ~x513 & ~x528 & ~x555 & ~x567 & ~x594 & ~x633 & ~x672 & ~x756 & ~x774 & ~x795 & ~x813 & ~x852;
assign c0246 =  x5 &  x8 &  x11 &  x14 &  x17 &  x23 &  x26 &  x29 &  x32 &  x35 &  x41 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x77 &  x80 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x113 &  x116 &  x119 &  x125 &  x128 &  x137 &  x143 &  x146 &  x149 &  x152 &  x155 &  x164 &  x167 &  x170 &  x173 &  x176 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x218 &  x221 &  x227 &  x230 &  x233 &  x248 &  x251 &  x257 &  x266 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x317 &  x320 &  x326 &  x332 &  x338 &  x344 &  x347 &  x350 &  x353 &  x356 &  x365 &  x368 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x395 &  x398 &  x404 &  x407 &  x410 &  x413 &  x419 &  x422 &  x428 &  x431 &  x437 &  x440 &  x446 &  x449 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x485 &  x488 &  x491 &  x494 &  x503 &  x506 &  x524 &  x530 &  x533 &  x536 &  x539 &  x548 &  x551 &  x554 &  x560 &  x563 &  x569 &  x578 &  x581 &  x584 &  x590 &  x593 &  x596 &  x599 &  x602 &  x611 &  x614 &  x617 &  x626 &  x629 &  x632 &  x635 &  x641 &  x644 &  x647 &  x650 &  x656 &  x659 &  x662 &  x674 &  x677 &  x686 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x749 &  x758 &  x761 &  x764 &  x770 &  x773 &  x779 &  x782 &  x785 &  x788 &  x791 &  x800 &  x803 &  x806 &  x809 &  x815 &  x821 &  x824 &  x827 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x872 &  x875 &  x878 &  x890 &  x893 &  x896 &  x899 &  x905 &  x908 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x950 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1058 &  x1061 &  x1067 &  x1079 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1127 &  x1130 & ~x6 & ~x51 & ~x66 & ~x84 & ~x90 & ~x123 & ~x126 & ~x129 & ~x168 & ~x216 & ~x255 & ~x294 & ~x852 & ~x963 & ~x969 & ~x1008 & ~x1041 & ~x1047;
assign c0248 =  x2 &  x5 &  x8 &  x11 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x107 &  x110 &  x116 &  x119 &  x122 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x155 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x206 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x390 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x429 &  x430 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x455 &  x458 &  x461 &  x464 &  x467 &  x469 &  x470 &  x476 &  x479 &  x482 &  x485 &  x488 &  x497 &  x500 &  x506 &  x508 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x547 &  x548 &  x551 &  x554 &  x560 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x625 &  x626 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x656 &  x659 &  x664 &  x665 &  x667 &  x668 &  x671 &  x674 &  x677 &  x680 &  x686 &  x689 &  x692 &  x701 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x731 &  x734 &  x737 &  x740 &  x743 &  x745 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x860 &  x863 &  x866 &  x869 &  x875 &  x878 &  x881 &  x884 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x913 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x947 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1070 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x396 & ~x435 & ~x474 & ~x513 & ~x555;
assign c0250 =  x8 &  x11 &  x14 &  x20 &  x23 &  x38 &  x47 &  x53 &  x59 &  x65 &  x68 &  x71 &  x80 &  x92 &  x95 &  x101 &  x110 &  x113 &  x131 &  x143 &  x158 &  x161 &  x164 &  x170 &  x176 &  x182 &  x185 &  x188 &  x194 &  x197 &  x200 &  x206 &  x209 &  x215 &  x218 &  x227 &  x242 &  x245 &  x248 &  x254 &  x280 &  x284 &  x286 &  x293 &  x296 &  x302 &  x305 &  x314 &  x320 &  x325 &  x326 &  x329 &  x332 &  x341 &  x344 &  x356 &  x368 &  x386 &  x392 &  x404 &  x407 &  x413 &  x422 &  x434 &  x437 &  x440 &  x458 &  x467 &  x470 &  x473 &  x476 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x506 &  x515 &  x527 &  x530 &  x533 &  x536 &  x542 &  x548 &  x560 &  x563 &  x569 &  x575 &  x587 &  x590 &  x593 &  x596 &  x599 &  x608 &  x614 &  x620 &  x626 &  x638 &  x647 &  x656 &  x659 &  x662 &  x665 &  x671 &  x677 &  x683 &  x689 &  x698 &  x703 &  x704 &  x707 &  x725 &  x728 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x781 &  x785 &  x788 &  x794 &  x803 &  x806 &  x812 &  x815 &  x818 &  x824 &  x830 &  x836 &  x839 &  x842 &  x845 &  x860 &  x863 &  x869 &  x872 &  x881 &  x887 &  x890 &  x893 &  x896 &  x899 &  x901 &  x902 &  x911 &  x917 &  x926 &  x935 &  x939 &  x941 &  x944 &  x959 &  x968 &  x974 &  x977 &  x979 &  x980 &  x983 &  x986 &  x995 &  x1007 &  x1013 &  x1018 &  x1022 &  x1028 &  x1046 &  x1049 &  x1058 &  x1061 &  x1067 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1109 &  x1112 &  x1115 &  x1124 &  x1127 &  x1130 & ~x306 & ~x351 & ~x528 & ~x591;
assign c0252 =  x11 &  x23 &  x26 &  x29 &  x32 &  x38 &  x50 &  x56 &  x59 &  x68 &  x74 &  x77 &  x86 &  x89 &  x95 &  x98 &  x116 &  x125 &  x128 &  x131 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x194 &  x197 &  x200 &  x203 &  x206 &  x218 &  x221 &  x227 &  x230 &  x233 &  x239 &  x263 &  x278 &  x287 &  x293 &  x296 &  x302 &  x323 &  x326 &  x329 &  x338 &  x344 &  x347 &  x350 &  x365 &  x374 &  x377 &  x380 &  x386 &  x392 &  x394 &  x395 &  x419 &  x422 &  x428 &  x433 &  x440 &  x446 &  x449 &  x452 &  x458 &  x464 &  x467 &  x472 &  x473 &  x482 &  x494 &  x497 &  x506 &  x518 &  x533 &  x539 &  x542 &  x551 &  x569 &  x572 &  x584 &  x590 &  x593 &  x599 &  x611 &  x620 &  x623 &  x626 &  x629 &  x638 &  x641 &  x650 &  x653 &  x656 &  x659 &  x662 &  x674 &  x680 &  x682 &  x686 &  x689 &  x695 &  x707 &  x710 &  x713 &  x716 &  x722 &  x728 &  x734 &  x740 &  x746 &  x758 &  x760 &  x764 &  x776 &  x779 &  x788 &  x791 &  x794 &  x799 &  x800 &  x803 &  x812 &  x815 &  x824 &  x827 &  x842 &  x845 &  x848 &  x851 &  x863 &  x869 &  x875 &  x877 &  x881 &  x884 &  x887 &  x893 &  x896 &  x917 &  x926 &  x932 &  x941 &  x944 &  x947 &  x965 &  x968 &  x971 &  x974 &  x986 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1019 &  x1025 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1067 &  x1073 &  x1076 &  x1088 &  x1091 &  x1094 &  x1109 &  x1118 &  x1121 &  x1127 &  x1130 & ~x24 & ~x30 & ~x702 & ~x780 & ~x819 & ~x945 & ~x984 & ~x1059;
assign c0254 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x26 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x244 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x272 &  x274 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x312 &  x313 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x351 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x391 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x430 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x464 &  x467 &  x469 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x508 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x547 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x279 & ~x318 & ~x319 & ~x357 & ~x358 & ~x396 & ~x435 & ~x480 & ~x519 & ~x780 & ~x819;
assign c0256 =  x5 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x197 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x470 &  x473 &  x476 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x562 &  x566 &  x569 &  x572 &  x575 &  x578 &  x584 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x702 &  x703 &  x704 &  x707 &  x710 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x737 &  x740 &  x742 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x779 &  x780 &  x781 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x819 &  x820 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x858 &  x859 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x893 &  x896 &  x897 &  x898 &  x902 &  x905 &  x908 &  x911 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x936 &  x937 &  x938 &  x940 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x976 &  x977 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1054 &  x1055 &  x1057 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x351 & ~x354 & ~x393 & ~x432 & ~x471 & ~x510 & ~x549 & ~x669 & ~x708 & ~x747 & ~x870;
assign c0258 =  x2 &  x8 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x44 &  x50 &  x53 &  x56 &  x59 &  x65 &  x74 &  x77 &  x83 &  x86 &  x89 &  x95 &  x107 &  x110 &  x113 &  x122 &  x134 &  x152 &  x155 &  x161 &  x164 &  x170 &  x173 &  x179 &  x182 &  x185 &  x191 &  x194 &  x197 &  x218 &  x221 &  x227 &  x233 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x266 &  x272 &  x275 &  x278 &  x280 &  x281 &  x287 &  x290 &  x298 &  x302 &  x311 &  x317 &  x320 &  x323 &  x326 &  x329 &  x335 &  x338 &  x341 &  x353 &  x362 &  x364 &  x365 &  x371 &  x380 &  x389 &  x395 &  x401 &  x416 &  x419 &  x422 &  x425 &  x431 &  x434 &  x437 &  x440 &  x443 &  x452 &  x455 &  x467 &  x476 &  x479 &  x491 &  x494 &  x497 &  x500 &  x503 &  x512 &  x518 &  x527 &  x530 &  x539 &  x554 &  x560 &  x563 &  x572 &  x575 &  x578 &  x584 &  x590 &  x593 &  x596 &  x601 &  x602 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x640 &  x641 &  x644 &  x650 &  x659 &  x662 &  x664 &  x665 &  x671 &  x680 &  x686 &  x689 &  x695 &  x698 &  x701 &  x704 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x731 &  x734 &  x743 &  x749 &  x752 &  x755 &  x758 &  x764 &  x767 &  x770 &  x776 &  x782 &  x785 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x820 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x859 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x893 &  x898 &  x902 &  x905 &  x908 &  x911 &  x917 &  x926 &  x929 &  x932 &  x938 &  x944 &  x947 &  x956 &  x962 &  x965 &  x968 &  x971 &  x976 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1043 &  x1049 &  x1054 &  x1055 &  x1057 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1093 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1124 &  x1130 & ~x354 & ~x393 & ~x471 & ~x708 & ~x747 & ~x786 & ~x831;
assign c0260 =  x2 &  x5 &  x8 &  x14 &  x23 &  x26 &  x32 &  x38 &  x53 &  x56 &  x59 &  x68 &  x71 &  x86 &  x92 &  x95 &  x98 &  x104 &  x107 &  x113 &  x116 &  x122 &  x128 &  x131 &  x134 &  x140 &  x146 &  x152 &  x155 &  x161 &  x164 &  x176 &  x185 &  x188 &  x191 &  x197 &  x200 &  x206 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x236 &  x239 &  x245 &  x251 &  x254 &  x266 &  x269 &  x272 &  x278 &  x281 &  x290 &  x293 &  x308 &  x311 &  x317 &  x323 &  x329 &  x332 &  x359 &  x362 &  x365 &  x371 &  x374 &  x380 &  x383 &  x386 &  x389 &  x394 &  x395 &  x398 &  x404 &  x407 &  x419 &  x422 &  x425 &  x428 &  x430 &  x440 &  x443 &  x452 &  x458 &  x461 &  x467 &  x473 &  x482 &  x485 &  x488 &  x491 &  x497 &  x500 &  x503 &  x509 &  x511 &  x512 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x542 &  x548 &  x550 &  x557 &  x560 &  x566 &  x569 &  x572 &  x575 &  x584 &  x599 &  x605 &  x608 &  x620 &  x623 &  x626 &  x632 &  x635 &  x638 &  x650 &  x653 &  x656 &  x668 &  x671 &  x674 &  x680 &  x683 &  x692 &  x695 &  x698 &  x701 &  x704 &  x710 &  x716 &  x719 &  x725 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x761 &  x764 &  x767 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x809 &  x811 &  x818 &  x824 &  x827 &  x830 &  x832 &  x833 &  x839 &  x845 &  x848 &  x854 &  x857 &  x863 &  x866 &  x877 &  x881 &  x884 &  x887 &  x893 &  x896 &  x905 &  x908 &  x910 &  x917 &  x923 &  x926 &  x944 &  x947 &  x949 &  x950 &  x959 &  x962 &  x971 &  x977 &  x983 &  x988 &  x989 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1019 &  x1027 &  x1028 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1064 &  x1066 &  x1070 &  x1073 &  x1076 &  x1079 &  x1091 &  x1094 &  x1103 &  x1106 &  x1112 &  x1121 &  x1124 &  x1130 & ~x99 & ~x144 & ~x183 & ~x222 & ~x294 & ~x741 & ~x780 & ~x819 & ~x858 & ~x897 & ~x936 & ~x975 & ~x1053;
assign c0262 =  x2 &  x5 &  x8 &  x14 &  x23 &  x26 &  x29 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x59 &  x62 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x149 &  x155 &  x158 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x197 &  x200 &  x203 &  x206 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x239 &  x242 &  x245 &  x248 &  x254 &  x263 &  x266 &  x269 &  x272 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x314 &  x317 &  x320 &  x326 &  x329 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x377 &  x383 &  x386 &  x389 &  x392 &  x395 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x428 &  x431 &  x434 &  x440 &  x446 &  x449 &  x452 &  x455 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x488 &  x491 &  x494 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x566 &  x572 &  x578 &  x584 &  x587 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x701 &  x703 &  x704 &  x707 &  x710 &  x713 &  x716 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x764 &  x770 &  x776 &  x779 &  x781 &  x785 &  x788 &  x794 &  x803 &  x812 &  x815 &  x818 &  x820 &  x821 &  x824 &  x827 &  x830 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x898 &  x899 &  x902 &  x905 &  x908 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x936 &  x938 &  x940 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x962 &  x965 &  x968 &  x974 &  x975 &  x976 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1015 &  x1016 &  x1018 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1054 &  x1055 &  x1057 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x393 & ~x432 & ~x474 & ~x513 & ~x549 & ~x837 & ~x972 & ~x1011 & ~x1050;
assign c0264 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x47 &  x53 &  x59 &  x62 &  x68 &  x74 &  x77 &  x80 &  x86 &  x89 &  x95 &  x98 &  x101 &  x104 &  x107 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x134 &  x143 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x170 &  x173 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x209 &  x212 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x254 &  x257 &  x263 &  x266 &  x269 &  x275 &  x278 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x325 &  x326 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x356 &  x359 &  x362 &  x365 &  x374 &  x377 &  x380 &  x383 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x557 &  x560 &  x563 &  x566 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x632 &  x635 &  x638 &  x641 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x703 &  x707 &  x710 &  x713 &  x716 &  x722 &  x725 &  x728 &  x731 &  x737 &  x740 &  x743 &  x749 &  x755 &  x758 &  x764 &  x767 &  x773 &  x776 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x820 &  x821 &  x823 &  x824 &  x830 &  x833 &  x836 &  x842 &  x845 &  x848 &  x851 &  x854 &  x859 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x896 &  x899 &  x901 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x929 &  x935 &  x937 &  x938 &  x939 &  x940 &  x941 &  x956 &  x959 &  x974 &  x976 &  x979 &  x983 &  x986 &  x992 &  x994 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1033 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1057 &  x1058 &  x1061 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1111 &  x1112 &  x1118 &  x1127 &  x1130 & ~x648;
assign c0266 =  x2 &  x5 &  x8 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x312 &  x313 &  x314 &  x317 &  x320 &  x323 &  x332 &  x335 &  x344 &  x347 &  x350 &  x351 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x404 &  x410 &  x413 &  x419 &  x422 &  x425 &  x430 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x455 &  x458 &  x461 &  x464 &  x467 &  x469 &  x470 &  x473 &  x479 &  x485 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x508 &  x509 &  x512 &  x515 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x581 &  x584 &  x590 &  x593 &  x596 &  x602 &  x605 &  x608 &  x617 &  x620 &  x626 &  x629 &  x632 &  x638 &  x644 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x667 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x698 &  x701 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x731 &  x734 &  x737 &  x740 &  x743 &  x745 &  x749 &  x752 &  x755 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x827 &  x836 &  x839 &  x842 &  x845 &  x848 &  x857 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x908 &  x914 &  x916 &  x917 &  x920 &  x923 &  x929 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x977 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x336 & ~x357 & ~x477 & ~x555;
assign c0268 =  x14 &  x17 &  x20 &  x23 &  x29 &  x32 &  x35 &  x38 &  x41 &  x50 &  x56 &  x59 &  x62 &  x71 &  x77 &  x80 &  x83 &  x86 &  x92 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x125 &  x137 &  x143 &  x146 &  x149 &  x152 &  x155 &  x164 &  x170 &  x182 &  x188 &  x191 &  x194 &  x197 &  x203 &  x206 &  x209 &  x212 &  x221 &  x224 &  x227 &  x236 &  x239 &  x251 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x284 &  x287 &  x290 &  x296 &  x305 &  x308 &  x311 &  x317 &  x323 &  x326 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x377 &  x380 &  x383 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x419 &  x431 &  x440 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x472 &  x473 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x511 &  x512 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x542 &  x545 &  x548 &  x549 &  x550 &  x551 &  x557 &  x563 &  x566 &  x578 &  x581 &  x584 &  x587 &  x589 &  x590 &  x596 &  x599 &  x611 &  x620 &  x623 &  x627 &  x628 &  x629 &  x632 &  x635 &  x638 &  x641 &  x650 &  x656 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x686 &  x689 &  x695 &  x701 &  x707 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x749 &  x752 &  x754 &  x758 &  x764 &  x767 &  x773 &  x779 &  x782 &  x785 &  x788 &  x791 &  x800 &  x806 &  x809 &  x812 &  x818 &  x821 &  x824 &  x830 &  x832 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x916 &  x929 &  x932 &  x935 &  x941 &  x947 &  x950 &  x953 &  x955 &  x956 &  x959 &  x962 &  x968 &  x971 &  x977 &  x983 &  x986 &  x989 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1130 & ~x318 & ~x333 & ~x357 & ~x702;
assign c0270 =  x2 &  x4 &  x8 &  x10 &  x11 &  x17 &  x20 &  x26 &  x32 &  x38 &  x43 &  x44 &  x47 &  x59 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x94 &  x98 &  x113 &  x116 &  x119 &  x122 &  x125 &  x131 &  x133 &  x134 &  x137 &  x146 &  x149 &  x155 &  x157 &  x158 &  x161 &  x164 &  x167 &  x173 &  x179 &  x182 &  x188 &  x191 &  x197 &  x200 &  x206 &  x212 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x251 &  x254 &  x257 &  x263 &  x266 &  x269 &  x272 &  x275 &  x281 &  x296 &  x302 &  x305 &  x311 &  x314 &  x317 &  x320 &  x329 &  x332 &  x335 &  x341 &  x350 &  x365 &  x371 &  x377 &  x380 &  x383 &  x386 &  x392 &  x395 &  x398 &  x407 &  x416 &  x433 &  x434 &  x437 &  x443 &  x446 &  x449 &  x458 &  x461 &  x464 &  x467 &  x470 &  x472 &  x476 &  x479 &  x482 &  x485 &  x488 &  x494 &  x497 &  x500 &  x503 &  x506 &  x511 &  x515 &  x518 &  x521 &  x529 &  x530 &  x536 &  x539 &  x545 &  x551 &  x554 &  x560 &  x568 &  x569 &  x572 &  x575 &  x581 &  x584 &  x590 &  x593 &  x596 &  x614 &  x623 &  x626 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x689 &  x692 &  x695 &  x698 &  x710 &  x719 &  x722 &  x725 &  x728 &  x731 &  x737 &  x740 &  x743 &  x746 &  x757 &  x767 &  x770 &  x776 &  x782 &  x785 &  x791 &  x794 &  x797 &  x803 &  x809 &  x812 &  x815 &  x818 &  x821 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x899 &  x905 &  x914 &  x917 &  x929 &  x935 &  x941 &  x944 &  x947 &  x965 &  x968 &  x977 &  x980 &  x986 &  x989 &  x995 &  x998 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1030 &  x1031 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1073 &  x1075 &  x1076 &  x1079 &  x1088 &  x1090 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1108 &  x1114 &  x1118 &  x1124 &  x1130;
assign c0272 =  x2 &  x5 &  x8 &  x17 &  x20 &  x29 &  x32 &  x35 &  x38 &  x44 &  x47 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x86 &  x92 &  x101 &  x113 &  x119 &  x125 &  x131 &  x134 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x257 &  x260 &  x266 &  x269 &  x272 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x326 &  x329 &  x335 &  x338 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x383 &  x386 &  x395 &  x404 &  x407 &  x413 &  x416 &  x419 &  x422 &  x428 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x497 &  x500 &  x506 &  x509 &  x518 &  x521 &  x527 &  x530 &  x536 &  x539 &  x545 &  x547 &  x548 &  x557 &  x560 &  x569 &  x572 &  x575 &  x578 &  x580 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x617 &  x619 &  x620 &  x623 &  x625 &  x632 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x703 &  x704 &  x707 &  x710 &  x713 &  x716 &  x722 &  x725 &  x731 &  x734 &  x737 &  x740 &  x742 &  x746 &  x752 &  x755 &  x758 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x797 &  x803 &  x808 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x893 &  x902 &  x908 &  x914 &  x917 &  x923 &  x926 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x956 &  x965 &  x968 &  x971 &  x974 &  x980 &  x983 &  x992 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1046 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1127 &  x1130 & ~x81 & ~x120 & ~x159 & ~x276 & ~x315 & ~x393 & ~x432 & ~x489 & ~x552 & ~x591;
assign c0274 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x23 &  x29 &  x32 &  x35 &  x41 &  x44 &  x47 &  x53 &  x55 &  x56 &  x59 &  x62 &  x65 &  x68 &  x77 &  x80 &  x92 &  x95 &  x98 &  x101 &  x107 &  x110 &  x112 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x143 &  x146 &  x149 &  x151 &  x152 &  x158 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x191 &  x194 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x230 &  x236 &  x239 &  x242 &  x245 &  x257 &  x263 &  x266 &  x272 &  x278 &  x281 &  x284 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x317 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x350 &  x353 &  x356 &  x359 &  x362 &  x371 &  x380 &  x383 &  x386 &  x389 &  x398 &  x401 &  x404 &  x407 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x455 &  x464 &  x470 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x523 &  x524 &  x536 &  x539 &  x542 &  x548 &  x554 &  x557 &  x560 &  x562 &  x566 &  x569 &  x574 &  x575 &  x578 &  x584 &  x590 &  x593 &  x596 &  x599 &  x602 &  x608 &  x614 &  x617 &  x623 &  x629 &  x632 &  x635 &  x638 &  x640 &  x641 &  x644 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x679 &  x680 &  x683 &  x686 &  x695 &  x698 &  x701 &  x704 &  x707 &  x713 &  x718 &  x719 &  x725 &  x728 &  x730 &  x731 &  x737 &  x746 &  x749 &  x755 &  x757 &  x758 &  x761 &  x764 &  x769 &  x773 &  x776 &  x779 &  x785 &  x791 &  x797 &  x800 &  x803 &  x806 &  x808 &  x809 &  x812 &  x814 &  x818 &  x821 &  x824 &  x827 &  x833 &  x839 &  x842 &  x845 &  x848 &  x854 &  x857 &  x860 &  x863 &  x866 &  x872 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x905 &  x908 &  x917 &  x920 &  x923 &  x924 &  x925 &  x926 &  x932 &  x935 &  x938 &  x950 &  x953 &  x956 &  x959 &  x964 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x998 &  x1001 &  x1004 &  x1010 &  x1016 &  x1019 &  x1022 &  x1028 &  x1031 &  x1037 &  x1040 &  x1042 &  x1043 &  x1046 &  x1049 &  x1058 &  x1061 &  x1067 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1112 &  x1118 &  x1124 &  x1127 &  x1130;
assign c0276 =  x8 &  x14 &  x50 &  x53 &  x59 &  x62 &  x101 &  x104 &  x110 &  x113 &  x119 &  x128 &  x146 &  x155 &  x161 &  x164 &  x170 &  x173 &  x188 &  x191 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x221 &  x239 &  x245 &  x257 &  x278 &  x290 &  x299 &  x302 &  x308 &  x317 &  x329 &  x347 &  x350 &  x359 &  x365 &  x368 &  x383 &  x389 &  x392 &  x398 &  x407 &  x410 &  x431 &  x443 &  x481 &  x484 &  x494 &  x509 &  x515 &  x518 &  x521 &  x523 &  x524 &  x527 &  x542 &  x551 &  x554 &  x557 &  x560 &  x562 &  x566 &  x572 &  x578 &  x587 &  x599 &  x602 &  x611 &  x614 &  x620 &  x623 &  x629 &  x647 &  x656 &  x662 &  x663 &  x665 &  x674 &  x680 &  x686 &  x703 &  x707 &  x710 &  x725 &  x728 &  x737 &  x749 &  x752 &  x755 &  x779 &  x782 &  x794 &  x800 &  x812 &  x836 &  x842 &  x848 &  x851 &  x857 &  x878 &  x893 &  x900 &  x902 &  x908 &  x911 &  x923 &  x929 &  x938 &  x939 &  x940 &  x941 &  x944 &  x962 &  x965 &  x971 &  x976 &  x986 &  x998 &  x1007 &  x1010 &  x1013 &  x1017 &  x1019 &  x1022 &  x1025 &  x1037 &  x1040 &  x1046 &  x1057 &  x1058 &  x1073 &  x1076 &  x1079 &  x1096 &  x1109 &  x1115 &  x1121 & ~x669 & ~x708;
assign c0278 =  x11 &  x17 &  x20 &  x23 &  x29 &  x32 &  x35 &  x44 &  x47 &  x50 &  x53 &  x65 &  x68 &  x77 &  x86 &  x95 &  x98 &  x104 &  x107 &  x113 &  x122 &  x125 &  x128 &  x131 &  x137 &  x140 &  x152 &  x155 &  x157 &  x160 &  x164 &  x167 &  x173 &  x179 &  x185 &  x188 &  x191 &  x194 &  x195 &  x196 &  x197 &  x200 &  x206 &  x209 &  x215 &  x218 &  x227 &  x230 &  x238 &  x239 &  x242 &  x254 &  x257 &  x260 &  x269 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x323 &  x326 &  x329 &  x335 &  x338 &  x341 &  x347 &  x350 &  x352 &  x353 &  x356 &  x365 &  x371 &  x377 &  x383 &  x386 &  x389 &  x392 &  x394 &  x398 &  x413 &  x425 &  x433 &  x434 &  x437 &  x440 &  x443 &  x446 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x472 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x512 &  x515 &  x518 &  x524 &  x530 &  x533 &  x536 &  x539 &  x545 &  x548 &  x551 &  x557 &  x563 &  x566 &  x572 &  x578 &  x581 &  x584 &  x587 &  x593 &  x596 &  x602 &  x617 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x647 &  x653 &  x656 &  x659 &  x671 &  x679 &  x680 &  x683 &  x689 &  x698 &  x707 &  x716 &  x718 &  x719 &  x722 &  x728 &  x731 &  x734 &  x737 &  x740 &  x752 &  x755 &  x758 &  x767 &  x770 &  x776 &  x785 &  x788 &  x803 &  x806 &  x809 &  x815 &  x821 &  x824 &  x833 &  x836 &  x839 &  x842 &  x845 &  x851 &  x863 &  x866 &  x881 &  x887 &  x890 &  x896 &  x899 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x932 &  x935 &  x938 &  x950 &  x956 &  x959 &  x971 &  x974 &  x980 &  x983 &  x986 &  x989 &  x995 &  x998 &  x1004 &  x1019 &  x1022 &  x1034 &  x1043 &  x1046 &  x1049 &  x1058 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1112 &  x1115 &  x1118 &  x1130 & ~x240 & ~x999 & ~x1083;
assign c0280 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x245 &  x251 &  x254 &  x257 &  x260 &  x266 &  x272 &  x275 &  x281 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x314 &  x317 &  x320 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x472 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x511 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x550 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x713 &  x716 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x854 &  x857 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x901 &  x902 &  x905 &  x908 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x935 &  x938 &  x940 &  x941 &  x944 &  x947 &  x950 &  x956 &  x959 &  x962 &  x968 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x27 & ~x66 & ~x105 & ~x168 & ~x201 & ~x207 & ~x210 & ~x249 & ~x495;
assign c0282 =  x5 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x80 &  x82 &  x83 &  x86 &  x89 &  x92 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x118 &  x122 &  x128 &  x134 &  x140 &  x143 &  x146 &  x149 &  x155 &  x156 &  x157 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x188 &  x191 &  x194 &  x195 &  x196 &  x197 &  x199 &  x200 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x235 &  x236 &  x238 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x272 &  x274 &  x275 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x317 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x355 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x380 &  x383 &  x386 &  x389 &  x392 &  x393 &  x395 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x431 &  x432 &  x433 &  x434 &  x437 &  x440 &  x443 &  x446 &  x455 &  x461 &  x464 &  x467 &  x470 &  x472 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x511 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x542 &  x550 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x656 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x698 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x728 &  x731 &  x734 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x760 &  x761 &  x764 &  x767 &  x770 &  x776 &  x779 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x827 &  x836 &  x839 &  x842 &  x845 &  x848 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x920 &  x923 &  x929 &  x932 &  x935 &  x941 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x983 &  x986 &  x989 &  x992 &  x998 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1124 &  x1127 &  x1130 & ~x546 & ~x585 & ~x663 & ~x819;
assign c0284 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x413 &  x416 &  x422 &  x425 &  x428 &  x430 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x467 &  x469 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x508 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x547 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x613 &  x614 &  x617 &  x620 &  x623 &  x625 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x667 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x698 &  x701 &  x703 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x742 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x198 & ~x237 & ~x453 & ~x474 & ~x492 & ~x513 & ~x531 & ~x552 & ~x570 & ~x591;
assign c0286 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x83 &  x86 &  x89 &  x92 &  x98 &  x101 &  x107 &  x110 &  x113 &  x119 &  x122 &  x128 &  x131 &  x134 &  x137 &  x140 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x227 &  x230 &  x236 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x263 &  x278 &  x281 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x320 &  x326 &  x332 &  x338 &  x341 &  x344 &  x352 &  x353 &  x356 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x391 &  x394 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x433 &  x440 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x470 &  x472 &  x476 &  x479 &  x482 &  x488 &  x494 &  x500 &  x503 &  x506 &  x509 &  x511 &  x512 &  x518 &  x521 &  x527 &  x533 &  x536 &  x538 &  x542 &  x545 &  x551 &  x557 &  x560 &  x566 &  x569 &  x575 &  x578 &  x581 &  x587 &  x589 &  x590 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x626 &  x628 &  x631 &  x632 &  x635 &  x641 &  x644 &  x647 &  x649 &  x656 &  x662 &  x665 &  x667 &  x670 &  x671 &  x674 &  x677 &  x680 &  x683 &  x685 &  x686 &  x689 &  x692 &  x698 &  x709 &  x710 &  x713 &  x716 &  x719 &  x728 &  x731 &  x734 &  x737 &  x743 &  x746 &  x749 &  x755 &  x758 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x785 &  x787 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x805 &  x806 &  x811 &  x812 &  x815 &  x818 &  x824 &  x826 &  x832 &  x833 &  x836 &  x839 &  x844 &  x845 &  x848 &  x851 &  x854 &  x860 &  x866 &  x871 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x949 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x988 &  x992 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1027 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1079 &  x1085 &  x1094 &  x1097 &  x1100 &  x1105 &  x1106 &  x1109 &  x1115 &  x1121 &  x1127;
assign c0288 =  x2 &  x5 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x134 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x383 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x410 &  x413 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x584 &  x587 &  x590 &  x596 &  x599 &  x602 &  x605 &  x611 &  x614 &  x617 &  x620 &  x623 &  x625 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x667 &  x668 &  x671 &  x674 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x701 &  x703 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x742 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x781 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x820 &  x821 &  x822 &  x823 &  x824 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x854 &  x857 &  x860 &  x861 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x898 &  x899 &  x900 &  x901 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x937 &  x938 &  x939 &  x940 &  x941 &  x944 &  x947 &  x950 &  x953 &  x959 &  x962 &  x968 &  x971 &  x974 &  x976 &  x977 &  x978 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1015 &  x1016 &  x1017 &  x1018 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1056 &  x1057 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1096 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x354 & ~x393 & ~x432 & ~x642 & ~x648;
assign c0290 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x56 &  x59 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x188 &  x191 &  x194 &  x197 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x242 &  x245 &  x248 &  x251 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x365 &  x368 &  x371 &  x374 &  x377 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x584 &  x585 &  x586 &  x587 &  x590 &  x593 &  x605 &  x611 &  x614 &  x617 &  x619 &  x620 &  x623 &  x624 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x659 &  x662 &  x663 &  x664 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x689 &  x692 &  x695 &  x701 &  x703 &  x707 &  x713 &  x719 &  x722 &  x728 &  x731 &  x734 &  x737 &  x742 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x764 &  x767 &  x769 &  x770 &  x773 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x808 &  x809 &  x812 &  x818 &  x820 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x851 &  x854 &  x859 &  x860 &  x862 &  x863 &  x866 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x914 &  x917 &  x920 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x977 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1028 &  x1034 &  x1037 &  x1040 &  x1046 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x537 & ~x792 & ~x831;
assign c0292 =  x41 &  x53 &  x182 &  x222 &  x335 &  x341 &  x344 &  x416 &  x445 &  x485 &  x502 &  x629 &  x680 &  x716 &  x761 &  x773 &  x776 &  x785 &  x812 &  x854 &  x863 &  x908 &  x1053 &  x1100 & ~x51 & ~x432 & ~x471 & ~x474;
assign c0294 =  x5 &  x8 &  x11 &  x14 &  x20 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x53 &  x56 &  x59 &  x73 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x101 &  x107 &  x110 &  x112 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x151 &  x152 &  x155 &  x158 &  x161 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x188 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x287 &  x293 &  x296 &  x302 &  x305 &  x314 &  x317 &  x320 &  x326 &  x329 &  x332 &  x335 &  x338 &  x344 &  x347 &  x350 &  x356 &  x362 &  x365 &  x371 &  x374 &  x377 &  x383 &  x386 &  x389 &  x395 &  x398 &  x407 &  x410 &  x413 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x452 &  x455 &  x458 &  x460 &  x461 &  x467 &  x473 &  x475 &  x476 &  x481 &  x485 &  x488 &  x491 &  x494 &  x497 &  x499 &  x500 &  x502 &  x503 &  x506 &  x512 &  x515 &  x520 &  x521 &  x524 &  x527 &  x533 &  x536 &  x541 &  x542 &  x545 &  x548 &  x554 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x580 &  x587 &  x590 &  x593 &  x598 &  x599 &  x602 &  x605 &  x611 &  x614 &  x617 &  x620 &  x629 &  x632 &  x635 &  x638 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x679 &  x683 &  x686 &  x695 &  x698 &  x707 &  x710 &  x713 &  x716 &  x718 &  x719 &  x731 &  x734 &  x737 &  x739 &  x740 &  x743 &  x746 &  x752 &  x758 &  x760 &  x761 &  x767 &  x770 &  x773 &  x775 &  x776 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x799 &  x800 &  x809 &  x815 &  x818 &  x824 &  x830 &  x833 &  x836 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x866 &  x872 &  x878 &  x881 &  x887 &  x890 &  x893 &  x899 &  x902 &  x905 &  x920 &  x926 &  x929 &  x932 &  x938 &  x944 &  x947 &  x950 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x986 &  x989 &  x992 &  x998 &  x1001 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1070 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1118 &  x1124;
assign c0296 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x390 &  x391 &  x392 &  x394 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x430 &  x431 &  x433 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x469 &  x470 &  x472 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x508 &  x509 &  x511 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x547 &  x548 &  x550 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x589 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x623 &  x626 &  x628 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x667 &  x668 &  x671 &  x674 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x731 &  x734 &  x737 &  x740 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x782 &  x785 &  x788 &  x791 &  x793 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x832 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x926 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x357 & ~x375 & ~x396 & ~x435 & ~x516 & ~x555;
assign c0298 =  x2 &  x5 &  x8 &  x14 &  x17 &  x23 &  x26 &  x29 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x71 &  x74 &  x77 &  x83 &  x89 &  x92 &  x95 &  x98 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x140 &  x146 &  x152 &  x155 &  x161 &  x167 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x242 &  x248 &  x251 &  x260 &  x266 &  x269 &  x272 &  x278 &  x287 &  x290 &  x293 &  x296 &  x299 &  x305 &  x314 &  x317 &  x320 &  x323 &  x326 &  x335 &  x341 &  x344 &  x347 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x406 &  x407 &  x416 &  x422 &  x428 &  x431 &  x437 &  x445 &  x446 &  x449 &  x452 &  x458 &  x464 &  x467 &  x470 &  x476 &  x479 &  x482 &  x488 &  x491 &  x494 &  x497 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x533 &  x539 &  x542 &  x545 &  x547 &  x551 &  x554 &  x557 &  x560 &  x562 &  x566 &  x569 &  x575 &  x581 &  x584 &  x585 &  x586 &  x587 &  x590 &  x596 &  x599 &  x602 &  x608 &  x614 &  x620 &  x623 &  x624 &  x625 &  x629 &  x632 &  x635 &  x638 &  x641 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x663 &  x668 &  x671 &  x674 &  x677 &  x686 &  x695 &  x698 &  x701 &  x703 &  x707 &  x710 &  x713 &  x719 &  x722 &  x725 &  x728 &  x737 &  x740 &  x742 &  x746 &  x749 &  x752 &  x755 &  x761 &  x764 &  x770 &  x776 &  x779 &  x781 &  x782 &  x785 &  x797 &  x803 &  x806 &  x809 &  x812 &  x815 &  x820 &  x821 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x859 &  x860 &  x866 &  x869 &  x872 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x898 &  x899 &  x901 &  x902 &  x905 &  x911 &  x917 &  x920 &  x923 &  x935 &  x938 &  x950 &  x953 &  x959 &  x962 &  x965 &  x971 &  x974 &  x979 &  x983 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1013 &  x1015 &  x1018 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1052 &  x1054 &  x1055 &  x1058 &  x1061 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x432 & ~x471 & ~x630 & ~x669;
assign c01 =  x8 &  x11 &  x100 &  x116 &  x179 &  x181 &  x194 &  x338 &  x359 &  x376 &  x389 &  x536 &  x599 &  x617 &  x653 &  x779 &  x818 &  x860 &  x868 &  x896 &  x983 &  x1091 & ~x660 & ~x843;
assign c03 =  x17 &  x20 &  x23 &  x50 &  x83 &  x101 &  x116 &  x140 &  x146 &  x167 &  x170 &  x173 &  x203 &  x206 &  x209 &  x218 &  x236 &  x242 &  x245 &  x254 &  x275 &  x281 &  x296 &  x299 &  x323 &  x332 &  x347 &  x356 &  x359 &  x374 &  x431 &  x437 &  x461 &  x467 &  x500 &  x503 &  x518 &  x521 &  x533 &  x536 &  x545 &  x551 &  x554 &  x560 &  x572 &  x595 &  x629 &  x632 &  x634 &  x635 &  x647 &  x665 &  x671 &  x740 &  x743 &  x746 &  x758 &  x764 &  x776 &  x794 &  x800 &  x809 &  x821 &  x827 &  x830 &  x851 &  x860 &  x863 &  x869 &  x884 &  x917 &  x929 &  x935 &  x953 &  x989 &  x992 &  x998 &  x1025 &  x1037 &  x1043 &  x1049 &  x1067 &  x1097 &  x1100 &  x1106 &  x1118 &  x1124 &  x1127 &  x1130 & ~x273 & ~x312 & ~x936 & ~x1098;
assign c05 =  x122 &  x485 &  x614 &  x745 &  x779 &  x800 &  x911 &  x1054 &  x1067 & ~x156 & ~x507 & ~x966 & ~x1104;
assign c07 =  x2 &  x17 &  x23 &  x26 &  x35 &  x44 &  x47 &  x68 &  x71 &  x74 &  x80 &  x92 &  x110 &  x113 &  x116 &  x140 &  x149 &  x152 &  x170 &  x179 &  x185 &  x194 &  x203 &  x206 &  x209 &  x221 &  x224 &  x233 &  x245 &  x251 &  x254 &  x269 &  x275 &  x278 &  x293 &  x308 &  x314 &  x320 &  x326 &  x332 &  x335 &  x338 &  x344 &  x347 &  x350 &  x353 &  x362 &  x365 &  x374 &  x380 &  x392 &  x401 &  x407 &  x422 &  x425 &  x428 &  x440 &  x443 &  x448 &  x455 &  x458 &  x461 &  x470 &  x476 &  x482 &  x485 &  x497 &  x503 &  x509 &  x512 &  x518 &  x539 &  x545 &  x554 &  x557 &  x563 &  x569 &  x575 &  x593 &  x602 &  x608 &  x611 &  x617 &  x641 &  x644 &  x659 &  x667 &  x677 &  x692 &  x698 &  x701 &  x713 &  x737 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x767 &  x776 &  x782 &  x785 &  x797 &  x803 &  x806 &  x809 &  x815 &  x821 &  x824 &  x833 &  x836 &  x845 &  x851 &  x854 &  x857 &  x866 &  x869 &  x875 &  x878 &  x881 &  x893 &  x899 &  x923 &  x926 &  x935 &  x950 &  x959 &  x983 &  x992 &  x1013 &  x1016 &  x1019 &  x1031 &  x1046 &  x1049 &  x1067 &  x1070 &  x1073 &  x1076 &  x1085 &  x1088 &  x1100 &  x1106 &  x1112 &  x1115 &  x1118 & ~x156 & ~x234 & ~x915 & ~x1035 & ~x1038;
assign c09 =  x104 &  x107 &  x140 &  x194 &  x203 &  x272 &  x359 &  x583 &  x632 &  x668 &  x788 &  x811 &  x947 &  x1070 &  x1124 & ~x372 & ~x663 & ~x666 & ~x834;
assign c011 =  x29 &  x44 &  x100 &  x101 &  x113 &  x116 &  x119 &  x125 &  x143 &  x152 &  x176 &  x179 &  x230 &  x266 &  x275 &  x281 &  x284 &  x316 &  x338 &  x356 &  x368 &  x416 &  x446 &  x488 &  x512 &  x518 &  x527 &  x548 &  x569 &  x572 &  x605 &  x620 &  x623 &  x632 &  x689 &  x767 &  x770 &  x797 &  x806 &  x815 &  x851 &  x857 &  x935 &  x1010 &  x1037 &  x1064 &  x1100 &  x1109 & ~x327 & ~x450 & ~x627 & ~x705;
assign c013 =  x56 &  x62 &  x74 &  x131 &  x349 &  x380 &  x437 &  x515 &  x599 &  x689 &  x710 &  x755 &  x758 &  x868 &  x905 &  x908 &  x946 &  x977 &  x1034 & ~x117 & ~x429 & ~x468 & ~x507 & ~x810;
assign c015 =  x47 &  x59 &  x168 &  x797 &  x920 & ~x399 & ~x438 & ~x585 & ~x756 & ~x885;
assign c017 = ~x251;
assign c019 =  x134 &  x206 &  x356 &  x413 &  x425 &  x620 &  x680 &  x774 &  x941 &  x1001 &  x1088 &  x1115 & ~x543 & ~x621 & ~x714;
assign c021 =  x5 &  x41 &  x44 &  x59 &  x68 &  x104 &  x110 &  x119 &  x131 &  x142 &  x158 &  x188 &  x233 &  x290 &  x302 &  x308 &  x344 &  x350 &  x356 &  x359 &  x362 &  x395 &  x422 &  x428 &  x440 &  x446 &  x448 &  x452 &  x458 &  x470 &  x476 &  x485 &  x497 &  x503 &  x524 &  x542 &  x548 &  x554 &  x563 &  x602 &  x608 &  x632 &  x635 &  x638 &  x650 &  x665 &  x680 &  x683 &  x695 &  x722 &  x728 &  x737 &  x743 &  x749 &  x785 &  x797 &  x857 &  x890 &  x935 &  x938 &  x962 &  x1025 &  x1040 &  x1043 &  x1046 &  x1049 &  x1064 &  x1085 &  x1094 &  x1106 &  x1109 &  x1115 &  x1130 & ~x195 & ~x234 & ~x312 & ~x1017;
assign c023 =  x8 &  x23 &  x32 &  x50 &  x83 &  x98 &  x104 &  x125 &  x142 &  x149 &  x164 &  x179 &  x200 &  x253 &  x292 &  x331 &  x332 &  x347 &  x386 &  x410 &  x428 &  x448 &  x449 &  x461 &  x464 &  x497 &  x530 &  x560 &  x620 &  x635 &  x641 &  x644 &  x650 &  x656 &  x722 &  x746 &  x755 &  x761 &  x806 &  x815 &  x866 &  x905 &  x1007 &  x1016 &  x1049 &  x1076 &  x1079 & ~x1017;
assign c025 =  x292 &  x418 & ~x0 & ~x978;
assign c027 =  x32 &  x40 &  x50 &  x59 &  x68 &  x80 &  x125 &  x139 &  x149 &  x167 &  x182 &  x191 &  x224 &  x269 &  x287 &  x311 &  x355 &  x362 &  x365 &  x368 &  x395 &  x440 &  x455 &  x482 &  x560 &  x566 &  x575 &  x584 &  x643 &  x647 &  x650 &  x716 &  x740 &  x746 &  x758 &  x779 &  x785 &  x791 &  x814 &  x818 &  x827 &  x838 &  x842 &  x844 &  x883 &  x890 &  x923 &  x941 &  x950 &  x974 &  x983 &  x1039 &  x1084 &  x1094;
assign c029 =  x23 &  x107 &  x176 &  x185 &  x284 &  x287 &  x335 &  x374 &  x391 &  x517 &  x893 &  x917 &  x1040 &  x1066 &  x1072 &  x1105 & ~x309 & ~x783 & ~x1053;
assign c031 = ~x39 & ~x165 & ~x321 & ~x660 & ~x699;
assign c033 =  x116 &  x439 &  x688 &  x758 &  x778 &  x893 &  x1109 & ~x642 & ~x717 & ~x984;
assign c035 =  x99 &  x210 &  x334 &  x529 & ~x888;
assign c037 =  x5 &  x11 &  x23 &  x38 &  x50 &  x53 &  x59 &  x80 &  x83 &  x92 &  x113 &  x116 &  x137 &  x140 &  x149 &  x200 &  x206 &  x218 &  x221 &  x248 &  x254 &  x257 &  x263 &  x272 &  x290 &  x296 &  x326 &  x341 &  x344 &  x371 &  x380 &  x386 &  x389 &  x395 &  x401 &  x404 &  x410 &  x419 &  x440 &  x452 &  x464 &  x467 &  x470 &  x482 &  x512 &  x515 &  x521 &  x533 &  x557 &  x578 &  x596 &  x599 &  x623 &  x644 &  x656 &  x665 &  x671 &  x674 &  x692 &  x695 &  x698 &  x707 &  x710 &  x713 &  x722 &  x734 &  x755 &  x764 &  x776 &  x785 &  x803 &  x824 &  x830 &  x839 &  x851 &  x863 &  x893 &  x896 &  x905 &  x935 &  x950 &  x959 &  x962 &  x980 &  x986 &  x1019 &  x1025 &  x1028 &  x1031 &  x1046 &  x1049 &  x1052 &  x1061 &  x1070 &  x1076 &  x1100 &  x1106 &  x1112 &  x1115 &  x1130 & ~x156 & ~x351 & ~x468 & ~x507 & ~x951 & ~x993 & ~x1104;
assign c039 =  x529 & ~x384 & ~x952 & ~x1114;
assign c041 =  x92 &  x581 & ~x265 & ~x706;
assign c043 =  x32 &  x38 &  x56 &  x77 &  x92 &  x98 &  x101 &  x122 &  x125 &  x131 &  x194 &  x200 &  x218 &  x220 &  x308 &  x329 &  x350 &  x370 &  x380 &  x392 &  x409 &  x434 &  x449 &  x458 &  x467 &  x470 &  x485 &  x503 &  x527 &  x575 &  x584 &  x614 &  x641 &  x644 &  x686 &  x701 &  x722 &  x755 &  x761 &  x773 &  x803 &  x845 &  x881 &  x1010 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 & ~x726 & ~x804 & ~x1056;
assign c045 =  x8 &  x928 & ~x403 & ~x678 & ~x681;
assign c047 =  x215 &  x389 &  x416 &  x455 &  x728 &  x817 &  x923 &  x1049 &  x1058 & ~x465 & ~x642 & ~x861 & ~x978;
assign c049 = ~x374;
assign c051 =  x224 &  x341 &  x367 &  x470 &  x499 &  x833 &  x907 &  x946 &  x977 & ~x429 & ~x850 & ~x966;
assign c053 =  x22 &  x74 &  x101 &  x217 &  x233 &  x407 &  x419 &  x551 &  x595 &  x683 &  x689 &  x698 &  x839 &  x853 &  x931 &  x932 &  x935 &  x968 &  x974 &  x983 &  x1043 &  x1046 &  x1075 &  x1108 &  x1126 & ~x939;
assign c055 = ~x315 & ~x390 & ~x559;
assign c057 =  x26 &  x38 &  x80 &  x86 &  x89 &  x98 &  x146 &  x173 &  x176 &  x293 &  x341 &  x347 &  x395 &  x494 &  x578 &  x584 &  x596 &  x611 &  x659 &  x674 &  x803 &  x806 &  x815 &  x821 &  x863 &  x872 &  x899 &  x935 &  x941 &  x992 &  x1118 & ~x111 & ~x156 & ~x537 & ~x741 & ~x822;
assign c059 =  x508 & ~x609 & ~x667;
assign c061 =  x38 &  x65 &  x121 &  x236 &  x241 &  x245 &  x344 &  x431 &  x589 &  x620 &  x1058 &  x1076 &  x1124 &  x1127 & ~x429 & ~x981;
assign c063 =  x227 &  x263 &  x278 &  x284 &  x302 &  x326 &  x335 &  x350 &  x362 &  x377 &  x380 &  x389 &  x443 &  x446 &  x458 &  x475 &  x485 &  x524 &  x545 &  x548 &  x551 &  x575 &  x581 &  x599 &  x662 &  x689 &  x695 &  x785 &  x881 &  x887 &  x911 &  x971 &  x983 &  x992 &  x1004 &  x1015 &  x1057 &  x1061 &  x1085 & ~x546 & ~x633 & ~x711 & ~x714 & ~x771;
assign c065 =  x293 &  x386 &  x434 &  x664 &  x703 &  x746 &  x829 & ~x429 & ~x468 & ~x639 & ~x960 & ~x999;
assign c067 = ~x843 & ~x940;
assign c069 =  x8 &  x121 &  x164 &  x344 &  x398 &  x461 &  x554 &  x578 &  x611 &  x710 &  x718 &  x776 &  x860 &  x869 &  x1046 &  x1103 &  x1115 & ~x318 & ~x357 & ~x667 & ~x744;
assign c071 =  x203 &  x511 &  x739 &  x1040 & ~x156 & ~x783;
assign c073 =  x198 &  x1084 &  x1120 & ~x114 & ~x549;
assign c075 = ~x312 & ~x655 & ~x678 & ~x699 & ~x876;
assign c077 =  x11 &  x14 &  x23 &  x50 &  x65 &  x83 &  x86 &  x113 &  x119 &  x152 &  x158 &  x161 &  x188 &  x221 &  x224 &  x236 &  x266 &  x280 &  x287 &  x302 &  x311 &  x320 &  x338 &  x365 &  x380 &  x386 &  x392 &  x398 &  x413 &  x416 &  x419 &  x500 &  x524 &  x596 &  x617 &  x671 &  x677 &  x683 &  x692 &  x734 &  x746 &  x770 &  x794 &  x803 &  x833 &  x836 &  x908 &  x932 &  x941 &  x953 &  x980 &  x986 &  x1001 &  x1010 &  x1013 &  x1028 &  x1037 &  x1049 &  x1070 &  x1088 &  x1124 & ~x231 & ~x232 & ~x783 & ~x822 & ~x861;
assign c079 =  x95 &  x404 &  x409 &  x628 &  x728 &  x773 &  x868 & ~x351 & ~x810 & ~x960 & ~x999;
assign c081 =  x47 &  x50 &  x77 &  x119 &  x122 &  x125 &  x146 &  x188 &  x233 &  x235 &  x254 &  x302 &  x383 &  x389 &  x392 &  x440 &  x452 &  x475 &  x527 &  x563 &  x605 &  x632 &  x668 &  x689 &  x707 &  x815 &  x914 &  x923 &  x928 &  x938 &  x956 &  x971 &  x977 &  x1016 &  x1127 & ~x558 & ~x597 & ~x819 & ~x834;
assign c083 =  x257 &  x262 &  x263 &  x604 & ~x612 & ~x739;
assign c085 =  x239 & ~x660 & ~x916 & ~x993 & ~x1032 & ~x1065;
assign c087 =  x115 &  x220 &  x259 &  x409 & ~x843 & ~x1095;
assign c089 =  x610 & ~x7 & ~x423 & ~x477 & ~x1113;
assign c091 =  x107 &  x209 &  x251 &  x428 &  x506 &  x617 &  x710 &  x1085 & ~x156 & ~x273 & ~x360 & ~x399 & ~x478;
assign c093 = ~x598 & ~x831;
assign c095 =  x100 &  x107 &  x302 &  x533 &  x587 &  x617 &  x764 &  x782 &  x803 &  x823 &  x827 &  x869 &  x901 & ~x705 & ~x822 & ~x936;
assign c097 = ~x156 & ~x1105;
assign c099 =  x800 & ~x492 & ~x706;
assign c0101 = ~x465 & ~x642 & ~x862;
assign c0103 = ~x116;
assign c0105 =  x50 &  x119 &  x128 &  x167 &  x191 &  x215 &  x224 &  x230 &  x253 &  x275 &  x292 &  x296 &  x341 &  x419 &  x461 &  x521 &  x584 &  x599 &  x608 &  x707 &  x782 &  x785 &  x788 &  x824 &  x842 &  x881 &  x950 &  x956 &  x992 &  x1016 &  x1019 &  x1067 &  x1115 &  x1127 & ~x729 & ~x840 & ~x978;
assign c0107 =  x17 &  x23 &  x59 &  x116 &  x122 &  x161 &  x188 &  x227 &  x233 &  x260 &  x281 &  x341 &  x350 &  x356 &  x455 &  x482 &  x500 &  x503 &  x506 &  x530 &  x551 &  x554 &  x560 &  x571 &  x581 &  x584 &  x599 &  x605 &  x617 &  x635 &  x653 &  x671 &  x689 &  x710 &  x722 &  x725 &  x728 &  x755 &  x758 &  x776 &  x779 &  x791 &  x911 &  x929 &  x938 &  x968 &  x971 &  x983 &  x1013 &  x1019 &  x1037 &  x1058 &  x1070 &  x1076 &  x1103 &  x1127 &  x1130 & ~x312 & ~x351 & ~x390 & ~x912 & ~x915 & ~x990 & ~x1074 & ~x1113;
assign c0109 =  x41 &  x329 &  x343 &  x346 &  x424 &  x527 &  x568 & ~x102 & ~x135 & ~x285 & ~x324 & ~x363 & ~x993 & ~x1071;
assign c0111 =  x436 & ~x640 & ~x939;
assign c0113 =  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x38 &  x41 &  x47 &  x50 &  x53 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x91 &  x92 &  x95 &  x98 &  x104 &  x110 &  x113 &  x119 &  x122 &  x125 &  x128 &  x134 &  x136 &  x137 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x212 &  x224 &  x227 &  x233 &  x236 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x275 &  x278 &  x281 &  x287 &  x290 &  x293 &  x299 &  x305 &  x311 &  x314 &  x317 &  x323 &  x329 &  x335 &  x338 &  x341 &  x344 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x389 &  x391 &  x395 &  x398 &  x401 &  x407 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x434 &  x440 &  x443 &  x446 &  x452 &  x455 &  x464 &  x470 &  x476 &  x479 &  x482 &  x485 &  x488 &  x494 &  x497 &  x500 &  x503 &  x509 &  x512 &  x515 &  x517 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x542 &  x545 &  x548 &  x551 &  x554 &  x556 &  x557 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x587 &  x593 &  x595 &  x608 &  x611 &  x614 &  x617 &  x623 &  x629 &  x632 &  x635 &  x638 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x665 &  x668 &  x674 &  x677 &  x680 &  x683 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x719 &  x722 &  x725 &  x728 &  x731 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x764 &  x770 &  x773 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x827 &  x833 &  x836 &  x839 &  x842 &  x851 &  x857 &  x863 &  x869 &  x872 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x980 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1088 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1124 &  x1127 &  x1130 & ~x381 & ~x537;
assign c0115 =  x337 & ~x36 & ~x922 & ~x1071;
assign c0117 =  x2 &  x8 &  x23 &  x50 &  x74 &  x80 &  x92 &  x98 &  x122 &  x128 &  x142 &  x182 &  x197 &  x209 &  x227 &  x254 &  x257 &  x296 &  x317 &  x332 &  x383 &  x407 &  x425 &  x428 &  x437 &  x446 &  x452 &  x467 &  x470 &  x482 &  x497 &  x509 &  x512 &  x524 &  x545 &  x560 &  x581 &  x638 &  x644 &  x662 &  x668 &  x686 &  x695 &  x707 &  x722 &  x785 &  x812 &  x827 &  x839 &  x884 &  x896 &  x911 &  x920 &  x929 &  x962 &  x1010 &  x1019 &  x1022 &  x1046 &  x1052 &  x1109 &  x1112 &  x1124 & ~x306 & ~x384 & ~x684 & ~x762 & ~x939 & ~x1017;
assign c0119 =  x136 & ~x282 & ~x462 & ~x1017;
assign c0121 =  x28 &  x80 &  x155 &  x331 &  x335 &  x548 &  x567 &  x607 &  x646 &  x1078;
assign c0123 = ~x164;
assign c0125 =  x5 &  x8 &  x29 &  x32 &  x41 &  x47 &  x56 &  x65 &  x74 &  x86 &  x116 &  x119 &  x122 &  x128 &  x134 &  x137 &  x140 &  x146 &  x152 &  x173 &  x179 &  x194 &  x200 &  x242 &  x245 &  x248 &  x257 &  x263 &  x272 &  x275 &  x278 &  x296 &  x311 &  x323 &  x341 &  x344 &  x347 &  x350 &  x356 &  x365 &  x374 &  x383 &  x389 &  x398 &  x410 &  x413 &  x416 &  x431 &  x446 &  x461 &  x503 &  x529 &  x533 &  x539 &  x545 &  x554 &  x566 &  x572 &  x590 &  x605 &  x611 &  x626 &  x647 &  x656 &  x680 &  x686 &  x689 &  x692 &  x707 &  x716 &  x731 &  x743 &  x758 &  x761 &  x764 &  x776 &  x785 &  x800 &  x812 &  x818 &  x833 &  x839 &  x851 &  x857 &  x860 &  x869 &  x875 &  x881 &  x890 &  x902 &  x911 &  x923 &  x935 &  x938 &  x947 &  x953 &  x956 &  x962 &  x965 &  x971 &  x983 &  x989 &  x992 &  x998 &  x1013 &  x1019 &  x1022 &  x1025 &  x1064 &  x1070 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1115 & ~x0 & ~x468 & ~x549 & ~x975;
assign c0127 =  x41 &  x44 &  x47 &  x53 &  x56 &  x59 &  x65 &  x68 &  x80 &  x83 &  x110 &  x122 &  x125 &  x134 &  x143 &  x167 &  x215 &  x242 &  x275 &  x281 &  x299 &  x305 &  x377 &  x401 &  x407 &  x422 &  x428 &  x434 &  x440 &  x473 &  x479 &  x485 &  x533 &  x548 &  x557 &  x560 &  x572 &  x653 &  x671 &  x686 &  x689 &  x701 &  x719 &  x722 &  x728 &  x737 &  x776 &  x779 &  x785 &  x818 &  x839 &  x941 &  x959 &  x962 &  x965 &  x974 &  x983 &  x986 &  x1007 &  x1010 &  x1049 &  x1091 &  x1100 &  x1103 &  x1124 &  x1127 & ~x0 & ~x507 & ~x627 & ~x975 & ~x1014;
assign c0129 = ~x492 & ~x628 & ~x1014;
assign c0131 =  x2 &  x8 &  x59 &  x65 &  x74 &  x146 &  x158 &  x161 &  x179 &  x200 &  x221 &  x326 &  x329 &  x332 &  x335 &  x341 &  x347 &  x350 &  x356 &  x425 &  x467 &  x488 &  x491 &  x497 &  x506 &  x509 &  x572 &  x589 &  x593 &  x596 &  x623 &  x635 &  x641 &  x686 &  x719 &  x725 &  x755 &  x767 &  x782 &  x791 &  x797 &  x824 &  x866 &  x881 &  x893 &  x911 &  x974 &  x1085 &  x1121 & ~x36 & ~x312 & ~x693 & ~x732 & ~x768 & ~x771 & ~x810;
assign c0133 =  x177 &  x250 &  x255 &  x892 & ~x1095;
assign c0135 = ~x681 & ~x715;
assign c0137 =  x19 &  x38 &  x80 &  x175 &  x595 &  x602 &  x620 &  x638 &  x715 &  x941 &  x986 &  x1055 &  x1078 & ~x813 & ~x1035;
assign c0139 =  x142 &  x181 &  x259 &  x544 &  x946 & ~x810 & ~x960;
assign c0141 =  x868 &  x872 & ~x654 & ~x772 & ~x1032;
assign c0143 =  x242 &  x251 &  x263 &  x365 &  x494 &  x644 &  x719 &  x857 &  x872 &  x1001 &  x1040 & ~x78 & ~x285 & ~x705 & ~x939;
assign c0145 =  x8 &  x86 &  x170 &  x188 &  x191 &  x194 &  x418 &  x422 &  x446 &  x482 &  x521 &  x617 &  x728 &  x731 &  x776 &  x812 &  x875 &  x881 &  x926 &  x940 &  x1013 &  x1052 &  x1094 &  x1109 & ~x204 & ~x282 & ~x360 & ~x399 & ~x556 & ~x594;
assign c0147 =  x65 &  x155 &  x179 &  x194 &  x254 &  x266 &  x272 &  x290 &  x293 &  x338 &  x371 &  x374 &  x383 &  x386 &  x398 &  x446 &  x506 &  x512 &  x539 &  x557 &  x563 &  x572 &  x602 &  x614 &  x620 &  x626 &  x628 &  x659 &  x668 &  x767 &  x782 &  x794 &  x827 &  x836 &  x848 &  x857 &  x881 &  x890 &  x926 &  x932 &  x938 &  x986 &  x992 &  x1007 &  x1043 &  x1061 &  x1094 & ~x312 & ~x525 & ~x861;
assign c0149 =  x5 &  x8 &  x11 &  x14 &  x26 &  x29 &  x32 &  x38 &  x41 &  x59 &  x62 &  x65 &  x68 &  x71 &  x83 &  x95 &  x104 &  x107 &  x113 &  x119 &  x125 &  x134 &  x140 &  x149 &  x152 &  x158 &  x170 &  x176 &  x179 &  x185 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x218 &  x227 &  x239 &  x248 &  x251 &  x254 &  x257 &  x281 &  x284 &  x293 &  x299 &  x302 &  x308 &  x326 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x371 &  x380 &  x386 &  x392 &  x395 &  x398 &  x401 &  x404 &  x416 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x449 &  x455 &  x467 &  x476 &  x479 &  x494 &  x497 &  x500 &  x503 &  x512 &  x518 &  x533 &  x539 &  x548 &  x551 &  x557 &  x563 &  x572 &  x575 &  x584 &  x593 &  x599 &  x602 &  x614 &  x620 &  x626 &  x629 &  x632 &  x638 &  x641 &  x647 &  x650 &  x656 &  x662 &  x665 &  x668 &  x671 &  x677 &  x686 &  x701 &  x704 &  x713 &  x716 &  x722 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x749 &  x755 &  x761 &  x764 &  x767 &  x770 &  x776 &  x779 &  x785 &  x794 &  x803 &  x806 &  x815 &  x818 &  x842 &  x848 &  x857 &  x860 &  x863 &  x866 &  x875 &  x881 &  x893 &  x899 &  x902 &  x905 &  x911 &  x914 &  x917 &  x920 &  x938 &  x944 &  x950 &  x956 &  x962 &  x971 &  x980 &  x986 &  x989 &  x992 &  x1010 &  x1013 &  x1016 &  x1028 &  x1034 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1064 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1115 &  x1127 &  x1130 & ~x585 & ~x628 & ~x1092;
assign c0151 =  x128 &  x184 &  x269 &  x404 &  x602 &  x1067 & ~x336 & ~x348 & ~x690 & ~x792 & ~x807;
assign c0153 = ~x503;
assign c0155 =  x152 &  x457 &  x631 &  x669 &  x950 &  x992 & ~x705 & ~x711 & ~x750;
assign c0157 = ~x91 & ~x225 & ~x261 & ~x381 & ~x627;
assign c0159 = ~x545;
assign c0163 =  x203 &  x397 &  x608 &  x1019 &  x1073 &  x1127 & ~x520 & ~x636 & ~x714;
assign c0165 =  x269 &  x398 &  x674 &  x797 &  x908 &  x1067 & ~x234 & ~x399 & ~x654 & ~x699 & ~x732 & ~x1074 & ~x1104;
assign c0167 =  x5 &  x17 &  x29 &  x32 &  x53 &  x68 &  x74 &  x80 &  x86 &  x89 &  x92 &  x107 &  x110 &  x113 &  x119 &  x125 &  x131 &  x140 &  x146 &  x149 &  x155 &  x158 &  x167 &  x176 &  x191 &  x203 &  x206 &  x218 &  x221 &  x224 &  x230 &  x242 &  x245 &  x257 &  x275 &  x284 &  x287 &  x293 &  x305 &  x311 &  x320 &  x323 &  x332 &  x341 &  x350 &  x356 &  x359 &  x368 &  x374 &  x389 &  x392 &  x401 &  x404 &  x416 &  x419 &  x422 &  x425 &  x431 &  x440 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x506 &  x512 &  x518 &  x527 &  x533 &  x536 &  x539 &  x542 &  x554 &  x560 &  x563 &  x572 &  x575 &  x584 &  x590 &  x596 &  x602 &  x605 &  x608 &  x614 &  x617 &  x629 &  x631 &  x632 &  x635 &  x641 &  x647 &  x650 &  x659 &  x665 &  x677 &  x686 &  x698 &  x701 &  x707 &  x713 &  x725 &  x728 &  x734 &  x743 &  x746 &  x752 &  x770 &  x773 &  x776 &  x785 &  x788 &  x791 &  x803 &  x812 &  x827 &  x830 &  x833 &  x836 &  x839 &  x848 &  x851 &  x860 &  x866 &  x869 &  x872 &  x875 &  x884 &  x896 &  x902 &  x905 &  x908 &  x917 &  x929 &  x935 &  x941 &  x944 &  x956 &  x959 &  x986 &  x992 &  x998 &  x1001 &  x1013 &  x1016 &  x1034 &  x1052 &  x1055 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1091 &  x1097 &  x1100 &  x1106 &  x1127 & ~x147 & ~x381 & ~x420 & ~x459 & ~x549 & ~x711;
assign c0169 =  x2 &  x8 &  x20 &  x23 &  x47 &  x65 &  x116 &  x137 &  x140 &  x146 &  x152 &  x164 &  x176 &  x185 &  x188 &  x191 &  x194 &  x197 &  x203 &  x206 &  x215 &  x269 &  x272 &  x275 &  x281 &  x302 &  x317 &  x320 &  x341 &  x365 &  x404 &  x422 &  x443 &  x470 &  x476 &  x479 &  x509 &  x512 &  x536 &  x551 &  x554 &  x566 &  x571 &  x587 &  x602 &  x611 &  x635 &  x644 &  x650 &  x680 &  x688 &  x698 &  x700 &  x701 &  x704 &  x710 &  x725 &  x737 &  x761 &  x767 &  x779 &  x785 &  x797 &  x824 &  x833 &  x839 &  x844 &  x845 &  x851 &  x856 &  x863 &  x884 &  x899 &  x902 &  x935 &  x947 &  x980 &  x989 &  x1025 &  x1045 &  x1052 &  x1055 &  x1061 &  x1067 &  x1082 &  x1091 &  x1100 &  x1109 & ~x246 & ~x525;
assign c0171 =  x184 &  x616 & ~x117 & ~x468 & ~x469 & ~x507 & ~x1113;
assign c0173 =  x29 &  x116 &  x160 &  x185 &  x218 &  x224 &  x239 &  x304 &  x310 &  x407 &  x415 &  x433 &  x458 &  x503 &  x554 &  x560 &  x581 &  x587 &  x683 &  x794 &  x875 &  x1028 & ~x195;
assign c0175 =  x17 &  x20 &  x23 &  x29 &  x32 &  x35 &  x44 &  x47 &  x50 &  x62 &  x65 &  x71 &  x77 &  x83 &  x86 &  x92 &  x95 &  x98 &  x104 &  x107 &  x110 &  x116 &  x119 &  x122 &  x125 &  x131 &  x140 &  x143 &  x146 &  x149 &  x161 &  x164 &  x173 &  x176 &  x182 &  x191 &  x203 &  x209 &  x212 &  x215 &  x224 &  x227 &  x230 &  x233 &  x254 &  x269 &  x275 &  x278 &  x281 &  x284 &  x293 &  x296 &  x299 &  x320 &  x323 &  x329 &  x332 &  x335 &  x341 &  x350 &  x356 &  x359 &  x365 &  x374 &  x383 &  x389 &  x398 &  x404 &  x410 &  x413 &  x419 &  x431 &  x440 &  x443 &  x449 &  x452 &  x461 &  x464 &  x470 &  x476 &  x482 &  x485 &  x497 &  x503 &  x512 &  x515 &  x521 &  x527 &  x530 &  x533 &  x536 &  x542 &  x545 &  x548 &  x554 &  x563 &  x566 &  x569 &  x572 &  x575 &  x584 &  x587 &  x590 &  x593 &  x599 &  x602 &  x605 &  x611 &  x617 &  x620 &  x623 &  x632 &  x635 &  x638 &  x641 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x680 &  x689 &  x692 &  x701 &  x704 &  x713 &  x716 &  x722 &  x725 &  x728 &  x743 &  x746 &  x758 &  x764 &  x773 &  x791 &  x800 &  x806 &  x809 &  x818 &  x830 &  x845 &  x848 &  x857 &  x860 &  x863 &  x866 &  x878 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x917 &  x920 &  x926 &  x929 &  x935 &  x938 &  x941 &  x944 &  x947 &  x956 &  x965 &  x971 &  x980 &  x986 &  x989 &  x992 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1034 &  x1046 &  x1052 &  x1055 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1097 &  x1100 &  x1109 &  x1112 &  x1118 &  x1130 & ~x753 & ~x759 & ~x792 & ~x798 & ~x831 & ~x909 & ~x948 & ~x949 & ~x954 & ~x988 & ~x1026 & ~x1065 & ~x1066;
assign c0177 =  x17 &  x35 &  x61 &  x83 &  x248 &  x307 &  x334 &  x346 &  x451 &  x490 &  x542 &  x547 &  x560 &  x662 &  x707 &  x710 &  x829 &  x931 &  x971 &  x1025 &  x1078;
assign c0179 =  x2 &  x26 &  x95 &  x215 &  x236 &  x305 &  x325 &  x338 &  x404 &  x410 &  x500 &  x506 &  x535 &  x584 &  x590 &  x593 &  x601 &  x604 &  x605 &  x607 &  x617 &  x635 &  x643 &  x668 &  x688 &  x721 &  x749 &  x764 &  x767 &  x776 &  x779 &  x803 &  x830 &  x887 &  x935 &  x938 &  x940 &  x971 &  x995 &  x998 &  x1067;
assign c0181 =  x5 &  x17 &  x41 &  x44 &  x53 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x119 &  x140 &  x143 &  x155 &  x161 &  x167 &  x173 &  x179 &  x182 &  x209 &  x221 &  x230 &  x242 &  x245 &  x262 &  x266 &  x281 &  x290 &  x299 &  x302 &  x305 &  x311 &  x343 &  x353 &  x365 &  x376 &  x377 &  x398 &  x425 &  x428 &  x437 &  x449 &  x452 &  x461 &  x467 &  x470 &  x479 &  x482 &  x485 &  x491 &  x536 &  x551 &  x560 &  x584 &  x590 &  x599 &  x602 &  x611 &  x620 &  x626 &  x629 &  x656 &  x662 &  x674 &  x683 &  x686 &  x701 &  x707 &  x713 &  x716 &  x719 &  x728 &  x734 &  x737 &  x752 &  x758 &  x761 &  x770 &  x782 &  x797 &  x800 &  x829 &  x830 &  x833 &  x842 &  x862 &  x875 &  x881 &  x884 &  x890 &  x893 &  x896 &  x899 &  x905 &  x926 &  x932 &  x941 &  x944 &  x946 &  x959 &  x968 &  x977 &  x989 &  x1004 &  x1019 &  x1025 &  x1040 &  x1046 &  x1052 &  x1061 &  x1076 &  x1079 &  x1082 &  x1094 &  x1097 &  x1100 &  x1112 &  x1118 &  x1124 &  x1127 &  x1130 & ~x195 & ~x234 & ~x390 & ~x429 & ~x468;
assign c0183 = ~x1001;
assign c0185 =  x35 &  x41 &  x152 &  x212 &  x248 &  x317 &  x374 &  x377 &  x404 &  x425 &  x557 &  x560 &  x571 &  x572 &  x593 &  x610 &  x611 &  x686 &  x713 &  x719 &  x815 &  x830 &  x869 &  x971 &  x995 &  x1076 &  x1091 &  x1100 & ~x411 & ~x423 & ~x625 & ~x711 & ~x750 & ~x828;
assign c0187 =  x20 &  x41 &  x89 &  x95 &  x128 &  x140 &  x173 &  x209 &  x224 &  x278 &  x314 &  x338 &  x371 &  x374 &  x380 &  x395 &  x425 &  x452 &  x476 &  x521 &  x539 &  x557 &  x590 &  x608 &  x617 &  x623 &  x638 &  x680 &  x695 &  x707 &  x710 &  x719 &  x743 &  x764 &  x770 &  x776 &  x791 &  x839 &  x869 &  x881 &  x890 &  x902 &  x941 &  x973 &  x980 &  x1001 &  x1028 &  x1043 &  x1070 & ~x324 & ~x363 & ~x381 & ~x408 & ~x447 & ~x465 & ~x564 & ~x603 & ~x642;
assign c0189 = ~x620;
assign c0191 =  x269 &  x296 &  x317 &  x476 &  x500 &  x568 &  x803 &  x806 &  x856 &  x895 &  x896 &  x923 &  x938 &  x971 &  x995 &  x1037 &  x1067 &  x1088 &  x1124 & ~x402 & ~x642 & ~x996;
assign c0193 =  x17 &  x65 &  x92 &  x128 &  x176 &  x212 &  x218 &  x245 &  x275 &  x371 &  x395 &  x410 &  x440 &  x449 &  x503 &  x506 &  x551 &  x572 &  x620 &  x644 &  x647 &  x662 &  x688 &  x752 &  x755 &  x788 &  x860 &  x923 &  x931 &  x932 &  x949 &  x953 &  x959 &  x965 &  x977 &  x988 &  x1013 &  x1019 &  x1058 &  x1111 &  x1117 &  x1118 & ~x627 & ~x744 & ~x783 & ~x936;
assign c0195 =  x631 & ~x304 & ~x705 & ~x936;
assign c0197 = ~x533;
assign c0199 =  x64 &  x155 &  x230 &  x277 &  x347 &  x395 &  x560 &  x626 &  x740 &  x764 &  x769 &  x938 &  x1010 &  x1070 & ~x546 & ~x627 & ~x936;
assign c0201 =  x5 &  x17 &  x74 &  x113 &  x131 &  x179 &  x182 &  x188 &  x257 &  x275 &  x287 &  x359 &  x368 &  x527 &  x539 &  x550 &  x563 &  x584 &  x605 &  x653 &  x665 &  x719 &  x791 &  x824 &  x851 &  x869 &  x956 &  x977 &  x983 &  x1004 &  x1007 &  x1013 &  x1037 &  x1076 &  x1079 &  x1106 &  x1115 &  x1121 &  x1130 & ~x195 & ~x765 & ~x804 & ~x900;
assign c0203 =  x5 &  x14 &  x32 &  x35 &  x38 &  x56 &  x64 &  x101 &  x103 &  x104 &  x110 &  x122 &  x128 &  x131 &  x140 &  x146 &  x158 &  x164 &  x176 &  x182 &  x197 &  x206 &  x209 &  x218 &  x221 &  x224 &  x227 &  x230 &  x239 &  x248 &  x259 &  x260 &  x275 &  x293 &  x305 &  x308 &  x320 &  x326 &  x329 &  x332 &  x356 &  x359 &  x362 &  x365 &  x368 &  x380 &  x389 &  x395 &  x401 &  x446 &  x464 &  x470 &  x476 &  x488 &  x491 &  x494 &  x503 &  x509 &  x515 &  x524 &  x527 &  x530 &  x560 &  x581 &  x584 &  x587 &  x593 &  x596 &  x635 &  x638 &  x653 &  x659 &  x665 &  x674 &  x695 &  x698 &  x710 &  x713 &  x716 &  x731 &  x734 &  x743 &  x746 &  x752 &  x764 &  x788 &  x803 &  x824 &  x827 &  x830 &  x833 &  x842 &  x860 &  x863 &  x881 &  x893 &  x902 &  x905 &  x917 &  x923 &  x947 &  x962 &  x968 &  x971 &  x980 &  x986 &  x989 &  x1004 &  x1016 &  x1028 &  x1031 &  x1034 &  x1040 &  x1051 &  x1067 &  x1078 &  x1085 &  x1091 &  x1094 &  x1097 &  x1115 &  x1127 & ~x186;
assign c0205 =  x239 &  x293 &  x368 &  x553 &  x773 & ~x394 & ~x414 & ~x492;
assign c0207 =  x178 &  x1126 & ~x660 & ~x915 & ~x924;
assign c0209 =  x97 &  x155 & ~x0 & ~x195 & ~x351 & ~x921 & ~x993;
assign c0211 =  x173 &  x181 &  x206 &  x212 &  x239 &  x248 &  x254 &  x302 &  x359 &  x452 &  x545 &  x644 &  x667 &  x704 &  x857 &  x869 &  x977 &  x1001 &  x1037 &  x1079 & ~x537 & ~x576 & ~x654 & ~x732 & ~x939;
assign c0213 =  x23 &  x250 &  x254 &  x256 &  x280 &  x346 &  x359 &  x536 &  x571 &  x581 &  x595 &  x758 &  x862 &  x866 &  x868 &  x893 &  x905 &  x907 &  x1061;
assign c0215 =  x5 &  x122 &  x152 &  x314 &  x350 &  x419 &  x467 &  x581 &  x623 &  x701 &  x800 &  x884 &  x928 &  x932 &  x964 &  x967 &  x1051 &  x1129 & ~x759 & ~x837 & ~x936;
assign c0217 =  x281 &  x377 &  x398 &  x643 &  x650 &  x749 &  x842 & ~x795 & ~x813 & ~x912 & ~x913 & ~x969 & ~x991 & ~x1107 & ~x1113;
assign c0219 =  x124 &  x315 & ~x627;
assign c0221 =  x44 &  x47 &  x80 &  x140 &  x152 &  x227 &  x299 &  x455 &  x472 &  x503 &  x509 &  x511 &  x629 &  x761 &  x806 &  x863 &  x908 &  x965 &  x1094 & ~x156 & ~x537 & ~x783;
assign c0223 =  x2 &  x11 &  x26 &  x32 &  x65 &  x71 &  x83 &  x89 &  x95 &  x107 &  x128 &  x146 &  x152 &  x167 &  x179 &  x227 &  x230 &  x235 &  x239 &  x248 &  x260 &  x272 &  x274 &  x275 &  x290 &  x329 &  x332 &  x335 &  x338 &  x425 &  x428 &  x440 &  x446 &  x488 &  x497 &  x500 &  x506 &  x518 &  x542 &  x545 &  x551 &  x557 &  x560 &  x569 &  x575 &  x590 &  x593 &  x635 &  x644 &  x650 &  x695 &  x704 &  x707 &  x710 &  x719 &  x740 &  x764 &  x770 &  x778 &  x817 &  x827 &  x842 &  x844 &  x856 &  x875 &  x881 &  x883 &  x884 &  x920 &  x923 &  x928 &  x929 &  x941 &  x944 &  x947 &  x959 &  x977 &  x980 &  x983 &  x989 &  x992 &  x1049 &  x1064 &  x1073 &  x1085 &  x1091 &  x1094 &  x1100 &  x1115 & ~x270 & ~x603;
assign c0225 =  x280 &  x568 &  x607 &  x895 & ~x679;
assign c0227 =  x865 &  x1083 &  x1117 & ~x126 & ~x657;
assign c0229 =  x5 &  x8 &  x14 &  x17 &  x26 &  x29 &  x32 &  x35 &  x41 &  x44 &  x50 &  x53 &  x56 &  x65 &  x68 &  x71 &  x80 &  x89 &  x92 &  x101 &  x107 &  x116 &  x119 &  x128 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x155 &  x158 &  x161 &  x167 &  x170 &  x179 &  x182 &  x185 &  x194 &  x197 &  x200 &  x203 &  x212 &  x221 &  x233 &  x236 &  x239 &  x245 &  x248 &  x251 &  x254 &  x260 &  x266 &  x269 &  x281 &  x284 &  x290 &  x296 &  x299 &  x302 &  x308 &  x314 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x377 &  x383 &  x386 &  x392 &  x395 &  x398 &  x404 &  x407 &  x410 &  x413 &  x422 &  x425 &  x428 &  x434 &  x437 &  x446 &  x449 &  x458 &  x461 &  x467 &  x472 &  x473 &  x476 &  x482 &  x488 &  x491 &  x494 &  x503 &  x515 &  x521 &  x524 &  x533 &  x542 &  x548 &  x560 &  x563 &  x575 &  x578 &  x581 &  x587 &  x590 &  x593 &  x596 &  x602 &  x605 &  x611 &  x626 &  x632 &  x635 &  x638 &  x641 &  x647 &  x650 &  x656 &  x659 &  x661 &  x662 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x692 &  x698 &  x707 &  x710 &  x713 &  x716 &  x719 &  x725 &  x734 &  x737 &  x740 &  x743 &  x758 &  x761 &  x770 &  x773 &  x779 &  x782 &  x788 &  x791 &  x800 &  x803 &  x806 &  x815 &  x818 &  x821 &  x824 &  x833 &  x839 &  x842 &  x848 &  x854 &  x860 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x890 &  x893 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x935 &  x944 &  x953 &  x959 &  x965 &  x971 &  x977 &  x980 &  x983 &  x995 &  x998 &  x1001 &  x1010 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1079 &  x1088 &  x1094 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x225 & ~x342 & ~x381 & ~x405 & ~x444 & ~x483 & ~x522 & ~x603 & ~x642;
assign c0231 =  x392 &  x659 &  x674 &  x947 & ~x9 & ~x669 & ~x792 & ~x939 & ~x1017;
assign c0233 =  x250 &  x340 &  x380 &  x563 &  x568 &  x815 & ~x438 & ~x757;
assign c0235 =  x2 &  x23 &  x38 &  x47 &  x50 &  x56 &  x59 &  x68 &  x71 &  x80 &  x92 &  x101 &  x122 &  x125 &  x128 &  x131 &  x143 &  x161 &  x170 &  x173 &  x215 &  x224 &  x257 &  x302 &  x317 &  x323 &  x332 &  x338 &  x350 &  x359 &  x365 &  x377 &  x380 &  x383 &  x398 &  x401 &  x428 &  x434 &  x437 &  x443 &  x449 &  x458 &  x461 &  x470 &  x482 &  x491 &  x506 &  x512 &  x524 &  x578 &  x584 &  x590 &  x593 &  x614 &  x620 &  x623 &  x629 &  x638 &  x641 &  x659 &  x662 &  x674 &  x680 &  x701 &  x707 &  x710 &  x743 &  x752 &  x785 &  x797 &  x809 &  x812 &  x815 &  x821 &  x833 &  x836 &  x839 &  x842 &  x869 &  x875 &  x896 &  x902 &  x905 &  x923 &  x944 &  x959 &  x980 &  x986 &  x992 &  x1010 &  x1016 &  x1022 &  x1028 &  x1031 &  x1037 &  x1040 &  x1061 &  x1094 &  x1103 &  x1109 &  x1118 &  x1124 &  x1127 &  x1130 & ~x465 & ~x642 & ~x783 & ~x822 & ~x861 & ~x862 & ~x939 & ~x978;
assign c0237 =  x35 &  x41 &  x44 &  x50 &  x62 &  x68 &  x83 &  x98 &  x104 &  x121 &  x122 &  x128 &  x146 &  x152 &  x155 &  x158 &  x182 &  x212 &  x227 &  x230 &  x242 &  x257 &  x278 &  x281 &  x287 &  x290 &  x293 &  x299 &  x308 &  x353 &  x359 &  x374 &  x389 &  x404 &  x416 &  x422 &  x425 &  x467 &  x476 &  x494 &  x500 &  x518 &  x542 &  x578 &  x593 &  x596 &  x599 &  x614 &  x617 &  x620 &  x626 &  x629 &  x635 &  x659 &  x662 &  x671 &  x677 &  x689 &  x692 &  x698 &  x701 &  x704 &  x719 &  x725 &  x731 &  x761 &  x764 &  x772 &  x776 &  x785 &  x791 &  x806 &  x818 &  x827 &  x848 &  x869 &  x887 &  x893 &  x896 &  x899 &  x905 &  x929 &  x938 &  x941 &  x965 &  x968 &  x977 &  x992 &  x995 &  x1010 &  x1016 &  x1019 &  x1025 &  x1028 &  x1034 &  x1061 &  x1073 &  x1082 &  x1085 &  x1091 & ~x609 & ~x681 & ~x822;
assign c0239 =  x11 &  x53 &  x65 &  x86 &  x95 &  x119 &  x173 &  x176 &  x305 &  x320 &  x386 &  x404 &  x409 &  x464 &  x473 &  x485 &  x500 &  x503 &  x545 &  x548 &  x578 &  x614 &  x635 &  x725 &  x743 &  x746 &  x764 &  x851 &  x944 &  x962 &  x986 &  x1016 &  x1034 &  x1052 &  x1058 &  x1064 &  x1067 &  x1076 &  x1079 & ~x156 & ~x954 & ~x1038 & ~x1074 & ~x1113;
assign c0241 =  x620 &  x1004 & ~x195 & ~x285 & ~x483 & ~x861;
assign c0243 =  x20 &  x22 &  x35 &  x50 &  x74 &  x101 &  x164 &  x200 &  x218 &  x289 &  x292 &  x302 &  x452 &  x476 &  x527 &  x587 &  x602 &  x626 &  x647 &  x656 &  x683 &  x734 &  x746 &  x815 &  x823 &  x829 &  x884 &  x985 &  x1034 & ~x468;
assign c0245 =  x98 &  x110 &  x137 &  x143 &  x242 &  x482 &  x509 &  x700 &  x758 &  x881 &  x934 &  x1052 &  x1064 &  x1085 &  x1094 & ~x420 & ~x525 & ~x783 & ~x936;
assign c0247 =  x152 &  x280 &  x1043 &  x1064 & ~x442 & ~x597;
assign c0249 =  x33 &  x196 &  x356 &  x526 &  x620 &  x724 &  x1042 & ~x714;
assign c0251 = ~x940;
assign c0253 =  x89 &  x215 &  x250 &  x301 &  x307 &  x346 &  x358 &  x422 &  x526 &  x590 &  x593 &  x698 &  x758 &  x848 &  x946 &  x1081 &  x1085;
assign c0255 =  x2 &  x5 &  x11 &  x20 &  x29 &  x35 &  x38 &  x47 &  x50 &  x53 &  x65 &  x68 &  x71 &  x86 &  x89 &  x100 &  x110 &  x116 &  x134 &  x139 &  x140 &  x145 &  x149 &  x173 &  x178 &  x185 &  x188 &  x200 &  x206 &  x212 &  x215 &  x217 &  x224 &  x230 &  x242 &  x245 &  x254 &  x272 &  x281 &  x287 &  x296 &  x302 &  x331 &  x335 &  x341 &  x347 &  x383 &  x398 &  x413 &  x416 &  x419 &  x434 &  x440 &  x452 &  x458 &  x464 &  x470 &  x476 &  x479 &  x482 &  x488 &  x503 &  x524 &  x529 &  x530 &  x542 &  x548 &  x554 &  x557 &  x566 &  x568 &  x569 &  x578 &  x584 &  x587 &  x593 &  x606 &  x607 &  x626 &  x635 &  x646 &  x647 &  x653 &  x659 &  x662 &  x668 &  x674 &  x680 &  x689 &  x707 &  x710 &  x713 &  x724 &  x725 &  x743 &  x746 &  x749 &  x761 &  x770 &  x776 &  x779 &  x791 &  x803 &  x806 &  x818 &  x821 &  x839 &  x848 &  x854 &  x869 &  x884 &  x896 &  x920 &  x959 &  x962 &  x986 &  x998 &  x1001 &  x1010 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1036 &  x1049 &  x1070 &  x1082 &  x1088 &  x1100 &  x1118 &  x1121 &  x1127 &  x1130;
assign c0257 =  x20 &  x29 &  x47 &  x50 &  x59 &  x71 &  x86 &  x101 &  x110 &  x119 &  x125 &  x134 &  x155 &  x158 &  x173 &  x203 &  x212 &  x218 &  x242 &  x257 &  x260 &  x263 &  x308 &  x311 &  x332 &  x335 &  x338 &  x380 &  x392 &  x403 &  x404 &  x410 &  x416 &  x437 &  x446 &  x452 &  x467 &  x473 &  x494 &  x497 &  x503 &  x509 &  x539 &  x542 &  x569 &  x587 &  x629 &  x644 &  x650 &  x667 &  x668 &  x695 &  x728 &  x731 &  x734 &  x737 &  x773 &  x812 &  x824 &  x863 &  x911 &  x923 &  x935 &  x947 &  x953 &  x959 &  x965 &  x968 &  x977 &  x983 &  x992 &  x1001 &  x1004 &  x1007 &  x1010 &  x1049 &  x1058 &  x1064 &  x1067 &  x1073 &  x1106 &  x1112 &  x1130 & ~x273 & ~x732 & ~x771 & ~x810 & ~x960 & ~x993;
assign c0259 = ~x251;
assign c0261 =  x77 &  x139 &  x220 &  x256 &  x331 &  x490 &  x529 &  x634 &  x970 &  x1078;
assign c0263 =  x58 & ~x492 & ~x745;
assign c0265 = ~x992;
assign c0267 =  x113 &  x149 &  x260 &  x263 &  x404 &  x443 &  x449 &  x452 &  x458 &  x560 &  x575 &  x620 &  x692 &  x716 &  x758 &  x797 &  x827 &  x875 &  x931 &  x932 &  x944 &  x1049 &  x1100 &  x1118 &  x1124 & ~x312 & ~x651 & ~x1056;
assign c0269 =  x185 &  x251 &  x254 &  x275 &  x305 &  x326 &  x343 &  x353 &  x392 &  x407 &  x521 &  x659 &  x686 &  x704 &  x767 &  x884 &  x896 &  x956 &  x965 & ~x354 & ~x390 & ~x429 & ~x468 & ~x507 & ~x633 & ~x660 & ~x966;
assign c0271 =  x171 &  x178 &  x1033 & ~x831 & ~x939;
assign c0273 =  x44 &  x70 &  x122 &  x131 &  x149 &  x173 &  x187 &  x239 &  x331 &  x401 &  x425 &  x446 &  x458 &  x485 &  x491 &  x521 &  x526 &  x548 &  x788 &  x829 &  x863 &  x989 &  x1055;
assign c0275 = ~x564 & ~x636 & ~x976 & ~x1074;
assign c0277 =  x269 &  x293 &  x437 &  x452 &  x677 &  x1052 & ~x369 & ~x588 & ~x936 & ~x976;
assign c0279 = ~x233;
assign c0281 =  x5 &  x14 &  x164 &  x170 &  x236 &  x248 &  x254 &  x260 &  x275 &  x278 &  x311 &  x344 &  x371 &  x434 &  x446 &  x494 &  x500 &  x503 &  x512 &  x518 &  x533 &  x539 &  x593 &  x608 &  x617 &  x638 &  x641 &  x644 &  x695 &  x701 &  x719 &  x725 &  x746 &  x787 &  x800 &  x809 &  x815 &  x817 &  x854 &  x908 &  x989 &  x1019 &  x1028 &  x1031 &  x1088 &  x1091 &  x1100 &  x1105 &  x1124 &  x1130 & ~x153 & ~x231 & ~x564 & ~x603 & ~x705;
assign c0283 =  x5 &  x11 &  x23 &  x26 &  x29 &  x32 &  x35 &  x41 &  x44 &  x47 &  x56 &  x62 &  x68 &  x74 &  x77 &  x80 &  x83 &  x95 &  x98 &  x101 &  x116 &  x122 &  x125 &  x128 &  x131 &  x134 &  x140 &  x143 &  x152 &  x158 &  x161 &  x164 &  x176 &  x182 &  x188 &  x191 &  x221 &  x230 &  x251 &  x254 &  x257 &  x263 &  x275 &  x290 &  x299 &  x311 &  x317 &  x323 &  x326 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x359 &  x362 &  x374 &  x377 &  x380 &  x383 &  x389 &  x392 &  x404 &  x407 &  x413 &  x422 &  x425 &  x428 &  x434 &  x440 &  x452 &  x458 &  x473 &  x476 &  x482 &  x485 &  x491 &  x497 &  x506 &  x509 &  x512 &  x524 &  x539 &  x545 &  x566 &  x569 &  x572 &  x578 &  x581 &  x590 &  x602 &  x617 &  x623 &  x629 &  x644 &  x647 &  x650 &  x656 &  x661 &  x662 &  x665 &  x674 &  x683 &  x692 &  x704 &  x728 &  x746 &  x755 &  x764 &  x766 &  x767 &  x773 &  x776 &  x785 &  x794 &  x815 &  x827 &  x830 &  x836 &  x839 &  x848 &  x851 &  x856 &  x893 &  x895 &  x896 &  x905 &  x914 &  x920 &  x923 &  x926 &  x938 &  x944 &  x950 &  x959 &  x971 &  x973 &  x974 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1007 &  x1016 &  x1019 &  x1025 &  x1028 &  x1034 &  x1046 &  x1052 &  x1055 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1094 &  x1097 &  x1100 &  x1112 &  x1118 &  x1121 &  x1127 & ~x207 & ~x246 & ~x285 & ~x525;
assign c0285 =  x41 &  x101 &  x119 &  x143 &  x161 &  x173 &  x179 &  x188 &  x200 &  x227 &  x238 &  x275 &  x365 &  x380 &  x404 &  x482 &  x524 &  x548 &  x554 &  x590 &  x596 &  x665 &  x673 &  x674 &  x698 &  x712 &  x716 &  x818 &  x857 &  x887 &  x923 &  x965 &  x1097 &  x1100 & ~x234 & ~x312 & ~x780;
assign c0287 =  x11 &  x177 &  x211 &  x256 &  x529 &  x607 &  x892;
assign c0289 =  x61 &  x139 &  x142 &  x172 &  x173 &  x182 &  x200 &  x203 &  x211 &  x254 &  x275 &  x284 &  x290 &  x296 &  x331 &  x334 &  x335 &  x389 &  x407 &  x443 &  x529 &  x638 &  x662 &  x668 &  x674 &  x727 &  x734 &  x761 &  x791 &  x860 &  x863 &  x902 &  x917 &  x932 &  x965 &  x1010 &  x1040 &  x1064 &  x1118;
assign c0291 =  x286 &  x643 & ~x430 & ~x660 & ~x885;
assign c0293 =  x12 &  x311 &  x350 &  x353 &  x397 &  x446 &  x476 &  x536 &  x574 &  x704 &  x722 &  x914 &  x950 &  x980 &  x1106;
assign c0295 =  x121 &  x352 &  x440 &  x668 &  x736 &  x905 & ~x447 & ~x667;
assign c0297 = ~x685 & ~x729 & ~x898;
assign c0299 =  x29 &  x56 &  x59 &  x71 &  x101 &  x104 &  x131 &  x167 &  x197 &  x200 &  x224 &  x233 &  x245 &  x248 &  x260 &  x284 &  x287 &  x317 &  x329 &  x335 &  x338 &  x353 &  x359 &  x401 &  x404 &  x410 &  x413 &  x425 &  x434 &  x440 &  x461 &  x470 &  x473 &  x500 &  x503 &  x515 &  x542 &  x548 &  x557 &  x560 &  x589 &  x599 &  x608 &  x626 &  x628 &  x671 &  x683 &  x713 &  x728 &  x761 &  x797 &  x812 &  x839 &  x845 &  x875 &  x899 &  x908 &  x965 &  x977 &  x1013 &  x1016 &  x1031 &  x1043 &  x1067 &  x1082 &  x1097 &  x1100 & ~x312 & ~x909 & ~x939;
assign c10 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x227 &  x233 &  x239 &  x242 &  x245 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x659 &  x662 &  x664 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x701 &  x703 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x742 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x776 &  x779 &  x781 &  x782 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x820 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x859 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x893 &  x896 &  x898 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x940 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x976 &  x977 &  x979 &  x980 &  x983 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1018 &  x1019 &  x1021 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1057 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x312 & ~x351 & ~x390 & ~x429 & ~x477 & ~x591 & ~x630;
assign c12 =  x14 &  x17 &  x20 &  x23 &  x29 &  x32 &  x35 &  x38 &  x41 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x89 &  x101 &  x107 &  x110 &  x116 &  x119 &  x122 &  x131 &  x134 &  x137 &  x143 &  x146 &  x152 &  x155 &  x161 &  x164 &  x173 &  x176 &  x182 &  x191 &  x200 &  x203 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x269 &  x272 &  x278 &  x281 &  x284 &  x290 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x317 &  x326 &  x332 &  x335 &  x341 &  x347 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x395 &  x407 &  x410 &  x413 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x446 &  x452 &  x455 &  x461 &  x467 &  x476 &  x479 &  x482 &  x485 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x512 &  x515 &  x521 &  x524 &  x527 &  x533 &  x536 &  x542 &  x545 &  x548 &  x557 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x587 &  x593 &  x596 &  x599 &  x605 &  x608 &  x611 &  x617 &  x620 &  x626 &  x629 &  x635 &  x638 &  x650 &  x653 &  x656 &  x665 &  x668 &  x671 &  x674 &  x680 &  x692 &  x698 &  x701 &  x707 &  x710 &  x713 &  x716 &  x722 &  x725 &  x737 &  x743 &  x746 &  x749 &  x752 &  x755 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x809 &  x812 &  x815 &  x821 &  x823 &  x824 &  x833 &  x836 &  x839 &  x851 &  x857 &  x866 &  x872 &  x875 &  x878 &  x884 &  x893 &  x896 &  x899 &  x905 &  x908 &  x911 &  x914 &  x917 &  x926 &  x929 &  x932 &  x938 &  x941 &  x944 &  x950 &  x953 &  x956 &  x959 &  x962 &  x968 &  x971 &  x980 &  x982 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1060 &  x1061 &  x1079 &  x1085 &  x1091 &  x1094 &  x1097 &  x1099 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 &  x1130 & ~x48 & ~x87 & ~x126 & ~x228 & ~x384 & ~x919 & ~x951 & ~x957 & ~x990 & ~x996 & ~x1029 & ~x1074;
assign c14 =  x2 &  x11 &  x23 &  x35 &  x41 &  x47 &  x50 &  x53 &  x89 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x119 &  x122 &  x125 &  x140 &  x143 &  x149 &  x158 &  x173 &  x182 &  x185 &  x194 &  x203 &  x215 &  x224 &  x227 &  x233 &  x236 &  x245 &  x248 &  x251 &  x257 &  x260 &  x284 &  x290 &  x299 &  x305 &  x314 &  x316 &  x317 &  x320 &  x326 &  x332 &  x341 &  x344 &  x353 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x377 &  x386 &  x389 &  x392 &  x404 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x446 &  x452 &  x458 &  x461 &  x464 &  x473 &  x476 &  x488 &  x500 &  x503 &  x509 &  x515 &  x521 &  x524 &  x527 &  x533 &  x539 &  x545 &  x548 &  x551 &  x557 &  x560 &  x566 &  x578 &  x584 &  x595 &  x599 &  x605 &  x608 &  x614 &  x620 &  x623 &  x626 &  x634 &  x635 &  x638 &  x644 &  x650 &  x656 &  x659 &  x662 &  x668 &  x669 &  x671 &  x677 &  x680 &  x689 &  x695 &  x704 &  x707 &  x709 &  x710 &  x713 &  x716 &  x722 &  x725 &  x737 &  x748 &  x749 &  x752 &  x755 &  x761 &  x764 &  x767 &  x773 &  x776 &  x779 &  x788 &  x791 &  x794 &  x797 &  x815 &  x818 &  x830 &  x839 &  x842 &  x851 &  x857 &  x860 &  x869 &  x872 &  x875 &  x884 &  x887 &  x890 &  x896 &  x899 &  x905 &  x908 &  x911 &  x917 &  x920 &  x926 &  x929 &  x932 &  x938 &  x941 &  x947 &  x965 &  x968 &  x974 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1010 &  x1013 &  x1019 &  x1028 &  x1033 &  x1037 &  x1040 &  x1049 &  x1052 &  x1058 &  x1067 &  x1070 &  x1073 &  x1085 &  x1088 &  x1097 &  x1100 &  x1103 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x486 & ~x600 & ~x624 & ~x663 & ~x702 & ~x741 & ~x780 & ~x819 & ~x858 & ~x900 & ~x936 & ~x939 & ~x975;
assign c16 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x29 &  x35 &  x38 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x125 &  x128 &  x137 &  x140 &  x143 &  x146 &  x152 &  x158 &  x161 &  x164 &  x167 &  x179 &  x188 &  x191 &  x194 &  x197 &  x203 &  x206 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x287 &  x290 &  x293 &  x296 &  x308 &  x311 &  x317 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x353 &  x356 &  x359 &  x371 &  x377 &  x380 &  x383 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x418 &  x419 &  x422 &  x425 &  x434 &  x437 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x460 &  x461 &  x464 &  x466 &  x467 &  x470 &  x476 &  x479 &  x485 &  x488 &  x497 &  x499 &  x503 &  x506 &  x512 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x545 &  x548 &  x557 &  x559 &  x560 &  x563 &  x565 &  x569 &  x572 &  x584 &  x587 &  x590 &  x593 &  x599 &  x602 &  x604 &  x605 &  x608 &  x611 &  x614 &  x620 &  x626 &  x629 &  x635 &  x640 &  x644 &  x647 &  x653 &  x656 &  x662 &  x668 &  x671 &  x674 &  x679 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x701 &  x713 &  x716 &  x718 &  x719 &  x722 &  x725 &  x731 &  x737 &  x743 &  x746 &  x749 &  x755 &  x758 &  x764 &  x767 &  x770 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x797 &  x800 &  x803 &  x809 &  x812 &  x821 &  x827 &  x830 &  x833 &  x839 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x875 &  x878 &  x881 &  x884 &  x887 &  x893 &  x896 &  x897 &  x898 &  x899 &  x902 &  x905 &  x908 &  x920 &  x923 &  x926 &  x935 &  x937 &  x941 &  x944 &  x947 &  x956 &  x959 &  x965 &  x968 &  x971 &  x977 &  x983 &  x986 &  x989 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1015 &  x1019 &  x1022 &  x1031 &  x1034 &  x1037 &  x1043 &  x1049 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1093 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 & ~x315 & ~x354 & ~x393 & ~x432 & ~x471 & ~x510 & ~x549 & ~x588 & ~x627 & ~x633;
assign c18 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x269 &  x272 &  x275 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x314 &  x317 &  x320 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x376 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x414 &  x415 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x454 &  x455 &  x458 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x493 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x526 &  x527 &  x530 &  x532 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x571 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x610 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x649 &  x650 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x688 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x727 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x766 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x965 &  x968 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x390 & ~x657 & ~x762 & ~x801 & ~x840;
assign c110 =  x5 &  x8 &  x11 &  x14 &  x20 &  x23 &  x32 &  x35 &  x38 &  x41 &  x50 &  x53 &  x62 &  x68 &  x74 &  x80 &  x82 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x116 &  x119 &  x122 &  x125 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x164 &  x167 &  x173 &  x182 &  x185 &  x191 &  x194 &  x197 &  x203 &  x206 &  x215 &  x218 &  x221 &  x230 &  x233 &  x236 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x277 &  x278 &  x281 &  x287 &  x293 &  x296 &  x299 &  x302 &  x317 &  x320 &  x326 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x355 &  x356 &  x359 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x386 &  x392 &  x395 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x436 &  x437 &  x440 &  x443 &  x446 &  x452 &  x455 &  x467 &  x475 &  x479 &  x491 &  x494 &  x500 &  x503 &  x512 &  x514 &  x515 &  x518 &  x521 &  x524 &  x527 &  x539 &  x545 &  x551 &  x553 &  x554 &  x557 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x592 &  x593 &  x596 &  x605 &  x608 &  x611 &  x614 &  x616 &  x620 &  x623 &  x626 &  x629 &  x635 &  x638 &  x641 &  x644 &  x653 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x710 &  x715 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x743 &  x746 &  x749 &  x752 &  x764 &  x766 &  x772 &  x776 &  x779 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x805 &  x806 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x854 &  x871 &  x872 &  x875 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x908 &  x910 &  x911 &  x914 &  x929 &  x932 &  x935 &  x938 &  x941 &  x949 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x980 &  x983 &  x986 &  x989 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1028 &  x1034 &  x1046 &  x1049 &  x1058 &  x1061 &  x1064 &  x1076 &  x1079 &  x1082 &  x1085 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 & ~x99 & ~x444 & ~x705;
assign c112 =  x1 &  x5 &  x11 &  x14 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x50 &  x56 &  x62 &  x65 &  x68 &  x71 &  x77 &  x80 &  x86 &  x92 &  x95 &  x98 &  x101 &  x107 &  x110 &  x113 &  x119 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x161 &  x164 &  x170 &  x176 &  x182 &  x185 &  x191 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x227 &  x236 &  x239 &  x245 &  x248 &  x251 &  x254 &  x260 &  x266 &  x269 &  x277 &  x284 &  x299 &  x302 &  x308 &  x311 &  x313 &  x314 &  x316 &  x317 &  x320 &  x326 &  x329 &  x332 &  x335 &  x338 &  x347 &  x350 &  x353 &  x355 &  x356 &  x359 &  x362 &  x368 &  x377 &  x380 &  x383 &  x389 &  x392 &  x394 &  x398 &  x410 &  x416 &  x419 &  x425 &  x428 &  x434 &  x440 &  x446 &  x449 &  x455 &  x464 &  x470 &  x472 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x497 &  x500 &  x509 &  x515 &  x518 &  x524 &  x530 &  x533 &  x536 &  x539 &  x545 &  x548 &  x551 &  x557 &  x560 &  x566 &  x569 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x596 &  x605 &  x611 &  x614 &  x620 &  x623 &  x629 &  x632 &  x635 &  x641 &  x644 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x680 &  x688 &  x689 &  x692 &  x698 &  x701 &  x704 &  x710 &  x713 &  x719 &  x725 &  x727 &  x728 &  x731 &  x734 &  x739 &  x746 &  x755 &  x761 &  x764 &  x766 &  x767 &  x776 &  x778 &  x779 &  x782 &  x788 &  x791 &  x794 &  x797 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x842 &  x845 &  x848 &  x851 &  x857 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x883 &  x884 &  x887 &  x890 &  x893 &  x896 &  x902 &  x905 &  x911 &  x917 &  x923 &  x929 &  x935 &  x938 &  x941 &  x944 &  x947 &  x953 &  x959 &  x961 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x998 &  x1001 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1040 &  x1043 &  x1045 &  x1049 &  x1051 &  x1052 &  x1055 &  x1058 &  x1061 &  x1067 &  x1070 &  x1073 &  x1076 &  x1078 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1112 &  x1121 &  x1124 &  x1127 & ~x6 & ~x45 & ~x123 & ~x741 & ~x780 & ~x819 & ~x858;
assign c114 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x91 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x119 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x458 &  x461 &  x464 &  x467 &  x470 &  x472 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x511 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x542 &  x545 &  x548 &  x550 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x623 &  x626 &  x628 &  x629 &  x632 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x667 &  x668 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x758 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x842 &  x845 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x962 &  x965 &  x968 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x333 & ~x372 & ~x450 & ~x459 & ~x489 & ~x498 & ~x528 & ~x723 & ~x918 & ~x957 & ~x990 & ~x996 & ~x1035;
assign c116 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x185 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x239 &  x242 &  x245 &  x248 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x337 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x395 &  x404 &  x407 &  x410 &  x413 &  x415 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x683 &  x686 &  x689 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x764 &  x770 &  x773 &  x776 &  x779 &  x782 &  x784 &  x785 &  x788 &  x794 &  x797 &  x800 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x943 &  x944 &  x947 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x977 &  x980 &  x982 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1021 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1060 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x117 & ~x156 & ~x195 & ~x234 & ~x312 & ~x795 & ~x873 & ~x912 & ~x951 & ~x996 & ~x999 & ~x1014 & ~x1053 & ~x1092;
assign c118 =  x2 &  x11 &  x17 &  x26 &  x41 &  x44 &  x47 &  x50 &  x53 &  x62 &  x83 &  x86 &  x92 &  x98 &  x101 &  x104 &  x113 &  x116 &  x122 &  x125 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x152 &  x155 &  x161 &  x173 &  x176 &  x182 &  x191 &  x194 &  x200 &  x203 &  x212 &  x218 &  x224 &  x227 &  x233 &  x236 &  x245 &  x251 &  x254 &  x257 &  x259 &  x260 &  x263 &  x266 &  x272 &  x275 &  x278 &  x284 &  x290 &  x292 &  x293 &  x296 &  x299 &  x302 &  x304 &  x311 &  x317 &  x323 &  x335 &  x337 &  x344 &  x353 &  x356 &  x359 &  x368 &  x371 &  x374 &  x383 &  x392 &  x398 &  x407 &  x413 &  x419 &  x422 &  x428 &  x431 &  x434 &  x437 &  x440 &  x446 &  x449 &  x458 &  x464 &  x470 &  x473 &  x476 &  x485 &  x491 &  x497 &  x500 &  x509 &  x512 &  x518 &  x524 &  x527 &  x530 &  x545 &  x554 &  x560 &  x563 &  x566 &  x581 &  x584 &  x593 &  x596 &  x611 &  x623 &  x626 &  x632 &  x638 &  x641 &  x644 &  x647 &  x656 &  x668 &  x677 &  x680 &  x689 &  x695 &  x701 &  x707 &  x716 &  x719 &  x725 &  x728 &  x734 &  x737 &  x743 &  x746 &  x749 &  x755 &  x761 &  x770 &  x773 &  x784 &  x788 &  x794 &  x797 &  x800 &  x803 &  x809 &  x812 &  x815 &  x821 &  x823 &  x829 &  x833 &  x839 &  x842 &  x845 &  x851 &  x862 &  x863 &  x872 &  x875 &  x884 &  x887 &  x899 &  x901 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x935 &  x938 &  x944 &  x947 &  x953 &  x959 &  x974 &  x977 &  x979 &  x980 &  x985 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1016 &  x1018 &  x1019 &  x1028 &  x1034 &  x1040 &  x1046 &  x1049 &  x1055 &  x1057 &  x1063 &  x1064 &  x1067 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x195 & ~x234 & ~x273 & ~x276 & ~x354 & ~x393 & ~x432 & ~x618;
assign c120 =  x14 &  x17 &  x20 &  x38 &  x41 &  x62 &  x68 &  x71 &  x74 &  x86 &  x89 &  x107 &  x116 &  x119 &  x122 &  x125 &  x155 &  x164 &  x167 &  x173 &  x176 &  x185 &  x188 &  x206 &  x209 &  x217 &  x218 &  x224 &  x227 &  x230 &  x245 &  x263 &  x266 &  x284 &  x290 &  x296 &  x311 &  x329 &  x331 &  x334 &  x335 &  x350 &  x356 &  x359 &  x368 &  x371 &  x376 &  x380 &  x383 &  x389 &  x395 &  x398 &  x415 &  x421 &  x427 &  x428 &  x440 &  x467 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x494 &  x497 &  x503 &  x530 &  x536 &  x539 &  x548 &  x557 &  x560 &  x578 &  x584 &  x593 &  x596 &  x598 &  x605 &  x608 &  x611 &  x626 &  x629 &  x641 &  x665 &  x671 &  x680 &  x695 &  x701 &  x707 &  x710 &  x716 &  x725 &  x731 &  x740 &  x749 &  x752 &  x758 &  x767 &  x779 &  x788 &  x806 &  x809 &  x815 &  x821 &  x827 &  x830 &  x845 &  x848 &  x857 &  x862 &  x863 &  x869 &  x872 &  x881 &  x893 &  x896 &  x899 &  x901 &  x908 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x941 &  x947 &  x953 &  x956 &  x962 &  x965 &  x968 &  x976 &  x979 &  x986 &  x989 &  x995 &  x998 &  x1004 &  x1010 &  x1016 &  x1018 &  x1019 &  x1022 &  x1025 &  x1057 &  x1063 &  x1073 &  x1079 &  x1088 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1127 & ~x393 & ~x660;
assign c122 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x263 &  x266 &  x272 &  x275 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x422 &  x425 &  x431 &  x437 &  x440 &  x443 &  x446 &  x449 &  x455 &  x458 &  x461 &  x464 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x584 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x623 &  x626 &  x629 &  x632 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x704 &  x707 &  x710 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x800 &  x803 &  x806 &  x809 &  x812 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x866 &  x869 &  x872 &  x875 &  x881 &  x884 &  x890 &  x893 &  x896 &  x899 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x938 &  x940 &  x941 &  x943 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x982 &  x983 &  x986 &  x989 &  x992 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1021 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x399 & ~x438 & ~x558 & ~x834 & ~x873 & ~x874 & ~x912 & ~x913 & ~x951;
assign c124 =  x5 &  x8 &  x11 &  x14 &  x17 &  x22 &  x26 &  x29 &  x32 &  x35 &  x38 &  x44 &  x50 &  x53 &  x56 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x89 &  x92 &  x95 &  x98 &  x100 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x239 &  x242 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x287 &  x289 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x323 &  x326 &  x328 &  x332 &  x335 &  x341 &  x344 &  x347 &  x350 &  x356 &  x359 &  x362 &  x365 &  x366 &  x367 &  x368 &  x371 &  x377 &  x380 &  x383 &  x392 &  x401 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x437 &  x443 &  x445 &  x446 &  x452 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x479 &  x482 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x560 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x593 &  x599 &  x605 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x641 &  x644 &  x653 &  x662 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x701 &  x704 &  x707 &  x710 &  x716 &  x719 &  x722 &  x728 &  x731 &  x734 &  x737 &  x740 &  x745 &  x746 &  x752 &  x755 &  x758 &  x761 &  x764 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x872 &  x878 &  x884 &  x887 &  x890 &  x893 &  x896 &  x902 &  x911 &  x917 &  x920 &  x923 &  x926 &  x935 &  x953 &  x956 &  x959 &  x962 &  x965 &  x971 &  x974 &  x980 &  x983 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1034 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1115 &  x1121 &  x1127 & ~x738 & ~x777 & ~x870 & ~x909 & ~x948;
assign c126 =  x2 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x152 &  x155 &  x158 &  x161 &  x164 &  x170 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x226 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x263 &  x265 &  x266 &  x269 &  x272 &  x275 &  x281 &  x284 &  x286 &  x287 &  x290 &  x292 &  x293 &  x296 &  x299 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x331 &  x332 &  x335 &  x338 &  x341 &  x343 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x370 &  x371 &  x374 &  x376 &  x380 &  x382 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x409 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x443 &  x446 &  x448 &  x449 &  x452 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x713 &  x716 &  x719 &  x725 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x788 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x815 &  x818 &  x823 &  x824 &  x827 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x901 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x938 &  x940 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x977 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1018 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 &  x1130 & ~x198 & ~x237 & ~x276 & ~x315 & ~x354 & ~x594 & ~x918;
assign c128 =  x5 &  x8 &  x11 &  x17 &  x23 &  x29 &  x32 &  x35 &  x41 &  x44 &  x47 &  x53 &  x56 &  x62 &  x71 &  x74 &  x77 &  x89 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x134 &  x140 &  x143 &  x146 &  x149 &  x158 &  x161 &  x164 &  x167 &  x173 &  x185 &  x188 &  x191 &  x194 &  x203 &  x206 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x245 &  x248 &  x251 &  x260 &  x263 &  x266 &  x272 &  x281 &  x284 &  x287 &  x290 &  x293 &  x299 &  x302 &  x305 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x338 &  x344 &  x347 &  x350 &  x359 &  x365 &  x368 &  x377 &  x380 &  x383 &  x389 &  x392 &  x395 &  x398 &  x404 &  x406 &  x407 &  x410 &  x413 &  x416 &  x419 &  x431 &  x434 &  x437 &  x440 &  x446 &  x452 &  x455 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x485 &  x497 &  x500 &  x503 &  x509 &  x512 &  x518 &  x521 &  x524 &  x530 &  x533 &  x536 &  x539 &  x545 &  x548 &  x551 &  x566 &  x569 &  x572 &  x575 &  x584 &  x586 &  x590 &  x599 &  x605 &  x608 &  x617 &  x625 &  x626 &  x629 &  x632 &  x647 &  x653 &  x656 &  x659 &  x662 &  x664 &  x668 &  x671 &  x674 &  x677 &  x683 &  x689 &  x692 &  x695 &  x698 &  x701 &  x707 &  x712 &  x713 &  x719 &  x728 &  x731 &  x734 &  x740 &  x742 &  x749 &  x752 &  x755 &  x764 &  x767 &  x770 &  x776 &  x779 &  x782 &  x784 &  x788 &  x790 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x818 &  x824 &  x827 &  x828 &  x830 &  x833 &  x836 &  x839 &  x845 &  x848 &  x851 &  x854 &  x860 &  x862 &  x868 &  x869 &  x872 &  x875 &  x887 &  x890 &  x893 &  x896 &  x902 &  x904 &  x905 &  x908 &  x911 &  x914 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x965 &  x971 &  x977 &  x986 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1052 &  x1055 &  x1061 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1115 &  x1118 &  x1121 &  x1130 & ~x576 & ~x615 & ~x771 & ~x876;
assign c130 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x56 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x254 &  x257 &  x259 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x320 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x491 &  x494 &  x497 &  x503 &  x506 &  x512 &  x515 &  x518 &  x524 &  x527 &  x530 &  x533 &  x536 &  x542 &  x545 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x671 &  x674 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x833 &  x836 &  x842 &  x845 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x883 &  x884 &  x887 &  x890 &  x896 &  x899 &  x902 &  x908 &  x911 &  x914 &  x920 &  x922 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x961 &  x962 &  x968 &  x971 &  x974 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1000 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x276 & ~x435 & ~x474 & ~x684 & ~x723 & ~x777;
assign c132 =  x14 &  x17 &  x56 &  x62 &  x68 &  x77 &  x80 &  x86 &  x107 &  x110 &  x122 &  x128 &  x131 &  x152 &  x164 &  x197 &  x209 &  x212 &  x218 &  x221 &  x227 &  x230 &  x242 &  x266 &  x278 &  x284 &  x287 &  x293 &  x299 &  x302 &  x329 &  x347 &  x353 &  x362 &  x365 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x395 &  x398 &  x401 &  x404 &  x407 &  x425 &  x430 &  x431 &  x434 &  x440 &  x455 &  x461 &  x467 &  x470 &  x479 &  x482 &  x485 &  x488 &  x497 &  x503 &  x506 &  x509 &  x511 &  x524 &  x527 &  x533 &  x536 &  x542 &  x554 &  x560 &  x563 &  x566 &  x572 &  x578 &  x596 &  x602 &  x605 &  x617 &  x623 &  x626 &  x628 &  x629 &  x635 &  x638 &  x650 &  x653 &  x662 &  x665 &  x668 &  x670 &  x680 &  x683 &  x686 &  x695 &  x698 &  x701 &  x709 &  x710 &  x713 &  x716 &  x722 &  x728 &  x731 &  x740 &  x748 &  x755 &  x758 &  x785 &  x788 &  x791 &  x794 &  x803 &  x812 &  x824 &  x826 &  x827 &  x833 &  x839 &  x845 &  x848 &  x851 &  x865 &  x869 &  x872 &  x881 &  x884 &  x905 &  x908 &  x911 &  x920 &  x935 &  x938 &  x953 &  x959 &  x977 &  x983 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1022 &  x1034 &  x1043 &  x1052 &  x1055 &  x1079 &  x1085 &  x1109 &  x1115 & ~x459 & ~x1008 & ~x1029 & ~x1068 & ~x1086 & ~x1102;
assign c134 =  x1 &  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x22 &  x23 &  x26 &  x29 &  x32 &  x38 &  x40 &  x41 &  x44 &  x47 &  x50 &  x53 &  x55 &  x56 &  x59 &  x61 &  x62 &  x65 &  x68 &  x71 &  x74 &  x79 &  x80 &  x83 &  x86 &  x89 &  x92 &  x94 &  x95 &  x98 &  x100 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x118 &  x119 &  x122 &  x125 &  x131 &  x133 &  x134 &  x139 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x161 &  x164 &  x167 &  x170 &  x172 &  x176 &  x178 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x211 &  x212 &  x215 &  x217 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x250 &  x251 &  x256 &  x257 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x289 &  x290 &  x293 &  x295 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x328 &  x329 &  x331 &  x332 &  x334 &  x335 &  x338 &  x341 &  x343 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x367 &  x368 &  x371 &  x374 &  x377 &  x380 &  x382 &  x383 &  x386 &  x389 &  x392 &  x398 &  x401 &  x404 &  x406 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x445 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x484 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x562 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x601 &  x602 &  x605 &  x608 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x809 &  x812 &  x815 &  x818 &  x820 &  x821 &  x823 &  x824 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x898 &  x899 &  x901 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x937 &  x938 &  x940 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1015 &  x1016 &  x1018 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x954;
assign c136 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x47 &  x49 &  x56 &  x59 &  x62 &  x68 &  x71 &  x77 &  x83 &  x86 &  x89 &  x92 &  x93 &  x94 &  x95 &  x98 &  x101 &  x107 &  x110 &  x116 &  x119 &  x122 &  x125 &  x128 &  x132 &  x133 &  x137 &  x140 &  x143 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x172 &  x173 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x203 &  x206 &  x209 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x239 &  x242 &  x245 &  x251 &  x254 &  x257 &  x259 &  x263 &  x272 &  x275 &  x284 &  x287 &  x290 &  x293 &  x296 &  x298 &  x299 &  x305 &  x308 &  x314 &  x317 &  x320 &  x329 &  x332 &  x335 &  x338 &  x344 &  x347 &  x350 &  x356 &  x359 &  x362 &  x368 &  x374 &  x377 &  x386 &  x389 &  x392 &  x395 &  x398 &  x404 &  x407 &  x413 &  x416 &  x419 &  x425 &  x428 &  x434 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x464 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x503 &  x506 &  x509 &  x518 &  x521 &  x524 &  x527 &  x530 &  x539 &  x545 &  x548 &  x554 &  x560 &  x563 &  x572 &  x575 &  x578 &  x584 &  x587 &  x590 &  x592 &  x599 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x626 &  x631 &  x632 &  x635 &  x638 &  x644 &  x650 &  x656 &  x659 &  x662 &  x665 &  x668 &  x670 &  x671 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x707 &  x710 &  x713 &  x716 &  x722 &  x725 &  x728 &  x731 &  x734 &  x743 &  x746 &  x749 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x782 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x827 &  x830 &  x833 &  x845 &  x848 &  x857 &  x860 &  x863 &  x865 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x950 &  x956 &  x959 &  x962 &  x965 &  x971 &  x977 &  x983 &  x986 &  x989 &  x998 &  x1001 &  x1004 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1064 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127;
assign c138 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x154 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x317 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x349 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x388 &  x389 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x428 &  x431 &  x434 &  x437 &  x440 &  x446 &  x449 &  x452 &  x458 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x544 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x703 &  x704 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x742 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x773 &  x776 &  x779 &  x781 &  x782 &  x784 &  x785 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x898 &  x901 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x940 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x979 &  x980 &  x982 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1018 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x312 & ~x699;
assign c140 =  x2 &  x5 &  x14 &  x17 &  x20 &  x26 &  x32 &  x35 &  x41 &  x44 &  x47 &  x53 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x146 &  x149 &  x152 &  x158 &  x161 &  x167 &  x170 &  x173 &  x176 &  x182 &  x185 &  x188 &  x191 &  x203 &  x206 &  x215 &  x218 &  x224 &  x230 &  x233 &  x236 &  x242 &  x251 &  x254 &  x257 &  x272 &  x278 &  x284 &  x287 &  x290 &  x293 &  x296 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x350 &  x353 &  x359 &  x362 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x386 &  x392 &  x395 &  x398 &  x401 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x476 &  x479 &  x482 &  x485 &  x491 &  x494 &  x497 &  x500 &  x503 &  x509 &  x511 &  x515 &  x524 &  x527 &  x530 &  x536 &  x542 &  x545 &  x547 &  x548 &  x551 &  x554 &  x560 &  x566 &  x569 &  x572 &  x578 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x614 &  x620 &  x623 &  x626 &  x628 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x659 &  x665 &  x667 &  x668 &  x671 &  x674 &  x677 &  x680 &  x686 &  x689 &  x692 &  x704 &  x709 &  x710 &  x713 &  x716 &  x719 &  x722 &  x728 &  x731 &  x743 &  x748 &  x752 &  x755 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x787 &  x794 &  x797 &  x800 &  x803 &  x809 &  x812 &  x818 &  x824 &  x827 &  x833 &  x839 &  x842 &  x845 &  x848 &  x857 &  x860 &  x863 &  x865 &  x866 &  x869 &  x872 &  x875 &  x878 &  x887 &  x890 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x938 &  x941 &  x944 &  x947 &  x950 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x989 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1088 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x195 & ~x543 & ~x606 & ~x639 & ~x645 & ~x678 & ~x858 & ~x897 & ~x936 & ~x975 & ~x1014 & ~x1053;
assign c142 =  x2 &  x8 &  x17 &  x26 &  x35 &  x38 &  x41 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x89 &  x92 &  x98 &  x101 &  x113 &  x121 &  x122 &  x125 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x158 &  x160 &  x161 &  x164 &  x167 &  x170 &  x182 &  x188 &  x191 &  x200 &  x206 &  x209 &  x212 &  x221 &  x224 &  x227 &  x230 &  x233 &  x242 &  x245 &  x248 &  x257 &  x260 &  x263 &  x269 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x302 &  x316 &  x320 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x353 &  x356 &  x359 &  x368 &  x374 &  x377 &  x386 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x422 &  x428 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x455 &  x458 &  x461 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x488 &  x494 &  x500 &  x506 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x551 &  x554 &  x566 &  x569 &  x575 &  x578 &  x581 &  x593 &  x599 &  x608 &  x611 &  x629 &  x632 &  x638 &  x650 &  x656 &  x659 &  x662 &  x665 &  x671 &  x674 &  x676 &  x683 &  x686 &  x692 &  x698 &  x701 &  x713 &  x715 &  x725 &  x731 &  x740 &  x746 &  x749 &  x752 &  x758 &  x761 &  x767 &  x776 &  x779 &  x782 &  x788 &  x797 &  x803 &  x805 &  x809 &  x812 &  x824 &  x832 &  x836 &  x838 &  x844 &  x845 &  x848 &  x857 &  x860 &  x863 &  x866 &  x869 &  x881 &  x883 &  x884 &  x887 &  x893 &  x896 &  x899 &  x902 &  x905 &  x911 &  x917 &  x920 &  x922 &  x923 &  x926 &  x935 &  x947 &  x953 &  x956 &  x959 &  x968 &  x971 &  x974 &  x983 &  x989 &  x998 &  x1000 &  x1001 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1046 &  x1052 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1121 &  x1124 &  x1130 & ~x303 & ~x342 & ~x384 & ~x501 & ~x780 & ~x819;
assign c144 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x35 &  x41 &  x44 &  x47 &  x50 &  x53 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x122 &  x125 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x227 &  x236 &  x239 &  x242 &  x245 &  x248 &  x254 &  x263 &  x269 &  x275 &  x284 &  x290 &  x299 &  x305 &  x311 &  x326 &  x332 &  x335 &  x341 &  x344 &  x350 &  x353 &  x359 &  x368 &  x371 &  x376 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x410 &  x415 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x443 &  x449 &  x455 &  x458 &  x464 &  x467 &  x470 &  x476 &  x479 &  x482 &  x485 &  x488 &  x493 &  x494 &  x497 &  x500 &  x503 &  x509 &  x512 &  x518 &  x521 &  x536 &  x539 &  x542 &  x545 &  x551 &  x554 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x599 &  x602 &  x605 &  x611 &  x617 &  x620 &  x626 &  x629 &  x641 &  x650 &  x653 &  x656 &  x662 &  x665 &  x668 &  x671 &  x680 &  x683 &  x689 &  x692 &  x695 &  x698 &  x704 &  x713 &  x716 &  x722 &  x725 &  x731 &  x734 &  x737 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x767 &  x776 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x803 &  x806 &  x809 &  x812 &  x815 &  x821 &  x827 &  x830 &  x836 &  x839 &  x842 &  x845 &  x847 &  x851 &  x854 &  x857 &  x860 &  x863 &  x878 &  x881 &  x884 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x956 &  x959 &  x965 &  x968 &  x971 &  x977 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1013 &  x1016 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1097 &  x1100 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x684 & ~x738 & ~x777 & ~x813 & ~x912;
assign c146 =  x2 &  x8 &  x14 &  x17 &  x26 &  x29 &  x32 &  x38 &  x41 &  x47 &  x53 &  x65 &  x83 &  x89 &  x92 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x143 &  x146 &  x149 &  x155 &  x164 &  x167 &  x179 &  x182 &  x188 &  x191 &  x194 &  x197 &  x209 &  x212 &  x215 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x272 &  x275 &  x277 &  x281 &  x284 &  x287 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x323 &  x326 &  x332 &  x335 &  x338 &  x341 &  x355 &  x356 &  x362 &  x365 &  x377 &  x383 &  x389 &  x394 &  x395 &  x398 &  x401 &  x407 &  x410 &  x413 &  x419 &  x422 &  x425 &  x428 &  x431 &  x433 &  x434 &  x440 &  x443 &  x449 &  x452 &  x458 &  x467 &  x476 &  x478 &  x479 &  x482 &  x485 &  x497 &  x506 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x542 &  x553 &  x554 &  x560 &  x563 &  x566 &  x572 &  x575 &  x584 &  x587 &  x592 &  x596 &  x605 &  x608 &  x617 &  x620 &  x629 &  x638 &  x647 &  x650 &  x653 &  x655 &  x662 &  x665 &  x668 &  x671 &  x674 &  x680 &  x683 &  x686 &  x688 &  x689 &  x694 &  x695 &  x701 &  x710 &  x713 &  x719 &  x722 &  x725 &  x727 &  x728 &  x733 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x758 &  x764 &  x767 &  x770 &  x772 &  x779 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x806 &  x811 &  x815 &  x818 &  x821 &  x827 &  x830 &  x836 &  x839 &  x845 &  x848 &  x857 &  x863 &  x866 &  x869 &  x872 &  x878 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x908 &  x911 &  x914 &  x922 &  x923 &  x926 &  x941 &  x944 &  x947 &  x950 &  x959 &  x965 &  x971 &  x986 &  x989 &  x992 &  x995 &  x1007 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1127 & ~x303 & ~x405 & ~x444 & ~x546 & ~x624 & ~x625 & ~x663 & ~x702 & ~x703 & ~x741 & ~x742 & ~x780 & ~x819 & ~x858 & ~x897 & ~x936;
assign c148 =  x17 &  x20 &  x26 &  x35 &  x44 &  x68 &  x77 &  x83 &  x86 &  x95 &  x98 &  x107 &  x110 &  x128 &  x143 &  x146 &  x179 &  x191 &  x194 &  x197 &  x200 &  x251 &  x254 &  x266 &  x272 &  x284 &  x314 &  x338 &  x350 &  x353 &  x356 &  x358 &  x362 &  x365 &  x374 &  x380 &  x397 &  x398 &  x404 &  x407 &  x428 &  x437 &  x443 &  x461 &  x467 &  x470 &  x473 &  x475 &  x476 &  x494 &  x497 &  x500 &  x518 &  x542 &  x548 &  x554 &  x563 &  x572 &  x581 &  x593 &  x608 &  x614 &  x620 &  x632 &  x635 &  x638 &  x641 &  x644 &  x653 &  x662 &  x665 &  x671 &  x686 &  x689 &  x692 &  x701 &  x710 &  x722 &  x734 &  x737 &  x740 &  x752 &  x755 &  x779 &  x785 &  x797 &  x808 &  x812 &  x827 &  x851 &  x854 &  x860 &  x884 &  x893 &  x896 &  x902 &  x914 &  x932 &  x941 &  x944 &  x953 &  x980 &  x1004 &  x1007 &  x1010 &  x1037 &  x1043 &  x1058 &  x1061 &  x1067 &  x1070 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1100 &  x1115 &  x1124 & ~x67 & ~x105 & ~x249 & ~x468 & ~x483;
assign c150 =  x5 &  x8 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x53 &  x56 &  x59 &  x62 &  x67 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x104 &  x107 &  x113 &  x116 &  x119 &  x128 &  x134 &  x137 &  x140 &  x143 &  x152 &  x155 &  x161 &  x164 &  x173 &  x176 &  x179 &  x188 &  x191 &  x197 &  x206 &  x209 &  x218 &  x227 &  x233 &  x239 &  x242 &  x248 &  x251 &  x260 &  x269 &  x272 &  x275 &  x278 &  x290 &  x293 &  x295 &  x302 &  x305 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x347 &  x350 &  x356 &  x362 &  x368 &  x374 &  x380 &  x386 &  x389 &  x398 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x427 &  x434 &  x440 &  x443 &  x446 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x494 &  x500 &  x503 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x545 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x590 &  x593 &  x602 &  x605 &  x608 &  x614 &  x617 &  x623 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x659 &  x662 &  x664 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x689 &  x692 &  x695 &  x698 &  x701 &  x703 &  x704 &  x713 &  x716 &  x722 &  x725 &  x734 &  x740 &  x742 &  x743 &  x749 &  x755 &  x758 &  x761 &  x767 &  x770 &  x773 &  x776 &  x782 &  x791 &  x797 &  x800 &  x803 &  x809 &  x815 &  x818 &  x821 &  x823 &  x827 &  x833 &  x839 &  x842 &  x845 &  x848 &  x859 &  x860 &  x863 &  x866 &  x869 &  x872 &  x878 &  x881 &  x884 &  x887 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x938 &  x941 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1058 &  x1061 &  x1070 &  x1073 &  x1076 &  x1082 &  x1088 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x276 & ~x354 & ~x432 & ~x588 & ~x753 & ~x915 & ~x954 & ~x993 & ~x1032 & ~x1065 & ~x1104;
assign c152 =  x5 &  x11 &  x16 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x44 &  x55 &  x56 &  x65 &  x71 &  x74 &  x83 &  x86 &  x88 &  x89 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x134 &  x137 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x176 &  x179 &  x182 &  x188 &  x194 &  x197 &  x203 &  x206 &  x218 &  x221 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x257 &  x266 &  x269 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x314 &  x317 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x353 &  x359 &  x362 &  x365 &  x368 &  x371 &  x380 &  x383 &  x386 &  x389 &  x392 &  x401 &  x404 &  x407 &  x413 &  x416 &  x419 &  x425 &  x431 &  x434 &  x437 &  x440 &  x443 &  x449 &  x461 &  x464 &  x470 &  x473 &  x479 &  x485 &  x488 &  x491 &  x494 &  x497 &  x506 &  x512 &  x515 &  x521 &  x524 &  x530 &  x536 &  x539 &  x542 &  x545 &  x548 &  x554 &  x556 &  x557 &  x563 &  x566 &  x569 &  x572 &  x578 &  x584 &  x587 &  x596 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x638 &  x641 &  x644 &  x647 &  x650 &  x656 &  x659 &  x665 &  x668 &  x674 &  x677 &  x683 &  x686 &  x692 &  x698 &  x707 &  x710 &  x713 &  x728 &  x731 &  x734 &  x737 &  x742 &  x743 &  x746 &  x751 &  x752 &  x764 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x794 &  x797 &  x800 &  x806 &  x815 &  x818 &  x824 &  x827 &  x830 &  x836 &  x842 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x868 &  x872 &  x878 &  x881 &  x884 &  x890 &  x893 &  x898 &  x899 &  x908 &  x911 &  x914 &  x920 &  x926 &  x929 &  x935 &  x937 &  x938 &  x941 &  x946 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x964 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x985 &  x986 &  x992 &  x998 &  x1001 &  x1004 &  x1013 &  x1016 &  x1019 &  x1024 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1042 &  x1043 &  x1046 &  x1055 &  x1063 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1081 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1120 &  x1121 &  x1124 &  x1127 &  x1130 & ~x543 & ~x621 & ~x660 & ~x777;
assign c154 =  x5 &  x8 &  x17 &  x20 &  x35 &  x44 &  x53 &  x56 &  x68 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x92 &  x98 &  x110 &  x113 &  x116 &  x119 &  x125 &  x143 &  x152 &  x155 &  x158 &  x173 &  x176 &  x179 &  x182 &  x185 &  x197 &  x203 &  x209 &  x212 &  x221 &  x227 &  x233 &  x236 &  x242 &  x245 &  x251 &  x257 &  x266 &  x269 &  x284 &  x293 &  x302 &  x317 &  x341 &  x347 &  x350 &  x356 &  x359 &  x365 &  x374 &  x386 &  x389 &  x392 &  x395 &  x398 &  x404 &  x407 &  x410 &  x413 &  x419 &  x422 &  x425 &  x431 &  x433 &  x443 &  x449 &  x452 &  x455 &  x470 &  x472 &  x476 &  x479 &  x482 &  x485 &  x491 &  x497 &  x511 &  x521 &  x536 &  x539 &  x542 &  x545 &  x548 &  x550 &  x551 &  x557 &  x560 &  x566 &  x572 &  x578 &  x581 &  x587 &  x593 &  x599 &  x602 &  x605 &  x614 &  x626 &  x641 &  x653 &  x656 &  x659 &  x668 &  x674 &  x680 &  x686 &  x695 &  x701 &  x704 &  x707 &  x709 &  x719 &  x731 &  x737 &  x743 &  x746 &  x748 &  x749 &  x752 &  x755 &  x764 &  x773 &  x776 &  x788 &  x791 &  x794 &  x797 &  x800 &  x806 &  x812 &  x818 &  x821 &  x826 &  x827 &  x830 &  x839 &  x857 &  x863 &  x869 &  x875 &  x878 &  x881 &  x899 &  x905 &  x908 &  x911 &  x914 &  x916 &  x920 &  x929 &  x932 &  x938 &  x950 &  x953 &  x955 &  x956 &  x959 &  x962 &  x965 &  x977 &  x980 &  x986 &  x989 &  x994 &  x995 &  x998 &  x1028 &  x1032 &  x1034 &  x1037 &  x1049 &  x1055 &  x1058 &  x1061 &  x1067 &  x1070 &  x1071 &  x1082 &  x1088 &  x1091 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 & ~x528 & ~x780 & ~x819 & ~x858 & ~x936 & ~x975;
assign c156 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x50 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x82 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x113 &  x119 &  x122 &  x128 &  x131 &  x137 &  x140 &  x143 &  x158 &  x164 &  x170 &  x173 &  x176 &  x179 &  x182 &  x191 &  x194 &  x199 &  x206 &  x209 &  x212 &  x218 &  x224 &  x227 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x277 &  x278 &  x281 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x308 &  x311 &  x314 &  x317 &  x320 &  x326 &  x329 &  x332 &  x335 &  x338 &  x347 &  x350 &  x353 &  x355 &  x356 &  x359 &  x362 &  x371 &  x374 &  x380 &  x383 &  x386 &  x389 &  x395 &  x398 &  x400 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x437 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x467 &  x470 &  x476 &  x482 &  x485 &  x491 &  x494 &  x497 &  x509 &  x512 &  x514 &  x515 &  x527 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x553 &  x557 &  x566 &  x569 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x605 &  x608 &  x610 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x649 &  x650 &  x653 &  x655 &  x656 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x688 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x727 &  x730 &  x731 &  x734 &  x737 &  x740 &  x743 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x766 &  x767 &  x769 &  x773 &  x779 &  x785 &  x788 &  x794 &  x800 &  x803 &  x805 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x836 &  x839 &  x842 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x905 &  x911 &  x920 &  x922 &  x923 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x977 &  x980 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x468 & ~x507 & ~x522 & ~x585 & ~x624 & ~x663 & ~x741;
assign c158 =  x8 &  x11 &  x14 &  x23 &  x35 &  x38 &  x47 &  x62 &  x65 &  x68 &  x74 &  x80 &  x89 &  x104 &  x107 &  x122 &  x125 &  x155 &  x158 &  x167 &  x170 &  x173 &  x185 &  x191 &  x197 &  x206 &  x212 &  x215 &  x218 &  x221 &  x227 &  x233 &  x236 &  x238 &  x242 &  x245 &  x248 &  x260 &  x272 &  x277 &  x281 &  x290 &  x293 &  x296 &  x305 &  x308 &  x316 &  x320 &  x323 &  x332 &  x338 &  x341 &  x347 &  x350 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x383 &  x386 &  x389 &  x392 &  x394 &  x395 &  x404 &  x413 &  x416 &  x419 &  x425 &  x437 &  x443 &  x446 &  x449 &  x452 &  x458 &  x461 &  x470 &  x472 &  x473 &  x485 &  x488 &  x494 &  x497 &  x503 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x545 &  x554 &  x557 &  x560 &  x563 &  x572 &  x578 &  x584 &  x587 &  x596 &  x599 &  x605 &  x611 &  x614 &  x617 &  x623 &  x626 &  x632 &  x637 &  x638 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x670 &  x680 &  x686 &  x689 &  x695 &  x701 &  x707 &  x710 &  x715 &  x716 &  x722 &  x728 &  x734 &  x746 &  x758 &  x764 &  x770 &  x773 &  x778 &  x779 &  x782 &  x785 &  x788 &  x791 &  x793 &  x800 &  x803 &  x806 &  x809 &  x812 &  x821 &  x824 &  x832 &  x833 &  x836 &  x839 &  x845 &  x857 &  x860 &  x866 &  x871 &  x872 &  x881 &  x883 &  x884 &  x887 &  x896 &  x899 &  x902 &  x910 &  x922 &  x923 &  x929 &  x935 &  x941 &  x947 &  x950 &  x953 &  x961 &  x974 &  x977 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1006 &  x1007 &  x1013 &  x1016 &  x1022 &  x1025 &  x1031 &  x1045 &  x1046 &  x1052 &  x1058 &  x1061 &  x1067 &  x1076 &  x1078 &  x1079 &  x1088 &  x1090 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1117 &  x1118 & ~x303 & ~x525 & ~x780 & ~x858 & ~x936 & ~x975;
assign c160 =  x2 &  x5 &  x8 &  x14 &  x17 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x74 &  x76 &  x77 &  x83 &  x86 &  x89 &  x92 &  x104 &  x107 &  x110 &  x116 &  x122 &  x125 &  x128 &  x131 &  x137 &  x140 &  x143 &  x149 &  x154 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x181 &  x182 &  x185 &  x188 &  x193 &  x194 &  x203 &  x206 &  x212 &  x218 &  x221 &  x226 &  x230 &  x233 &  x236 &  x242 &  x245 &  x248 &  x251 &  x254 &  x256 &  x257 &  x260 &  x265 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x293 &  x296 &  x299 &  x304 &  x308 &  x320 &  x323 &  x326 &  x329 &  x332 &  x338 &  x341 &  x343 &  x344 &  x347 &  x353 &  x356 &  x359 &  x365 &  x368 &  x371 &  x377 &  x383 &  x392 &  x395 &  x398 &  x404 &  x407 &  x413 &  x419 &  x425 &  x428 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x470 &  x476 &  x479 &  x482 &  x494 &  x497 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x539 &  x545 &  x551 &  x554 &  x560 &  x563 &  x566 &  x569 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x659 &  x662 &  x665 &  x668 &  x671 &  x680 &  x683 &  x686 &  x692 &  x698 &  x701 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x731 &  x734 &  x737 &  x740 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x784 &  x785 &  x788 &  x794 &  x797 &  x800 &  x803 &  x806 &  x812 &  x815 &  x821 &  x823 &  x824 &  x830 &  x836 &  x842 &  x848 &  x851 &  x854 &  x857 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x893 &  x896 &  x899 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x944 &  x947 &  x950 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1000 &  x1001 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1039 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1067 &  x1070 &  x1073 &  x1076 &  x1078 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1112 &  x1115 &  x1117 &  x1118 &  x1121 &  x1127 &  x1130 & ~x195 & ~x234 & ~x273 & ~x312 & ~x351 & ~x354;
assign c162 =  x2 &  x11 &  x20 &  x23 &  x32 &  x35 &  x38 &  x44 &  x50 &  x56 &  x62 &  x68 &  x71 &  x74 &  x77 &  x110 &  x116 &  x121 &  x128 &  x134 &  x140 &  x146 &  x155 &  x160 &  x161 &  x164 &  x170 &  x182 &  x188 &  x191 &  x194 &  x199 &  x200 &  x209 &  x215 &  x218 &  x221 &  x227 &  x230 &  x239 &  x242 &  x245 &  x257 &  x263 &  x266 &  x277 &  x278 &  x281 &  x290 &  x293 &  x302 &  x314 &  x316 &  x338 &  x344 &  x350 &  x353 &  x355 &  x365 &  x371 &  x374 &  x383 &  x386 &  x394 &  x398 &  x401 &  x413 &  x416 &  x431 &  x436 &  x440 &  x443 &  x461 &  x464 &  x473 &  x474 &  x478 &  x479 &  x485 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x512 &  x513 &  x514 &  x515 &  x517 &  x518 &  x521 &  x524 &  x530 &  x536 &  x539 &  x542 &  x548 &  x553 &  x554 &  x557 &  x560 &  x566 &  x569 &  x572 &  x578 &  x581 &  x584 &  x587 &  x590 &  x592 &  x593 &  x596 &  x602 &  x605 &  x608 &  x616 &  x620 &  x631 &  x635 &  x638 &  x644 &  x647 &  x650 &  x656 &  x659 &  x662 &  x670 &  x674 &  x683 &  x686 &  x698 &  x704 &  x707 &  x713 &  x716 &  x719 &  x731 &  x740 &  x752 &  x761 &  x764 &  x776 &  x782 &  x785 &  x788 &  x791 &  x794 &  x812 &  x818 &  x821 &  x827 &  x836 &  x839 &  x842 &  x857 &  x860 &  x866 &  x875 &  x884 &  x887 &  x899 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x938 &  x941 &  x944 &  x947 &  x950 &  x956 &  x962 &  x971 &  x974 &  x1001 &  x1010 &  x1016 &  x1019 &  x1022 &  x1031 &  x1034 &  x1037 &  x1043 &  x1061 &  x1067 &  x1070 &  x1079 &  x1082 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1130 & ~x444 & ~x705 & ~x744 & ~x783;
assign c164 =  x2 &  x5 &  x8 &  x11 &  x17 &  x23 &  x26 &  x29 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x116 &  x125 &  x134 &  x140 &  x143 &  x146 &  x155 &  x158 &  x161 &  x167 &  x170 &  x173 &  x182 &  x185 &  x188 &  x190 &  x191 &  x197 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x224 &  x230 &  x233 &  x245 &  x248 &  x251 &  x254 &  x260 &  x263 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x320 &  x323 &  x338 &  x341 &  x344 &  x356 &  x359 &  x365 &  x380 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x437 &  x440 &  x443 &  x445 &  x446 &  x449 &  x452 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x521 &  x524 &  x527 &  x533 &  x539 &  x548 &  x551 &  x554 &  x557 &  x563 &  x569 &  x575 &  x578 &  x581 &  x586 &  x593 &  x596 &  x605 &  x611 &  x614 &  x617 &  x620 &  x623 &  x625 &  x626 &  x629 &  x632 &  x635 &  x638 &  x644 &  x650 &  x656 &  x659 &  x662 &  x664 &  x665 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x703 &  x707 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x740 &  x742 &  x743 &  x746 &  x752 &  x755 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x791 &  x794 &  x797 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x833 &  x836 &  x839 &  x842 &  x848 &  x857 &  x863 &  x866 &  x872 &  x878 &  x884 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x953 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1046 &  x1049 &  x1058 &  x1061 &  x1064 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1118 &  x1121 & ~x237 & ~x276 & ~x315 & ~x354 & ~x360 & ~x399 & ~x435 & ~x438 & ~x474 & ~x513 & ~x552 & ~x597 & ~x636;
assign c166 =  x5 &  x14 &  x20 &  x23 &  x29 &  x32 &  x35 &  x47 &  x50 &  x53 &  x56 &  x59 &  x68 &  x74 &  x83 &  x95 &  x98 &  x104 &  x110 &  x113 &  x116 &  x119 &  x125 &  x128 &  x134 &  x149 &  x152 &  x161 &  x167 &  x170 &  x182 &  x185 &  x194 &  x206 &  x212 &  x218 &  x230 &  x239 &  x242 &  x245 &  x248 &  x254 &  x260 &  x263 &  x269 &  x272 &  x275 &  x281 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x323 &  x326 &  x329 &  x332 &  x338 &  x341 &  x347 &  x350 &  x353 &  x362 &  x382 &  x389 &  x392 &  x398 &  x404 &  x407 &  x410 &  x413 &  x415 &  x416 &  x421 &  x422 &  x425 &  x428 &  x431 &  x437 &  x440 &  x443 &  x446 &  x448 &  x452 &  x455 &  x461 &  x473 &  x476 &  x479 &  x482 &  x485 &  x487 &  x500 &  x503 &  x509 &  x512 &  x518 &  x521 &  x530 &  x533 &  x536 &  x542 &  x548 &  x551 &  x554 &  x560 &  x563 &  x565 &  x566 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x602 &  x605 &  x611 &  x614 &  x617 &  x623 &  x632 &  x635 &  x638 &  x641 &  x647 &  x662 &  x665 &  x671 &  x689 &  x692 &  x701 &  x704 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x746 &  x749 &  x752 &  x755 &  x758 &  x764 &  x773 &  x785 &  x794 &  x797 &  x800 &  x809 &  x812 &  x815 &  x818 &  x820 &  x821 &  x827 &  x836 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x859 &  x860 &  x863 &  x875 &  x878 &  x881 &  x884 &  x896 &  x902 &  x908 &  x911 &  x914 &  x920 &  x926 &  x935 &  x937 &  x940 &  x941 &  x950 &  x953 &  x956 &  x962 &  x977 &  x979 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1010 &  x1016 &  x1019 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1057 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1082 &  x1085 &  x1094 &  x1097 &  x1100 &  x1103 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x126 & ~x282 & ~x360 & ~x399 & ~x432 & ~x438 & ~x471 & ~x477 & ~x594 & ~x699;
assign c168 =  x2 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x107 &  x113 &  x116 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x265 &  x266 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x343 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x409 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x448 &  x449 &  x452 &  x455 &  x458 &  x464 &  x467 &  x470 &  x473 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x509 &  x512 &  x515 &  x518 &  x521 &  x523 &  x524 &  x527 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x710 &  x713 &  x716 &  x722 &  x725 &  x728 &  x734 &  x737 &  x740 &  x743 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x971 &  x974 &  x977 &  x983 &  x986 &  x989 &  x992 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x360 & ~x399 & ~x438 & ~x477 & ~x516 & ~x555 & ~x594 & ~x660 & ~x699 & ~x711 & ~x777 & ~x816 & ~x855;
assign c170 =  x2 &  x5 &  x14 &  x17 &  x20 &  x22 &  x23 &  x29 &  x32 &  x38 &  x50 &  x53 &  x60 &  x68 &  x71 &  x74 &  x86 &  x89 &  x92 &  x94 &  x95 &  x107 &  x113 &  x116 &  x119 &  x122 &  x125 &  x131 &  x134 &  x143 &  x145 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x172 &  x173 &  x182 &  x184 &  x188 &  x194 &  x203 &  x205 &  x206 &  x211 &  x212 &  x215 &  x218 &  x221 &  x223 &  x233 &  x236 &  x239 &  x242 &  x245 &  x250 &  x251 &  x254 &  x257 &  x260 &  x262 &  x263 &  x266 &  x269 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x301 &  x302 &  x304 &  x305 &  x311 &  x314 &  x320 &  x323 &  x329 &  x332 &  x335 &  x338 &  x340 &  x341 &  x344 &  x350 &  x353 &  x356 &  x362 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x395 &  x401 &  x406 &  x407 &  x410 &  x413 &  x419 &  x422 &  x425 &  x428 &  x440 &  x443 &  x446 &  x455 &  x461 &  x464 &  x467 &  x473 &  x479 &  x482 &  x485 &  x488 &  x494 &  x497 &  x500 &  x503 &  x506 &  x512 &  x515 &  x527 &  x530 &  x533 &  x545 &  x551 &  x554 &  x557 &  x563 &  x569 &  x572 &  x575 &  x578 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x611 &  x614 &  x620 &  x623 &  x632 &  x635 &  x644 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x674 &  x677 &  x680 &  x692 &  x716 &  x722 &  x725 &  x728 &  x734 &  x740 &  x743 &  x758 &  x770 &  x779 &  x782 &  x788 &  x791 &  x794 &  x800 &  x806 &  x809 &  x812 &  x815 &  x821 &  x827 &  x829 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x857 &  x860 &  x863 &  x869 &  x878 &  x881 &  x887 &  x890 &  x896 &  x899 &  x905 &  x908 &  x914 &  x917 &  x923 &  x926 &  x929 &  x935 &  x938 &  x947 &  x950 &  x956 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1052 &  x1055 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1124;
assign c172 =  x2 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x184 &  x185 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x368 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x431 &  x434 &  x437 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x497 &  x500 &  x503 &  x509 &  x511 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x550 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x665 &  x668 &  x670 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x698 &  x704 &  x706 &  x707 &  x709 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x740 &  x743 &  x746 &  x747 &  x748 &  x752 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x786 &  x787 &  x791 &  x794 &  x797 &  x806 &  x809 &  x812 &  x815 &  x821 &  x824 &  x826 &  x827 &  x830 &  x836 &  x842 &  x845 &  x854 &  x857 &  x865 &  x866 &  x869 &  x875 &  x878 &  x881 &  x884 &  x890 &  x893 &  x896 &  x899 &  x904 &  x905 &  x908 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1010 &  x1016 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x156 & ~x195 & ~x639 & ~x678 & ~x741 & ~x780 & ~x819 & ~x897 & ~x936 & ~x975 & ~x1053;
assign c174 =  x2 &  x8 &  x11 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x113 &  x116 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x194 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x230 &  x236 &  x238 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x277 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x316 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x355 &  x359 &  x362 &  x365 &  x368 &  x371 &  x380 &  x383 &  x389 &  x392 &  x394 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x428 &  x431 &  x433 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x497 &  x500 &  x503 &  x506 &  x509 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x548 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x662 &  x665 &  x671 &  x674 &  x677 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x709 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x740 &  x743 &  x746 &  x748 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x766 &  x767 &  x770 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x800 &  x803 &  x805 &  x806 &  x809 &  x812 &  x815 &  x818 &  x824 &  x827 &  x830 &  x833 &  x836 &  x842 &  x845 &  x848 &  x854 &  x857 &  x860 &  x866 &  x869 &  x872 &  x875 &  x881 &  x883 &  x884 &  x887 &  x890 &  x893 &  x896 &  x905 &  x908 &  x911 &  x917 &  x920 &  x922 &  x923 &  x926 &  x928 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x967 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1000 &  x1001 &  x1004 &  x1007 &  x1010 &  x1012 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1067 &  x1070 &  x1072 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x342 & ~x561 & ~x600 & ~x639 & ~x723 & ~x741 & ~x780 & ~x858 & ~x897 & ~x936 & ~x975;
assign c176 =  x2 &  x8 &  x17 &  x26 &  x35 &  x38 &  x40 &  x47 &  x53 &  x65 &  x68 &  x74 &  x86 &  x89 &  x92 &  x98 &  x107 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x149 &  x164 &  x170 &  x173 &  x176 &  x185 &  x197 &  x203 &  x206 &  x215 &  x224 &  x230 &  x257 &  x269 &  x272 &  x275 &  x278 &  x281 &  x290 &  x299 &  x302 &  x305 &  x311 &  x317 &  x338 &  x341 &  x344 &  x350 &  x353 &  x356 &  x359 &  x368 &  x371 &  x374 &  x380 &  x383 &  x410 &  x419 &  x428 &  x431 &  x437 &  x440 &  x443 &  x446 &  x452 &  x473 &  x479 &  x482 &  x503 &  x515 &  x518 &  x533 &  x539 &  x542 &  x548 &  x551 &  x557 &  x563 &  x569 &  x575 &  x578 &  x584 &  x590 &  x593 &  x596 &  x599 &  x602 &  x614 &  x617 &  x626 &  x638 &  x641 &  x644 &  x647 &  x653 &  x665 &  x668 &  x671 &  x674 &  x683 &  x686 &  x704 &  x710 &  x719 &  x722 &  x734 &  x737 &  x740 &  x749 &  x755 &  x770 &  x776 &  x782 &  x785 &  x794 &  x797 &  x800 &  x809 &  x815 &  x818 &  x824 &  x827 &  x839 &  x842 &  x872 &  x881 &  x884 &  x887 &  x890 &  x902 &  x908 &  x911 &  x914 &  x920 &  x926 &  x929 &  x941 &  x947 &  x953 &  x956 &  x965 &  x971 &  x977 &  x983 &  x986 &  x995 &  x1007 &  x1010 &  x1013 &  x1019 &  x1031 &  x1037 &  x1052 &  x1055 &  x1058 &  x1064 &  x1070 &  x1076 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x6 & ~x378 & ~x417 & ~x426 & ~x783 & ~x822 & ~x861 & ~x948 & ~x987;
assign c178 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x509 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x628 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x667 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x156 & ~x195 & ~x435 & ~x474 & ~x582 & ~x723 & ~x951 & ~x990 & ~x1029 & ~x1068;
assign c180 =  x2 &  x5 &  x11 &  x20 &  x26 &  x29 &  x32 &  x41 &  x44 &  x47 &  x50 &  x53 &  x59 &  x62 &  x65 &  x89 &  x92 &  x95 &  x98 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x128 &  x134 &  x137 &  x140 &  x146 &  x149 &  x155 &  x158 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x188 &  x194 &  x197 &  x200 &  x203 &  x209 &  x215 &  x221 &  x224 &  x227 &  x233 &  x236 &  x242 &  x251 &  x257 &  x260 &  x266 &  x272 &  x275 &  x281 &  x287 &  x290 &  x293 &  x299 &  x302 &  x305 &  x311 &  x314 &  x317 &  x323 &  x326 &  x338 &  x341 &  x347 &  x350 &  x359 &  x362 &  x371 &  x374 &  x377 &  x380 &  x389 &  x395 &  x401 &  x404 &  x407 &  x410 &  x413 &  x422 &  x425 &  x428 &  x433 &  x434 &  x437 &  x440 &  x443 &  x449 &  x458 &  x467 &  x470 &  x472 &  x476 &  x485 &  x491 &  x497 &  x500 &  x511 &  x512 &  x515 &  x521 &  x524 &  x536 &  x539 &  x545 &  x554 &  x557 &  x560 &  x566 &  x569 &  x572 &  x575 &  x581 &  x584 &  x587 &  x589 &  x593 &  x596 &  x599 &  x614 &  x617 &  x626 &  x628 &  x629 &  x632 &  x638 &  x650 &  x653 &  x656 &  x668 &  x671 &  x674 &  x680 &  x686 &  x695 &  x698 &  x704 &  x706 &  x707 &  x709 &  x710 &  x716 &  x722 &  x725 &  x728 &  x743 &  x746 &  x747 &  x758 &  x764 &  x773 &  x779 &  x782 &  x785 &  x791 &  x794 &  x800 &  x803 &  x809 &  x812 &  x815 &  x821 &  x826 &  x827 &  x833 &  x839 &  x842 &  x845 &  x854 &  x857 &  x860 &  x863 &  x865 &  x866 &  x872 &  x875 &  x878 &  x883 &  x887 &  x890 &  x896 &  x899 &  x904 &  x905 &  x908 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x943 &  x944 &  x953 &  x956 &  x959 &  x961 &  x962 &  x971 &  x974 &  x989 &  x992 &  x995 &  x1000 &  x1004 &  x1007 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1039 &  x1046 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1085 &  x1088 &  x1097 &  x1100 &  x1103 &  x1109 &  x1115 &  x1117 &  x1130 & ~x255 & ~x618 & ~x657 & ~x663 & ~x741 & ~x819 & ~x858 & ~x897 & ~x975 & ~x1014;
assign c182 =  x2 &  x5 &  x8 &  x11 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x155 &  x158 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x206 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x239 &  x242 &  x245 &  x248 &  x251 &  x257 &  x260 &  x263 &  x272 &  x275 &  x278 &  x281 &  x284 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x380 &  x382 &  x386 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x421 &  x422 &  x425 &  x431 &  x434 &  x440 &  x446 &  x448 &  x449 &  x452 &  x454 &  x455 &  x458 &  x460 &  x461 &  x464 &  x467 &  x473 &  x479 &  x482 &  x485 &  x487 &  x488 &  x491 &  x493 &  x494 &  x497 &  x500 &  x509 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x551 &  x554 &  x557 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x596 &  x599 &  x601 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x640 &  x641 &  x644 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x679 &  x683 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x779 &  x782 &  x785 &  x788 &  x794 &  x797 &  x803 &  x809 &  x812 &  x818 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x872 &  x878 &  x884 &  x887 &  x890 &  x893 &  x902 &  x905 &  x911 &  x914 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x937 &  x940 &  x941 &  x944 &  x947 &  x956 &  x962 &  x965 &  x968 &  x971 &  x974 &  x976 &  x979 &  x980 &  x983 &  x986 &  x989 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1015 &  x1016 &  x1018 &  x1019 &  x1022 &  x1025 &  x1034 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1057 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1096 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x351 & ~x354 & ~x429 & ~x432 & ~x549 & ~x588 & ~x594 & ~x1071;
assign c184 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x47 &  x50 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x140 &  x143 &  x146 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x227 &  x230 &  x233 &  x236 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x550 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x584 &  x587 &  x589 &  x590 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x626 &  x628 &  x629 &  x632 &  x635 &  x638 &  x644 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x667 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x743 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x904 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x935 &  x938 &  x941 &  x943 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x345 & ~x357 & ~x435 & ~x858 & ~x897 & ~x918 & ~x936 & ~x957 & ~x975 & ~x990 & ~x996 & ~x1008 & ~x1014 & ~x1029 & ~x1035 & ~x1047 & ~x1062 & ~x1068 & ~x1101;
assign c186 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x55 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x167 &  x170 &  x173 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x230 &  x233 &  x239 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x323 &  x326 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x458 &  x461 &  x464 &  x473 &  x476 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x593 &  x596 &  x599 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x698 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x731 &  x734 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x797 &  x800 &  x803 &  x815 &  x818 &  x824 &  x826 &  x827 &  x829 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x865 &  x866 &  x868 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x905 &  x907 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x945 &  x946 &  x947 &  x950 &  x953 &  x962 &  x968 &  x971 &  x974 &  x977 &  x980 &  x982 &  x983 &  x985 &  x986 &  x989 &  x992 &  x1001 &  x1004 &  x1007 &  x1016 &  x1019 &  x1021 &  x1024 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1061 &  x1063 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x351;
assign c188 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x41 &  x44 &  x50 &  x52 &  x56 &  x65 &  x68 &  x71 &  x74 &  x77 &  x83 &  x98 &  x107 &  x116 &  x119 &  x122 &  x130 &  x131 &  x137 &  x140 &  x146 &  x149 &  x152 &  x155 &  x164 &  x167 &  x179 &  x182 &  x188 &  x197 &  x202 &  x203 &  x206 &  x208 &  x212 &  x221 &  x224 &  x230 &  x241 &  x247 &  x248 &  x254 &  x272 &  x280 &  x286 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x317 &  x320 &  x325 &  x326 &  x332 &  x335 &  x338 &  x341 &  x344 &  x350 &  x353 &  x356 &  x359 &  x362 &  x374 &  x376 &  x377 &  x380 &  x382 &  x383 &  x389 &  x395 &  x398 &  x401 &  x404 &  x407 &  x413 &  x416 &  x422 &  x425 &  x434 &  x437 &  x446 &  x449 &  x455 &  x461 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x494 &  x497 &  x503 &  x512 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x545 &  x551 &  x554 &  x557 &  x581 &  x584 &  x587 &  x590 &  x593 &  x602 &  x605 &  x608 &  x614 &  x623 &  x626 &  x629 &  x632 &  x638 &  x641 &  x647 &  x650 &  x656 &  x662 &  x665 &  x668 &  x671 &  x674 &  x676 &  x680 &  x686 &  x698 &  x701 &  x704 &  x707 &  x713 &  x715 &  x716 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x746 &  x752 &  x764 &  x770 &  x773 &  x776 &  x782 &  x785 &  x788 &  x791 &  x797 &  x803 &  x809 &  x815 &  x824 &  x827 &  x833 &  x836 &  x845 &  x848 &  x851 &  x854 &  x860 &  x869 &  x878 &  x881 &  x884 &  x887 &  x890 &  x899 &  x904 &  x911 &  x914 &  x917 &  x923 &  x938 &  x940 &  x944 &  x950 &  x956 &  x965 &  x968 &  x971 &  x979 &  x980 &  x983 &  x986 &  x992 &  x1007 &  x1013 &  x1019 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1085 &  x1097 &  x1103 &  x1106 &  x1112 &  x1115;
assign c190 =  x2 &  x8 &  x14 &  x17 &  x23 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x230 &  x233 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x341 &  x344 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x389 &  x392 &  x395 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x434 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x506 &  x509 &  x512 &  x515 &  x518 &  x527 &  x530 &  x533 &  x536 &  x542 &  x545 &  x551 &  x557 &  x563 &  x566 &  x569 &  x572 &  x574 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x599 &  x602 &  x605 &  x611 &  x613 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x652 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x689 &  x690 &  x691 &  x695 &  x698 &  x701 &  x704 &  x707 &  x713 &  x715 &  x719 &  x722 &  x725 &  x728 &  x730 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x754 &  x755 &  x758 &  x761 &  x764 &  x767 &  x769 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x866 &  x869 &  x871 &  x872 &  x878 &  x881 &  x884 &  x887 &  x893 &  x896 &  x902 &  x905 &  x908 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x977 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1058 &  x1061 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x888;
assign c192 =  x2 &  x5 &  x11 &  x14 &  x17 &  x20 &  x23 &  x38 &  x41 &  x44 &  x50 &  x53 &  x56 &  x65 &  x74 &  x80 &  x83 &  x86 &  x95 &  x98 &  x101 &  x107 &  x116 &  x125 &  x131 &  x134 &  x137 &  x146 &  x149 &  x164 &  x167 &  x173 &  x176 &  x182 &  x185 &  x194 &  x197 &  x200 &  x212 &  x215 &  x227 &  x233 &  x239 &  x245 &  x260 &  x269 &  x278 &  x281 &  x284 &  x293 &  x302 &  x310 &  x320 &  x325 &  x332 &  x338 &  x341 &  x344 &  x362 &  x374 &  x377 &  x380 &  x388 &  x389 &  x395 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x428 &  x440 &  x442 &  x455 &  x476 &  x485 &  x488 &  x494 &  x497 &  x500 &  x503 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x548 &  x551 &  x560 &  x569 &  x575 &  x578 &  x587 &  x590 &  x593 &  x596 &  x605 &  x608 &  x617 &  x623 &  x626 &  x629 &  x635 &  x638 &  x647 &  x656 &  x659 &  x665 &  x668 &  x677 &  x686 &  x695 &  x698 &  x704 &  x707 &  x713 &  x725 &  x734 &  x737 &  x742 &  x745 &  x749 &  x755 &  x764 &  x776 &  x782 &  x784 &  x788 &  x791 &  x794 &  x800 &  x809 &  x824 &  x830 &  x836 &  x839 &  x854 &  x859 &  x866 &  x869 &  x875 &  x878 &  x887 &  x890 &  x896 &  x899 &  x901 &  x908 &  x911 &  x914 &  x917 &  x938 &  x940 &  x941 &  x959 &  x965 &  x968 &  x971 &  x974 &  x979 &  x983 &  x985 &  x992 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1021 &  x1022 &  x1025 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1058 &  x1061 &  x1063 &  x1070 &  x1097 &  x1103 &  x1115 &  x1124 & ~x312 & ~x915 & ~x966;
assign c194 =  x14 &  x17 &  x32 &  x41 &  x47 &  x53 &  x59 &  x70 &  x71 &  x77 &  x83 &  x86 &  x92 &  x95 &  x101 &  x104 &  x107 &  x109 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x148 &  x149 &  x158 &  x161 &  x167 &  x170 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x206 &  x215 &  x218 &  x221 &  x224 &  x230 &  x239 &  x245 &  x248 &  x251 &  x254 &  x257 &  x266 &  x275 &  x278 &  x281 &  x284 &  x290 &  x305 &  x311 &  x317 &  x320 &  x323 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x395 &  x404 &  x407 &  x410 &  x416 &  x422 &  x425 &  x428 &  x430 &  x431 &  x440 &  x449 &  x452 &  x461 &  x472 &  x476 &  x488 &  x494 &  x503 &  x509 &  x511 &  x512 &  x521 &  x524 &  x536 &  x542 &  x545 &  x551 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x584 &  x589 &  x593 &  x596 &  x599 &  x605 &  x614 &  x617 &  x623 &  x628 &  x635 &  x638 &  x641 &  x644 &  x656 &  x659 &  x662 &  x667 &  x668 &  x671 &  x674 &  x677 &  x683 &  x698 &  x701 &  x710 &  x713 &  x722 &  x725 &  x728 &  x737 &  x746 &  x748 &  x749 &  x752 &  x755 &  x758 &  x761 &  x770 &  x773 &  x776 &  x779 &  x782 &  x788 &  x791 &  x794 &  x806 &  x809 &  x818 &  x821 &  x826 &  x830 &  x833 &  x842 &  x845 &  x848 &  x854 &  x857 &  x860 &  x866 &  x869 &  x872 &  x875 &  x893 &  x905 &  x911 &  x917 &  x920 &  x929 &  x932 &  x935 &  x938 &  x944 &  x950 &  x956 &  x959 &  x962 &  x965 &  x971 &  x983 &  x992 &  x995 &  x998 &  x1000 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1025 &  x1031 &  x1034 &  x1039 &  x1040 &  x1043 &  x1045 &  x1058 &  x1067 &  x1073 &  x1078 &  x1082 &  x1084 &  x1085 &  x1088 &  x1091 &  x1103 &  x1105 &  x1109 &  x1115 &  x1117 &  x1127 & ~x501 & ~x639 & ~x741 & ~x897 & ~x975 & ~x1014 & ~x1053;
assign c196 =  x2 &  x5 &  x20 &  x23 &  x32 &  x38 &  x41 &  x43 &  x59 &  x62 &  x68 &  x71 &  x74 &  x77 &  x82 &  x83 &  x89 &  x92 &  x95 &  x98 &  x101 &  x107 &  x110 &  x119 &  x122 &  x131 &  x134 &  x140 &  x143 &  x146 &  x152 &  x155 &  x160 &  x164 &  x166 &  x176 &  x185 &  x191 &  x194 &  x197 &  x206 &  x215 &  x218 &  x227 &  x236 &  x238 &  x245 &  x254 &  x269 &  x274 &  x283 &  x284 &  x290 &  x299 &  x305 &  x308 &  x311 &  x313 &  x314 &  x317 &  x322 &  x323 &  x329 &  x341 &  x347 &  x352 &  x353 &  x368 &  x371 &  x374 &  x380 &  x386 &  x389 &  x392 &  x398 &  x404 &  x407 &  x416 &  x422 &  x434 &  x437 &  x443 &  x452 &  x455 &  x458 &  x461 &  x473 &  x478 &  x482 &  x488 &  x500 &  x503 &  x511 &  x512 &  x515 &  x518 &  x524 &  x527 &  x530 &  x542 &  x557 &  x560 &  x563 &  x566 &  x572 &  x575 &  x578 &  x584 &  x587 &  x590 &  x602 &  x605 &  x617 &  x620 &  x626 &  x635 &  x641 &  x644 &  x659 &  x662 &  x665 &  x674 &  x686 &  x692 &  x695 &  x707 &  x710 &  x719 &  x731 &  x743 &  x752 &  x758 &  x767 &  x776 &  x782 &  x785 &  x788 &  x791 &  x794 &  x803 &  x812 &  x818 &  x833 &  x836 &  x845 &  x851 &  x860 &  x866 &  x875 &  x878 &  x884 &  x893 &  x896 &  x899 &  x902 &  x911 &  x917 &  x920 &  x922 &  x926 &  x932 &  x938 &  x944 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x967 &  x971 &  x974 &  x980 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1006 &  x1007 &  x1010 &  x1016 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1055 &  x1058 &  x1073 &  x1076 &  x1085 &  x1094 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 & ~x186;
assign c198 =  x2 &  x5 &  x11 &  x14 &  x17 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x65 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x92 &  x101 &  x104 &  x107 &  x110 &  x116 &  x119 &  x125 &  x134 &  x140 &  x143 &  x152 &  x155 &  x161 &  x167 &  x173 &  x176 &  x179 &  x181 &  x182 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x206 &  x209 &  x212 &  x221 &  x224 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x269 &  x272 &  x275 &  x281 &  x284 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x326 &  x329 &  x332 &  x341 &  x350 &  x353 &  x356 &  x365 &  x368 &  x371 &  x374 &  x380 &  x383 &  x389 &  x395 &  x398 &  x401 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x431 &  x433 &  x434 &  x440 &  x443 &  x446 &  x452 &  x458 &  x461 &  x467 &  x470 &  x472 &  x473 &  x476 &  x479 &  x482 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x509 &  x511 &  x512 &  x515 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x593 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x626 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x677 &  x683 &  x686 &  x689 &  x695 &  x698 &  x701 &  x707 &  x710 &  x713 &  x716 &  x719 &  x725 &  x728 &  x734 &  x740 &  x747 &  x748 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x776 &  x779 &  x782 &  x785 &  x786 &  x787 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x826 &  x830 &  x833 &  x836 &  x839 &  x842 &  x844 &  x845 &  x854 &  x857 &  x860 &  x863 &  x865 &  x869 &  x872 &  x875 &  x878 &  x881 &  x883 &  x884 &  x887 &  x893 &  x899 &  x902 &  x904 &  x905 &  x908 &  x911 &  x914 &  x917 &  x922 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x950 &  x953 &  x956 &  x962 &  x965 &  x968 &  x971 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1010 &  x1012 &  x1019 &  x1022 &  x1025 &  x1031 &  x1037 &  x1040 &  x1043 &  x1045 &  x1049 &  x1055 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1084 &  x1085 &  x1088 &  x1090 &  x1091 &  x1094 &  x1097 &  x1103 &  x1115 &  x1121 &  x1127 &  x1129 & ~x663 & ~x741 & ~x780 & ~x858;
assign c1100 =  x2 &  x5 &  x8 &  x17 &  x20 &  x29 &  x32 &  x35 &  x38 &  x41 &  x50 &  x56 &  x59 &  x62 &  x68 &  x71 &  x77 &  x80 &  x82 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x113 &  x116 &  x119 &  x121 &  x122 &  x125 &  x128 &  x137 &  x149 &  x152 &  x160 &  x164 &  x167 &  x170 &  x176 &  x179 &  x182 &  x188 &  x191 &  x194 &  x197 &  x203 &  x215 &  x230 &  x236 &  x238 &  x239 &  x242 &  x245 &  x248 &  x260 &  x269 &  x274 &  x277 &  x278 &  x281 &  x284 &  x290 &  x293 &  x296 &  x308 &  x317 &  x320 &  x323 &  x335 &  x341 &  x344 &  x347 &  x350 &  x355 &  x356 &  x359 &  x368 &  x374 &  x383 &  x386 &  x389 &  x392 &  x394 &  x395 &  x397 &  x401 &  x404 &  x407 &  x410 &  x416 &  x419 &  x425 &  x436 &  x437 &  x440 &  x443 &  x449 &  x452 &  x455 &  x464 &  x467 &  x470 &  x473 &  x476 &  x482 &  x485 &  x488 &  x491 &  x500 &  x503 &  x506 &  x509 &  x512 &  x514 &  x515 &  x521 &  x527 &  x533 &  x542 &  x545 &  x551 &  x553 &  x554 &  x563 &  x569 &  x572 &  x578 &  x581 &  x584 &  x587 &  x592 &  x605 &  x608 &  x611 &  x617 &  x623 &  x629 &  x631 &  x632 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x671 &  x674 &  x677 &  x680 &  x686 &  x692 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x722 &  x725 &  x728 &  x731 &  x743 &  x746 &  x758 &  x766 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x812 &  x818 &  x821 &  x827 &  x830 &  x833 &  x836 &  x839 &  x845 &  x848 &  x851 &  x857 &  x863 &  x869 &  x875 &  x878 &  x884 &  x899 &  x905 &  x908 &  x911 &  x917 &  x920 &  x926 &  x932 &  x947 &  x950 &  x953 &  x956 &  x968 &  x971 &  x980 &  x992 &  x995 &  x998 &  x1013 &  x1016 &  x1025 &  x1028 &  x1034 &  x1055 &  x1058 &  x1061 &  x1070 &  x1073 &  x1079 &  x1088 &  x1091 &  x1094 &  x1097 &  x1106 &  x1112 &  x1115 &  x1130 & ~x114 & ~x303 & ~x366 & ~x444 & ~x624 & ~x663 & ~x741 & ~x780 & ~x819;
assign c1102 =  x2 &  x8 &  x11 &  x17 &  x23 &  x26 &  x29 &  x41 &  x47 &  x50 &  x53 &  x65 &  x74 &  x80 &  x95 &  x101 &  x104 &  x110 &  x116 &  x125 &  x128 &  x140 &  x146 &  x155 &  x158 &  x161 &  x167 &  x173 &  x176 &  x188 &  x200 &  x206 &  x209 &  x212 &  x221 &  x227 &  x230 &  x236 &  x239 &  x248 &  x254 &  x257 &  x266 &  x272 &  x275 &  x278 &  x281 &  x287 &  x290 &  x299 &  x308 &  x317 &  x323 &  x335 &  x344 &  x347 &  x350 &  x362 &  x371 &  x380 &  x383 &  x398 &  x401 &  x404 &  x407 &  x422 &  x428 &  x434 &  x452 &  x454 &  x458 &  x464 &  x470 &  x476 &  x482 &  x488 &  x491 &  x493 &  x494 &  x497 &  x503 &  x512 &  x514 &  x515 &  x524 &  x527 &  x530 &  x532 &  x533 &  x536 &  x539 &  x548 &  x551 &  x553 &  x557 &  x560 &  x571 &  x572 &  x575 &  x587 &  x590 &  x593 &  x602 &  x605 &  x608 &  x610 &  x616 &  x617 &  x623 &  x626 &  x635 &  x652 &  x668 &  x671 &  x677 &  x680 &  x686 &  x689 &  x691 &  x692 &  x698 &  x704 &  x707 &  x710 &  x713 &  x715 &  x719 &  x725 &  x728 &  x730 &  x734 &  x743 &  x749 &  x755 &  x758 &  x761 &  x770 &  x772 &  x779 &  x782 &  x791 &  x794 &  x803 &  x806 &  x809 &  x812 &  x818 &  x827 &  x836 &  x851 &  x857 &  x887 &  x890 &  x899 &  x905 &  x908 &  x923 &  x938 &  x950 &  x956 &  x959 &  x962 &  x980 &  x983 &  x992 &  x995 &  x1010 &  x1016 &  x1019 &  x1025 &  x1031 &  x1034 &  x1040 &  x1046 &  x1055 &  x1058 &  x1064 &  x1070 &  x1076 &  x1079 &  x1085 &  x1091 &  x1094 &  x1112 &  x1115 &  x1127 &  x1130 & ~x45 & ~x627 & ~x666 & ~x903;
assign c1104 =  x8 &  x17 &  x20 &  x29 &  x32 &  x35 &  x38 &  x44 &  x47 &  x50 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x82 &  x83 &  x86 &  x89 &  x98 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x125 &  x131 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x155 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x227 &  x230 &  x233 &  x238 &  x239 &  x257 &  x260 &  x263 &  x266 &  x272 &  x275 &  x277 &  x278 &  x281 &  x284 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x316 &  x317 &  x323 &  x326 &  x329 &  x335 &  x338 &  x341 &  x350 &  x353 &  x359 &  x362 &  x365 &  x371 &  x383 &  x386 &  x389 &  x394 &  x404 &  x410 &  x413 &  x419 &  x422 &  x425 &  x428 &  x434 &  x436 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x470 &  x475 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x503 &  x506 &  x512 &  x514 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x545 &  x548 &  x551 &  x553 &  x554 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x605 &  x608 &  x614 &  x616 &  x617 &  x623 &  x626 &  x632 &  x638 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x668 &  x671 &  x674 &  x680 &  x683 &  x689 &  x692 &  x698 &  x707 &  x710 &  x713 &  x716 &  x722 &  x731 &  x737 &  x740 &  x746 &  x749 &  x752 &  x755 &  x761 &  x764 &  x767 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x803 &  x806 &  x815 &  x821 &  x827 &  x836 &  x842 &  x845 &  x848 &  x851 &  x860 &  x869 &  x872 &  x881 &  x884 &  x887 &  x890 &  x893 &  x902 &  x905 &  x908 &  x917 &  x926 &  x929 &  x938 &  x941 &  x944 &  x953 &  x959 &  x965 &  x968 &  x974 &  x977 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1055 &  x1058 &  x1061 &  x1067 &  x1070 &  x1073 &  x1076 &  x1088 &  x1091 &  x1094 &  x1103 &  x1109 &  x1115 &  x1121 &  x1127 & ~x444 & ~x447 & ~x483 & ~x525 & ~x546 & ~x663 & ~x822 & ~x861 & ~x900 & ~x939 & ~x978;
assign c1106 =  x2 &  x5 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x328 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x367 &  x368 &  x370 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x893 &  x896 &  x899 &  x901 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x940 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x3 & ~x159 & ~x606 & ~x654 & ~x693 & ~x732 & ~x733;
assign c1108 =  x2 &  x14 &  x20 &  x23 &  x26 &  x29 &  x35 &  x38 &  x41 &  x44 &  x50 &  x53 &  x56 &  x62 &  x65 &  x77 &  x83 &  x89 &  x101 &  x104 &  x107 &  x110 &  x116 &  x122 &  x137 &  x140 &  x143 &  x152 &  x155 &  x160 &  x167 &  x179 &  x182 &  x188 &  x191 &  x194 &  x200 &  x206 &  x209 &  x218 &  x221 &  x230 &  x235 &  x251 &  x254 &  x260 &  x266 &  x269 &  x275 &  x277 &  x278 &  x281 &  x284 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x316 &  x317 &  x323 &  x326 &  x332 &  x335 &  x341 &  x344 &  x353 &  x355 &  x356 &  x371 &  x374 &  x380 &  x398 &  x401 &  x413 &  x419 &  x422 &  x425 &  x436 &  x440 &  x449 &  x452 &  x455 &  x458 &  x467 &  x473 &  x475 &  x482 &  x488 &  x491 &  x494 &  x506 &  x509 &  x512 &  x514 &  x524 &  x533 &  x539 &  x542 &  x545 &  x551 &  x554 &  x566 &  x569 &  x572 &  x575 &  x581 &  x587 &  x590 &  x592 &  x593 &  x602 &  x605 &  x611 &  x626 &  x629 &  x635 &  x641 &  x665 &  x674 &  x686 &  x688 &  x695 &  x704 &  x707 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x748 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x773 &  x779 &  x797 &  x800 &  x812 &  x818 &  x821 &  x824 &  x833 &  x836 &  x839 &  x860 &  x872 &  x875 &  x878 &  x881 &  x890 &  x896 &  x899 &  x914 &  x920 &  x929 &  x932 &  x935 &  x941 &  x947 &  x950 &  x956 &  x959 &  x983 &  x989 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1022 &  x1034 &  x1046 &  x1049 &  x1055 &  x1067 &  x1079 &  x1085 &  x1091 &  x1097 &  x1121 &  x1127 & ~x207 & ~x303 & ~x366 & ~x405 & ~x507 & ~x624 & ~x663 & ~x702 & ~x741 & ~x951;
assign c1110 =  x2 &  x5 &  x8 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x41 &  x44 &  x47 &  x50 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x89 &  x92 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x122 &  x125 &  x128 &  x134 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x185 &  x191 &  x197 &  x200 &  x203 &  x206 &  x215 &  x218 &  x224 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x256 &  x257 &  x260 &  x263 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x295 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x326 &  x329 &  x332 &  x334 &  x335 &  x338 &  x347 &  x353 &  x356 &  x358 &  x359 &  x362 &  x365 &  x368 &  x371 &  x373 &  x377 &  x380 &  x383 &  x386 &  x389 &  x395 &  x398 &  x401 &  x407 &  x410 &  x412 &  x413 &  x422 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x463 &  x464 &  x470 &  x473 &  x479 &  x488 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x545 &  x548 &  x551 &  x554 &  x557 &  x569 &  x572 &  x578 &  x581 &  x587 &  x590 &  x593 &  x596 &  x599 &  x601 &  x602 &  x605 &  x608 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x668 &  x674 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x725 &  x728 &  x731 &  x734 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x773 &  x785 &  x788 &  x794 &  x800 &  x803 &  x806 &  x809 &  x815 &  x818 &  x821 &  x823 &  x827 &  x829 &  x830 &  x833 &  x836 &  x842 &  x845 &  x848 &  x851 &  x857 &  x862 &  x863 &  x868 &  x869 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x901 &  x902 &  x905 &  x907 &  x908 &  x911 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x940 &  x944 &  x946 &  x947 &  x950 &  x953 &  x956 &  x962 &  x968 &  x971 &  x974 &  x979 &  x980 &  x983 &  x985 &  x986 &  x989 &  x992 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1018 &  x1019 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1058 &  x1063 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1121 &  x1130 & ~x429 & ~x468 & ~x1083;
assign c1112 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x29 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x122 &  x128 &  x137 &  x140 &  x143 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x209 &  x215 &  x218 &  x221 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x254 &  x257 &  x260 &  x263 &  x269 &  x275 &  x277 &  x278 &  x287 &  x290 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x316 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x397 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x436 &  x437 &  x440 &  x443 &  x449 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x475 &  x476 &  x479 &  x482 &  x485 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x553 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x592 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x617 &  x620 &  x623 &  x626 &  x629 &  x631 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x659 &  x662 &  x665 &  x668 &  x670 &  x671 &  x674 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x709 &  x710 &  x713 &  x715 &  x716 &  x722 &  x725 &  x727 &  x728 &  x731 &  x737 &  x740 &  x743 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x766 &  x767 &  x770 &  x773 &  x776 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x836 &  x842 &  x845 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x914 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x977 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x309 & ~x387 & ~x388 & ~x426 & ~x585 & ~x624 & ~x663 & ~x702 & ~x741;
assign c1114 =  x2 &  x8 &  x23 &  x26 &  x35 &  x38 &  x44 &  x50 &  x53 &  x56 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x104 &  x107 &  x113 &  x116 &  x119 &  x122 &  x131 &  x134 &  x137 &  x140 &  x146 &  x149 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x209 &  x218 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x275 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x308 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x350 &  x353 &  x356 &  x362 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x389 &  x392 &  x398 &  x404 &  x407 &  x419 &  x422 &  x425 &  x431 &  x434 &  x437 &  x440 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x479 &  x488 &  x491 &  x494 &  x506 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x548 &  x551 &  x554 &  x563 &  x566 &  x569 &  x572 &  x578 &  x584 &  x587 &  x590 &  x593 &  x601 &  x614 &  x617 &  x623 &  x629 &  x635 &  x638 &  x640 &  x641 &  x644 &  x647 &  x650 &  x656 &  x662 &  x665 &  x668 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x703 &  x710 &  x713 &  x734 &  x737 &  x740 &  x758 &  x767 &  x770 &  x773 &  x776 &  x779 &  x781 &  x782 &  x785 &  x788 &  x791 &  x794 &  x809 &  x812 &  x818 &  x821 &  x823 &  x827 &  x830 &  x842 &  x848 &  x851 &  x854 &  x857 &  x859 &  x860 &  x866 &  x869 &  x872 &  x875 &  x881 &  x887 &  x890 &  x896 &  x898 &  x902 &  x905 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x941 &  x944 &  x947 &  x950 &  x956 &  x959 &  x965 &  x968 &  x974 &  x976 &  x979 &  x980 &  x983 &  x986 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1018 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1067 &  x1070 &  x1073 &  x1079 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x198 & ~x276 & ~x315 & ~x351 & ~x390 & ~x399 & ~x438 & ~x471 & ~x477 & ~x510 & ~x549 & ~x954 & ~x993 & ~x1032;
assign c1116 =  x2 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x65 &  x68 &  x71 &  x74 &  x77 &  x86 &  x89 &  x92 &  x95 &  x101 &  x104 &  x107 &  x110 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x197 &  x203 &  x212 &  x215 &  x218 &  x230 &  x236 &  x239 &  x245 &  x248 &  x251 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x308 &  x311 &  x314 &  x317 &  x320 &  x326 &  x329 &  x332 &  x335 &  x338 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x389 &  x392 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x419 &  x422 &  x428 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x491 &  x494 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x626 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x713 &  x719 &  x722 &  x725 &  x731 &  x734 &  x737 &  x742 &  x743 &  x749 &  x752 &  x755 &  x758 &  x764 &  x767 &  x770 &  x773 &  x779 &  x781 &  x782 &  x785 &  x788 &  x791 &  x794 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x820 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x845 &  x851 &  x854 &  x857 &  x859 &  x860 &  x863 &  x866 &  x869 &  x875 &  x878 &  x884 &  x896 &  x899 &  x902 &  x905 &  x908 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x937 &  x938 &  x941 &  x944 &  x947 &  x956 &  x962 &  x965 &  x968 &  x971 &  x974 &  x980 &  x983 &  x992 &  x995 &  x1001 &  x1018 &  x1019 &  x1025 &  x1028 &  x1031 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1057 &  x1060 &  x1061 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1097 &  x1099 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 &  x1130 & ~x315 & ~x354 & ~x432 & ~x555 & ~x840 & ~x990 & ~x1029 & ~x1107;
assign c1118 =  x2 &  x5 &  x8 &  x11 &  x14 &  x23 &  x26 &  x38 &  x47 &  x53 &  x56 &  x62 &  x65 &  x68 &  x83 &  x89 &  x92 &  x95 &  x104 &  x113 &  x116 &  x122 &  x125 &  x131 &  x140 &  x143 &  x152 &  x158 &  x167 &  x173 &  x176 &  x188 &  x191 &  x197 &  x200 &  x203 &  x212 &  x215 &  x218 &  x221 &  x227 &  x230 &  x233 &  x236 &  x245 &  x250 &  x254 &  x257 &  x272 &  x281 &  x293 &  x296 &  x299 &  x305 &  x323 &  x326 &  x328 &  x329 &  x335 &  x341 &  x347 &  x353 &  x356 &  x365 &  x367 &  x368 &  x371 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x410 &  x416 &  x422 &  x428 &  x431 &  x449 &  x455 &  x461 &  x467 &  x476 &  x479 &  x482 &  x485 &  x500 &  x512 &  x515 &  x530 &  x536 &  x539 &  x545 &  x548 &  x560 &  x563 &  x581 &  x584 &  x587 &  x590 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x620 &  x635 &  x650 &  x653 &  x659 &  x662 &  x664 &  x665 &  x668 &  x671 &  x674 &  x677 &  x686 &  x695 &  x698 &  x707 &  x710 &  x719 &  x722 &  x731 &  x737 &  x740 &  x742 &  x743 &  x746 &  x749 &  x755 &  x758 &  x761 &  x767 &  x770 &  x773 &  x781 &  x784 &  x788 &  x797 &  x800 &  x806 &  x809 &  x812 &  x818 &  x827 &  x833 &  x836 &  x839 &  x860 &  x863 &  x866 &  x869 &  x878 &  x881 &  x884 &  x887 &  x896 &  x901 &  x902 &  x905 &  x914 &  x920 &  x929 &  x938 &  x941 &  x950 &  x953 &  x956 &  x965 &  x968 &  x977 &  x983 &  x995 &  x1001 &  x1004 &  x1010 &  x1028 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1073 &  x1082 &  x1085 &  x1094 &  x1097 &  x1103 &  x1112 &  x1115 &  x1121 &  x1124 & ~x315 & ~x435 & ~x474 & ~x630 & ~x694;
assign c1120 =  x38 &  x44 &  x47 &  x59 &  x62 &  x68 &  x71 &  x74 &  x80 &  x95 &  x98 &  x101 &  x104 &  x116 &  x119 &  x125 &  x140 &  x143 &  x149 &  x155 &  x161 &  x173 &  x182 &  x185 &  x188 &  x194 &  x200 &  x206 &  x212 &  x218 &  x227 &  x248 &  x251 &  x269 &  x278 &  x281 &  x293 &  x296 &  x299 &  x311 &  x314 &  x317 &  x326 &  x329 &  x332 &  x335 &  x344 &  x347 &  x368 &  x374 &  x383 &  x386 &  x392 &  x398 &  x401 &  x407 &  x416 &  x419 &  x428 &  x437 &  x452 &  x458 &  x470 &  x472 &  x485 &  x488 &  x491 &  x497 &  x503 &  x515 &  x524 &  x527 &  x530 &  x539 &  x548 &  x569 &  x572 &  x587 &  x596 &  x605 &  x608 &  x617 &  x623 &  x632 &  x638 &  x641 &  x653 &  x662 &  x683 &  x686 &  x695 &  x698 &  x716 &  x719 &  x722 &  x728 &  x731 &  x758 &  x767 &  x773 &  x776 &  x797 &  x809 &  x827 &  x836 &  x851 &  x857 &  x863 &  x869 &  x890 &  x905 &  x911 &  x920 &  x929 &  x935 &  x941 &  x950 &  x953 &  x961 &  x974 &  x986 &  x995 &  x998 &  x1004 &  x1016 &  x1022 &  x1025 &  x1037 &  x1046 &  x1049 &  x1061 &  x1076 &  x1078 &  x1097 &  x1100 &  x1112 &  x1124 & ~x72 & ~x177 & ~x495 & ~x678 & ~x756 & ~x897 & ~x936 & ~x975 & ~x1017 & ~x1053 & ~x1056 & ~x1095;
assign c1122 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x625 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x667 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x826 &  x827 &  x829 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x863 &  x865 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x901 &  x902 &  x904 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x357 & ~x534 & ~x558 & ~x597 & ~x636;
assign c1124 =  x8 &  x14 &  x17 &  x20 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x56 &  x62 &  x71 &  x74 &  x77 &  x80 &  x89 &  x92 &  x101 &  x107 &  x113 &  x116 &  x122 &  x125 &  x128 &  x131 &  x137 &  x143 &  x146 &  x149 &  x152 &  x155 &  x161 &  x164 &  x167 &  x170 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x212 &  x218 &  x221 &  x230 &  x236 &  x239 &  x242 &  x245 &  x260 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x296 &  x299 &  x305 &  x311 &  x314 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x362 &  x365 &  x371 &  x374 &  x377 &  x383 &  x389 &  x392 &  x398 &  x403 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x434 &  x440 &  x449 &  x452 &  x458 &  x461 &  x464 &  x467 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x521 &  x524 &  x530 &  x533 &  x536 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x575 &  x578 &  x581 &  x584 &  x587 &  x593 &  x596 &  x599 &  x605 &  x608 &  x611 &  x614 &  x626 &  x629 &  x632 &  x641 &  x644 &  x647 &  x656 &  x659 &  x662 &  x665 &  x671 &  x674 &  x677 &  x683 &  x686 &  x689 &  x695 &  x698 &  x704 &  x707 &  x710 &  x716 &  x719 &  x722 &  x725 &  x731 &  x734 &  x737 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x833 &  x836 &  x842 &  x848 &  x857 &  x869 &  x872 &  x878 &  x884 &  x887 &  x890 &  x896 &  x899 &  x902 &  x905 &  x908 &  x914 &  x917 &  x920 &  x932 &  x935 &  x941 &  x947 &  x950 &  x953 &  x959 &  x965 &  x971 &  x974 &  x977 &  x979 &  x980 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1018 &  x1019 &  x1022 &  x1028 &  x1034 &  x1043 &  x1052 &  x1055 &  x1058 &  x1061 &  x1070 &  x1073 &  x1076 &  x1079 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1130 & ~x555 & ~x810 & ~x811 & ~x849 & ~x912 & ~x960 & ~x966 & ~x990 & ~x999 & ~x1005;
assign c1126 =  x2 &  x5 &  x11 &  x14 &  x17 &  x20 &  x29 &  x32 &  x38 &  x56 &  x59 &  x62 &  x65 &  x74 &  x80 &  x82 &  x98 &  x101 &  x104 &  x107 &  x110 &  x119 &  x122 &  x128 &  x140 &  x146 &  x149 &  x158 &  x164 &  x167 &  x170 &  x173 &  x182 &  x188 &  x200 &  x206 &  x218 &  x221 &  x236 &  x239 &  x242 &  x245 &  x254 &  x257 &  x269 &  x275 &  x278 &  x281 &  x287 &  x296 &  x308 &  x311 &  x317 &  x323 &  x326 &  x332 &  x341 &  x344 &  x347 &  x350 &  x359 &  x361 &  x362 &  x374 &  x380 &  x386 &  x389 &  x392 &  x398 &  x401 &  x416 &  x419 &  x428 &  x431 &  x433 &  x434 &  x440 &  x452 &  x458 &  x461 &  x467 &  x472 &  x509 &  x512 &  x518 &  x521 &  x524 &  x533 &  x539 &  x542 &  x545 &  x548 &  x557 &  x569 &  x572 &  x578 &  x581 &  x587 &  x592 &  x599 &  x602 &  x608 &  x617 &  x620 &  x623 &  x631 &  x632 &  x638 &  x641 &  x644 &  x650 &  x659 &  x668 &  x671 &  x677 &  x692 &  x698 &  x707 &  x710 &  x713 &  x719 &  x728 &  x749 &  x752 &  x760 &  x761 &  x764 &  x767 &  x776 &  x785 &  x788 &  x799 &  x800 &  x808 &  x809 &  x824 &  x827 &  x836 &  x839 &  x845 &  x847 &  x851 &  x854 &  x860 &  x863 &  x872 &  x875 &  x877 &  x878 &  x887 &  x890 &  x893 &  x905 &  x908 &  x915 &  x916 &  x917 &  x920 &  x926 &  x929 &  x935 &  x941 &  x944 &  x947 &  x950 &  x955 &  x959 &  x968 &  x971 &  x974 &  x977 &  x983 &  x998 &  x1001 &  x1016 &  x1022 &  x1025 &  x1028 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1070 &  x1073 &  x1079 &  x1085 &  x1100 &  x1103 &  x1112 &  x1121 &  x1124 &  x1130 & ~x702;
assign c1128 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x35 &  x38 &  x41 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x212 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x272 &  x275 &  x278 &  x281 &  x284 &  x289 &  x290 &  x293 &  x296 &  x302 &  x305 &  x308 &  x311 &  x314 &  x323 &  x326 &  x328 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x365 &  x367 &  x368 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x398 &  x401 &  x404 &  x406 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x434 &  x437 &  x440 &  x446 &  x449 &  x452 &  x458 &  x464 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x557 &  x566 &  x569 &  x575 &  x578 &  x581 &  x586 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x625 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x659 &  x662 &  x664 &  x668 &  x671 &  x674 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x706 &  x707 &  x712 &  x713 &  x716 &  x725 &  x728 &  x731 &  x737 &  x740 &  x743 &  x745 &  x749 &  x751 &  x752 &  x755 &  x758 &  x761 &  x767 &  x770 &  x773 &  x779 &  x782 &  x784 &  x785 &  x788 &  x790 &  x791 &  x794 &  x797 &  x803 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x829 &  x830 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x857 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x896 &  x899 &  x905 &  x911 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1100 &  x1103 &  x1112 &  x1124 &  x1127 &  x1130 & ~x321 & ~x660 & ~x699 & ~x738 & ~x777;
assign c1130 =  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x35 &  x38 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x98 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x131 &  x134 &  x140 &  x146 &  x149 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x242 &  x248 &  x251 &  x257 &  x260 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x341 &  x344 &  x353 &  x356 &  x359 &  x362 &  x368 &  x371 &  x374 &  x376 &  x380 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x410 &  x415 &  x416 &  x419 &  x422 &  x425 &  x428 &  x434 &  x443 &  x449 &  x452 &  x454 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x488 &  x493 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x532 &  x536 &  x539 &  x542 &  x545 &  x548 &  x554 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x581 &  x584 &  x587 &  x596 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x626 &  x632 &  x638 &  x644 &  x650 &  x653 &  x656 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x689 &  x692 &  x695 &  x701 &  x710 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x743 &  x749 &  x752 &  x755 &  x758 &  x764 &  x767 &  x770 &  x773 &  x776 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x805 &  x806 &  x809 &  x815 &  x818 &  x821 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x893 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x923 &  x928 &  x929 &  x932 &  x941 &  x944 &  x947 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1084 &  x1085 &  x1088 &  x1097 &  x1100 &  x1103 &  x1115 &  x1118 &  x1121 &  x1123 &  x1124 &  x1127 &  x1130 & ~x411 & ~x507 & ~x546 & ~x606 & ~x645 & ~x663 & ~x741 & ~x780 & ~x858;
assign c1132 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x188 &  x191 &  x194 &  x197 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x341 &  x344 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x431 &  x437 &  x440 &  x446 &  x449 &  x452 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x339 & ~x363 & ~x378 & ~x379 & ~x402 & ~x417 & ~x418 & ~x456 & ~x457 & ~x495 & ~x496 & ~x519 & ~x558 & ~x636 & ~x702 & ~x741;
assign c1134 =  x2 &  x5 &  x8 &  x11 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x95 &  x98 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x251 &  x253 &  x254 &  x257 &  x263 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x353 &  x356 &  x359 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x389 &  x395 &  x398 &  x401 &  x404 &  x407 &  x409 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x448 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x524 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x593 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x273 & ~x312 & ~x927 & ~x966 & ~x1005 & ~x1030 & ~x1044 & ~x1068 & ~x1071 & ~x1086 & ~x1110;
assign c1136 =  x5 &  x11 &  x14 &  x23 &  x41 &  x44 &  x47 &  x50 &  x53 &  x74 &  x77 &  x80 &  x83 &  x86 &  x95 &  x98 &  x107 &  x113 &  x116 &  x119 &  x152 &  x155 &  x158 &  x164 &  x167 &  x173 &  x176 &  x179 &  x188 &  x191 &  x194 &  x206 &  x209 &  x212 &  x221 &  x224 &  x227 &  x230 &  x248 &  x263 &  x284 &  x287 &  x290 &  x302 &  x317 &  x320 &  x329 &  x338 &  x341 &  x359 &  x362 &  x377 &  x389 &  x394 &  x398 &  x410 &  x413 &  x422 &  x440 &  x449 &  x458 &  x464 &  x467 &  x476 &  x488 &  x500 &  x503 &  x506 &  x515 &  x517 &  x518 &  x530 &  x536 &  x557 &  x581 &  x590 &  x602 &  x623 &  x632 &  x680 &  x707 &  x713 &  x721 &  x731 &  x733 &  x734 &  x737 &  x740 &  x760 &  x767 &  x778 &  x782 &  x799 &  x800 &  x805 &  x806 &  x824 &  x833 &  x836 &  x839 &  x848 &  x851 &  x854 &  x860 &  x869 &  x878 &  x881 &  x883 &  x884 &  x893 &  x896 &  x902 &  x908 &  x916 &  x917 &  x920 &  x928 &  x929 &  x938 &  x965 &  x974 &  x983 &  x989 &  x998 &  x1001 &  x1004 &  x1007 &  x1033 &  x1034 &  x1040 &  x1058 &  x1064 &  x1073 &  x1076 &  x1084 &  x1088 &  x1094 &  x1100 &  x1106 &  x1127 & ~x486 & ~x663 & ~x703 & ~x742 & ~x819 & ~x900 & ~x936;
assign c1138 =  x8 &  x11 &  x14 &  x17 &  x35 &  x41 &  x44 &  x53 &  x62 &  x65 &  x68 &  x83 &  x89 &  x92 &  x101 &  x107 &  x110 &  x122 &  x134 &  x140 &  x146 &  x155 &  x167 &  x176 &  x179 &  x182 &  x188 &  x191 &  x197 &  x200 &  x212 &  x227 &  x230 &  x233 &  x238 &  x239 &  x242 &  x254 &  x260 &  x272 &  x275 &  x277 &  x278 &  x281 &  x290 &  x302 &  x305 &  x308 &  x311 &  x316 &  x323 &  x326 &  x329 &  x338 &  x344 &  x362 &  x365 &  x371 &  x383 &  x389 &  x392 &  x394 &  x401 &  x407 &  x425 &  x431 &  x437 &  x443 &  x452 &  x455 &  x464 &  x467 &  x479 &  x482 &  x503 &  x512 &  x515 &  x533 &  x536 &  x539 &  x548 &  x551 &  x554 &  x557 &  x563 &  x566 &  x572 &  x584 &  x587 &  x590 &  x599 &  x605 &  x614 &  x616 &  x617 &  x623 &  x629 &  x631 &  x632 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x661 &  x662 &  x670 &  x671 &  x674 &  x677 &  x680 &  x689 &  x692 &  x694 &  x695 &  x701 &  x704 &  x709 &  x731 &  x737 &  x740 &  x743 &  x748 &  x749 &  x752 &  x755 &  x761 &  x767 &  x778 &  x782 &  x785 &  x791 &  x794 &  x797 &  x806 &  x809 &  x836 &  x871 &  x875 &  x890 &  x902 &  x904 &  x910 &  x923 &  x929 &  x944 &  x947 &  x949 &  x950 &  x959 &  x962 &  x974 &  x980 &  x983 &  x995 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1031 &  x1034 &  x1040 &  x1046 &  x1049 &  x1052 &  x1058 &  x1067 &  x1070 &  x1079 &  x1091 &  x1100 &  x1118 &  x1121 &  x1124 &  x1130 & ~x303 & ~x405 & ~x444 & ~x741 & ~x780 & ~x858 & ~x897 & ~x936;
assign c1140 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x122 &  x128 &  x137 &  x140 &  x142 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x179 &  x182 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x251 &  x257 &  x266 &  x269 &  x281 &  x284 &  x287 &  x293 &  x299 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x437 &  x440 &  x449 &  x452 &  x455 &  x461 &  x464 &  x467 &  x473 &  x479 &  x485 &  x488 &  x494 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x587 &  x589 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x628 &  x632 &  x638 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x667 &  x668 &  x671 &  x674 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x704 &  x706 &  x707 &  x710 &  x713 &  x715 &  x716 &  x722 &  x734 &  x737 &  x743 &  x749 &  x752 &  x754 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x779 &  x782 &  x785 &  x788 &  x791 &  x792 &  x793 &  x794 &  x797 &  x800 &  x806 &  x809 &  x815 &  x818 &  x821 &  x824 &  x827 &  x832 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x871 &  x872 &  x875 &  x881 &  x884 &  x890 &  x893 &  x896 &  x899 &  x902 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x941 &  x944 &  x947 &  x950 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1027 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x657 & ~x819;
assign c1142 =  x2 &  x5 &  x14 &  x20 &  x26 &  x29 &  x32 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x77 &  x80 &  x86 &  x89 &  x92 &  x95 &  x101 &  x110 &  x122 &  x125 &  x128 &  x134 &  x140 &  x143 &  x146 &  x161 &  x164 &  x170 &  x173 &  x179 &  x182 &  x188 &  x194 &  x197 &  x200 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x230 &  x233 &  x242 &  x248 &  x251 &  x263 &  x266 &  x272 &  x275 &  x284 &  x287 &  x296 &  x317 &  x323 &  x326 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x353 &  x356 &  x362 &  x365 &  x368 &  x371 &  x377 &  x386 &  x389 &  x392 &  x395 &  x401 &  x407 &  x413 &  x416 &  x419 &  x425 &  x428 &  x434 &  x437 &  x446 &  x449 &  x455 &  x461 &  x464 &  x467 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x503 &  x518 &  x524 &  x527 &  x530 &  x533 &  x545 &  x551 &  x563 &  x575 &  x578 &  x581 &  x586 &  x587 &  x590 &  x593 &  x596 &  x602 &  x605 &  x611 &  x614 &  x617 &  x620 &  x623 &  x625 &  x626 &  x632 &  x635 &  x638 &  x641 &  x647 &  x650 &  x653 &  x662 &  x665 &  x667 &  x673 &  x674 &  x686 &  x692 &  x698 &  x701 &  x704 &  x706 &  x712 &  x722 &  x728 &  x731 &  x734 &  x740 &  x746 &  x752 &  x758 &  x761 &  x764 &  x776 &  x779 &  x782 &  x785 &  x787 &  x788 &  x791 &  x794 &  x800 &  x803 &  x815 &  x818 &  x823 &  x826 &  x833 &  x836 &  x839 &  x842 &  x851 &  x854 &  x857 &  x860 &  x866 &  x869 &  x872 &  x875 &  x878 &  x890 &  x893 &  x896 &  x899 &  x902 &  x904 &  x911 &  x914 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x941 &  x950 &  x953 &  x956 &  x962 &  x965 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x995 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1067 &  x1070 &  x1076 &  x1082 &  x1088 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1130 & ~x399 & ~x702 & ~x741 & ~x858;
assign c1144 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x44 &  x47 &  x50 &  x56 &  x65 &  x68 &  x74 &  x77 &  x80 &  x82 &  x86 &  x89 &  x92 &  x95 &  x101 &  x104 &  x107 &  x110 &  x119 &  x121 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x152 &  x155 &  x160 &  x164 &  x170 &  x173 &  x179 &  x182 &  x188 &  x191 &  x194 &  x199 &  x200 &  x203 &  x206 &  x209 &  x215 &  x221 &  x230 &  x233 &  x236 &  x238 &  x242 &  x245 &  x248 &  x251 &  x260 &  x272 &  x275 &  x277 &  x278 &  x284 &  x293 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x316 &  x317 &  x323 &  x326 &  x329 &  x335 &  x338 &  x341 &  x344 &  x350 &  x353 &  x355 &  x356 &  x359 &  x362 &  x365 &  x374 &  x380 &  x383 &  x386 &  x389 &  x392 &  x394 &  x395 &  x397 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x428 &  x431 &  x436 &  x440 &  x443 &  x452 &  x455 &  x458 &  x464 &  x470 &  x473 &  x475 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x503 &  x512 &  x514 &  x515 &  x518 &  x524 &  x527 &  x530 &  x532 &  x533 &  x539 &  x542 &  x545 &  x551 &  x553 &  x554 &  x557 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x590 &  x592 &  x593 &  x596 &  x598 &  x599 &  x608 &  x610 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x631 &  x632 &  x635 &  x637 &  x638 &  x641 &  x643 &  x650 &  x653 &  x659 &  x662 &  x665 &  x668 &  x670 &  x671 &  x677 &  x680 &  x686 &  x688 &  x692 &  x701 &  x704 &  x707 &  x709 &  x710 &  x713 &  x715 &  x719 &  x725 &  x728 &  x731 &  x734 &  x743 &  x746 &  x748 &  x749 &  x752 &  x754 &  x755 &  x758 &  x766 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x793 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x815 &  x821 &  x824 &  x827 &  x830 &  x832 &  x833 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x902 &  x905 &  x908 &  x911 &  x917 &  x923 &  x926 &  x929 &  x932 &  x938 &  x947 &  x953 &  x956 &  x959 &  x965 &  x968 &  x971 &  x977 &  x980 &  x983 &  x986 &  x995 &  x1004 &  x1007 &  x1010 &  x1013 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1055 &  x1058 &  x1061 &  x1067 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x483 & ~x546 & ~x585 & ~x624 & ~x741 & ~x780;
assign c1146 =  x2 &  x8 &  x14 &  x17 &  x26 &  x35 &  x38 &  x50 &  x59 &  x80 &  x89 &  x91 &  x92 &  x95 &  x104 &  x116 &  x119 &  x130 &  x143 &  x161 &  x164 &  x173 &  x185 &  x194 &  x197 &  x200 &  x206 &  x236 &  x239 &  x242 &  x248 &  x272 &  x281 &  x284 &  x293 &  x298 &  x305 &  x311 &  x317 &  x320 &  x329 &  x341 &  x350 &  x353 &  x356 &  x362 &  x365 &  x368 &  x374 &  x377 &  x383 &  x386 &  x389 &  x392 &  x407 &  x410 &  x413 &  x416 &  x428 &  x437 &  x440 &  x446 &  x452 &  x476 &  x479 &  x494 &  x500 &  x503 &  x509 &  x521 &  x527 &  x539 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x590 &  x593 &  x602 &  x605 &  x608 &  x611 &  x626 &  x629 &  x632 &  x644 &  x647 &  x653 &  x656 &  x662 &  x671 &  x674 &  x677 &  x680 &  x683 &  x689 &  x695 &  x701 &  x704 &  x710 &  x716 &  x719 &  x731 &  x734 &  x740 &  x746 &  x749 &  x758 &  x761 &  x773 &  x776 &  x785 &  x788 &  x797 &  x800 &  x803 &  x806 &  x815 &  x818 &  x821 &  x823 &  x824 &  x826 &  x827 &  x842 &  x848 &  x854 &  x857 &  x860 &  x862 &  x863 &  x865 &  x872 &  x884 &  x893 &  x896 &  x899 &  x903 &  x904 &  x911 &  x914 &  x926 &  x953 &  x956 &  x962 &  x968 &  x971 &  x974 &  x983 &  x986 &  x988 &  x992 &  x1001 &  x1007 &  x1019 &  x1022 &  x1027 &  x1028 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1066 &  x1073 &  x1085 &  x1088 &  x1091 &  x1094 &  x1103 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 & ~x156 & ~x276;
assign c1148 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x163 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x202 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x241 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x272 &  x275 &  x278 &  x280 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x343 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x761 &  x764 &  x767 &  x770 &  x773 &  x779 &  x782 &  x784 &  x785 &  x788 &  x790 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x827 &  x829 &  x830 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x863 &  x865 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x896 &  x899 &  x901 &  x902 &  x904 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x940 &  x941 &  x943 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x979 &  x980 &  x982 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1018 &  x1019 &  x1021 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x312 & ~x582 & ~x621;
assign c1150 =  x2 &  x5 &  x11 &  x14 &  x17 &  x20 &  x23 &  x32 &  x35 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x62 &  x65 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x92 &  x98 &  x104 &  x107 &  x110 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x137 &  x140 &  x146 &  x149 &  x152 &  x155 &  x158 &  x160 &  x161 &  x164 &  x167 &  x173 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x209 &  x212 &  x215 &  x221 &  x227 &  x235 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x257 &  x260 &  x263 &  x266 &  x269 &  x275 &  x277 &  x284 &  x287 &  x290 &  x293 &  x299 &  x302 &  x308 &  x311 &  x314 &  x316 &  x317 &  x320 &  x323 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x353 &  x355 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x377 &  x383 &  x386 &  x392 &  x394 &  x395 &  x398 &  x410 &  x413 &  x419 &  x422 &  x425 &  x433 &  x434 &  x437 &  x439 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x470 &  x472 &  x478 &  x479 &  x485 &  x491 &  x494 &  x500 &  x503 &  x506 &  x509 &  x511 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x551 &  x554 &  x556 &  x560 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x593 &  x595 &  x596 &  x602 &  x605 &  x611 &  x614 &  x623 &  x626 &  x629 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x671 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x719 &  x722 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x752 &  x761 &  x764 &  x767 &  x770 &  x776 &  x779 &  x782 &  x788 &  x791 &  x794 &  x797 &  x803 &  x806 &  x808 &  x809 &  x818 &  x821 &  x824 &  x827 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x866 &  x869 &  x872 &  x875 &  x878 &  x887 &  x889 &  x890 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x920 &  x922 &  x923 &  x926 &  x928 &  x929 &  x932 &  x935 &  x938 &  x941 &  x947 &  x950 &  x959 &  x962 &  x971 &  x977 &  x983 &  x986 &  x989 &  x992 &  x998 &  x1001 &  x1007 &  x1012 &  x1013 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1046 &  x1049 &  x1051 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1085 &  x1088 &  x1097 &  x1100 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x303 & ~x780 & ~x819;
assign c1152 =  x5 &  x8 &  x14 &  x20 &  x23 &  x26 &  x35 &  x38 &  x50 &  x53 &  x56 &  x62 &  x65 &  x74 &  x83 &  x86 &  x89 &  x92 &  x95 &  x101 &  x104 &  x110 &  x119 &  x122 &  x128 &  x137 &  x146 &  x164 &  x167 &  x170 &  x176 &  x179 &  x185 &  x191 &  x212 &  x227 &  x230 &  x251 &  x254 &  x266 &  x272 &  x275 &  x277 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x305 &  x311 &  x316 &  x317 &  x320 &  x323 &  x329 &  x335 &  x344 &  x350 &  x377 &  x380 &  x383 &  x386 &  x395 &  x404 &  x413 &  x416 &  x422 &  x425 &  x428 &  x433 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x470 &  x473 &  x479 &  x482 &  x500 &  x509 &  x515 &  x518 &  x521 &  x536 &  x545 &  x548 &  x551 &  x553 &  x554 &  x560 &  x566 &  x575 &  x590 &  x593 &  x596 &  x599 &  x602 &  x611 &  x614 &  x617 &  x623 &  x626 &  x631 &  x632 &  x641 &  x644 &  x653 &  x656 &  x659 &  x668 &  x670 &  x671 &  x680 &  x683 &  x695 &  x698 &  x710 &  x719 &  x725 &  x731 &  x737 &  x740 &  x755 &  x758 &  x761 &  x764 &  x773 &  x776 &  x782 &  x785 &  x794 &  x797 &  x803 &  x809 &  x812 &  x818 &  x824 &  x827 &  x836 &  x848 &  x851 &  x857 &  x860 &  x863 &  x866 &  x872 &  x881 &  x896 &  x908 &  x914 &  x920 &  x926 &  x929 &  x935 &  x938 &  x944 &  x947 &  x950 &  x959 &  x962 &  x965 &  x971 &  x980 &  x998 &  x1007 &  x1010 &  x1022 &  x1025 &  x1031 &  x1037 &  x1040 &  x1046 &  x1049 &  x1055 &  x1058 &  x1061 &  x1070 &  x1073 &  x1079 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1112 &  x1121 &  x1124 & ~x381 & ~x387 & ~x388 & ~x420 & ~x504 & ~x585 & ~x663 & ~x741 & ~x780;
assign c1154 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x196 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x235 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x274 &  x278 &  x281 &  x284 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x436 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x467 &  x470 &  x473 &  x475 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x493 &  x494 &  x500 &  x503 &  x506 &  x509 &  x512 &  x514 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x611 &  x614 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x653 &  x662 &  x665 &  x668 &  x671 &  x674 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x803 &  x806 &  x809 &  x812 &  x815 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 &  x1130 & ~x6 & ~x24 & ~x45 & ~x69 & ~x84 & ~x108 & ~x123 & ~x147 & ~x186 & ~x264 & ~x303 & ~x666 & ~x705;
assign c1156 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x667 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x806 &  x809 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x982 &  x983 &  x986 &  x992 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x87 & ~x126 & ~x165 & ~x183 & ~x204 & ~x399 & ~x720 & ~x801 & ~x840 & ~x879 & ~x990 & ~x996 & ~x1029 & ~x1035 & ~x1068;
assign c1158 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x262 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x301 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x326 &  x329 &  x332 &  x335 &  x338 &  x340 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x377 &  x379 &  x380 &  x383 &  x386 &  x392 &  x395 &  x398 &  x404 &  x407 &  x410 &  x413 &  x416 &  x418 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x446 &  x449 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x520 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x553 &  x554 &  x557 &  x559 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x592 &  x596 &  x598 &  x599 &  x602 &  x605 &  x608 &  x610 &  x614 &  x620 &  x623 &  x626 &  x629 &  x631 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x649 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x788 &  x791 &  x794 &  x796 &  x797 &  x800 &  x803 &  x806 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x835 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x866 &  x869 &  x872 &  x875 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x702 & ~x762;
assign c1160 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x47 &  x50 &  x56 &  x62 &  x68 &  x71 &  x74 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x107 &  x113 &  x116 &  x119 &  x125 &  x128 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x298 &  x299 &  x302 &  x305 &  x311 &  x314 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x371 &  x377 &  x380 &  x386 &  x392 &  x395 &  x398 &  x404 &  x413 &  x416 &  x419 &  x422 &  x437 &  x446 &  x449 &  x452 &  x455 &  x458 &  x464 &  x467 &  x470 &  x473 &  x476 &  x482 &  x485 &  x488 &  x494 &  x497 &  x500 &  x503 &  x506 &  x512 &  x518 &  x530 &  x539 &  x545 &  x548 &  x551 &  x563 &  x566 &  x569 &  x572 &  x575 &  x584 &  x587 &  x593 &  x599 &  x602 &  x608 &  x614 &  x623 &  x625 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x647 &  x650 &  x656 &  x662 &  x665 &  x668 &  x671 &  x674 &  x680 &  x686 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x713 &  x725 &  x728 &  x734 &  x737 &  x743 &  x745 &  x749 &  x752 &  x755 &  x761 &  x764 &  x767 &  x773 &  x776 &  x779 &  x784 &  x785 &  x788 &  x791 &  x794 &  x806 &  x809 &  x812 &  x815 &  x818 &  x823 &  x824 &  x833 &  x836 &  x839 &  x842 &  x845 &  x851 &  x857 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x890 &  x899 &  x901 &  x902 &  x905 &  x908 &  x917 &  x929 &  x935 &  x938 &  x940 &  x941 &  x947 &  x950 &  x953 &  x956 &  x962 &  x968 &  x971 &  x974 &  x980 &  x983 &  x985 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1097 &  x1100 &  x1117 &  x1123 &  x1124 &  x1130 & ~x123 & ~x162 & ~x240 & ~x876;
assign c1162 =  x2 &  x5 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x41 &  x44 &  x47 &  x50 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x116 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x188 &  x191 &  x194 &  x197 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x257 &  x263 &  x266 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x511 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x554 &  x557 &  x563 &  x566 &  x569 &  x572 &  x575 &  x581 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x628 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x656 &  x659 &  x662 &  x665 &  x667 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x758 &  x761 &  x770 &  x773 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x865 &  x866 &  x869 &  x875 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x904 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x9 & ~x48 & ~x87 & ~x126 & ~x204 & ~x639 & ~x657 & ~x678 & ~x717 & ~x780 & ~x795 & ~x819 & ~x858 & ~x897 & ~x936 & ~x1014 & ~x1029 & ~x1053 & ~x1062 & ~x1092 & ~x1101;
assign c1164 =  x2 &  x8 &  x17 &  x19 &  x29 &  x35 &  x41 &  x44 &  x47 &  x50 &  x56 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x122 &  x125 &  x131 &  x134 &  x140 &  x149 &  x161 &  x164 &  x173 &  x176 &  x179 &  x188 &  x191 &  x194 &  x200 &  x203 &  x206 &  x209 &  x212 &  x218 &  x233 &  x236 &  x238 &  x239 &  x242 &  x245 &  x248 &  x263 &  x269 &  x272 &  x277 &  x278 &  x281 &  x290 &  x293 &  x296 &  x314 &  x317 &  x329 &  x332 &  x335 &  x338 &  x344 &  x350 &  x352 &  x353 &  x355 &  x359 &  x365 &  x368 &  x371 &  x383 &  x386 &  x391 &  x392 &  x394 &  x398 &  x407 &  x413 &  x419 &  x428 &  x434 &  x437 &  x452 &  x458 &  x464 &  x467 &  x472 &  x479 &  x482 &  x497 &  x506 &  x511 &  x512 &  x530 &  x533 &  x539 &  x548 &  x551 &  x557 &  x560 &  x563 &  x572 &  x575 &  x578 &  x581 &  x587 &  x590 &  x592 &  x605 &  x608 &  x614 &  x617 &  x620 &  x626 &  x631 &  x638 &  x641 &  x644 &  x650 &  x653 &  x656 &  x662 &  x665 &  x668 &  x671 &  x692 &  x698 &  x701 &  x707 &  x708 &  x709 &  x713 &  x719 &  x725 &  x731 &  x740 &  x748 &  x758 &  x773 &  x776 &  x779 &  x782 &  x785 &  x787 &  x788 &  x794 &  x797 &  x800 &  x815 &  x824 &  x830 &  x836 &  x839 &  x842 &  x845 &  x848 &  x866 &  x869 &  x890 &  x899 &  x902 &  x905 &  x911 &  x914 &  x917 &  x922 &  x926 &  x929 &  x938 &  x941 &  x953 &  x956 &  x959 &  x961 &  x968 &  x974 &  x977 &  x986 &  x989 &  x994 &  x1000 &  x1001 &  x1004 &  x1013 &  x1022 &  x1034 &  x1043 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1091 &  x1097 &  x1100 &  x1103 &  x1112 &  x1130 & ~x381;
assign c1166 =  x5 &  x11 &  x17 &  x26 &  x29 &  x32 &  x35 &  x41 &  x44 &  x47 &  x50 &  x53 &  x59 &  x62 &  x74 &  x80 &  x83 &  x86 &  x89 &  x95 &  x98 &  x104 &  x107 &  x113 &  x116 &  x122 &  x125 &  x128 &  x131 &  x137 &  x140 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x173 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x248 &  x257 &  x260 &  x269 &  x275 &  x278 &  x281 &  x286 &  x290 &  x299 &  x302 &  x305 &  x308 &  x314 &  x317 &  x320 &  x323 &  x326 &  x335 &  x338 &  x344 &  x347 &  x350 &  x353 &  x356 &  x362 &  x371 &  x374 &  x377 &  x386 &  x389 &  x392 &  x395 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x437 &  x443 &  x446 &  x449 &  x452 &  x458 &  x461 &  x470 &  x473 &  x476 &  x479 &  x485 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x512 &  x515 &  x518 &  x521 &  x530 &  x533 &  x539 &  x545 &  x548 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x590 &  x593 &  x596 &  x602 &  x605 &  x608 &  x617 &  x620 &  x623 &  x629 &  x632 &  x641 &  x653 &  x656 &  x659 &  x665 &  x668 &  x677 &  x683 &  x686 &  x692 &  x698 &  x710 &  x716 &  x725 &  x734 &  x737 &  x740 &  x743 &  x745 &  x746 &  x749 &  x752 &  x761 &  x764 &  x770 &  x773 &  x776 &  x782 &  x788 &  x794 &  x803 &  x806 &  x809 &  x812 &  x818 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x845 &  x848 &  x851 &  x854 &  x860 &  x862 &  x863 &  x866 &  x872 &  x878 &  x881 &  x884 &  x887 &  x890 &  x896 &  x899 &  x908 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x941 &  x944 &  x953 &  x956 &  x959 &  x962 &  x968 &  x971 &  x974 &  x977 &  x983 &  x986 &  x989 &  x1001 &  x1010 &  x1016 &  x1019 &  x1025 &  x1028 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x126 & ~x321 & ~x360 & ~x435 & ~x474 & ~x513 & ~x552 & ~x771 & ~x795 & ~x849;
assign c1168 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x34 &  x38 &  x41 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x73 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x188 &  x191 &  x197 &  x200 &  x203 &  x206 &  x209 &  x218 &  x221 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x250 &  x251 &  x260 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x308 &  x311 &  x314 &  x320 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x365 &  x368 &  x380 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x430 &  x431 &  x437 &  x440 &  x443 &  x446 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x469 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x506 &  x508 &  x515 &  x521 &  x524 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x547 &  x548 &  x551 &  x557 &  x560 &  x566 &  x569 &  x572 &  x578 &  x581 &  x586 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x644 &  x647 &  x653 &  x656 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x683 &  x689 &  x692 &  x695 &  x698 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x797 &  x806 &  x809 &  x812 &  x818 &  x821 &  x824 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x851 &  x860 &  x863 &  x866 &  x869 &  x878 &  x881 &  x884 &  x890 &  x893 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x922 &  x926 &  x932 &  x935 &  x938 &  x941 &  x944 &  x950 &  x962 &  x965 &  x967 &  x968 &  x974 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1028 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1121 &  x1124 &  x1130 & ~x543 & ~x681 & ~x717;
assign c1170 =  x8 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x47 &  x50 &  x53 &  x56 &  x62 &  x65 &  x68 &  x71 &  x77 &  x83 &  x86 &  x89 &  x92 &  x98 &  x101 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x146 &  x152 &  x155 &  x158 &  x164 &  x167 &  x170 &  x182 &  x185 &  x188 &  x191 &  x193 &  x200 &  x203 &  x218 &  x221 &  x224 &  x232 &  x239 &  x248 &  x269 &  x272 &  x275 &  x278 &  x284 &  x287 &  x296 &  x302 &  x308 &  x314 &  x323 &  x332 &  x338 &  x341 &  x356 &  x359 &  x362 &  x371 &  x380 &  x386 &  x389 &  x392 &  x401 &  x404 &  x410 &  x416 &  x419 &  x422 &  x434 &  x446 &  x449 &  x452 &  x461 &  x473 &  x476 &  x479 &  x488 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x533 &  x542 &  x545 &  x551 &  x557 &  x560 &  x569 &  x578 &  x581 &  x584 &  x587 &  x590 &  x596 &  x605 &  x608 &  x617 &  x625 &  x632 &  x641 &  x656 &  x664 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x692 &  x695 &  x698 &  x704 &  x707 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x737 &  x740 &  x746 &  x749 &  x755 &  x758 &  x773 &  x776 &  x784 &  x785 &  x788 &  x794 &  x797 &  x809 &  x815 &  x821 &  x823 &  x827 &  x839 &  x845 &  x851 &  x863 &  x872 &  x875 &  x878 &  x884 &  x887 &  x893 &  x899 &  x908 &  x911 &  x917 &  x920 &  x923 &  x929 &  x935 &  x938 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x971 &  x974 &  x977 &  x980 &  x995 &  x998 &  x1013 &  x1022 &  x1028 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1058 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1100 &  x1103 &  x1106 &  x1109 &  x1121 &  x1127 &  x1130 & ~x654 & ~x717 & ~x733 & ~x756 & ~x795 & ~x798 & ~x834 & ~x873 & ~x918 & ~x951;
assign c1172 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x298 &  x299 &  x302 &  x305 &  x308 &  x310 &  x311 &  x314 &  x320 &  x323 &  x326 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x625 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1084 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1123 &  x1124 &  x1127 &  x1130 & ~x273 & ~x576 & ~x615 & ~x654 & ~x693 & ~x717 & ~x732 & ~x756 & ~x771 & ~x798;
assign c1174 =  x5 &  x8 &  x11 &  x20 &  x41 &  x44 &  x47 &  x56 &  x74 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x125 &  x134 &  x137 &  x140 &  x158 &  x161 &  x167 &  x185 &  x188 &  x197 &  x200 &  x209 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x242 &  x245 &  x248 &  x251 &  x257 &  x260 &  x263 &  x266 &  x269 &  x284 &  x290 &  x299 &  x302 &  x305 &  x308 &  x311 &  x317 &  x323 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x356 &  x368 &  x371 &  x383 &  x389 &  x395 &  x407 &  x416 &  x422 &  x425 &  x428 &  x434 &  x440 &  x443 &  x446 &  x455 &  x458 &  x461 &  x464 &  x467 &  x472 &  x479 &  x482 &  x488 &  x491 &  x494 &  x497 &  x503 &  x509 &  x511 &  x512 &  x515 &  x524 &  x530 &  x539 &  x557 &  x569 &  x575 &  x581 &  x584 &  x587 &  x596 &  x605 &  x614 &  x617 &  x620 &  x626 &  x629 &  x635 &  x638 &  x644 &  x671 &  x677 &  x686 &  x689 &  x695 &  x698 &  x704 &  x707 &  x710 &  x713 &  x715 &  x719 &  x728 &  x734 &  x746 &  x749 &  x754 &  x755 &  x761 &  x773 &  x776 &  x782 &  x791 &  x794 &  x800 &  x806 &  x809 &  x824 &  x832 &  x836 &  x842 &  x845 &  x851 &  x854 &  x863 &  x866 &  x871 &  x875 &  x878 &  x881 &  x893 &  x899 &  x902 &  x905 &  x909 &  x911 &  x923 &  x935 &  x938 &  x948 &  x950 &  x959 &  x968 &  x974 &  x977 &  x986 &  x987 &  x988 &  x989 &  x992 &  x1001 &  x1004 &  x1007 &  x1010 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1046 &  x1049 &  x1070 &  x1073 &  x1076 &  x1088 &  x1097 &  x1100 &  x1106 &  x1109 &  x1118 &  x1124 &  x1127 & ~x639 & ~x678 & ~x756 & ~x936 & ~x975;
assign c1176 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x62 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x92 &  x98 &  x101 &  x104 &  x110 &  x113 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x218 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x275 &  x278 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x304 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x343 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x380 &  x382 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x416 &  x419 &  x421 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x460 &  x461 &  x464 &  x467 &  x470 &  x473 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x499 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x538 &  x539 &  x542 &  x545 &  x548 &  x551 &  x557 &  x559 &  x560 &  x566 &  x569 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x611 &  x614 &  x617 &  x623 &  x626 &  x629 &  x632 &  x638 &  x640 &  x641 &  x644 &  x650 &  x653 &  x659 &  x662 &  x665 &  x668 &  x674 &  x677 &  x679 &  x680 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x737 &  x740 &  x743 &  x746 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x781 &  x785 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x820 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x859 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x893 &  x896 &  x898 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x937 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x965 &  x971 &  x974 &  x976 &  x977 &  x980 &  x983 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1018 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1057 &  x1058 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1096 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1121 &  x1127 &  x1130 & ~x354 & ~x393 & ~x432 & ~x549 & ~x588 & ~x954 & ~x955 & ~x993 & ~x1032;
assign c1178 =  x2 &  x5 &  x11 &  x17 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x74 &  x83 &  x86 &  x89 &  x91 &  x92 &  x95 &  x98 &  x101 &  x107 &  x110 &  x113 &  x122 &  x125 &  x128 &  x130 &  x131 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x155 &  x158 &  x161 &  x167 &  x170 &  x173 &  x176 &  x185 &  x191 &  x197 &  x200 &  x212 &  x218 &  x221 &  x224 &  x227 &  x239 &  x245 &  x251 &  x254 &  x257 &  x260 &  x263 &  x269 &  x275 &  x278 &  x284 &  x287 &  x290 &  x293 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x359 &  x365 &  x368 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x404 &  x410 &  x416 &  x419 &  x422 &  x428 &  x431 &  x434 &  x446 &  x449 &  x461 &  x464 &  x467 &  x470 &  x473 &  x479 &  x482 &  x488 &  x494 &  x500 &  x503 &  x506 &  x511 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x542 &  x545 &  x548 &  x551 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x581 &  x587 &  x589 &  x596 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x629 &  x635 &  x638 &  x647 &  x650 &  x653 &  x659 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x698 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x728 &  x731 &  x734 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x776 &  x779 &  x782 &  x788 &  x791 &  x794 &  x797 &  x800 &  x806 &  x809 &  x812 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x860 &  x863 &  x865 &  x866 &  x869 &  x872 &  x875 &  x878 &  x890 &  x893 &  x896 &  x899 &  x902 &  x904 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x956 &  x959 &  x962 &  x968 &  x971 &  x974 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1052 &  x1055 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1082 &  x1088 &  x1090 &  x1091 &  x1094 &  x1103 &  x1106 &  x1109 &  x1112 &  x1121 &  x1124 &  x1127 &  x1130 & ~x0 & ~x126 & ~x165 & ~x204 & ~x639 & ~x678 & ~x756 & ~x834 & ~x936 & ~x1029 & ~x1053 & ~x1092 & ~x1125;
assign c1180 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x29 &  x32 &  x38 &  x41 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x143 &  x146 &  x149 &  x152 &  x158 &  x167 &  x170 &  x173 &  x176 &  x179 &  x188 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x245 &  x254 &  x257 &  x263 &  x266 &  x269 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x328 &  x329 &  x332 &  x335 &  x341 &  x344 &  x350 &  x356 &  x359 &  x362 &  x368 &  x371 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x406 &  x407 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x440 &  x443 &  x445 &  x446 &  x452 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x581 &  x587 &  x593 &  x596 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x623 &  x629 &  x638 &  x641 &  x644 &  x650 &  x653 &  x656 &  x659 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x703 &  x704 &  x707 &  x710 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x742 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x764 &  x767 &  x776 &  x782 &  x785 &  x788 &  x791 &  x794 &  x800 &  x806 &  x809 &  x812 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x839 &  x842 &  x848 &  x851 &  x854 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x890 &  x893 &  x896 &  x899 &  x905 &  x911 &  x914 &  x920 &  x926 &  x932 &  x935 &  x937 &  x938 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x976 &  x977 &  x980 &  x983 &  x989 &  x995 &  x998 &  x1001 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1054 &  x1055 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x399 & ~x438 & ~x477 & ~x516 & ~x555 & ~x594 & ~x1029 & ~x1032 & ~x1068;
assign c1182 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x19 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x47 &  x50 &  x56 &  x58 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x104 &  x107 &  x116 &  x122 &  x125 &  x128 &  x131 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x167 &  x170 &  x182 &  x185 &  x191 &  x194 &  x197 &  x200 &  x203 &  x209 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x278 &  x281 &  x284 &  x287 &  x293 &  x299 &  x302 &  x311 &  x317 &  x320 &  x326 &  x329 &  x335 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x377 &  x380 &  x392 &  x398 &  x404 &  x413 &  x425 &  x428 &  x431 &  x433 &  x434 &  x437 &  x440 &  x446 &  x449 &  x452 &  x458 &  x464 &  x470 &  x472 &  x473 &  x482 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x511 &  x512 &  x515 &  x518 &  x521 &  x539 &  x542 &  x545 &  x548 &  x556 &  x563 &  x569 &  x575 &  x578 &  x584 &  x587 &  x592 &  x595 &  x596 &  x599 &  x602 &  x617 &  x629 &  x631 &  x632 &  x635 &  x638 &  x641 &  x647 &  x653 &  x662 &  x668 &  x670 &  x671 &  x677 &  x680 &  x692 &  x707 &  x709 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x743 &  x746 &  x749 &  x755 &  x758 &  x767 &  x773 &  x776 &  x779 &  x782 &  x787 &  x788 &  x791 &  x797 &  x806 &  x812 &  x815 &  x818 &  x821 &  x824 &  x826 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x851 &  x854 &  x857 &  x860 &  x866 &  x872 &  x875 &  x878 &  x887 &  x890 &  x893 &  x896 &  x902 &  x905 &  x914 &  x917 &  x923 &  x932 &  x941 &  x943 &  x944 &  x947 &  x950 &  x953 &  x956 &  x965 &  x974 &  x977 &  x980 &  x983 &  x986 &  x994 &  x995 &  x1004 &  x1007 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1066 &  x1067 &  x1070 &  x1079 &  x1085 &  x1088 &  x1094 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1127 &  x1130 & ~x483 & ~x585 & ~x624 & ~x645 & ~x702 & ~x780;
assign c1184 =  x1 &  x2 &  x5 &  x8 &  x10 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x40 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x79 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x137 &  x140 &  x143 &  x152 &  x155 &  x157 &  x158 &  x167 &  x170 &  x173 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x196 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x235 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x290 &  x293 &  x296 &  x302 &  x305 &  x308 &  x314 &  x317 &  x320 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x395 &  x398 &  x400 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x572 &  x578 &  x581 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x638 &  x641 &  x647 &  x650 &  x653 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x697 &  x698 &  x701 &  x710 &  x713 &  x719 &  x722 &  x728 &  x731 &  x734 &  x736 &  x740 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x775 &  x776 &  x779 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x812 &  x815 &  x818 &  x821 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1043 &  x1046 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x6 & ~x45 & ~x123 & ~x162 & ~x246 & ~x753 & ~x831 & ~x870 & ~x1032 & ~x1065 & ~x1071 & ~x1104;
assign c1186 =  x8 &  x14 &  x35 &  x38 &  x41 &  x44 &  x47 &  x53 &  x65 &  x68 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x107 &  x113 &  x122 &  x128 &  x137 &  x149 &  x158 &  x161 &  x164 &  x170 &  x182 &  x185 &  x188 &  x194 &  x197 &  x206 &  x209 &  x212 &  x233 &  x236 &  x239 &  x251 &  x260 &  x263 &  x269 &  x275 &  x284 &  x287 &  x293 &  x299 &  x305 &  x308 &  x323 &  x329 &  x332 &  x338 &  x341 &  x347 &  x350 &  x353 &  x356 &  x362 &  x368 &  x374 &  x380 &  x383 &  x389 &  x395 &  x398 &  x401 &  x404 &  x410 &  x416 &  x425 &  x428 &  x433 &  x437 &  x449 &  x452 &  x455 &  x458 &  x467 &  x470 &  x472 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x512 &  x515 &  x524 &  x533 &  x542 &  x548 &  x554 &  x557 &  x566 &  x575 &  x590 &  x593 &  x602 &  x605 &  x614 &  x617 &  x620 &  x626 &  x631 &  x632 &  x644 &  x647 &  x650 &  x656 &  x659 &  x668 &  x677 &  x692 &  x695 &  x704 &  x716 &  x731 &  x734 &  x737 &  x740 &  x748 &  x749 &  x761 &  x764 &  x767 &  x770 &  x776 &  x794 &  x797 &  x800 &  x821 &  x827 &  x833 &  x839 &  x845 &  x848 &  x851 &  x863 &  x872 &  x878 &  x881 &  x887 &  x890 &  x896 &  x899 &  x902 &  x905 &  x908 &  x917 &  x923 &  x935 &  x944 &  x947 &  x956 &  x962 &  x965 &  x968 &  x971 &  x983 &  x989 &  x1001 &  x1007 &  x1010 &  x1016 &  x1034 &  x1040 &  x1046 &  x1052 &  x1055 &  x1058 &  x1067 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1112 &  x1124 & ~x420 & ~x498 & ~x600 & ~x639 & ~x678 & ~x717 & ~x897 & ~x951 & ~x1014 & ~x1023 & ~x1053 & ~x1063 & ~x1101 & ~x1102;
assign c1188 =  x2 &  x11 &  x14 &  x17 &  x32 &  x35 &  x38 &  x44 &  x47 &  x50 &  x53 &  x56 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x107 &  x113 &  x116 &  x122 &  x128 &  x131 &  x134 &  x140 &  x146 &  x149 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x176 &  x179 &  x185 &  x188 &  x191 &  x197 &  x206 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x245 &  x251 &  x254 &  x257 &  x266 &  x269 &  x272 &  x275 &  x281 &  x290 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x317 &  x323 &  x326 &  x332 &  x335 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x362 &  x365 &  x368 &  x374 &  x377 &  x380 &  x386 &  x392 &  x395 &  x398 &  x401 &  x404 &  x410 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x449 &  x452 &  x458 &  x461 &  x464 &  x467 &  x470 &  x476 &  x479 &  x481 &  x482 &  x485 &  x488 &  x494 &  x497 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x569 &  x572 &  x578 &  x584 &  x593 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x626 &  x629 &  x635 &  x638 &  x644 &  x647 &  x653 &  x656 &  x659 &  x665 &  x668 &  x671 &  x674 &  x680 &  x686 &  x692 &  x695 &  x698 &  x704 &  x716 &  x722 &  x725 &  x728 &  x731 &  x743 &  x745 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x776 &  x779 &  x782 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x821 &  x823 &  x827 &  x830 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x860 &  x863 &  x866 &  x872 &  x878 &  x887 &  x890 &  x901 &  x902 &  x905 &  x908 &  x911 &  x917 &  x920 &  x923 &  x926 &  x929 &  x938 &  x940 &  x941 &  x944 &  x947 &  x950 &  x965 &  x971 &  x979 &  x980 &  x982 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1018 &  x1019 &  x1022 &  x1028 &  x1031 &  x1037 &  x1040 &  x1049 &  x1055 &  x1058 &  x1061 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1127 & ~x606 & ~x873 & ~x912 & ~x915 & ~x918 & ~x993 & ~x1029 & ~x1032 & ~x1068 & ~x1074 & ~x1113;
assign c1190 =  x2 &  x5 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x164 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x191 &  x194 &  x197 &  x200 &  x206 &  x209 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x341 &  x344 &  x347 &  x350 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x440 &  x443 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x605 &  x611 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x701 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x776 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x893 &  x896 &  x899 &  x901 &  x902 &  x905 &  x911 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1018 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1057 &  x1058 &  x1059 &  x1060 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1099 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130 & ~x732 & ~x772 & ~x810 & ~x811 & ~x849 & ~x850 & ~x888 & ~x927;
assign c1192 =  x2 &  x5 &  x8 &  x11 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x59 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x142 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x188 &  x191 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x220 &  x221 &  x230 &  x236 &  x239 &  x242 &  x248 &  x251 &  x253 &  x254 &  x259 &  x260 &  x263 &  x266 &  x269 &  x272 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x304 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x326 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x370 &  x371 &  x374 &  x377 &  x380 &  x383 &  x389 &  x392 &  x395 &  x398 &  x407 &  x410 &  x416 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x470 &  x473 &  x482 &  x485 &  x488 &  x491 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x542 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x611 &  x614 &  x620 &  x623 &  x626 &  x629 &  x635 &  x638 &  x644 &  x650 &  x656 &  x659 &  x665 &  x671 &  x674 &  x677 &  x680 &  x683 &  x689 &  x692 &  x695 &  x698 &  x701 &  x707 &  x710 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x749 &  x752 &  x755 &  x758 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x839 &  x842 &  x845 &  x854 &  x857 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1085 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 & ~x81 & ~x120 & ~x198 & ~x237 & ~x276 & ~x315 & ~x318 & ~x474 & ~x480 & ~x513 & ~x552;
assign c1194 =  x2 &  x5 &  x11 &  x14 &  x17 &  x23 &  x26 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x95 &  x104 &  x107 &  x113 &  x116 &  x119 &  x122 &  x128 &  x131 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x242 &  x245 &  x248 &  x251 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x278 &  x281 &  x284 &  x287 &  x290 &  x296 &  x299 &  x302 &  x308 &  x311 &  x314 &  x320 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x353 &  x356 &  x362 &  x368 &  x371 &  x374 &  x389 &  x392 &  x398 &  x404 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x431 &  x434 &  x440 &  x443 &  x449 &  x455 &  x458 &  x461 &  x464 &  x470 &  x473 &  x476 &  x479 &  x482 &  x488 &  x494 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x524 &  x527 &  x530 &  x533 &  x539 &  x542 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x572 &  x575 &  x581 &  x587 &  x590 &  x596 &  x599 &  x604 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x629 &  x632 &  x635 &  x638 &  x641 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x671 &  x680 &  x683 &  x692 &  x695 &  x698 &  x701 &  x704 &  x706 &  x710 &  x716 &  x719 &  x725 &  x731 &  x734 &  x740 &  x746 &  x752 &  x755 &  x761 &  x764 &  x767 &  x773 &  x779 &  x784 &  x788 &  x791 &  x794 &  x803 &  x806 &  x812 &  x821 &  x823 &  x824 &  x827 &  x830 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x893 &  x899 &  x901 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x956 &  x962 &  x965 &  x968 &  x971 &  x974 &  x979 &  x980 &  x983 &  x985 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1016 &  x1031 &  x1034 &  x1040 &  x1043 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1115 &  x1121 &  x1124 &  x1127 & ~x195 & ~x234 & ~x552 & ~x657 & ~x669;
assign c1196 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x116 &  x119 &  x122 &  x125 &  x128 &  x130 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x290 &  x293 &  x296 &  x299 &  x302 &  x304 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x338 &  x341 &  x343 &  x344 &  x350 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x380 &  x382 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x470 &  x473 &  x476 &  x482 &  x485 &  x488 &  x491 &  x494 &  x506 &  x509 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x587 &  x590 &  x596 &  x599 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x683 &  x686 &  x689 &  x692 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x728 &  x731 &  x740 &  x743 &  x746 &  x749 &  x752 &  x758 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x812 &  x815 &  x821 &  x823 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x868 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x901 &  x902 &  x905 &  x907 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x940 &  x941 &  x946 &  x947 &  x950 &  x953 &  x959 &  x962 &  x968 &  x971 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1013 &  x1016 &  x1018 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1057 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1127 & ~x738 & ~x739 & ~x777;
assign c1198 =  x1 &  x5 &  x8 &  x11 &  x17 &  x29 &  x32 &  x35 &  x41 &  x47 &  x50 &  x53 &  x56 &  x62 &  x71 &  x74 &  x77 &  x80 &  x83 &  x89 &  x95 &  x107 &  x113 &  x122 &  x125 &  x131 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x155 &  x158 &  x164 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x227 &  x230 &  x236 &  x242 &  x245 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x335 &  x341 &  x347 &  x350 &  x353 &  x356 &  x359 &  x368 &  x371 &  x380 &  x383 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x443 &  x449 &  x452 &  x455 &  x461 &  x464 &  x467 &  x470 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x506 &  x512 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x539 &  x545 &  x548 &  x551 &  x560 &  x562 &  x563 &  x569 &  x575 &  x593 &  x596 &  x602 &  x605 &  x608 &  x614 &  x620 &  x623 &  x626 &  x635 &  x638 &  x641 &  x647 &  x653 &  x656 &  x662 &  x665 &  x677 &  x680 &  x683 &  x686 &  x689 &  x695 &  x701 &  x704 &  x707 &  x713 &  x716 &  x719 &  x725 &  x728 &  x734 &  x737 &  x743 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x779 &  x782 &  x788 &  x791 &  x797 &  x800 &  x803 &  x809 &  x812 &  x815 &  x818 &  x820 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x845 &  x848 &  x851 &  x854 &  x857 &  x859 &  x863 &  x869 &  x872 &  x875 &  x881 &  x884 &  x887 &  x890 &  x896 &  x898 &  x899 &  x905 &  x911 &  x914 &  x917 &  x923 &  x926 &  x932 &  x937 &  x938 &  x941 &  x944 &  x947 &  x956 &  x959 &  x962 &  x976 &  x977 &  x980 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1054 &  x1064 &  x1067 &  x1073 &  x1079 &  x1085 &  x1091 &  x1094 &  x1100 &  x1103 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x180 & ~x219 & ~x393 & ~x510 & ~x660 & ~x1005 & ~x1032 & ~x1065 & ~x1071 & ~x1077 & ~x1089;
assign c1200 =  x2 &  x5 &  x8 &  x14 &  x17 &  x23 &  x29 &  x35 &  x38 &  x44 &  x47 &  x56 &  x59 &  x62 &  x65 &  x68 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x101 &  x104 &  x107 &  x113 &  x116 &  x119 &  x122 &  x128 &  x131 &  x137 &  x140 &  x149 &  x155 &  x160 &  x161 &  x164 &  x170 &  x176 &  x179 &  x182 &  x185 &  x188 &  x194 &  x197 &  x199 &  x206 &  x209 &  x215 &  x218 &  x224 &  x227 &  x230 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x266 &  x269 &  x272 &  x277 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x314 &  x316 &  x317 &  x323 &  x326 &  x329 &  x338 &  x344 &  x347 &  x350 &  x355 &  x359 &  x361 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x394 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x419 &  x422 &  x428 &  x431 &  x433 &  x440 &  x446 &  x449 &  x452 &  x458 &  x461 &  x464 &  x470 &  x473 &  x479 &  x482 &  x491 &  x494 &  x497 &  x503 &  x512 &  x514 &  x521 &  x527 &  x530 &  x533 &  x536 &  x545 &  x551 &  x553 &  x557 &  x560 &  x566 &  x569 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x626 &  x629 &  x632 &  x641 &  x650 &  x653 &  x659 &  x665 &  x671 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x704 &  x710 &  x713 &  x716 &  x722 &  x725 &  x727 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x758 &  x767 &  x770 &  x772 &  x773 &  x776 &  x779 &  x782 &  x788 &  x791 &  x794 &  x805 &  x806 &  x811 &  x812 &  x815 &  x821 &  x824 &  x833 &  x836 &  x842 &  x844 &  x845 &  x848 &  x854 &  x857 &  x860 &  x863 &  x872 &  x875 &  x883 &  x884 &  x887 &  x890 &  x896 &  x911 &  x914 &  x917 &  x926 &  x929 &  x932 &  x941 &  x947 &  x953 &  x956 &  x961 &  x962 &  x965 &  x971 &  x974 &  x977 &  x980 &  x986 &  x998 &  x1001 &  x1010 &  x1016 &  x1022 &  x1034 &  x1040 &  x1043 &  x1049 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 & ~x483 & ~x507 & ~x546 & ~x561 & ~x606 & ~x624 & ~x645 & ~x663 & ~x702 & ~x741 & ~x780 & ~x858;
assign c1202 =  x2 &  x8 &  x17 &  x23 &  x26 &  x29 &  x35 &  x38 &  x44 &  x53 &  x56 &  x71 &  x74 &  x77 &  x89 &  x95 &  x107 &  x110 &  x113 &  x116 &  x122 &  x128 &  x131 &  x134 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x179 &  x182 &  x188 &  x191 &  x194 &  x197 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x230 &  x233 &  x236 &  x239 &  x245 &  x251 &  x257 &  x269 &  x272 &  x275 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x317 &  x323 &  x326 &  x335 &  x338 &  x341 &  x344 &  x350 &  x353 &  x377 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x433 &  x434 &  x437 &  x440 &  x443 &  x449 &  x452 &  x461 &  x467 &  x476 &  x479 &  x482 &  x488 &  x491 &  x494 &  x497 &  x506 &  x509 &  x512 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x557 &  x560 &  x566 &  x572 &  x575 &  x578 &  x584 &  x587 &  x590 &  x593 &  x605 &  x614 &  x617 &  x620 &  x623 &  x626 &  x632 &  x635 &  x647 &  x653 &  x656 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x701 &  x704 &  x709 &  x710 &  x713 &  x716 &  x722 &  x725 &  x731 &  x734 &  x737 &  x743 &  x749 &  x767 &  x773 &  x785 &  x787 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x854 &  x857 &  x865 &  x866 &  x869 &  x872 &  x877 &  x878 &  x881 &  x887 &  x893 &  x896 &  x899 &  x908 &  x914 &  x917 &  x923 &  x932 &  x944 &  x947 &  x950 &  x953 &  x955 &  x956 &  x959 &  x962 &  x968 &  x974 &  x977 &  x983 &  x986 &  x995 &  x1004 &  x1007 &  x1016 &  x1019 &  x1027 &  x1028 &  x1031 &  x1033 &  x1037 &  x1040 &  x1043 &  x1046 &  x1055 &  x1058 &  x1061 &  x1066 &  x1067 &  x1073 &  x1076 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1115 &  x1121 &  x1127 & ~x420 & ~x459 & ~x460 & ~x537 & ~x936 & ~x1017 & ~x1056;
assign c1204 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x26 &  x29 &  x41 &  x47 &  x50 &  x53 &  x56 &  x62 &  x65 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x122 &  x128 &  x131 &  x134 &  x140 &  x143 &  x146 &  x152 &  x158 &  x161 &  x164 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x209 &  x212 &  x215 &  x221 &  x224 &  x233 &  x236 &  x239 &  x242 &  x248 &  x254 &  x257 &  x263 &  x266 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x296 &  x302 &  x305 &  x311 &  x314 &  x317 &  x320 &  x329 &  x335 &  x338 &  x343 &  x344 &  x353 &  x359 &  x362 &  x365 &  x371 &  x374 &  x380 &  x382 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x404 &  x407 &  x415 &  x416 &  x419 &  x422 &  x425 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x455 &  x460 &  x473 &  x476 &  x479 &  x482 &  x488 &  x494 &  x497 &  x503 &  x506 &  x512 &  x515 &  x518 &  x521 &  x524 &  x526 &  x530 &  x533 &  x536 &  x539 &  x548 &  x557 &  x560 &  x563 &  x565 &  x566 &  x569 &  x572 &  x578 &  x584 &  x587 &  x593 &  x596 &  x601 &  x605 &  x617 &  x626 &  x629 &  x632 &  x635 &  x640 &  x641 &  x647 &  x653 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x704 &  x710 &  x716 &  x725 &  x728 &  x731 &  x734 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x764 &  x767 &  x776 &  x779 &  x782 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x815 &  x818 &  x824 &  x827 &  x833 &  x836 &  x839 &  x842 &  x845 &  x851 &  x854 &  x860 &  x862 &  x863 &  x866 &  x872 &  x875 &  x884 &  x887 &  x893 &  x896 &  x898 &  x899 &  x901 &  x902 &  x905 &  x911 &  x914 &  x917 &  x920 &  x929 &  x932 &  x937 &  x938 &  x941 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x976 &  x980 &  x983 &  x986 &  x995 &  x998 &  x1001 &  x1015 &  x1016 &  x1017 &  x1022 &  x1031 &  x1034 &  x1043 &  x1046 &  x1049 &  x1052 &  x1054 &  x1055 &  x1057 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1096 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x198 & ~x237 & ~x276 & ~x312 & ~x315 & ~x351 & ~x354 & ~x393 & ~x429 & ~x432 & ~x510 & ~x549 & ~x1032 & ~x1071;
assign c1206 =  x2 &  x5 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x107 &  x110 &  x113 &  x122 &  x125 &  x137 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x242 &  x245 &  x248 &  x251 &  x254 &  x260 &  x263 &  x266 &  x269 &  x271 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x292 &  x293 &  x296 &  x299 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x344 &  x346 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x428 &  x431 &  x434 &  x437 &  x443 &  x449 &  x452 &  x455 &  x458 &  x464 &  x467 &  x470 &  x476 &  x479 &  x482 &  x485 &  x487 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x548 &  x551 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x611 &  x614 &  x617 &  x620 &  x625 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x647 &  x653 &  x656 &  x659 &  x662 &  x668 &  x671 &  x674 &  x689 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x745 &  x746 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x773 &  x776 &  x779 &  x782 &  x784 &  x785 &  x788 &  x791 &  x800 &  x803 &  x818 &  x821 &  x823 &  x824 &  x829 &  x833 &  x836 &  x842 &  x845 &  x848 &  x851 &  x857 &  x863 &  x869 &  x872 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x947 &  x950 &  x953 &  x959 &  x962 &  x965 &  x971 &  x977 &  x980 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1058 &  x1061 &  x1067 &  x1070 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x237 & ~x276 & ~x315 & ~x354 & ~x513 & ~x552;
assign c1208 =  x2 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x35 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x97 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x136 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x164 &  x167 &  x170 &  x173 &  x175 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x197 &  x200 &  x203 &  x209 &  x212 &  x214 &  x215 &  x218 &  x221 &  x224 &  x227 &  x236 &  x239 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x326 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x353 &  x356 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x584 &  x590 &  x593 &  x596 &  x599 &  x605 &  x608 &  x611 &  x614 &  x626 &  x632 &  x638 &  x641 &  x644 &  x647 &  x656 &  x662 &  x665 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x713 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x746 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x779 &  x782 &  x791 &  x794 &  x800 &  x803 &  x806 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x854 &  x857 &  x863 &  x866 &  x872 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x929 &  x932 &  x935 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x977 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1070 &  x1073 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1130 & ~x336 & ~x660 & ~x699 & ~x816 & ~x855 & ~x912 & ~x951 & ~x990 & ~x1029 & ~x1068 & ~x1107;
assign c1210 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x50 &  x53 &  x56 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x104 &  x107 &  x110 &  x116 &  x122 &  x128 &  x131 &  x134 &  x137 &  x143 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x191 &  x194 &  x197 &  x200 &  x206 &  x209 &  x212 &  x218 &  x221 &  x227 &  x230 &  x233 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x290 &  x296 &  x302 &  x305 &  x308 &  x311 &  x320 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x404 &  x407 &  x409 &  x410 &  x413 &  x416 &  x434 &  x437 &  x440 &  x443 &  x446 &  x448 &  x449 &  x452 &  x458 &  x461 &  x464 &  x467 &  x470 &  x476 &  x479 &  x487 &  x488 &  x491 &  x497 &  x503 &  x509 &  x512 &  x515 &  x518 &  x524 &  x525 &  x526 &  x527 &  x530 &  x536 &  x539 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x565 &  x566 &  x569 &  x572 &  x578 &  x581 &  x584 &  x587 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x656 &  x659 &  x662 &  x665 &  x668 &  x674 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x703 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x731 &  x734 &  x737 &  x740 &  x742 &  x746 &  x749 &  x752 &  x758 &  x761 &  x764 &  x770 &  x773 &  x776 &  x782 &  x785 &  x788 &  x791 &  x800 &  x803 &  x806 &  x809 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x854 &  x857 &  x866 &  x869 &  x872 &  x875 &  x878 &  x884 &  x887 &  x890 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x923 &  x926 &  x932 &  x935 &  x938 &  x940 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1043 &  x1046 &  x1049 &  x1055 &  x1060 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x78 & ~x117 & ~x156 & ~x195 & ~x273 & ~x312 & ~x351 & ~x354 & ~x393 & ~x438;
assign c1212 =  x2 &  x5 &  x11 &  x14 &  x20 &  x25 &  x26 &  x29 &  x32 &  x35 &  x37 &  x41 &  x47 &  x52 &  x53 &  x56 &  x59 &  x62 &  x64 &  x68 &  x76 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x103 &  x107 &  x119 &  x122 &  x131 &  x134 &  x137 &  x146 &  x152 &  x155 &  x158 &  x161 &  x164 &  x170 &  x188 &  x191 &  x194 &  x197 &  x206 &  x209 &  x215 &  x221 &  x224 &  x227 &  x230 &  x242 &  x245 &  x248 &  x254 &  x266 &  x269 &  x275 &  x293 &  x296 &  x308 &  x320 &  x326 &  x329 &  x332 &  x338 &  x344 &  x347 &  x353 &  x359 &  x362 &  x365 &  x368 &  x389 &  x392 &  x401 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x428 &  x437 &  x446 &  x449 &  x452 &  x455 &  x461 &  x470 &  x476 &  x482 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x511 &  x515 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x542 &  x545 &  x554 &  x557 &  x560 &  x572 &  x575 &  x581 &  x584 &  x593 &  x596 &  x599 &  x602 &  x608 &  x614 &  x617 &  x626 &  x632 &  x650 &  x653 &  x659 &  x662 &  x665 &  x667 &  x668 &  x674 &  x677 &  x680 &  x692 &  x695 &  x698 &  x706 &  x707 &  x716 &  x722 &  x725 &  x728 &  x731 &  x734 &  x740 &  x746 &  x749 &  x752 &  x755 &  x761 &  x764 &  x770 &  x773 &  x782 &  x785 &  x788 &  x794 &  x800 &  x806 &  x809 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x854 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x890 &  x893 &  x896 &  x899 &  x902 &  x904 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x967 &  x977 &  x980 &  x995 &  x998 &  x1001 &  x1013 &  x1016 &  x1025 &  x1028 &  x1031 &  x1037 &  x1043 &  x1049 &  x1051 &  x1058 &  x1061 &  x1064 &  x1073 &  x1076 &  x1088 &  x1090 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1127 &  x1129 & ~x918 & ~x936 & ~x957 & ~x1014 & ~x1092;
assign c1214 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x101 &  x107 &  x110 &  x113 &  x119 &  x122 &  x128 &  x131 &  x134 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x161 &  x164 &  x170 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x275 &  x278 &  x281 &  x284 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x371 &  x374 &  x376 &  x377 &  x380 &  x382 &  x383 &  x389 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x415 &  x416 &  x421 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x448 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x491 &  x494 &  x497 &  x500 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x526 &  x530 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x562 &  x563 &  x565 &  x566 &  x569 &  x572 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x599 &  x601 &  x602 &  x604 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x719 &  x722 &  x725 &  x728 &  x734 &  x737 &  x740 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x901 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x938 &  x940 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x977 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1018 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x9 & ~x126 & ~x432 & ~x657 & ~x813;
assign c1216 =  x2 &  x5 &  x8 &  x11 &  x20 &  x26 &  x29 &  x38 &  x41 &  x44 &  x62 &  x65 &  x68 &  x70 &  x71 &  x74 &  x77 &  x83 &  x95 &  x98 &  x101 &  x119 &  x122 &  x128 &  x134 &  x137 &  x140 &  x143 &  x152 &  x155 &  x161 &  x167 &  x170 &  x173 &  x182 &  x188 &  x206 &  x209 &  x212 &  x215 &  x227 &  x230 &  x233 &  x245 &  x248 &  x254 &  x257 &  x260 &  x269 &  x275 &  x278 &  x281 &  x284 &  x287 &  x289 &  x290 &  x296 &  x305 &  x308 &  x314 &  x323 &  x326 &  x329 &  x335 &  x338 &  x341 &  x350 &  x371 &  x374 &  x376 &  x382 &  x383 &  x386 &  x389 &  x406 &  x407 &  x413 &  x415 &  x422 &  x434 &  x443 &  x446 &  x455 &  x461 &  x467 &  x470 &  x473 &  x479 &  x482 &  x485 &  x488 &  x497 &  x506 &  x512 &  x518 &  x524 &  x527 &  x530 &  x533 &  x539 &  x545 &  x548 &  x551 &  x560 &  x562 &  x563 &  x569 &  x575 &  x584 &  x590 &  x596 &  x599 &  x601 &  x605 &  x617 &  x623 &  x629 &  x632 &  x640 &  x641 &  x659 &  x671 &  x680 &  x692 &  x701 &  x704 &  x710 &  x713 &  x716 &  x740 &  x743 &  x746 &  x755 &  x758 &  x761 &  x767 &  x776 &  x779 &  x782 &  x788 &  x794 &  x803 &  x806 &  x809 &  x812 &  x815 &  x824 &  x827 &  x842 &  x857 &  x860 &  x869 &  x875 &  x890 &  x899 &  x902 &  x908 &  x914 &  x917 &  x923 &  x929 &  x932 &  x935 &  x937 &  x941 &  x947 &  x950 &  x953 &  x956 &  x959 &  x974 &  x980 &  x989 &  x992 &  x995 &  x1004 &  x1007 &  x1010 &  x1022 &  x1028 &  x1031 &  x1034 &  x1046 &  x1049 &  x1052 &  x1061 &  x1064 &  x1070 &  x1073 &  x1088 &  x1091 &  x1100 &  x1106 &  x1118 &  x1121 &  x1124 &  x1130 & ~x390 & ~x915 & ~x951 & ~x993;
assign c1218 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x53 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x89 &  x92 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x188 &  x191 &  x194 &  x197 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x257 &  x263 &  x266 &  x269 &  x272 &  x281 &  x284 &  x287 &  x289 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x328 &  x329 &  x332 &  x335 &  x338 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x367 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x547 &  x548 &  x554 &  x557 &  x560 &  x566 &  x569 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x614 &  x617 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x656 &  x659 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x812 &  x815 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x842 &  x845 &  x848 &  x854 &  x857 &  x860 &  x866 &  x869 &  x872 &  x875 &  x878 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x983 &  x986 &  x989 &  x992 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 & ~x81 & ~x120 & ~x159 & ~x198 & ~x282 & ~x321 & ~x357 & ~x474 & ~x513 & ~x681;
assign c1220 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x275 &  x278 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x391 &  x392 &  x394 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x433 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x511 &  x512 &  x515 &  x517 &  x518 &  x521 &  x524 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x556 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x595 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x629 &  x633 &  x634 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x673 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x709 &  x710 &  x712 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x748 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x785 &  x787 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x815 &  x818 &  x821 &  x824 &  x826 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x381 & ~x420 & ~x459 & ~x741;
assign c1222 =  x1 &  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x40 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x547 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x667 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x784 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1006 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x321 & ~x360 & ~x435 & ~x474 & ~x513 & ~x552 & ~x720;
assign c1224 =  x2 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x50 &  x59 &  x77 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x116 &  x119 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x155 &  x158 &  x160 &  x161 &  x173 &  x179 &  x182 &  x185 &  x191 &  x194 &  x197 &  x199 &  x212 &  x215 &  x221 &  x224 &  x230 &  x233 &  x236 &  x238 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x266 &  x272 &  x277 &  x281 &  x284 &  x287 &  x290 &  x293 &  x299 &  x305 &  x308 &  x311 &  x314 &  x323 &  x335 &  x338 &  x350 &  x355 &  x362 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x398 &  x401 &  x404 &  x407 &  x410 &  x428 &  x431 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x464 &  x470 &  x476 &  x479 &  x485 &  x488 &  x500 &  x503 &  x506 &  x512 &  x515 &  x518 &  x521 &  x527 &  x533 &  x539 &  x542 &  x545 &  x551 &  x553 &  x554 &  x557 &  x563 &  x572 &  x578 &  x581 &  x590 &  x596 &  x599 &  x605 &  x611 &  x614 &  x620 &  x623 &  x631 &  x632 &  x647 &  x653 &  x656 &  x659 &  x668 &  x670 &  x671 &  x674 &  x676 &  x677 &  x680 &  x689 &  x692 &  x698 &  x701 &  x710 &  x713 &  x716 &  x728 &  x734 &  x746 &  x749 &  x752 &  x776 &  x782 &  x785 &  x794 &  x800 &  x803 &  x805 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x881 &  x884 &  x887 &  x893 &  x896 &  x899 &  x902 &  x908 &  x914 &  x920 &  x929 &  x932 &  x947 &  x950 &  x959 &  x968 &  x974 &  x980 &  x992 &  x995 &  x1004 &  x1007 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1034 &  x1037 &  x1043 &  x1046 &  x1058 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1094 &  x1106 &  x1118 &  x1121 &  x1130 & ~x99 & ~x309 & ~x405 & ~x444 & ~x483 & ~x546 & ~x585 & ~x624 & ~x663 & ~x702 & ~x741 & ~x780 & ~x819 & ~x858;
assign c1226 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x122 &  x125 &  x131 &  x134 &  x137 &  x140 &  x146 &  x149 &  x152 &  x155 &  x161 &  x164 &  x167 &  x170 &  x176 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x212 &  x218 &  x224 &  x233 &  x236 &  x239 &  x245 &  x248 &  x251 &  x254 &  x257 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x344 &  x350 &  x353 &  x359 &  x362 &  x365 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x394 &  x395 &  x398 &  x401 &  x404 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x433 &  x437 &  x446 &  x449 &  x455 &  x458 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x530 &  x533 &  x545 &  x548 &  x551 &  x554 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x611 &  x614 &  x617 &  x620 &  x632 &  x634 &  x638 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x665 &  x673 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x701 &  x704 &  x707 &  x710 &  x712 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x734 &  x737 &  x740 &  x743 &  x746 &  x748 &  x749 &  x751 &  x752 &  x755 &  x761 &  x764 &  x770 &  x773 &  x776 &  x779 &  x785 &  x787 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x818 &  x821 &  x824 &  x826 &  x830 &  x833 &  x836 &  x845 &  x848 &  x851 &  x854 &  x860 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x893 &  x899 &  x902 &  x905 &  x908 &  x914 &  x917 &  x920 &  x922 &  x926 &  x928 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x953 &  x959 &  x961 &  x962 &  x965 &  x967 &  x968 &  x971 &  x973 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x994 &  x995 &  x998 &  x1000 &  x1001 &  x1004 &  x1006 &  x1007 &  x1010 &  x1013 &  x1022 &  x1027 &  x1031 &  x1033 &  x1034 &  x1037 &  x1045 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1072 &  x1073 &  x1076 &  x1078 &  x1079 &  x1082 &  x1085 &  x1088 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1124 &  x1130 & ~x606 & ~x645 & ~x741 & ~x819 & ~x858 & ~x897 & ~x975 & ~x1053 & ~x1092;
assign c1228 =  x2 &  x8 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x74 &  x77 &  x80 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x188 &  x191 &  x194 &  x197 &  x203 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x257 &  x260 &  x269 &  x275 &  x278 &  x284 &  x287 &  x290 &  x296 &  x299 &  x305 &  x308 &  x314 &  x317 &  x320 &  x326 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x413 &  x415 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x488 &  x491 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x836 &  x839 &  x842 &  x845 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x968 &  x971 &  x974 &  x977 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1018 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x0 & ~x39 & ~x156 & ~x234 & ~x273 & ~x618 & ~x849 & ~x873 & ~x1029 & ~x1030 & ~x1068 & ~x1107 & ~x1113;
assign c1230 =  x2 &  x17 &  x32 &  x38 &  x53 &  x56 &  x68 &  x80 &  x89 &  x95 &  x98 &  x113 &  x116 &  x122 &  x137 &  x149 &  x161 &  x176 &  x196 &  x199 &  x209 &  x218 &  x221 &  x233 &  x238 &  x242 &  x277 &  x287 &  x290 &  x293 &  x296 &  x311 &  x316 &  x320 &  x335 &  x341 &  x356 &  x359 &  x365 &  x374 &  x377 &  x380 &  x383 &  x389 &  x392 &  x398 &  x401 &  x404 &  x410 &  x413 &  x428 &  x433 &  x434 &  x440 &  x443 &  x452 &  x467 &  x476 &  x479 &  x485 &  x488 &  x491 &  x503 &  x506 &  x509 &  x527 &  x530 &  x533 &  x539 &  x542 &  x545 &  x554 &  x566 &  x581 &  x598 &  x608 &  x614 &  x616 &  x617 &  x623 &  x626 &  x631 &  x641 &  x653 &  x656 &  x665 &  x671 &  x677 &  x683 &  x700 &  x704 &  x719 &  x722 &  x725 &  x734 &  x737 &  x740 &  x748 &  x761 &  x767 &  x773 &  x782 &  x788 &  x794 &  x797 &  x809 &  x812 &  x818 &  x824 &  x833 &  x836 &  x839 &  x848 &  x851 &  x865 &  x869 &  x875 &  x884 &  x899 &  x904 &  x911 &  x914 &  x923 &  x926 &  x938 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x973 &  x977 &  x980 &  x983 &  x988 &  x998 &  x1004 &  x1019 &  x1022 &  x1025 &  x1034 &  x1043 &  x1046 &  x1070 &  x1088 &  x1091 &  x1097 &  x1103 &  x1106 &  x1127 &  x1130 & ~x303 & ~x897 & ~x936;
assign c1232 =  x5 &  x8 &  x14 &  x20 &  x23 &  x26 &  x29 &  x38 &  x41 &  x44 &  x47 &  x56 &  x59 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x92 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x131 &  x134 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x167 &  x170 &  x176 &  x179 &  x182 &  x185 &  x194 &  x203 &  x206 &  x209 &  x212 &  x218 &  x221 &  x227 &  x230 &  x233 &  x236 &  x239 &  x245 &  x251 &  x263 &  x266 &  x269 &  x272 &  x278 &  x281 &  x284 &  x290 &  x293 &  x296 &  x305 &  x308 &  x311 &  x314 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x343 &  x344 &  x353 &  x362 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x407 &  x410 &  x413 &  x425 &  x428 &  x431 &  x437 &  x446 &  x458 &  x467 &  x470 &  x473 &  x482 &  x485 &  x488 &  x494 &  x500 &  x503 &  x506 &  x515 &  x518 &  x521 &  x524 &  x533 &  x536 &  x539 &  x545 &  x548 &  x557 &  x563 &  x569 &  x572 &  x575 &  x578 &  x584 &  x587 &  x590 &  x593 &  x596 &  x601 &  x602 &  x608 &  x611 &  x614 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x644 &  x650 &  x653 &  x656 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x695 &  x698 &  x703 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x728 &  x734 &  x737 &  x740 &  x742 &  x749 &  x752 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x784 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x812 &  x815 &  x818 &  x823 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x854 &  x857 &  x862 &  x863 &  x866 &  x869 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x899 &  x900 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x935 &  x939 &  x940 &  x947 &  x956 &  x962 &  x965 &  x971 &  x977 &  x979 &  x980 &  x983 &  x992 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1061 &  x1070 &  x1073 &  x1082 &  x1085 &  x1088 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1130 & ~x657 & ~x660 & ~x699 & ~x777;
assign c1234 =  x5 &  x14 &  x17 &  x32 &  x38 &  x56 &  x59 &  x80 &  x83 &  x86 &  x92 &  x95 &  x101 &  x113 &  x122 &  x125 &  x128 &  x131 &  x143 &  x149 &  x155 &  x158 &  x161 &  x167 &  x176 &  x182 &  x185 &  x188 &  x215 &  x221 &  x224 &  x233 &  x242 &  x245 &  x251 &  x254 &  x257 &  x263 &  x266 &  x272 &  x275 &  x293 &  x296 &  x311 &  x317 &  x320 &  x323 &  x329 &  x335 &  x338 &  x347 &  x353 &  x356 &  x362 &  x365 &  x392 &  x401 &  x403 &  x428 &  x440 &  x443 &  x458 &  x461 &  x467 &  x473 &  x479 &  x488 &  x500 &  x509 &  x527 &  x536 &  x539 &  x548 &  x551 &  x554 &  x557 &  x560 &  x581 &  x584 &  x586 &  x590 &  x593 &  x596 &  x599 &  x620 &  x635 &  x638 &  x653 &  x656 &  x662 &  x665 &  x668 &  x674 &  x686 &  x695 &  x704 &  x707 &  x725 &  x731 &  x734 &  x740 &  x742 &  x743 &  x761 &  x764 &  x776 &  x782 &  x785 &  x788 &  x797 &  x800 &  x823 &  x827 &  x833 &  x836 &  x860 &  x863 &  x872 &  x875 &  x884 &  x899 &  x901 &  x902 &  x920 &  x923 &  x938 &  x941 &  x944 &  x950 &  x953 &  x956 &  x965 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x1004 &  x1007 &  x1013 &  x1025 &  x1028 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1079 &  x1094 &  x1097 &  x1109 &  x1124 &  x1127 & ~x315 & ~x393 & ~x432 & ~x555 & ~x594 & ~x636 & ~x714 & ~x951;
assign c1236 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x44 &  x47 &  x50 &  x56 &  x59 &  x65 &  x68 &  x71 &  x74 &  x77 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x104 &  x107 &  x110 &  x113 &  x119 &  x122 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x284 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x319 &  x323 &  x329 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x389 &  x392 &  x395 &  x397 &  x398 &  x403 &  x404 &  x407 &  x413 &  x416 &  x419 &  x422 &  x425 &  x431 &  x434 &  x440 &  x442 &  x443 &  x446 &  x452 &  x455 &  x461 &  x467 &  x470 &  x473 &  x475 &  x476 &  x479 &  x482 &  x485 &  x488 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x520 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x542 &  x545 &  x548 &  x551 &  x553 &  x554 &  x557 &  x560 &  x563 &  x572 &  x578 &  x581 &  x587 &  x590 &  x593 &  x596 &  x598 &  x602 &  x605 &  x608 &  x614 &  x617 &  x620 &  x623 &  x626 &  x632 &  x635 &  x638 &  x647 &  x650 &  x656 &  x659 &  x662 &  x668 &  x671 &  x674 &  x676 &  x677 &  x680 &  x683 &  x686 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x715 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x752 &  x755 &  x758 &  x761 &  x766 &  x767 &  x770 &  x773 &  x778 &  x779 &  x785 &  x788 &  x793 &  x794 &  x797 &  x800 &  x805 &  x806 &  x812 &  x818 &  x821 &  x827 &  x832 &  x833 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x869 &  x871 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x899 &  x902 &  x905 &  x908 &  x914 &  x920 &  x923 &  x926 &  x932 &  x938 &  x941 &  x944 &  x947 &  x949 &  x950 &  x953 &  x956 &  x959 &  x962 &  x968 &  x974 &  x977 &  x980 &  x983 &  x988 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 & ~x450;
assign c1238 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x338 &  x344 &  x347 &  x350 &  x356 &  x359 &  x362 &  x365 &  x368 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x404 &  x407 &  x410 &  x413 &  x415 &  x416 &  x419 &  x421 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x518 &  x521 &  x523 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x662 &  x665 &  x667 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x703 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x742 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x770 &  x773 &  x779 &  x781 &  x784 &  x785 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x820 &  x821 &  x823 &  x824 &  x827 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x859 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x898 &  x899 &  x901 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x940 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x234 & ~x273 & ~x312 & ~x351 & ~x390 & ~x477 & ~x591 & ~x630 & ~x669 & ~x759 & ~x798;
assign c1240 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x508 &  x509 &  x511 &  x512 &  x518 &  x521 &  x527 &  x533 &  x536 &  x539 &  x542 &  x545 &  x547 &  x548 &  x550 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x590 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x628 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x745 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x318 & ~x357 & ~x360 & ~x396 & ~x435 & ~x498 & ~x795 & ~x858 & ~x897;
assign c1242 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x112 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x151 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x190 &  x191 &  x194 &  x197 &  x200 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x284 &  x286 &  x287 &  x290 &  x293 &  x296 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x380 &  x383 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x626 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x722 &  x725 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x782 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x823 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x901 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x938 &  x940 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x977 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1021 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x234 & ~x273 & ~x654 & ~x693 & ~x732 & ~x733 & ~x771 & ~x795 & ~x834 & ~x873;
assign c1244 =  x2 &  x5 &  x11 &  x17 &  x20 &  x23 &  x26 &  x32 &  x35 &  x38 &  x44 &  x47 &  x56 &  x59 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x122 &  x128 &  x131 &  x134 &  x137 &  x143 &  x146 &  x149 &  x152 &  x155 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x181 &  x182 &  x185 &  x188 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x220 &  x221 &  x224 &  x227 &  x230 &  x232 &  x233 &  x236 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x259 &  x260 &  x263 &  x266 &  x271 &  x272 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x311 &  x317 &  x320 &  x323 &  x326 &  x329 &  x335 &  x344 &  x347 &  x350 &  x353 &  x368 &  x371 &  x374 &  x383 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x440 &  x443 &  x446 &  x455 &  x458 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x530 &  x533 &  x536 &  x539 &  x542 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x605 &  x608 &  x611 &  x620 &  x626 &  x629 &  x632 &  x638 &  x644 &  x647 &  x653 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x758 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x794 &  x797 &  x803 &  x812 &  x815 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x851 &  x854 &  x857 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x893 &  x899 &  x901 &  x902 &  x905 &  x908 &  x917 &  x920 &  x926 &  x929 &  x935 &  x938 &  x940 &  x941 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1019 &  x1021 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1088 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130 & ~x165 & ~x195 & ~x204 & ~x234 & ~x273 & ~x282 & ~x312 & ~x321 & ~x351 & ~x360 & ~x399 & ~x516 & ~x912 & ~x951 & ~x990 & ~x1029;
assign c1246 =  x2 &  x5 &  x8 &  x11 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x41 &  x44 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x91 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x122 &  x125 &  x128 &  x130 &  x131 &  x134 &  x140 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x169 &  x170 &  x173 &  x176 &  x182 &  x185 &  x191 &  x194 &  x197 &  x203 &  x206 &  x209 &  x212 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x350 &  x359 &  x362 &  x365 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x533 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x563 &  x566 &  x569 &  x572 &  x575 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x626 &  x628 &  x629 &  x632 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x743 &  x745 &  x749 &  x752 &  x758 &  x761 &  x764 &  x770 &  x773 &  x776 &  x779 &  x782 &  x784 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x809 &  x812 &  x815 &  x818 &  x821 &  x823 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x865 &  x866 &  x869 &  x872 &  x875 &  x878 &  x884 &  x890 &  x893 &  x896 &  x899 &  x903 &  x904 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x929 &  x932 &  x935 &  x941 &  x942 &  x943 &  x944 &  x947 &  x950 &  x953 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x117 & ~x156 & ~x195 & ~x858 & ~x897 & ~x918 & ~x936 & ~x975 & ~x1014 & ~x1053 & ~x1092;
assign c1248 =  x2 &  x8 &  x11 &  x14 &  x17 &  x20 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x89 &  x92 &  x101 &  x107 &  x113 &  x119 &  x125 &  x128 &  x134 &  x149 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x176 &  x179 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x215 &  x218 &  x221 &  x224 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x293 &  x296 &  x299 &  x305 &  x308 &  x314 &  x317 &  x326 &  x329 &  x335 &  x344 &  x350 &  x356 &  x359 &  x362 &  x365 &  x368 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x401 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x449 &  x464 &  x472 &  x479 &  x482 &  x491 &  x500 &  x503 &  x512 &  x517 &  x518 &  x521 &  x527 &  x530 &  x533 &  x539 &  x542 &  x545 &  x548 &  x557 &  x560 &  x563 &  x569 &  x575 &  x578 &  x584 &  x587 &  x593 &  x595 &  x596 &  x599 &  x605 &  x611 &  x623 &  x632 &  x644 &  x650 &  x656 &  x659 &  x665 &  x671 &  x677 &  x680 &  x683 &  x692 &  x698 &  x704 &  x707 &  x710 &  x716 &  x722 &  x727 &  x734 &  x740 &  x746 &  x749 &  x758 &  x761 &  x766 &  x770 &  x785 &  x794 &  x797 &  x800 &  x803 &  x805 &  x806 &  x812 &  x815 &  x818 &  x821 &  x824 &  x842 &  x845 &  x848 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x878 &  x881 &  x884 &  x893 &  x896 &  x899 &  x902 &  x908 &  x911 &  x917 &  x920 &  x929 &  x938 &  x941 &  x949 &  x953 &  x956 &  x965 &  x968 &  x977 &  x980 &  x988 &  x989 &  x992 &  x998 &  x1004 &  x1016 &  x1019 &  x1022 &  x1034 &  x1037 &  x1040 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1067 &  x1070 &  x1076 &  x1082 &  x1094 &  x1097 &  x1103 &  x1112 &  x1121 &  x1127 &  x1130 & ~x420 & ~x459 & ~x528 & ~x780 & ~x819;
assign c1250 =  x5 &  x8 &  x11 &  x14 &  x23 &  x29 &  x32 &  x38 &  x50 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x98 &  x101 &  x104 &  x107 &  x110 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x155 &  x158 &  x161 &  x164 &  x170 &  x176 &  x185 &  x188 &  x191 &  x197 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x224 &  x227 &  x230 &  x236 &  x239 &  x242 &  x245 &  x248 &  x254 &  x257 &  x263 &  x269 &  x275 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x380 &  x386 &  x389 &  x395 &  x404 &  x410 &  x413 &  x419 &  x422 &  x425 &  x428 &  x431 &  x437 &  x443 &  x449 &  x452 &  x458 &  x464 &  x467 &  x473 &  x476 &  x485 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x530 &  x533 &  x539 &  x542 &  x545 &  x551 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x584 &  x587 &  x593 &  x596 &  x602 &  x605 &  x614 &  x617 &  x620 &  x623 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x671 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x725 &  x728 &  x731 &  x734 &  x737 &  x743 &  x752 &  x758 &  x764 &  x767 &  x776 &  x782 &  x785 &  x794 &  x797 &  x800 &  x803 &  x806 &  x818 &  x821 &  x824 &  x833 &  x836 &  x839 &  x842 &  x848 &  x851 &  x857 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x905 &  x914 &  x917 &  x923 &  x932 &  x938 &  x940 &  x944 &  x947 &  x950 &  x953 &  x956 &  x965 &  x971 &  x977 &  x979 &  x980 &  x983 &  x989 &  x992 &  x995 &  x1004 &  x1007 &  x1010 &  x1013 &  x1018 &  x1019 &  x1022 &  x1025 &  x1031 &  x1040 &  x1043 &  x1049 &  x1052 &  x1057 &  x1061 &  x1064 &  x1067 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1100 &  x1103 &  x1121 &  x1124 &  x1127 &  x1130 & ~x273 & ~x846 & ~x855 & ~x894 & ~x909 & ~x933 & ~x934 & ~x948 & ~x973 & ~x1011 & ~x1029 & ~x1050 & ~x1068;
assign c1252 =  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x305 &  x308 &  x311 &  x314 &  x317 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x415 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x454 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x518 &  x520 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x559 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x611 &  x614 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x662 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x863 &  x866 &  x869 &  x875 &  x878 &  x881 &  x887 &  x890 &  x893 &  x896 &  x899 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x87 & ~x390 & ~x429 & ~x468 & ~x507 & ~x528 & ~x585 & ~x645 & ~x723 & ~x762 & ~x801 & ~x840 & ~x879 & ~x918 & ~x957 & ~x996 & ~x1029 & ~x1035 & ~x1068 & ~x1074 & ~x1113;
assign c1254 =  x2 &  x5 &  x8 &  x11 &  x17 &  x20 &  x26 &  x29 &  x35 &  x38 &  x41 &  x44 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x80 &  x89 &  x92 &  x95 &  x101 &  x104 &  x107 &  x113 &  x116 &  x119 &  x122 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x191 &  x194 &  x197 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x230 &  x233 &  x245 &  x248 &  x251 &  x254 &  x257 &  x266 &  x269 &  x275 &  x278 &  x281 &  x284 &  x287 &  x293 &  x299 &  x308 &  x311 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x341 &  x344 &  x347 &  x350 &  x353 &  x355 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x380 &  x383 &  x389 &  x392 &  x394 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x446 &  x449 &  x455 &  x458 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x524 &  x527 &  x530 &  x533 &  x539 &  x542 &  x545 &  x548 &  x554 &  x557 &  x560 &  x563 &  x569 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x602 &  x605 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x638 &  x641 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x740 &  x743 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x770 &  x773 &  x776 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x812 &  x815 &  x821 &  x824 &  x827 &  x830 &  x833 &  x839 &  x848 &  x860 &  x866 &  x869 &  x878 &  x883 &  x887 &  x890 &  x893 &  x899 &  x902 &  x905 &  x908 &  x914 &  x920 &  x922 &  x923 &  x929 &  x935 &  x941 &  x947 &  x950 &  x956 &  x959 &  x962 &  x965 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x995 &  x1001 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x381 & ~x459 & ~x501 & ~x540 & ~x579 & ~x600 & ~x618 & ~x657 & ~x678 & ~x741 & ~x780 & ~x795 & ~x819 & ~x834 & ~x858 & ~x873 & ~x897 & ~x975 & ~x1068;
assign c1256 =  x1 &  x2 &  x5 &  x8 &  x14 &  x17 &  x29 &  x41 &  x47 &  x50 &  x53 &  x59 &  x65 &  x68 &  x74 &  x86 &  x98 &  x100 &  x101 &  x104 &  x113 &  x119 &  x122 &  x128 &  x131 &  x137 &  x139 &  x143 &  x146 &  x152 &  x164 &  x167 &  x170 &  x173 &  x182 &  x185 &  x188 &  x200 &  x206 &  x215 &  x227 &  x236 &  x245 &  x254 &  x257 &  x275 &  x278 &  x287 &  x290 &  x293 &  x296 &  x302 &  x305 &  x308 &  x311 &  x317 &  x332 &  x335 &  x338 &  x347 &  x353 &  x356 &  x365 &  x368 &  x374 &  x383 &  x389 &  x392 &  x395 &  x398 &  x403 &  x425 &  x427 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x452 &  x458 &  x464 &  x470 &  x476 &  x482 &  x485 &  x500 &  x506 &  x521 &  x530 &  x533 &  x545 &  x548 &  x551 &  x554 &  x557 &  x563 &  x572 &  x578 &  x581 &  x584 &  x590 &  x599 &  x602 &  x605 &  x608 &  x617 &  x620 &  x626 &  x629 &  x635 &  x638 &  x641 &  x647 &  x650 &  x653 &  x656 &  x662 &  x683 &  x692 &  x701 &  x706 &  x707 &  x713 &  x722 &  x725 &  x731 &  x742 &  x743 &  x746 &  x752 &  x755 &  x767 &  x770 &  x773 &  x779 &  x797 &  x800 &  x809 &  x812 &  x836 &  x854 &  x857 &  x859 &  x862 &  x863 &  x872 &  x875 &  x887 &  x896 &  x901 &  x905 &  x908 &  x911 &  x917 &  x926 &  x935 &  x938 &  x940 &  x947 &  x959 &  x962 &  x977 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x998 &  x1004 &  x1010 &  x1013 &  x1016 &  x1018 &  x1024 &  x1028 &  x1034 &  x1037 &  x1046 &  x1049 &  x1052 &  x1054 &  x1058 &  x1064 &  x1076 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1112 &  x1118 &  x1127 &  x1130 & ~x393 & ~x588 & ~x954 & ~x993 & ~x1032;
assign c1258 =  x2 &  x5 &  x8 &  x11 &  x14 &  x23 &  x35 &  x38 &  x47 &  x50 &  x59 &  x74 &  x77 &  x80 &  x89 &  x95 &  x98 &  x101 &  x104 &  x110 &  x119 &  x134 &  x137 &  x167 &  x173 &  x176 &  x182 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x218 &  x221 &  x224 &  x227 &  x230 &  x245 &  x251 &  x254 &  x257 &  x260 &  x263 &  x269 &  x281 &  x284 &  x287 &  x290 &  x293 &  x299 &  x302 &  x311 &  x317 &  x323 &  x326 &  x335 &  x338 &  x341 &  x344 &  x350 &  x353 &  x356 &  x359 &  x371 &  x377 &  x383 &  x392 &  x395 &  x401 &  x404 &  x410 &  x428 &  x434 &  x437 &  x443 &  x449 &  x458 &  x464 &  x482 &  x485 &  x488 &  x503 &  x518 &  x527 &  x530 &  x542 &  x554 &  x557 &  x560 &  x569 &  x575 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x608 &  x614 &  x617 &  x623 &  x638 &  x641 &  x647 &  x650 &  x659 &  x662 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x707 &  x710 &  x713 &  x716 &  x728 &  x731 &  x734 &  x737 &  x740 &  x746 &  x749 &  x761 &  x764 &  x767 &  x770 &  x776 &  x779 &  x784 &  x785 &  x788 &  x797 &  x800 &  x803 &  x809 &  x815 &  x821 &  x823 &  x824 &  x830 &  x839 &  x851 &  x854 &  x862 &  x863 &  x866 &  x875 &  x881 &  x902 &  x905 &  x917 &  x926 &  x929 &  x932 &  x938 &  x940 &  x944 &  x947 &  x950 &  x953 &  x956 &  x965 &  x977 &  x979 &  x980 &  x983 &  x995 &  x1001 &  x1004 &  x1007 &  x1016 &  x1018 &  x1019 &  x1022 &  x1025 &  x1031 &  x1037 &  x1043 &  x1052 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1100 &  x1112 &  x1118 &  x1130 & ~x195 & ~x234 & ~x261 & ~x273 & ~x300 & ~x339 & ~x378 & ~x456 & ~x855 & ~x894 & ~x972 & ~x973;
assign c1260 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x709 &  x710 &  x712 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x736 &  x737 &  x740 &  x743 &  x746 &  x748 &  x749 &  x751 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x775 &  x776 &  x782 &  x785 &  x787 &  x788 &  x790 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x829 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x868 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x907 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x946 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x985 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1024 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1063 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x582 & ~x621 & ~x684;
assign c1262 =  x2 &  x8 &  x11 &  x38 &  x41 &  x47 &  x59 &  x62 &  x71 &  x77 &  x86 &  x95 &  x101 &  x119 &  x122 &  x125 &  x131 &  x134 &  x152 &  x167 &  x170 &  x173 &  x182 &  x194 &  x206 &  x227 &  x236 &  x248 &  x260 &  x275 &  x281 &  x296 &  x305 &  x308 &  x326 &  x341 &  x344 &  x362 &  x365 &  x368 &  x371 &  x380 &  x386 &  x395 &  x404 &  x407 &  x428 &  x431 &  x434 &  x437 &  x440 &  x449 &  x458 &  x467 &  x482 &  x485 &  x491 &  x494 &  x503 &  x506 &  x515 &  x518 &  x521 &  x523 &  x524 &  x527 &  x542 &  x562 &  x563 &  x584 &  x587 &  x596 &  x601 &  x602 &  x608 &  x614 &  x617 &  x620 &  x629 &  x632 &  x635 &  x638 &  x644 &  x647 &  x653 &  x665 &  x671 &  x680 &  x683 &  x692 &  x701 &  x704 &  x707 &  x710 &  x722 &  x728 &  x731 &  x749 &  x755 &  x758 &  x764 &  x767 &  x770 &  x806 &  x809 &  x821 &  x833 &  x836 &  x851 &  x854 &  x857 &  x863 &  x872 &  x875 &  x878 &  x887 &  x890 &  x899 &  x901 &  x905 &  x917 &  x932 &  x935 &  x940 &  x947 &  x950 &  x953 &  x959 &  x965 &  x977 &  x986 &  x995 &  x1001 &  x1007 &  x1010 &  x1016 &  x1018 &  x1025 &  x1031 &  x1043 &  x1056 &  x1070 &  x1073 &  x1082 &  x1091 &  x1099 &  x1100 &  x1109 &  x1118 &  x1124 & ~x273 & ~x855 & ~x996;
assign c1264 =  x8 &  x29 &  x35 &  x44 &  x47 &  x53 &  x65 &  x68 &  x71 &  x80 &  x86 &  x95 &  x98 &  x101 &  x107 &  x110 &  x119 &  x122 &  x134 &  x143 &  x146 &  x152 &  x155 &  x179 &  x185 &  x188 &  x194 &  x203 &  x221 &  x236 &  x239 &  x251 &  x263 &  x266 &  x281 &  x287 &  x296 &  x302 &  x308 &  x311 &  x317 &  x323 &  x326 &  x338 &  x341 &  x344 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x386 &  x392 &  x407 &  x413 &  x419 &  x431 &  x434 &  x440 &  x449 &  x452 &  x458 &  x461 &  x464 &  x476 &  x479 &  x485 &  x497 &  x500 &  x514 &  x518 &  x520 &  x527 &  x530 &  x536 &  x539 &  x548 &  x553 &  x557 &  x559 &  x569 &  x572 &  x584 &  x587 &  x596 &  x599 &  x602 &  x605 &  x608 &  x610 &  x614 &  x620 &  x626 &  x629 &  x632 &  x635 &  x638 &  x647 &  x649 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x680 &  x688 &  x701 &  x704 &  x715 &  x716 &  x719 &  x725 &  x727 &  x728 &  x731 &  x734 &  x740 &  x743 &  x746 &  x749 &  x755 &  x761 &  x767 &  x776 &  x785 &  x788 &  x791 &  x806 &  x815 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x848 &  x860 &  x863 &  x872 &  x875 &  x881 &  x890 &  x902 &  x908 &  x911 &  x917 &  x920 &  x926 &  x935 &  x950 &  x956 &  x962 &  x968 &  x974 &  x977 &  x983 &  x995 &  x1001 &  x1004 &  x1007 &  x1016 &  x1028 &  x1043 &  x1046 &  x1052 &  x1055 &  x1067 &  x1079 &  x1082 &  x1091 &  x1097 &  x1109 &  x1112 &  x1115 &  x1118 &  x1127 &  x1130 & ~x165 & ~x189 & ~x228 & ~x585 & ~x625 & ~x657 & ~x663 & ~x664;
assign c1266 =  x2 &  x14 &  x35 &  x44 &  x53 &  x59 &  x68 &  x83 &  x86 &  x89 &  x95 &  x98 &  x113 &  x119 &  x122 &  x125 &  x131 &  x140 &  x146 &  x149 &  x152 &  x155 &  x161 &  x164 &  x173 &  x176 &  x179 &  x191 &  x197 &  x200 &  x209 &  x212 &  x215 &  x224 &  x227 &  x230 &  x233 &  x242 &  x251 &  x257 &  x266 &  x269 &  x275 &  x278 &  x281 &  x284 &  x293 &  x296 &  x302 &  x305 &  x314 &  x317 &  x326 &  x332 &  x341 &  x347 &  x356 &  x359 &  x371 &  x376 &  x383 &  x389 &  x398 &  x404 &  x416 &  x422 &  x425 &  x428 &  x434 &  x443 &  x452 &  x455 &  x461 &  x464 &  x467 &  x476 &  x479 &  x484 &  x485 &  x491 &  x494 &  x500 &  x515 &  x518 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x560 &  x563 &  x572 &  x578 &  x584 &  x587 &  x593 &  x614 &  x617 &  x620 &  x626 &  x635 &  x638 &  x641 &  x644 &  x647 &  x656 &  x665 &  x668 &  x698 &  x703 &  x719 &  x722 &  x728 &  x731 &  x734 &  x737 &  x740 &  x752 &  x761 &  x767 &  x776 &  x788 &  x794 &  x818 &  x821 &  x823 &  x827 &  x830 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x869 &  x875 &  x887 &  x896 &  x901 &  x905 &  x914 &  x917 &  x920 &  x926 &  x929 &  x938 &  x944 &  x950 &  x959 &  x962 &  x965 &  x974 &  x983 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1022 &  x1037 &  x1055 &  x1058 &  x1064 &  x1070 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1100 &  x1106 &  x1109 &  x1115 &  x1118 &  x1130 & ~x351 & ~x390 & ~x594 & ~x732 & ~x810 & ~x873 & ~x894 & ~x933;
assign c1268 =  x11 &  x14 &  x17 &  x23 &  x26 &  x29 &  x35 &  x41 &  x47 &  x56 &  x62 &  x86 &  x89 &  x95 &  x107 &  x113 &  x116 &  x131 &  x137 &  x140 &  x155 &  x158 &  x164 &  x170 &  x176 &  x188 &  x197 &  x203 &  x206 &  x215 &  x218 &  x221 &  x224 &  x242 &  x248 &  x275 &  x277 &  x281 &  x287 &  x290 &  x299 &  x314 &  x316 &  x323 &  x332 &  x341 &  x344 &  x355 &  x356 &  x365 &  x368 &  x371 &  x374 &  x377 &  x383 &  x392 &  x398 &  x404 &  x410 &  x428 &  x433 &  x446 &  x449 &  x461 &  x470 &  x473 &  x479 &  x485 &  x491 &  x494 &  x497 &  x503 &  x518 &  x524 &  x533 &  x545 &  x548 &  x554 &  x557 &  x563 &  x569 &  x575 &  x581 &  x592 &  x596 &  x599 &  x608 &  x623 &  x631 &  x638 &  x650 &  x656 &  x665 &  x668 &  x670 &  x671 &  x680 &  x692 &  x704 &  x713 &  x716 &  x725 &  x748 &  x749 &  x755 &  x758 &  x770 &  x776 &  x778 &  x785 &  x791 &  x797 &  x809 &  x821 &  x830 &  x836 &  x842 &  x851 &  x854 &  x860 &  x869 &  x872 &  x881 &  x884 &  x890 &  x893 &  x896 &  x920 &  x935 &  x944 &  x950 &  x953 &  x959 &  x989 &  x994 &  x995 &  x1001 &  x1013 &  x1016 &  x1031 &  x1033 &  x1034 &  x1037 &  x1040 &  x1043 &  x1052 &  x1055 &  x1064 &  x1076 &  x1082 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1111 &  x1115 &  x1121 &  x1127 &  x1130 & ~x606 & ~x645 & ~x663 & ~x703 & ~x741 & ~x780 & ~x781 & ~x819 & ~x820 & ~x858 & ~x898 & ~x900 & ~x975 & ~x978 & ~x1015 & ~x1017 & ~x1092;
assign c1270 =  x2 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x35 &  x38 &  x41 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x131 &  x134 &  x137 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x164 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x227 &  x233 &  x236 &  x242 &  x245 &  x248 &  x251 &  x254 &  x263 &  x266 &  x272 &  x274 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x317 &  x320 &  x323 &  x329 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x517 &  x518 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x556 &  x557 &  x566 &  x569 &  x572 &  x575 &  x578 &  x584 &  x590 &  x593 &  x595 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x629 &  x632 &  x635 &  x638 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x670 &  x671 &  x674 &  x676 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x704 &  x707 &  x709 &  x710 &  x713 &  x716 &  x719 &  x725 &  x727 &  x731 &  x734 &  x737 &  x740 &  x746 &  x748 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x793 &  x794 &  x796 &  x799 &  x800 &  x803 &  x805 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x827 &  x830 &  x833 &  x835 &  x836 &  x838 &  x839 &  x848 &  x851 &  x854 &  x857 &  x860 &  x866 &  x871 &  x872 &  x875 &  x877 &  x878 &  x881 &  x884 &  x890 &  x896 &  x899 &  x905 &  x908 &  x910 &  x911 &  x917 &  x923 &  x929 &  x932 &  x935 &  x938 &  x941 &  x947 &  x949 &  x950 &  x953 &  x955 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x309 & ~x822 & ~x939 & ~x978 & ~x1017;
assign c1272 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x155 &  x157 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x196 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x235 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x274 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x391 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x458 &  x461 &  x464 &  x467 &  x470 &  x476 &  x479 &  x482 &  x485 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x709 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x730 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x748 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x769 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x808 &  x809 &  x812 &  x815 &  x818 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x850 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130 & ~x162 & ~x201 & ~x309 & ~x744 & ~x783 & ~x822 & ~x900 & ~x939 & ~x942 & ~x981 & ~x1020 & ~x1059 & ~x1098;
assign c1274 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x413 &  x416 &  x419 &  x422 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x511 &  x512 &  x515 &  x518 &  x524 &  x527 &  x530 &  x536 &  x539 &  x542 &  x545 &  x548 &  x550 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x673 &  x674 &  x676 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x712 &  x713 &  x715 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x754 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x776 &  x779 &  x782 &  x785 &  x791 &  x793 &  x794 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x832 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x856 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x949 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x980 &  x983 &  x986 &  x988 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x639 & ~x678 & ~x702 & ~x741 & ~x780 & ~x819 & ~x858 & ~x897 & ~x936 & ~x975 & ~x1014 & ~x1017;
assign c1276 =  x23 &  x35 &  x41 &  x47 &  x50 &  x71 &  x98 &  x110 &  x113 &  x116 &  x119 &  x122 &  x128 &  x131 &  x137 &  x188 &  x191 &  x194 &  x199 &  x203 &  x215 &  x224 &  x230 &  x233 &  x260 &  x266 &  x278 &  x293 &  x299 &  x302 &  x305 &  x317 &  x344 &  x350 &  x353 &  x355 &  x362 &  x371 &  x374 &  x380 &  x383 &  x389 &  x394 &  x395 &  x397 &  x404 &  x422 &  x436 &  x449 &  x452 &  x474 &  x497 &  x514 &  x524 &  x545 &  x554 &  x569 &  x575 &  x581 &  x592 &  x599 &  x602 &  x614 &  x620 &  x631 &  x641 &  x644 &  x659 &  x670 &  x674 &  x707 &  x722 &  x725 &  x731 &  x749 &  x752 &  x767 &  x785 &  x791 &  x803 &  x806 &  x809 &  x824 &  x833 &  x836 &  x842 &  x844 &  x848 &  x860 &  x881 &  x890 &  x893 &  x899 &  x917 &  x923 &  x926 &  x929 &  x932 &  x938 &  x947 &  x955 &  x974 &  x1007 &  x1013 &  x1016 &  x1028 &  x1031 &  x1040 &  x1055 &  x1064 &  x1076 &  x1079 &  x1088 &  x1091 &  x1097 &  x1115 &  x1127 & ~x303 & ~x405 & ~x444 & ~x507 & ~x624 & ~x663 & ~x741 & ~x858 & ~x897;
assign c1278 =  x2 &  x5 &  x14 &  x26 &  x29 &  x41 &  x44 &  x50 &  x59 &  x65 &  x68 &  x74 &  x77 &  x83 &  x89 &  x95 &  x98 &  x101 &  x107 &  x110 &  x116 &  x128 &  x131 &  x134 &  x140 &  x143 &  x155 &  x176 &  x179 &  x182 &  x185 &  x194 &  x200 &  x203 &  x209 &  x212 &  x215 &  x218 &  x221 &  x227 &  x230 &  x239 &  x242 &  x245 &  x248 &  x254 &  x263 &  x266 &  x269 &  x281 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x314 &  x317 &  x320 &  x323 &  x326 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x353 &  x356 &  x359 &  x365 &  x374 &  x377 &  x383 &  x386 &  x394 &  x398 &  x410 &  x413 &  x416 &  x419 &  x425 &  x431 &  x433 &  x437 &  x440 &  x443 &  x446 &  x464 &  x472 &  x473 &  x476 &  x482 &  x488 &  x491 &  x497 &  x512 &  x518 &  x530 &  x536 &  x539 &  x548 &  x557 &  x581 &  x584 &  x587 &  x605 &  x608 &  x611 &  x614 &  x617 &  x623 &  x632 &  x650 &  x656 &  x662 &  x668 &  x671 &  x680 &  x686 &  x692 &  x701 &  x704 &  x707 &  x716 &  x722 &  x725 &  x731 &  x734 &  x737 &  x743 &  x746 &  x749 &  x758 &  x761 &  x764 &  x773 &  x782 &  x788 &  x791 &  x794 &  x803 &  x809 &  x815 &  x818 &  x830 &  x833 &  x842 &  x844 &  x848 &  x863 &  x872 &  x878 &  x881 &  x884 &  x887 &  x893 &  x896 &  x902 &  x905 &  x908 &  x917 &  x922 &  x932 &  x935 &  x947 &  x953 &  x961 &  x962 &  x968 &  x971 &  x977 &  x980 &  x992 &  x995 &  x1004 &  x1007 &  x1010 &  x1013 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1051 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1070 &  x1078 &  x1082 &  x1091 &  x1094 &  x1103 &  x1112 &  x1115 &  x1117 &  x1118 &  x1127 &  x1130 & ~x87 & ~x126 & ~x204 & ~x585 & ~x663 & ~x702 & ~x741 & ~x819 & ~x858 & ~x984;
assign c1280 =  x2 &  x5 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x41 &  x44 &  x53 &  x77 &  x95 &  x101 &  x110 &  x113 &  x116 &  x119 &  x125 &  x134 &  x137 &  x149 &  x152 &  x161 &  x167 &  x176 &  x179 &  x182 &  x188 &  x191 &  x200 &  x203 &  x209 &  x215 &  x218 &  x221 &  x227 &  x230 &  x239 &  x242 &  x245 &  x251 &  x257 &  x260 &  x266 &  x269 &  x272 &  x275 &  x277 &  x281 &  x290 &  x296 &  x305 &  x308 &  x314 &  x317 &  x320 &  x326 &  x332 &  x335 &  x344 &  x350 &  x355 &  x356 &  x359 &  x371 &  x374 &  x386 &  x389 &  x392 &  x394 &  x395 &  x398 &  x404 &  x410 &  x422 &  x425 &  x428 &  x431 &  x434 &  x446 &  x449 &  x458 &  x461 &  x464 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x497 &  x500 &  x503 &  x509 &  x512 &  x515 &  x533 &  x539 &  x542 &  x545 &  x548 &  x551 &  x572 &  x575 &  x578 &  x593 &  x596 &  x599 &  x614 &  x626 &  x632 &  x644 &  x659 &  x662 &  x665 &  x668 &  x671 &  x677 &  x680 &  x683 &  x701 &  x704 &  x710 &  x716 &  x722 &  x725 &  x728 &  x733 &  x739 &  x740 &  x746 &  x758 &  x761 &  x764 &  x776 &  x779 &  x785 &  x791 &  x797 &  x800 &  x803 &  x809 &  x812 &  x815 &  x817 &  x821 &  x824 &  x832 &  x839 &  x844 &  x851 &  x854 &  x856 &  x860 &  x866 &  x871 &  x872 &  x881 &  x883 &  x890 &  x895 &  x902 &  x908 &  x910 &  x914 &  x916 &  x917 &  x920 &  x922 &  x926 &  x932 &  x934 &  x935 &  x944 &  x947 &  x949 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x977 &  x980 &  x998 &  x1016 &  x1019 &  x1031 &  x1034 &  x1040 &  x1049 &  x1052 &  x1055 &  x1058 &  x1073 &  x1079 &  x1082 &  x1085 &  x1100 &  x1103 &  x1115 &  x1121 &  x1124 &  x1127 & ~x303 & ~x447 & ~x486 & ~x525 & ~x624 & ~x663 & ~x702 & ~x858 & ~x861 & ~x900 & ~x939 & ~x975 & ~x978;
assign c1282 =  x11 &  x38 &  x41 &  x65 &  x98 &  x104 &  x116 &  x119 &  x122 &  x131 &  x140 &  x164 &  x173 &  x176 &  x185 &  x212 &  x215 &  x221 &  x239 &  x254 &  x272 &  x275 &  x290 &  x305 &  x308 &  x317 &  x329 &  x335 &  x341 &  x344 &  x359 &  x371 &  x376 &  x388 &  x395 &  x409 &  x415 &  x422 &  x434 &  x443 &  x452 &  x470 &  x476 &  x488 &  x509 &  x512 &  x524 &  x527 &  x548 &  x560 &  x575 &  x581 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x641 &  x650 &  x662 &  x665 &  x674 &  x683 &  x695 &  x698 &  x716 &  x731 &  x746 &  x749 &  x752 &  x764 &  x776 &  x779 &  x782 &  x797 &  x824 &  x827 &  x842 &  x845 &  x878 &  x881 &  x896 &  x899 &  x905 &  x914 &  x929 &  x935 &  x941 &  x944 &  x959 &  x971 &  x974 &  x977 &  x980 &  x983 &  x992 &  x1004 &  x1013 &  x1016 &  x1018 &  x1028 &  x1034 &  x1040 &  x1046 &  x1061 &  x1064 &  x1088 &  x1091 &  x1094 &  x1097 &  x1109 &  x1118 &  x1121 & ~x198 & ~x273 & ~x432 & ~x438 & ~x738 & ~x846 & ~x954 & ~x990;
assign c1284 =  x2 &  x5 &  x8 &  x11 &  x17 &  x23 &  x29 &  x32 &  x38 &  x41 &  x47 &  x53 &  x56 &  x59 &  x68 &  x71 &  x74 &  x80 &  x83 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x134 &  x137 &  x140 &  x143 &  x146 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x185 &  x191 &  x197 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x227 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x254 &  x257 &  x263 &  x269 &  x275 &  x278 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x308 &  x314 &  x320 &  x323 &  x326 &  x329 &  x335 &  x338 &  x341 &  x344 &  x353 &  x356 &  x359 &  x362 &  x368 &  x371 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x418 &  x419 &  x422 &  x428 &  x431 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x464 &  x467 &  x470 &  x476 &  x479 &  x481 &  x482 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x511 &  x515 &  x520 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x542 &  x548 &  x550 &  x551 &  x554 &  x557 &  x558 &  x559 &  x560 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x596 &  x598 &  x602 &  x605 &  x608 &  x614 &  x623 &  x632 &  x635 &  x637 &  x638 &  x641 &  x647 &  x656 &  x659 &  x671 &  x674 &  x676 &  x680 &  x689 &  x692 &  x695 &  x698 &  x704 &  x707 &  x710 &  x713 &  x715 &  x716 &  x722 &  x725 &  x731 &  x734 &  x737 &  x743 &  x746 &  x749 &  x758 &  x761 &  x767 &  x770 &  x776 &  x791 &  x794 &  x797 &  x800 &  x806 &  x809 &  x815 &  x818 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x869 &  x875 &  x878 &  x884 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x917 &  x920 &  x926 &  x929 &  x932 &  x935 &  x941 &  x944 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x971 &  x974 &  x980 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1058 &  x1061 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1100 &  x1106 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 &  x1130 & ~x741 & ~x780 & ~x858 & ~x936 & ~x975;
assign c1286 =  x2 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x53 &  x56 &  x68 &  x71 &  x74 &  x77 &  x80 &  x92 &  x98 &  x113 &  x116 &  x122 &  x128 &  x131 &  x137 &  x140 &  x143 &  x149 &  x152 &  x154 &  x158 &  x164 &  x167 &  x170 &  x176 &  x182 &  x185 &  x188 &  x191 &  x197 &  x200 &  x203 &  x206 &  x209 &  x218 &  x224 &  x227 &  x233 &  x239 &  x242 &  x245 &  x251 &  x257 &  x260 &  x263 &  x269 &  x278 &  x284 &  x296 &  x305 &  x311 &  x317 &  x326 &  x332 &  x335 &  x344 &  x350 &  x353 &  x362 &  x365 &  x368 &  x374 &  x377 &  x389 &  x392 &  x398 &  x401 &  x404 &  x410 &  x413 &  x419 &  x422 &  x425 &  x434 &  x443 &  x449 &  x455 &  x458 &  x464 &  x473 &  x476 &  x479 &  x485 &  x491 &  x494 &  x497 &  x500 &  x503 &  x509 &  x512 &  x515 &  x518 &  x530 &  x533 &  x542 &  x548 &  x554 &  x557 &  x560 &  x563 &  x569 &  x572 &  x581 &  x584 &  x587 &  x590 &  x593 &  x599 &  x602 &  x608 &  x611 &  x617 &  x620 &  x623 &  x626 &  x629 &  x635 &  x641 &  x644 &  x656 &  x662 &  x665 &  x671 &  x695 &  x701 &  x707 &  x710 &  x713 &  x719 &  x722 &  x734 &  x737 &  x740 &  x743 &  x746 &  x752 &  x773 &  x794 &  x803 &  x806 &  x815 &  x818 &  x821 &  x827 &  x833 &  x836 &  x845 &  x857 &  x863 &  x866 &  x869 &  x872 &  x878 &  x884 &  x887 &  x893 &  x896 &  x899 &  x911 &  x914 &  x923 &  x926 &  x929 &  x932 &  x941 &  x944 &  x959 &  x965 &  x968 &  x974 &  x977 &  x980 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1019 &  x1025 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1070 &  x1073 &  x1076 &  x1091 &  x1094 &  x1100 &  x1112 &  x1130 & ~x171 & ~x324 & ~x333 & ~x372 & ~x441 & ~x891 & ~x948 & ~x1107;
assign c1288 =  x5 &  x26 &  x35 &  x47 &  x56 &  x62 &  x65 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x107 &  x113 &  x116 &  x119 &  x134 &  x143 &  x155 &  x161 &  x170 &  x173 &  x176 &  x185 &  x188 &  x197 &  x206 &  x224 &  x227 &  x230 &  x233 &  x245 &  x251 &  x254 &  x263 &  x269 &  x272 &  x305 &  x308 &  x344 &  x347 &  x359 &  x362 &  x365 &  x374 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x404 &  x407 &  x422 &  x425 &  x428 &  x443 &  x467 &  x476 &  x479 &  x485 &  x488 &  x503 &  x518 &  x521 &  x524 &  x530 &  x533 &  x551 &  x554 &  x557 &  x563 &  x566 &  x575 &  x578 &  x584 &  x587 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x626 &  x629 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x662 &  x665 &  x668 &  x680 &  x686 &  x689 &  x698 &  x701 &  x710 &  x713 &  x716 &  x728 &  x731 &  x734 &  x740 &  x743 &  x752 &  x758 &  x761 &  x764 &  x767 &  x773 &  x776 &  x778 &  x779 &  x788 &  x793 &  x794 &  x803 &  x806 &  x809 &  x818 &  x824 &  x839 &  x845 &  x848 &  x851 &  x856 &  x860 &  x869 &  x871 &  x872 &  x877 &  x881 &  x887 &  x890 &  x893 &  x895 &  x899 &  x902 &  x905 &  x910 &  x914 &  x916 &  x920 &  x923 &  x926 &  x947 &  x953 &  x956 &  x968 &  x983 &  x986 &  x989 &  x992 &  x994 &  x998 &  x1001 &  x1010 &  x1013 &  x1019 &  x1022 &  x1031 &  x1040 &  x1049 &  x1055 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1112 &  x1115 &  x1121 &  x1124 &  x1129 & ~x426 & ~x465 & ~x780 & ~x981 & ~x1059 & ~x1098;
assign c1290 =  x2 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x70 &  x71 &  x74 &  x76 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x101 &  x107 &  x109 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x136 &  x137 &  x140 &  x143 &  x146 &  x148 &  x149 &  x152 &  x154 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x175 &  x179 &  x182 &  x185 &  x187 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x214 &  x215 &  x218 &  x221 &  x224 &  x226 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x253 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x298 &  x299 &  x302 &  x305 &  x308 &  x310 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x641 &  x644 &  x647 &  x650 &  x656 &  x659 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x943 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x977 &  x980 &  x982 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1021 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x156 & ~x195 & ~x234 & ~x273 & ~x276 & ~x879;
assign c1292 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x104 &  x110 &  x113 &  x116 &  x119 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x203 &  x206 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x251 &  x254 &  x257 &  x260 &  x263 &  x269 &  x271 &  x272 &  x278 &  x281 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x310 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x359 &  x362 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x389 &  x392 &  x395 &  x398 &  x404 &  x406 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x445 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x484 &  x485 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x524 &  x527 &  x533 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x584 &  x586 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x625 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x668 &  x671 &  x674 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x779 &  x782 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x827 &  x833 &  x836 &  x839 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x890 &  x893 &  x896 &  x899 &  x901 &  x902 &  x905 &  x908 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x941 &  x944 &  x950 &  x953 &  x959 &  x962 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x234 & ~x273 & ~x516 & ~x654 & ~x655 & ~x693;
assign c1294 =  x50 &  x62 &  x77 &  x86 &  x95 &  x101 &  x110 &  x116 &  x131 &  x134 &  x137 &  x140 &  x149 &  x182 &  x188 &  x194 &  x200 &  x212 &  x221 &  x260 &  x278 &  x302 &  x305 &  x335 &  x344 &  x356 &  x401 &  x404 &  x410 &  x419 &  x425 &  x434 &  x446 &  x452 &  x476 &  x484 &  x488 &  x500 &  x509 &  x518 &  x523 &  x554 &  x557 &  x562 &  x584 &  x593 &  x602 &  x608 &  x620 &  x650 &  x671 &  x695 &  x698 &  x701 &  x713 &  x719 &  x725 &  x731 &  x737 &  x740 &  x773 &  x794 &  x803 &  x809 &  x815 &  x818 &  x824 &  x830 &  x833 &  x836 &  x845 &  x860 &  x866 &  x869 &  x884 &  x890 &  x893 &  x905 &  x908 &  x911 &  x923 &  x929 &  x935 &  x938 &  x941 &  x947 &  x979 &  x1001 &  x1018 &  x1025 &  x1049 &  x1061 &  x1073 &  x1082 &  x1085 &  x1091 &  x1099 &  x1100 &  x1112 &  x1115 & ~x633 & ~x870 & ~x990 & ~x1068 & ~x1086;
assign c1296 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x359 &  x362 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x406 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x440 &  x443 &  x445 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x542 &  x545 &  x548 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x644 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x784 &  x785 &  x788 &  x791 &  x797 &  x800 &  x803 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x865 &  x866 &  x869 &  x872 &  x878 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x904 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 & ~x435 & ~x474 & ~x576 & ~x615 & ~x616 & ~x654 & ~x693 & ~x732 & ~x756 & ~x795;
assign c1298 =  x2 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x29 &  x32 &  x41 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x104 &  x107 &  x113 &  x119 &  x122 &  x125 &  x128 &  x131 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x191 &  x194 &  x197 &  x203 &  x206 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x257 &  x260 &  x263 &  x266 &  x269 &  x275 &  x278 &  x281 &  x284 &  x290 &  x293 &  x296 &  x299 &  x302 &  x308 &  x311 &  x314 &  x320 &  x329 &  x332 &  x341 &  x344 &  x350 &  x353 &  x356 &  x368 &  x371 &  x374 &  x377 &  x386 &  x392 &  x394 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x433 &  x434 &  x436 &  x437 &  x439 &  x440 &  x443 &  x452 &  x455 &  x458 &  x461 &  x464 &  x472 &  x475 &  x476 &  x479 &  x482 &  x485 &  x494 &  x497 &  x500 &  x503 &  x506 &  x512 &  x514 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x542 &  x548 &  x551 &  x553 &  x554 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x584 &  x587 &  x590 &  x593 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x680 &  x686 &  x689 &  x695 &  x698 &  x704 &  x707 &  x710 &  x713 &  x715 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x794 &  x800 &  x806 &  x818 &  x821 &  x824 &  x830 &  x836 &  x842 &  x845 &  x848 &  x854 &  x857 &  x860 &  x866 &  x869 &  x875 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x905 &  x908 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x968 &  x971 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1103 &  x1106 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x489 & ~x528 & ~x529 & ~x567;
assign c11 = ~x59 & ~x365;
assign c13 =  x46 &  x730 &  x941 &  x1013 & ~x258 & ~x297 & ~x675;
assign c15 =  x48 &  x312;
assign c17 =  x936 & ~x796 & ~x904;
assign c19 =  x334 &  x589 & ~x156 & ~x669 & ~x747;
assign c113 =  x53 &  x353 &  x394 &  x410 &  x443 &  x472 &  x536 &  x542 &  x602 &  x679 &  x695 &  x887 &  x896 &  x986 &  x1016 &  x1025 & ~x63 & ~x474 & ~x822 & ~x900;
assign c115 =  x583 & ~x387 & ~x570 & ~x687;
assign c117 =  x38 &  x95 &  x98 &  x265 &  x269 &  x368 &  x397 &  x436 &  x500 &  x521 &  x734 &  x827 &  x836 &  x857 &  x887 &  x899 &  x956 &  x962 & ~x351 & ~x726 & ~x903 & ~x942 & ~x981 & ~x1098;
assign c119 =  x514 &  x703 &  x742 & ~x468 & ~x1060;
assign c121 = ~x710;
assign c123 =  x624 & ~x865;
assign c125 =  x158 &  x317 &  x332 &  x458 &  x470 &  x535 &  x665 &  x695 &  x770 &  x866 &  x1060 &  x1070 &  x1124 & ~x672 & ~x1053;
assign c127 =  x67 &  x184 &  x476 &  x560 &  x574 &  x622 &  x685 &  x724 &  x860 &  x895 &  x931;
assign c129 =  x990;
assign c131 =  x289 &  x320 &  x328 &  x357 &  x449 &  x605 &  x674 &  x794;
assign c133 =  x77 &  x262 &  x691 &  x703 & ~x715;
assign c135 =  x6 &  x892 &  x928;
assign c137 = ~x514;
assign c139 = ~x787 & ~x801 & ~x1011 & ~x1117;
assign c141 =  x703 &  x738 &  x739 & ~x204 & ~x669;
assign c143 =  x717 &  x912 &  x1087;
assign c145 =  x756 &  x912 & ~x649;
assign c147 =  x428 &  x457 &  x620 &  x803 & ~x447 & ~x559;
assign c149 =  x46 &  x53 &  x212 &  x263 &  x269 &  x305 &  x457 &  x554 &  x902 &  x923 &  x932 &  x1052 &  x1061 &  x1091 & ~x327 & ~x861 & ~x885;
assign c151 =  x718 &  x1030 &  x1105 & ~x784;
assign c153 =  x207 &  x574 &  x613 &  x1108;
assign c155 =  x7 &  x41 &  x392 &  x739 &  x857 &  x872 &  x977 &  x1058 &  x1070 &  x1099 &  x1117 & ~x0 & ~x480 & ~x516;
assign c157 = ~x596;
assign c159 =  x754 &  x967 & ~x219 & ~x258 & ~x453 & ~x741 & ~x744;
assign c161 =  x241 & ~x156 & ~x525 & ~x597 & ~x1090;
assign c163 = ~x359 & ~x560 & ~x563;
assign c165 =  x87 &  x165 &  x753;
assign c167 = ~x272;
assign c169 =  x477 &  x624;
assign c171 =  x424 &  x529 &  x1033 & ~x159 & ~x486;
assign c173 =  x385 & ~x259 & ~x1080;
assign c175 = ~x842;
assign c177 =  x2 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x44 &  x50 &  x56 &  x59 &  x65 &  x74 &  x77 &  x83 &  x92 &  x95 &  x98 &  x107 &  x113 &  x116 &  x119 &  x122 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x155 &  x158 &  x161 &  x164 &  x167 &  x173 &  x179 &  x182 &  x185 &  x191 &  x194 &  x197 &  x209 &  x212 &  x215 &  x218 &  x224 &  x230 &  x242 &  x245 &  x248 &  x251 &  x263 &  x266 &  x272 &  x275 &  x278 &  x284 &  x287 &  x296 &  x299 &  x302 &  x305 &  x308 &  x317 &  x320 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x395 &  x398 &  x401 &  x404 &  x410 &  x413 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x451 &  x452 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x485 &  x488 &  x491 &  x494 &  x497 &  x506 &  x509 &  x512 &  x518 &  x521 &  x527 &  x533 &  x536 &  x542 &  x548 &  x551 &  x557 &  x560 &  x563 &  x566 &  x578 &  x581 &  x584 &  x587 &  x589 &  x590 &  x596 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x626 &  x628 &  x629 &  x632 &  x638 &  x644 &  x647 &  x650 &  x653 &  x656 &  x665 &  x668 &  x671 &  x683 &  x686 &  x689 &  x692 &  x695 &  x701 &  x704 &  x707 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x739 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x764 &  x767 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x833 &  x836 &  x845 &  x848 &  x851 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x878 &  x881 &  x884 &  x893 &  x896 &  x899 &  x902 &  x908 &  x911 &  x914 &  x920 &  x923 &  x926 &  x929 &  x932 &  x941 &  x944 &  x950 &  x956 &  x959 &  x965 &  x968 &  x977 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1028 &  x1034 &  x1040 &  x1046 &  x1049 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1079 &  x1082 &  x1088 &  x1094 &  x1097 &  x1100 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 &  x1130 & ~x522 & ~x669 & ~x693;
assign c179 =  x185 &  x280 &  x311 &  x319 &  x528 &  x529 &  x931 & ~x243;
assign c181 =  x46 &  x59 &  x71 &  x224 &  x284 &  x305 &  x322 &  x398 &  x434 &  x485 &  x569 &  x581 &  x587 &  x647 &  x695 &  x722 &  x788 &  x872 &  x935 &  x1031 &  x1043 &  x1091 & ~x27 & ~x39 & ~x300 & ~x306 & ~x672;
assign c183 = ~x530;
assign c185 =  x347 &  x470 &  x480 &  x523 &  x560 &  x647 &  x668 &  x734 &  x763 &  x764 &  x785 &  x788 &  x853 &  x893 &  x1049 &  x1076;
assign c187 =  x270 &  x349 &  x439 &  x454 & ~x945;
assign c189 = ~x3 & ~x331 & ~x441 & ~x672;
assign c191 =  x5 &  x7 &  x17 &  x20 &  x44 &  x56 &  x62 &  x68 &  x71 &  x74 &  x77 &  x89 &  x98 &  x107 &  x110 &  x116 &  x122 &  x128 &  x131 &  x140 &  x170 &  x173 &  x209 &  x212 &  x215 &  x218 &  x242 &  x245 &  x260 &  x263 &  x272 &  x278 &  x296 &  x311 &  x314 &  x320 &  x323 &  x326 &  x335 &  x338 &  x353 &  x362 &  x380 &  x383 &  x389 &  x392 &  x407 &  x413 &  x416 &  x419 &  x425 &  x428 &  x437 &  x443 &  x458 &  x464 &  x467 &  x503 &  x506 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x533 &  x539 &  x551 &  x581 &  x590 &  x596 &  x605 &  x611 &  x628 &  x629 &  x632 &  x635 &  x638 &  x656 &  x667 &  x668 &  x680 &  x692 &  x719 &  x740 &  x746 &  x749 &  x773 &  x782 &  x785 &  x788 &  x803 &  x812 &  x821 &  x824 &  x845 &  x851 &  x881 &  x911 &  x917 &  x920 &  x929 &  x944 &  x956 &  x959 &  x965 &  x971 &  x980 &  x983 &  x992 &  x1001 &  x1004 &  x1025 &  x1028 &  x1040 &  x1052 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1085 &  x1094 &  x1106 &  x1109 &  x1121 &  x1130 & ~x561 & ~x639 & ~x669 & ~x792;
assign c193 =  x424 &  x518 &  x1091 & ~x220 & ~x906 & ~x1080 & ~x1119;
assign c195 = ~x410;
assign c197 =  x840 & ~x234 & ~x483;
assign c199 =  x13 &  x26 &  x38 &  x41 &  x50 &  x125 &  x149 &  x173 &  x209 &  x248 &  x319 &  x332 &  x392 &  x419 &  x451 &  x491 &  x521 &  x527 &  x529 &  x539 &  x653 &  x662 &  x692 &  x707 &  x749 &  x806 &  x839 &  x848 &  x875 &  x896 &  x911 &  x941 &  x950 &  x989 &  x1028 & ~x792 & ~x831;
assign c1101 =  x154 &  x344 &  x544 &  x616 &  x676 &  x1006 &  x1111 & ~x132;
assign c1103 =  x656 &  x776 & ~x57 & ~x292 & ~x331 & ~x447 & ~x564;
assign c1105 = ~x78 & ~x786 & ~x1057;
assign c1107 =  x289 &  x295 &  x396 & ~x636;
assign c1109 =  x629 &  x705 &  x1079 & ~x393 & ~x715;
assign c1111 = ~x326;
assign c1113 = ~x428;
assign c1115 =  x7 &  x59 &  x344 &  x377 &  x475 &  x863 &  x932 &  x1033 &  x1046 &  x1052 &  x1058 & ~x240 & ~x249 & ~x345;
assign c1117 =  x298 &  x1014 & ~x717 & ~x835;
assign c1119 = ~x436 & ~x784;
assign c1121 =  x7 &  x46 &  x124 &  x840 &  x1036;
assign c1123 =  x204 & ~x358;
assign c1125 =  x343 &  x409 &  x439 &  x625 &  x661 & ~x747;
assign c1127 =  x432 &  x471 & ~x670;
assign c1129 =  x602 &  x620 &  x707 &  x941 & ~x39 & ~x327 & ~x669 & ~x939;
assign c1131 =  x87 &  x234 &  x1027 & ~x220;
assign c1133 =  x477 & ~x351 & ~x384 & ~x390 & ~x933;
assign c1135 =  x574 &  x724 &  x763 &  x814 &  x841 & ~x321 & ~x429;
assign c1137 =  x198 & ~x93 & ~x250 & ~x745;
assign c1141 = ~x893;
assign c1143 =  x625 &  x733 & ~x600 & ~x631;
assign c1145 =  x26 &  x59 &  x68 &  x71 &  x101 &  x197 &  x221 &  x242 &  x362 &  x545 &  x596 &  x605 &  x629 &  x659 &  x707 &  x779 &  x911 &  x938 &  x944 &  x1013 &  x1040 &  x1070 &  x1087 &  x1097 &  x1121 & ~x522 & ~x531 & ~x648 & ~x687;
assign c1147 =  x47 &  x260 &  x284 &  x360 &  x547 &  x703 &  x752 &  x830 &  x884 &  x896 &  x1007 & ~x453;
assign c1149 =  x5 &  x8 &  x17 &  x23 &  x44 &  x56 &  x68 &  x71 &  x77 &  x89 &  x104 &  x119 &  x161 &  x200 &  x203 &  x227 &  x230 &  x251 &  x257 &  x275 &  x278 &  x287 &  x293 &  x308 &  x344 &  x368 &  x374 &  x401 &  x431 &  x440 &  x470 &  x494 &  x500 &  x515 &  x521 &  x524 &  x533 &  x554 &  x575 &  x578 &  x629 &  x641 &  x659 &  x665 &  x671 &  x677 &  x698 &  x710 &  x719 &  x728 &  x731 &  x770 &  x797 &  x806 &  x821 &  x824 &  x833 &  x836 &  x845 &  x866 &  x869 &  x890 &  x935 &  x938 &  x950 &  x977 &  x989 &  x992 &  x995 &  x1013 &  x1016 &  x1022 &  x1025 &  x1034 &  x1043 &  x1046 &  x1064 &  x1070 &  x1112 & ~x0 & ~x630 & ~x861 & ~x939;
assign c1151 =  x28 &  x248 &  x278 &  x314 &  x418 &  x613 &  x632 &  x696 &  x853 &  x1049 &  x1090;
assign c1153 =  x490 &  x580 & ~x132 & ~x976 & ~x1053;
assign c1155 =  x379 & ~x403 & ~x555;
assign c1157 =  x236 &  x530 &  x590 &  x620 &  x638 &  x692 &  x710 &  x740 &  x848 &  x872 &  x920 &  x1111 & ~x288 & ~x445 & ~x474 & ~x897 & ~x936;
assign c1159 =  x537 &  x857 & ~x93 & ~x906 & ~x1074;
assign c1161 = ~x827;
assign c1163 = ~x722;
assign c1165 =  x218 &  x418 &  x514 &  x745 &  x758 &  x976 & ~x198 & ~x639 & ~x747;
assign c1167 =  x1029 & ~x747;
assign c1169 =  x7 &  x23 &  x275 &  x688 &  x722 &  x733 &  x802 &  x821 & ~x555 & ~x885;
assign c1171 = ~x281;
assign c1173 =  x241 &  x287 &  x305 &  x622 &  x1107;
assign c1175 =  x204 & ~x0 & ~x261;
assign c1177 = ~x935;
assign c1179 =  x23 &  x35 &  x65 &  x173 &  x206 &  x251 &  x287 &  x323 &  x374 &  x377 &  x386 &  x401 &  x407 &  x413 &  x422 &  x464 &  x476 &  x482 &  x500 &  x512 &  x530 &  x551 &  x554 &  x572 &  x704 &  x737 &  x764 &  x773 &  x779 &  x788 &  x818 &  x824 &  x830 &  x833 &  x944 &  x1049 &  x1052 &  x1055 & ~x273 & ~x786 & ~x834 & ~x835 & ~x873 & ~x942 & ~x981;
assign c1181 =  x172 &  x307 &  x446 &  x622 &  x662 &  x739 &  x923 & ~x972 & ~x1059;
assign c1183 = ~x1041 & ~x1117;
assign c1185 =  x165;
assign c1187 =  x2 &  x5 &  x14 &  x17 &  x20 &  x23 &  x29 &  x32 &  x41 &  x44 &  x46 &  x47 &  x50 &  x53 &  x62 &  x65 &  x68 &  x71 &  x74 &  x83 &  x89 &  x92 &  x95 &  x104 &  x107 &  x113 &  x116 &  x119 &  x122 &  x125 &  x131 &  x134 &  x146 &  x149 &  x164 &  x167 &  x176 &  x179 &  x182 &  x185 &  x188 &  x197 &  x212 &  x215 &  x224 &  x227 &  x230 &  x233 &  x236 &  x242 &  x248 &  x251 &  x257 &  x266 &  x278 &  x281 &  x284 &  x287 &  x290 &  x296 &  x302 &  x311 &  x317 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x344 &  x350 &  x353 &  x359 &  x362 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x404 &  x407 &  x410 &  x419 &  x422 &  x425 &  x428 &  x434 &  x440 &  x452 &  x458 &  x464 &  x467 &  x473 &  x476 &  x479 &  x485 &  x488 &  x491 &  x494 &  x497 &  x506 &  x512 &  x515 &  x521 &  x524 &  x530 &  x533 &  x535 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x563 &  x568 &  x569 &  x574 &  x575 &  x581 &  x596 &  x599 &  x602 &  x605 &  x608 &  x614 &  x616 &  x617 &  x620 &  x626 &  x629 &  x632 &  x638 &  x647 &  x650 &  x653 &  x655 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x701 &  x704 &  x716 &  x728 &  x737 &  x743 &  x755 &  x758 &  x761 &  x764 &  x767 &  x773 &  x776 &  x779 &  x785 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x818 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x896 &  x899 &  x923 &  x926 &  x932 &  x938 &  x953 &  x956 &  x965 &  x968 &  x974 &  x980 &  x983 &  x986 &  x989 &  x992 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1034 &  x1049 &  x1058 &  x1061 &  x1064 &  x1067 &  x1076 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x756 & ~x834 & ~x870 & ~x873;
assign c1189 = ~x728;
assign c1191 =  x29 &  x89 &  x104 &  x164 &  x212 &  x305 &  x332 &  x383 &  x392 &  x395 &  x412 &  x451 &  x490 &  x500 &  x506 &  x512 &  x518 &  x529 &  x566 &  x572 &  x584 &  x596 &  x608 &  x660 &  x661 &  x695 &  x788 &  x860 &  x878 &  x1004;
assign c1193 =  x274 &  x739 &  x1026 & ~x474;
assign c1195 =  x382 & ~x805 & ~x979;
assign c1197 =  x38 &  x62 &  x68 &  x74 &  x77 &  x86 &  x128 &  x131 &  x134 &  x161 &  x179 &  x188 &  x209 &  x215 &  x224 &  x254 &  x263 &  x269 &  x275 &  x278 &  x287 &  x290 &  x293 &  x332 &  x338 &  x341 &  x362 &  x386 &  x404 &  x437 &  x497 &  x503 &  x512 &  x518 &  x521 &  x527 &  x539 &  x545 &  x548 &  x551 &  x587 &  x608 &  x614 &  x622 &  x629 &  x683 &  x692 &  x731 &  x752 &  x761 &  x782 &  x791 &  x803 &  x827 &  x830 &  x842 &  x845 &  x848 &  x854 &  x857 &  x875 &  x881 &  x884 &  x890 &  x893 &  x902 &  x926 &  x941 &  x944 &  x951 &  x983 &  x990 &  x1030 &  x1031 &  x1040 &  x1048 &  x1052 &  x1061 &  x1070 &  x1079 &  x1097 &  x1100 &  x1112 &  x1121 &  x1127;
assign c1199 =  x820 & ~x40 & ~x378 & ~x573 & ~x981;
assign c1201 =  x351 &  x1021 &  x1077;
assign c1203 =  x778 & ~x492 & ~x571 & ~x669;
assign c1205 =  x859 &  x1069 & ~x687 & ~x726 & ~x864;
assign c1207 =  x87 &  x967 & ~x181;
assign c1209 = ~x297 & ~x357 & ~x667 & ~x706;
assign c1211 =  x278 &  x281 &  x679 &  x878 &  x1021 &  x1105 & ~x474 & ~x783;
assign c1213 =  x237 & ~x96 & ~x280 & ~x288;
assign c1215 =  x82 &  x970 &  x1028 &  x1118 & ~x351 & ~x648 & ~x687;
assign c1217 = ~x784;
assign c1219 = ~x533;
assign c1221 =  x45 &  x908 & ~x222 & ~x822 & ~x861 & ~x900;
assign c1223 =  x46 &  x47 &  x109 &  x185 &  x227 &  x251 &  x275 &  x307 &  x325 &  x403 &  x655 &  x707 &  x758 &  x839 &  x881 &  x944 &  x1085 &  x1097 &  x1115;
assign c1225 =  x499 &  x913 &  x1027 & ~x15 & ~x93 & ~x915;
assign c1227 =  x1029 &  x1068 & ~x922;
assign c1229 =  x167 &  x305 &  x344 &  x358 &  x397 &  x572 &  x605 &  x734 &  x860 &  x884 &  x1076 & ~x159 & ~x273 & ~x312 & ~x906 & ~x1020 & ~x1098;
assign c1231 =  x1105 & ~x433 & ~x945;
assign c1233 = ~x297 & ~x376 & ~x885;
assign c1235 = ~x839;
assign c1237 =  x627 &  x702;
assign c1239 =  x757 &  x835 & ~x273 & ~x570 & ~x726 & ~x882 & ~x900;
assign c1241 = ~x436 & ~x667 & ~x745;
assign c1243 =  x35 &  x38 &  x68 &  x80 &  x92 &  x95 &  x161 &  x191 &  x193 &  x206 &  x239 &  x260 &  x290 &  x302 &  x326 &  x332 &  x389 &  x425 &  x440 &  x452 &  x461 &  x464 &  x485 &  x538 &  x548 &  x551 &  x572 &  x641 &  x647 &  x653 &  x656 &  x674 &  x680 &  x683 &  x707 &  x710 &  x716 &  x737 &  x755 &  x779 &  x785 &  x815 &  x863 &  x899 &  x905 &  x929 &  x941 &  x965 &  x968 &  x974 &  x995 &  x1030 &  x1031 &  x1043 &  x1064 &  x1085 &  x1097 &  x1109 & ~x39 & ~x366;
assign c1245 =  x403 & ~x93 & ~x267 & ~x366;
assign c1247 =  x165 &  x312 & ~x891;
assign c1249 =  x265 &  x457 &  x505 &  x969 & ~x903;
assign c1251 = ~x554;
assign c1253 =  x717 &  x1012 & ~x783;
assign c1255 =  x353 &  x455 &  x466 &  x470 &  x575 &  x767 & ~x525 & ~x561 & ~x604;
assign c1257 = ~x77;
assign c1259 =  x45 &  x1077 & ~x258;
assign c1261 = ~x525 & ~x748;
assign c1263 =  x7 & ~x16 & ~x55 & ~x106;
assign c1265 = ~x965;
assign c1267 =  x5 &  x26 &  x62 &  x77 &  x92 &  x101 &  x107 &  x122 &  x128 &  x140 &  x155 &  x161 &  x173 &  x176 &  x179 &  x182 &  x188 &  x191 &  x197 &  x200 &  x203 &  x221 &  x227 &  x233 &  x236 &  x242 &  x248 &  x293 &  x308 &  x311 &  x323 &  x335 &  x347 &  x353 &  x365 &  x374 &  x377 &  x398 &  x407 &  x410 &  x428 &  x452 &  x473 &  x497 &  x503 &  x518 &  x521 &  x548 &  x554 &  x560 &  x566 &  x578 &  x587 &  x590 &  x596 &  x605 &  x608 &  x617 &  x620 &  x626 &  x632 &  x641 &  x665 &  x668 &  x680 &  x681 &  x683 &  x704 &  x707 &  x710 &  x713 &  x719 &  x734 &  x739 &  x758 &  x764 &  x779 &  x782 &  x785 &  x800 &  x806 &  x809 &  x818 &  x824 &  x827 &  x830 &  x836 &  x839 &  x856 &  x905 &  x908 &  x911 &  x926 &  x935 &  x938 &  x941 &  x944 &  x953 &  x956 &  x965 &  x977 &  x1001 &  x1004 &  x1007 &  x1010 &  x1012 &  x1019 &  x1025 &  x1028 &  x1037 &  x1043 &  x1046 &  x1052 &  x1055 &  x1070 &  x1076 &  x1079 &  x1091 &  x1103 &  x1106 &  x1130 & ~x438;
assign c1269 =  x739 & ~x42 & ~x370 & ~x672;
assign c1271 =  x652 & ~x604 & ~x633;
assign c1273 =  x205 &  x725 & ~x183 & ~x438 & ~x741 & ~x783 & ~x1047 & ~x1107;
assign c1275 =  x242 &  x550 &  x578 &  x710 &  x874 &  x998 & ~x117 & ~x150 & ~x183 & ~x339 & ~x366;
assign c1277 =  x44 &  x49 &  x125 &  x127 &  x152 &  x176 &  x200 &  x236 &  x245 &  x254 &  x266 &  x269 &  x275 &  x281 &  x299 &  x302 &  x314 &  x317 &  x350 &  x388 &  x398 &  x404 &  x422 &  x434 &  x437 &  x452 &  x505 &  x560 &  x575 &  x605 &  x698 &  x701 &  x739 &  x749 &  x770 &  x791 &  x842 &  x854 &  x875 &  x953 &  x971 &  x1028 &  x1058 &  x1127 & ~x249;
assign c1279 =  x128 &  x514 &  x741 & ~x747 & ~x825 & ~x864;
assign c1281 =  x26 &  x242 &  x358 &  x398 &  x425 &  x446 &  x485 &  x574 &  x812 &  x863 &  x872 &  x953 &  x1022 &  x1034 &  x1043 &  x1109 & ~x636 & ~x676;
assign c1283 =  x325 &  x538 & ~x522 & ~x649;
assign c1285 =  x349 &  x568 &  x760 &  x931 &  x934;
assign c1287 =  x307 &  x415 &  x529 &  x532 &  x1006 & ~x1119;
assign c1289 =  x624 & ~x571;
assign c1291 =  x38 &  x47 &  x431 &  x485 &  x491 &  x644 &  x649 &  x662 &  x701 &  x704 &  x943 &  x989 &  x1033 & ~x183 & ~x480 & ~x516;
assign c1293 =  x2 &  x5 &  x23 &  x29 &  x38 &  x47 &  x89 &  x92 &  x125 &  x143 &  x170 &  x173 &  x179 &  x206 &  x221 &  x227 &  x254 &  x257 &  x276 &  x277 &  x356 &  x371 &  x401 &  x413 &  x422 &  x428 &  x434 &  x455 &  x461 &  x476 &  x485 &  x518 &  x530 &  x551 &  x560 &  x563 &  x572 &  x590 &  x614 &  x629 &  x644 &  x695 &  x701 &  x704 &  x779 &  x803 &  x812 &  x818 &  x839 &  x842 &  x905 &  x908 &  x920 &  x938 &  x944 &  x959 &  x1052 &  x1064 &  x1073 &  x1082 &  x1118 & ~x357 & ~x396 & ~x435 & ~x588;
assign c1295 =  x163 &  x319 &  x547 & ~x442 & ~x828;
assign c1297 =  x317 &  x443 &  x536 &  x554 &  x572 &  x641 &  x694 &  x842 &  x929 &  x1022 &  x1082 & ~x282 & ~x531 & ~x708 & ~x1080;
assign c1299 =  x17 &  x41 &  x44 &  x119 &  x131 &  x161 &  x164 &  x191 &  x203 &  x206 &  x218 &  x281 &  x287 &  x311 &  x398 &  x428 &  x632 &  x662 &  x674 &  x686 &  x719 &  x773 &  x782 &  x800 &  x803 &  x827 &  x860 &  x866 &  x884 &  x910 &  x926 &  x953 &  x955 &  x956 &  x992 &  x1034 &  x1037 &  x1052 &  x1058 &  x1091 &  x1097 &  x1099 &  x1100 &  x1109 &  x1130 & ~x402 & ~x672 & ~x702 & ~x897 & ~x936 & ~x1053;
assign c20 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x59 &  x62 &  x65 &  x71 &  x74 &  x83 &  x86 &  x89 &  x92 &  x98 &  x104 &  x107 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x134 &  x137 &  x140 &  x146 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x218 &  x221 &  x224 &  x230 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x320 &  x323 &  x326 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x464 &  x467 &  x473 &  x476 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x545 &  x548 &  x554 &  x557 &  x560 &  x563 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x704 &  x710 &  x716 &  x722 &  x725 &  x728 &  x731 &  x734 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x776 &  x779 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x824 &  x830 &  x833 &  x836 &  x839 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x869 &  x872 &  x875 &  x878 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x911 &  x920 &  x923 &  x932 &  x935 &  x938 &  x941 &  x947 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x976 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x234 & ~x651 & ~x786 & ~x825 & ~x864 & ~x870 & ~x882 & ~x1020 & ~x1098 & ~x1116;
assign c22 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x248 &  x251 &  x260 &  x263 &  x269 &  x272 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x352 &  x353 &  x356 &  x362 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x386 &  x389 &  x391 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x614 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x785 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x896 &  x899 &  x905 &  x908 &  x911 &  x914 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x977 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x378 & ~x438 & ~x477 & ~x492 & ~x510 & ~x513 & ~x531 & ~x552 & ~x570 & ~x627 & ~x648 & ~x666 & ~x705 & ~x744;
assign c24 =  x2 &  x5 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x62 &  x68 &  x71 &  x77 &  x83 &  x86 &  x89 &  x92 &  x95 &  x101 &  x104 &  x107 &  x110 &  x116 &  x119 &  x122 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x182 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x257 &  x260 &  x263 &  x266 &  x272 &  x275 &  x278 &  x283 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x353 &  x356 &  x361 &  x362 &  x365 &  x368 &  x374 &  x377 &  x380 &  x383 &  x389 &  x392 &  x395 &  x404 &  x416 &  x419 &  x422 &  x428 &  x431 &  x437 &  x443 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x488 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x518 &  x521 &  x524 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x584 &  x593 &  x596 &  x599 &  x605 &  x611 &  x614 &  x617 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x662 &  x665 &  x668 &  x671 &  x674 &  x683 &  x686 &  x689 &  x692 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x758 &  x764 &  x767 &  x770 &  x776 &  x779 &  x782 &  x785 &  x788 &  x797 &  x800 &  x803 &  x806 &  x809 &  x815 &  x818 &  x821 &  x827 &  x830 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x860 &  x863 &  x866 &  x869 &  x878 &  x881 &  x884 &  x887 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x947 &  x950 &  x953 &  x956 &  x959 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1052 &  x1055 &  x1058 &  x1061 &  x1067 &  x1073 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x33 & ~x222 & ~x495 & ~x726 & ~x747 & ~x861 & ~x900 & ~x939 & ~x978 & ~x1080 & ~x1119;
assign c26 =  x5 &  x23 &  x29 &  x38 &  x50 &  x59 &  x62 &  x116 &  x122 &  x146 &  x149 &  x161 &  x176 &  x179 &  x188 &  x194 &  x197 &  x206 &  x215 &  x221 &  x239 &  x257 &  x269 &  x275 &  x284 &  x296 &  x308 &  x317 &  x320 &  x326 &  x338 &  x344 &  x347 &  x350 &  x353 &  x362 &  x364 &  x371 &  x410 &  x428 &  x431 &  x442 &  x446 &  x455 &  x461 &  x476 &  x482 &  x485 &  x487 &  x497 &  x503 &  x506 &  x512 &  x515 &  x518 &  x520 &  x532 &  x554 &  x559 &  x569 &  x571 &  x590 &  x596 &  x599 &  x607 &  x608 &  x632 &  x641 &  x650 &  x686 &  x716 &  x719 &  x725 &  x749 &  x755 &  x761 &  x776 &  x779 &  x782 &  x784 &  x785 &  x788 &  x791 &  x809 &  x824 &  x830 &  x851 &  x857 &  x866 &  x881 &  x884 &  x887 &  x941 &  x947 &  x950 &  x953 &  x977 &  x991 &  x998 &  x1013 &  x1034 &  x1049 &  x1061 &  x1076 &  x1085 &  x1091 &  x1106 &  x1124 &  x1127 & ~x885 & ~x921;
assign c28 =  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x41 &  x44 &  x47 &  x50 &  x53 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x230 &  x233 &  x236 &  x242 &  x245 &  x248 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x358 &  x359 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x401 &  x407 &  x410 &  x413 &  x415 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x454 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x542 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x596 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x677 &  x680 &  x686 &  x689 &  x695 &  x698 &  x703 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x872 &  x875 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x934 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x998 &  x1001 &  x1004 &  x1007 &  x1009 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1048 &  x1049 &  x1052 &  x1055 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x942 & ~x978;
assign c210 =  x5 &  x11 &  x14 &  x17 &  x23 &  x35 &  x38 &  x44 &  x50 &  x53 &  x56 &  x62 &  x65 &  x68 &  x74 &  x77 &  x80 &  x86 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x119 &  x122 &  x134 &  x137 &  x140 &  x142 &  x143 &  x152 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x181 &  x182 &  x188 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x224 &  x227 &  x236 &  x239 &  x245 &  x248 &  x251 &  x254 &  x260 &  x263 &  x266 &  x272 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x305 &  x308 &  x317 &  x320 &  x329 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x368 &  x374 &  x377 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x400 &  x401 &  x404 &  x410 &  x413 &  x419 &  x422 &  x425 &  x428 &  x437 &  x439 &  x443 &  x446 &  x449 &  x452 &  x458 &  x461 &  x467 &  x470 &  x473 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x506 &  x521 &  x527 &  x530 &  x533 &  x542 &  x548 &  x554 &  x557 &  x560 &  x566 &  x572 &  x578 &  x590 &  x593 &  x596 &  x602 &  x605 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x659 &  x665 &  x671 &  x674 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x731 &  x734 &  x737 &  x746 &  x749 &  x752 &  x755 &  x764 &  x770 &  x773 &  x776 &  x782 &  x788 &  x791 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x830 &  x836 &  x839 &  x842 &  x845 &  x854 &  x857 &  x860 &  x866 &  x875 &  x878 &  x881 &  x884 &  x887 &  x893 &  x908 &  x911 &  x914 &  x917 &  x920 &  x926 &  x932 &  x938 &  x944 &  x953 &  x959 &  x962 &  x965 &  x968 &  x971 &  x977 &  x980 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1094 &  x1097 &  x1100 &  x1103 &  x1118 &  x1121 &  x1130 & ~x654 & ~x903 & ~x904 & ~x942 & ~x981 & ~x1020 & ~x1038;
assign c212 =  x2 &  x8 &  x11 &  x14 &  x17 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x71 &  x74 &  x77 &  x80 &  x83 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x113 &  x116 &  x119 &  x125 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x54 & ~x93 & ~x522 & ~x561 & ~x600 & ~x639 & ~x648 & ~x687 & ~x688 & ~x726 & ~x765 & ~x786 & ~x804 & ~x825 & ~x843 & ~x870;
assign c214 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x50 &  x53 &  x56 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x92 &  x101 &  x107 &  x110 &  x113 &  x116 &  x121 &  x122 &  x128 &  x131 &  x134 &  x143 &  x146 &  x149 &  x152 &  x158 &  x160 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x199 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x224 &  x227 &  x230 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x272 &  x275 &  x278 &  x284 &  x290 &  x293 &  x296 &  x299 &  x302 &  x311 &  x313 &  x314 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x344 &  x347 &  x350 &  x352 &  x353 &  x359 &  x365 &  x371 &  x380 &  x383 &  x389 &  x392 &  x395 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x423 &  x424 &  x428 &  x431 &  x437 &  x443 &  x449 &  x458 &  x461 &  x462 &  x463 &  x464 &  x473 &  x476 &  x491 &  x494 &  x497 &  x500 &  x501 &  x502 &  x503 &  x506 &  x512 &  x515 &  x518 &  x521 &  x527 &  x530 &  x539 &  x542 &  x545 &  x551 &  x557 &  x560 &  x566 &  x572 &  x575 &  x580 &  x581 &  x584 &  x587 &  x593 &  x599 &  x601 &  x605 &  x611 &  x614 &  x617 &  x620 &  x626 &  x632 &  x635 &  x638 &  x640 &  x641 &  x644 &  x647 &  x650 &  x656 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x679 &  x680 &  x683 &  x686 &  x692 &  x701 &  x704 &  x707 &  x713 &  x716 &  x718 &  x719 &  x722 &  x725 &  x728 &  x731 &  x737 &  x743 &  x749 &  x752 &  x758 &  x761 &  x764 &  x773 &  x776 &  x779 &  x782 &  x785 &  x800 &  x806 &  x812 &  x815 &  x818 &  x821 &  x827 &  x830 &  x836 &  x842 &  x845 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x872 &  x875 &  x878 &  x881 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x926 &  x929 &  x932 &  x941 &  x944 &  x950 &  x959 &  x965 &  x968 &  x971 &  x974 &  x977 &  x986 &  x989 &  x998 &  x1001 &  x1004 &  x1010 &  x1019 &  x1028 &  x1031 &  x1037 &  x1043 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x396 & ~x435 & ~x513;
assign c216 =  x2 &  x5 &  x8 &  x11 &  x17 &  x23 &  x26 &  x32 &  x35 &  x38 &  x41 &  x44 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x74 &  x92 &  x101 &  x104 &  x107 &  x110 &  x119 &  x122 &  x125 &  x137 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x176 &  x179 &  x185 &  x191 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x214 &  x215 &  x218 &  x220 &  x221 &  x227 &  x233 &  x236 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x269 &  x272 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x362 &  x377 &  x383 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x437 &  x439 &  x440 &  x443 &  x446 &  x449 &  x455 &  x458 &  x467 &  x470 &  x472 &  x473 &  x476 &  x479 &  x482 &  x485 &  x491 &  x497 &  x500 &  x503 &  x509 &  x512 &  x515 &  x521 &  x524 &  x530 &  x533 &  x542 &  x547 &  x551 &  x554 &  x560 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x596 &  x599 &  x605 &  x608 &  x611 &  x614 &  x617 &  x623 &  x625 &  x626 &  x629 &  x632 &  x635 &  x641 &  x644 &  x647 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x683 &  x686 &  x698 &  x701 &  x704 &  x707 &  x713 &  x716 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x770 &  x773 &  x776 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x815 &  x818 &  x821 &  x824 &  x836 &  x839 &  x842 &  x848 &  x857 &  x860 &  x866 &  x869 &  x872 &  x875 &  x878 &  x887 &  x890 &  x893 &  x899 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x953 &  x956 &  x962 &  x965 &  x968 &  x977 &  x983 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1031 &  x1037 &  x1040 &  x1043 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x591 & ~x630 & ~x669 & ~x708 & ~x786 & ~x822 & ~x861 & ~x900;
assign c218 =  x2 &  x5 &  x11 &  x14 &  x17 &  x20 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x80 &  x83 &  x86 &  x89 &  x98 &  x101 &  x104 &  x113 &  x121 &  x122 &  x125 &  x128 &  x131 &  x134 &  x143 &  x146 &  x149 &  x155 &  x160 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x185 &  x188 &  x189 &  x191 &  x197 &  x199 &  x200 &  x206 &  x209 &  x212 &  x227 &  x229 &  x230 &  x233 &  x236 &  x238 &  x239 &  x242 &  x248 &  x251 &  x260 &  x266 &  x269 &  x272 &  x278 &  x284 &  x287 &  x290 &  x299 &  x302 &  x305 &  x311 &  x314 &  x317 &  x320 &  x323 &  x329 &  x332 &  x335 &  x338 &  x347 &  x353 &  x356 &  x371 &  x377 &  x383 &  x389 &  x392 &  x398 &  x401 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x437 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x473 &  x479 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x524 &  x527 &  x530 &  x536 &  x542 &  x545 &  x548 &  x551 &  x554 &  x560 &  x566 &  x569 &  x575 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x640 &  x641 &  x647 &  x650 &  x653 &  x656 &  x659 &  x665 &  x668 &  x671 &  x677 &  x679 &  x683 &  x701 &  x718 &  x719 &  x722 &  x728 &  x731 &  x734 &  x737 &  x740 &  x749 &  x755 &  x757 &  x758 &  x761 &  x764 &  x770 &  x773 &  x779 &  x782 &  x785 &  x791 &  x794 &  x797 &  x800 &  x803 &  x809 &  x815 &  x818 &  x824 &  x827 &  x839 &  x842 &  x845 &  x848 &  x851 &  x860 &  x863 &  x866 &  x869 &  x872 &  x878 &  x881 &  x884 &  x890 &  x893 &  x899 &  x902 &  x905 &  x911 &  x920 &  x926 &  x929 &  x935 &  x938 &  x941 &  x944 &  x950 &  x953 &  x956 &  x959 &  x962 &  x968 &  x971 &  x974 &  x980 &  x983 &  x986 &  x989 &  x995 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1034 &  x1037 &  x1039 &  x1043 &  x1049 &  x1055 &  x1058 &  x1064 &  x1067 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130 & ~x627 & ~x666 & ~x705 & ~x744 & ~x783 & ~x936;
assign c220 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x205 &  x206 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x242 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x283 &  x287 &  x293 &  x295 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x316 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x419 &  x425 &  x428 &  x430 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x464 &  x467 &  x469 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x560 &  x563 &  x566 &  x569 &  x575 &  x578 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x601 &  x602 &  x611 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x794 &  x797 &  x800 &  x806 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x381 & ~x420 & ~x421 & ~x459 & ~x498 & ~x705 & ~x744 & ~x783;
assign c222 =  x5 &  x8 &  x11 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x47 &  x50 &  x53 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x89 &  x92 &  x98 &  x101 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x296 &  x298 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x358 &  x362 &  x364 &  x368 &  x374 &  x377 &  x383 &  x386 &  x389 &  x392 &  x395 &  x397 &  x398 &  x401 &  x404 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x436 &  x437 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x512 &  x518 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x542 &  x548 &  x551 &  x554 &  x557 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x587 &  x590 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x626 &  x629 &  x635 &  x638 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x701 &  x710 &  x713 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x746 &  x749 &  x752 &  x761 &  x764 &  x767 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x818 &  x821 &  x824 &  x827 &  x833 &  x836 &  x839 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x875 &  x878 &  x881 &  x884 &  x887 &  x892 &  x893 &  x896 &  x899 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x944 &  x947 &  x959 &  x962 &  x965 &  x971 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1130 & ~x675 & ~x726 & ~x825 & ~x864 & ~x882 & ~x903 & ~x921 & ~x1038 & ~x1077 & ~x1116;
assign c224 =  x2 &  x5 &  x8 &  x11 &  x14 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x104 &  x107 &  x113 &  x119 &  x122 &  x125 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x152 &  x155 &  x158 &  x161 &  x164 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x197 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x240 &  x241 &  x242 &  x248 &  x251 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x314 &  x315 &  x317 &  x320 &  x322 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x355 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x391 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x433 &  x434 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x467 &  x469 &  x470 &  x473 &  x476 &  x479 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x641 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x689 &  x692 &  x701 &  x704 &  x707 &  x710 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x785 &  x788 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x851 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x947 &  x950 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x783;
assign c226 =  x2 &  x8 &  x14 &  x17 &  x26 &  x29 &  x32 &  x38 &  x50 &  x56 &  x59 &  x65 &  x74 &  x89 &  x92 &  x101 &  x122 &  x128 &  x134 &  x137 &  x140 &  x146 &  x149 &  x164 &  x170 &  x173 &  x182 &  x206 &  x209 &  x224 &  x227 &  x230 &  x233 &  x242 &  x254 &  x257 &  x269 &  x290 &  x293 &  x299 &  x305 &  x311 &  x317 &  x326 &  x329 &  x335 &  x338 &  x341 &  x347 &  x350 &  x362 &  x368 &  x374 &  x389 &  x392 &  x398 &  x404 &  x416 &  x421 &  x425 &  x431 &  x443 &  x449 &  x452 &  x455 &  x459 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x503 &  x509 &  x512 &  x530 &  x533 &  x539 &  x545 &  x548 &  x551 &  x557 &  x560 &  x563 &  x572 &  x584 &  x587 &  x596 &  x599 &  x605 &  x611 &  x614 &  x626 &  x638 &  x641 &  x644 &  x647 &  x650 &  x656 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x692 &  x695 &  x701 &  x710 &  x713 &  x716 &  x722 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x752 &  x755 &  x758 &  x764 &  x770 &  x773 &  x776 &  x782 &  x797 &  x800 &  x806 &  x809 &  x812 &  x818 &  x833 &  x836 &  x842 &  x848 &  x851 &  x857 &  x863 &  x878 &  x887 &  x890 &  x893 &  x905 &  x908 &  x914 &  x920 &  x923 &  x932 &  x938 &  x944 &  x947 &  x950 &  x953 &  x959 &  x962 &  x965 &  x968 &  x971 &  x973 &  x977 &  x980 &  x986 &  x989 &  x992 &  x1001 &  x1013 &  x1019 &  x1028 &  x1034 &  x1052 &  x1058 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1097 &  x1100 &  x1109 &  x1115 &  x1124 &  x1127 & ~x165 & ~x321 & ~x663;
assign c228 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x41 &  x47 &  x59 &  x62 &  x65 &  x68 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x101 &  x110 &  x113 &  x119 &  x122 &  x125 &  x131 &  x137 &  x140 &  x143 &  x146 &  x152 &  x155 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x215 &  x224 &  x227 &  x230 &  x233 &  x236 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x266 &  x269 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x299 &  x302 &  x305 &  x308 &  x311 &  x317 &  x319 &  x320 &  x326 &  x329 &  x335 &  x338 &  x341 &  x344 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x380 &  x383 &  x389 &  x395 &  x397 &  x398 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x452 &  x458 &  x461 &  x467 &  x470 &  x476 &  x485 &  x487 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x512 &  x515 &  x521 &  x527 &  x530 &  x533 &  x536 &  x542 &  x545 &  x551 &  x566 &  x569 &  x572 &  x575 &  x581 &  x590 &  x592 &  x593 &  x596 &  x602 &  x611 &  x623 &  x626 &  x632 &  x635 &  x641 &  x647 &  x650 &  x653 &  x665 &  x671 &  x677 &  x680 &  x683 &  x686 &  x689 &  x695 &  x698 &  x701 &  x707 &  x713 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x745 &  x746 &  x749 &  x755 &  x758 &  x764 &  x770 &  x785 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x830 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x872 &  x875 &  x881 &  x884 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x920 &  x923 &  x926 &  x938 &  x941 &  x944 &  x947 &  x953 &  x962 &  x968 &  x971 &  x974 &  x977 &  x980 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1064 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1112 &  x1121 &  x1130 & ~x276 & ~x312 & ~x315 & ~x351 & ~x390 & ~x429 & ~x942 & ~x1056;
assign c230 =  x5 &  x14 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x44 &  x47 &  x50 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x86 &  x92 &  x95 &  x101 &  x104 &  x110 &  x113 &  x125 &  x128 &  x131 &  x134 &  x143 &  x146 &  x149 &  x155 &  x163 &  x164 &  x167 &  x170 &  x173 &  x179 &  x182 &  x188 &  x191 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x227 &  x239 &  x242 &  x245 &  x251 &  x254 &  x257 &  x260 &  x263 &  x272 &  x277 &  x281 &  x284 &  x287 &  x290 &  x296 &  x302 &  x305 &  x308 &  x313 &  x314 &  x316 &  x317 &  x320 &  x323 &  x326 &  x335 &  x344 &  x347 &  x352 &  x353 &  x355 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x391 &  x394 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x430 &  x431 &  x437 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x469 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x491 &  x494 &  x497 &  x506 &  x508 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x566 &  x569 &  x578 &  x581 &  x584 &  x587 &  x590 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x620 &  x623 &  x626 &  x632 &  x635 &  x638 &  x641 &  x647 &  x650 &  x659 &  x662 &  x665 &  x668 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x770 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x812 &  x815 &  x818 &  x821 &  x827 &  x830 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x866 &  x872 &  x881 &  x884 &  x890 &  x893 &  x905 &  x911 &  x914 &  x920 &  x923 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x950 &  x959 &  x965 &  x971 &  x977 &  x989 &  x992 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1049 &  x1052 &  x1058 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130 & ~x474 & ~x513 & ~x552 & ~x555 & ~x588 & ~x594 & ~x666 & ~x744 & ~x783;
assign c232 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x80 &  x83 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x166 &  x167 &  x170 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x218 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x244 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x272 &  x275 &  x281 &  x284 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x314 &  x316 &  x320 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x391 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x424 &  x425 &  x428 &  x434 &  x437 &  x440 &  x443 &  x446 &  x452 &  x461 &  x464 &  x466 &  x467 &  x470 &  x473 &  x476 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x502 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x688 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x713 &  x716 &  x719 &  x722 &  x725 &  x727 &  x728 &  x731 &  x734 &  x740 &  x743 &  x746 &  x749 &  x752 &  x758 &  x761 &  x764 &  x767 &  x770 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x893 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x932 &  x935 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x375 & ~x414;
assign c234 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x113 &  x116 &  x119 &  x122 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x197 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x377 &  x380 &  x383 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x455 &  x461 &  x464 &  x467 &  x470 &  x476 &  x479 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x814 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x863 &  x866 &  x869 &  x872 &  x878 &  x881 &  x884 &  x887 &  x890 &  x892 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x931 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x970 &  x971 &  x974 &  x980 &  x983 &  x986 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1009 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1048 &  x1049 &  x1055 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x243 & ~x282 & ~x321 & ~x390 & ~x468 & ~x507 & ~x508 & ~x546 & ~x585 & ~x729 & ~x768;
assign c236 =  x11 &  x17 &  x32 &  x44 &  x50 &  x56 &  x62 &  x74 &  x77 &  x95 &  x101 &  x104 &  x110 &  x113 &  x116 &  x131 &  x149 &  x164 &  x200 &  x203 &  x209 &  x212 &  x218 &  x224 &  x227 &  x233 &  x242 &  x245 &  x254 &  x257 &  x272 &  x281 &  x299 &  x302 &  x317 &  x323 &  x359 &  x371 &  x395 &  x401 &  x434 &  x437 &  x440 &  x446 &  x449 &  x455 &  x458 &  x461 &  x462 &  x464 &  x467 &  x470 &  x473 &  x479 &  x482 &  x488 &  x494 &  x512 &  x524 &  x533 &  x554 &  x563 &  x569 &  x590 &  x593 &  x599 &  x617 &  x618 &  x619 &  x629 &  x638 &  x641 &  x644 &  x647 &  x653 &  x659 &  x662 &  x671 &  x677 &  x698 &  x704 &  x716 &  x718 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x736 &  x761 &  x773 &  x796 &  x803 &  x809 &  x815 &  x824 &  x835 &  x854 &  x857 &  x863 &  x869 &  x874 &  x875 &  x884 &  x890 &  x902 &  x920 &  x923 &  x935 &  x950 &  x953 &  x956 &  x971 &  x974 &  x980 &  x998 &  x1010 &  x1019 &  x1022 &  x1028 &  x1043 &  x1052 &  x1061 &  x1070 &  x1079 &  x1088 &  x1094 &  x1097 &  x1103 &  x1121 & ~x372;
assign c238 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x29 &  x32 &  x35 &  x41 &  x50 &  x53 &  x56 &  x62 &  x65 &  x71 &  x74 &  x77 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x107 &  x110 &  x119 &  x125 &  x128 &  x131 &  x134 &  x137 &  x143 &  x146 &  x149 &  x155 &  x161 &  x164 &  x167 &  x170 &  x176 &  x179 &  x182 &  x188 &  x194 &  x197 &  x212 &  x215 &  x221 &  x227 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x272 &  x275 &  x278 &  x281 &  x284 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x314 &  x317 &  x323 &  x326 &  x329 &  x338 &  x341 &  x344 &  x347 &  x350 &  x356 &  x358 &  x365 &  x374 &  x380 &  x383 &  x386 &  x389 &  x395 &  x398 &  x401 &  x419 &  x425 &  x428 &  x446 &  x449 &  x455 &  x472 &  x473 &  x476 &  x479 &  x485 &  x488 &  x491 &  x503 &  x506 &  x511 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x542 &  x545 &  x554 &  x557 &  x566 &  x572 &  x575 &  x581 &  x584 &  x587 &  x593 &  x599 &  x608 &  x614 &  x626 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x658 &  x659 &  x662 &  x665 &  x674 &  x680 &  x686 &  x689 &  x697 &  x701 &  x704 &  x710 &  x716 &  x725 &  x734 &  x743 &  x749 &  x752 &  x755 &  x758 &  x761 &  x767 &  x770 &  x775 &  x776 &  x779 &  x788 &  x794 &  x800 &  x809 &  x812 &  x813 &  x814 &  x815 &  x818 &  x821 &  x827 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x853 &  x854 &  x857 &  x860 &  x884 &  x887 &  x892 &  x893 &  x896 &  x899 &  x908 &  x911 &  x914 &  x917 &  x923 &  x932 &  x935 &  x938 &  x941 &  x947 &  x953 &  x959 &  x962 &  x965 &  x974 &  x977 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1037 &  x1040 &  x1043 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1082 &  x1085 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x519 & ~x792;
assign c240 =  x5 &  x6 &  x7 &  x14 &  x29 &  x35 &  x38 &  x41 &  x53 &  x56 &  x62 &  x65 &  x68 &  x77 &  x80 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x116 &  x119 &  x122 &  x128 &  x131 &  x134 &  x140 &  x143 &  x146 &  x158 &  x164 &  x170 &  x173 &  x176 &  x191 &  x194 &  x197 &  x212 &  x215 &  x224 &  x230 &  x233 &  x236 &  x239 &  x251 &  x254 &  x257 &  x269 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x316 &  x317 &  x326 &  x329 &  x332 &  x335 &  x341 &  x347 &  x350 &  x353 &  x356 &  x359 &  x365 &  x371 &  x377 &  x383 &  x389 &  x395 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x443 &  x455 &  x467 &  x470 &  x479 &  x482 &  x485 &  x491 &  x494 &  x497 &  x503 &  x506 &  x512 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x545 &  x551 &  x554 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x593 &  x602 &  x605 &  x608 &  x614 &  x620 &  x623 &  x635 &  x638 &  x641 &  x644 &  x647 &  x653 &  x659 &  x662 &  x665 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x701 &  x704 &  x707 &  x710 &  x716 &  x719 &  x728 &  x731 &  x734 &  x737 &  x743 &  x752 &  x757 &  x758 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x809 &  x821 &  x824 &  x827 &  x833 &  x835 &  x842 &  x848 &  x857 &  x860 &  x863 &  x866 &  x869 &  x881 &  x884 &  x892 &  x893 &  x899 &  x908 &  x914 &  x917 &  x920 &  x923 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x953 &  x956 &  x965 &  x968 &  x974 &  x977 &  x980 &  x986 &  x989 &  x995 &  x1001 &  x1004 &  x1007 &  x1019 &  x1022 &  x1025 &  x1028 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1067 &  x1070 &  x1082 &  x1088 &  x1097 &  x1100 &  x1118 &  x1121 &  x1130 & ~x783 & ~x861 & ~x957;
assign c242 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x29 &  x32 &  x38 &  x41 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x107 &  x110 &  x113 &  x119 &  x125 &  x128 &  x131 &  x137 &  x140 &  x146 &  x149 &  x152 &  x155 &  x161 &  x164 &  x167 &  x170 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x251 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x305 &  x308 &  x311 &  x314 &  x320 &  x323 &  x326 &  x332 &  x335 &  x341 &  x344 &  x347 &  x350 &  x353 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x380 &  x383 &  x389 &  x392 &  x395 &  x398 &  x401 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x464 &  x467 &  x470 &  x479 &  x482 &  x485 &  x488 &  x491 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x662 &  x668 &  x671 &  x674 &  x677 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x725 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x797 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x833 &  x836 &  x839 &  x842 &  x845 &  x851 &  x854 &  x857 &  x860 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x920 &  x926 &  x929 &  x935 &  x938 &  x941 &  x944 &  x947 &  x953 &  x959 &  x962 &  x965 &  x968 &  x971 &  x977 &  x980 &  x983 &  x986 &  x989 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 & ~x72 & ~x90 & ~x144 & ~x183 & ~x363 & ~x519 & ~x558 & ~x570 & ~x636 & ~x648 & ~x900 & ~x939 & ~x978 & ~x1017 & ~x1056;
assign c244 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x163 &  x164 &  x167 &  x169 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x202 &  x203 &  x206 &  x208 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x241 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x280 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x319 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x397 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x631 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x892 &  x893 &  x896 &  x898 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x923 &  x926 &  x929 &  x931 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x970 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x991 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1009 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x687;
assign c246 =  x2 &  x5 &  x14 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x143 &  x155 &  x158 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x272 &  x275 &  x281 &  x284 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x389 &  x392 &  x395 &  x398 &  x404 &  x410 &  x413 &  x416 &  x419 &  x422 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x449 &  x452 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x485 &  x488 &  x491 &  x494 &  x497 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x548 &  x551 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x611 &  x617 &  x623 &  x632 &  x635 &  x644 &  x647 &  x656 &  x659 &  x665 &  x668 &  x671 &  x674 &  x677 &  x683 &  x686 &  x692 &  x698 &  x701 &  x704 &  x710 &  x716 &  x719 &  x725 &  x728 &  x731 &  x734 &  x737 &  x743 &  x752 &  x761 &  x767 &  x770 &  x773 &  x779 &  x782 &  x791 &  x794 &  x800 &  x803 &  x806 &  x809 &  x812 &  x818 &  x821 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x893 &  x902 &  x905 &  x908 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x980 &  x983 &  x986 &  x989 &  x995 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1130 & ~x195 & ~x339 & ~x492 & ~x495 & ~x531 & ~x534 & ~x570 & ~x609 & ~x648 & ~x669 & ~x687 & ~x708 & ~x726 & ~x765 & ~x864 & ~x882 & ~x981;
assign c248 =  x2 &  x5 &  x8 &  x11 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x319 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x358 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x395 &  x397 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x449 &  x452 &  x455 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x488 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x550 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x587 &  x589 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x611 &  x614 &  x617 &  x620 &  x623 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x710 &  x713 &  x716 &  x722 &  x725 &  x728 &  x731 &  x734 &  x736 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x775 &  x776 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x814 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x852 &  x853 &  x854 &  x860 &  x866 &  x869 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x892 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x926 &  x929 &  x931 &  x932 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1063 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x273 & ~x312 & ~x351;
assign c250 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x44 &  x50 &  x59 &  x62 &  x65 &  x74 &  x86 &  x89 &  x92 &  x101 &  x104 &  x119 &  x125 &  x137 &  x143 &  x146 &  x149 &  x152 &  x158 &  x170 &  x185 &  x194 &  x197 &  x203 &  x209 &  x212 &  x230 &  x242 &  x245 &  x251 &  x257 &  x260 &  x272 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x317 &  x323 &  x329 &  x338 &  x341 &  x344 &  x347 &  x353 &  x359 &  x362 &  x368 &  x371 &  x380 &  x383 &  x389 &  x392 &  x395 &  x413 &  x422 &  x428 &  x431 &  x443 &  x446 &  x449 &  x458 &  x464 &  x470 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x497 &  x506 &  x521 &  x524 &  x527 &  x533 &  x539 &  x542 &  x548 &  x551 &  x557 &  x563 &  x575 &  x578 &  x590 &  x602 &  x608 &  x611 &  x617 &  x623 &  x629 &  x635 &  x647 &  x650 &  x653 &  x656 &  x659 &  x668 &  x671 &  x680 &  x686 &  x689 &  x692 &  x698 &  x701 &  x704 &  x707 &  x722 &  x725 &  x728 &  x731 &  x743 &  x746 &  x749 &  x758 &  x767 &  x770 &  x773 &  x779 &  x782 &  x788 &  x800 &  x812 &  x815 &  x827 &  x830 &  x836 &  x848 &  x857 &  x863 &  x869 &  x875 &  x881 &  x887 &  x890 &  x896 &  x899 &  x902 &  x911 &  x920 &  x926 &  x932 &  x938 &  x941 &  x944 &  x947 &  x953 &  x959 &  x962 &  x965 &  x968 &  x974 &  x977 &  x980 &  x983 &  x986 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1019 &  x1022 &  x1031 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1070 &  x1082 &  x1109 &  x1118 &  x1121 &  x1124 & ~x15 & ~x99 & ~x495 & ~x726 & ~x747 & ~x768 & ~x807 & ~x846 & ~x885 & ~x900 & ~x939 & ~x978 & ~x1017 & ~x1056 & ~x1080;
assign c252 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x19 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x694 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x733 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x27 & ~x66 & ~x183 & ~x300 & ~x339 & ~x378 & ~x417 & ~x495 & ~x708 & ~x864;
assign c254 =  x17 &  x20 &  x29 &  x32 &  x44 &  x47 &  x56 &  x62 &  x71 &  x74 &  x77 &  x89 &  x98 &  x101 &  x128 &  x140 &  x143 &  x146 &  x149 &  x170 &  x173 &  x185 &  x188 &  x194 &  x197 &  x209 &  x218 &  x245 &  x257 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x287 &  x296 &  x302 &  x305 &  x308 &  x311 &  x316 &  x323 &  x326 &  x329 &  x353 &  x356 &  x359 &  x362 &  x368 &  x371 &  x380 &  x383 &  x385 &  x395 &  x410 &  x425 &  x428 &  x431 &  x458 &  x461 &  x470 &  x473 &  x476 &  x485 &  x487 &  x491 &  x494 &  x497 &  x503 &  x515 &  x521 &  x526 &  x542 &  x557 &  x563 &  x572 &  x590 &  x596 &  x602 &  x611 &  x620 &  x626 &  x640 &  x641 &  x656 &  x659 &  x665 &  x668 &  x674 &  x689 &  x692 &  x698 &  x707 &  x713 &  x722 &  x725 &  x737 &  x746 &  x749 &  x757 &  x758 &  x767 &  x773 &  x779 &  x782 &  x785 &  x796 &  x812 &  x818 &  x839 &  x848 &  x866 &  x872 &  x875 &  x887 &  x904 &  x905 &  x929 &  x932 &  x938 &  x950 &  x953 &  x956 &  x962 &  x965 &  x974 &  x986 &  x989 &  x994 &  x998 &  x1004 &  x1016 &  x1022 &  x1040 &  x1049 &  x1061 &  x1067 &  x1070 &  x1079 &  x1091 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 & ~x339 & ~x936;
assign c256 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x251 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x788 &  x791 &  x794 &  x797 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x950 &  x953 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x156 & ~x195 & ~x300 & ~x339 & ~x378 & ~x417 & ~x418 & ~x669 & ~x708 & ~x726 & ~x900 & ~x1056 & ~x1095;
assign c258 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x316 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x355 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x394 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x433 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x472 &  x473 &  x476 &  x479 &  x482 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x671 &  x674 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x890 &  x896 &  x899 &  x902 &  x905 &  x908 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x78 & ~x117 & ~x156 & ~x195 & ~x300 & ~x339 & ~x594 & ~x627 & ~x633 & ~x843;
assign c260 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x80 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x128 &  x131 &  x134 &  x137 &  x140 &  x146 &  x149 &  x152 &  x158 &  x161 &  x164 &  x167 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x245 &  x248 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x341 &  x353 &  x356 &  x359 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x398 &  x401 &  x404 &  x407 &  x410 &  x416 &  x422 &  x425 &  x428 &  x433 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x455 &  x461 &  x464 &  x470 &  x472 &  x473 &  x476 &  x479 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x548 &  x551 &  x554 &  x560 &  x563 &  x569 &  x572 &  x575 &  x581 &  x584 &  x599 &  x602 &  x605 &  x608 &  x611 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x656 &  x659 &  x662 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x722 &  x725 &  x728 &  x731 &  x737 &  x740 &  x743 &  x746 &  x752 &  x755 &  x758 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x809 &  x812 &  x815 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x845 &  x854 &  x857 &  x860 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x893 &  x896 &  x899 &  x902 &  x905 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1130 & ~x0 & ~x39 & ~x78 & ~x570 & ~x591 & ~x630 & ~x636 & ~x750 & ~x765 & ~x804 & ~x861 & ~x900 & ~x939;
assign c262 =  x2 &  x5 &  x29 &  x35 &  x38 &  x41 &  x56 &  x62 &  x65 &  x71 &  x83 &  x101 &  x110 &  x116 &  x122 &  x125 &  x131 &  x134 &  x137 &  x140 &  x149 &  x161 &  x167 &  x176 &  x179 &  x188 &  x197 &  x206 &  x212 &  x224 &  x227 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x266 &  x272 &  x275 &  x287 &  x293 &  x299 &  x305 &  x317 &  x320 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x356 &  x359 &  x368 &  x371 &  x374 &  x377 &  x380 &  x389 &  x392 &  x398 &  x401 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x437 &  x440 &  x449 &  x458 &  x461 &  x470 &  x473 &  x478 &  x479 &  x482 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x545 &  x554 &  x557 &  x560 &  x563 &  x575 &  x578 &  x581 &  x587 &  x599 &  x605 &  x608 &  x611 &  x617 &  x620 &  x623 &  x626 &  x629 &  x647 &  x671 &  x674 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x707 &  x710 &  x719 &  x734 &  x740 &  x746 &  x749 &  x758 &  x767 &  x770 &  x791 &  x794 &  x797 &  x800 &  x806 &  x818 &  x821 &  x830 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x860 &  x866 &  x869 &  x875 &  x896 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x929 &  x938 &  x944 &  x947 &  x953 &  x956 &  x962 &  x965 &  x971 &  x980 &  x995 &  x1004 &  x1007 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1040 &  x1043 &  x1049 &  x1058 &  x1061 &  x1063 &  x1073 &  x1079 &  x1085 &  x1088 &  x1100 &  x1103 &  x1109 &  x1115 &  x1118 &  x1130 & ~x717 & ~x747 & ~x756 & ~x786 & ~x825 & ~x864 & ~x978 & ~x981 & ~x1059;
assign c264 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x137 &  x140 &  x143 &  x152 &  x155 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x227 &  x233 &  x236 &  x239 &  x242 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x281 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x331 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x359 &  x364 &  x365 &  x368 &  x371 &  x374 &  x377 &  x383 &  x386 &  x395 &  x398 &  x401 &  x403 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x464 &  x470 &  x473 &  x475 &  x476 &  x479 &  x482 &  x485 &  x491 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x542 &  x545 &  x548 &  x557 &  x560 &  x566 &  x569 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x629 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x758 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x820 &  x821 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x892 &  x893 &  x898 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x931 &  x932 &  x935 &  x937 &  x938 &  x941 &  x947 &  x953 &  x956 &  x959 &  x965 &  x968 &  x970 &  x971 &  x974 &  x976 &  x980 &  x983 &  x986 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1009 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1069 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1093 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1118 &  x1121 &  x1130 & ~x156 & ~x195 & ~x234 & ~x273 & ~x351 & ~x390 & ~x882 & ~x903 & ~x942;
assign c266 =  x2 &  x5 &  x8 &  x11 &  x17 &  x26 &  x29 &  x32 &  x35 &  x41 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x77 &  x80 &  x83 &  x89 &  x92 &  x95 &  x98 &  x107 &  x113 &  x116 &  x122 &  x128 &  x134 &  x137 &  x146 &  x149 &  x155 &  x158 &  x161 &  x170 &  x173 &  x182 &  x185 &  x203 &  x206 &  x209 &  x212 &  x218 &  x221 &  x227 &  x236 &  x242 &  x245 &  x251 &  x260 &  x266 &  x269 &  x275 &  x278 &  x281 &  x284 &  x286 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x317 &  x319 &  x320 &  x326 &  x332 &  x350 &  x353 &  x356 &  x358 &  x362 &  x365 &  x374 &  x377 &  x383 &  x392 &  x407 &  x410 &  x413 &  x419 &  x422 &  x425 &  x431 &  x437 &  x440 &  x443 &  x446 &  x449 &  x455 &  x458 &  x461 &  x467 &  x470 &  x473 &  x479 &  x485 &  x491 &  x503 &  x518 &  x521 &  x526 &  x527 &  x530 &  x542 &  x545 &  x548 &  x551 &  x557 &  x560 &  x565 &  x566 &  x572 &  x575 &  x581 &  x587 &  x590 &  x593 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x629 &  x632 &  x635 &  x641 &  x647 &  x656 &  x662 &  x665 &  x671 &  x674 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x701 &  x710 &  x713 &  x716 &  x719 &  x722 &  x728 &  x731 &  x734 &  x737 &  x740 &  x746 &  x755 &  x764 &  x767 &  x779 &  x785 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x821 &  x830 &  x833 &  x839 &  x845 &  x848 &  x860 &  x863 &  x866 &  x875 &  x881 &  x884 &  x902 &  x905 &  x911 &  x914 &  x926 &  x929 &  x938 &  x944 &  x947 &  x953 &  x956 &  x962 &  x965 &  x968 &  x971 &  x986 &  x992 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1025 &  x1028 &  x1034 &  x1040 &  x1046 &  x1049 &  x1061 &  x1064 &  x1070 &  x1073 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1121 &  x1130 & ~x612 & ~x726 & ~x882 & ~x945 & ~x1038;
assign c268 =  x2 &  x8 &  x11 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x43 &  x44 &  x53 &  x56 &  x59 &  x62 &  x68 &  x74 &  x80 &  x81 &  x83 &  x89 &  x92 &  x104 &  x107 &  x110 &  x113 &  x120 &  x121 &  x122 &  x125 &  x131 &  x137 &  x146 &  x152 &  x158 &  x159 &  x161 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x206 &  x212 &  x218 &  x221 &  x224 &  x230 &  x233 &  x239 &  x245 &  x248 &  x263 &  x266 &  x269 &  x275 &  x287 &  x293 &  x296 &  x302 &  x305 &  x308 &  x314 &  x323 &  x329 &  x335 &  x338 &  x347 &  x362 &  x365 &  x380 &  x383 &  x386 &  x389 &  x392 &  x398 &  x404 &  x407 &  x416 &  x419 &  x422 &  x424 &  x425 &  x428 &  x431 &  x434 &  x440 &  x452 &  x461 &  x470 &  x473 &  x488 &  x491 &  x494 &  x497 &  x509 &  x518 &  x521 &  x523 &  x524 &  x539 &  x542 &  x545 &  x548 &  x560 &  x569 &  x575 &  x578 &  x584 &  x587 &  x596 &  x602 &  x605 &  x611 &  x623 &  x626 &  x635 &  x638 &  x644 &  x647 &  x656 &  x668 &  x674 &  x677 &  x686 &  x695 &  x701 &  x707 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x740 &  x746 &  x749 &  x752 &  x755 &  x761 &  x764 &  x767 &  x770 &  x773 &  x779 &  x788 &  x791 &  x794 &  x797 &  x806 &  x818 &  x821 &  x824 &  x830 &  x842 &  x848 &  x851 &  x854 &  x860 &  x863 &  x869 &  x872 &  x875 &  x881 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x935 &  x938 &  x941 &  x944 &  x950 &  x956 &  x962 &  x968 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1031 &  x1034 &  x1040 &  x1046 &  x1049 &  x1052 &  x1061 &  x1070 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1106 &  x1118 &  x1124 &  x1127 &  x1130 & ~x297 & ~x396 & ~x936 & ~x975 & ~x1014;
assign c270 =  x2 &  x14 &  x17 &  x20 &  x26 &  x29 &  x50 &  x53 &  x56 &  x59 &  x65 &  x74 &  x107 &  x116 &  x119 &  x121 &  x122 &  x131 &  x137 &  x140 &  x146 &  x149 &  x152 &  x158 &  x160 &  x164 &  x167 &  x170 &  x179 &  x182 &  x185 &  x188 &  x191 &  x197 &  x203 &  x212 &  x221 &  x224 &  x227 &  x230 &  x233 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x269 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x305 &  x308 &  x311 &  x314 &  x326 &  x329 &  x332 &  x335 &  x347 &  x352 &  x356 &  x359 &  x362 &  x368 &  x371 &  x374 &  x386 &  x389 &  x392 &  x395 &  x404 &  x407 &  x413 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x443 &  x446 &  x452 &  x461 &  x473 &  x479 &  x485 &  x494 &  x500 &  x503 &  x506 &  x518 &  x521 &  x524 &  x536 &  x545 &  x548 &  x560 &  x566 &  x569 &  x572 &  x575 &  x584 &  x608 &  x611 &  x620 &  x626 &  x629 &  x632 &  x647 &  x668 &  x674 &  x680 &  x692 &  x695 &  x698 &  x704 &  x716 &  x725 &  x728 &  x731 &  x737 &  x743 &  x746 &  x752 &  x755 &  x758 &  x761 &  x785 &  x788 &  x797 &  x800 &  x803 &  x806 &  x812 &  x815 &  x821 &  x824 &  x830 &  x833 &  x836 &  x848 &  x860 &  x863 &  x866 &  x872 &  x875 &  x884 &  x887 &  x896 &  x899 &  x902 &  x905 &  x907 &  x917 &  x923 &  x926 &  x929 &  x932 &  x938 &  x947 &  x956 &  x959 &  x962 &  x968 &  x974 &  x983 &  x986 &  x995 &  x998 &  x1013 &  x1016 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1043 &  x1049 &  x1058 &  x1064 &  x1067 &  x1076 &  x1082 &  x1088 &  x1094 &  x1097 &  x1103 &  x1115 &  x1124 &  x1127 & ~x297 & ~x336 & ~x357 & ~x375 & ~x432 & ~x435 & ~x510 & ~x550 & ~x588 & ~x627 & ~x666;
assign c272 =  x2 &  x5 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x98 &  x101 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x137 &  x143 &  x149 &  x152 &  x155 &  x158 &  x160 &  x164 &  x167 &  x170 &  x173 &  x179 &  x182 &  x185 &  x191 &  x194 &  x196 &  x199 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x230 &  x233 &  x235 &  x236 &  x238 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x269 &  x272 &  x274 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x308 &  x311 &  x313 &  x317 &  x323 &  x326 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x395 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x431 &  x434 &  x437 &  x440 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x533 &  x539 &  x542 &  x545 &  x548 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x605 &  x611 &  x614 &  x617 &  x619 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x689 &  x692 &  x695 &  x698 &  x704 &  x710 &  x713 &  x718 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x757 &  x758 &  x761 &  x764 &  x770 &  x773 &  x776 &  x779 &  x785 &  x788 &  x794 &  x797 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x878 &  x881 &  x884 &  x887 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1000 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1039 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1078 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x396 & ~x435 & ~x474 & ~x513 & ~x627 & ~x666 & ~x744 & ~x783 & ~x822 & ~x861 & ~x936;
assign c274 =  x2 &  x8 &  x11 &  x14 &  x20 &  x26 &  x35 &  x44 &  x47 &  x50 &  x56 &  x59 &  x62 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x104 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x131 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x200 &  x203 &  x206 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x239 &  x242 &  x248 &  x251 &  x263 &  x266 &  x269 &  x272 &  x275 &  x281 &  x284 &  x287 &  x293 &  x296 &  x302 &  x308 &  x311 &  x317 &  x320 &  x323 &  x332 &  x341 &  x344 &  x350 &  x352 &  x356 &  x359 &  x362 &  x368 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x412 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x434 &  x446 &  x452 &  x458 &  x464 &  x476 &  x479 &  x485 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x524 &  x527 &  x530 &  x536 &  x557 &  x563 &  x575 &  x578 &  x581 &  x584 &  x590 &  x593 &  x596 &  x599 &  x601 &  x602 &  x605 &  x608 &  x614 &  x620 &  x626 &  x629 &  x632 &  x638 &  x639 &  x650 &  x653 &  x659 &  x665 &  x671 &  x683 &  x692 &  x704 &  x707 &  x710 &  x725 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x761 &  x763 &  x770 &  x773 &  x779 &  x782 &  x791 &  x797 &  x800 &  x802 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x827 &  x830 &  x836 &  x839 &  x847 &  x848 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x938 &  x941 &  x947 &  x950 &  x956 &  x959 &  x962 &  x968 &  x971 &  x977 &  x980 &  x983 &  x986 &  x995 &  x1007 &  x1013 &  x1019 &  x1022 &  x1031 &  x1034 &  x1043 &  x1061 &  x1064 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1097 &  x1100 &  x1106 &  x1115 &  x1121 &  x1127 &  x1130 & ~x324 & ~x363 & ~x519 & ~x588 & ~x627;
assign c276 =  x2 &  x5 &  x8 &  x11 &  x17 &  x20 &  x23 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x116 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x194 &  x197 &  x200 &  x202 &  x203 &  x206 &  x212 &  x218 &  x221 &  x227 &  x230 &  x233 &  x239 &  x241 &  x242 &  x245 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x316 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x352 &  x355 &  x356 &  x359 &  x362 &  x368 &  x371 &  x374 &  x377 &  x383 &  x386 &  x389 &  x391 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x464 &  x467 &  x469 &  x473 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x509 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x614 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x689 &  x692 &  x698 &  x701 &  x704 &  x707 &  x710 &  x716 &  x719 &  x722 &  x725 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x782 &  x785 &  x788 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x821 &  x824 &  x827 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x869 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x0 & ~x39 & ~x78 & ~x117 & ~x363 & ~x402 & ~x441 & ~x480 & ~x519 & ~x627 & ~x666 & ~x705 & ~x783 & ~x822;
assign c278 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x26 &  x29 &  x35 &  x47 &  x50 &  x53 &  x59 &  x62 &  x65 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x116 &  x125 &  x128 &  x137 &  x140 &  x143 &  x146 &  x149 &  x154 &  x155 &  x161 &  x167 &  x182 &  x185 &  x187 &  x188 &  x191 &  x194 &  x197 &  x200 &  x202 &  x203 &  x209 &  x214 &  x215 &  x218 &  x220 &  x224 &  x226 &  x227 &  x236 &  x241 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x269 &  x272 &  x278 &  x287 &  x296 &  x299 &  x305 &  x308 &  x311 &  x317 &  x319 &  x326 &  x329 &  x337 &  x341 &  x350 &  x353 &  x358 &  x365 &  x377 &  x380 &  x392 &  x395 &  x407 &  x409 &  x410 &  x413 &  x419 &  x425 &  x431 &  x440 &  x443 &  x449 &  x455 &  x461 &  x464 &  x470 &  x479 &  x482 &  x488 &  x491 &  x497 &  x500 &  x503 &  x506 &  x512 &  x515 &  x518 &  x530 &  x533 &  x551 &  x554 &  x563 &  x566 &  x572 &  x593 &  x596 &  x599 &  x602 &  x605 &  x611 &  x614 &  x617 &  x623 &  x626 &  x629 &  x635 &  x641 &  x644 &  x650 &  x656 &  x659 &  x668 &  x671 &  x683 &  x692 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x724 &  x728 &  x737 &  x743 &  x746 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x779 &  x782 &  x785 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x821 &  x824 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x872 &  x877 &  x878 &  x881 &  x884 &  x887 &  x902 &  x905 &  x908 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x935 &  x941 &  x944 &  x947 &  x956 &  x959 &  x962 &  x971 &  x980 &  x986 &  x989 &  x992 &  x998 &  x1001 &  x1013 &  x1022 &  x1025 &  x1046 &  x1052 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1109 &  x1115 &  x1121 &  x1124 &  x1130 & ~x195 & ~x234 & ~x273 & ~x312;
assign c280 =  x2 &  x5 &  x14 &  x17 &  x20 &  x23 &  x32 &  x47 &  x50 &  x53 &  x56 &  x62 &  x65 &  x71 &  x74 &  x83 &  x86 &  x89 &  x98 &  x101 &  x116 &  x119 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x155 &  x158 &  x161 &  x164 &  x182 &  x194 &  x212 &  x221 &  x224 &  x227 &  x236 &  x242 &  x245 &  x254 &  x260 &  x275 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x305 &  x308 &  x311 &  x316 &  x326 &  x329 &  x338 &  x341 &  x350 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x380 &  x383 &  x389 &  x392 &  x401 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x430 &  x437 &  x440 &  x446 &  x449 &  x461 &  x464 &  x469 &  x473 &  x479 &  x482 &  x497 &  x503 &  x508 &  x523 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x551 &  x557 &  x572 &  x578 &  x584 &  x593 &  x601 &  x617 &  x620 &  x623 &  x626 &  x632 &  x638 &  x640 &  x647 &  x653 &  x659 &  x665 &  x679 &  x683 &  x689 &  x692 &  x695 &  x710 &  x713 &  x716 &  x718 &  x719 &  x728 &  x731 &  x734 &  x743 &  x746 &  x749 &  x770 &  x779 &  x782 &  x788 &  x796 &  x797 &  x800 &  x809 &  x812 &  x815 &  x827 &  x833 &  x835 &  x839 &  x842 &  x851 &  x854 &  x860 &  x875 &  x890 &  x908 &  x911 &  x914 &  x920 &  x929 &  x935 &  x938 &  x941 &  x944 &  x953 &  x959 &  x965 &  x968 &  x974 &  x989 &  x1004 &  x1013 &  x1016 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1052 &  x1055 &  x1064 &  x1067 &  x1070 &  x1076 &  x1082 &  x1088 &  x1103 &  x1106 &  x1118 &  x1121 &  x1124 &  x1130 & ~x519 & ~x558 & ~x591 & ~x630 & ~x669 & ~x714 & ~x753;
assign c282 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x43 &  x44 &  x47 &  x49 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x79 &  x80 &  x82 &  x83 &  x86 &  x88 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x121 &  x122 &  x125 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x157 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x196 &  x197 &  x200 &  x203 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x230 &  x233 &  x235 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x274 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x305 &  x308 &  x311 &  x313 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x346 &  x347 &  x350 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x380 &  x383 &  x385 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x674 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x69 & ~x108 & ~x129 & ~x147 & ~x168 & ~x207 & ~x246 & ~x285 & ~x297 & ~x627 & ~x666 & ~x705 & ~x744 & ~x939;
assign c284 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x257 &  x260 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x511 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x549 &  x550 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x589 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x697 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x736 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x775 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130 & ~x156 & ~x195 & ~x234 & ~x273 & ~x648 & ~x687 & ~x726 & ~x765;
assign c286 =  x2 &  x29 &  x44 &  x50 &  x59 &  x62 &  x74 &  x77 &  x80 &  x83 &  x110 &  x125 &  x131 &  x140 &  x149 &  x152 &  x158 &  x164 &  x179 &  x191 &  x194 &  x206 &  x212 &  x224 &  x227 &  x242 &  x245 &  x251 &  x254 &  x257 &  x260 &  x266 &  x269 &  x275 &  x278 &  x287 &  x293 &  x296 &  x299 &  x308 &  x317 &  x326 &  x332 &  x335 &  x344 &  x347 &  x350 &  x356 &  x359 &  x365 &  x368 &  x383 &  x386 &  x416 &  x419 &  x428 &  x437 &  x443 &  x446 &  x452 &  x455 &  x458 &  x463 &  x479 &  x494 &  x502 &  x503 &  x506 &  x509 &  x515 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x545 &  x548 &  x554 &  x560 &  x563 &  x566 &  x569 &  x578 &  x593 &  x602 &  x605 &  x608 &  x620 &  x626 &  x629 &  x632 &  x635 &  x638 &  x644 &  x647 &  x656 &  x662 &  x677 &  x680 &  x686 &  x695 &  x707 &  x718 &  x725 &  x728 &  x734 &  x743 &  x746 &  x749 &  x757 &  x758 &  x764 &  x782 &  x785 &  x788 &  x796 &  x797 &  x806 &  x815 &  x833 &  x845 &  x848 &  x866 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x914 &  x923 &  x929 &  x941 &  x947 &  x953 &  x962 &  x968 &  x971 &  x977 &  x980 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1022 &  x1025 &  x1028 &  x1031 &  x1043 &  x1067 & ~x66 & ~x105 & ~x184 & ~x222 & ~x300;
assign c288 =  x5 &  x8 &  x11 &  x14 &  x17 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x44 &  x47 &  x50 &  x56 &  x59 &  x62 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x401 &  x404 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x601 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x640 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x677 &  x679 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x718 &  x719 &  x722 &  x725 &  x728 &  x731 &  x733 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x757 &  x758 &  x761 &  x764 &  x767 &  x770 &  x771 &  x772 &  x773 &  x776 &  x779 &  x782 &  x788 &  x791 &  x794 &  x796 &  x797 &  x800 &  x803 &  x806 &  x809 &  x811 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x835 &  x836 &  x839 &  x842 &  x848 &  x850 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x874 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x441 & ~x480 & ~x675;
assign c290 =  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x77 &  x83 &  x86 &  x89 &  x92 &  x98 &  x101 &  x107 &  x110 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x137 &  x140 &  x143 &  x146 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x176 &  x179 &  x182 &  x185 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x224 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x299 &  x302 &  x308 &  x314 &  x317 &  x320 &  x323 &  x329 &  x335 &  x338 &  x341 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x464 &  x467 &  x470 &  x472 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x503 &  x509 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x545 &  x550 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x701 &  x704 &  x707 &  x710 &  x713 &  x719 &  x725 &  x731 &  x734 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x773 &  x776 &  x782 &  x785 &  x794 &  x806 &  x809 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x845 &  x848 &  x851 &  x854 &  x863 &  x866 &  x872 &  x875 &  x878 &  x884 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x944 &  x947 &  x950 &  x953 &  x959 &  x962 &  x965 &  x968 &  x980 &  x983 &  x989 &  x998 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1130 & ~x492 & ~x531 & ~x571 & ~x594 & ~x609 & ~x633 & ~x672 & ~x687 & ~x726 & ~x765 & ~x804 & ~x843 & ~x861 & ~x882 & ~x900 & ~x921;
assign c292 =  x2 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x107 &  x110 &  x116 &  x122 &  x125 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x164 &  x167 &  x170 &  x176 &  x179 &  x182 &  x185 &  x191 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x227 &  x230 &  x233 &  x242 &  x245 &  x248 &  x251 &  x257 &  x263 &  x266 &  x275 &  x278 &  x281 &  x290 &  x293 &  x296 &  x299 &  x305 &  x308 &  x311 &  x314 &  x320 &  x323 &  x326 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x362 &  x371 &  x374 &  x377 &  x380 &  x389 &  x395 &  x398 &  x401 &  x404 &  x419 &  x422 &  x425 &  x428 &  x434 &  x440 &  x446 &  x449 &  x455 &  x461 &  x464 &  x467 &  x470 &  x473 &  x479 &  x482 &  x485 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x548 &  x554 &  x557 &  x560 &  x569 &  x572 &  x578 &  x581 &  x584 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x650 &  x653 &  x659 &  x662 &  x665 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x689 &  x695 &  x704 &  x710 &  x713 &  x716 &  x725 &  x728 &  x731 &  x740 &  x743 &  x746 &  x752 &  x755 &  x758 &  x764 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x803 &  x809 &  x812 &  x815 &  x818 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x848 &  x851 &  x857 &  x860 &  x863 &  x869 &  x872 &  x884 &  x887 &  x890 &  x893 &  x896 &  x908 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x950 &  x956 &  x959 &  x965 &  x968 &  x971 &  x977 &  x980 &  x983 &  x992 &  x998 &  x1001 &  x1007 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1046 &  x1055 &  x1061 &  x1064 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1091 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x396 & ~x510 & ~x546 & ~x549 & ~x585 & ~x645 & ~x646 & ~x804;
assign c294 =  x2 &  x11 &  x14 &  x17 &  x20 &  x23 &  x29 &  x32 &  x35 &  x38 &  x41 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x83 &  x86 &  x89 &  x92 &  x98 &  x104 &  x107 &  x110 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x179 &  x182 &  x185 &  x188 &  x191 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x316 &  x317 &  x320 &  x323 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x389 &  x391 &  x392 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x437 &  x440 &  x443 &  x446 &  x452 &  x458 &  x461 &  x464 &  x467 &  x473 &  x476 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x542 &  x545 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x584 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x611 &  x614 &  x617 &  x620 &  x623 &  x632 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x794 &  x800 &  x803 &  x806 &  x809 &  x812 &  x818 &  x821 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x845 &  x848 &  x854 &  x857 &  x860 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x902 &  x914 &  x917 &  x920 &  x926 &  x929 &  x932 &  x938 &  x944 &  x947 &  x953 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1043 &  x1046 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x261 & ~x300 & ~x339 & ~x375 & ~x378 & ~x414 & ~x453 & ~x492 & ~x531 & ~x585 & ~x624 & ~x666 & ~x705 & ~x726 & ~x744 & ~x783 & ~x822 & ~x975 & ~x1014 & ~x1086;
assign c296 =  x2 &  x5 &  x6 &  x7 &  x8 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x45 &  x46 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x85 &  x86 &  x88 &  x89 &  x92 &  x95 &  x98 &  x104 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x127 &  x128 &  x131 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x238 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x272 &  x275 &  x277 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x316 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x355 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x398 &  x401 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x593 &  x596 &  x599 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x640 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x679 &  x680 &  x683 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x718 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x757 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x775 &  x776 &  x779 &  x782 &  x785 &  x788 &  x794 &  x796 &  x797 &  x800 &  x803 &  x809 &  x812 &  x814 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x835 &  x836 &  x839 &  x842 &  x845 &  x848 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x874 &  x875 &  x878 &  x884 &  x887 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x913 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130;
assign c298 =  x2 &  x8 &  x11 &  x17 &  x23 &  x32 &  x35 &  x47 &  x50 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x77 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x122 &  x125 &  x131 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x170 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x197 &  x200 &  x203 &  x206 &  x212 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x251 &  x254 &  x257 &  x263 &  x266 &  x269 &  x272 &  x275 &  x281 &  x283 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x308 &  x314 &  x316 &  x317 &  x326 &  x329 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x368 &  x371 &  x377 &  x380 &  x383 &  x386 &  x389 &  x391 &  x392 &  x395 &  x398 &  x401 &  x404 &  x410 &  x422 &  x425 &  x428 &  x430 &  x431 &  x434 &  x437 &  x443 &  x449 &  x452 &  x455 &  x458 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x491 &  x497 &  x500 &  x502 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x545 &  x548 &  x557 &  x560 &  x563 &  x569 &  x578 &  x581 &  x584 &  x587 &  x590 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x623 &  x626 &  x629 &  x635 &  x637 &  x644 &  x647 &  x650 &  x653 &  x656 &  x658 &  x659 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x704 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x764 &  x767 &  x770 &  x782 &  x785 &  x794 &  x797 &  x806 &  x809 &  x812 &  x821 &  x824 &  x827 &  x833 &  x836 &  x851 &  x866 &  x869 &  x872 &  x875 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x920 &  x923 &  x926 &  x929 &  x935 &  x938 &  x941 &  x944 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1019 &  x1025 &  x1034 &  x1037 &  x1043 &  x1049 &  x1055 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x381 & ~x382 & ~x420 & ~x498 & ~x783;
assign c2100 =  x2 &  x5 &  x7 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x46 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x85 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x124 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x39 & ~x78 & ~x117 & ~x690 & ~x729 & ~x840 & ~x879 & ~x918 & ~x957 & ~x958 & ~x996 & ~x999 & ~x1035 & ~x1113;
assign c2102 =  x2 &  x3 &  x4 &  x5 &  x8 &  x10 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x41 &  x42 &  x43 &  x44 &  x47 &  x49 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x77 &  x80 &  x82 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x119 &  x121 &  x122 &  x125 &  x128 &  x134 &  x137 &  x140 &  x152 &  x158 &  x160 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x197 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x278 &  x281 &  x284 &  x290 &  x293 &  x296 &  x299 &  x302 &  x308 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x338 &  x344 &  x347 &  x350 &  x353 &  x359 &  x362 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x410 &  x413 &  x419 &  x422 &  x425 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x458 &  x461 &  x464 &  x467 &  x470 &  x476 &  x479 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x524 &  x530 &  x533 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x560 &  x563 &  x566 &  x572 &  x575 &  x578 &  x581 &  x587 &  x593 &  x599 &  x602 &  x605 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x638 &  x641 &  x647 &  x650 &  x653 &  x659 &  x662 &  x665 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x695 &  x698 &  x704 &  x707 &  x710 &  x716 &  x719 &  x725 &  x728 &  x731 &  x734 &  x743 &  x746 &  x749 &  x752 &  x758 &  x764 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x797 &  x800 &  x812 &  x815 &  x818 &  x824 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x878 &  x881 &  x884 &  x887 &  x890 &  x899 &  x902 &  x905 &  x911 &  x914 &  x920 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x950 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x977 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1052 &  x1055 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1130 & ~x471 & ~x510 & ~x549 & ~x550 & ~x588 & ~x627 & ~x666 & ~x702 & ~x705 & ~x741;
assign c2104 =  x5 &  x8 &  x11 &  x26 &  x28 &  x29 &  x44 &  x47 &  x50 &  x53 &  x55 &  x59 &  x62 &  x65 &  x80 &  x88 &  x89 &  x94 &  x98 &  x100 &  x101 &  x119 &  x122 &  x127 &  x128 &  x131 &  x133 &  x134 &  x137 &  x143 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x182 &  x184 &  x188 &  x191 &  x203 &  x212 &  x230 &  x236 &  x239 &  x241 &  x245 &  x248 &  x260 &  x278 &  x281 &  x284 &  x287 &  x295 &  x302 &  x308 &  x311 &  x314 &  x320 &  x329 &  x338 &  x341 &  x356 &  x362 &  x365 &  x368 &  x374 &  x380 &  x383 &  x386 &  x395 &  x398 &  x401 &  x404 &  x407 &  x413 &  x416 &  x431 &  x434 &  x437 &  x443 &  x458 &  x461 &  x467 &  x479 &  x485 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x512 &  x515 &  x518 &  x521 &  x527 &  x536 &  x551 &  x554 &  x557 &  x569 &  x575 &  x584 &  x587 &  x590 &  x596 &  x602 &  x611 &  x614 &  x620 &  x623 &  x626 &  x629 &  x635 &  x644 &  x653 &  x665 &  x668 &  x671 &  x674 &  x680 &  x692 &  x695 &  x698 &  x710 &  x716 &  x722 &  x725 &  x731 &  x734 &  x740 &  x746 &  x755 &  x758 &  x764 &  x773 &  x779 &  x782 &  x794 &  x797 &  x800 &  x806 &  x809 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x851 &  x857 &  x874 &  x875 &  x878 &  x881 &  x890 &  x892 &  x893 &  x896 &  x908 &  x913 &  x914 &  x917 &  x923 &  x932 &  x935 &  x944 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x977 &  x980 &  x986 &  x989 &  x991 &  x992 &  x1003 &  x1004 &  x1010 &  x1016 &  x1019 &  x1034 &  x1040 &  x1046 &  x1055 &  x1058 &  x1061 &  x1076 &  x1091 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1127 &  x1130 & ~x480 & ~x861;
assign c2106 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x143 &  x146 &  x149 &  x155 &  x161 &  x164 &  x167 &  x170 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x317 &  x319 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x353 &  x356 &  x359 &  x374 &  x377 &  x380 &  x383 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x464 &  x467 &  x470 &  x473 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x509 &  x511 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x542 &  x545 &  x548 &  x550 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x635 &  x638 &  x644 &  x647 &  x650 &  x656 &  x659 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x770 &  x773 &  x776 &  x779 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x9 & ~x48 & ~x156 & ~x195 & ~x306 & ~x558 & ~x597 & ~x753 & ~x900;
assign c2108 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x433 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x476 &  x479 &  x482 &  x485 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x156 & ~x195 & ~x234 & ~x453 & ~x492 & ~x531 & ~x534 & ~x570 & ~x609 & ~x648 & ~x687 & ~x747 & ~x765 & ~x804 & ~x843 & ~x900;
assign c2110 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x43 &  x47 &  x50 &  x56 &  x59 &  x62 &  x65 &  x68 &  x74 &  x77 &  x80 &  x82 &  x86 &  x92 &  x101 &  x104 &  x107 &  x113 &  x116 &  x119 &  x121 &  x122 &  x125 &  x128 &  x131 &  x137 &  x140 &  x149 &  x152 &  x155 &  x160 &  x164 &  x170 &  x173 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x196 &  x197 &  x200 &  x206 &  x209 &  x212 &  x215 &  x221 &  x227 &  x233 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x305 &  x307 &  x308 &  x311 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x345 &  x346 &  x347 &  x350 &  x353 &  x362 &  x371 &  x374 &  x380 &  x383 &  x384 &  x385 &  x386 &  x389 &  x392 &  x398 &  x401 &  x407 &  x410 &  x413 &  x416 &  x422 &  x423 &  x424 &  x431 &  x437 &  x440 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x463 &  x464 &  x467 &  x470 &  x476 &  x479 &  x485 &  x488 &  x491 &  x494 &  x500 &  x506 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x548 &  x554 &  x557 &  x563 &  x566 &  x569 &  x572 &  x581 &  x584 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x620 &  x629 &  x632 &  x635 &  x638 &  x641 &  x650 &  x656 &  x662 &  x671 &  x674 &  x686 &  x689 &  x704 &  x707 &  x722 &  x728 &  x731 &  x737 &  x749 &  x752 &  x755 &  x758 &  x761 &  x767 &  x770 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x806 &  x809 &  x812 &  x815 &  x818 &  x833 &  x839 &  x845 &  x851 &  x854 &  x860 &  x863 &  x869 &  x872 &  x875 &  x878 &  x884 &  x887 &  x890 &  x896 &  x902 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x938 &  x941 &  x947 &  x950 &  x953 &  x968 &  x977 &  x986 &  x989 &  x992 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1022 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1055 &  x1061 &  x1064 &  x1073 &  x1076 &  x1082 &  x1094 &  x1106 &  x1112 &  x1118 &  x1121 &  x1124 &  x1130 & ~x54 & ~x549 & ~x627;
assign c2112 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x277 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x314 &  x316 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x542 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x375 & ~x396 & ~x414 & ~x438 & ~x453 & ~x477 & ~x516 & ~x552 & ~x627 & ~x666 & ~x705 & ~x744 & ~x783 & ~x822 & ~x936 & ~x975 & ~x1014 & ~x1092;
assign c2114 =  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x131 &  x134 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x167 &  x170 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x430 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x476 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x635 &  x640 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x757 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x796 &  x797 &  x800 &  x806 &  x809 &  x812 &  x815 &  x818 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x902 &  x905 &  x908 &  x911 &  x913 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x952 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x989 &  x991 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1028 &  x1030 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x402 & ~x403 & ~x480 & ~x519 & ~x627 & ~x666 & ~x667 & ~x705 & ~x706 & ~x783 & ~x822 & ~x861;
assign c2116 =  x2 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x59 &  x65 &  x74 &  x80 &  x83 &  x86 &  x92 &  x98 &  x119 &  x125 &  x128 &  x134 &  x137 &  x140 &  x149 &  x155 &  x161 &  x164 &  x170 &  x179 &  x200 &  x209 &  x218 &  x221 &  x233 &  x236 &  x239 &  x242 &  x245 &  x251 &  x257 &  x266 &  x272 &  x275 &  x278 &  x290 &  x299 &  x302 &  x305 &  x310 &  x320 &  x326 &  x329 &  x335 &  x344 &  x347 &  x350 &  x364 &  x374 &  x377 &  x383 &  x386 &  x389 &  x401 &  x403 &  x407 &  x410 &  x416 &  x422 &  x425 &  x431 &  x434 &  x437 &  x442 &  x449 &  x452 &  x461 &  x473 &  x476 &  x481 &  x482 &  x487 &  x488 &  x491 &  x494 &  x497 &  x500 &  x505 &  x515 &  x520 &  x524 &  x526 &  x530 &  x533 &  x539 &  x545 &  x548 &  x557 &  x559 &  x560 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x587 &  x593 &  x598 &  x602 &  x605 &  x617 &  x626 &  x629 &  x632 &  x638 &  x643 &  x644 &  x647 &  x656 &  x668 &  x674 &  x676 &  x677 &  x680 &  x689 &  x698 &  x707 &  x710 &  x712 &  x719 &  x722 &  x728 &  x746 &  x749 &  x752 &  x758 &  x761 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x794 &  x797 &  x800 &  x803 &  x809 &  x815 &  x821 &  x824 &  x827 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x863 &  x866 &  x869 &  x872 &  x878 &  x881 &  x884 &  x887 &  x899 &  x902 &  x914 &  x917 &  x920 &  x926 &  x929 &  x932 &  x944 &  x947 &  x953 &  x956 &  x959 &  x962 &  x968 &  x971 &  x986 &  x989 &  x992 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1055 &  x1058 &  x1067 &  x1070 &  x1076 &  x1079 &  x1088 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1130 & ~x222 & ~x261 & ~x624 & ~x663;
assign c2118 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x35 &  x38 &  x41 &  x44 &  x47 &  x53 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x104 &  x107 &  x110 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x209 &  x212 &  x215 &  x218 &  x220 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x251 &  x254 &  x257 &  x263 &  x266 &  x269 &  x272 &  x275 &  x284 &  x287 &  x290 &  x296 &  x302 &  x305 &  x308 &  x311 &  x320 &  x323 &  x326 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x365 &  x371 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x407 &  x409 &  x413 &  x416 &  x422 &  x425 &  x431 &  x437 &  x439 &  x443 &  x452 &  x458 &  x461 &  x464 &  x470 &  x473 &  x478 &  x479 &  x482 &  x485 &  x488 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x707 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x740 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x779 &  x782 &  x785 &  x791 &  x794 &  x797 &  x803 &  x806 &  x809 &  x812 &  x818 &  x820 &  x821 &  x824 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x898 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x937 &  x938 &  x944 &  x950 &  x953 &  x956 &  x968 &  x971 &  x974 &  x977 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1073 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x903 & ~x942 & ~x1020 & ~x1021 & ~x1038 & ~x1077 & ~x1116;
assign c2120 =  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x41 &  x44 &  x47 &  x50 &  x56 &  x62 &  x65 &  x68 &  x71 &  x74 &  x83 &  x86 &  x89 &  x98 &  x101 &  x113 &  x116 &  x119 &  x128 &  x131 &  x137 &  x140 &  x143 &  x149 &  x152 &  x155 &  x164 &  x167 &  x170 &  x176 &  x182 &  x185 &  x188 &  x197 &  x209 &  x215 &  x218 &  x221 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x244 &  x245 &  x248 &  x251 &  x260 &  x263 &  x269 &  x272 &  x275 &  x284 &  x287 &  x296 &  x302 &  x305 &  x308 &  x313 &  x314 &  x316 &  x320 &  x323 &  x329 &  x338 &  x344 &  x347 &  x352 &  x365 &  x374 &  x380 &  x383 &  x389 &  x391 &  x392 &  x401 &  x404 &  x407 &  x410 &  x416 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x470 &  x476 &  x479 &  x482 &  x488 &  x491 &  x494 &  x497 &  x503 &  x506 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x545 &  x551 &  x554 &  x557 &  x560 &  x569 &  x572 &  x578 &  x581 &  x599 &  x602 &  x611 &  x617 &  x620 &  x629 &  x635 &  x641 &  x647 &  x650 &  x653 &  x656 &  x668 &  x671 &  x674 &  x680 &  x686 &  x689 &  x695 &  x698 &  x704 &  x716 &  x719 &  x722 &  x725 &  x734 &  x737 &  x740 &  x749 &  x758 &  x761 &  x770 &  x776 &  x779 &  x785 &  x788 &  x794 &  x797 &  x803 &  x821 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x854 &  x860 &  x863 &  x866 &  x878 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x941 &  x944 &  x959 &  x971 &  x977 &  x980 &  x983 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1127 &  x1130 & ~x261 & ~x300 & ~x301 & ~x339 & ~x340 & ~x705 & ~x744 & ~x975 & ~x1002 & ~x1008 & ~x1014 & ~x1041 & ~x1047 & ~x1125;
assign c2122 =  x5 &  x8 &  x11 &  x17 &  x23 &  x26 &  x32 &  x35 &  x38 &  x41 &  x47 &  x50 &  x53 &  x56 &  x62 &  x71 &  x74 &  x80 &  x83 &  x85 &  x92 &  x95 &  x101 &  x104 &  x110 &  x119 &  x122 &  x124 &  x125 &  x128 &  x131 &  x134 &  x137 &  x146 &  x152 &  x155 &  x158 &  x161 &  x163 &  x167 &  x170 &  x173 &  x179 &  x185 &  x188 &  x199 &  x200 &  x201 &  x202 &  x203 &  x206 &  x209 &  x212 &  x215 &  x227 &  x236 &  x238 &  x239 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x269 &  x272 &  x278 &  x281 &  x284 &  x287 &  x290 &  x296 &  x302 &  x305 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x344 &  x353 &  x355 &  x359 &  x362 &  x365 &  x374 &  x383 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x449 &  x455 &  x458 &  x461 &  x467 &  x470 &  x473 &  x476 &  x485 &  x488 &  x494 &  x497 &  x500 &  x503 &  x512 &  x515 &  x518 &  x524 &  x533 &  x539 &  x542 &  x545 &  x548 &  x554 &  x557 &  x560 &  x566 &  x569 &  x572 &  x581 &  x590 &  x596 &  x599 &  x605 &  x611 &  x614 &  x620 &  x623 &  x629 &  x640 &  x641 &  x644 &  x653 &  x662 &  x665 &  x674 &  x677 &  x689 &  x694 &  x695 &  x698 &  x704 &  x707 &  x710 &  x713 &  x719 &  x722 &  x725 &  x728 &  x731 &  x733 &  x734 &  x737 &  x740 &  x749 &  x755 &  x758 &  x761 &  x767 &  x772 &  x773 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x809 &  x811 &  x812 &  x818 &  x821 &  x833 &  x842 &  x848 &  x854 &  x857 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x935 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x971 &  x974 &  x977 &  x986 &  x989 &  x992 &  x998 &  x1013 &  x1016 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1091 &  x1094 &  x1097 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 & ~x741;
assign c2124 =  x2 &  x11 &  x14 &  x17 &  x26 &  x29 &  x32 &  x41 &  x47 &  x50 &  x56 &  x62 &  x68 &  x77 &  x83 &  x89 &  x110 &  x113 &  x119 &  x125 &  x128 &  x134 &  x146 &  x149 &  x152 &  x155 &  x158 &  x160 &  x161 &  x164 &  x167 &  x176 &  x188 &  x191 &  x197 &  x200 &  x209 &  x215 &  x221 &  x233 &  x238 &  x242 &  x248 &  x254 &  x260 &  x263 &  x272 &  x277 &  x281 &  x293 &  x296 &  x302 &  x305 &  x311 &  x326 &  x332 &  x335 &  x338 &  x341 &  x347 &  x356 &  x370 &  x371 &  x380 &  x383 &  x392 &  x395 &  x398 &  x404 &  x410 &  x413 &  x416 &  x425 &  x428 &  x434 &  x437 &  x440 &  x446 &  x448 &  x452 &  x458 &  x464 &  x467 &  x470 &  x476 &  x479 &  x481 &  x482 &  x500 &  x503 &  x506 &  x509 &  x512 &  x518 &  x520 &  x521 &  x524 &  x526 &  x536 &  x539 &  x542 &  x548 &  x554 &  x557 &  x566 &  x575 &  x578 &  x581 &  x584 &  x593 &  x596 &  x605 &  x614 &  x617 &  x629 &  x637 &  x641 &  x643 &  x644 &  x647 &  x653 &  x656 &  x659 &  x677 &  x680 &  x682 &  x689 &  x692 &  x698 &  x707 &  x713 &  x719 &  x724 &  x728 &  x737 &  x749 &  x755 &  x767 &  x770 &  x773 &  x776 &  x782 &  x785 &  x788 &  x791 &  x809 &  x812 &  x818 &  x821 &  x827 &  x830 &  x842 &  x845 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x878 &  x887 &  x902 &  x908 &  x911 &  x917 &  x923 &  x929 &  x932 &  x941 &  x944 &  x947 &  x953 &  x959 &  x962 &  x968 &  x980 &  x992 &  x998 &  x1001 &  x1010 &  x1013 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1052 &  x1058 &  x1061 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1100 &  x1103 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x1113;
assign c2126 =  x20 &  x32 &  x35 &  x40 &  x53 &  x71 &  x74 &  x77 &  x110 &  x113 &  x121 &  x125 &  x128 &  x143 &  x158 &  x164 &  x170 &  x179 &  x194 &  x200 &  x203 &  x215 &  x224 &  x230 &  x233 &  x245 &  x251 &  x260 &  x272 &  x281 &  x284 &  x302 &  x307 &  x313 &  x323 &  x326 &  x329 &  x341 &  x344 &  x345 &  x346 &  x350 &  x356 &  x359 &  x362 &  x371 &  x374 &  x385 &  x401 &  x407 &  x413 &  x425 &  x434 &  x449 &  x452 &  x473 &  x482 &  x485 &  x500 &  x503 &  x518 &  x521 &  x533 &  x545 &  x548 &  x575 &  x581 &  x593 &  x605 &  x623 &  x626 &  x629 &  x635 &  x656 &  x674 &  x689 &  x701 &  x704 &  x710 &  x716 &  x719 &  x722 &  x734 &  x743 &  x749 &  x755 &  x767 &  x788 &  x812 &  x836 &  x851 &  x857 &  x860 &  x863 &  x869 &  x872 &  x874 &  x884 &  x887 &  x890 &  x896 &  x905 &  x908 &  x917 &  x920 &  x926 &  x932 &  x938 &  x941 &  x952 &  x956 &  x962 &  x965 &  x974 &  x977 &  x980 &  x983 &  x988 &  x992 &  x1007 &  x1013 &  x1025 &  x1027 &  x1028 &  x1030 &  x1046 &  x1049 &  x1052 &  x1058 &  x1064 &  x1067 &  x1069 &  x1073 &  x1091 &  x1094 &  x1097 &  x1103 &  x1118 &  x1130 & ~x297 & ~x627 & ~x744 & ~x783;
assign c2128 =  x2 &  x5 &  x11 &  x14 &  x38 &  x47 &  x59 &  x74 &  x86 &  x95 &  x98 &  x101 &  x113 &  x122 &  x125 &  x134 &  x137 &  x140 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x173 &  x176 &  x188 &  x194 &  x200 &  x209 &  x212 &  x215 &  x218 &  x221 &  x230 &  x233 &  x236 &  x239 &  x248 &  x254 &  x257 &  x263 &  x269 &  x272 &  x275 &  x293 &  x296 &  x299 &  x302 &  x317 &  x319 &  x323 &  x326 &  x329 &  x338 &  x359 &  x383 &  x392 &  x398 &  x401 &  x404 &  x407 &  x425 &  x428 &  x431 &  x437 &  x446 &  x449 &  x461 &  x473 &  x491 &  x494 &  x497 &  x512 &  x524 &  x533 &  x542 &  x545 &  x548 &  x554 &  x560 &  x575 &  x581 &  x584 &  x596 &  x608 &  x620 &  x623 &  x626 &  x629 &  x638 &  x641 &  x650 &  x659 &  x686 &  x692 &  x701 &  x704 &  x713 &  x722 &  x728 &  x743 &  x749 &  x752 &  x758 &  x761 &  x770 &  x773 &  x776 &  x785 &  x809 &  x815 &  x827 &  x830 &  x842 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x872 &  x881 &  x896 &  x899 &  x902 &  x905 &  x917 &  x929 &  x938 &  x941 &  x944 &  x950 &  x965 &  x968 &  x971 &  x977 &  x989 &  x1001 &  x1025 &  x1028 &  x1034 &  x1040 &  x1043 &  x1061 &  x1073 &  x1088 &  x1100 &  x1109 &  x1121 &  x1124 & ~x198 & ~x558 & ~x648 & ~x669 & ~x675 & ~x792 & ~x900 & ~x939 & ~x978 & ~x981 & ~x1056;
assign c2130 =  x5 &  x14 &  x17 &  x20 &  x29 &  x41 &  x43 &  x47 &  x50 &  x53 &  x56 &  x59 &  x65 &  x68 &  x71 &  x77 &  x82 &  x83 &  x86 &  x98 &  x110 &  x119 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x152 &  x160 &  x167 &  x170 &  x176 &  x179 &  x185 &  x191 &  x196 &  x197 &  x200 &  x206 &  x209 &  x212 &  x218 &  x221 &  x227 &  x236 &  x242 &  x245 &  x248 &  x254 &  x257 &  x260 &  x263 &  x269 &  x272 &  x275 &  x284 &  x299 &  x308 &  x311 &  x317 &  x320 &  x323 &  x329 &  x338 &  x353 &  x356 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x401 &  x406 &  x407 &  x413 &  x425 &  x434 &  x437 &  x443 &  x445 &  x446 &  x449 &  x458 &  x461 &  x464 &  x473 &  x479 &  x484 &  x485 &  x491 &  x497 &  x503 &  x512 &  x518 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x554 &  x572 &  x575 &  x578 &  x584 &  x593 &  x596 &  x599 &  x605 &  x608 &  x617 &  x620 &  x623 &  x626 &  x632 &  x638 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x677 &  x680 &  x686 &  x692 &  x695 &  x707 &  x710 &  x713 &  x719 &  x731 &  x734 &  x737 &  x740 &  x746 &  x749 &  x755 &  x761 &  x767 &  x770 &  x773 &  x779 &  x782 &  x788 &  x794 &  x797 &  x800 &  x806 &  x815 &  x821 &  x848 &  x854 &  x857 &  x860 &  x866 &  x869 &  x872 &  x875 &  x878 &  x884 &  x890 &  x892 &  x893 &  x902 &  x905 &  x908 &  x911 &  x929 &  x931 &  x932 &  x938 &  x944 &  x953 &  x955 &  x956 &  x968 &  x971 &  x977 &  x980 &  x986 &  x989 &  x992 &  x998 &  x1001 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1058 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1097 &  x1103 &  x1112 &  x1115 &  x1127 & ~x207 & ~x246 & ~x279 & ~x285 & ~x507;
assign c2132 =  x2 &  x5 &  x11 &  x14 &  x20 &  x23 &  x29 &  x35 &  x38 &  x41 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x116 &  x119 &  x122 &  x125 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x361 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x400 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x439 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x478 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x542 &  x547 &  x548 &  x551 &  x554 &  x557 &  x560 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x590 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x625 &  x626 &  x629 &  x632 &  x635 &  x638 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x734 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x761 &  x764 &  x767 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x842 &  x845 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x878 &  x881 &  x884 &  x890 &  x893 &  x896 &  x899 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x977 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x495 & ~x498 & ~x537 & ~x861 & ~x888 & ~x900 & ~x927 & ~x978 & ~x1017;
assign c2134 =  x2 &  x8 &  x11 &  x14 &  x20 &  x23 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x62 &  x65 &  x68 &  x77 &  x80 &  x83 &  x89 &  x95 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x122 &  x125 &  x128 &  x134 &  x140 &  x143 &  x146 &  x149 &  x155 &  x158 &  x161 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x251 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x290 &  x293 &  x299 &  x302 &  x305 &  x308 &  x317 &  x320 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x350 &  x356 &  x358 &  x359 &  x362 &  x365 &  x368 &  x377 &  x383 &  x395 &  x397 &  x398 &  x401 &  x404 &  x407 &  x410 &  x419 &  x422 &  x428 &  x431 &  x434 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x473 &  x476 &  x479 &  x482 &  x488 &  x494 &  x500 &  x503 &  x509 &  x512 &  x518 &  x521 &  x536 &  x539 &  x545 &  x548 &  x551 &  x554 &  x557 &  x563 &  x566 &  x572 &  x578 &  x581 &  x584 &  x587 &  x590 &  x599 &  x602 &  x608 &  x611 &  x614 &  x623 &  x626 &  x628 &  x629 &  x632 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x683 &  x686 &  x689 &  x692 &  x698 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x725 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x782 &  x785 &  x788 &  x794 &  x797 &  x800 &  x803 &  x809 &  x812 &  x815 &  x818 &  x820 &  x824 &  x827 &  x830 &  x833 &  x836 &  x848 &  x851 &  x857 &  x860 &  x866 &  x869 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x892 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x914 &  x920 &  x923 &  x926 &  x932 &  x937 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x976 &  x977 &  x980 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1013 &  x1022 &  x1025 &  x1031 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x234 & ~x273 & ~x312 & ~x351 & ~x390 & ~x573 & ~x825 & ~x981;
assign c2136 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x89 &  x92 &  x95 &  x101 &  x104 &  x107 &  x110 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x278 &  x281 &  x284 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x383 &  x386 &  x389 &  x392 &  x394 &  x395 &  x398 &  x400 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x470 &  x473 &  x476 &  x479 &  x482 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x884 &  x887 &  x890 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x117 & ~x156 & ~x195 & ~x441 & ~x480 & ~x726 & ~x744 & ~x765 & ~x780;
assign c2138 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x44 &  x47 &  x50 &  x53 &  x56 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x86 &  x89 &  x95 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x236 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x283 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x305 &  x308 &  x314 &  x317 &  x320 &  x323 &  x329 &  x335 &  x341 &  x347 &  x350 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x395 &  x401 &  x404 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x752 &  x755 &  x761 &  x764 &  x767 &  x770 &  x776 &  x779 &  x785 &  x791 &  x794 &  x797 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x893 &  x899 &  x902 &  x905 &  x908 &  x911 &  x917 &  x920 &  x923 &  x929 &  x932 &  x938 &  x941 &  x944 &  x947 &  x950 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 & ~x378 & ~x396 & ~x513 & ~x588 & ~x627 & ~x666 & ~x667 & ~x705 & ~x744 & ~x783 & ~x819 & ~x822 & ~x825 & ~x864;
assign c2140 =  x2 &  x8 &  x17 &  x38 &  x44 &  x50 &  x59 &  x65 &  x68 &  x71 &  x74 &  x83 &  x86 &  x104 &  x110 &  x116 &  x119 &  x128 &  x137 &  x140 &  x143 &  x146 &  x152 &  x155 &  x158 &  x161 &  x164 &  x194 &  x197 &  x203 &  x206 &  x212 &  x218 &  x221 &  x224 &  x230 &  x236 &  x242 &  x251 &  x257 &  x272 &  x281 &  x287 &  x296 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x326 &  x329 &  x341 &  x344 &  x350 &  x353 &  x356 &  x359 &  x371 &  x374 &  x377 &  x380 &  x386 &  x392 &  x395 &  x401 &  x410 &  x422 &  x428 &  x437 &  x440 &  x443 &  x446 &  x449 &  x455 &  x458 &  x461 &  x467 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x506 &  x509 &  x512 &  x521 &  x527 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x563 &  x572 &  x575 &  x581 &  x584 &  x596 &  x599 &  x605 &  x608 &  x614 &  x620 &  x629 &  x632 &  x635 &  x638 &  x647 &  x653 &  x659 &  x662 &  x665 &  x668 &  x671 &  x692 &  x695 &  x701 &  x704 &  x707 &  x713 &  x716 &  x725 &  x728 &  x734 &  x737 &  x743 &  x749 &  x758 &  x761 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x797 &  x803 &  x806 &  x815 &  x824 &  x827 &  x839 &  x842 &  x854 &  x887 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x926 &  x929 &  x944 &  x953 &  x965 &  x971 &  x974 &  x977 &  x980 &  x983 &  x1001 &  x1004 &  x1010 &  x1013 &  x1022 &  x1025 &  x1037 &  x1040 &  x1043 &  x1049 &  x1064 &  x1070 &  x1073 &  x1082 &  x1085 &  x1091 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1127 & ~x99 & ~x456 & ~x669 & ~x702 & ~x843 & ~x879 & ~x880 & ~x885;
assign c2142 =  x8 &  x14 &  x17 &  x20 &  x23 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x74 &  x77 &  x86 &  x89 &  x95 &  x98 &  x101 &  x107 &  x110 &  x113 &  x116 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x155 &  x173 &  x176 &  x182 &  x185 &  x188 &  x194 &  x197 &  x206 &  x209 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x251 &  x254 &  x260 &  x263 &  x266 &  x275 &  x277 &  x281 &  x284 &  x287 &  x293 &  x296 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x332 &  x338 &  x347 &  x350 &  x353 &  x356 &  x359 &  x368 &  x371 &  x374 &  x377 &  x389 &  x392 &  x395 &  x401 &  x416 &  x419 &  x422 &  x428 &  x430 &  x434 &  x437 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x469 &  x470 &  x473 &  x476 &  x479 &  x482 &  x488 &  x497 &  x500 &  x506 &  x508 &  x509 &  x512 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x539 &  x545 &  x548 &  x554 &  x557 &  x560 &  x563 &  x566 &  x575 &  x578 &  x581 &  x587 &  x593 &  x596 &  x599 &  x605 &  x617 &  x620 &  x623 &  x629 &  x632 &  x638 &  x641 &  x647 &  x659 &  x662 &  x665 &  x671 &  x677 &  x680 &  x683 &  x686 &  x704 &  x707 &  x713 &  x716 &  x719 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x770 &  x773 &  x776 &  x785 &  x791 &  x794 &  x800 &  x803 &  x809 &  x812 &  x818 &  x824 &  x827 &  x830 &  x833 &  x845 &  x848 &  x851 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x884 &  x890 &  x893 &  x896 &  x902 &  x905 &  x908 &  x911 &  x917 &  x920 &  x926 &  x929 &  x932 &  x935 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x971 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1067 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x402 & ~x441 & ~x474 & ~x480 & ~x519 & ~x525 & ~x552 & ~x591 & ~x681 & ~x708 & ~x720 & ~x753 & ~x759;
assign c2144 =  x2 &  x5 &  x8 &  x17 &  x20 &  x23 &  x38 &  x41 &  x44 &  x50 &  x53 &  x56 &  x59 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x92 &  x101 &  x104 &  x107 &  x119 &  x125 &  x131 &  x140 &  x146 &  x149 &  x152 &  x155 &  x161 &  x167 &  x176 &  x179 &  x182 &  x185 &  x191 &  x194 &  x203 &  x206 &  x209 &  x212 &  x221 &  x227 &  x230 &  x232 &  x239 &  x242 &  x245 &  x257 &  x260 &  x263 &  x269 &  x272 &  x278 &  x284 &  x290 &  x302 &  x314 &  x317 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x353 &  x359 &  x362 &  x368 &  x374 &  x377 &  x380 &  x389 &  x392 &  x395 &  x401 &  x404 &  x407 &  x413 &  x419 &  x422 &  x425 &  x428 &  x434 &  x437 &  x449 &  x452 &  x458 &  x461 &  x470 &  x479 &  x482 &  x488 &  x491 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x581 &  x587 &  x593 &  x596 &  x602 &  x605 &  x611 &  x614 &  x623 &  x632 &  x644 &  x650 &  x659 &  x665 &  x674 &  x680 &  x686 &  x692 &  x695 &  x698 &  x716 &  x722 &  x725 &  x728 &  x734 &  x737 &  x743 &  x746 &  x755 &  x758 &  x764 &  x767 &  x770 &  x773 &  x776 &  x782 &  x791 &  x800 &  x803 &  x806 &  x812 &  x815 &  x818 &  x827 &  x830 &  x836 &  x839 &  x845 &  x851 &  x860 &  x869 &  x872 &  x875 &  x878 &  x887 &  x893 &  x896 &  x899 &  x902 &  x908 &  x917 &  x920 &  x929 &  x935 &  x941 &  x944 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x980 &  x983 &  x985 &  x986 &  x989 &  x998 &  x1001 &  x1004 &  x1016 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1049 &  x1055 &  x1064 &  x1067 &  x1070 &  x1088 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1130 & ~x402 & ~x441 & ~x861 & ~x900 & ~x939 & ~x1017 & ~x1038 & ~x1050;
assign c2146 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x29 &  x35 &  x41 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x80 &  x83 &  x89 &  x92 &  x98 &  x104 &  x107 &  x110 &  x113 &  x119 &  x122 &  x125 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x181 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x209 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x284 &  x290 &  x293 &  x299 &  x305 &  x311 &  x314 &  x320 &  x323 &  x326 &  x329 &  x338 &  x341 &  x347 &  x350 &  x353 &  x356 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x419 &  x422 &  x425 &  x431 &  x437 &  x440 &  x446 &  x449 &  x452 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x497 &  x500 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x590 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x686 &  x692 &  x695 &  x698 &  x701 &  x704 &  x710 &  x713 &  x716 &  x719 &  x722 &  x728 &  x731 &  x734 &  x737 &  x743 &  x746 &  x749 &  x755 &  x764 &  x767 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x794 &  x797 &  x800 &  x803 &  x806 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x839 &  x842 &  x845 &  x848 &  x854 &  x857 &  x860 &  x866 &  x869 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x908 &  x911 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x992 &  x1001 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x234 & ~x402 & ~x441 & ~x480 & ~x636 & ~x666 & ~x831 & ~x861 & ~x900 & ~x939 & ~x948;
assign c2148 =  x2 &  x5 &  x11 &  x14 &  x20 &  x23 &  x26 &  x32 &  x35 &  x41 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x98 &  x107 &  x110 &  x116 &  x119 &  x122 &  x125 &  x128 &  x134 &  x140 &  x146 &  x152 &  x155 &  x158 &  x161 &  x164 &  x173 &  x179 &  x185 &  x188 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x218 &  x221 &  x224 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x266 &  x275 &  x278 &  x281 &  x287 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x326 &  x329 &  x335 &  x338 &  x341 &  x344 &  x350 &  x353 &  x355 &  x359 &  x361 &  x362 &  x365 &  x368 &  x371 &  x380 &  x383 &  x386 &  x389 &  x392 &  x400 &  x401 &  x404 &  x407 &  x413 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x452 &  x455 &  x458 &  x461 &  x467 &  x469 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x494 &  x497 &  x500 &  x506 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x542 &  x545 &  x547 &  x548 &  x551 &  x554 &  x557 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x587 &  x590 &  x593 &  x596 &  x599 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x635 &  x638 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x728 &  x731 &  x734 &  x737 &  x740 &  x742 &  x743 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x806 &  x809 &  x812 &  x815 &  x818 &  x824 &  x827 &  x833 &  x836 &  x842 &  x845 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x872 &  x875 &  x881 &  x884 &  x887 &  x893 &  x899 &  x902 &  x905 &  x911 &  x917 &  x920 &  x926 &  x929 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x983 &  x992 &  x1001 &  x1007 &  x1013 &  x1016 &  x1019 &  x1025 &  x1031 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 & ~x342 & ~x381 & ~x441 & ~x480 & ~x783 & ~x822;
assign c2150 =  x2 &  x8 &  x11 &  x17 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x86 &  x89 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x160 &  x161 &  x167 &  x170 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x197 &  x199 &  x200 &  x206 &  x209 &  x212 &  x218 &  x221 &  x224 &  x227 &  x236 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x274 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x302 &  x305 &  x311 &  x313 &  x314 &  x317 &  x326 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x365 &  x368 &  x374 &  x377 &  x380 &  x383 &  x386 &  x392 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x464 &  x467 &  x470 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x524 &  x527 &  x530 &  x533 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x587 &  x590 &  x596 &  x599 &  x602 &  x605 &  x608 &  x620 &  x626 &  x629 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x665 &  x668 &  x671 &  x674 &  x677 &  x683 &  x695 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x788 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x851 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x893 &  x896 &  x899 &  x905 &  x908 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x947 &  x950 &  x953 &  x956 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 & ~x54 & ~x55 & ~x93 & ~x396 & ~x435 & ~x585 & ~x624 & ~x627 & ~x663 & ~x702 & ~x741 & ~x780 & ~x1062;
assign c2152 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x310 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x349 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x99 & ~x339 & ~x495 & ~x534 & ~x573 & ~x612 & ~x651 & ~x652 & ~x690 & ~x691 & ~x729 & ~x768 & ~x807 & ~x846 & ~x885 & ~x1002 & ~x1119;
assign c2154 =  x5 &  x11 &  x14 &  x17 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x59 &  x62 &  x68 &  x71 &  x83 &  x92 &  x98 &  x101 &  x107 &  x110 &  x113 &  x116 &  x119 &  x121 &  x122 &  x125 &  x127 &  x128 &  x134 &  x140 &  x152 &  x158 &  x161 &  x167 &  x173 &  x191 &  x200 &  x203 &  x206 &  x209 &  x212 &  x218 &  x221 &  x227 &  x230 &  x233 &  x235 &  x236 &  x242 &  x248 &  x251 &  x257 &  x260 &  x263 &  x266 &  x275 &  x278 &  x281 &  x284 &  x287 &  x293 &  x296 &  x302 &  x308 &  x311 &  x313 &  x314 &  x320 &  x323 &  x329 &  x341 &  x344 &  x350 &  x353 &  x356 &  x365 &  x374 &  x389 &  x392 &  x398 &  x407 &  x410 &  x413 &  x419 &  x422 &  x424 &  x437 &  x440 &  x443 &  x446 &  x455 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x485 &  x491 &  x494 &  x497 &  x500 &  x503 &  x512 &  x521 &  x539 &  x542 &  x545 &  x560 &  x569 &  x572 &  x575 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x620 &  x623 &  x635 &  x647 &  x650 &  x656 &  x665 &  x668 &  x671 &  x674 &  x680 &  x683 &  x686 &  x692 &  x698 &  x710 &  x722 &  x725 &  x731 &  x740 &  x743 &  x755 &  x758 &  x770 &  x773 &  x776 &  x779 &  x782 &  x791 &  x797 &  x800 &  x806 &  x812 &  x815 &  x818 &  x821 &  x830 &  x833 &  x836 &  x839 &  x842 &  x851 &  x854 &  x860 &  x863 &  x866 &  x869 &  x871 &  x872 &  x875 &  x878 &  x887 &  x896 &  x902 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x959 &  x962 &  x977 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1061 &  x1067 &  x1076 &  x1079 &  x1100 &  x1103 &  x1106 &  x1118 &  x1121 &  x1124 & ~x279 & ~x510 & ~x552 & ~x627 & ~x744 & ~x975 & ~x1014;
assign c2156 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x44 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x134 &  x137 &  x143 &  x146 &  x149 &  x152 &  x155 &  x161 &  x167 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x218 &  x224 &  x227 &  x230 &  x236 &  x239 &  x245 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x317 &  x320 &  x326 &  x329 &  x332 &  x335 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x425 &  x431 &  x434 &  x437 &  x440 &  x443 &  x449 &  x452 &  x455 &  x458 &  x461 &  x470 &  x473 &  x476 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x626 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x668 &  x671 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x703 &  x707 &  x710 &  x716 &  x719 &  x725 &  x731 &  x734 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x806 &  x809 &  x812 &  x815 &  x818 &  x824 &  x827 &  x833 &  x836 &  x839 &  x842 &  x845 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1046 &  x1049 &  x1055 &  x1058 &  x1061 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 & ~x126 & ~x165 & ~x195 & ~x234 & ~x273 & ~x558 & ~x597 & ~x636 & ~x669 & ~x675 & ~x714 & ~x747 & ~x753 & ~x786 & ~x792 & ~x939 & ~x978 & ~x1017;
assign c2158 =  x2 &  x5 &  x8 &  x11 &  x17 &  x20 &  x29 &  x32 &  x38 &  x41 &  x44 &  x50 &  x56 &  x59 &  x65 &  x71 &  x74 &  x77 &  x86 &  x89 &  x92 &  x98 &  x107 &  x110 &  x116 &  x119 &  x122 &  x125 &  x134 &  x137 &  x140 &  x146 &  x149 &  x155 &  x158 &  x161 &  x164 &  x167 &  x176 &  x188 &  x191 &  x194 &  x203 &  x206 &  x212 &  x221 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x257 &  x260 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x302 &  x305 &  x308 &  x311 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x368 &  x370 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x395 &  x398 &  x401 &  x404 &  x407 &  x413 &  x422 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x452 &  x455 &  x461 &  x467 &  x473 &  x476 &  x479 &  x482 &  x491 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x527 &  x533 &  x539 &  x551 &  x554 &  x563 &  x566 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x598 &  x599 &  x602 &  x605 &  x611 &  x623 &  x626 &  x635 &  x638 &  x641 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x667 &  x671 &  x674 &  x677 &  x680 &  x686 &  x692 &  x695 &  x698 &  x707 &  x713 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x761 &  x764 &  x767 &  x770 &  x773 &  x779 &  x782 &  x785 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x821 &  x839 &  x842 &  x845 &  x851 &  x854 &  x857 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x941 &  x944 &  x947 &  x950 &  x953 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x989 &  x992 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1061 &  x1070 &  x1073 &  x1079 &  x1088 &  x1091 &  x1094 &  x1100 &  x1106 &  x1109 &  x1112 &  x1118 &  x1124 &  x1127 &  x1130 & ~x810 & ~x882 & ~x921 & ~x981 & ~x1038 & ~x1116;
assign c2160 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x46 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x85 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x124 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x316 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x355 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x718 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x757 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x796 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x835 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x874 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x516 & ~x687 & ~x702 & ~x726 & ~x744 & ~x783;
assign c2162 =  x8 &  x11 &  x14 &  x20 &  x23 &  x32 &  x38 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x71 &  x77 &  x80 &  x86 &  x98 &  x101 &  x107 &  x110 &  x116 &  x122 &  x125 &  x128 &  x134 &  x137 &  x140 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x170 &  x176 &  x185 &  x188 &  x191 &  x197 &  x203 &  x206 &  x209 &  x215 &  x218 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x266 &  x269 &  x275 &  x278 &  x281 &  x290 &  x293 &  x296 &  x299 &  x305 &  x311 &  x317 &  x320 &  x323 &  x338 &  x341 &  x350 &  x353 &  x362 &  x380 &  x386 &  x389 &  x392 &  x401 &  x410 &  x413 &  x431 &  x434 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x467 &  x470 &  x473 &  x476 &  x485 &  x491 &  x503 &  x509 &  x512 &  x524 &  x527 &  x530 &  x533 &  x539 &  x542 &  x551 &  x554 &  x557 &  x563 &  x566 &  x575 &  x578 &  x581 &  x584 &  x587 &  x596 &  x599 &  x602 &  x608 &  x611 &  x626 &  x632 &  x638 &  x641 &  x644 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x668 &  x677 &  x680 &  x683 &  x689 &  x692 &  x698 &  x703 &  x719 &  x722 &  x728 &  x731 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x770 &  x773 &  x779 &  x782 &  x788 &  x794 &  x800 &  x803 &  x806 &  x812 &  x815 &  x818 &  x821 &  x833 &  x836 &  x839 &  x842 &  x848 &  x854 &  x857 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x890 &  x896 &  x899 &  x920 &  x926 &  x941 &  x947 &  x953 &  x965 &  x974 &  x980 &  x983 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1013 &  x1016 &  x1022 &  x1025 &  x1031 &  x1043 &  x1046 &  x1049 &  x1058 &  x1070 &  x1076 &  x1082 &  x1085 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1121 &  x1124 &  x1127 & ~x558 & ~x636 & ~x669 & ~x676 & ~x714 & ~x747 & ~x792 & ~x864 & ~x939 & ~x978;
assign c2164 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x277 &  x278 &  x283 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x316 &  x317 &  x320 &  x322 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x355 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x391 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x430 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x469 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x508 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x547 &  x548 &  x551 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x366 & ~x405 & ~x630 & ~x705 & ~x744 & ~x783 & ~x822 & ~x861 & ~x900;
assign c2166 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x59 &  x62 &  x65 &  x71 &  x74 &  x77 &  x80 &  x83 &  x92 &  x95 &  x98 &  x101 &  x104 &  x113 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x149 &  x152 &  x155 &  x158 &  x161 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x209 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x278 &  x281 &  x284 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x325 &  x326 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x356 &  x359 &  x362 &  x364 &  x365 &  x368 &  x370 &  x371 &  x374 &  x380 &  x389 &  x398 &  x404 &  x407 &  x409 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x455 &  x458 &  x461 &  x470 &  x473 &  x476 &  x479 &  x481 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x518 &  x520 &  x521 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x548 &  x551 &  x563 &  x565 &  x566 &  x569 &  x572 &  x578 &  x581 &  x584 &  x590 &  x602 &  x604 &  x605 &  x608 &  x611 &  x614 &  x617 &  x623 &  x626 &  x632 &  x635 &  x643 &  x644 &  x647 &  x650 &  x656 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x680 &  x681 &  x682 &  x683 &  x686 &  x689 &  x695 &  x701 &  x704 &  x707 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x779 &  x782 &  x785 &  x791 &  x794 &  x797 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x857 &  x860 &  x863 &  x866 &  x872 &  x874 &  x875 &  x881 &  x884 &  x887 &  x890 &  x893 &  x902 &  x908 &  x911 &  x914 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x944 &  x947 &  x950 &  x953 &  x962 &  x965 &  x968 &  x974 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1034 &  x1037 &  x1040 &  x1046 &  x1058 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x144 & ~x183;
assign c2168 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x26 &  x29 &  x32 &  x38 &  x44 &  x47 &  x50 &  x53 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x101 &  x113 &  x116 &  x119 &  x122 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x152 &  x161 &  x164 &  x167 &  x170 &  x173 &  x182 &  x185 &  x188 &  x191 &  x197 &  x203 &  x206 &  x212 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x242 &  x251 &  x260 &  x269 &  x275 &  x284 &  x290 &  x296 &  x302 &  x305 &  x314 &  x320 &  x323 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x368 &  x371 &  x374 &  x377 &  x383 &  x386 &  x389 &  x398 &  x401 &  x404 &  x407 &  x410 &  x416 &  x422 &  x425 &  x428 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x464 &  x467 &  x472 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x497 &  x500 &  x503 &  x509 &  x511 &  x512 &  x521 &  x524 &  x530 &  x533 &  x542 &  x545 &  x547 &  x551 &  x560 &  x569 &  x572 &  x581 &  x586 &  x590 &  x593 &  x596 &  x599 &  x602 &  x608 &  x611 &  x617 &  x620 &  x623 &  x625 &  x626 &  x632 &  x638 &  x643 &  x644 &  x650 &  x653 &  x656 &  x659 &  x665 &  x668 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x707 &  x713 &  x724 &  x725 &  x731 &  x737 &  x749 &  x758 &  x761 &  x763 &  x764 &  x773 &  x776 &  x782 &  x788 &  x791 &  x797 &  x799 &  x800 &  x802 &  x803 &  x806 &  x809 &  x812 &  x821 &  x827 &  x830 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x896 &  x899 &  x905 &  x911 &  x932 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x989 &  x992 &  x995 &  x998 &  x1007 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1028 &  x1034 &  x1037 &  x1040 &  x1043 &  x1055 &  x1058 &  x1067 &  x1073 &  x1079 &  x1085 &  x1112 &  x1121 &  x1124 &  x1127 & ~x459 & ~x498 & ~x849;
assign c2170 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x26 &  x44 &  x47 &  x50 &  x53 &  x56 &  x62 &  x65 &  x68 &  x71 &  x77 &  x80 &  x83 &  x86 &  x89 &  x98 &  x104 &  x113 &  x116 &  x119 &  x125 &  x128 &  x131 &  x134 &  x137 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x173 &  x179 &  x182 &  x191 &  x194 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x233 &  x248 &  x260 &  x269 &  x278 &  x281 &  x284 &  x290 &  x302 &  x305 &  x308 &  x317 &  x320 &  x323 &  x326 &  x332 &  x335 &  x347 &  x353 &  x356 &  x362 &  x368 &  x377 &  x383 &  x386 &  x389 &  x395 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x431 &  x434 &  x440 &  x446 &  x449 &  x464 &  x473 &  x479 &  x482 &  x485 &  x488 &  x491 &  x497 &  x506 &  x509 &  x512 &  x515 &  x518 &  x524 &  x527 &  x533 &  x536 &  x539 &  x542 &  x545 &  x551 &  x554 &  x557 &  x563 &  x566 &  x569 &  x578 &  x587 &  x590 &  x593 &  x596 &  x602 &  x608 &  x623 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x656 &  x662 &  x677 &  x680 &  x692 &  x695 &  x698 &  x704 &  x710 &  x713 &  x719 &  x731 &  x740 &  x743 &  x746 &  x749 &  x752 &  x758 &  x776 &  x785 &  x788 &  x791 &  x806 &  x809 &  x812 &  x818 &  x821 &  x824 &  x827 &  x833 &  x845 &  x848 &  x851 &  x854 &  x860 &  x863 &  x866 &  x869 &  x878 &  x881 &  x893 &  x896 &  x899 &  x920 &  x926 &  x932 &  x935 &  x941 &  x944 &  x950 &  x956 &  x968 &  x971 &  x980 &  x983 &  x986 &  x992 &  x1001 &  x1004 &  x1007 &  x1010 &  x1019 &  x1022 &  x1025 &  x1037 &  x1040 &  x1043 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1091 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 & ~x570 & ~x675 & ~x687 & ~x714 & ~x727 & ~x747 & ~x753 & ~x765 & ~x786 & ~x831 & ~x978 & ~x999 & ~x1038;
assign c2172 =  x2 &  x14 &  x23 &  x32 &  x41 &  x44 &  x47 &  x50 &  x56 &  x59 &  x80 &  x92 &  x98 &  x101 &  x107 &  x113 &  x116 &  x131 &  x134 &  x146 &  x149 &  x164 &  x170 &  x173 &  x182 &  x185 &  x191 &  x194 &  x197 &  x206 &  x209 &  x218 &  x224 &  x233 &  x236 &  x239 &  x245 &  x251 &  x254 &  x263 &  x266 &  x272 &  x278 &  x281 &  x284 &  x287 &  x293 &  x296 &  x314 &  x326 &  x329 &  x332 &  x335 &  x341 &  x374 &  x377 &  x389 &  x407 &  x419 &  x422 &  x437 &  x440 &  x443 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x476 &  x487 &  x494 &  x509 &  x515 &  x521 &  x524 &  x530 &  x533 &  x539 &  x548 &  x554 &  x560 &  x565 &  x569 &  x575 &  x578 &  x587 &  x590 &  x599 &  x602 &  x629 &  x632 &  x635 &  x640 &  x662 &  x671 &  x679 &  x680 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x707 &  x710 &  x718 &  x722 &  x728 &  x740 &  x746 &  x752 &  x756 &  x757 &  x758 &  x761 &  x770 &  x773 &  x776 &  x794 &  x796 &  x800 &  x803 &  x806 &  x809 &  x815 &  x827 &  x833 &  x835 &  x836 &  x839 &  x845 &  x848 &  x851 &  x854 &  x863 &  x874 &  x875 &  x878 &  x887 &  x890 &  x905 &  x908 &  x911 &  x932 &  x938 &  x941 &  x950 &  x953 &  x956 &  x974 &  x989 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1013 &  x1025 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1082 &  x1085 &  x1088 &  x1097 &  x1100 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 & ~x510 & ~x549 & ~x552 & ~x589 & ~x627 & ~x666 & ~x705;
assign c2174 =  x2 &  x5 &  x8 &  x20 &  x26 &  x29 &  x35 &  x47 &  x56 &  x59 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x104 &  x107 &  x110 &  x122 &  x131 &  x134 &  x135 &  x137 &  x140 &  x146 &  x149 &  x152 &  x155 &  x170 &  x176 &  x182 &  x185 &  x188 &  x191 &  x197 &  x203 &  x206 &  x209 &  x218 &  x230 &  x236 &  x239 &  x242 &  x251 &  x254 &  x257 &  x260 &  x269 &  x272 &  x275 &  x278 &  x290 &  x296 &  x302 &  x305 &  x311 &  x314 &  x320 &  x329 &  x332 &  x335 &  x341 &  x344 &  x347 &  x350 &  x356 &  x365 &  x368 &  x386 &  x392 &  x398 &  x404 &  x407 &  x409 &  x410 &  x416 &  x419 &  x424 &  x425 &  x428 &  x431 &  x434 &  x443 &  x449 &  x458 &  x464 &  x470 &  x473 &  x476 &  x479 &  x482 &  x487 &  x503 &  x512 &  x515 &  x521 &  x536 &  x539 &  x548 &  x560 &  x572 &  x578 &  x584 &  x587 &  x596 &  x599 &  x602 &  x617 &  x623 &  x626 &  x629 &  x632 &  x638 &  x644 &  x647 &  x653 &  x671 &  x680 &  x692 &  x695 &  x701 &  x704 &  x713 &  x716 &  x722 &  x725 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x761 &  x764 &  x779 &  x782 &  x797 &  x799 &  x809 &  x815 &  x821 &  x830 &  x838 &  x839 &  x842 &  x848 &  x854 &  x863 &  x866 &  x869 &  x890 &  x893 &  x896 &  x905 &  x908 &  x911 &  x920 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x953 &  x956 &  x959 &  x962 &  x965 &  x974 &  x977 &  x980 &  x989 &  x995 &  x1004 &  x1010 &  x1019 &  x1028 &  x1037 &  x1040 &  x1052 &  x1058 &  x1061 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1112 &  x1115 &  x1121 & ~x378 & ~x702 & ~x819;
assign c2176 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x397 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x434 &  x436 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x117 & ~x156 & ~x195 & ~x339 & ~x417 & ~x456 & ~x792 & ~x831 & ~x882 & ~x921 & ~x1056 & ~x1095;
assign c2178 =  x5 &  x8 &  x11 &  x14 &  x17 &  x32 &  x44 &  x62 &  x68 &  x71 &  x77 &  x80 &  x83 &  x86 &  x89 &  x101 &  x104 &  x107 &  x113 &  x131 &  x137 &  x140 &  x143 &  x149 &  x152 &  x155 &  x158 &  x164 &  x170 &  x173 &  x176 &  x179 &  x185 &  x197 &  x200 &  x203 &  x206 &  x215 &  x221 &  x224 &  x233 &  x245 &  x251 &  x254 &  x257 &  x260 &  x278 &  x287 &  x290 &  x293 &  x305 &  x308 &  x311 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x350 &  x359 &  x362 &  x368 &  x370 &  x377 &  x383 &  x398 &  x406 &  x410 &  x425 &  x427 &  x428 &  x440 &  x443 &  x446 &  x447 &  x449 &  x455 &  x470 &  x479 &  x482 &  x485 &  x494 &  x500 &  x503 &  x515 &  x521 &  x523 &  x524 &  x526 &  x530 &  x536 &  x539 &  x542 &  x554 &  x563 &  x566 &  x569 &  x575 &  x581 &  x596 &  x605 &  x620 &  x629 &  x640 &  x641 &  x644 &  x653 &  x656 &  x662 &  x668 &  x677 &  x679 &  x680 &  x689 &  x698 &  x701 &  x712 &  x713 &  x716 &  x731 &  x734 &  x746 &  x749 &  x752 &  x760 &  x761 &  x764 &  x767 &  x797 &  x803 &  x809 &  x812 &  x815 &  x821 &  x827 &  x839 &  x845 &  x854 &  x857 &  x860 &  x863 &  x878 &  x881 &  x887 &  x890 &  x896 &  x908 &  x914 &  x916 &  x920 &  x923 &  x929 &  x932 &  x935 &  x947 &  x959 &  x965 &  x968 &  x971 &  x983 &  x989 &  x1001 &  x1004 &  x1010 &  x1016 &  x1019 &  x1022 &  x1028 &  x1064 &  x1073 &  x1076 &  x1097 &  x1106 &  x1109 &  x1115 &  x1130;
assign c2180 =  x5 &  x11 &  x23 &  x26 &  x50 &  x56 &  x77 &  x80 &  x83 &  x95 &  x98 &  x101 &  x143 &  x149 &  x161 &  x167 &  x170 &  x176 &  x188 &  x227 &  x236 &  x257 &  x281 &  x284 &  x296 &  x299 &  x302 &  x305 &  x314 &  x317 &  x332 &  x338 &  x341 &  x344 &  x356 &  x365 &  x380 &  x386 &  x404 &  x407 &  x431 &  x440 &  x470 &  x473 &  x479 &  x482 &  x491 &  x494 &  x503 &  x509 &  x527 &  x530 &  x539 &  x557 &  x566 &  x572 &  x584 &  x592 &  x611 &  x629 &  x632 &  x635 &  x647 &  x653 &  x656 &  x668 &  x674 &  x677 &  x680 &  x689 &  x706 &  x713 &  x719 &  x728 &  x737 &  x749 &  x776 &  x797 &  x803 &  x827 &  x833 &  x848 &  x851 &  x860 &  x869 &  x872 &  x878 &  x881 &  x893 &  x896 &  x908 &  x920 &  x929 &  x944 &  x953 &  x1004 &  x1016 &  x1031 &  x1034 &  x1067 &  x1070 &  x1079 &  x1085 &  x1088 &  x1094 &  x1103 &  x1121 &  x1127 &  x1130 & ~x123 & ~x162 & ~x240 & ~x351 & ~x717 & ~x729 & ~x1020;
assign c2182 =  x5 &  x11 &  x20 &  x26 &  x29 &  x44 &  x47 &  x50 &  x59 &  x77 &  x83 &  x95 &  x98 &  x104 &  x107 &  x113 &  x119 &  x122 &  x134 &  x137 &  x146 &  x152 &  x158 &  x164 &  x170 &  x185 &  x191 &  x197 &  x206 &  x209 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x269 &  x287 &  x290 &  x299 &  x314 &  x320 &  x329 &  x332 &  x335 &  x338 &  x344 &  x347 &  x353 &  x362 &  x368 &  x374 &  x377 &  x380 &  x383 &  x389 &  x392 &  x395 &  x404 &  x410 &  x412 &  x437 &  x446 &  x452 &  x461 &  x473 &  x489 &  x490 &  x494 &  x503 &  x512 &  x524 &  x527 &  x529 &  x530 &  x533 &  x545 &  x575 &  x581 &  x586 &  x593 &  x602 &  x607 &  x617 &  x620 &  x623 &  x625 &  x629 &  x638 &  x662 &  x665 &  x671 &  x686 &  x692 &  x701 &  x707 &  x713 &  x719 &  x746 &  x755 &  x758 &  x776 &  x781 &  x782 &  x785 &  x788 &  x806 &  x820 &  x824 &  x827 &  x839 &  x841 &  x845 &  x859 &  x863 &  x866 &  x878 &  x884 &  x896 &  x898 &  x902 &  x914 &  x917 &  x920 &  x935 &  x937 &  x938 &  x944 &  x983 &  x989 &  x998 &  x1007 &  x1010 &  x1013 &  x1022 &  x1025 &  x1028 &  x1040 &  x1043 &  x1052 &  x1061 &  x1070 &  x1079 &  x1088 &  x1091 &  x1097 &  x1109 &  x1115 &  x1124 & ~x981 & ~x1026 & ~x1038 & ~x1065;
assign c2184 =  x8 &  x14 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x80 &  x83 &  x92 &  x98 &  x101 &  x104 &  x107 &  x119 &  x121 &  x122 &  x125 &  x131 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x161 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x194 &  x196 &  x197 &  x200 &  x212 &  x218 &  x221 &  x224 &  x227 &  x230 &  x235 &  x236 &  x242 &  x245 &  x248 &  x254 &  x257 &  x260 &  x266 &  x269 &  x272 &  x274 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x296 &  x299 &  x302 &  x308 &  x311 &  x313 &  x314 &  x317 &  x323 &  x329 &  x332 &  x344 &  x350 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x401 &  x404 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x458 &  x464 &  x467 &  x470 &  x479 &  x482 &  x491 &  x500 &  x503 &  x509 &  x512 &  x515 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x545 &  x548 &  x554 &  x557 &  x560 &  x566 &  x569 &  x575 &  x578 &  x581 &  x584 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x698 &  x704 &  x713 &  x716 &  x718 &  x719 &  x722 &  x728 &  x731 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x757 &  x758 &  x761 &  x764 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x809 &  x815 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x842 &  x848 &  x851 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x932 &  x938 &  x941 &  x944 &  x950 &  x959 &  x962 &  x965 &  x968 &  x971 &  x980 &  x983 &  x986 &  x988 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1066 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1100 &  x1103 &  x1106 &  x1109 &  x1111 &  x1112 &  x1118 &  x1124 &  x1127 &  x1130 & ~x318 & ~x357 & ~x396 & ~x435 & ~x438 & ~x474 & ~x513 & ~x627 & ~x666 & ~x705;
assign c2186 =  x2 &  x5 &  x8 &  x11 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x140 &  x143 &  x146 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x290 &  x293 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x356 &  x359 &  x362 &  x364 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x458 &  x461 &  x464 &  x470 &  x473 &  x475 &  x476 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x628 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x659 &  x662 &  x664 &  x667 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x698 &  x701 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x742 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x781 &  x782 &  x785 &  x788 &  x791 &  x794 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x820 &  x821 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x896 &  x898 &  x899 &  x902 &  x905 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x937 &  x944 &  x947 &  x950 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x976 &  x977 &  x983 &  x986 &  x989 &  x992 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1093 &  x1094 &  x1097 &  x1100 &  x1103 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x234 & ~x273 & ~x312 & ~x351 & ~x390 & ~x429 & ~x942 & ~x978 & ~x1017;
assign c2188 =  x2 &  x8 &  x11 &  x23 &  x32 &  x35 &  x41 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x122 &  x131 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x167 &  x179 &  x182 &  x185 &  x188 &  x194 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x257 &  x260 &  x263 &  x275 &  x284 &  x287 &  x293 &  x302 &  x308 &  x311 &  x314 &  x317 &  x319 &  x320 &  x329 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x380 &  x386 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x436 &  x437 &  x440 &  x446 &  x449 &  x458 &  x461 &  x464 &  x467 &  x470 &  x475 &  x485 &  x491 &  x494 &  x497 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x539 &  x548 &  x551 &  x554 &  x560 &  x566 &  x569 &  x572 &  x575 &  x578 &  x590 &  x596 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x626 &  x629 &  x635 &  x638 &  x641 &  x647 &  x656 &  x665 &  x671 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x704 &  x710 &  x713 &  x716 &  x722 &  x725 &  x728 &  x731 &  x737 &  x743 &  x745 &  x749 &  x752 &  x758 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x797 &  x800 &  x803 &  x809 &  x815 &  x818 &  x824 &  x827 &  x836 &  x839 &  x842 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x914 &  x923 &  x926 &  x938 &  x941 &  x947 &  x959 &  x965 &  x968 &  x971 &  x974 &  x976 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1016 &  x1025 &  x1028 &  x1046 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1082 &  x1085 &  x1088 &  x1093 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x234 & ~x273 & ~x312 & ~x351 & ~x390 & ~x429 & ~x507 & ~x807 & ~x906 & ~x1020 & ~x1038 & ~x1059 & ~x1098;
assign c2190 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x83 &  x86 &  x89 &  x92 &  x95 &  x104 &  x107 &  x110 &  x113 &  x119 &  x122 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x161 &  x167 &  x170 &  x173 &  x176 &  x179 &  x188 &  x194 &  x197 &  x202 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x266 &  x269 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x320 &  x323 &  x329 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x365 &  x368 &  x371 &  x374 &  x386 &  x392 &  x395 &  x398 &  x404 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x434 &  x437 &  x440 &  x446 &  x449 &  x452 &  x455 &  x458 &  x464 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x509 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x560 &  x563 &  x566 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x599 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x629 &  x632 &  x644 &  x647 &  x653 &  x656 &  x659 &  x668 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x704 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x830 &  x833 &  x836 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x935 &  x938 &  x941 &  x944 &  x947 &  x953 &  x956 &  x962 &  x965 &  x971 &  x974 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1049 &  x1052 &  x1055 &  x1058 &  x1067 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1124 &  x1127 &  x1130 & ~x117 & ~x156 & ~x726 & ~x867 & ~x942 & ~x943 & ~x981 & ~x1038 & ~x1059;
assign c2192 =  x5 &  x17 &  x20 &  x26 &  x38 &  x68 &  x77 &  x83 &  x89 &  x98 &  x101 &  x116 &  x128 &  x131 &  x137 &  x143 &  x152 &  x167 &  x176 &  x188 &  x191 &  x200 &  x203 &  x206 &  x209 &  x212 &  x221 &  x224 &  x230 &  x233 &  x239 &  x242 &  x245 &  x248 &  x257 &  x272 &  x290 &  x293 &  x296 &  x299 &  x305 &  x308 &  x311 &  x314 &  x329 &  x332 &  x335 &  x344 &  x352 &  x356 &  x365 &  x368 &  x371 &  x377 &  x380 &  x385 &  x392 &  x395 &  x413 &  x416 &  x423 &  x424 &  x425 &  x431 &  x434 &  x443 &  x449 &  x452 &  x455 &  x458 &  x463 &  x467 &  x479 &  x485 &  x491 &  x494 &  x497 &  x500 &  x502 &  x503 &  x512 &  x521 &  x524 &  x527 &  x530 &  x542 &  x551 &  x557 &  x575 &  x584 &  x590 &  x596 &  x608 &  x617 &  x641 &  x650 &  x653 &  x662 &  x665 &  x674 &  x692 &  x701 &  x710 &  x713 &  x728 &  x737 &  x740 &  x743 &  x749 &  x758 &  x764 &  x767 &  x770 &  x782 &  x791 &  x794 &  x797 &  x800 &  x806 &  x809 &  x818 &  x827 &  x830 &  x833 &  x845 &  x848 &  x851 &  x857 &  x860 &  x866 &  x869 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x905 &  x929 &  x938 &  x947 &  x950 &  x953 &  x959 &  x965 &  x974 &  x977 &  x989 &  x995 &  x998 &  x1007 &  x1019 &  x1022 &  x1034 &  x1049 &  x1052 &  x1061 &  x1064 &  x1070 &  x1076 &  x1079 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 & ~x435 & ~x663 & ~x702 & ~x705 & ~x706 & ~x744;
assign c2194 =  x2 &  x5 &  x8 &  x11 &  x17 &  x20 &  x26 &  x32 &  x47 &  x50 &  x65 &  x71 &  x77 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x155 &  x167 &  x179 &  x185 &  x209 &  x215 &  x221 &  x230 &  x233 &  x236 &  x242 &  x245 &  x254 &  x257 &  x263 &  x266 &  x269 &  x275 &  x293 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x320 &  x323 &  x325 &  x329 &  x332 &  x341 &  x347 &  x350 &  x353 &  x356 &  x359 &  x365 &  x371 &  x392 &  x395 &  x404 &  x407 &  x410 &  x412 &  x419 &  x422 &  x425 &  x428 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x464 &  x476 &  x485 &  x491 &  x497 &  x500 &  x503 &  x506 &  x518 &  x521 &  x530 &  x536 &  x542 &  x548 &  x551 &  x557 &  x560 &  x566 &  x575 &  x578 &  x584 &  x587 &  x589 &  x593 &  x596 &  x599 &  x602 &  x608 &  x611 &  x620 &  x623 &  x629 &  x632 &  x635 &  x638 &  x641 &  x647 &  x650 &  x656 &  x659 &  x662 &  x674 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x710 &  x716 &  x725 &  x731 &  x734 &  x740 &  x746 &  x749 &  x752 &  x758 &  x764 &  x767 &  x770 &  x773 &  x776 &  x785 &  x791 &  x800 &  x809 &  x815 &  x824 &  x842 &  x845 &  x848 &  x851 &  x857 &  x860 &  x863 &  x869 &  x872 &  x875 &  x893 &  x896 &  x905 &  x908 &  x914 &  x917 &  x920 &  x929 &  x941 &  x947 &  x950 &  x953 &  x962 &  x965 &  x968 &  x971 &  x977 &  x980 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1037 &  x1040 &  x1048 &  x1049 &  x1055 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1088 &  x1093 &  x1094 &  x1097 &  x1100 &  x1109 &  x1115 &  x1121 &  x1127 &  x1130 & ~x18 & ~x882 & ~x921 & ~x1000 & ~x1038 & ~x1039 & ~x1116;
assign c2196 =  x11 &  x17 &  x26 &  x38 &  x44 &  x50 &  x56 &  x59 &  x62 &  x65 &  x74 &  x83 &  x86 &  x89 &  x98 &  x110 &  x113 &  x122 &  x125 &  x134 &  x137 &  x140 &  x143 &  x148 &  x161 &  x170 &  x173 &  x179 &  x182 &  x185 &  x187 &  x200 &  x203 &  x221 &  x227 &  x233 &  x236 &  x239 &  x251 &  x254 &  x257 &  x263 &  x266 &  x272 &  x275 &  x284 &  x287 &  x290 &  x293 &  x296 &  x314 &  x323 &  x332 &  x338 &  x341 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x374 &  x380 &  x386 &  x389 &  x398 &  x401 &  x413 &  x416 &  x425 &  x431 &  x434 &  x437 &  x446 &  x455 &  x458 &  x467 &  x470 &  x479 &  x485 &  x488 &  x491 &  x494 &  x497 &  x503 &  x506 &  x509 &  x515 &  x518 &  x524 &  x527 &  x530 &  x536 &  x545 &  x551 &  x554 &  x557 &  x560 &  x578 &  x581 &  x584 &  x587 &  x593 &  x599 &  x605 &  x614 &  x617 &  x620 &  x626 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x683 &  x686 &  x692 &  x695 &  x698 &  x704 &  x719 &  x734 &  x737 &  x746 &  x755 &  x758 &  x761 &  x764 &  x770 &  x776 &  x779 &  x788 &  x791 &  x800 &  x803 &  x806 &  x815 &  x818 &  x827 &  x830 &  x836 &  x839 &  x842 &  x845 &  x863 &  x869 &  x872 &  x878 &  x881 &  x884 &  x887 &  x902 &  x914 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x959 &  x962 &  x965 &  x971 &  x986 &  x1001 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1043 &  x1052 &  x1067 &  x1088 &  x1091 &  x1097 &  x1103 &  x1121 &  x1127 & ~x156 & ~x195 & ~x234 & ~x273 & ~x306 & ~x558 & ~x648 & ~x669 & ~x675 & ~x687 & ~x714 & ~x726 & ~x753 & ~x900 & ~x939;
assign c2198 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x125 &  x131 &  x134 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x181 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x227 &  x230 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x269 &  x272 &  x275 &  x278 &  x281 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x331 &  x332 &  x335 &  x338 &  x341 &  x347 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x409 &  x410 &  x413 &  x416 &  x422 &  x425 &  x431 &  x434 &  x440 &  x443 &  x446 &  x449 &  x455 &  x458 &  x461 &  x464 &  x466 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x491 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x559 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x587 &  x593 &  x596 &  x598 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x637 &  x638 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x722 &  x724 &  x725 &  x728 &  x731 &  x734 &  x737 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x763 &  x764 &  x767 &  x770 &  x773 &  x776 &  x782 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1048 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x885;
assign c2200 =  x2 &  x5 &  x11 &  x23 &  x35 &  x47 &  x50 &  x56 &  x59 &  x62 &  x68 &  x74 &  x89 &  x92 &  x95 &  x98 &  x101 &  x107 &  x110 &  x113 &  x119 &  x121 &  x125 &  x134 &  x137 &  x143 &  x146 &  x152 &  x170 &  x173 &  x185 &  x188 &  x191 &  x197 &  x206 &  x227 &  x230 &  x236 &  x238 &  x239 &  x248 &  x260 &  x263 &  x277 &  x281 &  x284 &  x287 &  x290 &  x308 &  x326 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x365 &  x368 &  x377 &  x380 &  x395 &  x407 &  x410 &  x428 &  x431 &  x434 &  x437 &  x443 &  x446 &  x464 &  x476 &  x488 &  x500 &  x503 &  x509 &  x518 &  x521 &  x527 &  x533 &  x536 &  x545 &  x551 &  x554 &  x560 &  x563 &  x566 &  x572 &  x599 &  x605 &  x611 &  x614 &  x638 &  x644 &  x662 &  x674 &  x680 &  x692 &  x695 &  x713 &  x719 &  x728 &  x731 &  x740 &  x743 &  x746 &  x761 &  x764 &  x776 &  x782 &  x797 &  x800 &  x803 &  x806 &  x809 &  x818 &  x824 &  x827 &  x833 &  x839 &  x842 &  x845 &  x857 &  x875 &  x878 &  x881 &  x896 &  x914 &  x920 &  x923 &  x929 &  x938 &  x944 &  x959 &  x962 &  x968 &  x974 &  x986 &  x998 &  x1004 &  x1010 &  x1013 &  x1022 &  x1027 &  x1028 &  x1043 &  x1049 &  x1058 &  x1064 &  x1066 &  x1067 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1109 &  x1112 &  x1121 &  x1130 & ~x144 & ~x183 & ~x184 & ~x222 & ~x378 & ~x432 & ~x510;
assign c2202 =  x8 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x47 &  x50 &  x53 &  x59 &  x62 &  x65 &  x71 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x158 &  x161 &  x164 &  x170 &  x173 &  x176 &  x179 &  x182 &  x188 &  x191 &  x194 &  x197 &  x203 &  x215 &  x218 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x251 &  x254 &  x257 &  x260 &  x269 &  x272 &  x275 &  x278 &  x281 &  x290 &  x296 &  x299 &  x305 &  x308 &  x314 &  x317 &  x323 &  x332 &  x335 &  x338 &  x344 &  x347 &  x350 &  x353 &  x359 &  x365 &  x380 &  x383 &  x389 &  x392 &  x398 &  x401 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x434 &  x440 &  x443 &  x455 &  x458 &  x461 &  x464 &  x467 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x503 &  x506 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x545 &  x554 &  x557 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x599 &  x605 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x647 &  x650 &  x656 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x713 &  x716 &  x719 &  x722 &  x725 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x752 &  x755 &  x761 &  x764 &  x767 &  x770 &  x773 &  x779 &  x785 &  x788 &  x794 &  x797 &  x809 &  x812 &  x818 &  x821 &  x824 &  x842 &  x845 &  x848 &  x851 &  x860 &  x869 &  x872 &  x875 &  x878 &  x881 &  x893 &  x896 &  x899 &  x902 &  x911 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x968 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1100 &  x1103 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130 & ~x192 & ~x480 & ~x531 & ~x636 & ~x648 & ~x669 & ~x675 & ~x687 & ~x708 & ~x714 & ~x831 & ~x861 & ~x900 & ~x939 & ~x954 & ~x993 & ~x1017;
assign c2204 =  x5 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x47 &  x50 &  x56 &  x59 &  x62 &  x65 &  x74 &  x77 &  x80 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x128 &  x131 &  x134 &  x137 &  x149 &  x152 &  x155 &  x158 &  x161 &  x167 &  x170 &  x173 &  x176 &  x182 &  x185 &  x188 &  x191 &  x197 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x263 &  x266 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x305 &  x308 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x383 &  x386 &  x392 &  x395 &  x401 &  x404 &  x410 &  x413 &  x416 &  x419 &  x422 &  x428 &  x431 &  x434 &  x440 &  x443 &  x449 &  x452 &  x458 &  x467 &  x470 &  x473 &  x476 &  x482 &  x485 &  x488 &  x490 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x527 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x671 &  x674 &  x677 &  x680 &  x689 &  x692 &  x698 &  x704 &  x707 &  x710 &  x713 &  x716 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x743 &  x746 &  x749 &  x752 &  x755 &  x761 &  x764 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x800 &  x803 &  x812 &  x815 &  x818 &  x821 &  x827 &  x830 &  x833 &  x836 &  x839 &  x845 &  x851 &  x857 &  x860 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x914 &  x917 &  x920 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x947 &  x953 &  x959 &  x962 &  x965 &  x971 &  x974 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1055 &  x1058 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x252 & ~x573 & ~x612 & ~x613 & ~x729 & ~x768 & ~x882 & ~x999;
assign c2206 =  x2 &  x8 &  x11 &  x14 &  x20 &  x29 &  x35 &  x41 &  x44 &  x50 &  x65 &  x68 &  x71 &  x74 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x194 &  x212 &  x215 &  x218 &  x230 &  x233 &  x236 &  x238 &  x242 &  x245 &  x248 &  x254 &  x257 &  x263 &  x266 &  x269 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x296 &  x299 &  x302 &  x308 &  x311 &  x314 &  x316 &  x317 &  x320 &  x326 &  x329 &  x332 &  x341 &  x347 &  x353 &  x355 &  x356 &  x359 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x395 &  x398 &  x404 &  x407 &  x413 &  x416 &  x425 &  x428 &  x434 &  x446 &  x449 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x479 &  x482 &  x485 &  x491 &  x494 &  x497 &  x506 &  x509 &  x512 &  x518 &  x521 &  x524 &  x533 &  x536 &  x542 &  x551 &  x554 &  x560 &  x566 &  x575 &  x578 &  x584 &  x587 &  x590 &  x593 &  x599 &  x608 &  x611 &  x614 &  x623 &  x626 &  x632 &  x638 &  x644 &  x647 &  x650 &  x653 &  x659 &  x662 &  x665 &  x671 &  x674 &  x677 &  x683 &  x686 &  x692 &  x698 &  x701 &  x704 &  x707 &  x713 &  x719 &  x722 &  x725 &  x728 &  x731 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x761 &  x764 &  x770 &  x776 &  x782 &  x785 &  x788 &  x791 &  x794 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x845 &  x848 &  x851 &  x857 &  x863 &  x866 &  x872 &  x875 &  x881 &  x887 &  x890 &  x899 &  x908 &  x911 &  x914 &  x917 &  x923 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x953 &  x956 &  x962 &  x968 &  x977 &  x980 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1013 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1049 &  x1052 &  x1058 &  x1061 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x0 & ~x261 & ~x474 & ~x555 & ~x585 & ~x624 & ~x627 & ~x663 & ~x666 & ~x705 & ~x744 & ~x1041 & ~x1080;
assign c2208 =  x2 &  x5 &  x7 &  x8 &  x11 &  x14 &  x17 &  x23 &  x26 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x86 &  x89 &  x92 &  x95 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x194 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x224 &  x233 &  x236 &  x239 &  x242 &  x245 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x284 &  x287 &  x290 &  x296 &  x299 &  x308 &  x311 &  x313 &  x317 &  x323 &  x326 &  x329 &  x335 &  x338 &  x341 &  x344 &  x350 &  x353 &  x356 &  x359 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x386 &  x392 &  x395 &  x401 &  x404 &  x410 &  x413 &  x416 &  x422 &  x425 &  x431 &  x434 &  x437 &  x440 &  x449 &  x452 &  x458 &  x461 &  x467 &  x476 &  x479 &  x491 &  x494 &  x497 &  x500 &  x502 &  x503 &  x509 &  x512 &  x515 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x557 &  x560 &  x569 &  x572 &  x575 &  x578 &  x581 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x614 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x671 &  x674 &  x677 &  x680 &  x683 &  x691 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x713 &  x716 &  x718 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x767 &  x773 &  x776 &  x779 &  x782 &  x788 &  x794 &  x797 &  x800 &  x803 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x845 &  x854 &  x863 &  x866 &  x869 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1046 &  x1049 &  x1055 &  x1061 &  x1064 &  x1067 &  x1073 &  x1079 &  x1082 &  x1085 &  x1091 &  x1100 &  x1103 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x324 & ~x363 & ~x375 & ~x402 & ~x435 & ~x474 & ~x627 & ~x666 & ~x744;
assign c2210 =  x2 &  x8 &  x23 &  x26 &  x41 &  x43 &  x44 &  x50 &  x53 &  x56 &  x59 &  x65 &  x68 &  x74 &  x77 &  x80 &  x81 &  x83 &  x92 &  x95 &  x101 &  x110 &  x113 &  x120 &  x122 &  x134 &  x137 &  x143 &  x146 &  x149 &  x152 &  x158 &  x159 &  x160 &  x161 &  x164 &  x170 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x212 &  x218 &  x221 &  x224 &  x230 &  x233 &  x238 &  x239 &  x242 &  x248 &  x251 &  x257 &  x260 &  x263 &  x269 &  x278 &  x284 &  x290 &  x293 &  x305 &  x308 &  x314 &  x316 &  x320 &  x323 &  x326 &  x329 &  x335 &  x338 &  x341 &  x344 &  x350 &  x356 &  x359 &  x365 &  x368 &  x371 &  x374 &  x377 &  x386 &  x389 &  x395 &  x398 &  x401 &  x425 &  x428 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x470 &  x479 &  x497 &  x500 &  x503 &  x506 &  x518 &  x530 &  x533 &  x539 &  x551 &  x557 &  x560 &  x575 &  x578 &  x584 &  x587 &  x596 &  x599 &  x602 &  x605 &  x608 &  x614 &  x617 &  x620 &  x623 &  x638 &  x653 &  x656 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x683 &  x686 &  x689 &  x701 &  x704 &  x707 &  x713 &  x716 &  x719 &  x734 &  x737 &  x746 &  x749 &  x752 &  x757 &  x758 &  x764 &  x770 &  x773 &  x782 &  x788 &  x794 &  x803 &  x812 &  x815 &  x821 &  x824 &  x830 &  x836 &  x842 &  x845 &  x848 &  x857 &  x863 &  x869 &  x884 &  x887 &  x890 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x929 &  x935 &  x938 &  x940 &  x941 &  x950 &  x953 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x979 &  x980 &  x998 &  x1004 &  x1007 &  x1016 &  x1017 &  x1018 &  x1019 &  x1025 &  x1037 &  x1043 &  x1049 &  x1052 &  x1061 &  x1073 &  x1079 &  x1082 &  x1085 &  x1091 &  x1096 &  x1106 &  x1109 &  x1112 &  x1121 &  x1127 & ~x702 & ~x780;
assign c2212 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x358 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x439 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x539 &  x542 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x614 &  x617 &  x620 &  x623 &  x625 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x758 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x860 &  x863 &  x866 &  x869 &  x872 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x612 & ~x786 & ~x825 & ~x831 & ~x864 & ~x870 & ~x900 & ~x903 & ~x939 & ~x978;
assign c2214 =  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x29 &  x32 &  x35 &  x41 &  x44 &  x47 &  x50 &  x56 &  x59 &  x65 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x97 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x122 &  x125 &  x128 &  x131 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x320 &  x323 &  x326 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x392 &  x395 &  x398 &  x401 &  x404 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x434 &  x437 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x530 &  x533 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x583 &  x584 &  x590 &  x596 &  x599 &  x601 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x622 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x656 &  x659 &  x662 &  x671 &  x674 &  x677 &  x679 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x713 &  x716 &  x718 &  x719 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x757 &  x758 &  x761 &  x764 &  x770 &  x773 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x796 &  x797 &  x800 &  x803 &  x806 &  x809 &  x814 &  x818 &  x821 &  x827 &  x834 &  x835 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x853 &  x857 &  x860 &  x863 &  x866 &  x868 &  x869 &  x874 &  x875 &  x878 &  x884 &  x887 &  x890 &  x892 &  x893 &  x899 &  x902 &  x913 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x931 &  x932 &  x935 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x983 &  x986 &  x989 &  x991 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1030 &  x1031 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1127;
assign c2216 =  x2 &  x11 &  x17 &  x23 &  x35 &  x38 &  x44 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x119 &  x122 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x164 &  x173 &  x176 &  x179 &  x188 &  x194 &  x197 &  x203 &  x206 &  x209 &  x212 &  x218 &  x224 &  x233 &  x239 &  x242 &  x245 &  x248 &  x254 &  x257 &  x260 &  x266 &  x269 &  x278 &  x281 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x314 &  x317 &  x323 &  x326 &  x329 &  x332 &  x335 &  x341 &  x347 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x431 &  x437 &  x440 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x470 &  x476 &  x479 &  x482 &  x485 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x527 &  x530 &  x533 &  x536 &  x545 &  x548 &  x553 &  x554 &  x557 &  x560 &  x563 &  x572 &  x575 &  x581 &  x584 &  x587 &  x593 &  x599 &  x605 &  x608 &  x617 &  x629 &  x635 &  x638 &  x641 &  x653 &  x656 &  x659 &  x662 &  x665 &  x671 &  x674 &  x677 &  x686 &  x692 &  x698 &  x701 &  x707 &  x710 &  x712 &  x713 &  x716 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x743 &  x746 &  x749 &  x758 &  x764 &  x767 &  x773 &  x779 &  x782 &  x788 &  x794 &  x797 &  x800 &  x803 &  x806 &  x812 &  x815 &  x824 &  x827 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x854 &  x857 &  x858 &  x860 &  x863 &  x869 &  x878 &  x887 &  x890 &  x896 &  x898 &  x902 &  x905 &  x908 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x937 &  x941 &  x944 &  x947 &  x950 &  x956 &  x959 &  x968 &  x971 &  x974 &  x975 &  x976 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1048 &  x1052 &  x1053 &  x1054 &  x1058 &  x1061 &  x1064 &  x1070 &  x1076 &  x1085 &  x1088 &  x1091 &  x1093 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x354 & ~x393 & ~x549 & ~x903 & ~x1020 & ~x1059 & ~x1098 & ~x1116;
assign c2218 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x128 &  x131 &  x137 &  x140 &  x143 &  x146 &  x152 &  x158 &  x161 &  x167 &  x170 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x433 &  x434 &  x440 &  x443 &  x446 &  x449 &  x455 &  x458 &  x464 &  x467 &  x470 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x581 &  x584 &  x590 &  x593 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x632 &  x638 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x697 &  x698 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x731 &  x734 &  x736 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x117 & ~x156 & ~x195 & ~x234 & ~x273 & ~x648 & ~x687 & ~x726 & ~x747 & ~x786 & ~x900 & ~x939 & ~x978;
assign c2220 =  x2 &  x5 &  x8 &  x11 &  x17 &  x29 &  x32 &  x38 &  x44 &  x47 &  x53 &  x59 &  x62 &  x65 &  x70 &  x71 &  x74 &  x77 &  x86 &  x95 &  x104 &  x113 &  x116 &  x119 &  x128 &  x131 &  x134 &  x137 &  x143 &  x146 &  x152 &  x155 &  x170 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x212 &  x215 &  x218 &  x221 &  x224 &  x242 &  x245 &  x251 &  x254 &  x263 &  x266 &  x269 &  x272 &  x284 &  x287 &  x293 &  x299 &  x302 &  x311 &  x314 &  x317 &  x319 &  x320 &  x326 &  x329 &  x331 &  x332 &  x335 &  x341 &  x344 &  x353 &  x358 &  x359 &  x362 &  x368 &  x371 &  x383 &  x386 &  x392 &  x395 &  x398 &  x407 &  x410 &  x413 &  x416 &  x419 &  x428 &  x434 &  x446 &  x449 &  x461 &  x464 &  x470 &  x476 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x518 &  x524 &  x536 &  x539 &  x545 &  x548 &  x551 &  x557 &  x566 &  x572 &  x575 &  x581 &  x587 &  x590 &  x593 &  x596 &  x599 &  x608 &  x611 &  x614 &  x617 &  x626 &  x629 &  x641 &  x644 &  x659 &  x662 &  x665 &  x668 &  x674 &  x683 &  x689 &  x695 &  x701 &  x710 &  x722 &  x731 &  x737 &  x740 &  x743 &  x758 &  x767 &  x776 &  x788 &  x800 &  x809 &  x818 &  x821 &  x824 &  x827 &  x830 &  x836 &  x842 &  x845 &  x848 &  x853 &  x854 &  x857 &  x860 &  x863 &  x869 &  x872 &  x875 &  x884 &  x887 &  x890 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x920 &  x923 &  x932 &  x935 &  x937 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x968 &  x971 &  x974 &  x976 &  x991 &  x992 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1022 &  x1028 &  x1037 &  x1043 &  x1052 &  x1055 &  x1058 &  x1061 &  x1063 &  x1064 &  x1067 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1093 &  x1097 &  x1100 &  x1103 &  x1109 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x675;
assign c2222 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x140 &  x143 &  x146 &  x149 &  x152 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x188 &  x191 &  x194 &  x197 &  x203 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x236 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x266 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x296 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x322 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x353 &  x355 &  x356 &  x359 &  x361 &  x362 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x433 &  x434 &  x437 &  x440 &  x446 &  x449 &  x455 &  x458 &  x461 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x545 &  x554 &  x563 &  x566 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x638 &  x641 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x761 &  x764 &  x770 &  x773 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x860 &  x863 &  x866 &  x869 &  x872 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x926 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1100 &  x1103 &  x1109 &  x1115 &  x1127 &  x1130 & ~x156 & ~x195 & ~x378 & ~x381 & ~x417 & ~x513 & ~x534 & ~x552 & ~x783;
assign c2224 =  x2 &  x11 &  x17 &  x20 &  x26 &  x29 &  x32 &  x38 &  x47 &  x56 &  x59 &  x62 &  x68 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x98 &  x101 &  x107 &  x113 &  x116 &  x122 &  x125 &  x128 &  x134 &  x137 &  x142 &  x146 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x184 &  x185 &  x188 &  x191 &  x194 &  x197 &  x203 &  x209 &  x212 &  x215 &  x224 &  x230 &  x233 &  x236 &  x239 &  x251 &  x266 &  x272 &  x275 &  x284 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x320 &  x323 &  x326 &  x335 &  x347 &  x353 &  x356 &  x359 &  x365 &  x368 &  x371 &  x374 &  x377 &  x383 &  x389 &  x407 &  x410 &  x416 &  x422 &  x425 &  x428 &  x434 &  x437 &  x440 &  x443 &  x449 &  x455 &  x458 &  x461 &  x464 &  x467 &  x488 &  x491 &  x500 &  x503 &  x506 &  x511 &  x512 &  x515 &  x518 &  x533 &  x536 &  x542 &  x550 &  x551 &  x557 &  x560 &  x563 &  x572 &  x584 &  x587 &  x590 &  x593 &  x596 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x635 &  x641 &  x647 &  x656 &  x659 &  x668 &  x671 &  x701 &  x704 &  x707 &  x713 &  x734 &  x737 &  x743 &  x746 &  x755 &  x761 &  x764 &  x770 &  x773 &  x776 &  x779 &  x785 &  x791 &  x797 &  x809 &  x812 &  x818 &  x821 &  x827 &  x830 &  x836 &  x842 &  x845 &  x848 &  x851 &  x866 &  x878 &  x890 &  x905 &  x911 &  x914 &  x917 &  x926 &  x929 &  x932 &  x938 &  x944 &  x947 &  x950 &  x962 &  x965 &  x971 &  x980 &  x983 &  x986 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1025 &  x1031 &  x1034 &  x1037 &  x1049 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1091 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1130 & ~x519 & ~x558 & ~x675 & ~x792 & ~x843 & ~x882 & ~x909;
assign c2226 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x260 &  x263 &  x266 &  x269 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x781 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x815 &  x818 &  x820 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x893 &  x896 &  x899 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x441 & ~x480 & ~x519 & ~x753 & ~x792 & ~x831 & ~x832 & ~x870 & ~x871 & ~x882 & ~x909 & ~x921 & ~x948 & ~x1056 & ~x1095;
assign c2228 =  x2 &  x8 &  x17 &  x20 &  x23 &  x26 &  x29 &  x35 &  x38 &  x47 &  x50 &  x59 &  x65 &  x68 &  x77 &  x83 &  x86 &  x89 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x128 &  x131 &  x134 &  x137 &  x143 &  x146 &  x149 &  x152 &  x155 &  x161 &  x164 &  x170 &  x173 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x206 &  x212 &  x215 &  x218 &  x221 &  x230 &  x251 &  x260 &  x266 &  x272 &  x278 &  x284 &  x287 &  x290 &  x293 &  x305 &  x311 &  x313 &  x314 &  x317 &  x323 &  x326 &  x329 &  x332 &  x338 &  x341 &  x344 &  x350 &  x353 &  x362 &  x365 &  x371 &  x377 &  x380 &  x386 &  x392 &  x398 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x428 &  x431 &  x434 &  x443 &  x446 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x524 &  x530 &  x536 &  x542 &  x545 &  x551 &  x557 &  x560 &  x566 &  x572 &  x575 &  x578 &  x581 &  x584 &  x593 &  x596 &  x599 &  x611 &  x617 &  x620 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x647 &  x653 &  x656 &  x659 &  x662 &  x671 &  x674 &  x680 &  x683 &  x686 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x722 &  x725 &  x728 &  x737 &  x740 &  x743 &  x752 &  x758 &  x761 &  x764 &  x767 &  x770 &  x779 &  x782 &  x785 &  x797 &  x800 &  x803 &  x809 &  x812 &  x815 &  x824 &  x836 &  x839 &  x842 &  x845 &  x851 &  x854 &  x857 &  x860 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x950 &  x953 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x983 &  x989 &  x992 &  x1000 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1039 &  x1043 &  x1046 &  x1051 &  x1052 &  x1058 &  x1064 &  x1070 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x435 & ~x453 & ~x474 & ~x513 & ~x552 & ~x585 & ~x627 & ~x666 & ~x705 & ~x744 & ~x822 & ~x861 & ~x897 & ~x900 & ~x936 & ~x939 & ~x975 & ~x1014 & ~x1053 & ~x1092;
assign c2230 =  x5 &  x8 &  x11 &  x17 &  x20 &  x23 &  x32 &  x35 &  x44 &  x50 &  x53 &  x56 &  x59 &  x62 &  x71 &  x77 &  x83 &  x86 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x116 &  x122 &  x125 &  x128 &  x137 &  x155 &  x158 &  x164 &  x170 &  x182 &  x188 &  x191 &  x194 &  x197 &  x206 &  x209 &  x212 &  x218 &  x221 &  x227 &  x230 &  x233 &  x236 &  x242 &  x248 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x326 &  x329 &  x335 &  x338 &  x341 &  x344 &  x350 &  x353 &  x359 &  x365 &  x371 &  x374 &  x377 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x430 &  x431 &  x433 &  x440 &  x446 &  x455 &  x458 &  x467 &  x469 &  x476 &  x479 &  x482 &  x494 &  x497 &  x500 &  x503 &  x508 &  x512 &  x521 &  x524 &  x527 &  x533 &  x536 &  x542 &  x545 &  x547 &  x548 &  x554 &  x560 &  x563 &  x572 &  x575 &  x578 &  x581 &  x586 &  x593 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x625 &  x629 &  x632 &  x635 &  x638 &  x644 &  x647 &  x653 &  x656 &  x665 &  x668 &  x674 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x710 &  x716 &  x728 &  x731 &  x734 &  x737 &  x749 &  x761 &  x767 &  x773 &  x779 &  x782 &  x785 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x842 &  x845 &  x848 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x887 &  x899 &  x902 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x956 &  x959 &  x968 &  x971 &  x974 &  x977 &  x980 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1067 &  x1073 &  x1076 &  x1082 &  x1088 &  x1100 &  x1106 &  x1109 &  x1112 &  x1121 &  x1124 &  x1127 & ~x342 & ~x381 & ~x420 & ~x513 & ~x552 & ~x630 & ~x633 & ~x783 & ~x822 & ~x825 & ~x864;
assign c2232 =  x2 &  x5 &  x11 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x41 &  x47 &  x50 &  x56 &  x59 &  x65 &  x71 &  x74 &  x77 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x119 &  x122 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x164 &  x167 &  x170 &  x173 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x233 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x281 &  x287 &  x290 &  x293 &  x296 &  x302 &  x305 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x335 &  x338 &  x341 &  x344 &  x347 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x416 &  x422 &  x425 &  x428 &  x431 &  x434 &  x440 &  x443 &  x452 &  x455 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x506 &  x509 &  x512 &  x518 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x545 &  x551 &  x554 &  x557 &  x560 &  x566 &  x572 &  x575 &  x578 &  x581 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x629 &  x638 &  x641 &  x647 &  x650 &  x653 &  x656 &  x659 &  x665 &  x668 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x704 &  x710 &  x713 &  x716 &  x719 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x797 &  x800 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x911 &  x914 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x950 &  x962 &  x968 &  x971 &  x974 &  x977 &  x983 &  x989 &  x992 &  x995 &  x1001 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1073 &  x1079 &  x1082 &  x1088 &  x1097 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x402 & ~x441 & ~x480 & ~x519 & ~x570 & ~x609 & ~x648 & ~x675 & ~x687 & ~x747 & ~x765 & ~x792 & ~x804 & ~x843 & ~x861 & ~x882 & ~x900 & ~x939 & ~x978 & ~x1095;
assign c2234 =  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x92 &  x98 &  x104 &  x107 &  x110 &  x119 &  x122 &  x128 &  x131 &  x134 &  x140 &  x143 &  x146 &  x152 &  x155 &  x158 &  x161 &  x167 &  x170 &  x173 &  x176 &  x179 &  x188 &  x191 &  x197 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x293 &  x296 &  x299 &  x302 &  x305 &  x311 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x344 &  x347 &  x350 &  x353 &  x356 &  x362 &  x368 &  x370 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x479 &  x482 &  x485 &  x491 &  x494 &  x497 &  x500 &  x503 &  x509 &  x512 &  x515 &  x518 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x566 &  x569 &  x572 &  x575 &  x581 &  x584 &  x587 &  x590 &  x593 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x629 &  x632 &  x635 &  x641 &  x647 &  x650 &  x653 &  x659 &  x662 &  x665 &  x671 &  x674 &  x680 &  x686 &  x692 &  x695 &  x698 &  x704 &  x707 &  x710 &  x716 &  x722 &  x725 &  x728 &  x731 &  x737 &  x743 &  x746 &  x752 &  x755 &  x758 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x794 &  x797 &  x803 &  x809 &  x812 &  x815 &  x818 &  x821 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x872 &  x875 &  x878 &  x881 &  x887 &  x893 &  x896 &  x899 &  x905 &  x908 &  x911 &  x913 &  x914 &  x917 &  x920 &  x929 &  x932 &  x935 &  x937 &  x938 &  x944 &  x946 &  x947 &  x950 &  x952 &  x953 &  x956 &  x959 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x991 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1069 &  x1070 &  x1073 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130 & ~x942 & ~x948 & ~x987 & ~x988 & ~x1065;
assign c2236 =  x17 &  x23 &  x32 &  x35 &  x47 &  x50 &  x56 &  x65 &  x71 &  x83 &  x86 &  x101 &  x113 &  x116 &  x131 &  x137 &  x146 &  x158 &  x170 &  x173 &  x185 &  x203 &  x209 &  x227 &  x230 &  x251 &  x254 &  x257 &  x272 &  x293 &  x302 &  x308 &  x317 &  x320 &  x332 &  x335 &  x341 &  x353 &  x356 &  x358 &  x362 &  x365 &  x377 &  x386 &  x392 &  x401 &  x407 &  x419 &  x425 &  x437 &  x440 &  x446 &  x452 &  x455 &  x458 &  x461 &  x470 &  x473 &  x475 &  x482 &  x488 &  x497 &  x500 &  x503 &  x509 &  x512 &  x515 &  x518 &  x524 &  x530 &  x533 &  x539 &  x548 &  x557 &  x560 &  x566 &  x569 &  x581 &  x593 &  x599 &  x605 &  x608 &  x614 &  x620 &  x641 &  x647 &  x650 &  x659 &  x662 &  x665 &  x668 &  x680 &  x689 &  x692 &  x698 &  x701 &  x707 &  x713 &  x716 &  x719 &  x731 &  x737 &  x743 &  x764 &  x770 &  x782 &  x788 &  x800 &  x806 &  x812 &  x818 &  x820 &  x821 &  x824 &  x842 &  x845 &  x848 &  x857 &  x860 &  x872 &  x881 &  x890 &  x893 &  x905 &  x908 &  x920 &  x923 &  x926 &  x929 &  x956 &  x962 &  x965 &  x974 &  x980 &  x986 &  x1001 &  x1007 &  x1037 &  x1049 &  x1061 &  x1064 &  x1073 &  x1076 &  x1085 &  x1088 &  x1097 &  x1103 &  x1109 &  x1118 &  x1121 &  x1127 & ~x198 & ~x276 & ~x765 & ~x870 & ~x904 & ~x942 & ~x1056;
assign c2238 =  x2 &  x5 &  x8 &  x11 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x128 &  x131 &  x134 &  x137 &  x143 &  x146 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x680 &  x683 &  x686 &  x689 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x722 &  x725 &  x728 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x878 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x995 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x285 & ~x324 & ~x363 & ~x402 & ~x441 & ~x480 & ~x519 & ~x531 & ~x564 & ~x570 & ~x603 & ~x609 & ~x648 & ~x675 & ~x687 & ~x714 & ~x831 & ~x861 & ~x870 & ~x900 & ~x939 & ~x978 & ~x1017;
assign c2240 =  x8 &  x11 &  x14 &  x17 &  x23 &  x26 &  x32 &  x35 &  x38 &  x41 &  x44 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x116 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x185 &  x191 &  x194 &  x197 &  x200 &  x203 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x476 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x580 &  x581 &  x584 &  x587 &  x593 &  x596 &  x599 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x622 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x658 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x683 &  x689 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x812 &  x815 &  x818 &  x821 &  x824 &  x830 &  x833 &  x835 &  x836 &  x839 &  x842 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x920 &  x923 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x950 &  x953 &  x965 &  x968 &  x971 &  x980 &  x989 &  x1001 &  x1007 &  x1010 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1103 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x0 & ~x33 & ~x72 & ~x171;
assign c2242 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x35 &  x38 &  x41 &  x50 &  x53 &  x62 &  x65 &  x68 &  x74 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x107 &  x110 &  x113 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x158 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x203 &  x206 &  x209 &  x212 &  x218 &  x221 &  x224 &  x227 &  x230 &  x232 &  x233 &  x236 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x293 &  x299 &  x302 &  x305 &  x308 &  x310 &  x311 &  x314 &  x317 &  x320 &  x323 &  x329 &  x332 &  x335 &  x341 &  x344 &  x349 &  x350 &  x356 &  x359 &  x362 &  x371 &  x374 &  x376 &  x377 &  x380 &  x386 &  x389 &  x392 &  x395 &  x397 &  x398 &  x401 &  x404 &  x407 &  x413 &  x416 &  x422 &  x425 &  x431 &  x434 &  x436 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x470 &  x473 &  x475 &  x476 &  x478 &  x479 &  x482 &  x488 &  x494 &  x497 &  x500 &  x503 &  x506 &  x515 &  x518 &  x521 &  x527 &  x530 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x575 &  x578 &  x593 &  x596 &  x602 &  x605 &  x608 &  x614 &  x617 &  x620 &  x623 &  x629 &  x632 &  x635 &  x638 &  x644 &  x647 &  x650 &  x656 &  x659 &  x662 &  x665 &  x671 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x713 &  x719 &  x722 &  x725 &  x728 &  x731 &  x737 &  x740 &  x743 &  x746 &  x749 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x788 &  x791 &  x794 &  x797 &  x806 &  x809 &  x818 &  x821 &  x824 &  x827 &  x833 &  x836 &  x839 &  x842 &  x851 &  x853 &  x854 &  x856 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x878 &  x881 &  x890 &  x892 &  x893 &  x896 &  x899 &  x905 &  x908 &  x911 &  x914 &  x920 &  x929 &  x931 &  x932 &  x938 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x968 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1034 &  x1037 &  x1046 &  x1048 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1087 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 & ~x312 & ~x351 & ~x390 & ~x429;
assign c2244 =  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x44 &  x47 &  x50 &  x53 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x166 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x203 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x244 &  x245 &  x248 &  x254 &  x257 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x283 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x314 &  x317 &  x320 &  x322 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x361 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x383 &  x386 &  x389 &  x391 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x430 &  x431 &  x434 &  x437 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x601 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x623 &  x629 &  x632 &  x635 &  x640 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x988 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1027 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1066 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x396 & ~x435 & ~x474 & ~x513 & ~x552 & ~x975 & ~x1014;
assign c2246 =  x2 &  x5 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x83 &  x86 &  x89 &  x92 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x121 &  x125 &  x128 &  x131 &  x134 &  x140 &  x146 &  x149 &  x155 &  x158 &  x160 &  x161 &  x164 &  x167 &  x176 &  x179 &  x182 &  x185 &  x191 &  x194 &  x199 &  x200 &  x203 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x263 &  x269 &  x272 &  x275 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x355 &  x356 &  x362 &  x368 &  x371 &  x374 &  x377 &  x380 &  x386 &  x392 &  x395 &  x404 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x473 &  x476 &  x479 &  x482 &  x485 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x557 &  x563 &  x569 &  x575 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x614 &  x617 &  x620 &  x623 &  x626 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x656 &  x659 &  x662 &  x671 &  x674 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x776 &  x779 &  x782 &  x785 &  x791 &  x794 &  x797 &  x800 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x872 &  x878 &  x881 &  x884 &  x887 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x917 &  x920 &  x923 &  x926 &  x929 &  x935 &  x938 &  x950 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1028 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1061 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x258 & ~x298 & ~x336 & ~x337 & ~x375 & ~x414 & ~x453 & ~x510 & ~x513 & ~x627 & ~x666 & ~x705 & ~x744;
assign c2248 =  x5 &  x11 &  x14 &  x17 &  x23 &  x26 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x59 &  x62 &  x68 &  x80 &  x83 &  x86 &  x89 &  x95 &  x98 &  x101 &  x107 &  x113 &  x119 &  x128 &  x131 &  x137 &  x146 &  x149 &  x152 &  x161 &  x164 &  x170 &  x178 &  x179 &  x191 &  x194 &  x197 &  x209 &  x212 &  x218 &  x221 &  x224 &  x233 &  x236 &  x239 &  x242 &  x245 &  x254 &  x256 &  x257 &  x266 &  x269 &  x272 &  x275 &  x278 &  x284 &  x287 &  x290 &  x296 &  x299 &  x305 &  x311 &  x314 &  x317 &  x320 &  x329 &  x332 &  x344 &  x347 &  x350 &  x359 &  x368 &  x371 &  x373 &  x374 &  x377 &  x380 &  x383 &  x389 &  x392 &  x404 &  x407 &  x413 &  x422 &  x425 &  x428 &  x431 &  x437 &  x440 &  x443 &  x449 &  x452 &  x461 &  x467 &  x470 &  x473 &  x476 &  x485 &  x488 &  x494 &  x500 &  x503 &  x509 &  x512 &  x518 &  x521 &  x524 &  x527 &  x536 &  x539 &  x542 &  x545 &  x551 &  x557 &  x560 &  x563 &  x566 &  x572 &  x578 &  x584 &  x587 &  x590 &  x599 &  x605 &  x608 &  x611 &  x617 &  x623 &  x632 &  x644 &  x647 &  x653 &  x656 &  x659 &  x665 &  x668 &  x674 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x704 &  x713 &  x719 &  x731 &  x734 &  x736 &  x758 &  x761 &  x770 &  x773 &  x775 &  x785 &  x788 &  x791 &  x794 &  x800 &  x803 &  x809 &  x812 &  x815 &  x824 &  x835 &  x836 &  x842 &  x845 &  x848 &  x851 &  x854 &  x860 &  x872 &  x875 &  x878 &  x884 &  x887 &  x890 &  x892 &  x893 &  x896 &  x905 &  x911 &  x913 &  x920 &  x926 &  x929 &  x935 &  x941 &  x944 &  x947 &  x950 &  x959 &  x962 &  x971 &  x974 &  x977 &  x983 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1069 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1088 &  x1094 &  x1097 &  x1103 &  x1109 &  x1112 &  x1124 &  x1127 & ~x531 & ~x570 & ~x609 & ~x633 & ~x648 & ~x822;
assign c2250 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x188 &  x191 &  x194 &  x197 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x256 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x332 &  x334 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x373 &  x374 &  x377 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x419 &  x422 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x542 &  x545 &  x548 &  x554 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x622 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x653 &  x656 &  x659 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x685 &  x686 &  x689 &  x692 &  x695 &  x701 &  x704 &  x709 &  x710 &  x713 &  x716 &  x718 &  x722 &  x724 &  x725 &  x727 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x752 &  x755 &  x757 &  x758 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x796 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x830 &  x833 &  x835 &  x836 &  x839 &  x842 &  x845 &  x854 &  x857 &  x860 &  x866 &  x869 &  x872 &  x874 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x905 &  x911 &  x913 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x994 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1072 &  x1073 &  x1076 &  x1079 &  x1088 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x93;
assign c2252 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x35 &  x44 &  x47 &  x53 &  x56 &  x62 &  x65 &  x68 &  x71 &  x73 &  x74 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x137 &  x140 &  x143 &  x149 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x176 &  x182 &  x187 &  x188 &  x191 &  x197 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x226 &  x227 &  x230 &  x236 &  x239 &  x242 &  x245 &  x251 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x359 &  x371 &  x374 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x464 &  x467 &  x473 &  x476 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x542 &  x545 &  x551 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x626 &  x629 &  x635 &  x638 &  x644 &  x650 &  x653 &  x656 &  x659 &  x662 &  x668 &  x671 &  x689 &  x692 &  x695 &  x698 &  x704 &  x707 &  x713 &  x716 &  x719 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x773 &  x776 &  x782 &  x785 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x839 &  x842 &  x845 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x938 &  x941 &  x944 &  x947 &  x953 &  x959 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x992 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1048 &  x1049 &  x1052 &  x1054 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1085 &  x1091 &  x1093 &  x1100 &  x1103 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 & ~x234 & ~x273 & ~x312 & ~x351 & ~x390 & ~x837 & ~x843 & ~x882 & ~x942 & ~x999 & ~x1038;
assign c2254 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x310 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x415 &  x416 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x454 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x521 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x66 & ~x573 & ~x615 & ~x654 & ~x768 & ~x906;
assign c2256 =  x2 &  x11 &  x14 &  x35 &  x38 &  x43 &  x59 &  x65 &  x68 &  x74 &  x82 &  x86 &  x95 &  x110 &  x116 &  x119 &  x140 &  x143 &  x146 &  x170 &  x173 &  x185 &  x197 &  x206 &  x218 &  x224 &  x242 &  x245 &  x251 &  x254 &  x260 &  x269 &  x284 &  x287 &  x296 &  x302 &  x308 &  x320 &  x329 &  x350 &  x353 &  x365 &  x374 &  x386 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x434 &  x440 &  x446 &  x467 &  x470 &  x473 &  x479 &  x482 &  x497 &  x521 &  x536 &  x545 &  x548 &  x551 &  x560 &  x590 &  x617 &  x629 &  x635 &  x641 &  x650 &  x680 &  x683 &  x686 &  x692 &  x698 &  x710 &  x725 &  x728 &  x731 &  x734 &  x737 &  x743 &  x746 &  x752 &  x755 &  x767 &  x775 &  x776 &  x782 &  x788 &  x800 &  x816 &  x830 &  x839 &  x842 &  x845 &  x851 &  x854 &  x860 &  x863 &  x866 &  x875 &  x887 &  x911 &  x920 &  x929 &  x935 &  x941 &  x953 &  x956 &  x959 &  x965 &  x977 &  x986 &  x989 &  x998 &  x1016 &  x1019 &  x1022 &  x1037 &  x1046 &  x1058 &  x1063 &  x1067 &  x1079 &  x1085 &  x1088 &  x1091 &  x1100 &  x1109 &  x1112 &  x1121 & ~x753;
assign c2258 =  x2 &  x8 &  x11 &  x14 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x42 &  x43 &  x44 &  x50 &  x56 &  x59 &  x62 &  x65 &  x71 &  x74 &  x77 &  x80 &  x81 &  x82 &  x83 &  x86 &  x89 &  x92 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x120 &  x121 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x155 &  x158 &  x160 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x197 &  x203 &  x209 &  x218 &  x221 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x275 &  x278 &  x284 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x317 &  x320 &  x323 &  x329 &  x332 &  x344 &  x346 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x392 &  x395 &  x401 &  x407 &  x410 &  x413 &  x422 &  x425 &  x428 &  x431 &  x440 &  x443 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x470 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x542 &  x545 &  x548 &  x554 &  x557 &  x563 &  x566 &  x569 &  x572 &  x575 &  x581 &  x584 &  x587 &  x593 &  x596 &  x599 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x626 &  x629 &  x641 &  x644 &  x656 &  x659 &  x662 &  x665 &  x671 &  x674 &  x677 &  x680 &  x683 &  x689 &  x692 &  x698 &  x701 &  x704 &  x707 &  x713 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x743 &  x746 &  x749 &  x752 &  x758 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x788 &  x794 &  x797 &  x803 &  x809 &  x812 &  x815 &  x818 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x887 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x917 &  x920 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x986 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1100 &  x1103 &  x1109 &  x1115 &  x1124 &  x1127 &  x1130 & ~x219 & ~x261 & ~x390 & ~x507 & ~x768;
assign c2260 =  x11 &  x14 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x47 &  x50 &  x59 &  x65 &  x71 &  x77 &  x83 &  x86 &  x89 &  x95 &  x98 &  x101 &  x107 &  x116 &  x119 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x155 &  x158 &  x161 &  x164 &  x170 &  x173 &  x179 &  x182 &  x188 &  x191 &  x194 &  x197 &  x200 &  x206 &  x209 &  x215 &  x218 &  x224 &  x230 &  x236 &  x239 &  x242 &  x248 &  x254 &  x266 &  x269 &  x278 &  x281 &  x284 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x320 &  x326 &  x329 &  x335 &  x341 &  x344 &  x353 &  x356 &  x364 &  x365 &  x368 &  x377 &  x383 &  x386 &  x389 &  x392 &  x398 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x458 &  x467 &  x470 &  x475 &  x476 &  x479 &  x485 &  x491 &  x494 &  x497 &  x503 &  x506 &  x509 &  x512 &  x518 &  x527 &  x533 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x560 &  x563 &  x572 &  x578 &  x587 &  x590 &  x593 &  x596 &  x599 &  x608 &  x611 &  x614 &  x623 &  x629 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x659 &  x665 &  x668 &  x671 &  x674 &  x677 &  x683 &  x695 &  x698 &  x707 &  x716 &  x722 &  x731 &  x740 &  x743 &  x746 &  x749 &  x752 &  x770 &  x776 &  x782 &  x785 &  x788 &  x791 &  x797 &  x800 &  x803 &  x809 &  x812 &  x824 &  x827 &  x836 &  x839 &  x845 &  x851 &  x857 &  x863 &  x866 &  x869 &  x872 &  x878 &  x884 &  x890 &  x893 &  x896 &  x899 &  x905 &  x917 &  x923 &  x926 &  x929 &  x932 &  x941 &  x944 &  x950 &  x956 &  x965 &  x971 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1016 &  x1022 &  x1028 &  x1037 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1106 &  x1109 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x135 & ~x273 & ~x312 & ~x351 & ~x468 & ~x942 & ~x948 & ~x1017 & ~x1065;
assign c2262 =  x2 &  x8 &  x14 &  x17 &  x20 &  x29 &  x32 &  x44 &  x53 &  x56 &  x62 &  x77 &  x80 &  x83 &  x86 &  x89 &  x101 &  x107 &  x110 &  x113 &  x116 &  x119 &  x125 &  x128 &  x131 &  x137 &  x140 &  x143 &  x146 &  x155 &  x158 &  x170 &  x173 &  x182 &  x188 &  x191 &  x197 &  x206 &  x215 &  x218 &  x227 &  x230 &  x245 &  x248 &  x254 &  x260 &  x263 &  x275 &  x281 &  x284 &  x293 &  x299 &  x302 &  x311 &  x314 &  x320 &  x326 &  x329 &  x338 &  x341 &  x344 &  x347 &  x353 &  x359 &  x362 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x394 &  x395 &  x401 &  x407 &  x410 &  x416 &  x419 &  x422 &  x425 &  x431 &  x434 &  x437 &  x440 &  x446 &  x449 &  x452 &  x455 &  x464 &  x467 &  x469 &  x470 &  x476 &  x479 &  x482 &  x485 &  x488 &  x494 &  x515 &  x518 &  x524 &  x530 &  x533 &  x536 &  x542 &  x548 &  x551 &  x560 &  x563 &  x569 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x590 &  x593 &  x596 &  x602 &  x608 &  x614 &  x617 &  x620 &  x623 &  x629 &  x632 &  x638 &  x641 &  x647 &  x650 &  x656 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x680 &  x686 &  x689 &  x692 &  x701 &  x704 &  x725 &  x728 &  x737 &  x740 &  x749 &  x761 &  x764 &  x767 &  x773 &  x776 &  x782 &  x797 &  x803 &  x809 &  x812 &  x815 &  x818 &  x821 &  x827 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x860 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x896 &  x899 &  x902 &  x917 &  x920 &  x923 &  x926 &  x935 &  x941 &  x944 &  x947 &  x953 &  x962 &  x968 &  x974 &  x977 &  x983 &  x986 &  x989 &  x1001 &  x1004 &  x1007 &  x1019 &  x1025 &  x1028 &  x1034 &  x1037 &  x1043 &  x1049 &  x1055 &  x1058 &  x1061 &  x1067 &  x1070 &  x1079 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1121 &  x1130 & ~x156 & ~x552 & ~x558 & ~x591 & ~x630 & ~x636 & ~x669 & ~x675 & ~x708 & ~x747 & ~x753 & ~x900 & ~x939;
assign c2264 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x82 &  x83 &  x86 &  x88 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x121 &  x122 &  x125 &  x128 &  x134 &  x137 &  x139 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x157 &  x158 &  x160 &  x161 &  x164 &  x166 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x191 &  x194 &  x196 &  x197 &  x203 &  x205 &  x206 &  x209 &  x215 &  x218 &  x224 &  x227 &  x233 &  x235 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x274 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x311 &  x313 &  x314 &  x317 &  x320 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x398 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x548 &  x551 &  x554 &  x557 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x629 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x809 &  x812 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x988 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1013 &  x1016 &  x1019 &  x1025 &  x1027 &  x1028 &  x1031 &  x1034 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1066 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x258 & ~x297 & ~x492;
assign c2266 =  x2 &  x5 &  x8 &  x11 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x98 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x131 &  x134 &  x146 &  x149 &  x152 &  x155 &  x164 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x227 &  x230 &  x233 &  x236 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x266 &  x269 &  x272 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x320 &  x323 &  x326 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x362 &  x365 &  x368 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x395 &  x401 &  x404 &  x407 &  x410 &  x412 &  x416 &  x419 &  x425 &  x428 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x490 &  x494 &  x497 &  x500 &  x503 &  x506 &  x512 &  x515 &  x518 &  x521 &  x527 &  x533 &  x542 &  x545 &  x548 &  x551 &  x554 &  x556 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x584 &  x587 &  x590 &  x595 &  x596 &  x599 &  x602 &  x607 &  x608 &  x611 &  x614 &  x617 &  x620 &  x626 &  x629 &  x632 &  x638 &  x641 &  x644 &  x646 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x776 &  x779 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x839 &  x841 &  x842 &  x845 &  x848 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x875 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x911 &  x914 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x953 &  x962 &  x965 &  x968 &  x971 &  x974 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1070 &  x1076 &  x1079 &  x1082 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1118 &  x1121 &  x1124 & ~x924 & ~x942 & ~x981 & ~x1059 & ~x1095;
assign c2268 =  x5 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x35 &  x41 &  x44 &  x47 &  x56 &  x62 &  x65 &  x71 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x104 &  x107 &  x110 &  x113 &  x119 &  x122 &  x125 &  x128 &  x131 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x161 &  x167 &  x170 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x200 &  x212 &  x215 &  x221 &  x227 &  x230 &  x233 &  x242 &  x245 &  x248 &  x251 &  x254 &  x260 &  x266 &  x269 &  x272 &  x275 &  x277 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x302 &  x305 &  x308 &  x313 &  x314 &  x317 &  x323 &  x326 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x356 &  x359 &  x362 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x391 &  x392 &  x395 &  x398 &  x404 &  x407 &  x413 &  x416 &  x419 &  x422 &  x428 &  x430 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x469 &  x470 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x509 &  x512 &  x515 &  x518 &  x527 &  x530 &  x533 &  x536 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x578 &  x584 &  x587 &  x590 &  x593 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x626 &  x629 &  x632 &  x638 &  x650 &  x653 &  x659 &  x662 &  x671 &  x674 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x710 &  x713 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x761 &  x770 &  x773 &  x776 &  x782 &  x785 &  x788 &  x791 &  x800 &  x809 &  x815 &  x818 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x854 &  x857 &  x860 &  x863 &  x866 &  x872 &  x875 &  x878 &  x881 &  x884 &  x890 &  x893 &  x896 &  x902 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x474 & ~x531 & ~x570 & ~x609 & ~x726 & ~x744 & ~x786 & ~x822 & ~x861 & ~x862 & ~x900;
assign c2270 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x23 &  x26 &  x29 &  x35 &  x38 &  x41 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x80 &  x83 &  x89 &  x92 &  x98 &  x104 &  x107 &  x113 &  x119 &  x122 &  x125 &  x128 &  x134 &  x137 &  x143 &  x146 &  x155 &  x161 &  x167 &  x170 &  x179 &  x182 &  x185 &  x188 &  x191 &  x197 &  x200 &  x203 &  x212 &  x218 &  x221 &  x224 &  x230 &  x233 &  x236 &  x239 &  x248 &  x251 &  x254 &  x260 &  x266 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x341 &  x344 &  x347 &  x350 &  x353 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x383 &  x386 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x431 &  x437 &  x440 &  x443 &  x446 &  x452 &  x455 &  x458 &  x464 &  x470 &  x473 &  x479 &  x482 &  x485 &  x488 &  x494 &  x497 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x530 &  x539 &  x542 &  x548 &  x551 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x584 &  x587 &  x590 &  x596 &  x599 &  x602 &  x608 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x659 &  x662 &  x668 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x764 &  x767 &  x770 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x800 &  x809 &  x815 &  x818 &  x824 &  x827 &  x833 &  x836 &  x842 &  x845 &  x851 &  x857 &  x860 &  x863 &  x869 &  x872 &  x875 &  x878 &  x884 &  x887 &  x893 &  x899 &  x902 &  x905 &  x908 &  x914 &  x917 &  x929 &  x935 &  x938 &  x941 &  x944 &  x953 &  x956 &  x959 &  x962 &  x965 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1034 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 &  x1130 & ~x222 & ~x223 & ~x261 & ~x456 & ~x495 & ~x496 & ~x534 & ~x535 & ~x573 & ~x574 & ~x609 & ~x612 & ~x711;
assign c2272 =  x5 &  x11 &  x14 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x224 &  x227 &  x230 &  x239 &  x242 &  x248 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x320 &  x326 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x359 &  x362 &  x365 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x440 &  x443 &  x446 &  x449 &  x452 &  x454 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x626 &  x632 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x667 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x784 &  x785 &  x791 &  x794 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x851 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x898 &  x902 &  x905 &  x908 &  x911 &  x917 &  x923 &  x926 &  x929 &  x935 &  x938 &  x941 &  x950 &  x953 &  x956 &  x962 &  x965 &  x968 &  x971 &  x974 &  x976 &  x977 &  x980 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x273 & ~x312 & ~x351 & ~x390 & ~x429 & ~x468 & ~x846 & ~x960 & ~x961 & ~x981 & ~x999 & ~x1020 & ~x1038 & ~x1059;
assign c2274 =  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x26 &  x29 &  x32 &  x41 &  x44 &  x47 &  x49 &  x53 &  x59 &  x62 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x107 &  x110 &  x113 &  x116 &  x121 &  x122 &  x125 &  x128 &  x131 &  x137 &  x140 &  x143 &  x146 &  x149 &  x155 &  x157 &  x158 &  x160 &  x161 &  x166 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x196 &  x197 &  x199 &  x200 &  x203 &  x205 &  x206 &  x209 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x234 &  x235 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x263 &  x266 &  x274 &  x275 &  x278 &  x281 &  x284 &  x290 &  x296 &  x299 &  x305 &  x311 &  x314 &  x317 &  x320 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x350 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x377 &  x380 &  x389 &  x391 &  x392 &  x401 &  x404 &  x407 &  x413 &  x416 &  x419 &  x422 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x503 &  x506 &  x512 &  x515 &  x521 &  x524 &  x533 &  x539 &  x548 &  x551 &  x554 &  x557 &  x563 &  x566 &  x569 &  x575 &  x578 &  x584 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x623 &  x626 &  x629 &  x632 &  x635 &  x641 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x695 &  x701 &  x704 &  x710 &  x713 &  x716 &  x719 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x857 &  x860 &  x863 &  x866 &  x872 &  x875 &  x878 &  x884 &  x887 &  x890 &  x893 &  x896 &  x908 &  x911 &  x914 &  x917 &  x920 &  x926 &  x929 &  x932 &  x935 &  x941 &  x944 &  x947 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x980 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1034 &  x1037 &  x1040 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x186 & ~x225 & ~x264 & ~x279 & ~x318 & ~x474 & ~x588 & ~x627;
assign c2276 =  x8 &  x14 &  x20 &  x23 &  x26 &  x35 &  x38 &  x41 &  x46 &  x50 &  x59 &  x71 &  x74 &  x77 &  x80 &  x83 &  x85 &  x86 &  x89 &  x101 &  x104 &  x107 &  x140 &  x146 &  x170 &  x173 &  x179 &  x188 &  x191 &  x200 &  x206 &  x212 &  x224 &  x227 &  x233 &  x251 &  x254 &  x260 &  x266 &  x269 &  x272 &  x275 &  x278 &  x287 &  x290 &  x311 &  x317 &  x320 &  x323 &  x326 &  x332 &  x335 &  x338 &  x344 &  x353 &  x359 &  x365 &  x368 &  x383 &  x386 &  x389 &  x395 &  x407 &  x416 &  x419 &  x425 &  x449 &  x455 &  x458 &  x461 &  x470 &  x473 &  x479 &  x482 &  x487 &  x506 &  x509 &  x515 &  x518 &  x521 &  x526 &  x527 &  x533 &  x536 &  x544 &  x545 &  x563 &  x565 &  x566 &  x572 &  x581 &  x587 &  x593 &  x601 &  x605 &  x614 &  x623 &  x629 &  x635 &  x638 &  x641 &  x644 &  x653 &  x659 &  x662 &  x668 &  x671 &  x674 &  x680 &  x683 &  x686 &  x698 &  x701 &  x707 &  x713 &  x722 &  x724 &  x725 &  x731 &  x734 &  x743 &  x746 &  x749 &  x752 &  x755 &  x764 &  x770 &  x779 &  x782 &  x788 &  x797 &  x806 &  x812 &  x818 &  x821 &  x824 &  x833 &  x836 &  x838 &  x839 &  x851 &  x854 &  x860 &  x863 &  x869 &  x875 &  x878 &  x881 &  x890 &  x899 &  x902 &  x905 &  x907 &  x908 &  x911 &  x914 &  x916 &  x917 &  x920 &  x926 &  x929 &  x938 &  x944 &  x947 &  x950 &  x962 &  x971 &  x974 &  x980 &  x983 &  x989 &  x992 &  x994 &  x995 &  x1007 &  x1016 &  x1019 &  x1025 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1058 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1100 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 & ~x624;
assign c2278 =  x2 &  x10 &  x11 &  x14 &  x17 &  x20 &  x23 &  x29 &  x32 &  x35 &  x38 &  x41 &  x43 &  x44 &  x47 &  x50 &  x53 &  x56 &  x62 &  x65 &  x68 &  x71 &  x77 &  x80 &  x82 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x107 &  x110 &  x113 &  x116 &  x118 &  x119 &  x121 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x146 &  x149 &  x152 &  x155 &  x157 &  x158 &  x160 &  x161 &  x164 &  x167 &  x170 &  x173 &  x182 &  x185 &  x194 &  x196 &  x197 &  x199 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x260 &  x269 &  x272 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x299 &  x305 &  x307 &  x308 &  x314 &  x317 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x346 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x377 &  x380 &  x383 &  x389 &  x395 &  x398 &  x401 &  x404 &  x407 &  x413 &  x419 &  x422 &  x424 &  x425 &  x428 &  x434 &  x437 &  x440 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x467 &  x470 &  x473 &  x482 &  x485 &  x488 &  x494 &  x500 &  x512 &  x515 &  x518 &  x524 &  x527 &  x533 &  x539 &  x548 &  x551 &  x554 &  x557 &  x560 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x587 &  x595 &  x602 &  x605 &  x611 &  x617 &  x623 &  x626 &  x629 &  x632 &  x634 &  x635 &  x638 &  x644 &  x647 &  x650 &  x656 &  x665 &  x668 &  x671 &  x674 &  x677 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x716 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x743 &  x746 &  x752 &  x755 &  x758 &  x761 &  x764 &  x773 &  x776 &  x779 &  x782 &  x788 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x839 &  x845 &  x848 &  x851 &  x857 &  x860 &  x863 &  x869 &  x872 &  x881 &  x884 &  x887 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x941 &  x944 &  x947 &  x950 &  x956 &  x959 &  x962 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1019 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1046 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1073 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1121 &  x1124 &  x1127 & ~x321 & ~x432 & ~x471 & ~x510 & ~x729;
assign c2280 =  x8 &  x11 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x56 &  x59 &  x62 &  x68 &  x77 &  x80 &  x86 &  x92 &  x101 &  x104 &  x107 &  x110 &  x116 &  x119 &  x122 &  x128 &  x131 &  x137 &  x140 &  x143 &  x146 &  x152 &  x155 &  x158 &  x164 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x197 &  x206 &  x209 &  x212 &  x218 &  x221 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x254 &  x257 &  x263 &  x266 &  x272 &  x278 &  x281 &  x284 &  x290 &  x296 &  x299 &  x302 &  x308 &  x311 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x365 &  x368 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x398 &  x401 &  x407 &  x413 &  x416 &  x422 &  x428 &  x431 &  x440 &  x443 &  x446 &  x449 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x476 &  x482 &  x491 &  x494 &  x497 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x539 &  x542 &  x547 &  x548 &  x551 &  x554 &  x557 &  x563 &  x575 &  x581 &  x584 &  x590 &  x593 &  x602 &  x605 &  x614 &  x620 &  x625 &  x626 &  x629 &  x632 &  x644 &  x647 &  x650 &  x662 &  x665 &  x668 &  x674 &  x680 &  x686 &  x692 &  x695 &  x698 &  x703 &  x704 &  x710 &  x713 &  x728 &  x737 &  x743 &  x746 &  x755 &  x761 &  x764 &  x767 &  x770 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x812 &  x815 &  x818 &  x821 &  x824 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x857 &  x860 &  x863 &  x866 &  x872 &  x875 &  x878 &  x881 &  x896 &  x902 &  x905 &  x908 &  x911 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x977 &  x980 &  x983 &  x986 &  x1001 &  x1004 &  x1007 &  x1016 &  x1022 &  x1025 &  x1037 &  x1046 &  x1055 &  x1058 &  x1061 &  x1073 &  x1076 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 & ~x441 & ~x519 & ~x534 & ~x558 & ~x669 & ~x708 & ~x744 & ~x792 & ~x861 & ~x939 & ~x978;
assign c2282 =  x1 &  x8 &  x14 &  x20 &  x23 &  x29 &  x32 &  x38 &  x41 &  x44 &  x53 &  x56 &  x59 &  x65 &  x80 &  x83 &  x86 &  x92 &  x95 &  x110 &  x128 &  x134 &  x140 &  x143 &  x149 &  x155 &  x158 &  x161 &  x167 &  x170 &  x173 &  x176 &  x182 &  x191 &  x197 &  x200 &  x206 &  x212 &  x221 &  x227 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x250 &  x251 &  x275 &  x281 &  x287 &  x296 &  x299 &  x308 &  x311 &  x323 &  x326 &  x328 &  x329 &  x335 &  x341 &  x353 &  x359 &  x365 &  x368 &  x383 &  x389 &  x395 &  x398 &  x419 &  x434 &  x437 &  x440 &  x443 &  x455 &  x458 &  x461 &  x464 &  x473 &  x475 &  x482 &  x503 &  x506 &  x515 &  x521 &  x527 &  x530 &  x533 &  x539 &  x554 &  x560 &  x572 &  x578 &  x581 &  x584 &  x596 &  x599 &  x602 &  x608 &  x614 &  x617 &  x620 &  x623 &  x629 &  x635 &  x638 &  x641 &  x653 &  x656 &  x659 &  x662 &  x665 &  x671 &  x674 &  x677 &  x683 &  x686 &  x689 &  x692 &  x698 &  x701 &  x703 &  x707 &  x713 &  x716 &  x722 &  x725 &  x728 &  x734 &  x743 &  x746 &  x749 &  x767 &  x770 &  x776 &  x779 &  x788 &  x791 &  x806 &  x812 &  x815 &  x820 &  x821 &  x824 &  x827 &  x830 &  x833 &  x839 &  x845 &  x848 &  x851 &  x857 &  x859 &  x860 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x890 &  x892 &  x898 &  x899 &  x905 &  x908 &  x911 &  x929 &  x931 &  x932 &  x935 &  x937 &  x938 &  x941 &  x947 &  x950 &  x952 &  x953 &  x956 &  x962 &  x968 &  x971 &  x980 &  x983 &  x986 &  x991 &  x995 &  x998 &  x1004 &  x1009 &  x1010 &  x1015 &  x1025 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1061 &  x1073 &  x1088 &  x1093 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1127 &  x1130 & ~x675 & ~x837 & ~x876 & ~x882 & ~x1077;
assign c2284 =  x2 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x242 &  x245 &  x248 &  x251 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x311 &  x317 &  x320 &  x323 &  x329 &  x332 &  x335 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x391 &  x392 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x434 &  x437 &  x440 &  x443 &  x449 &  x452 &  x455 &  x458 &  x461 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x584 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x640 &  x641 &  x644 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x710 &  x716 &  x719 &  x725 &  x728 &  x731 &  x734 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x757 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x842 &  x845 &  x848 &  x851 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x938 &  x941 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x983 &  x986 &  x989 &  x992 &  x998 &  x1001 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1129 &  x1130 & ~x261 & ~x435 & ~x663 & ~x705 & ~x744 & ~x975 & ~x1008 & ~x1014 & ~x1047 & ~x1053 & ~x1092 & ~x1125;
assign c2286 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x38 &  x41 &  x44 &  x47 &  x53 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x104 &  x107 &  x110 &  x113 &  x116 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x146 &  x149 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x218 &  x221 &  x227 &  x230 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x272 &  x275 &  x278 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x380 &  x383 &  x389 &  x395 &  x398 &  x401 &  x407 &  x410 &  x413 &  x416 &  x425 &  x428 &  x431 &  x437 &  x446 &  x449 &  x452 &  x455 &  x458 &  x464 &  x467 &  x473 &  x476 &  x479 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x514 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x563 &  x566 &  x572 &  x575 &  x578 &  x584 &  x587 &  x590 &  x593 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x638 &  x644 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x674 &  x677 &  x680 &  x686 &  x689 &  x695 &  x698 &  x701 &  x703 &  x704 &  x710 &  x719 &  x722 &  x725 &  x728 &  x731 &  x737 &  x740 &  x742 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x779 &  x781 &  x782 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x818 &  x820 &  x824 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x854 &  x859 &  x860 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x905 &  x911 &  x914 &  x917 &  x920 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x950 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x986 &  x989 &  x992 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1130 & ~x315 & ~x612 & ~x669 & ~x864 & ~x900 & ~x903 & ~x939 & ~x942 & ~x978 & ~x981;
assign c2288 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x56 &  x59 &  x62 &  x65 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x92 &  x95 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x170 &  x173 &  x176 &  x179 &  x182 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x233 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x356 &  x358 &  x359 &  x362 &  x371 &  x377 &  x380 &  x389 &  x392 &  x395 &  x397 &  x401 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x434 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x464 &  x467 &  x470 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x533 &  x539 &  x542 &  x551 &  x554 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x602 &  x614 &  x617 &  x620 &  x623 &  x626 &  x632 &  x635 &  x644 &  x647 &  x650 &  x653 &  x659 &  x662 &  x665 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x736 &  x737 &  x740 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x770 &  x773 &  x775 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x842 &  x845 &  x848 &  x851 &  x857 &  x860 &  x863 &  x869 &  x875 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x905 &  x908 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x959 &  x962 &  x965 &  x968 &  x977 &  x986 &  x989 &  x992 &  x995 &  x1007 &  x1016 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x273 & ~x558 & ~x636 & ~x753 & ~x900 & ~x939 & ~x978;
assign c2290 =  x2 &  x5 &  x8 &  x11 &  x17 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x83 &  x89 &  x92 &  x95 &  x101 &  x110 &  x113 &  x131 &  x134 &  x137 &  x140 &  x149 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x191 &  x194 &  x197 &  x203 &  x209 &  x218 &  x224 &  x227 &  x236 &  x239 &  x245 &  x251 &  x254 &  x257 &  x263 &  x266 &  x269 &  x272 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x305 &  x317 &  x323 &  x326 &  x329 &  x335 &  x341 &  x344 &  x350 &  x353 &  x356 &  x359 &  x362 &  x368 &  x371 &  x373 &  x374 &  x377 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x403 &  x404 &  x407 &  x410 &  x412 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x442 &  x446 &  x452 &  x458 &  x461 &  x464 &  x470 &  x473 &  x476 &  x491 &  x497 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x539 &  x542 &  x548 &  x551 &  x556 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x584 &  x587 &  x590 &  x596 &  x602 &  x605 &  x608 &  x617 &  x620 &  x623 &  x629 &  x638 &  x644 &  x647 &  x650 &  x653 &  x659 &  x668 &  x674 &  x677 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x722 &  x728 &  x731 &  x734 &  x737 &  x746 &  x752 &  x758 &  x761 &  x770 &  x773 &  x776 &  x788 &  x791 &  x794 &  x797 &  x800 &  x806 &  x818 &  x827 &  x836 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x872 &  x881 &  x884 &  x890 &  x893 &  x896 &  x899 &  x905 &  x908 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x938 &  x941 &  x944 &  x947 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x983 &  x992 &  x995 &  x998 &  x1001 &  x1013 &  x1019 &  x1025 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1103 &  x1106 &  x1109 &  x1124 & ~x693 & ~x768 & ~x786 & ~x807 & ~x942 & ~x1020 & ~x1056;
assign c2292 =  x8 &  x17 &  x20 &  x26 &  x29 &  x32 &  x53 &  x59 &  x65 &  x83 &  x86 &  x92 &  x104 &  x110 &  x122 &  x152 &  x170 &  x173 &  x176 &  x185 &  x200 &  x203 &  x206 &  x227 &  x236 &  x242 &  x278 &  x296 &  x302 &  x305 &  x310 &  x314 &  x317 &  x326 &  x349 &  x374 &  x388 &  x389 &  x407 &  x419 &  x434 &  x437 &  x440 &  x461 &  x470 &  x473 &  x476 &  x491 &  x494 &  x497 &  x509 &  x512 &  x527 &  x530 &  x554 &  x566 &  x584 &  x587 &  x608 &  x617 &  x647 &  x653 &  x656 &  x659 &  x668 &  x674 &  x710 &  x746 &  x767 &  x773 &  x779 &  x782 &  x788 &  x794 &  x797 &  x800 &  x803 &  x809 &  x815 &  x818 &  x830 &  x851 &  x860 &  x866 &  x911 &  x938 &  x941 &  x953 &  x956 &  x959 &  x965 &  x971 &  x986 &  x992 &  x1004 &  x1049 &  x1058 &  x1061 &  x1064 &  x1076 &  x1088 &  x1112 &  x1124 &  x1127 & ~x579 & ~x618 & ~x657 & ~x658 & ~x735 & ~x882 & ~x909 & ~x948;
assign c2294 =  x2 &  x5 &  x11 &  x14 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x47 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x77 &  x83 &  x86 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x146 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x206 &  x209 &  x212 &  x215 &  x217 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x358 &  x359 &  x362 &  x365 &  x371 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x401 &  x407 &  x410 &  x419 &  x422 &  x428 &  x431 &  x434 &  x437 &  x443 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x629 &  x635 &  x641 &  x644 &  x647 &  x650 &  x662 &  x665 &  x668 &  x671 &  x674 &  x680 &  x682 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x758 &  x767 &  x770 &  x773 &  x776 &  x779 &  x781 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x820 &  x821 &  x824 &  x827 &  x830 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x853 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x874 &  x875 &  x878 &  x881 &  x890 &  x892 &  x893 &  x896 &  x898 &  x899 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x931 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x952 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x983 &  x986 &  x989 &  x991 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1009 &  x1010 &  x1013 &  x1016 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x273 & ~x312 & ~x882;
assign c2296 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x53 &  x56 &  x62 &  x65 &  x68 &  x71 &  x80 &  x83 &  x92 &  x95 &  x98 &  x104 &  x107 &  x110 &  x113 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x139 &  x140 &  x143 &  x146 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x176 &  x178 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x209 &  x212 &  x217 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x287 &  x290 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x358 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x395 &  x397 &  x398 &  x400 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x436 &  x437 &  x439 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x472 &  x473 &  x476 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x511 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x547 &  x548 &  x550 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x614 &  x617 &  x620 &  x625 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x710 &  x713 &  x716 &  x719 &  x725 &  x728 &  x731 &  x734 &  x737 &  x742 &  x743 &  x746 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x776 &  x779 &  x782 &  x785 &  x788 &  x794 &  x797 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x845 &  x854 &  x857 &  x860 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x935 &  x941 &  x944 &  x947 &  x950 &  x953 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x861 & ~x978;
assign c2298 =  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x47 &  x50 &  x53 &  x56 &  x59 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x104 &  x107 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x155 &  x160 &  x167 &  x173 &  x179 &  x182 &  x196 &  x203 &  x209 &  x212 &  x221 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x260 &  x263 &  x269 &  x274 &  x278 &  x281 &  x284 &  x287 &  x296 &  x299 &  x311 &  x313 &  x326 &  x329 &  x332 &  x335 &  x341 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x449 &  x452 &  x455 &  x458 &  x461 &  x473 &  x488 &  x491 &  x494 &  x503 &  x512 &  x515 &  x521 &  x527 &  x530 &  x539 &  x542 &  x545 &  x551 &  x554 &  x557 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x593 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x662 &  x665 &  x671 &  x674 &  x680 &  x683 &  x686 &  x701 &  x704 &  x707 &  x710 &  x722 &  x725 &  x731 &  x734 &  x743 &  x749 &  x752 &  x755 &  x758 &  x767 &  x770 &  x776 &  x779 &  x791 &  x797 &  x800 &  x803 &  x812 &  x818 &  x821 &  x833 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x890 &  x896 &  x902 &  x905 &  x908 &  x911 &  x914 &  x920 &  x923 &  x926 &  x932 &  x935 &  x941 &  x950 &  x953 &  x962 &  x965 &  x968 &  x971 &  x974 &  x980 &  x983 &  x986 &  x992 &  x998 &  x1001 &  x1007 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1046 &  x1049 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x246 & ~x285 & ~x324 & ~x357 & ~x363 & ~x402 & ~x441 & ~x453 & ~x480 & ~x588 & ~x627 & ~x628 & ~x666 & ~x705 & ~x744 & ~x780 & ~x858 & ~x897 & ~x936 & ~x975 & ~x1014;
assign c21 =  x37 &  x76 &  x702 &  x932 & ~x510 & ~x891;
assign c23 =  x5 &  x68 &  x86 &  x92 &  x98 &  x101 &  x107 &  x167 &  x290 &  x296 &  x308 &  x344 &  x353 &  x401 &  x419 &  x431 &  x515 &  x539 &  x545 &  x550 &  x674 &  x719 &  x755 &  x770 &  x911 &  x929 &  x977 &  x986 &  x989 &  x1001 &  x1022 &  x1061 &  x1067 &  x1073 &  x1094 & ~x561 & ~x723 & ~x735 & ~x762 & ~x774 & ~x775;
assign c25 =  x5 &  x17 &  x23 &  x26 &  x41 &  x56 &  x71 &  x80 &  x83 &  x110 &  x122 &  x137 &  x176 &  x221 &  x224 &  x233 &  x239 &  x244 &  x263 &  x266 &  x275 &  x296 &  x305 &  x308 &  x323 &  x335 &  x395 &  x407 &  x413 &  x422 &  x452 &  x455 &  x473 &  x527 &  x554 &  x572 &  x581 &  x596 &  x611 &  x623 &  x629 &  x671 &  x680 &  x691 &  x692 &  x731 &  x755 &  x764 &  x767 &  x779 &  x782 &  x794 &  x806 &  x833 &  x845 &  x848 &  x860 &  x866 &  x878 &  x881 &  x893 &  x896 &  x956 &  x958 &  x983 &  x992 &  x998 &  x1004 &  x1031 &  x1049 &  x1088 &  x1115 & ~x750 & ~x816 & ~x984 & ~x1062;
assign c27 =  x552 &  x591 &  x638 & ~x447 & ~x486 & ~x936 & ~x1092;
assign c29 =  x550 &  x867 & ~x582 & ~x771;
assign c211 =  x337 &  x421 &  x460 &  x551 &  x703 &  x937 &  x989 & ~x1086;
assign c213 =  x2 &  x38 &  x71 &  x440 &  x506 &  x512 &  x590 &  x659 &  x698 &  x784 &  x848 &  x854 &  x940 &  x1001 &  x1025 &  x1070 &  x1100 & ~x441 & ~x519 & ~x600 & ~x636;
assign c215 =  x197 &  x223 &  x481 &  x703 &  x731 &  x1021 & ~x393 & ~x771 & ~x915;
assign c217 =  x455 &  x472 & ~x405 & ~x820 & ~x1014 & ~x1017;
assign c219 =  x50 &  x248 &  x312 &  x410 &  x449 &  x686 & ~x126 & ~x165 & ~x900 & ~x1095;
assign c221 =  x8 &  x11 &  x14 &  x29 &  x41 &  x47 &  x80 &  x92 &  x98 &  x101 &  x113 &  x122 &  x137 &  x143 &  x152 &  x188 &  x200 &  x203 &  x206 &  x212 &  x230 &  x239 &  x257 &  x260 &  x266 &  x284 &  x302 &  x305 &  x314 &  x320 &  x323 &  x344 &  x371 &  x377 &  x404 &  x407 &  x422 &  x428 &  x437 &  x440 &  x443 &  x452 &  x458 &  x461 &  x467 &  x476 &  x479 &  x488 &  x494 &  x500 &  x512 &  x518 &  x536 &  x554 &  x557 &  x560 &  x575 &  x590 &  x614 &  x620 &  x626 &  x629 &  x632 &  x647 &  x650 &  x656 &  x671 &  x674 &  x692 &  x704 &  x706 &  x710 &  x716 &  x728 &  x745 &  x746 &  x755 &  x758 &  x764 &  x785 &  x788 &  x803 &  x818 &  x824 &  x836 &  x848 &  x862 &  x866 &  x869 &  x878 &  x884 &  x890 &  x896 &  x905 &  x911 &  x917 &  x926 &  x938 &  x944 &  x979 &  x992 &  x1001 &  x1004 &  x1018 &  x1028 &  x1031 &  x1043 &  x1049 &  x1067 &  x1079 &  x1088 &  x1112 &  x1115 & ~x597 & ~x636 & ~x639;
assign c223 =  x2 &  x17 &  x65 &  x296 &  x317 &  x320 &  x359 &  x445 &  x560 &  x940 &  x1004 &  x1007 &  x1010 & ~x78 & ~x315 & ~x795 & ~x813;
assign c225 =  x37 &  x236 &  x292 &  x437 &  x803 & ~x159 & ~x852;
assign c227 =  x2 &  x59 &  x68 &  x71 &  x86 &  x101 &  x113 &  x176 &  x188 &  x194 &  x233 &  x245 &  x251 &  x263 &  x311 &  x341 &  x347 &  x362 &  x389 &  x419 &  x422 &  x467 &  x485 &  x497 &  x511 &  x530 &  x533 &  x548 &  x584 &  x617 &  x626 &  x632 &  x647 &  x653 &  x677 &  x680 &  x683 &  x707 &  x761 &  x776 &  x794 &  x811 &  x845 &  x881 &  x893 &  x896 &  x929 &  x944 &  x953 &  x962 &  x968 &  x1034 &  x1039 &  x1046 &  x1097 &  x1115 & ~x858 & ~x936;
assign c229 =  x152 &  x197 &  x289 &  x596 &  x755 &  x901 &  x937 &  x1057 & ~x120 & ~x159 & ~x510 & ~x903;
assign c231 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x29 &  x38 &  x41 &  x74 &  x80 &  x110 &  x119 &  x128 &  x131 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x173 &  x176 &  x194 &  x197 &  x233 &  x242 &  x254 &  x269 &  x278 &  x287 &  x293 &  x299 &  x305 &  x323 &  x326 &  x329 &  x335 &  x341 &  x344 &  x347 &  x362 &  x368 &  x392 &  x398 &  x404 &  x416 &  x428 &  x430 &  x434 &  x437 &  x440 &  x455 &  x458 &  x473 &  x479 &  x482 &  x488 &  x491 &  x503 &  x508 &  x539 &  x547 &  x557 &  x563 &  x586 &  x589 &  x614 &  x626 &  x628 &  x632 &  x635 &  x647 &  x650 &  x662 &  x677 &  x683 &  x686 &  x695 &  x704 &  x706 &  x710 &  x712 &  x713 &  x743 &  x746 &  x751 &  x770 &  x773 &  x776 &  x782 &  x800 &  x809 &  x812 &  x821 &  x842 &  x866 &  x875 &  x884 &  x887 &  x893 &  x896 &  x902 &  x917 &  x923 &  x932 &  x938 &  x941 &  x953 &  x962 &  x995 &  x998 &  x1004 &  x1010 &  x1022 &  x1025 &  x1028 &  x1040 &  x1067 &  x1073 &  x1076 &  x1094 &  x1100 &  x1112 &  x1118 &  x1121 &  x1124 &  x1130 & ~x474 & ~x513 & ~x552;
assign c233 =  x320 &  x432 &  x550 & ~x522 & ~x624 & ~x858 & ~x984;
assign c235 =  x29 &  x50 &  x53 &  x59 &  x95 &  x221 &  x398 &  x419 &  x497 &  x514 &  x553 &  x629 &  x662 &  x677 &  x685 &  x731 &  x785 &  x791 &  x839 &  x872 &  x917 &  x980 &  x1010 &  x1109 &  x1127 &  x1130 & ~x84 & ~x162 & ~x663 & ~x822 & ~x942 & ~x981;
assign c237 =  x167 &  x206 &  x380 &  x401 &  x473 &  x620 &  x638 &  x652 &  x736 &  x812 &  x842 &  x958 &  x965 & ~x660 & ~x699 & ~x1068;
assign c239 = ~x316 & ~x708;
assign c241 =  x113 &  x122 &  x164 &  x167 &  x281 &  x296 &  x317 &  x335 &  x416 &  x431 &  x472 &  x557 &  x631 &  x632 &  x662 &  x670 &  x683 &  x692 &  x821 &  x863 &  x1013 &  x1064 &  x1085 &  x1097 &  x1118 &  x1121 & ~x279 & ~x858 & ~x897 & ~x1077;
assign c243 =  x77 &  x89 &  x116 &  x203 &  x221 &  x245 &  x257 &  x287 &  x314 &  x374 &  x440 &  x452 &  x476 &  x494 &  x545 &  x644 &  x646 &  x650 &  x686 &  x713 &  x731 &  x824 &  x962 &  x980 &  x992 &  x1109 & ~x45 & ~x331 & ~x369 & ~x819;
assign c245 = ~x709;
assign c247 =  x741 &  x867 & ~x390 & ~x709;
assign c249 =  x513 &  x535 & ~x348 & ~x858;
assign c251 =  x686 &  x853 &  x859 &  x885 & ~x201 & ~x1056;
assign c253 =  x2 &  x8 &  x14 &  x32 &  x37 &  x53 &  x59 &  x74 &  x80 &  x140 &  x146 &  x167 &  x176 &  x179 &  x194 &  x200 &  x203 &  x218 &  x224 &  x226 &  x227 &  x233 &  x242 &  x248 &  x251 &  x269 &  x302 &  x308 &  x310 &  x311 &  x350 &  x359 &  x392 &  x398 &  x401 &  x407 &  x416 &  x425 &  x464 &  x476 &  x488 &  x503 &  x506 &  x536 &  x542 &  x566 &  x578 &  x581 &  x584 &  x587 &  x596 &  x605 &  x608 &  x632 &  x638 &  x641 &  x644 &  x674 &  x680 &  x689 &  x695 &  x707 &  x713 &  x716 &  x722 &  x737 &  x758 &  x767 &  x770 &  x776 &  x797 &  x821 &  x824 &  x830 &  x842 &  x845 &  x854 &  x860 &  x863 &  x875 &  x884 &  x893 &  x905 &  x914 &  x935 &  x944 &  x950 &  x962 &  x971 &  x986 &  x1013 &  x1019 &  x1028 &  x1058 &  x1061 &  x1067 &  x1085 &  x1088 &  x1106 &  x1109 &  x1130 & ~x81 & ~x240 & ~x513 & ~x552 & ~x591;
assign c255 =  x17 &  x134 &  x143 &  x170 &  x211 &  x524 &  x536 &  x706 &  x746 &  x791 &  x857 &  x862 &  x914 &  x938 &  x1001 &  x1013 &  x1096 & ~x237 & ~x276 & ~x816;
assign c257 =  x17 &  x29 &  x47 &  x71 &  x155 &  x218 &  x248 &  x254 &  x296 &  x311 &  x340 &  x347 &  x374 &  x389 &  x485 &  x547 &  x557 &  x602 &  x683 &  x728 &  x731 &  x878 &  x881 &  x977 &  x1043 &  x1052 & ~x513 & ~x693 & ~x765 & ~x777 & ~x816 & ~x1065;
assign c259 =  x196 &  x206 &  x242 &  x248 &  x458 &  x670 &  x844 &  x854 &  x1103 &  x1124 & ~x124 & ~x828 & ~x1098;
assign c261 =  x134 &  x140 &  x148 &  x188 &  x227 &  x290 &  x323 &  x407 &  x413 &  x481 &  x484 &  x485 &  x488 &  x560 &  x665 &  x683 &  x767 &  x776 &  x800 &  x836 &  x859 &  x898 &  x904 &  x962 &  x998 &  x1010 &  x1054 &  x1058 &  x1120 &  x1130 & ~x588;
assign c263 =  x76 &  x445 &  x646 &  x808 & ~x738;
assign c265 =  x110 &  x419 &  x446 &  x626 &  x689 &  x823 &  x862 &  x875 & ~x237 & ~x594 & ~x747 & ~x981;
assign c267 =  x485 &  x508 &  x547 &  x698 &  x845 &  x905 &  x926 &  x995 &  x1028 & ~x159 & ~x399 & ~x400 & ~x615;
assign c269 =  x64 &  x170 &  x175 &  x226 &  x253 &  x269 &  x419 &  x425 &  x467 &  x491 &  x569 &  x641 &  x659 &  x728 &  x742 &  x866 &  x875 &  x953 & ~x411 & ~x816 & ~x849;
assign c271 =  x550 &  x687 & ~x861;
assign c273 =  x550 & ~x601 & ~x774 & ~x858;
assign c275 =  x65 &  x140 &  x325 &  x380 &  x404 &  x434 &  x479 &  x638 &  x692 &  x869 &  x926 &  x938 &  x1060 &  x1099 &  x1124 & ~x234 & ~x354 & ~x393 & ~x798;
assign c277 =  x5 &  x29 &  x44 &  x47 &  x53 &  x137 &  x188 &  x197 &  x242 &  x245 &  x260 &  x299 &  x359 &  x440 &  x445 &  x452 &  x455 &  x497 &  x512 &  x527 &  x585 &  x587 &  x593 &  x596 &  x644 &  x647 &  x659 &  x662 &  x686 &  x701 &  x710 &  x716 &  x722 &  x731 &  x755 &  x764 &  x781 &  x791 &  x806 &  x809 &  x836 &  x884 &  x902 &  x905 &  x926 &  x941 &  x947 &  x1025 &  x1112 & ~x474 & ~x513 & ~x615 & ~x870;
assign c279 =  x11 &  x47 &  x56 &  x79 &  x92 &  x122 &  x146 &  x167 &  x227 &  x278 &  x281 &  x296 &  x323 &  x344 &  x389 &  x425 &  x476 &  x488 &  x491 &  x530 &  x572 &  x590 &  x593 &  x608 &  x629 &  x671 &  x674 &  x710 &  x727 &  x737 &  x791 &  x811 &  x812 &  x860 &  x922 &  x926 &  x977 &  x980 &  x995 &  x998 &  x1019 &  x1037 &  x1043 &  x1058 &  x1064 &  x1078 &  x1127 & ~x102 & ~x162 & ~x942;
assign c281 =  x352 &  x510 & ~x240 & ~x663;
assign c283 =  x26 &  x32 &  x47 &  x86 &  x122 &  x131 &  x143 &  x170 &  x203 &  x251 &  x302 &  x326 &  x362 &  x368 &  x413 &  x455 &  x458 &  x470 &  x479 &  x644 &  x674 &  x683 &  x743 &  x788 &  x806 &  x818 &  x824 &  x905 &  x914 &  x932 &  x956 &  x992 &  x1001 &  x1013 &  x1064 & ~x3 & ~x132 & ~x217 & ~x462;
assign c285 =  x697 &  x724 &  x808 & ~x705 & ~x828 & ~x855 & ~x1056;
assign c287 =  x14 &  x194 &  x302 &  x404 &  x667 &  x862 &  x1094 & ~x237 & ~x354 & ~x597 & ~x636;
assign c289 =  x23 &  x91 &  x125 &  x173 &  x398 &  x407 &  x419 &  x671 &  x747 &  x908 &  x926 &  x1031 & ~x411 & ~x1092;
assign c291 =  x8 &  x20 &  x29 &  x38 &  x47 &  x53 &  x56 &  x71 &  x80 &  x83 &  x89 &  x95 &  x104 &  x113 &  x125 &  x128 &  x140 &  x143 &  x152 &  x155 &  x158 &  x164 &  x176 &  x185 &  x191 &  x212 &  x215 &  x221 &  x251 &  x254 &  x260 &  x269 &  x284 &  x299 &  x305 &  x311 &  x329 &  x332 &  x344 &  x347 &  x353 &  x359 &  x362 &  x377 &  x392 &  x407 &  x422 &  x425 &  x428 &  x431 &  x449 &  x452 &  x470 &  x473 &  x500 &  x509 &  x542 &  x551 &  x554 &  x563 &  x566 &  x569 &  x587 &  x605 &  x653 &  x668 &  x689 &  x692 &  x698 &  x701 &  x728 &  x734 &  x737 &  x785 &  x812 &  x818 &  x833 &  x842 &  x857 &  x860 &  x862 &  x869 &  x872 &  x875 &  x881 &  x890 &  x923 &  x929 &  x932 &  x938 &  x953 &  x962 &  x974 &  x1007 &  x1022 &  x1031 &  x1040 &  x1049 &  x1058 &  x1061 &  x1067 &  x1085 &  x1097 &  x1112 & ~x30 & ~x213 & ~x516 & ~x555 & ~x597 & ~x942;
assign c293 =  x71 &  x134 &  x140 &  x218 &  x248 &  x353 &  x394 &  x401 &  x434 &  x500 &  x648 &  x687 &  x695 &  x748 &  x785 &  x824 &  x833 &  x871 &  x944 &  x1079 &  x1082 & ~x822;
assign c295 =  x748 &  x967 &  x1006 & ~x42 & ~x486 & ~x525;
assign c297 =  x1096 & ~x871 & ~x912;
assign c299 =  x35 &  x47 &  x83 &  x104 &  x107 &  x113 &  x146 &  x155 &  x200 &  x212 &  x236 &  x239 &  x254 &  x269 &  x287 &  x305 &  x311 &  x323 &  x328 &  x395 &  x398 &  x431 &  x443 &  x446 &  x461 &  x464 &  x512 &  x539 &  x542 &  x545 &  x563 &  x590 &  x638 &  x647 &  x656 &  x683 &  x689 &  x692 &  x695 &  x701 &  x770 &  x818 &  x824 &  x833 &  x890 &  x902 &  x917 &  x931 &  x932 &  x941 &  x947 &  x962 &  x1004 &  x1013 &  x1019 &  x1055 &  x1058 &  x1106 & ~x396 & ~x435 & ~x474 & ~x816 & ~x972 & ~x1044 & ~x1104;
assign c2101 =  x288 &  x1074 &  x1113 & ~x738;
assign c2103 =  x742 &  x790 &  x1067 & ~x156 & ~x799;
assign c2105 =  x10 &  x23 &  x28 &  x86 &  x101 &  x113 &  x119 &  x134 &  x167 &  x172 &  x188 &  x215 &  x242 &  x251 &  x347 &  x359 &  x386 &  x428 &  x446 &  x449 &  x452 &  x506 &  x557 &  x611 &  x656 &  x719 &  x728 &  x773 &  x791 &  x794 &  x809 &  x812 &  x836 &  x851 &  x890 &  x899 &  x902 &  x920 &  x929 &  x958 &  x959 &  x968 &  x997 &  x1007 &  x1091 &  x1124 & ~x582 & ~x816;
assign c2107 =  x421 &  x616 &  x898 &  x1035 &  x1113;
assign c2109 =  x25 &  x304 &  x305 &  x365 &  x674 &  x710 &  x983 &  x998 &  x1016 & ~x399 & ~x1092;
assign c2111 =  x5 &  x17 &  x20 &  x23 &  x32 &  x47 &  x62 &  x65 &  x68 &  x83 &  x89 &  x95 &  x116 &  x143 &  x158 &  x194 &  x197 &  x212 &  x215 &  x218 &  x236 &  x251 &  x260 &  x263 &  x272 &  x275 &  x287 &  x299 &  x302 &  x308 &  x335 &  x353 &  x359 &  x362 &  x365 &  x371 &  x374 &  x377 &  x407 &  x413 &  x422 &  x425 &  x428 &  x437 &  x440 &  x470 &  x476 &  x485 &  x491 &  x500 &  x503 &  x518 &  x536 &  x542 &  x548 &  x551 &  x554 &  x557 &  x569 &  x578 &  x593 &  x596 &  x602 &  x611 &  x623 &  x629 &  x632 &  x635 &  x644 &  x647 &  x662 &  x665 &  x671 &  x677 &  x689 &  x733 &  x740 &  x758 &  x766 &  x767 &  x770 &  x776 &  x785 &  x805 &  x815 &  x821 &  x844 &  x845 &  x860 &  x881 &  x908 &  x917 &  x920 &  x971 &  x977 &  x986 &  x995 &  x998 &  x1013 &  x1022 &  x1052 &  x1070 &  x1091 &  x1094 &  x1097 &  x1103 &  x1115 &  x1118 &  x1127 & ~x447 & ~x486 & ~x828 & ~x1020 & ~x1059;
assign c2113 =  x2 &  x25 &  x50 &  x53 &  x80 &  x107 &  x146 &  x179 &  x218 &  x224 &  x233 &  x242 &  x257 &  x266 &  x278 &  x281 &  x296 &  x329 &  x347 &  x350 &  x356 &  x362 &  x401 &  x413 &  x431 &  x452 &  x455 &  x470 &  x482 &  x494 &  x500 &  x509 &  x527 &  x536 &  x551 &  x560 &  x566 &  x572 &  x608 &  x635 &  x638 &  x647 &  x668 &  x671 &  x683 &  x698 &  x722 &  x764 &  x770 &  x782 &  x788 &  x791 &  x794 &  x803 &  x806 &  x812 &  x821 &  x824 &  x845 &  x851 &  x872 &  x878 &  x884 &  x890 &  x893 &  x914 &  x920 &  x932 &  x956 &  x962 &  x965 &  x977 &  x980 &  x995 &  x1001 &  x1004 &  x1010 &  x1025 &  x1031 &  x1040 &  x1076 &  x1084 &  x1094 &  x1097 &  x1100 &  x1115 & ~x240 & ~x357 & ~x462;
assign c2115 =  x80 &  x188 &  x311 &  x368 &  x392 &  x545 &  x671 &  x869 &  x920 &  x1061 &  x1067 & ~x3 & ~x162 & ~x174 & ~x258 & ~x318 & ~x1023 & ~x1101;
assign c2117 =  x62 &  x95 &  x107 &  x113 &  x215 &  x245 &  x257 &  x299 &  x314 &  x395 &  x416 &  x476 &  x635 &  x680 &  x764 &  x866 &  x881 &  x908 &  x932 &  x941 &  x974 &  x983 &  x992 &  x1010 &  x1046 &  x1078 &  x1088 & ~x30 & ~x267 & ~x423 & ~x915;
assign c2119 =  x786 & ~x582 & ~x799;
assign c2121 =  x10 &  x82 &  x88 &  x98 &  x149 &  x236 &  x287 &  x350 &  x413 &  x461 &  x521 &  x557 &  x701 &  x728 &  x842 &  x851 &  x958 &  x983 &  x998 &  x1061 &  x1067 & ~x699 & ~x816 & ~x933;
assign c2123 =  x5 &  x14 &  x38 &  x74 &  x86 &  x95 &  x104 &  x125 &  x155 &  x203 &  x224 &  x233 &  x254 &  x260 &  x269 &  x278 &  x305 &  x314 &  x317 &  x335 &  x341 &  x347 &  x362 &  x383 &  x397 &  x410 &  x431 &  x434 &  x443 &  x446 &  x449 &  x452 &  x461 &  x488 &  x506 &  x515 &  x539 &  x545 &  x566 &  x635 &  x650 &  x656 &  x665 &  x668 &  x680 &  x683 &  x686 &  x692 &  x698 &  x707 &  x731 &  x734 &  x755 &  x758 &  x785 &  x794 &  x803 &  x818 &  x824 &  x827 &  x851 &  x872 &  x887 &  x902 &  x917 &  x926 &  x950 &  x959 &  x971 &  x995 &  x998 &  x1004 &  x1019 &  x1025 &  x1034 &  x1046 &  x1061 &  x1064 &  x1070 &  x1091 &  x1115 &  x1127 &  x1130 & ~x90 & ~x333 & ~x390 & ~x477 & ~x930;
assign c2125 =  x226 &  x702 &  x741 & ~x471 & ~x474 & ~x510;
assign c2127 =  x445 &  x901 &  x906 &  x940;
assign c2129 =  x861 & ~x709;
assign c2131 =  x2 &  x8 &  x11 &  x14 &  x17 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x56 &  x62 &  x65 &  x68 &  x74 &  x80 &  x86 &  x92 &  x95 &  x98 &  x104 &  x110 &  x122 &  x125 &  x128 &  x134 &  x140 &  x143 &  x146 &  x149 &  x155 &  x164 &  x167 &  x173 &  x176 &  x179 &  x182 &  x206 &  x215 &  x221 &  x224 &  x230 &  x242 &  x245 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x274 &  x281 &  x284 &  x287 &  x290 &  x302 &  x305 &  x313 &  x314 &  x329 &  x332 &  x335 &  x341 &  x344 &  x350 &  x352 &  x353 &  x359 &  x368 &  x371 &  x374 &  x377 &  x392 &  x395 &  x401 &  x404 &  x407 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x433 &  x434 &  x440 &  x443 &  x446 &  x449 &  x455 &  x461 &  x470 &  x473 &  x479 &  x482 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x509 &  x511 &  x512 &  x524 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x560 &  x590 &  x593 &  x596 &  x605 &  x608 &  x611 &  x614 &  x620 &  x632 &  x634 &  x635 &  x638 &  x641 &  x644 &  x650 &  x656 &  x659 &  x662 &  x677 &  x689 &  x695 &  x704 &  x707 &  x716 &  x737 &  x740 &  x743 &  x752 &  x758 &  x767 &  x776 &  x782 &  x785 &  x794 &  x809 &  x815 &  x836 &  x839 &  x842 &  x848 &  x851 &  x860 &  x863 &  x869 &  x881 &  x884 &  x887 &  x890 &  x896 &  x899 &  x902 &  x905 &  x911 &  x917 &  x920 &  x923 &  x926 &  x929 &  x935 &  x941 &  x944 &  x953 &  x965 &  x971 &  x983 &  x986 &  x992 &  x998 &  x1004 &  x1007 &  x1013 &  x1019 &  x1031 &  x1040 &  x1049 &  x1055 &  x1067 &  x1073 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1115 &  x1118 &  x1121 &  x1127 & ~x483 & ~x741 & ~x780 & ~x819 & ~x858;
assign c2133 =  x394 &  x709 &  x811 &  x895 &  x1000 &  x1033 &  x1051;
assign c2135 =  x176 &  x185 &  x226 &  x628 &  x875 &  x988 & ~x477 & ~x963;
assign c2137 =  x909 & ~x775 & ~x892;
assign c2139 =  x407 &  x670 &  x766 &  x811 &  x910 & ~x333 & ~x334 & ~x342;
assign c2141 =  x77 &  x86 &  x158 &  x182 &  x203 &  x215 &  x293 &  x317 &  x323 &  x329 &  x395 &  x407 &  x524 &  x602 &  x611 &  x742 &  x781 &  x803 &  x818 &  x848 &  x863 &  x914 &  x935 &  x943 &  x962 &  x982 &  x995 &  x1004 &  x1010 &  x1031 &  x1055 &  x1112 & ~x237 & ~x916 & ~x954;
assign c2143 =  x742 &  x1020 & ~x915;
assign c2145 =  x11 &  x29 &  x38 &  x44 &  x65 &  x68 &  x74 &  x86 &  x89 &  x92 &  x95 &  x116 &  x119 &  x131 &  x134 &  x137 &  x158 &  x164 &  x167 &  x170 &  x176 &  x182 &  x188 &  x191 &  x194 &  x197 &  x203 &  x206 &  x209 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x251 &  x254 &  x263 &  x281 &  x287 &  x290 &  x302 &  x305 &  x308 &  x320 &  x332 &  x338 &  x344 &  x347 &  x359 &  x362 &  x365 &  x374 &  x380 &  x383 &  x386 &  x389 &  x392 &  x398 &  x404 &  x410 &  x419 &  x425 &  x446 &  x452 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x494 &  x497 &  x506 &  x515 &  x518 &  x521 &  x524 &  x527 &  x533 &  x557 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x593 &  x596 &  x602 &  x611 &  x617 &  x623 &  x626 &  x635 &  x638 &  x641 &  x650 &  x653 &  x671 &  x674 &  x677 &  x686 &  x692 &  x701 &  x704 &  x710 &  x719 &  x722 &  x728 &  x731 &  x742 &  x743 &  x746 &  x749 &  x752 &  x761 &  x764 &  x773 &  x776 &  x779 &  x781 &  x785 &  x788 &  x797 &  x815 &  x823 &  x827 &  x851 &  x860 &  x863 &  x866 &  x881 &  x887 &  x899 &  x901 &  x902 &  x911 &  x917 &  x920 &  x923 &  x926 &  x937 &  x940 &  x950 &  x953 &  x968 &  x971 &  x974 &  x980 &  x983 &  x989 &  x992 &  x995 &  x1007 &  x1010 &  x1013 &  x1016 &  x1018 &  x1019 &  x1025 &  x1031 &  x1037 &  x1040 &  x1049 &  x1055 &  x1058 &  x1061 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1100 &  x1103 &  x1109 &  x1118 &  x1124 &  x1130 & ~x510 & ~x597 & ~x636;
assign c2147 =  x70 &  x148 &  x753 &  x925 &  x964;
assign c2149 =  x103 &  x266 & ~x198 & ~x240 & ~x397;
assign c2151 =  x23 &  x32 &  x35 &  x47 &  x68 &  x98 &  x164 &  x185 &  x203 &  x206 &  x221 &  x233 &  x278 &  x329 &  x332 &  x350 &  x416 &  x419 &  x472 &  x473 &  x488 &  x497 &  x500 &  x527 &  x536 &  x550 &  x566 &  x581 &  x626 &  x668 &  x674 &  x695 &  x704 &  x707 &  x713 &  x719 &  x731 &  x746 &  x755 &  x767 &  x803 &  x851 &  x854 &  x860 &  x869 &  x878 &  x902 &  x908 &  x910 &  x950 &  x986 &  x995 &  x1000 &  x1025 &  x1052 &  x1067 &  x1091 &  x1112 & ~x1008 & ~x1014;
assign c2153 =  x14 &  x23 &  x35 &  x44 &  x62 &  x89 &  x92 &  x134 &  x137 &  x158 &  x176 &  x179 &  x206 &  x212 &  x221 &  x242 &  x251 &  x260 &  x278 &  x290 &  x302 &  x313 &  x344 &  x389 &  x419 &  x422 &  x443 &  x464 &  x467 &  x476 &  x503 &  x509 &  x536 &  x545 &  x551 &  x578 &  x593 &  x596 &  x605 &  x608 &  x611 &  x620 &  x635 &  x653 &  x659 &  x665 &  x670 &  x674 &  x685 &  x686 &  x707 &  x710 &  x713 &  x722 &  x728 &  x731 &  x743 &  x755 &  x761 &  x767 &  x787 &  x800 &  x827 &  x836 &  x848 &  x860 &  x872 &  x881 &  x899 &  x926 &  x929 &  x938 &  x941 &  x947 &  x950 &  x971 &  x974 &  x1013 &  x1019 &  x1022 &  x1025 &  x1076 &  x1088 &  x1118 &  x1124 & ~x447 & ~x663 & ~x741 & ~x819 & ~x1104;
assign c2155 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x155 &  x158 &  x164 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x239 &  x242 &  x248 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x278 &  x281 &  x284 &  x287 &  x290 &  x296 &  x305 &  x308 &  x311 &  x317 &  x320 &  x323 &  x326 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x365 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x398 &  x401 &  x407 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x455 &  x458 &  x461 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x524 &  x527 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x632 &  x635 &  x638 &  x641 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x734 &  x736 &  x740 &  x743 &  x746 &  x748 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x775 &  x776 &  x785 &  x787 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x896 &  x899 &  x902 &  x905 &  x911 &  x914 &  x917 &  x926 &  x929 &  x932 &  x935 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x961 &  x962 &  x964 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1000 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1030 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x6 & ~x45;
assign c2157 =  x319 &  x337 &  x652 &  x692 &  x806 &  x1010 &  x1085 & ~x393 & ~x816 & ~x1050;
assign c2159 =  x858 &  x1017 &  x1056 & ~x1083;
assign c2161 =  x56 &  x80 &  x113 &  x146 &  x395 &  x407 &  x443 &  x533 &  x545 &  x610 &  x616 &  x680 &  x688 &  x755 &  x761 &  x814 &  x967 &  x1088 &  x1109 &  x1118 & ~x45 & ~x123;
assign c2163 =  x275 &  x382 &  x431 &  x665 &  x683 & ~x42 & ~x553 & ~x654;
assign c2165 =  x290 &  x727 &  x803 & ~x3 & ~x213 & ~x486 & ~x912 & ~x1029;
assign c2167 =  x20 &  x230 &  x299 &  x407 &  x535 &  x601 &  x815 & ~x672 & ~x829 & ~x1089;
assign c2169 =  x2 &  x29 &  x35 &  x41 &  x62 &  x71 &  x117 &  x118 &  x125 &  x140 &  x157 &  x179 &  x197 &  x209 &  x224 &  x239 &  x242 &  x257 &  x263 &  x277 &  x284 &  x316 &  x323 &  x347 &  x355 &  x377 &  x389 &  x394 &  x395 &  x398 &  x419 &  x455 &  x461 &  x464 &  x472 &  x482 &  x497 &  x521 &  x533 &  x539 &  x563 &  x569 &  x584 &  x587 &  x590 &  x596 &  x608 &  x629 &  x686 &  x695 &  x701 &  x728 &  x752 &  x788 &  x794 &  x797 &  x800 &  x809 &  x815 &  x818 &  x824 &  x827 &  x836 &  x842 &  x854 &  x869 &  x878 &  x893 &  x896 &  x905 &  x911 &  x932 &  x938 &  x947 &  x956 &  x965 &  x968 &  x1001 &  x1004 &  x1022 &  x1031 &  x1037 &  x1040 &  x1049 &  x1055 &  x1070 &  x1073 &  x1100 &  x1112 &  x1130 & ~x741 & ~x780 & ~x819 & ~x861;
assign c2171 =  x8 &  x23 &  x26 &  x62 &  x122 &  x128 &  x197 &  x218 &  x305 &  x326 &  x335 &  x347 &  x386 &  x392 &  x413 &  x416 &  x422 &  x425 &  x430 &  x470 &  x476 &  x488 &  x491 &  x518 &  x542 &  x545 &  x548 &  x550 &  x554 &  x560 &  x593 &  x611 &  x667 &  x683 &  x737 &  x773 &  x833 &  x884 &  x899 &  x910 &  x923 &  x959 &  x961 &  x1019 &  x1028 &  x1034 &  x1040 &  x1115 & ~x663;
assign c2173 =  x406 &  x608 &  x677 &  x808 &  x1022 & ~x276 & ~x615 & ~x699 & ~x810;
assign c2175 =  x20 &  x32 &  x41 &  x47 &  x50 &  x56 &  x74 &  x95 &  x113 &  x131 &  x134 &  x143 &  x158 &  x161 &  x191 &  x194 &  x209 &  x227 &  x239 &  x245 &  x260 &  x266 &  x272 &  x278 &  x284 &  x299 &  x305 &  x308 &  x317 &  x332 &  x356 &  x377 &  x383 &  x395 &  x401 &  x404 &  x422 &  x428 &  x440 &  x458 &  x467 &  x476 &  x491 &  x494 &  x512 &  x521 &  x536 &  x575 &  x581 &  x589 &  x593 &  x596 &  x614 &  x617 &  x623 &  x628 &  x629 &  x638 &  x644 &  x650 &  x656 &  x667 &  x686 &  x725 &  x746 &  x761 &  x782 &  x800 &  x803 &  x839 &  x869 &  x884 &  x890 &  x893 &  x896 &  x905 &  x911 &  x917 &  x920 &  x929 &  x935 &  x938 &  x947 &  x959 &  x961 &  x998 &  x1019 &  x1027 &  x1028 &  x1039 &  x1040 &  x1072 &  x1085 &  x1091 &  x1094 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x897;
assign c2177 =  x25 &  x254 &  x628 &  x914 &  x961 &  x1000 & ~x813 & ~x852;
assign c2179 =  x196 &  x552 &  x590 &  x722 &  x782 &  x836 &  x905 & ~x408 & ~x447 & ~x897 & ~x936 & ~x978;
assign c2181 =  x981 & ~x234;
assign c2183 =  x592 &  x909 & ~x468 & ~x486;
assign c2185 =  x44 &  x50 &  x65 &  x86 &  x245 &  x257 &  x433 &  x511 &  x527 &  x557 &  x628 &  x707 &  x737 &  x844 &  x875 &  x883 &  x922 &  x989 & ~x483 & ~x936;
assign c2187 =  x57 &  x128 &  x244 &  x283 &  x340 &  x457 &  x1064;
assign c2189 =  x41 &  x86 &  x170 &  x218 &  x298 &  x299 &  x344 &  x362 &  x476 &  x493 &  x499 &  x545 &  x616 &  x788 &  x872 &  x917 &  x944 &  x1000 &  x1022 &  x1049 & ~x438 & ~x477;
assign c2191 =  x351 &  x469 &  x667 & ~x819 & ~x858;
assign c2193 =  x442 &  x491 &  x663 &  x668 & ~x354 & ~x510 & ~x591;
assign c2195 =  x74 &  x107 &  x518 &  x524 &  x644 &  x737 &  x808 &  x845 &  x863 &  x904 &  x910 &  x925 &  x980 & ~x564;
assign c2197 =  x89 &  x140 &  x323 &  x380 &  x389 &  x416 &  x527 &  x692 &  x752 &  x826 &  x865 & ~x81 & ~x117 & ~x609 & ~x642;
assign c2199 =  x748 &  x908 & ~x3 & ~x42 & ~x279 & ~x486 & ~x828;
assign c2201 =  x5 &  x8 &  x14 &  x17 &  x29 &  x32 &  x35 &  x41 &  x44 &  x53 &  x56 &  x59 &  x68 &  x77 &  x86 &  x89 &  x92 &  x95 &  x98 &  x107 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x134 &  x137 &  x149 &  x164 &  x173 &  x176 &  x182 &  x188 &  x197 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x227 &  x239 &  x248 &  x251 &  x257 &  x263 &  x266 &  x269 &  x272 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x308 &  x311 &  x317 &  x320 &  x326 &  x332 &  x335 &  x341 &  x349 &  x362 &  x368 &  x371 &  x377 &  x383 &  x388 &  x389 &  x392 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x437 &  x446 &  x455 &  x470 &  x476 &  x479 &  x482 &  x485 &  x491 &  x497 &  x500 &  x506 &  x509 &  x512 &  x515 &  x554 &  x563 &  x569 &  x572 &  x575 &  x593 &  x596 &  x611 &  x617 &  x626 &  x629 &  x638 &  x644 &  x650 &  x659 &  x665 &  x668 &  x671 &  x683 &  x689 &  x692 &  x698 &  x701 &  x742 &  x746 &  x749 &  x752 &  x755 &  x761 &  x779 &  x781 &  x782 &  x791 &  x800 &  x806 &  x815 &  x818 &  x820 &  x821 &  x824 &  x827 &  x830 &  x842 &  x845 &  x848 &  x859 &  x860 &  x881 &  x884 &  x887 &  x898 &  x908 &  x911 &  x917 &  x929 &  x932 &  x937 &  x940 &  x941 &  x947 &  x956 &  x962 &  x976 &  x977 &  x978 &  x986 &  x989 &  x998 &  x1001 &  x1007 &  x1010 &  x1017 &  x1018 &  x1022 &  x1025 &  x1046 &  x1052 &  x1055 &  x1056 &  x1058 &  x1061 &  x1064 &  x1067 &  x1076 &  x1082 &  x1088 &  x1096 &  x1097 &  x1103 &  x1115 &  x1121 &  x1124 &  x1127;
assign c2203 =  x1130 & ~x84 & ~x309 & ~x462 & ~x774 & ~x819 & ~x1059;
assign c2205 =  x41 &  x65 &  x86 &  x200 &  x206 &  x209 &  x350 &  x440 &  x509 &  x515 &  x572 &  x653 &  x788 &  x818 &  x871 &  x959 &  x1025 &  x1049 &  x1055 & ~x141 & ~x516 & ~x558 & ~x708 & ~x1020;
assign c2207 =  x8 &  x17 &  x50 &  x65 &  x68 &  x74 &  x92 &  x107 &  x110 &  x116 &  x131 &  x146 &  x164 &  x173 &  x182 &  x185 &  x188 &  x203 &  x221 &  x224 &  x245 &  x269 &  x284 &  x287 &  x296 &  x299 &  x302 &  x308 &  x314 &  x341 &  x359 &  x362 &  x371 &  x377 &  x380 &  x383 &  x392 &  x395 &  x398 &  x413 &  x422 &  x443 &  x458 &  x464 &  x479 &  x503 &  x506 &  x509 &  x518 &  x530 &  x539 &  x542 &  x551 &  x572 &  x581 &  x614 &  x650 &  x656 &  x698 &  x719 &  x725 &  x743 &  x755 &  x764 &  x779 &  x812 &  x824 &  x830 &  x854 &  x857 &  x881 &  x917 &  x926 &  x950 &  x965 &  x968 &  x992 &  x1004 &  x1022 &  x1025 &  x1028 &  x1034 &  x1046 &  x1052 &  x1060 &  x1064 &  x1079 &  x1082 &  x1091 &  x1099 &  x1100 &  x1115 & ~x204 & ~x423 & ~x513 & ~x771;
assign c2209 =  x79 & ~x84 & ~x97 & ~x309 & ~x381 & ~x615 & ~x783;
assign c2211 =  x14 &  x421 &  x613 &  x614 &  x632 &  x701 &  x937 &  x976 &  x1000;
assign c2213 =  x747 &  x904 & ~x334;
assign c2215 =  x980 &  x1007 & ~x276 & ~x660 & ~x969 & ~x1029 & ~x1068 & ~x1086;
assign c2217 =  x122 &  x254 &  x343 &  x585 &  x703 &  x1126 & ~x553 & ~x1065;
assign c2219 =  x580 & ~x526 & ~x661;
assign c2221 =  x2 &  x89 &  x104 &  x110 &  x158 &  x209 &  x233 &  x287 &  x290 &  x344 &  x359 &  x413 &  x461 &  x481 &  x482 &  x485 &  x497 &  x575 &  x650 &  x656 &  x662 &  x698 &  x710 &  x716 &  x718 &  x728 &  x731 &  x782 &  x788 &  x815 &  x824 &  x842 &  x878 &  x884 &  x911 &  x920 &  x932 &  x935 &  x968 &  x986 &  x992 &  x1001 &  x1055 &  x1082 & ~x348 & ~x384 & ~x423 & ~x489 & ~x744 & ~x783 & ~x822;
assign c2223 =  x858 &  x936 &  x1017 &  x1056 & ~x510;
assign c2225 =  x781 &  x940 &  x1096 & ~x871 & ~x913;
assign c2227 =  x223 &  x865 & ~x490 & ~x615;
assign c2229 =  x41 &  x53 &  x74 &  x140 &  x161 &  x167 &  x173 &  x182 &  x284 &  x337 &  x421 &  x452 &  x464 &  x485 &  x527 &  x626 &  x652 &  x713 &  x719 &  x734 &  x740 &  x749 &  x770 &  x773 &  x806 &  x812 &  x827 &  x859 &  x863 &  x869 &  x937 &  x980 &  x1000 &  x1010 &  x1028 &  x1064 &  x1097 &  x1103 &  x1115;
assign c2231 =  x41 &  x176 &  x346 &  x566 &  x586 &  x695 &  x701 &  x725 &  x734 &  x860 &  x979 &  x1019 &  x1028 &  x1052 & ~x516 & ~x597;
assign c2233 =  x897 &  x1020;
assign c2235 =  x77 &  x80 &  x95 &  x128 &  x191 &  x197 &  x254 &  x257 &  x305 &  x347 &  x362 &  x401 &  x437 &  x467 &  x472 &  x511 &  x530 &  x545 &  x548 &  x602 &  x668 &  x719 &  x812 &  x815 &  x1001 &  x1037 & ~x579 & ~x618 & ~x660 & ~x801 & ~x813;
assign c2237 =  x510 & ~x478;
assign c2239 =  x340 &  x392 &  x665 &  x741 & ~x513 & ~x630;
assign c2241 =  x442 &  x1096 & ~x832 & ~x849 & ~x871;
assign c2243 =  x32 &  x44 &  x71 &  x152 &  x158 &  x194 &  x212 &  x247 &  x272 &  x314 &  x374 &  x406 &  x431 &  x479 &  x524 &  x530 &  x560 &  x593 &  x599 &  x614 &  x625 &  x662 &  x701 &  x713 &  x725 &  x806 &  x815 &  x818 &  x826 &  x830 &  x842 &  x878 &  x908 &  x911 &  x929 &  x932 &  x944 &  x953 &  x959 &  x962 &  x965 &  x1001 &  x1022 &  x1058 &  x1073 &  x1115 &  x1121 & ~x738 & ~x816 & ~x1011;
assign c2245 =  x91 &  x546 & ~x315 & ~x474 & ~x636 & ~x675;
assign c2247 =  x72 &  x111 &  x458 & ~x108 & ~x252 & ~x894 & ~x933 & ~x1122;
assign c2249 = ~x333 & ~x874 & ~x969;
assign c2251 =  x29 &  x41 &  x44 &  x80 &  x92 &  x113 &  x131 &  x137 &  x140 &  x164 &  x182 &  x191 &  x194 &  x209 &  x218 &  x248 &  x260 &  x269 &  x278 &  x284 &  x296 &  x299 &  x302 &  x314 &  x320 &  x323 &  x347 &  x356 &  x368 &  x374 &  x389 &  x392 &  x401 &  x404 &  x422 &  x425 &  x476 &  x485 &  x488 &  x497 &  x506 &  x509 &  x515 &  x530 &  x536 &  x551 &  x563 &  x566 &  x572 &  x575 &  x578 &  x587 &  x590 &  x596 &  x623 &  x632 &  x641 &  x656 &  x662 &  x665 &  x668 &  x719 &  x731 &  x779 &  x797 &  x800 &  x806 &  x827 &  x830 &  x836 &  x839 &  x845 &  x851 &  x854 &  x863 &  x866 &  x869 &  x881 &  x887 &  x890 &  x893 &  x925 &  x947 &  x958 &  x986 &  x998 &  x1004 &  x1028 &  x1034 &  x1037 &  x1073 &  x1079 &  x1091 &  x1103 &  x1106 &  x1121 & ~x42 & ~x819;
assign c2253 =  x787 & ~x120 & ~x682;
assign c2255 =  x77 &  x116 &  x179 &  x343 &  x496 &  x656 &  x788 &  x818 &  x926 & ~x42 & ~x159 & ~x513 & ~x591 & ~x708;
assign c2257 =  x17 &  x23 &  x32 &  x35 &  x44 &  x47 &  x50 &  x68 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x113 &  x119 &  x128 &  x134 &  x140 &  x173 &  x176 &  x182 &  x188 &  x200 &  x203 &  x206 &  x209 &  x227 &  x230 &  x251 &  x263 &  x278 &  x284 &  x290 &  x302 &  x305 &  x308 &  x317 &  x344 &  x347 &  x356 &  x371 &  x374 &  x386 &  x398 &  x404 &  x410 &  x425 &  x428 &  x446 &  x458 &  x461 &  x467 &  x476 &  x488 &  x512 &  x545 &  x581 &  x587 &  x596 &  x614 &  x620 &  x632 &  x638 &  x647 &  x653 &  x656 &  x659 &  x677 &  x680 &  x692 &  x695 &  x698 &  x704 &  x707 &  x725 &  x734 &  x737 &  x743 &  x746 &  x761 &  x764 &  x776 &  x785 &  x791 &  x794 &  x815 &  x823 &  x830 &  x836 &  x845 &  x854 &  x857 &  x860 &  x862 &  x863 &  x872 &  x881 &  x929 &  x938 &  x940 &  x959 &  x968 &  x974 &  x979 &  x980 &  x995 &  x998 &  x1010 &  x1018 &  x1025 &  x1052 &  x1057 &  x1076 &  x1079 &  x1091 &  x1100 &  x1106 &  x1109 &  x1127 & ~x159 & ~x1047 & ~x1086;
assign c2259 =  x38 &  x65 &  x68 &  x83 &  x89 &  x95 &  x107 &  x173 &  x230 &  x263 &  x278 &  x287 &  x323 &  x326 &  x350 &  x395 &  x467 &  x476 &  x488 &  x497 &  x515 &  x536 &  x568 &  x593 &  x623 &  x631 &  x646 &  x650 &  x653 &  x656 &  x709 &  x710 &  x725 &  x737 &  x746 &  x755 &  x776 &  x787 &  x797 &  x818 &  x824 &  x890 &  x893 &  x911 &  x914 &  x950 &  x980 &  x983 &  x1016 &  x1049 &  x1070 &  x1118 & ~x549 & ~x981 & ~x1104 & ~x1107;
assign c2261 =  x14 &  x20 &  x65 &  x74 &  x77 &  x86 &  x92 &  x185 &  x191 &  x200 &  x215 &  x224 &  x266 &  x284 &  x293 &  x302 &  x317 &  x323 &  x347 &  x356 &  x413 &  x455 &  x470 &  x503 &  x509 &  x545 &  x557 &  x638 &  x641 &  x650 &  x680 &  x685 &  x689 &  x704 &  x719 &  x727 &  x733 &  x737 &  x749 &  x772 &  x779 &  x782 &  x788 &  x791 &  x800 &  x821 &  x827 &  x851 &  x860 &  x883 &  x893 &  x899 &  x911 &  x953 &  x961 &  x983 &  x1000 &  x1001 &  x1016 &  x1106 &  x1118 & ~x201 & ~x981 & ~x1020 & ~x1098;
assign c2263 =  x8 &  x14 &  x32 &  x44 &  x56 &  x77 &  x79 &  x80 &  x86 &  x98 &  x118 &  x119 &  x128 &  x131 &  x146 &  x157 &  x164 &  x167 &  x182 &  x191 &  x206 &  x209 &  x218 &  x221 &  x233 &  x236 &  x248 &  x257 &  x260 &  x266 &  x269 &  x272 &  x281 &  x299 &  x311 &  x316 &  x329 &  x338 &  x355 &  x362 &  x365 &  x374 &  x386 &  x394 &  x404 &  x410 &  x416 &  x425 &  x433 &  x440 &  x458 &  x470 &  x482 &  x488 &  x491 &  x494 &  x497 &  x512 &  x515 &  x518 &  x527 &  x530 &  x533 &  x536 &  x539 &  x545 &  x560 &  x569 &  x584 &  x587 &  x599 &  x602 &  x605 &  x629 &  x644 &  x665 &  x670 &  x671 &  x680 &  x686 &  x698 &  x701 &  x713 &  x716 &  x719 &  x721 &  x728 &  x746 &  x749 &  x752 &  x779 &  x782 &  x785 &  x787 &  x788 &  x794 &  x799 &  x800 &  x806 &  x815 &  x818 &  x824 &  x832 &  x848 &  x856 &  x869 &  x871 &  x878 &  x884 &  x887 &  x893 &  x902 &  x905 &  x910 &  x929 &  x938 &  x941 &  x944 &  x947 &  x956 &  x974 &  x980 &  x986 &  x989 &  x995 &  x998 &  x1016 &  x1028 &  x1040 &  x1052 &  x1070 &  x1085 &  x1091 &  x1094 &  x1103 &  x1109 &  x1118 &  x1124 &  x1127 & ~x702 & ~x783 & ~x900;
assign c2265 =  x181 &  x625 &  x783;
assign c2267 =  x11 &  x107 &  x110 &  x113 &  x125 &  x134 &  x200 &  x218 &  x260 &  x266 &  x272 &  x476 &  x510 &  x587 &  x623 &  x628 &  x773 &  x836 &  x899 &  x986 &  x1070 &  x1106 & ~x438 & ~x477 & ~x618;
assign c2269 =  x233 &  x346 &  x518 &  x617 &  x823 &  x901 &  x940 &  x1100 & ~x198 & ~x486 & ~x672;
assign c2271 =  x218 &  x235 &  x395 &  x513 &  x518 &  x815 &  x916 &  x998 & ~x447 & ~x741;
assign c2273 =  x56 &  x61 &  x62 &  x83 &  x92 &  x101 &  x110 &  x137 &  x140 &  x146 &  x155 &  x173 &  x215 &  x236 &  x239 &  x266 &  x275 &  x287 &  x293 &  x304 &  x311 &  x326 &  x335 &  x337 &  x359 &  x386 &  x404 &  x416 &  x421 &  x446 &  x452 &  x455 &  x458 &  x476 &  x497 &  x515 &  x533 &  x539 &  x554 &  x566 &  x587 &  x596 &  x620 &  x701 &  x713 &  x728 &  x737 &  x755 &  x757 &  x770 &  x809 &  x824 &  x836 &  x839 &  x845 &  x866 &  x881 &  x965 &  x989 &  x992 &  x998 &  x1007 &  x1025 &  x1031 &  x1037 &  x1043 &  x1079 &  x1082 &  x1084 &  x1091 &  x1121 & ~x471;
assign c2275 =  x382 &  x718 &  x897 &  x975;
assign c2277 =  x175 &  x226 &  x265 &  x1117 & ~x1069;
assign c2279 =  x11 &  x62 &  x311 &  x312 &  x748 &  x995 & ~x201 & ~x448;
assign c2281 =  x2 &  x14 &  x17 &  x47 &  x107 &  x131 &  x140 &  x143 &  x173 &  x188 &  x209 &  x266 &  x278 &  x356 &  x359 &  x368 &  x404 &  x416 &  x455 &  x464 &  x485 &  x515 &  x545 &  x551 &  x554 &  x611 &  x638 &  x647 &  x677 &  x701 &  x707 &  x716 &  x731 &  x770 &  x772 &  x773 &  x776 &  x779 &  x872 &  x884 &  x890 &  x893 &  x941 &  x959 &  x965 &  x983 &  x1019 &  x1031 &  x1043 &  x1067 &  x1070 &  x1091 &  x1115 &  x1130 & ~x45 & ~x108 & ~x618 & ~x774 & ~x1026;
assign c2283 =  x125 &  x421 &  x452 &  x484 &  x530 &  x575 &  x758 &  x769 &  x884 &  x885 &  x935 &  x937 &  x968 &  x1013 & ~x510;
assign c2285 =  x62 &  x65 &  x119 &  x122 &  x209 &  x227 &  x239 &  x260 &  x329 &  x368 &  x392 &  x395 &  x407 &  x431 &  x464 &  x476 &  x488 &  x524 &  x530 &  x539 &  x593 &  x602 &  x647 &  x653 &  x662 &  x745 &  x746 &  x752 &  x776 &  x791 &  x794 &  x818 &  x821 &  x884 &  x905 &  x923 &  x944 &  x953 &  x959 &  x965 &  x983 &  x998 &  x1016 &  x1021 &  x1049 &  x1060 &  x1061 &  x1106 & ~x81 & ~x600;
assign c2287 =  x960 & ~x373;
assign c2289 =  x2 &  x11 &  x86 &  x281 &  x320 &  x323 &  x341 &  x353 &  x394 &  x497 &  x527 &  x533 &  x560 &  x641 &  x755 &  x782 &  x794 &  x851 &  x878 &  x881 &  x902 &  x908 &  x956 &  x959 &  x1007 &  x1082 &  x1097 &  x1103 & ~x108 & ~x213 & ~x858 & ~x978 & ~x1020;
assign c2291 =  x292 &  x1056 & ~x312;
assign c2293 = ~x562 & ~x1024;
assign c2295 =  x2 &  x26 &  x71 &  x98 &  x146 &  x242 &  x260 &  x281 &  x305 &  x329 &  x557 &  x580 &  x641 &  x653 &  x704 &  x743 &  x773 &  x806 &  x848 &  x905 &  x926 &  x940 &  x944 &  x977 &  x1013 &  x1016 &  x1121 & ~x195 & ~x237 & ~x276 & ~x354 & ~x393 & ~x747;
assign c2297 =  x418 &  x678 & ~x688;
assign c2299 =  x71 &  x589 &  x983 &  x994 &  x1006 & ~x387 & ~x819;
assign c30 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x302 &  x305 &  x308 &  x314 &  x317 &  x320 &  x323 &  x325 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x364 &  x365 &  x368 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x403 &  x404 &  x407 &  x409 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x442 &  x443 &  x448 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x478 &  x479 &  x481 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x517 &  x518 &  x519 &  x520 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x556 &  x557 &  x559 &  x560 &  x563 &  x566 &  x569 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x595 &  x596 &  x599 &  x602 &  x605 &  x611 &  x614 &  x617 &  x620 &  x623 &  x628 &  x629 &  x632 &  x634 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x667 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x704 &  x707 &  x710 &  x716 &  x719 &  x725 &  x728 &  x734 &  x737 &  x740 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x784 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x901 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x940 &  x944 &  x946 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1018 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1057 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 &  x1130;
assign c32 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x26 &  x29 &  x41 &  x47 &  x56 &  x62 &  x71 &  x74 &  x77 &  x83 &  x86 &  x92 &  x95 &  x98 &  x107 &  x113 &  x119 &  x122 &  x128 &  x137 &  x161 &  x164 &  x170 &  x182 &  x185 &  x188 &  x194 &  x199 &  x200 &  x206 &  x212 &  x218 &  x224 &  x230 &  x233 &  x236 &  x238 &  x239 &  x248 &  x263 &  x266 &  x287 &  x290 &  x293 &  x302 &  x314 &  x316 &  x317 &  x326 &  x329 &  x341 &  x344 &  x355 &  x368 &  x380 &  x383 &  x389 &  x394 &  x395 &  x398 &  x401 &  x413 &  x419 &  x422 &  x425 &  x433 &  x440 &  x455 &  x464 &  x470 &  x472 &  x473 &  x482 &  x488 &  x494 &  x503 &  x509 &  x521 &  x530 &  x536 &  x545 &  x548 &  x551 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x593 &  x596 &  x599 &  x602 &  x605 &  x617 &  x623 &  x626 &  x631 &  x638 &  x641 &  x647 &  x662 &  x670 &  x674 &  x695 &  x701 &  x704 &  x707 &  x716 &  x746 &  x749 &  x752 &  x754 &  x758 &  x773 &  x776 &  x785 &  x788 &  x791 &  x793 &  x797 &  x803 &  x812 &  x821 &  x824 &  x830 &  x836 &  x842 &  x848 &  x854 &  x857 &  x866 &  x871 &  x875 &  x878 &  x883 &  x884 &  x899 &  x905 &  x908 &  x911 &  x916 &  x917 &  x932 &  x938 &  x947 &  x949 &  x956 &  x959 &  x962 &  x968 &  x974 &  x983 &  x988 &  x989 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1019 &  x1034 &  x1055 &  x1058 &  x1061 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1100 &  x1106 &  x1109 &  x1124 &  x1127 &  x1130 & ~x105 & ~x639 & ~x663 & ~x702 & ~x741 & ~x780 & ~x781 & ~x819 & ~x930 & ~x945 & ~x1023 & ~x1092;
assign c34 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x125 &  x128 &  x134 &  x137 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x448 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x614 &  x617 &  x620 &  x623 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x869 &  x875 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x901 &  x905 &  x911 &  x914 &  x920 &  x923 &  x926 &  x929 &  x935 &  x938 &  x940 &  x941 &  x944 &  x947 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x75 & ~x114 & ~x153 & ~x243 & ~x282 & ~x321 & ~x360 & ~x912 & ~x951 & ~x990 & ~x1029 & ~x1113;
assign c36 =  x2 &  x11 &  x14 &  x17 &  x32 &  x35 &  x38 &  x41 &  x44 &  x59 &  x68 &  x71 &  x80 &  x86 &  x92 &  x95 &  x116 &  x134 &  x140 &  x149 &  x155 &  x161 &  x164 &  x167 &  x176 &  x182 &  x185 &  x194 &  x197 &  x200 &  x203 &  x206 &  x215 &  x224 &  x236 &  x242 &  x248 &  x251 &  x263 &  x287 &  x289 &  x290 &  x293 &  x305 &  x307 &  x314 &  x332 &  x344 &  x347 &  x356 &  x367 &  x371 &  x374 &  x386 &  x389 &  x392 &  x395 &  x398 &  x403 &  x406 &  x407 &  x413 &  x422 &  x425 &  x442 &  x443 &  x446 &  x452 &  x464 &  x481 &  x482 &  x491 &  x497 &  x503 &  x512 &  x521 &  x523 &  x527 &  x530 &  x533 &  x536 &  x554 &  x560 &  x566 &  x581 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x607 &  x608 &  x614 &  x617 &  x620 &  x623 &  x629 &  x632 &  x635 &  x641 &  x653 &  x668 &  x671 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x701 &  x703 &  x704 &  x706 &  x710 &  x713 &  x722 &  x734 &  x737 &  x742 &  x743 &  x745 &  x746 &  x749 &  x764 &  x767 &  x776 &  x779 &  x782 &  x784 &  x785 &  x788 &  x794 &  x797 &  x803 &  x809 &  x812 &  x820 &  x821 &  x824 &  x836 &  x839 &  x842 &  x845 &  x848 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x878 &  x884 &  x890 &  x893 &  x896 &  x901 &  x902 &  x907 &  x911 &  x920 &  x923 &  x929 &  x932 &  x937 &  x938 &  x940 &  x946 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x985 &  x995 &  x998 &  x1001 &  x1010 &  x1019 &  x1022 &  x1025 &  x1034 &  x1040 &  x1043 &  x1055 &  x1057 &  x1070 &  x1073 &  x1085 &  x1088 &  x1091 &  x1100 &  x1103 &  x1106 &  x1112 &  x1124;
assign c38 =  x17 &  x20 &  x26 &  x29 &  x35 &  x38 &  x47 &  x53 &  x56 &  x59 &  x71 &  x83 &  x89 &  x101 &  x104 &  x107 &  x116 &  x125 &  x128 &  x143 &  x158 &  x161 &  x164 &  x167 &  x173 &  x176 &  x185 &  x197 &  x200 &  x203 &  x218 &  x221 &  x230 &  x236 &  x239 &  x247 &  x248 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x278 &  x290 &  x293 &  x296 &  x299 &  x302 &  x311 &  x326 &  x331 &  x347 &  x353 &  x356 &  x359 &  x371 &  x374 &  x380 &  x389 &  x392 &  x395 &  x398 &  x404 &  x407 &  x410 &  x413 &  x419 &  x425 &  x446 &  x449 &  x452 &  x467 &  x470 &  x482 &  x485 &  x491 &  x494 &  x497 &  x509 &  x524 &  x533 &  x539 &  x542 &  x545 &  x548 &  x550 &  x551 &  x557 &  x569 &  x572 &  x581 &  x589 &  x593 &  x596 &  x602 &  x608 &  x611 &  x617 &  x623 &  x626 &  x628 &  x632 &  x638 &  x641 &  x667 &  x680 &  x683 &  x695 &  x701 &  x707 &  x709 &  x719 &  x722 &  x745 &  x746 &  x747 &  x749 &  x752 &  x755 &  x758 &  x764 &  x767 &  x770 &  x776 &  x779 &  x784 &  x785 &  x797 &  x803 &  x812 &  x818 &  x821 &  x827 &  x830 &  x839 &  x851 &  x857 &  x860 &  x869 &  x878 &  x887 &  x890 &  x902 &  x920 &  x926 &  x929 &  x944 &  x956 &  x983 &  x986 &  x994 &  x1001 &  x1004 &  x1007 &  x1019 &  x1028 &  x1031 &  x1034 &  x1040 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1094 &  x1106 &  x1109 &  x1115 &  x1118 &  x1127 & ~x156 & ~x663 & ~x702 & ~x780 & ~x819 & ~x936;
assign c310 =  x5 &  x11 &  x14 &  x17 &  x20 &  x23 &  x29 &  x35 &  x38 &  x44 &  x50 &  x53 &  x56 &  x59 &  x65 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x119 &  x125 &  x128 &  x134 &  x137 &  x146 &  x152 &  x155 &  x161 &  x164 &  x170 &  x173 &  x176 &  x179 &  x182 &  x188 &  x191 &  x194 &  x206 &  x209 &  x215 &  x218 &  x221 &  x224 &  x226 &  x227 &  x230 &  x233 &  x236 &  x239 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x265 &  x266 &  x272 &  x275 &  x281 &  x284 &  x286 &  x287 &  x289 &  x290 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x317 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x353 &  x359 &  x362 &  x370 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x395 &  x398 &  x401 &  x403 &  x404 &  x407 &  x410 &  x413 &  x419 &  x431 &  x434 &  x437 &  x440 &  x442 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x464 &  x470 &  x476 &  x480 &  x481 &  x485 &  x494 &  x497 &  x503 &  x506 &  x512 &  x515 &  x518 &  x521 &  x524 &  x530 &  x536 &  x539 &  x542 &  x548 &  x554 &  x556 &  x560 &  x563 &  x566 &  x569 &  x575 &  x581 &  x587 &  x590 &  x593 &  x595 &  x596 &  x602 &  x614 &  x617 &  x623 &  x626 &  x629 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x674 &  x680 &  x683 &  x686 &  x689 &  x698 &  x704 &  x707 &  x716 &  x719 &  x722 &  x725 &  x731 &  x734 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x794 &  x800 &  x803 &  x806 &  x809 &  x815 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x872 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x902 &  x905 &  x908 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x941 &  x944 &  x950 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1061 &  x1067 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1109 &  x1115 &  x1118 &  x1121 &  x1127 & ~x390 & ~x813;
assign c312 =  x2 &  x5 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x35 &  x38 &  x41 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x395 &  x398 &  x401 &  x403 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x434 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x481 &  x482 &  x485 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x520 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x554 &  x557 &  x559 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x626 &  x629 &  x632 &  x635 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x776 &  x779 &  x782 &  x785 &  x788 &  x794 &  x797 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x836 &  x842 &  x845 &  x848 &  x851 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x901 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x940 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x979 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1018 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1057 &  x1058 &  x1061 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x3 & ~x42 & ~x81 & ~x117 & ~x156 & ~x195 & ~x234 & ~x273 & ~x312 & ~x390 & ~x429 & ~x996 & ~x1035 & ~x1074;
assign c314 =  x2 &  x8 &  x17 &  x23 &  x26 &  x35 &  x41 &  x44 &  x53 &  x65 &  x68 &  x77 &  x83 &  x86 &  x89 &  x92 &  x101 &  x110 &  x113 &  x116 &  x119 &  x122 &  x134 &  x137 &  x155 &  x160 &  x164 &  x167 &  x170 &  x176 &  x185 &  x188 &  x197 &  x199 &  x200 &  x203 &  x209 &  x212 &  x221 &  x236 &  x238 &  x239 &  x248 &  x251 &  x257 &  x260 &  x269 &  x272 &  x275 &  x281 &  x284 &  x290 &  x293 &  x296 &  x299 &  x305 &  x308 &  x314 &  x317 &  x320 &  x326 &  x329 &  x332 &  x335 &  x338 &  x344 &  x350 &  x355 &  x368 &  x371 &  x374 &  x380 &  x383 &  x394 &  x395 &  x407 &  x410 &  x413 &  x419 &  x422 &  x431 &  x433 &  x440 &  x443 &  x464 &  x467 &  x470 &  x476 &  x482 &  x485 &  x491 &  x506 &  x509 &  x511 &  x512 &  x527 &  x530 &  x536 &  x539 &  x548 &  x551 &  x560 &  x578 &  x581 &  x587 &  x589 &  x593 &  x596 &  x599 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x628 &  x635 &  x638 &  x650 &  x653 &  x665 &  x671 &  x677 &  x689 &  x692 &  x695 &  x698 &  x704 &  x722 &  x725 &  x728 &  x737 &  x740 &  x746 &  x752 &  x755 &  x764 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x830 &  x833 &  x836 &  x839 &  x851 &  x854 &  x857 &  x869 &  x875 &  x878 &  x881 &  x884 &  x896 &  x899 &  x905 &  x908 &  x914 &  x917 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x956 &  x962 &  x968 &  x971 &  x974 &  x992 &  x995 &  x1001 &  x1010 &  x1013 &  x1019 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1061 &  x1076 &  x1085 &  x1091 &  x1097 &  x1100 &  x1109 &  x1112 &  x1118 &  x1124 &  x1127 &  x1130 & ~x537 & ~x561 & ~x576 & ~x600 & ~x609 & ~x615 & ~x717 & ~x795 & ~x834;
assign c316 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x265 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x304 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x343 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x382 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x421 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x460 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x499 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x538 &  x539 &  x542 &  x545 &  x548 &  x551 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x577 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x616 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x643 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1018 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1054 &  x1055 &  x1057 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1096 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x1032 & ~x1038 & ~x1071 & ~x1072 & ~x1110 & ~x1128;
assign c318 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x134 &  x140 &  x143 &  x146 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x319 &  x320 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x358 &  x359 &  x362 &  x364 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x401 &  x403 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x442 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x470 &  x473 &  x476 &  x481 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x520 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x584 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x617 &  x620 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x770 &  x773 &  x776 &  x779 &  x781 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x820 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x836 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x859 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x898 &  x899 &  x901 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x940 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x976 &  x977 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1015 &  x1018 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1057 &  x1058 &  x1060 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1096 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x159 & ~x198 & ~x234 & ~x237 & ~x273 & ~x312 & ~x315 & ~x351 & ~x390 & ~x429 & ~x873 & ~x912 & ~x951;
assign c320 =  x8 &  x17 &  x26 &  x32 &  x44 &  x47 &  x53 &  x56 &  x59 &  x65 &  x71 &  x83 &  x86 &  x92 &  x95 &  x98 &  x107 &  x110 &  x116 &  x122 &  x137 &  x140 &  x143 &  x158 &  x173 &  x188 &  x191 &  x202 &  x206 &  x212 &  x215 &  x224 &  x227 &  x236 &  x242 &  x245 &  x251 &  x260 &  x265 &  x269 &  x272 &  x278 &  x284 &  x290 &  x293 &  x305 &  x308 &  x311 &  x320 &  x323 &  x335 &  x338 &  x347 &  x353 &  x356 &  x362 &  x368 &  x371 &  x376 &  x380 &  x383 &  x395 &  x404 &  x407 &  x416 &  x419 &  x428 &  x431 &  x434 &  x440 &  x446 &  x467 &  x470 &  x476 &  x479 &  x488 &  x491 &  x497 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x542 &  x548 &  x554 &  x563 &  x572 &  x575 &  x578 &  x584 &  x587 &  x605 &  x620 &  x629 &  x632 &  x638 &  x644 &  x650 &  x653 &  x659 &  x668 &  x671 &  x674 &  x686 &  x689 &  x698 &  x701 &  x704 &  x713 &  x719 &  x743 &  x761 &  x773 &  x779 &  x788 &  x800 &  x812 &  x821 &  x827 &  x839 &  x848 &  x851 &  x854 &  x860 &  x872 &  x875 &  x881 &  x884 &  x899 &  x901 &  x907 &  x914 &  x917 &  x923 &  x926 &  x929 &  x938 &  x944 &  x947 &  x950 &  x965 &  x971 &  x977 &  x980 &  x983 &  x986 &  x992 &  x995 &  x1004 &  x1019 &  x1043 &  x1046 &  x1049 &  x1058 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1097 &  x1100 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1130 & ~x156 & ~x159 & ~x234 & ~x351 & ~x657 & ~x697 & ~x735 & ~x774;
assign c322 =  x8 &  x29 &  x35 &  x41 &  x74 &  x77 &  x86 &  x92 &  x98 &  x110 &  x116 &  x128 &  x137 &  x158 &  x176 &  x179 &  x182 &  x197 &  x206 &  x209 &  x218 &  x230 &  x236 &  x248 &  x254 &  x260 &  x266 &  x269 &  x272 &  x275 &  x296 &  x302 &  x305 &  x308 &  x317 &  x320 &  x326 &  x335 &  x350 &  x353 &  x356 &  x359 &  x368 &  x374 &  x377 &  x380 &  x392 &  x395 &  x419 &  x431 &  x434 &  x443 &  x445 &  x446 &  x455 &  x461 &  x476 &  x482 &  x488 &  x497 &  x503 &  x524 &  x530 &  x542 &  x551 &  x557 &  x563 &  x566 &  x572 &  x578 &  x589 &  x590 &  x605 &  x623 &  x626 &  x628 &  x641 &  x656 &  x662 &  x674 &  x680 &  x683 &  x698 &  x707 &  x710 &  x713 &  x728 &  x736 &  x740 &  x742 &  x755 &  x758 &  x761 &  x764 &  x773 &  x774 &  x776 &  x788 &  x791 &  x797 &  x800 &  x803 &  x812 &  x821 &  x833 &  x845 &  x848 &  x851 &  x853 &  x857 &  x872 &  x878 &  x884 &  x887 &  x890 &  x892 &  x899 &  x902 &  x920 &  x923 &  x926 &  x937 &  x940 &  x944 &  x947 &  x968 &  x970 &  x971 &  x976 &  x977 &  x979 &  x980 &  x983 &  x989 &  x992 &  x1004 &  x1007 &  x1009 &  x1019 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1097 &  x1106 &  x1118 &  x1124 &  x1130;
assign c324 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x325 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x355 &  x356 &  x359 &  x362 &  x364 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x394 &  x395 &  x398 &  x401 &  x403 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x433 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x472 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x508 &  x509 &  x511 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x547 &  x548 &  x550 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x589 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x625 &  x626 &  x628 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x667 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x703 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x826 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x417;
assign c326 =  x2 &  x5 &  x8 &  x11 &  x17 &  x20 &  x26 &  x29 &  x35 &  x41 &  x44 &  x47 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x122 &  x128 &  x134 &  x137 &  x149 &  x152 &  x164 &  x167 &  x170 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x205 &  x209 &  x212 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x242 &  x248 &  x257 &  x260 &  x266 &  x269 &  x272 &  x275 &  x281 &  x287 &  x290 &  x293 &  x296 &  x302 &  x305 &  x308 &  x311 &  x317 &  x320 &  x323 &  x326 &  x335 &  x341 &  x347 &  x352 &  x356 &  x359 &  x368 &  x371 &  x374 &  x377 &  x389 &  x391 &  x394 &  x398 &  x401 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x433 &  x434 &  x437 &  x440 &  x443 &  x446 &  x452 &  x455 &  x458 &  x461 &  x464 &  x470 &  x472 &  x476 &  x479 &  x488 &  x491 &  x503 &  x506 &  x509 &  x511 &  x515 &  x521 &  x524 &  x530 &  x539 &  x542 &  x550 &  x551 &  x557 &  x560 &  x566 &  x569 &  x572 &  x581 &  x584 &  x589 &  x593 &  x596 &  x599 &  x602 &  x605 &  x614 &  x617 &  x626 &  x628 &  x629 &  x638 &  x650 &  x656 &  x668 &  x671 &  x674 &  x677 &  x683 &  x686 &  x689 &  x695 &  x698 &  x707 &  x709 &  x710 &  x713 &  x719 &  x722 &  x731 &  x740 &  x743 &  x755 &  x773 &  x776 &  x785 &  x787 &  x812 &  x815 &  x818 &  x821 &  x830 &  x833 &  x836 &  x845 &  x854 &  x857 &  x866 &  x869 &  x872 &  x881 &  x887 &  x893 &  x902 &  x905 &  x908 &  x914 &  x920 &  x929 &  x932 &  x935 &  x938 &  x944 &  x950 &  x953 &  x956 &  x959 &  x974 &  x977 &  x980 &  x983 &  x998 &  x1001 &  x1010 &  x1016 &  x1022 &  x1031 &  x1037 &  x1043 &  x1046 &  x1058 &  x1067 &  x1070 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1100 &  x1109 &  x1115 &  x1127 &  x1130 & ~x357 & ~x600 & ~x601 & ~x639 & ~x702 & ~x741 & ~x780 & ~x819 & ~x858;
assign c328 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x23 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x356 &  x359 &  x364 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x403 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x442 &  x443 &  x446 &  x448 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x473 &  x476 &  x479 &  x481 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x568 &  x569 &  x572 &  x575 &  x578 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x607 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x646 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x667 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x745 &  x746 &  x749 &  x752 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x781 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x820 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x836 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x859 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x878 &  x884 &  x887 &  x890 &  x893 &  x896 &  x898 &  x899 &  x901 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x937 &  x940 &  x941 &  x944 &  x947 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x976 &  x977 &  x979 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1015 &  x1016 &  x1019 &  x1021 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1057 &  x1058 &  x1060 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1096 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x195 & ~x234 & ~x312;
assign c330 =  x8 &  x14 &  x17 &  x20 &  x23 &  x26 &  x28 &  x29 &  x32 &  x35 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x61 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x86 &  x92 &  x95 &  x98 &  x100 &  x101 &  x104 &  x107 &  x110 &  x112 &  x116 &  x119 &  x122 &  x128 &  x131 &  x134 &  x137 &  x139 &  x140 &  x143 &  x145 &  x146 &  x149 &  x151 &  x152 &  x158 &  x161 &  x164 &  x167 &  x173 &  x178 &  x179 &  x182 &  x184 &  x185 &  x190 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x211 &  x212 &  x217 &  x218 &  x221 &  x224 &  x227 &  x229 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x250 &  x251 &  x254 &  x256 &  x257 &  x260 &  x262 &  x263 &  x266 &  x268 &  x269 &  x275 &  x278 &  x281 &  x284 &  x287 &  x289 &  x293 &  x295 &  x296 &  x299 &  x301 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x328 &  x329 &  x332 &  x334 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x362 &  x365 &  x368 &  x373 &  x374 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x406 &  x412 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x445 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x467 &  x470 &  x473 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x556 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x584 &  x587 &  x590 &  x593 &  x595 &  x596 &  x599 &  x602 &  x608 &  x614 &  x617 &  x620 &  x626 &  x629 &  x632 &  x635 &  x638 &  x650 &  x653 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x820 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x842 &  x851 &  x854 &  x859 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x898 &  x901 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x940 &  x941 &  x944 &  x946 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 &  x1130 & ~x549 & ~x627;
assign c332 =  x2 &  x5 &  x11 &  x14 &  x17 &  x20 &  x23 &  x29 &  x32 &  x41 &  x44 &  x50 &  x53 &  x56 &  x62 &  x65 &  x68 &  x71 &  x73 &  x74 &  x80 &  x86 &  x89 &  x92 &  x100 &  x101 &  x110 &  x112 &  x113 &  x119 &  x122 &  x125 &  x128 &  x131 &  x140 &  x143 &  x146 &  x151 &  x152 &  x158 &  x164 &  x167 &  x170 &  x172 &  x176 &  x179 &  x182 &  x185 &  x191 &  x197 &  x203 &  x206 &  x209 &  x211 &  x212 &  x221 &  x224 &  x227 &  x230 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x269 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x302 &  x308 &  x311 &  x320 &  x323 &  x326 &  x329 &  x332 &  x341 &  x347 &  x350 &  x353 &  x356 &  x362 &  x368 &  x373 &  x374 &  x380 &  x383 &  x386 &  x389 &  x392 &  x398 &  x401 &  x407 &  x410 &  x413 &  x416 &  x422 &  x428 &  x431 &  x434 &  x437 &  x440 &  x445 &  x449 &  x451 &  x452 &  x461 &  x464 &  x467 &  x470 &  x476 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x509 &  x512 &  x515 &  x518 &  x524 &  x530 &  x533 &  x536 &  x542 &  x545 &  x548 &  x556 &  x557 &  x566 &  x569 &  x572 &  x581 &  x584 &  x586 &  x587 &  x590 &  x593 &  x595 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x625 &  x626 &  x629 &  x632 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x668 &  x671 &  x680 &  x683 &  x686 &  x703 &  x704 &  x707 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x746 &  x752 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x781 &  x782 &  x785 &  x788 &  x790 &  x791 &  x794 &  x797 &  x806 &  x812 &  x818 &  x820 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x859 &  x860 &  x862 &  x863 &  x866 &  x869 &  x875 &  x878 &  x884 &  x887 &  x890 &  x893 &  x896 &  x902 &  x905 &  x908 &  x911 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x977 &  x980 &  x986 &  x989 &  x992 &  x1007 &  x1010 &  x1013 &  x1022 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1055 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x123;
assign c334 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x35 &  x38 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x92 &  x95 &  x98 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x152 &  x158 &  x161 &  x167 &  x170 &  x173 &  x176 &  x179 &  x185 &  x191 &  x194 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x272 &  x275 &  x281 &  x284 &  x286 &  x287 &  x290 &  x293 &  x296 &  x299 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x325 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x362 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x386 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x428 &  x431 &  x434 &  x437 &  x440 &  x446 &  x449 &  x452 &  x455 &  x461 &  x464 &  x467 &  x473 &  x476 &  x479 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x527 &  x533 &  x536 &  x545 &  x548 &  x550 &  x551 &  x554 &  x557 &  x560 &  x563 &  x572 &  x575 &  x578 &  x584 &  x587 &  x589 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x628 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x667 &  x668 &  x671 &  x674 &  x677 &  x683 &  x686 &  x692 &  x695 &  x701 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x745 &  x746 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x836 &  x842 &  x845 &  x848 &  x851 &  x854 &  x862 &  x863 &  x866 &  x869 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x956 &  x959 &  x962 &  x965 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x39 & ~x42 & ~x78 & ~x81 & ~x117 & ~x159 & ~x195 & ~x234 & ~x378 & ~x417 & ~x687 & ~x1053 & ~x1092;
assign c336 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x38 &  x41 &  x44 &  x50 &  x52 &  x56 &  x65 &  x68 &  x77 &  x80 &  x83 &  x89 &  x95 &  x98 &  x101 &  x113 &  x116 &  x119 &  x121 &  x122 &  x125 &  x134 &  x137 &  x143 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x170 &  x182 &  x191 &  x203 &  x206 &  x209 &  x215 &  x218 &  x227 &  x230 &  x238 &  x239 &  x242 &  x245 &  x251 &  x254 &  x260 &  x263 &  x266 &  x269 &  x275 &  x277 &  x278 &  x281 &  x284 &  x287 &  x296 &  x299 &  x302 &  x308 &  x311 &  x314 &  x316 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x341 &  x344 &  x347 &  x350 &  x353 &  x355 &  x356 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x383 &  x389 &  x392 &  x394 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x416 &  x428 &  x431 &  x433 &  x434 &  x443 &  x449 &  x452 &  x461 &  x467 &  x470 &  x472 &  x473 &  x482 &  x485 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x524 &  x530 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x553 &  x554 &  x563 &  x569 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x614 &  x617 &  x623 &  x629 &  x632 &  x638 &  x641 &  x647 &  x650 &  x656 &  x659 &  x662 &  x668 &  x674 &  x677 &  x680 &  x683 &  x692 &  x695 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x728 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x797 &  x803 &  x806 &  x812 &  x818 &  x830 &  x833 &  x836 &  x839 &  x845 &  x848 &  x851 &  x854 &  x857 &  x863 &  x872 &  x875 &  x881 &  x890 &  x893 &  x899 &  x905 &  x908 &  x914 &  x917 &  x923 &  x929 &  x935 &  x938 &  x941 &  x944 &  x947 &  x953 &  x956 &  x959 &  x962 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1043 &  x1052 &  x1058 &  x1061 &  x1070 &  x1073 &  x1076 &  x1091 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1127 & ~x507 & ~x546 & ~x585 & ~x663 & ~x672 & ~x702 & ~x783 & ~x789 & ~x819 & ~x822 & ~x828 & ~x858 & ~x900 & ~x939 & ~x945;
assign c338 =  x5 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x86 &  x89 &  x92 &  x98 &  x104 &  x110 &  x113 &  x116 &  x119 &  x131 &  x137 &  x140 &  x149 &  x152 &  x158 &  x161 &  x164 &  x170 &  x179 &  x182 &  x185 &  x188 &  x197 &  x203 &  x206 &  x209 &  x218 &  x220 &  x224 &  x242 &  x245 &  x248 &  x254 &  x272 &  x275 &  x281 &  x284 &  x287 &  x293 &  x296 &  x305 &  x311 &  x320 &  x323 &  x338 &  x344 &  x350 &  x362 &  x365 &  x368 &  x370 &  x377 &  x380 &  x386 &  x389 &  x407 &  x410 &  x425 &  x428 &  x431 &  x434 &  x440 &  x446 &  x449 &  x452 &  x455 &  x461 &  x467 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x497 &  x500 &  x503 &  x509 &  x512 &  x515 &  x518 &  x527 &  x533 &  x536 &  x539 &  x545 &  x548 &  x554 &  x557 &  x560 &  x566 &  x578 &  x584 &  x596 &  x602 &  x605 &  x611 &  x620 &  x623 &  x629 &  x632 &  x638 &  x641 &  x647 &  x650 &  x656 &  x668 &  x674 &  x680 &  x683 &  x686 &  x689 &  x695 &  x698 &  x706 &  x707 &  x716 &  x719 &  x725 &  x734 &  x743 &  x752 &  x755 &  x758 &  x761 &  x770 &  x773 &  x776 &  x779 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x827 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x857 &  x872 &  x878 &  x881 &  x887 &  x890 &  x893 &  x896 &  x899 &  x914 &  x917 &  x920 &  x929 &  x944 &  x947 &  x950 &  x965 &  x971 &  x974 &  x980 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1052 &  x1058 &  x1061 &  x1073 &  x1088 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 & ~x33 & ~x39 & ~x48 & ~x87 & ~x117 & ~x126 & ~x156 & ~x234 & ~x423 & ~x768 & ~x969 & ~x1074 & ~x1113;
assign c340 =  x5 &  x8 &  x11 &  x17 &  x20 &  x23 &  x26 &  x29 &  x35 &  x38 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x65 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x113 &  x119 &  x122 &  x128 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x188 &  x191 &  x193 &  x194 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x224 &  x230 &  x233 &  x239 &  x245 &  x248 &  x251 &  x254 &  x257 &  x263 &  x266 &  x272 &  x275 &  x281 &  x284 &  x286 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x308 &  x314 &  x320 &  x323 &  x325 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x362 &  x363 &  x364 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x389 &  x392 &  x395 &  x398 &  x407 &  x410 &  x419 &  x422 &  x428 &  x431 &  x434 &  x440 &  x446 &  x461 &  x464 &  x467 &  x470 &  x473 &  x479 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x527 &  x530 &  x536 &  x539 &  x545 &  x551 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x632 &  x635 &  x638 &  x644 &  x647 &  x650 &  x653 &  x662 &  x668 &  x674 &  x677 &  x683 &  x686 &  x689 &  x695 &  x701 &  x704 &  x707 &  x713 &  x716 &  x722 &  x725 &  x728 &  x740 &  x743 &  x746 &  x752 &  x755 &  x761 &  x770 &  x773 &  x776 &  x784 &  x785 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x823 &  x830 &  x833 &  x836 &  x839 &  x848 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x881 &  x884 &  x887 &  x890 &  x893 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x941 &  x944 &  x947 &  x953 &  x959 &  x962 &  x965 &  x968 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1078 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1118 &  x1121 &  x1124 &  x1130 & ~x0 & ~x117 & ~x156 & ~x195 & ~x234 & ~x312 & ~x795 & ~x834 & ~x975 & ~x1014 & ~x1053 & ~x1092;
assign c342 =  x5 &  x8 &  x11 &  x23 &  x32 &  x35 &  x41 &  x44 &  x53 &  x62 &  x65 &  x71 &  x77 &  x86 &  x92 &  x110 &  x116 &  x119 &  x140 &  x143 &  x149 &  x152 &  x167 &  x176 &  x188 &  x191 &  x197 &  x200 &  x203 &  x221 &  x224 &  x233 &  x248 &  x251 &  x269 &  x272 &  x277 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x308 &  x314 &  x316 &  x329 &  x355 &  x356 &  x365 &  x371 &  x380 &  x389 &  x392 &  x393 &  x398 &  x401 &  x413 &  x419 &  x425 &  x431 &  x432 &  x440 &  x443 &  x446 &  x458 &  x461 &  x464 &  x476 &  x488 &  x494 &  x497 &  x500 &  x503 &  x509 &  x515 &  x530 &  x533 &  x539 &  x542 &  x550 &  x557 &  x563 &  x572 &  x575 &  x581 &  x590 &  x593 &  x599 &  x608 &  x611 &  x626 &  x629 &  x635 &  x644 &  x650 &  x656 &  x659 &  x665 &  x668 &  x670 &  x674 &  x683 &  x686 &  x704 &  x707 &  x709 &  x710 &  x713 &  x722 &  x725 &  x728 &  x734 &  x740 &  x743 &  x746 &  x758 &  x773 &  x779 &  x782 &  x788 &  x800 &  x803 &  x809 &  x818 &  x824 &  x827 &  x830 &  x833 &  x836 &  x845 &  x863 &  x875 &  x878 &  x890 &  x893 &  x902 &  x922 &  x926 &  x932 &  x935 &  x941 &  x947 &  x961 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1019 &  x1025 &  x1034 &  x1043 &  x1055 &  x1058 &  x1070 &  x1073 &  x1082 &  x1094 &  x1097 &  x1100 &  x1106 &  x1118 &  x1124 &  x1127 & ~x261 & ~x600 & ~x702 & ~x741 & ~x756 & ~x819 & ~x840 & ~x891 & ~x1053;
assign c344 =  x11 &  x14 &  x23 &  x29 &  x32 &  x35 &  x38 &  x59 &  x65 &  x68 &  x77 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x107 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x146 &  x149 &  x152 &  x155 &  x158 &  x164 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x251 &  x254 &  x257 &  x266 &  x269 &  x277 &  x284 &  x286 &  x302 &  x305 &  x308 &  x311 &  x314 &  x316 &  x317 &  x320 &  x326 &  x329 &  x335 &  x338 &  x341 &  x362 &  x371 &  x377 &  x395 &  x401 &  x404 &  x407 &  x410 &  x413 &  x431 &  x433 &  x437 &  x446 &  x449 &  x452 &  x455 &  x464 &  x467 &  x470 &  x476 &  x488 &  x491 &  x497 &  x500 &  x506 &  x512 &  x515 &  x518 &  x527 &  x536 &  x542 &  x545 &  x550 &  x551 &  x554 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x584 &  x587 &  x596 &  x599 &  x602 &  x605 &  x608 &  x617 &  x620 &  x623 &  x626 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x667 &  x668 &  x674 &  x680 &  x683 &  x689 &  x695 &  x701 &  x706 &  x713 &  x722 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x752 &  x755 &  x758 &  x767 &  x773 &  x776 &  x785 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x818 &  x821 &  x824 &  x830 &  x833 &  x836 &  x842 &  x848 &  x851 &  x854 &  x857 &  x866 &  x869 &  x872 &  x878 &  x881 &  x899 &  x902 &  x905 &  x908 &  x911 &  x917 &  x920 &  x923 &  x929 &  x932 &  x938 &  x941 &  x947 &  x965 &  x974 &  x977 &  x986 &  x989 &  x998 &  x1001 &  x1007 &  x1010 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1052 &  x1058 &  x1061 &  x1067 &  x1076 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1127 &  x1130 & ~x342 & ~x381 & ~x420 & ~x421 & ~x459 & ~x498 & ~x499 & ~x576 & ~x600;
assign c346 =  x1 &  x5 &  x8 &  x11 &  x23 &  x26 &  x35 &  x38 &  x44 &  x47 &  x50 &  x65 &  x68 &  x71 &  x80 &  x95 &  x98 &  x107 &  x110 &  x113 &  x119 &  x125 &  x131 &  x140 &  x143 &  x152 &  x155 &  x158 &  x161 &  x167 &  x173 &  x182 &  x194 &  x197 &  x200 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x242 &  x245 &  x248 &  x251 &  x257 &  x272 &  x281 &  x284 &  x290 &  x293 &  x296 &  x302 &  x326 &  x329 &  x332 &  x335 &  x344 &  x347 &  x353 &  x355 &  x356 &  x359 &  x362 &  x371 &  x374 &  x377 &  x383 &  x386 &  x389 &  x391 &  x394 &  x395 &  x398 &  x410 &  x416 &  x422 &  x433 &  x437 &  x443 &  x446 &  x449 &  x452 &  x458 &  x461 &  x464 &  x467 &  x470 &  x472 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x503 &  x506 &  x511 &  x512 &  x518 &  x527 &  x536 &  x542 &  x554 &  x557 &  x560 &  x566 &  x572 &  x578 &  x581 &  x593 &  x596 &  x608 &  x614 &  x623 &  x629 &  x632 &  x635 &  x638 &  x641 &  x647 &  x659 &  x662 &  x668 &  x671 &  x677 &  x680 &  x683 &  x704 &  x722 &  x731 &  x740 &  x743 &  x755 &  x758 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x785 &  x788 &  x797 &  x800 &  x803 &  x809 &  x812 &  x814 &  x821 &  x830 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x857 &  x860 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x893 &  x896 &  x905 &  x911 &  x917 &  x920 &  x925 &  x926 &  x935 &  x938 &  x941 &  x953 &  x959 &  x965 &  x968 &  x970 &  x977 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1016 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1055 &  x1064 &  x1070 &  x1088 &  x1097 &  x1103 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x45 & ~x84 & ~x123 & ~x240 & ~x252;
assign c348 =  x11 &  x14 &  x17 &  x20 &  x26 &  x29 &  x35 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x74 &  x92 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x122 &  x131 &  x137 &  x149 &  x152 &  x158 &  x179 &  x188 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x230 &  x233 &  x245 &  x251 &  x254 &  x260 &  x275 &  x281 &  x284 &  x293 &  x299 &  x302 &  x305 &  x317 &  x326 &  x329 &  x332 &  x335 &  x347 &  x356 &  x362 &  x365 &  x371 &  x380 &  x386 &  x395 &  x401 &  x404 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x446 &  x452 &  x458 &  x473 &  x479 &  x482 &  x488 &  x491 &  x500 &  x518 &  x527 &  x530 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x557 &  x563 &  x566 &  x575 &  x581 &  x589 &  x590 &  x593 &  x599 &  x617 &  x623 &  x626 &  x632 &  x638 &  x641 &  x644 &  x653 &  x659 &  x662 &  x664 &  x668 &  x677 &  x686 &  x692 &  x703 &  x704 &  x706 &  x710 &  x713 &  x716 &  x734 &  x737 &  x752 &  x761 &  x770 &  x779 &  x781 &  x782 &  x785 &  x794 &  x797 &  x803 &  x812 &  x815 &  x836 &  x839 &  x842 &  x848 &  x851 &  x857 &  x860 &  x863 &  x866 &  x869 &  x878 &  x887 &  x890 &  x893 &  x896 &  x898 &  x899 &  x901 &  x905 &  x908 &  x920 &  x929 &  x935 &  x938 &  x947 &  x953 &  x962 &  x965 &  x968 &  x971 &  x977 &  x980 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1073 &  x1085 &  x1088 &  x1094 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 & ~x609 & ~x669 & ~x795 & ~x834 & ~x835 & ~x1104;
assign c350 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x38 &  x44 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x77 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x113 &  x116 &  x119 &  x125 &  x131 &  x137 &  x140 &  x143 &  x146 &  x149 &  x155 &  x161 &  x164 &  x167 &  x170 &  x173 &  x179 &  x182 &  x185 &  x191 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x275 &  x278 &  x284 &  x287 &  x290 &  x298 &  x299 &  x302 &  x305 &  x311 &  x314 &  x317 &  x320 &  x323 &  x335 &  x337 &  x338 &  x341 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x376 &  x377 &  x383 &  x392 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x434 &  x436 &  x437 &  x439 &  x440 &  x441 &  x442 &  x443 &  x446 &  x449 &  x455 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x481 &  x485 &  x491 &  x494 &  x497 &  x500 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x523 &  x524 &  x527 &  x530 &  x533 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x560 &  x563 &  x569 &  x575 &  x578 &  x581 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x626 &  x629 &  x632 &  x638 &  x641 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x680 &  x683 &  x689 &  x692 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x722 &  x728 &  x731 &  x734 &  x737 &  x740 &  x746 &  x749 &  x755 &  x764 &  x773 &  x776 &  x779 &  x788 &  x791 &  x797 &  x800 &  x806 &  x809 &  x815 &  x824 &  x827 &  x830 &  x833 &  x839 &  x845 &  x848 &  x854 &  x857 &  x866 &  x869 &  x875 &  x881 &  x884 &  x887 &  x890 &  x896 &  x899 &  x905 &  x908 &  x911 &  x914 &  x920 &  x923 &  x926 &  x929 &  x932 &  x941 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x980 &  x986 &  x989 &  x992 &  x1001 &  x1004 &  x1010 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1097 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x351 & ~x390 & ~x429 & ~x468 & ~x507 & ~x975 & ~x1014 & ~x1053 & ~x1092;
assign c352 =  x5 &  x14 &  x17 &  x26 &  x44 &  x47 &  x53 &  x56 &  x62 &  x65 &  x68 &  x74 &  x77 &  x83 &  x86 &  x89 &  x92 &  x95 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x131 &  x134 &  x136 &  x137 &  x143 &  x146 &  x149 &  x152 &  x155 &  x164 &  x170 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x212 &  x214 &  x215 &  x221 &  x230 &  x242 &  x248 &  x254 &  x257 &  x263 &  x269 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x305 &  x311 &  x314 &  x320 &  x329 &  x331 &  x332 &  x335 &  x338 &  x341 &  x347 &  x353 &  x356 &  x359 &  x365 &  x370 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x422 &  x428 &  x431 &  x443 &  x449 &  x452 &  x455 &  x458 &  x464 &  x467 &  x470 &  x485 &  x488 &  x491 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x563 &  x566 &  x575 &  x578 &  x587 &  x590 &  x596 &  x605 &  x608 &  x614 &  x617 &  x623 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x659 &  x665 &  x668 &  x674 &  x683 &  x686 &  x692 &  x698 &  x701 &  x710 &  x713 &  x725 &  x731 &  x737 &  x740 &  x743 &  x749 &  x751 &  x752 &  x755 &  x770 &  x776 &  x782 &  x784 &  x790 &  x791 &  x797 &  x800 &  x806 &  x812 &  x818 &  x821 &  x823 &  x824 &  x827 &  x829 &  x830 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x866 &  x869 &  x872 &  x881 &  x884 &  x887 &  x890 &  x899 &  x902 &  x905 &  x907 &  x911 &  x914 &  x917 &  x923 &  x929 &  x932 &  x935 &  x941 &  x944 &  x950 &  x953 &  x962 &  x965 &  x968 &  x971 &  x974 &  x982 &  x986 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1025 &  x1031 &  x1034 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1061 &  x1067 &  x1073 &  x1079 &  x1085 &  x1088 &  x1091 &  x1097 &  x1099 &  x1100 &  x1106 &  x1109 &  x1115 &  x1127 & ~x111 & ~x117 & ~x156 & ~x273 & ~x312;
assign c354 =  x23 &  x29 &  x32 &  x35 &  x38 &  x47 &  x56 &  x65 &  x80 &  x92 &  x95 &  x110 &  x116 &  x122 &  x125 &  x133 &  x143 &  x167 &  x172 &  x176 &  x182 &  x184 &  x185 &  x188 &  x194 &  x197 &  x221 &  x223 &  x227 &  x230 &  x236 &  x242 &  x245 &  x248 &  x251 &  x254 &  x256 &  x257 &  x259 &  x263 &  x269 &  x275 &  x281 &  x287 &  x293 &  x296 &  x302 &  x305 &  x307 &  x308 &  x314 &  x323 &  x328 &  x334 &  x335 &  x338 &  x341 &  x350 &  x371 &  x374 &  x380 &  x386 &  x389 &  x392 &  x395 &  x401 &  x403 &  x404 &  x407 &  x416 &  x425 &  x440 &  x442 &  x446 &  x452 &  x458 &  x461 &  x470 &  x473 &  x479 &  x485 &  x506 &  x509 &  x512 &  x521 &  x524 &  x545 &  x551 &  x557 &  x566 &  x569 &  x575 &  x581 &  x584 &  x590 &  x605 &  x608 &  x614 &  x617 &  x632 &  x638 &  x641 &  x644 &  x650 &  x671 &  x680 &  x683 &  x686 &  x695 &  x698 &  x701 &  x719 &  x722 &  x731 &  x743 &  x746 &  x752 &  x758 &  x767 &  x779 &  x781 &  x782 &  x785 &  x791 &  x794 &  x806 &  x812 &  x823 &  x824 &  x833 &  x836 &  x842 &  x851 &  x859 &  x862 &  x872 &  x875 &  x878 &  x884 &  x893 &  x898 &  x901 &  x911 &  x920 &  x929 &  x932 &  x937 &  x938 &  x941 &  x947 &  x965 &  x968 &  x971 &  x976 &  x989 &  x1001 &  x1018 &  x1019 &  x1031 &  x1034 &  x1040 &  x1043 &  x1049 &  x1055 &  x1064 &  x1070 &  x1076 &  x1094 &  x1103 &  x1118 &  x1121 & ~x201;
assign c356 =  x5 &  x8 &  x11 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x47 &  x50 &  x53 &  x56 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x95 &  x98 &  x101 &  x104 &  x107 &  x113 &  x119 &  x122 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x203 &  x206 &  x209 &  x212 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x314 &  x317 &  x320 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x350 &  x353 &  x356 &  x359 &  x365 &  x368 &  x374 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x407 &  x409 &  x410 &  x413 &  x416 &  x428 &  x434 &  x437 &  x446 &  x449 &  x452 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x485 &  x488 &  x491 &  x500 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x673 &  x674 &  x677 &  x683 &  x686 &  x692 &  x698 &  x701 &  x704 &  x707 &  x710 &  x712 &  x713 &  x716 &  x719 &  x722 &  x725 &  x731 &  x734 &  x737 &  x740 &  x746 &  x751 &  x752 &  x755 &  x758 &  x761 &  x764 &  x770 &  x772 &  x776 &  x779 &  x782 &  x788 &  x790 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x811 &  x812 &  x818 &  x820 &  x824 &  x827 &  x829 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x857 &  x860 &  x863 &  x868 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x977 &  x980 &  x986 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1121 &  x1124 &  x1127 & ~x159 & ~x198 & ~x237 & ~x276 & ~x315 & ~x393 & ~x471;
assign c358 =  x2 &  x5 &  x8 &  x17 &  x20 &  x23 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x167 &  x170 &  x173 &  x176 &  x178 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x275 &  x278 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x341 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x524 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x571 &  x572 &  x575 &  x578 &  x581 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x665 &  x668 &  x670 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x698 &  x701 &  x704 &  x707 &  x709 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x6 & ~x69 & ~x1005 & ~x1044 & ~x1062 & ~x1089 & ~x1101;
assign c360 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x128 &  x134 &  x137 &  x146 &  x149 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x206 &  x209 &  x212 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x356 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x448 &  x449 &  x452 &  x455 &  x457 &  x458 &  x461 &  x464 &  x467 &  x473 &  x476 &  x479 &  x482 &  x485 &  x487 &  x488 &  x491 &  x494 &  x496 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x524 &  x526 &  x527 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x559 &  x560 &  x563 &  x565 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x598 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x629 &  x632 &  x638 &  x641 &  x643 &  x644 &  x647 &  x650 &  x653 &  x656 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x682 &  x683 &  x686 &  x689 &  x692 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x806 &  x809 &  x812 &  x815 &  x820 &  x821 &  x823 &  x824 &  x833 &  x836 &  x839 &  x845 &  x848 &  x851 &  x854 &  x857 &  x859 &  x860 &  x862 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x896 &  x898 &  x901 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x937 &  x938 &  x940 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x962 &  x965 &  x968 &  x971 &  x974 &  x976 &  x977 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1015 &  x1016 &  x1018 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1054 &  x1057 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1093 &  x1094 &  x1096 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x351 & ~x843 & ~x882;
assign c362 =  x2 &  x5 &  x8 &  x17 &  x26 &  x38 &  x53 &  x56 &  x65 &  x77 &  x98 &  x107 &  x119 &  x125 &  x128 &  x131 &  x146 &  x155 &  x161 &  x173 &  x188 &  x212 &  x242 &  x245 &  x254 &  x260 &  x263 &  x275 &  x284 &  x287 &  x302 &  x305 &  x311 &  x338 &  x359 &  x377 &  x380 &  x386 &  x398 &  x419 &  x425 &  x440 &  x458 &  x464 &  x470 &  x476 &  x488 &  x491 &  x563 &  x572 &  x581 &  x584 &  x596 &  x620 &  x632 &  x656 &  x674 &  x677 &  x701 &  x704 &  x716 &  x728 &  x737 &  x755 &  x758 &  x767 &  x770 &  x797 &  x812 &  x821 &  x836 &  x845 &  x848 &  x851 &  x863 &  x872 &  x878 &  x884 &  x899 &  x901 &  x911 &  x914 &  x929 &  x932 &  x935 &  x986 &  x1007 &  x1025 &  x1028 &  x1037 &  x1046 &  x1052 &  x1064 &  x1079 &  x1085 &  x1103 &  x1109 &  x1124 &  x1130 & ~x30 & ~x795 & ~x796 & ~x804 & ~x835 & ~x843 & ~x873 & ~x990 & ~x1035;
assign c364 =  x2 &  x4 &  x26 &  x32 &  x35 &  x38 &  x40 &  x50 &  x53 &  x59 &  x65 &  x68 &  x80 &  x104 &  x107 &  x113 &  x116 &  x128 &  x149 &  x152 &  x155 &  x157 &  x161 &  x164 &  x170 &  x173 &  x179 &  x182 &  x188 &  x194 &  x200 &  x209 &  x212 &  x215 &  x224 &  x245 &  x251 &  x254 &  x257 &  x263 &  x266 &  x269 &  x275 &  x277 &  x281 &  x287 &  x290 &  x296 &  x314 &  x317 &  x326 &  x329 &  x332 &  x335 &  x344 &  x347 &  x350 &  x353 &  x362 &  x365 &  x371 &  x401 &  x404 &  x416 &  x419 &  x428 &  x431 &  x434 &  x437 &  x440 &  x446 &  x449 &  x464 &  x467 &  x473 &  x479 &  x503 &  x509 &  x512 &  x518 &  x524 &  x527 &  x533 &  x536 &  x539 &  x542 &  x545 &  x551 &  x563 &  x566 &  x569 &  x575 &  x578 &  x587 &  x608 &  x620 &  x629 &  x644 &  x647 &  x650 &  x656 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x689 &  x701 &  x704 &  x707 &  x713 &  x719 &  x746 &  x749 &  x755 &  x758 &  x767 &  x776 &  x800 &  x803 &  x809 &  x824 &  x827 &  x835 &  x839 &  x844 &  x845 &  x848 &  x857 &  x869 &  x881 &  x887 &  x893 &  x896 &  x902 &  x911 &  x914 &  x932 &  x944 &  x950 &  x953 &  x956 &  x962 &  x965 &  x968 &  x971 &  x977 &  x980 &  x986 &  x992 &  x998 &  x1001 &  x1004 &  x1019 &  x1024 &  x1031 &  x1037 &  x1040 &  x1043 &  x1052 &  x1070 &  x1085 &  x1088 &  x1091 &  x1097 &  x1130 & ~x141 & ~x309 & ~x348 & ~x624;
assign c366 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x65 &  x71 &  x77 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x188 &  x191 &  x200 &  x206 &  x209 &  x212 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x260 &  x263 &  x269 &  x272 &  x275 &  x278 &  x281 &  x287 &  x289 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x353 &  x356 &  x362 &  x364 &  x365 &  x368 &  x371 &  x374 &  x377 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x403 &  x404 &  x410 &  x413 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x442 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x547 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x584 &  x586 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x625 &  x626 &  x632 &  x635 &  x638 &  x641 &  x647 &  x650 &  x653 &  x659 &  x664 &  x665 &  x668 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x698 &  x701 &  x703 &  x707 &  x710 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x737 &  x740 &  x742 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x770 &  x773 &  x776 &  x779 &  x781 &  x782 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x851 &  x854 &  x857 &  x859 &  x862 &  x863 &  x866 &  x872 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x901 &  x902 &  x905 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x940 &  x941 &  x943 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1055 &  x1058 &  x1061 &  x1064 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x570 & ~x609 & ~x675 & ~x714 & ~x753 & ~x792;
assign c368 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x131 &  x137 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x167 &  x168 &  x169 &  x170 &  x173 &  x182 &  x185 &  x188 &  x194 &  x197 &  x200 &  x205 &  x206 &  x208 &  x209 &  x212 &  x215 &  x218 &  x221 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x391 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x470 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x503 &  x506 &  x509 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x542 &  x545 &  x548 &  x550 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x589 &  x593 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x628 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x748 &  x749 &  x752 &  x755 &  x758 &  x761 &  x767 &  x770 &  x773 &  x779 &  x782 &  x785 &  x787 &  x788 &  x791 &  x794 &  x797 &  x800 &  x806 &  x809 &  x812 &  x815 &  x818 &  x824 &  x826 &  x827 &  x830 &  x833 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1004 &  x1007 &  x1010 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x117 & ~x483 & ~x522 & ~x561 & ~x780;
assign c370 =  x8 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x53 &  x56 &  x59 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x130 &  x131 &  x134 &  x137 &  x140 &  x143 &  x149 &  x155 &  x158 &  x161 &  x164 &  x167 &  x169 &  x170 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x207 &  x208 &  x209 &  x212 &  x215 &  x218 &  x224 &  x227 &  x236 &  x238 &  x239 &  x248 &  x251 &  x254 &  x257 &  x266 &  x269 &  x272 &  x275 &  x277 &  x278 &  x281 &  x287 &  x290 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x316 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x344 &  x350 &  x352 &  x353 &  x355 &  x359 &  x365 &  x368 &  x377 &  x383 &  x392 &  x394 &  x395 &  x398 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x433 &  x434 &  x437 &  x443 &  x446 &  x449 &  x452 &  x458 &  x461 &  x464 &  x467 &  x470 &  x472 &  x473 &  x476 &  x482 &  x485 &  x491 &  x494 &  x497 &  x503 &  x506 &  x509 &  x511 &  x512 &  x515 &  x518 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x550 &  x554 &  x557 &  x560 &  x572 &  x578 &  x587 &  x590 &  x596 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x632 &  x635 &  x638 &  x641 &  x647 &  x650 &  x653 &  x656 &  x662 &  x671 &  x674 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x740 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x776 &  x779 &  x782 &  x797 &  x806 &  x812 &  x818 &  x821 &  x826 &  x827 &  x833 &  x839 &  x842 &  x848 &  x854 &  x857 &  x860 &  x865 &  x869 &  x872 &  x875 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x941 &  x944 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x971 &  x974 &  x977 &  x983 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1028 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 & ~x357 & ~x366 & ~x444 & ~x483 & ~x522 & ~x561 & ~x600;
assign c372 =  x5 &  x8 &  x11 &  x62 &  x65 &  x80 &  x83 &  x86 &  x89 &  x98 &  x104 &  x107 &  x121 &  x122 &  x125 &  x128 &  x134 &  x152 &  x158 &  x164 &  x167 &  x170 &  x173 &  x179 &  x182 &  x188 &  x194 &  x197 &  x199 &  x200 &  x203 &  x209 &  x221 &  x227 &  x238 &  x239 &  x242 &  x251 &  x257 &  x269 &  x277 &  x278 &  x281 &  x284 &  x290 &  x314 &  x316 &  x317 &  x326 &  x329 &  x332 &  x338 &  x341 &  x350 &  x353 &  x355 &  x356 &  x362 &  x377 &  x386 &  x394 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x431 &  x433 &  x434 &  x437 &  x443 &  x446 &  x452 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x500 &  x503 &  x521 &  x530 &  x536 &  x539 &  x542 &  x551 &  x557 &  x560 &  x566 &  x569 &  x572 &  x575 &  x599 &  x605 &  x608 &  x617 &  x620 &  x623 &  x626 &  x632 &  x635 &  x653 &  x659 &  x677 &  x695 &  x698 &  x704 &  x716 &  x725 &  x728 &  x731 &  x737 &  x746 &  x758 &  x764 &  x767 &  x770 &  x779 &  x794 &  x809 &  x812 &  x821 &  x827 &  x836 &  x839 &  x844 &  x860 &  x866 &  x869 &  x872 &  x875 &  x878 &  x884 &  x893 &  x902 &  x914 &  x922 &  x923 &  x926 &  x929 &  x935 &  x950 &  x956 &  x961 &  x968 &  x974 &  x977 &  x980 &  x983 &  x989 &  x995 &  x998 &  x1000 &  x1001 &  x1007 &  x1010 &  x1016 &  x1034 &  x1037 &  x1040 &  x1043 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1082 &  x1088 &  x1094 &  x1100 &  x1109 &  x1117 &  x1118 &  x1121 &  x1127 & ~x300 & ~x522 & ~x561 & ~x639 & ~x702 & ~x741 & ~x900 & ~x936 & ~x939 & ~x975 & ~x1014 & ~x1053 & ~x1056 & ~x1092;
assign c374 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x38 &  x44 &  x47 &  x59 &  x62 &  x71 &  x86 &  x95 &  x98 &  x101 &  x107 &  x110 &  x113 &  x116 &  x122 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x155 &  x158 &  x167 &  x170 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x212 &  x227 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x251 &  x257 &  x260 &  x278 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x317 &  x320 &  x321 &  x322 &  x326 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x355 &  x359 &  x361 &  x371 &  x377 &  x383 &  x386 &  x391 &  x392 &  x394 &  x395 &  x398 &  x404 &  x410 &  x413 &  x416 &  x425 &  x430 &  x433 &  x440 &  x446 &  x455 &  x458 &  x464 &  x467 &  x469 &  x472 &  x473 &  x482 &  x485 &  x491 &  x497 &  x503 &  x506 &  x509 &  x518 &  x524 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x589 &  x593 &  x595 &  x608 &  x611 &  x617 &  x623 &  x628 &  x629 &  x635 &  x638 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x716 &  x731 &  x737 &  x749 &  x752 &  x758 &  x761 &  x764 &  x773 &  x776 &  x782 &  x785 &  x788 &  x794 &  x797 &  x803 &  x809 &  x812 &  x821 &  x824 &  x826 &  x827 &  x830 &  x836 &  x839 &  x848 &  x851 &  x860 &  x863 &  x866 &  x875 &  x890 &  x893 &  x899 &  x902 &  x905 &  x908 &  x911 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x971 &  x974 &  x977 &  x980 &  x989 &  x995 &  x998 &  x1007 &  x1013 &  x1016 &  x1019 &  x1025 &  x1031 &  x1034 &  x1043 &  x1055 &  x1067 &  x1070 &  x1073 &  x1082 &  x1085 &  x1097 &  x1100 &  x1106 &  x1112 &  x1115 &  x1121 & ~x435 & ~x492 & ~x600;
assign c376 =  x2 &  x5 &  x8 &  x10 &  x11 &  x14 &  x17 &  x23 &  x29 &  x32 &  x35 &  x41 &  x47 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x80 &  x104 &  x113 &  x119 &  x125 &  x134 &  x140 &  x143 &  x152 &  x155 &  x161 &  x167 &  x170 &  x173 &  x179 &  x182 &  x200 &  x203 &  x206 &  x215 &  x227 &  x233 &  x245 &  x251 &  x260 &  x263 &  x266 &  x272 &  x275 &  x277 &  x278 &  x284 &  x287 &  x290 &  x296 &  x302 &  x317 &  x329 &  x350 &  x356 &  x365 &  x374 &  x377 &  x383 &  x386 &  x401 &  x416 &  x419 &  x425 &  x431 &  x433 &  x437 &  x443 &  x446 &  x449 &  x452 &  x458 &  x461 &  x467 &  x476 &  x485 &  x488 &  x494 &  x497 &  x506 &  x515 &  x518 &  x524 &  x527 &  x533 &  x539 &  x545 &  x548 &  x551 &  x557 &  x563 &  x572 &  x590 &  x592 &  x593 &  x599 &  x608 &  x611 &  x614 &  x617 &  x631 &  x635 &  x641 &  x644 &  x647 &  x650 &  x656 &  x662 &  x670 &  x671 &  x674 &  x677 &  x686 &  x692 &  x694 &  x701 &  x719 &  x722 &  x725 &  x728 &  x731 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x767 &  x770 &  x772 &  x773 &  x776 &  x788 &  x800 &  x809 &  x812 &  x821 &  x824 &  x826 &  x830 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x860 &  x869 &  x878 &  x881 &  x905 &  x917 &  x920 &  x929 &  x938 &  x944 &  x947 &  x956 &  x959 &  x962 &  x965 &  x986 &  x992 &  x1001 &  x1007 &  x1013 &  x1022 &  x1025 &  x1028 &  x1034 &  x1040 &  x1046 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1124 & ~x483 & ~x522 & ~x663 & ~x741 & ~x819 & ~x858 & ~x897 & ~x936 & ~x978 & ~x1014 & ~x1017 & ~x1092 & ~x1095;
assign c378 =  x5 &  x8 &  x26 &  x35 &  x41 &  x44 &  x59 &  x71 &  x80 &  x83 &  x95 &  x98 &  x104 &  x110 &  x119 &  x122 &  x128 &  x137 &  x140 &  x143 &  x146 &  x158 &  x161 &  x170 &  x176 &  x179 &  x182 &  x191 &  x197 &  x200 &  x203 &  x206 &  x212 &  x218 &  x224 &  x227 &  x230 &  x236 &  x242 &  x245 &  x251 &  x254 &  x257 &  x260 &  x263 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x343 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x365 &  x371 &  x377 &  x383 &  x386 &  x389 &  x392 &  x407 &  x409 &  x413 &  x416 &  x419 &  x422 &  x425 &  x434 &  x449 &  x452 &  x455 &  x461 &  x467 &  x470 &  x482 &  x487 &  x488 &  x494 &  x500 &  x503 &  x515 &  x520 &  x527 &  x530 &  x542 &  x557 &  x559 &  x565 &  x569 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x608 &  x617 &  x623 &  x626 &  x635 &  x638 &  x641 &  x643 &  x647 &  x650 &  x653 &  x665 &  x668 &  x674 &  x677 &  x680 &  x689 &  x698 &  x701 &  x707 &  x710 &  x713 &  x719 &  x728 &  x734 &  x740 &  x746 &  x749 &  x752 &  x755 &  x761 &  x764 &  x770 &  x776 &  x779 &  x781 &  x782 &  x785 &  x791 &  x800 &  x806 &  x809 &  x812 &  x815 &  x821 &  x824 &  x830 &  x836 &  x839 &  x845 &  x848 &  x851 &  x857 &  x860 &  x862 &  x863 &  x866 &  x875 &  x878 &  x884 &  x896 &  x898 &  x899 &  x901 &  x911 &  x917 &  x920 &  x932 &  x935 &  x937 &  x938 &  x947 &  x950 &  x959 &  x971 &  x974 &  x976 &  x977 &  x979 &  x980 &  x985 &  x986 &  x989 &  x992 &  x998 &  x1007 &  x1016 &  x1018 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1049 &  x1057 &  x1058 &  x1064 &  x1067 &  x1070 &  x1082 &  x1088 &  x1094 &  x1097 &  x1100 &  x1106 &  x1112 &  x1115 &  x1118 &  x1130 & ~x354 & ~x687 & ~x747 & ~x873;
assign c380 =  x2 &  x5 &  x8 &  x11 &  x17 &  x20 &  x23 &  x29 &  x35 &  x38 &  x47 &  x53 &  x56 &  x62 &  x65 &  x74 &  x77 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x119 &  x122 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x185 &  x191 &  x194 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x239 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x284 &  x290 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x397 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x467 &  x473 &  x476 &  x479 &  x485 &  x488 &  x494 &  x497 &  x500 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x538 &  x542 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x575 &  x577 &  x581 &  x584 &  x587 &  x590 &  x593 &  x599 &  x602 &  x605 &  x608 &  x611 &  x613 &  x615 &  x616 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x652 &  x653 &  x655 &  x656 &  x659 &  x662 &  x668 &  x671 &  x674 &  x680 &  x686 &  x689 &  x691 &  x692 &  x694 &  x698 &  x701 &  x704 &  x707 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x739 &  x743 &  x746 &  x749 &  x752 &  x755 &  x761 &  x764 &  x770 &  x773 &  x776 &  x778 &  x779 &  x782 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x817 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x851 &  x854 &  x856 &  x857 &  x860 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x908 &  x914 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x980 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x429 & ~x468;
assign c382 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x167 &  x173 &  x176 &  x179 &  x182 &  x185 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x263 &  x266 &  x269 &  x272 &  x275 &  x281 &  x284 &  x286 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x325 &  x326 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x364 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x403 &  x404 &  x410 &  x413 &  x416 &  x422 &  x433 &  x434 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x464 &  x467 &  x473 &  x482 &  x485 &  x488 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x527 &  x530 &  x539 &  x542 &  x545 &  x547 &  x548 &  x551 &  x554 &  x557 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x584 &  x586 &  x587 &  x590 &  x593 &  x596 &  x599 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x625 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x662 &  x664 &  x665 &  x671 &  x674 &  x677 &  x680 &  x683 &  x692 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x784 &  x785 &  x791 &  x794 &  x797 &  x800 &  x809 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x854 &  x860 &  x862 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x890 &  x899 &  x902 &  x908 &  x911 &  x914 &  x926 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x971 &  x977 &  x980 &  x986 &  x989 &  x992 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1021 &  x1022 &  x1025 &  x1028 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1091 &  x1094 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x234 & ~x273 & ~x552 & ~x609 & ~x648;
assign c384 =  x8 &  x11 &  x26 &  x41 &  x65 &  x68 &  x71 &  x88 &  x92 &  x101 &  x107 &  x113 &  x122 &  x127 &  x128 &  x131 &  x143 &  x155 &  x170 &  x182 &  x191 &  x205 &  x206 &  x209 &  x218 &  x221 &  x224 &  x230 &  x233 &  x239 &  x244 &  x245 &  x257 &  x266 &  x278 &  x281 &  x283 &  x305 &  x320 &  x323 &  x329 &  x332 &  x338 &  x365 &  x371 &  x377 &  x380 &  x395 &  x404 &  x410 &  x425 &  x428 &  x434 &  x440 &  x461 &  x467 &  x482 &  x497 &  x506 &  x512 &  x514 &  x515 &  x527 &  x536 &  x545 &  x551 &  x553 &  x554 &  x556 &  x557 &  x566 &  x569 &  x571 &  x584 &  x587 &  x590 &  x592 &  x593 &  x595 &  x596 &  x602 &  x610 &  x611 &  x614 &  x620 &  x622 &  x623 &  x626 &  x631 &  x635 &  x638 &  x650 &  x656 &  x662 &  x670 &  x686 &  x698 &  x701 &  x704 &  x710 &  x719 &  x725 &  x728 &  x734 &  x743 &  x746 &  x754 &  x764 &  x767 &  x776 &  x782 &  x791 &  x793 &  x800 &  x803 &  x806 &  x809 &  x818 &  x821 &  x827 &  x829 &  x833 &  x842 &  x857 &  x860 &  x866 &  x868 &  x869 &  x896 &  x905 &  x914 &  x920 &  x926 &  x929 &  x938 &  x953 &  x962 &  x965 &  x974 &  x977 &  x980 &  x998 &  x1010 &  x1028 &  x1037 &  x1055 &  x1064 &  x1079 &  x1082 &  x1094 &  x1100 &  x1112 &  x1118;
assign c386 =  x5 &  x11 &  x14 &  x17 &  x23 &  x26 &  x35 &  x38 &  x44 &  x47 &  x50 &  x56 &  x62 &  x65 &  x68 &  x71 &  x74 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x197 &  x200 &  x205 &  x206 &  x209 &  x215 &  x221 &  x227 &  x230 &  x233 &  x236 &  x238 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x260 &  x263 &  x269 &  x272 &  x274 &  x275 &  x277 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x302 &  x305 &  x308 &  x313 &  x314 &  x316 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x355 &  x356 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x394 &  x395 &  x398 &  x401 &  x407 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x433 &  x434 &  x440 &  x446 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x511 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x548 &  x551 &  x554 &  x557 &  x560 &  x566 &  x569 &  x572 &  x575 &  x581 &  x584 &  x587 &  x590 &  x593 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x623 &  x626 &  x629 &  x632 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x731 &  x734 &  x737 &  x743 &  x749 &  x752 &  x755 &  x758 &  x764 &  x767 &  x770 &  x773 &  x776 &  x785 &  x787 &  x788 &  x791 &  x794 &  x797 &  x803 &  x806 &  x809 &  x815 &  x818 &  x821 &  x824 &  x826 &  x827 &  x830 &  x833 &  x836 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x893 &  x896 &  x899 &  x902 &  x908 &  x911 &  x914 &  x920 &  x923 &  x926 &  x929 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x962 &  x965 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130 & ~x522 & ~x585 & ~x600 & ~x624 & ~x663 & ~x702 & ~x741 & ~x780 & ~x819 & ~x966;
assign c388 =  x2 &  x8 &  x17 &  x20 &  x32 &  x56 &  x74 &  x86 &  x92 &  x95 &  x104 &  x113 &  x122 &  x134 &  x155 &  x161 &  x164 &  x170 &  x173 &  x176 &  x182 &  x209 &  x221 &  x233 &  x244 &  x254 &  x260 &  x277 &  x287 &  x302 &  x305 &  x308 &  x323 &  x326 &  x353 &  x355 &  x359 &  x368 &  x380 &  x386 &  x389 &  x394 &  x395 &  x407 &  x434 &  x437 &  x446 &  x452 &  x458 &  x464 &  x470 &  x472 &  x503 &  x506 &  x515 &  x524 &  x530 &  x536 &  x545 &  x548 &  x550 &  x557 &  x578 &  x587 &  x589 &  x605 &  x620 &  x626 &  x628 &  x629 &  x632 &  x641 &  x644 &  x650 &  x674 &  x692 &  x695 &  x704 &  x722 &  x725 &  x731 &  x740 &  x749 &  x770 &  x815 &  x839 &  x869 &  x872 &  x878 &  x896 &  x911 &  x917 &  x920 &  x926 &  x932 &  x941 &  x953 &  x968 &  x989 &  x995 &  x1004 &  x1007 &  x1010 &  x1016 &  x1025 &  x1067 &  x1082 &  x1085 &  x1127 &  x1130 & ~x339 & ~x340 & ~x561 & ~x678 & ~x780 & ~x858;
assign c390 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x101 &  x104 &  x107 &  x119 &  x122 &  x125 &  x128 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x244 &  x245 &  x248 &  x251 &  x254 &  x257 &  x263 &  x266 &  x269 &  x272 &  x274 &  x275 &  x278 &  x281 &  x283 &  x284 &  x287 &  x290 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x314 &  x317 &  x320 &  x322 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x360 &  x361 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x400 &  x404 &  x407 &  x410 &  x413 &  x419 &  x425 &  x431 &  x433 &  x434 &  x437 &  x439 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x472 &  x473 &  x476 &  x478 &  x479 &  x482 &  x485 &  x488 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x668 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x727 &  x728 &  x731 &  x734 &  x740 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x787 &  x788 &  x791 &  x794 &  x800 &  x803 &  x806 &  x809 &  x818 &  x821 &  x824 &  x826 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x844 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x865 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x900 & ~x939 & ~x1095;
assign c392 =  x2 &  x14 &  x26 &  x29 &  x35 &  x52 &  x68 &  x71 &  x80 &  x89 &  x91 &  x110 &  x113 &  x152 &  x173 &  x194 &  x224 &  x230 &  x233 &  x248 &  x251 &  x257 &  x260 &  x287 &  x296 &  x313 &  x326 &  x329 &  x338 &  x347 &  x374 &  x394 &  x404 &  x410 &  x416 &  x433 &  x452 &  x455 &  x470 &  x473 &  x475 &  x476 &  x479 &  x500 &  x503 &  x515 &  x518 &  x524 &  x530 &  x542 &  x548 &  x551 &  x553 &  x563 &  x581 &  x584 &  x587 &  x593 &  x611 &  x617 &  x626 &  x631 &  x647 &  x674 &  x686 &  x689 &  x704 &  x709 &  x716 &  x737 &  x749 &  x752 &  x766 &  x767 &  x770 &  x782 &  x785 &  x787 &  x797 &  x803 &  x805 &  x827 &  x836 &  x844 &  x848 &  x850 &  x857 &  x869 &  x878 &  x883 &  x890 &  x899 &  x917 &  x941 &  x962 &  x965 &  x968 &  x982 &  x1007 &  x1013 &  x1016 &  x1058 &  x1067 &  x1076 &  x1088 &  x1099 &  x1103 &  x1109 &  x1115 &  x1124 & ~x444 & ~x546 & ~x663 & ~x702 & ~x780 & ~x819 & ~x1014 & ~x1053;
assign c394 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x89 &  x92 &  x98 &  x101 &  x110 &  x113 &  x116 &  x119 &  x125 &  x128 &  x131 &  x140 &  x143 &  x149 &  x152 &  x155 &  x158 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x191 &  x197 &  x200 &  x203 &  x206 &  x218 &  x221 &  x227 &  x233 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x290 &  x293 &  x296 &  x302 &  x305 &  x308 &  x317 &  x323 &  x326 &  x335 &  x338 &  x341 &  x344 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x380 &  x392 &  x395 &  x398 &  x401 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x437 &  x443 &  x446 &  x449 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x497 &  x503 &  x509 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x548 &  x551 &  x554 &  x560 &  x563 &  x566 &  x572 &  x575 &  x578 &  x581 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x626 &  x629 &  x632 &  x635 &  x641 &  x647 &  x650 &  x653 &  x656 &  x659 &  x665 &  x674 &  x677 &  x680 &  x683 &  x689 &  x692 &  x695 &  x698 &  x707 &  x710 &  x713 &  x716 &  x719 &  x725 &  x731 &  x734 &  x740 &  x743 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x773 &  x779 &  x782 &  x788 &  x791 &  x794 &  x797 &  x800 &  x806 &  x812 &  x815 &  x818 &  x821 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x854 &  x857 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x901 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1018 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1118 &  x1130 & ~x30 & ~x69 & ~x108 & ~x843 & ~x882 & ~x909 & ~x912 & ~x951 & ~x990 & ~x991 & ~x993 & ~x1029 & ~x1032 & ~x1068 & ~x1071 & ~x1113;
assign c396 =  x1 &  x2 &  x8 &  x11 &  x14 &  x20 &  x23 &  x50 &  x56 &  x59 &  x65 &  x79 &  x83 &  x101 &  x107 &  x113 &  x119 &  x122 &  x128 &  x134 &  x137 &  x143 &  x155 &  x158 &  x164 &  x167 &  x176 &  x179 &  x182 &  x194 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x236 &  x239 &  x245 &  x248 &  x254 &  x260 &  x263 &  x275 &  x287 &  x290 &  x293 &  x296 &  x302 &  x326 &  x341 &  x344 &  x356 &  x365 &  x383 &  x392 &  x398 &  x401 &  x407 &  x410 &  x413 &  x419 &  x425 &  x431 &  x449 &  x452 &  x455 &  x467 &  x476 &  x479 &  x485 &  x506 &  x521 &  x530 &  x533 &  x542 &  x548 &  x551 &  x554 &  x557 &  x563 &  x566 &  x569 &  x575 &  x599 &  x602 &  x605 &  x608 &  x614 &  x617 &  x626 &  x629 &  x632 &  x635 &  x638 &  x650 &  x653 &  x656 &  x659 &  x662 &  x668 &  x671 &  x683 &  x692 &  x698 &  x710 &  x713 &  x722 &  x728 &  x731 &  x734 &  x749 &  x758 &  x779 &  x782 &  x803 &  x809 &  x812 &  x818 &  x821 &  x833 &  x842 &  x845 &  x848 &  x851 &  x866 &  x869 &  x875 &  x887 &  x899 &  x902 &  x905 &  x911 &  x923 &  x932 &  x938 &  x941 &  x947 &  x950 &  x956 &  x971 &  x980 &  x992 &  x1001 &  x1007 &  x1010 &  x1025 &  x1028 &  x1031 &  x1052 &  x1055 &  x1058 &  x1070 &  x1082 &  x1085 &  x1109 &  x1115 &  x1118 &  x1130 & ~x30 & ~x201 & ~x837 & ~x948 & ~x993 & ~x1008 & ~x1032 & ~x1089 & ~x1098 & ~x1104;
assign c398 =  x13 &  x14 &  x26 &  x35 &  x43 &  x50 &  x53 &  x82 &  x88 &  x89 &  x98 &  x107 &  x113 &  x116 &  x119 &  x140 &  x143 &  x146 &  x152 &  x158 &  x167 &  x179 &  x191 &  x194 &  x209 &  x212 &  x215 &  x218 &  x224 &  x245 &  x254 &  x257 &  x266 &  x274 &  x275 &  x277 &  x278 &  x284 &  x296 &  x308 &  x311 &  x313 &  x314 &  x316 &  x317 &  x320 &  x347 &  x365 &  x368 &  x383 &  x395 &  x401 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x434 &  x446 &  x455 &  x458 &  x473 &  x479 &  x482 &  x485 &  x488 &  x509 &  x518 &  x527 &  x542 &  x557 &  x578 &  x587 &  x599 &  x602 &  x605 &  x608 &  x611 &  x613 &  x617 &  x620 &  x623 &  x626 &  x653 &  x656 &  x662 &  x671 &  x686 &  x689 &  x692 &  x695 &  x704 &  x707 &  x713 &  x746 &  x758 &  x761 &  x764 &  x793 &  x803 &  x821 &  x824 &  x830 &  x839 &  x848 &  x869 &  x875 &  x877 &  x890 &  x899 &  x929 &  x932 &  x935 &  x941 &  x944 &  x953 &  x956 &  x962 &  x977 &  x992 &  x1010 &  x1016 &  x1019 &  x1022 &  x1031 &  x1040 &  x1049 &  x1055 &  x1070 &  x1112 & ~x663 & ~x702 & ~x741 & ~x903 & ~x1098;
assign c3100 =  x2 &  x5 &  x8 &  x14 &  x20 &  x23 &  x29 &  x35 &  x38 &  x41 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x80 &  x83 &  x86 &  x92 &  x95 &  x101 &  x107 &  x110 &  x113 &  x116 &  x125 &  x137 &  x140 &  x143 &  x164 &  x173 &  x176 &  x179 &  x182 &  x188 &  x191 &  x194 &  x197 &  x200 &  x212 &  x215 &  x218 &  x221 &  x224 &  x230 &  x233 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x266 &  x272 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x320 &  x323 &  x326 &  x332 &  x335 &  x338 &  x344 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x403 &  x407 &  x410 &  x416 &  x419 &  x422 &  x428 &  x431 &  x437 &  x440 &  x442 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x470 &  x473 &  x476 &  x482 &  x485 &  x488 &  x500 &  x503 &  x506 &  x512 &  x515 &  x518 &  x519 &  x521 &  x527 &  x533 &  x536 &  x542 &  x545 &  x548 &  x550 &  x551 &  x554 &  x560 &  x563 &  x566 &  x578 &  x581 &  x584 &  x587 &  x589 &  x590 &  x593 &  x598 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x626 &  x628 &  x629 &  x635 &  x641 &  x644 &  x647 &  x653 &  x656 &  x662 &  x665 &  x667 &  x668 &  x671 &  x674 &  x677 &  x689 &  x692 &  x695 &  x701 &  x704 &  x706 &  x707 &  x710 &  x716 &  x719 &  x725 &  x728 &  x734 &  x737 &  x740 &  x743 &  x744 &  x746 &  x752 &  x755 &  x758 &  x764 &  x770 &  x776 &  x782 &  x784 &  x785 &  x788 &  x791 &  x806 &  x812 &  x815 &  x821 &  x823 &  x824 &  x830 &  x836 &  x842 &  x845 &  x851 &  x857 &  x860 &  x866 &  x872 &  x878 &  x881 &  x884 &  x887 &  x890 &  x896 &  x899 &  x901 &  x902 &  x905 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x938 &  x943 &  x947 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1055 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x234 & ~x273 & ~x312 & ~x429;
assign c3102 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x41 &  x44 &  x47 &  x49 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x77 &  x80 &  x86 &  x92 &  x95 &  x98 &  x104 &  x107 &  x110 &  x118 &  x119 &  x125 &  x128 &  x131 &  x134 &  x140 &  x146 &  x152 &  x155 &  x158 &  x167 &  x170 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x260 &  x266 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x296 &  x299 &  x305 &  x308 &  x311 &  x314 &  x317 &  x326 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x436 &  x437 &  x440 &  x443 &  x446 &  x449 &  x455 &  x461 &  x464 &  x470 &  x473 &  x476 &  x478 &  x479 &  x482 &  x485 &  x488 &  x491 &  x500 &  x503 &  x506 &  x509 &  x515 &  x517 &  x518 &  x520 &  x524 &  x527 &  x530 &  x533 &  x539 &  x542 &  x545 &  x551 &  x554 &  x556 &  x557 &  x559 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x593 &  x595 &  x596 &  x598 &  x599 &  x602 &  x611 &  x620 &  x626 &  x632 &  x638 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x682 &  x683 &  x686 &  x689 &  x692 &  x695 &  x704 &  x707 &  x710 &  x713 &  x719 &  x721 &  x725 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x758 &  x761 &  x767 &  x773 &  x776 &  x788 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x860 &  x863 &  x866 &  x872 &  x878 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x908 &  x911 &  x914 &  x920 &  x926 &  x932 &  x935 &  x938 &  x941 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x977 &  x983 &  x986 &  x989 &  x995 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1067 &  x1070 &  x1082 &  x1091 &  x1094 &  x1097 &  x1100 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130 & ~x30 & ~x69 & ~x84;
assign c3104 =  x8 &  x13 &  x20 &  x23 &  x35 &  x44 &  x47 &  x52 &  x62 &  x74 &  x77 &  x80 &  x86 &  x89 &  x95 &  x122 &  x125 &  x128 &  x134 &  x143 &  x146 &  x149 &  x155 &  x164 &  x179 &  x182 &  x191 &  x197 &  x199 &  x200 &  x224 &  x238 &  x245 &  x272 &  x277 &  x278 &  x281 &  x284 &  x302 &  x308 &  x311 &  x316 &  x317 &  x323 &  x329 &  x344 &  x350 &  x374 &  x377 &  x383 &  x398 &  x401 &  x419 &  x422 &  x428 &  x431 &  x437 &  x440 &  x449 &  x455 &  x461 &  x472 &  x476 &  x488 &  x491 &  x497 &  x512 &  x518 &  x524 &  x527 &  x539 &  x548 &  x554 &  x566 &  x575 &  x578 &  x581 &  x584 &  x596 &  x611 &  x617 &  x644 &  x656 &  x668 &  x670 &  x671 &  x674 &  x677 &  x680 &  x686 &  x692 &  x695 &  x709 &  x722 &  x725 &  x727 &  x728 &  x731 &  x740 &  x755 &  x767 &  x772 &  x773 &  x776 &  x782 &  x785 &  x797 &  x800 &  x812 &  x821 &  x833 &  x839 &  x848 &  x851 &  x866 &  x887 &  x893 &  x896 &  x911 &  x920 &  x923 &  x932 &  x935 &  x941 &  x962 &  x971 &  x974 &  x980 &  x989 &  x1001 &  x1007 &  x1019 &  x1022 &  x1034 &  x1037 &  x1043 &  x1046 &  x1052 &  x1055 &  x1064 &  x1067 &  x1085 &  x1091 &  x1100 &  x1109 &  x1130 & ~x336 & ~x579 & ~x663 & ~x703 & ~x783 & ~x858 & ~x1053;
assign c3106 =  x5 &  x8 &  x11 &  x17 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x47 &  x59 &  x65 &  x71 &  x77 &  x80 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x113 &  x116 &  x119 &  x122 &  x131 &  x134 &  x137 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x176 &  x179 &  x185 &  x191 &  x194 &  x197 &  x200 &  x203 &  x209 &  x215 &  x218 &  x224 &  x230 &  x239 &  x242 &  x248 &  x251 &  x257 &  x260 &  x263 &  x266 &  x275 &  x278 &  x281 &  x284 &  x287 &  x304 &  x308 &  x314 &  x323 &  x326 &  x329 &  x332 &  x335 &  x343 &  x347 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x380 &  x383 &  x386 &  x389 &  x395 &  x401 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x443 &  x446 &  x448 &  x449 &  x455 &  x458 &  x467 &  x470 &  x479 &  x485 &  x488 &  x491 &  x494 &  x500 &  x503 &  x509 &  x512 &  x515 &  x521 &  x527 &  x536 &  x542 &  x545 &  x548 &  x554 &  x575 &  x578 &  x581 &  x584 &  x590 &  x596 &  x605 &  x608 &  x611 &  x617 &  x623 &  x629 &  x635 &  x638 &  x641 &  x644 &  x650 &  x656 &  x662 &  x665 &  x674 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x703 &  x704 &  x707 &  x710 &  x719 &  x722 &  x725 &  x731 &  x737 &  x740 &  x743 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x781 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x806 &  x809 &  x812 &  x818 &  x820 &  x827 &  x830 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x859 &  x860 &  x862 &  x863 &  x869 &  x878 &  x881 &  x884 &  x890 &  x893 &  x896 &  x899 &  x901 &  x902 &  x907 &  x908 &  x911 &  x914 &  x920 &  x923 &  x926 &  x929 &  x932 &  x940 &  x941 &  x944 &  x946 &  x947 &  x959 &  x962 &  x965 &  x971 &  x979 &  x980 &  x983 &  x985 &  x986 &  x989 &  x992 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1018 &  x1019 &  x1034 &  x1040 &  x1049 &  x1052 &  x1055 &  x1057 &  x1058 &  x1064 &  x1076 &  x1082 &  x1085 &  x1088 &  x1094 &  x1097 &  x1106 &  x1109 &  x1118 &  x1121 &  x1130 & ~x669 & ~x687 & ~x726 & ~x792 & ~x795 & ~x831 & ~x834;
assign c3108 =  x2 &  x5 &  x8 &  x11 &  x17 &  x20 &  x23 &  x29 &  x32 &  x35 &  x44 &  x50 &  x56 &  x59 &  x71 &  x74 &  x77 &  x86 &  x107 &  x113 &  x116 &  x119 &  x122 &  x125 &  x131 &  x134 &  x137 &  x140 &  x143 &  x149 &  x155 &  x161 &  x167 &  x170 &  x173 &  x182 &  x185 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x239 &  x245 &  x248 &  x251 &  x254 &  x263 &  x266 &  x272 &  x275 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x319 &  x326 &  x329 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x365 &  x368 &  x374 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x401 &  x403 &  x406 &  x407 &  x409 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x445 &  x446 &  x449 &  x452 &  x458 &  x464 &  x467 &  x470 &  x476 &  x479 &  x482 &  x485 &  x488 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x511 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x584 &  x587 &  x589 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x623 &  x626 &  x628 &  x629 &  x632 &  x641 &  x644 &  x653 &  x659 &  x662 &  x664 &  x665 &  x667 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x701 &  x703 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x725 &  x731 &  x737 &  x740 &  x742 &  x743 &  x745 &  x746 &  x749 &  x755 &  x758 &  x761 &  x767 &  x770 &  x773 &  x776 &  x784 &  x785 &  x788 &  x794 &  x797 &  x800 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x827 &  x830 &  x836 &  x839 &  x845 &  x848 &  x854 &  x857 &  x860 &  x862 &  x866 &  x869 &  x872 &  x878 &  x881 &  x887 &  x890 &  x893 &  x899 &  x901 &  x905 &  x911 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x977 &  x983 &  x989 &  x992 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1043 &  x1049 &  x1058 &  x1061 &  x1064 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x12 & ~x1065 & ~x1104;
assign c3110 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x397 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x436 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x475 &  x476 &  x479 &  x482 &  x485 &  x488 &  x490 &  x491 &  x493 &  x494 &  x497 &  x499 &  x500 &  x503 &  x506 &  x509 &  x512 &  x514 &  x515 &  x518 &  x520 &  x521 &  x524 &  x526 &  x527 &  x529 &  x530 &  x532 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x553 &  x554 &  x556 &  x557 &  x559 &  x563 &  x565 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x595 &  x596 &  x598 &  x599 &  x602 &  x604 &  x605 &  x607 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x637 &  x638 &  x641 &  x644 &  x646 &  x647 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x676 &  x677 &  x680 &  x683 &  x685 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x715 &  x716 &  x719 &  x722 &  x724 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x754 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x985 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x390 & ~x429 & ~x468 & ~x507 & ~x546;
assign c3112 =  x41 &  x44 &  x47 &  x50 &  x56 &  x121 &  x140 &  x143 &  x155 &  x158 &  x161 &  x196 &  x200 &  x224 &  x230 &  x233 &  x235 &  x239 &  x245 &  x248 &  x251 &  x253 &  x266 &  x269 &  x272 &  x277 &  x281 &  x284 &  x287 &  x293 &  x311 &  x313 &  x316 &  x317 &  x326 &  x350 &  x355 &  x362 &  x386 &  x389 &  x392 &  x394 &  x398 &  x410 &  x413 &  x419 &  x434 &  x452 &  x464 &  x491 &  x497 &  x509 &  x512 &  x515 &  x524 &  x545 &  x551 &  x578 &  x584 &  x592 &  x605 &  x608 &  x626 &  x631 &  x632 &  x635 &  x641 &  x650 &  x653 &  x659 &  x665 &  x668 &  x670 &  x671 &  x695 &  x698 &  x704 &  x725 &  x727 &  x739 &  x740 &  x764 &  x778 &  x779 &  x785 &  x787 &  x791 &  x817 &  x818 &  x821 &  x826 &  x827 &  x832 &  x839 &  x845 &  x851 &  x856 &  x860 &  x872 &  x877 &  x887 &  x902 &  x905 &  x908 &  x923 &  x938 &  x944 &  x950 &  x956 &  x968 &  x980 &  x983 &  x1000 &  x1037 &  x1055 &  x1073 &  x1085 &  x1091 &  x1112;
assign c3114 =  x5 &  x8 &  x11 &  x17 &  x23 &  x26 &  x32 &  x35 &  x38 &  x47 &  x56 &  x68 &  x71 &  x80 &  x86 &  x92 &  x95 &  x101 &  x113 &  x119 &  x122 &  x125 &  x131 &  x137 &  x143 &  x167 &  x185 &  x188 &  x191 &  x197 &  x209 &  x212 &  x215 &  x242 &  x245 &  x263 &  x269 &  x272 &  x281 &  x296 &  x302 &  x308 &  x317 &  x320 &  x329 &  x341 &  x350 &  x368 &  x371 &  x374 &  x377 &  x386 &  x389 &  x398 &  x404 &  x407 &  x422 &  x437 &  x440 &  x443 &  x452 &  x473 &  x476 &  x482 &  x485 &  x494 &  x497 &  x506 &  x518 &  x520 &  x527 &  x545 &  x554 &  x559 &  x563 &  x572 &  x575 &  x581 &  x587 &  x589 &  x590 &  x593 &  x596 &  x608 &  x614 &  x617 &  x626 &  x635 &  x641 &  x647 &  x656 &  x659 &  x664 &  x665 &  x668 &  x677 &  x680 &  x686 &  x689 &  x692 &  x698 &  x702 &  x706 &  x707 &  x710 &  x713 &  x716 &  x722 &  x731 &  x734 &  x737 &  x740 &  x758 &  x764 &  x770 &  x781 &  x782 &  x788 &  x791 &  x794 &  x800 &  x803 &  x809 &  x833 &  x836 &  x839 &  x851 &  x857 &  x860 &  x862 &  x875 &  x881 &  x887 &  x890 &  x893 &  x898 &  x908 &  x911 &  x917 &  x923 &  x932 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x974 &  x977 &  x983 &  x995 &  x1016 &  x1018 &  x1034 &  x1043 &  x1046 &  x1067 &  x1073 &  x1082 &  x1088 &  x1100 &  x1106 &  x1118 & ~x351 & ~x429;
assign c3116 =  x2 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x64 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x89 &  x92 &  x95 &  x98 &  x104 &  x107 &  x110 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x230 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x292 &  x293 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x317 &  x323 &  x326 &  x329 &  x331 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x365 &  x370 &  x371 &  x374 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x413 &  x416 &  x419 &  x422 &  x425 &  x434 &  x440 &  x443 &  x449 &  x452 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x542 &  x548 &  x551 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x584 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x647 &  x650 &  x653 &  x656 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x712 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x740 &  x743 &  x745 &  x746 &  x750 &  x751 &  x752 &  x755 &  x758 &  x761 &  x767 &  x770 &  x776 &  x779 &  x782 &  x785 &  x788 &  x790 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x827 &  x829 &  x830 &  x833 &  x836 &  x842 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x868 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x45 & ~x84 & ~x195 & ~x234 & ~x273 & ~x312;
assign c3118 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x71 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x107 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x143 &  x146 &  x152 &  x155 &  x158 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x269 &  x272 &  x275 &  x287 &  x290 &  x296 &  x299 &  x305 &  x311 &  x314 &  x323 &  x326 &  x329 &  x331 &  x332 &  x335 &  x338 &  x341 &  x347 &  x353 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x434 &  x436 &  x437 &  x440 &  x442 &  x443 &  x446 &  x455 &  x458 &  x461 &  x467 &  x470 &  x473 &  x476 &  x479 &  x481 &  x482 &  x491 &  x494 &  x497 &  x500 &  x506 &  x509 &  x512 &  x515 &  x518 &  x519 &  x520 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x548 &  x550 &  x551 &  x554 &  x557 &  x559 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x589 &  x590 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x623 &  x628 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x703 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x731 &  x734 &  x737 &  x740 &  x742 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x764 &  x767 &  x770 &  x773 &  x776 &  x781 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x866 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x901 &  x902 &  x905 &  x908 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x943 &  x944 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1097 &  x1106 &  x1112 &  x1115 &  x1127 &  x1130 & ~x429;
assign c3120 =  x2 &  x5 &  x8 &  x13 &  x20 &  x23 &  x26 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x52 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x146 &  x152 &  x155 &  x158 &  x161 &  x164 &  x170 &  x173 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x236 &  x242 &  x245 &  x251 &  x254 &  x257 &  x266 &  x269 &  x272 &  x275 &  x277 &  x278 &  x281 &  x290 &  x293 &  x296 &  x299 &  x308 &  x311 &  x314 &  x316 &  x317 &  x320 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x355 &  x356 &  x365 &  x368 &  x371 &  x374 &  x377 &  x383 &  x392 &  x394 &  x395 &  x398 &  x407 &  x410 &  x416 &  x419 &  x425 &  x428 &  x433 &  x437 &  x440 &  x449 &  x452 &  x458 &  x461 &  x470 &  x472 &  x473 &  x476 &  x479 &  x482 &  x491 &  x503 &  x506 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x590 &  x593 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x662 &  x670 &  x671 &  x674 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x707 &  x709 &  x710 &  x713 &  x715 &  x716 &  x722 &  x725 &  x734 &  x737 &  x740 &  x743 &  x746 &  x752 &  x754 &  x755 &  x761 &  x764 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x793 &  x794 &  x797 &  x800 &  x803 &  x805 &  x806 &  x812 &  x818 &  x821 &  x827 &  x830 &  x832 &  x833 &  x836 &  x842 &  x845 &  x848 &  x854 &  x860 &  x866 &  x871 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x896 &  x905 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x986 &  x988 &  x989 &  x995 &  x998 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1034 &  x1040 &  x1043 &  x1046 &  x1055 &  x1058 &  x1061 &  x1064 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1127 &  x1130 & ~x600 & ~x663 & ~x702 & ~x741 & ~x819 & ~x840 & ~x897 & ~x898 & ~x900 & ~x937 & ~x939 & ~x976 & ~x1014 & ~x1092;
assign c3122 =  x2 &  x11 &  x14 &  x20 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x68 &  x74 &  x80 &  x83 &  x89 &  x101 &  x113 &  x116 &  x119 &  x122 &  x134 &  x140 &  x143 &  x146 &  x152 &  x155 &  x158 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x191 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x238 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x260 &  x263 &  x266 &  x272 &  x275 &  x277 &  x281 &  x287 &  x296 &  x299 &  x302 &  x308 &  x311 &  x314 &  x316 &  x317 &  x320 &  x323 &  x329 &  x338 &  x347 &  x355 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x392 &  x398 &  x401 &  x404 &  x410 &  x413 &  x422 &  x425 &  x428 &  x433 &  x434 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x527 &  x533 &  x536 &  x539 &  x548 &  x554 &  x557 &  x560 &  x566 &  x572 &  x575 &  x584 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x629 &  x632 &  x635 &  x638 &  x641 &  x647 &  x656 &  x662 &  x665 &  x668 &  x670 &  x671 &  x674 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x698 &  x704 &  x707 &  x709 &  x710 &  x719 &  x725 &  x728 &  x737 &  x743 &  x748 &  x749 &  x758 &  x761 &  x764 &  x770 &  x773 &  x776 &  x779 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x821 &  x827 &  x830 &  x833 &  x836 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x896 &  x899 &  x902 &  x905 &  x908 &  x920 &  x926 &  x929 &  x932 &  x938 &  x944 &  x947 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x977 &  x980 &  x986 &  x992 &  x995 &  x998 &  x1004 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x0 & ~x261 & ~x375 & ~x561 & ~x600 & ~x639 & ~x678 & ~x717 & ~x756 & ~x780 & ~x819 & ~x858 & ~x879 & ~x891 & ~x897 & ~x975 & ~x1014;
assign c3124 =  x38 &  x71 &  x74 &  x107 &  x113 &  x125 &  x170 &  x206 &  x227 &  x248 &  x261 &  x278 &  x434 &  x488 &  x491 &  x497 &  x542 &  x557 &  x578 &  x584 &  x668 &  x710 &  x743 &  x746 &  x782 &  x791 &  x830 &  x851 &  x857 &  x859 &  x866 &  x875 &  x881 &  x887 &  x896 &  x901 &  x905 &  x911 &  x941 &  x962 &  x983 &  x995 &  x1004 &  x1013 &  x1016 &  x1064 &  x1115 &  x1118 &  x1124 & ~x198 & ~x510 & ~x588;
assign c3126 =  x5 &  x11 &  x14 &  x17 &  x23 &  x26 &  x29 &  x35 &  x38 &  x41 &  x44 &  x53 &  x56 &  x62 &  x68 &  x74 &  x80 &  x83 &  x89 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x152 &  x155 &  x158 &  x164 &  x167 &  x170 &  x173 &  x182 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x242 &  x245 &  x248 &  x251 &  x253 &  x254 &  x257 &  x260 &  x263 &  x278 &  x281 &  x287 &  x290 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x323 &  x326 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x356 &  x359 &  x362 &  x365 &  x368 &  x370 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x395 &  x409 &  x410 &  x416 &  x419 &  x425 &  x428 &  x434 &  x440 &  x443 &  x452 &  x455 &  x461 &  x470 &  x473 &  x479 &  x481 &  x485 &  x491 &  x497 &  x500 &  x503 &  x506 &  x511 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x545 &  x548 &  x550 &  x551 &  x554 &  x557 &  x566 &  x572 &  x581 &  x584 &  x589 &  x590 &  x596 &  x599 &  x602 &  x605 &  x611 &  x614 &  x623 &  x628 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x656 &  x665 &  x668 &  x671 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x698 &  x704 &  x706 &  x707 &  x713 &  x719 &  x722 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x752 &  x755 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x869 &  x872 &  x878 &  x890 &  x893 &  x896 &  x899 &  x901 &  x908 &  x911 &  x914 &  x917 &  x920 &  x932 &  x935 &  x938 &  x941 &  x944 &  x953 &  x962 &  x974 &  x977 &  x983 &  x989 &  x992 &  x998 &  x1001 &  x1004 &  x1010 &  x1019 &  x1022 &  x1025 &  x1034 &  x1040 &  x1046 &  x1049 &  x1052 &  x1061 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x39 & ~x78 & ~x273 & ~x312 & ~x351 & ~x429 & ~x462 & ~x507 & ~x891;
assign c3128 =  x2 &  x5 &  x8 &  x14 &  x20 &  x23 &  x35 &  x38 &  x41 &  x50 &  x56 &  x59 &  x62 &  x68 &  x83 &  x95 &  x104 &  x107 &  x110 &  x113 &  x119 &  x122 &  x125 &  x128 &  x137 &  x140 &  x143 &  x146 &  x149 &  x164 &  x173 &  x176 &  x182 &  x185 &  x194 &  x203 &  x212 &  x221 &  x230 &  x233 &  x236 &  x251 &  x254 &  x257 &  x266 &  x269 &  x281 &  x287 &  x296 &  x305 &  x314 &  x317 &  x332 &  x335 &  x341 &  x347 &  x350 &  x353 &  x356 &  x371 &  x377 &  x383 &  x388 &  x389 &  x392 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x422 &  x428 &  x434 &  x437 &  x440 &  x443 &  x446 &  x448 &  x452 &  x467 &  x473 &  x476 &  x484 &  x494 &  x497 &  x500 &  x503 &  x518 &  x520 &  x527 &  x530 &  x533 &  x542 &  x545 &  x548 &  x557 &  x559 &  x560 &  x565 &  x569 &  x572 &  x575 &  x578 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x614 &  x617 &  x623 &  x626 &  x632 &  x635 &  x650 &  x656 &  x668 &  x674 &  x677 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x706 &  x710 &  x713 &  x716 &  x728 &  x740 &  x755 &  x758 &  x767 &  x770 &  x776 &  x779 &  x781 &  x782 &  x784 &  x785 &  x791 &  x803 &  x806 &  x812 &  x818 &  x820 &  x821 &  x827 &  x836 &  x839 &  x842 &  x859 &  x860 &  x866 &  x875 &  x878 &  x887 &  x890 &  x893 &  x896 &  x899 &  x901 &  x908 &  x914 &  x920 &  x929 &  x937 &  x938 &  x939 &  x941 &  x944 &  x947 &  x950 &  x956 &  x959 &  x962 &  x971 &  x977 &  x978 &  x980 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1010 &  x1016 &  x1017 &  x1022 &  x1025 &  x1031 &  x1040 &  x1055 &  x1056 &  x1058 &  x1064 &  x1076 &  x1088 &  x1091 &  x1094 &  x1095 &  x1096 &  x1103 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x282 & ~x312 & ~x315 & ~x354 & ~x390 & ~x429 & ~x468;
assign c3130 =  x11 &  x17 &  x23 &  x25 &  x26 &  x29 &  x35 &  x41 &  x47 &  x50 &  x53 &  x59 &  x65 &  x68 &  x74 &  x83 &  x95 &  x101 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x137 &  x158 &  x161 &  x167 &  x169 &  x170 &  x173 &  x179 &  x185 &  x188 &  x191 &  x203 &  x206 &  x207 &  x212 &  x215 &  x218 &  x233 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x263 &  x266 &  x269 &  x272 &  x275 &  x287 &  x293 &  x302 &  x323 &  x326 &  x329 &  x335 &  x338 &  x347 &  x350 &  x353 &  x356 &  x362 &  x365 &  x368 &  x371 &  x374 &  x380 &  x386 &  x398 &  x413 &  x419 &  x422 &  x431 &  x434 &  x437 &  x440 &  x446 &  x455 &  x461 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x488 &  x491 &  x494 &  x503 &  x506 &  x509 &  x515 &  x530 &  x533 &  x536 &  x542 &  x548 &  x550 &  x554 &  x557 &  x569 &  x572 &  x575 &  x578 &  x584 &  x589 &  x593 &  x596 &  x602 &  x608 &  x614 &  x620 &  x623 &  x626 &  x628 &  x635 &  x638 &  x650 &  x653 &  x656 &  x659 &  x665 &  x671 &  x674 &  x677 &  x686 &  x689 &  x692 &  x701 &  x704 &  x707 &  x710 &  x716 &  x725 &  x728 &  x731 &  x737 &  x740 &  x749 &  x755 &  x758 &  x764 &  x773 &  x779 &  x782 &  x785 &  x791 &  x797 &  x800 &  x818 &  x821 &  x824 &  x827 &  x839 &  x842 &  x850 &  x863 &  x866 &  x869 &  x878 &  x887 &  x890 &  x893 &  x896 &  x902 &  x905 &  x917 &  x920 &  x923 &  x932 &  x941 &  x944 &  x947 &  x953 &  x956 &  x959 &  x971 &  x974 &  x986 &  x992 &  x994 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1031 &  x1037 &  x1043 &  x1052 &  x1058 &  x1064 &  x1073 &  x1076 &  x1079 &  x1088 &  x1100 &  x1106 &  x1109 &  x1115 &  x1121 &  x1127 &  x1130 & ~x309 & ~x348 & ~x897 & ~x1092;
assign c3132 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x89 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x226 &  x227 &  x230 &  x233 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x260 &  x263 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x320 &  x326 &  x329 &  x332 &  x335 &  x341 &  x344 &  x347 &  x350 &  x353 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x431 &  x434 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x479 &  x482 &  x485 &  x488 &  x491 &  x497 &  x500 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x530 &  x533 &  x536 &  x539 &  x542 &  x548 &  x551 &  x554 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x608 &  x611 &  x617 &  x626 &  x628 &  x629 &  x632 &  x635 &  x641 &  x644 &  x650 &  x656 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x803 &  x806 &  x809 &  x812 &  x815 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x941 &  x944 &  x950 &  x953 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 &  x1130 & ~x48 & ~x126 & ~x165 & ~x312 & ~x351 & ~x390 & ~x429 & ~x1029 & ~x1047 & ~x1104 & ~x1107 & ~x1125;
assign c3134 =  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x47 &  x53 &  x56 &  x59 &  x68 &  x71 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x254 &  x257 &  x260 &  x263 &  x269 &  x272 &  x278 &  x281 &  x284 &  x287 &  x293 &  x299 &  x302 &  x305 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x359 &  x362 &  x365 &  x371 &  x374 &  x380 &  x383 &  x386 &  x389 &  x392 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x428 &  x431 &  x434 &  x440 &  x443 &  x446 &  x449 &  x452 &  x458 &  x461 &  x464 &  x470 &  x473 &  x476 &  x479 &  x482 &  x491 &  x494 &  x497 &  x503 &  x506 &  x512 &  x515 &  x518 &  x521 &  x524 &  x530 &  x533 &  x536 &  x542 &  x545 &  x548 &  x551 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x634 &  x635 &  x638 &  x644 &  x647 &  x650 &  x653 &  x659 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x719 &  x722 &  x725 &  x728 &  x734 &  x737 &  x740 &  x749 &  x755 &  x761 &  x764 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x797 &  x800 &  x803 &  x809 &  x812 &  x815 &  x818 &  x824 &  x827 &  x830 &  x842 &  x845 &  x848 &  x851 &  x857 &  x860 &  x863 &  x872 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x935 &  x938 &  x944 &  x947 &  x950 &  x953 &  x956 &  x962 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1091 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x45 & ~x876 & ~x894 & ~x909 & ~x915 & ~x987 & ~x993 & ~x1029 & ~x1035 & ~x1068;
assign c3136 =  x2 &  x5 &  x14 &  x23 &  x26 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x62 &  x77 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x125 &  x143 &  x149 &  x152 &  x158 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x239 &  x242 &  x245 &  x248 &  x251 &  x257 &  x263 &  x269 &  x272 &  x275 &  x281 &  x290 &  x311 &  x320 &  x322 &  x323 &  x329 &  x335 &  x338 &  x341 &  x347 &  x359 &  x362 &  x368 &  x374 &  x380 &  x400 &  x401 &  x407 &  x410 &  x413 &  x419 &  x431 &  x434 &  x439 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x464 &  x470 &  x476 &  x478 &  x479 &  x485 &  x494 &  x497 &  x500 &  x511 &  x521 &  x530 &  x539 &  x542 &  x548 &  x551 &  x554 &  x557 &  x563 &  x578 &  x584 &  x593 &  x596 &  x599 &  x602 &  x608 &  x617 &  x620 &  x626 &  x629 &  x632 &  x641 &  x644 &  x653 &  x656 &  x659 &  x668 &  x671 &  x683 &  x689 &  x692 &  x701 &  x707 &  x710 &  x713 &  x719 &  x722 &  x731 &  x737 &  x749 &  x755 &  x761 &  x764 &  x776 &  x779 &  x785 &  x788 &  x800 &  x809 &  x815 &  x824 &  x830 &  x839 &  x851 &  x854 &  x857 &  x860 &  x872 &  x875 &  x878 &  x884 &  x887 &  x890 &  x896 &  x905 &  x908 &  x911 &  x920 &  x923 &  x932 &  x935 &  x943 &  x947 &  x953 &  x962 &  x965 &  x974 &  x977 &  x986 &  x1001 &  x1004 &  x1010 &  x1016 &  x1025 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1064 &  x1079 &  x1082 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1124 & ~x936 & ~x993 & ~x1014 & ~x1053 & ~x1056 & ~x1092;
assign c3138 =  x5 &  x8 &  x11 &  x17 &  x20 &  x23 &  x26 &  x32 &  x41 &  x50 &  x77 &  x86 &  x98 &  x101 &  x104 &  x107 &  x110 &  x116 &  x128 &  x140 &  x143 &  x146 &  x149 &  x167 &  x170 &  x173 &  x176 &  x185 &  x188 &  x194 &  x203 &  x215 &  x218 &  x227 &  x230 &  x242 &  x245 &  x248 &  x254 &  x263 &  x272 &  x278 &  x281 &  x285 &  x293 &  x299 &  x305 &  x326 &  x332 &  x335 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x368 &  x371 &  x374 &  x377 &  x386 &  x389 &  x394 &  x395 &  x398 &  x401 &  x413 &  x422 &  x425 &  x431 &  x443 &  x446 &  x452 &  x458 &  x467 &  x470 &  x479 &  x494 &  x497 &  x503 &  x512 &  x527 &  x533 &  x539 &  x545 &  x548 &  x551 &  x554 &  x563 &  x575 &  x578 &  x581 &  x584 &  x589 &  x593 &  x608 &  x623 &  x626 &  x628 &  x638 &  x641 &  x647 &  x653 &  x656 &  x665 &  x668 &  x671 &  x677 &  x680 &  x686 &  x698 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x731 &  x752 &  x755 &  x773 &  x776 &  x787 &  x791 &  x803 &  x806 &  x809 &  x821 &  x830 &  x839 &  x842 &  x845 &  x851 &  x857 &  x866 &  x875 &  x878 &  x884 &  x887 &  x890 &  x893 &  x905 &  x920 &  x929 &  x944 &  x959 &  x965 &  x968 &  x974 &  x977 &  x998 &  x1004 &  x1010 &  x1013 &  x1019 &  x1025 &  x1028 &  x1034 &  x1052 &  x1064 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1109 &  x1112 &  x1118 &  x1121 &  x1127 & ~x117 & ~x195 & ~x228 & ~x657 & ~x780 & ~x858 & ~x897 & ~x936 & ~x975 & ~x1014 & ~x1053 & ~x1092;
assign c3140 =  x2 &  x4 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x38 &  x40 &  x41 &  x43 &  x44 &  x47 &  x50 &  x56 &  x59 &  x61 &  x62 &  x65 &  x71 &  x74 &  x77 &  x83 &  x86 &  x89 &  x92 &  x95 &  x101 &  x107 &  x110 &  x113 &  x116 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x235 &  x236 &  x239 &  x245 &  x248 &  x251 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x274 &  x275 &  x277 &  x281 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x314 &  x316 &  x317 &  x320 &  x326 &  x332 &  x335 &  x344 &  x347 &  x350 &  x353 &  x356 &  x362 &  x365 &  x368 &  x371 &  x374 &  x380 &  x383 &  x386 &  x389 &  x392 &  x394 &  x398 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x428 &  x431 &  x433 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x467 &  x470 &  x472 &  x473 &  x476 &  x482 &  x485 &  x488 &  x497 &  x500 &  x506 &  x509 &  x515 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x592 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x613 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x652 &  x656 &  x659 &  x662 &  x665 &  x668 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x709 &  x710 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x746 &  x749 &  x752 &  x755 &  x761 &  x767 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x821 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x866 &  x869 &  x872 &  x875 &  x878 &  x887 &  x890 &  x893 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x947 &  x950 &  x953 &  x956 &  x962 &  x965 &  x968 &  x977 &  x980 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x30 & ~x69 & ~x663 & ~x702 & ~x741 & ~x780;
assign c3142 =  x2 &  x17 &  x20 &  x23 &  x26 &  x29 &  x38 &  x41 &  x46 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x89 &  x92 &  x98 &  x104 &  x110 &  x113 &  x116 &  x119 &  x122 &  x128 &  x134 &  x137 &  x140 &  x143 &  x149 &  x155 &  x161 &  x164 &  x167 &  x170 &  x179 &  x191 &  x194 &  x197 &  x203 &  x209 &  x218 &  x224 &  x233 &  x236 &  x239 &  x245 &  x248 &  x251 &  x257 &  x263 &  x269 &  x272 &  x275 &  x278 &  x284 &  x287 &  x290 &  x299 &  x302 &  x311 &  x314 &  x316 &  x317 &  x323 &  x332 &  x335 &  x338 &  x341 &  x347 &  x355 &  x356 &  x359 &  x362 &  x368 &  x371 &  x377 &  x380 &  x386 &  x389 &  x394 &  x398 &  x401 &  x410 &  x416 &  x422 &  x425 &  x428 &  x433 &  x440 &  x443 &  x449 &  x458 &  x461 &  x464 &  x467 &  x470 &  x472 &  x479 &  x485 &  x491 &  x494 &  x503 &  x506 &  x512 &  x515 &  x518 &  x524 &  x527 &  x530 &  x533 &  x542 &  x545 &  x548 &  x550 &  x551 &  x554 &  x560 &  x563 &  x572 &  x575 &  x581 &  x587 &  x593 &  x599 &  x602 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x641 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x671 &  x683 &  x686 &  x692 &  x698 &  x701 &  x707 &  x713 &  x719 &  x731 &  x746 &  x752 &  x758 &  x761 &  x773 &  x782 &  x785 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x836 &  x851 &  x854 &  x860 &  x866 &  x869 &  x871 &  x872 &  x875 &  x878 &  x881 &  x902 &  x905 &  x911 &  x914 &  x920 &  x926 &  x932 &  x935 &  x944 &  x947 &  x953 &  x956 &  x962 &  x968 &  x971 &  x974 &  x977 &  x983 &  x986 &  x989 &  x992 &  x998 &  x1000 &  x1001 &  x1004 &  x1022 &  x1025 &  x1028 &  x1031 &  x1033 &  x1037 &  x1046 &  x1049 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1094 &  x1097 &  x1100 &  x1106 &  x1115 &  x1118 &  x1124 &  x1130 & ~x600 & ~x639 & ~x663 & ~x678 & ~x702 & ~x717 & ~x756 & ~x780 & ~x781 & ~x819 & ~x820 & ~x858 & ~x859 & ~x897 & ~x898 & ~x1014 & ~x1053 & ~x1092;
assign c3144 =  x8 &  x14 &  x23 &  x26 &  x29 &  x35 &  x38 &  x41 &  x44 &  x50 &  x53 &  x56 &  x62 &  x68 &  x74 &  x77 &  x80 &  x104 &  x107 &  x116 &  x122 &  x131 &  x134 &  x137 &  x143 &  x152 &  x155 &  x158 &  x164 &  x167 &  x170 &  x185 &  x191 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x233 &  x236 &  x242 &  x251 &  x257 &  x263 &  x269 &  x275 &  x284 &  x293 &  x296 &  x299 &  x302 &  x311 &  x320 &  x323 &  x326 &  x332 &  x335 &  x338 &  x344 &  x350 &  x359 &  x362 &  x365 &  x371 &  x383 &  x392 &  x394 &  x395 &  x398 &  x413 &  x428 &  x432 &  x433 &  x434 &  x440 &  x452 &  x471 &  x476 &  x479 &  x482 &  x485 &  x488 &  x494 &  x500 &  x509 &  x511 &  x515 &  x518 &  x521 &  x524 &  x530 &  x536 &  x548 &  x550 &  x557 &  x560 &  x566 &  x575 &  x581 &  x584 &  x593 &  x596 &  x605 &  x608 &  x623 &  x632 &  x641 &  x644 &  x656 &  x665 &  x668 &  x674 &  x680 &  x686 &  x689 &  x692 &  x707 &  x713 &  x716 &  x722 &  x731 &  x734 &  x740 &  x743 &  x748 &  x752 &  x758 &  x764 &  x767 &  x770 &  x773 &  x779 &  x785 &  x794 &  x797 &  x803 &  x815 &  x818 &  x824 &  x827 &  x833 &  x839 &  x845 &  x851 &  x857 &  x866 &  x869 &  x889 &  x905 &  x911 &  x917 &  x920 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x950 &  x968 &  x977 &  x980 &  x983 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1019 &  x1022 &  x1034 &  x1037 &  x1040 &  x1058 &  x1070 &  x1073 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x123 & ~x162 & ~x339 & ~x663 & ~x702 & ~x819 & ~x858;
assign c3146 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x104 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x350 &  x353 &  x359 &  x362 &  x364 &  x365 &  x368 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x403 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x428 &  x431 &  x434 &  x437 &  x442 &  x443 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x470 &  x473 &  x476 &  x479 &  x481 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x518 &  x520 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x559 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x584 &  x587 &  x590 &  x593 &  x596 &  x598 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x626 &  x632 &  x635 &  x637 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x794 &  x800 &  x806 &  x809 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x851 &  x854 &  x857 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x890 &  x893 &  x896 &  x902 &  x905 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x946 &  x947 &  x950 &  x953 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x976 &  x977 &  x980 &  x985 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1024 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x3 & ~x42 & ~x120 & ~x159 & ~x162 & ~x198 & ~x201 & ~x237 & ~x276 & ~x315 & ~x354 & ~x393 & ~x471;
assign c3148 =  x2 &  x5 &  x8 &  x13 &  x20 &  x29 &  x35 &  x41 &  x44 &  x47 &  x50 &  x56 &  x59 &  x65 &  x68 &  x80 &  x86 &  x92 &  x95 &  x101 &  x104 &  x107 &  x113 &  x119 &  x122 &  x125 &  x128 &  x131 &  x140 &  x143 &  x146 &  x149 &  x152 &  x167 &  x170 &  x176 &  x185 &  x188 &  x191 &  x194 &  x197 &  x199 &  x203 &  x209 &  x212 &  x215 &  x218 &  x221 &  x227 &  x233 &  x236 &  x238 &  x239 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x277 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x308 &  x316 &  x317 &  x326 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x355 &  x359 &  x365 &  x368 &  x371 &  x377 &  x380 &  x386 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x428 &  x431 &  x433 &  x440 &  x446 &  x449 &  x452 &  x461 &  x472 &  x479 &  x488 &  x494 &  x497 &  x503 &  x506 &  x509 &  x511 &  x512 &  x515 &  x518 &  x533 &  x536 &  x542 &  x545 &  x550 &  x554 &  x557 &  x560 &  x563 &  x566 &  x572 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x635 &  x638 &  x644 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x671 &  x674 &  x683 &  x686 &  x692 &  x698 &  x701 &  x707 &  x713 &  x716 &  x719 &  x725 &  x728 &  x734 &  x743 &  x749 &  x752 &  x755 &  x761 &  x764 &  x767 &  x770 &  x773 &  x785 &  x788 &  x794 &  x797 &  x800 &  x803 &  x806 &  x812 &  x821 &  x830 &  x833 &  x836 &  x839 &  x845 &  x854 &  x869 &  x875 &  x878 &  x881 &  x883 &  x893 &  x899 &  x902 &  x911 &  x914 &  x920 &  x923 &  x929 &  x932 &  x938 &  x941 &  x944 &  x947 &  x953 &  x956 &  x965 &  x968 &  x971 &  x974 &  x983 &  x992 &  x1025 &  x1027 &  x1028 &  x1031 &  x1034 &  x1043 &  x1055 &  x1061 &  x1064 &  x1070 &  x1082 &  x1085 &  x1091 &  x1100 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130 & ~x639 & ~x717 & ~x741 & ~x819 & ~x820 & ~x858 & ~x859 & ~x898 & ~x900 & ~x936 & ~x975 & ~x1092;
assign c3150 =  x5 &  x11 &  x13 &  x20 &  x29 &  x32 &  x35 &  x38 &  x47 &  x50 &  x56 &  x62 &  x65 &  x68 &  x74 &  x77 &  x83 &  x86 &  x98 &  x101 &  x104 &  x107 &  x113 &  x122 &  x125 &  x128 &  x134 &  x140 &  x149 &  x152 &  x164 &  x167 &  x182 &  x191 &  x199 &  x200 &  x203 &  x218 &  x221 &  x230 &  x238 &  x239 &  x242 &  x251 &  x260 &  x263 &  x266 &  x269 &  x277 &  x278 &  x281 &  x284 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x313 &  x314 &  x320 &  x323 &  x326 &  x332 &  x338 &  x341 &  x344 &  x350 &  x359 &  x362 &  x365 &  x371 &  x374 &  x395 &  x398 &  x401 &  x407 &  x410 &  x416 &  x419 &  x425 &  x428 &  x434 &  x443 &  x449 &  x455 &  x458 &  x467 &  x470 &  x476 &  x479 &  x482 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x527 &  x542 &  x551 &  x557 &  x566 &  x569 &  x572 &  x575 &  x578 &  x584 &  x596 &  x599 &  x605 &  x614 &  x620 &  x632 &  x650 &  x659 &  x674 &  x677 &  x680 &  x683 &  x692 &  x695 &  x698 &  x701 &  x707 &  x713 &  x728 &  x731 &  x737 &  x740 &  x743 &  x749 &  x755 &  x761 &  x770 &  x776 &  x779 &  x782 &  x788 &  x794 &  x800 &  x803 &  x812 &  x818 &  x830 &  x833 &  x836 &  x838 &  x844 &  x845 &  x851 &  x857 &  x866 &  x872 &  x883 &  x884 &  x887 &  x896 &  x905 &  x914 &  x922 &  x923 &  x926 &  x932 &  x938 &  x941 &  x947 &  x953 &  x956 &  x965 &  x980 &  x986 &  x998 &  x1007 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1043 &  x1055 &  x1058 &  x1061 &  x1064 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1127 & ~x105 & ~x144 & ~x300 & ~x339 & ~x444 & ~x624 & ~x780 & ~x819 & ~x858 & ~x897 & ~x906 & ~x975 & ~x984 & ~x1092;
assign c3152 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x35 &  x38 &  x41 &  x47 &  x50 &  x56 &  x59 &  x62 &  x65 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x98 &  x101 &  x116 &  x119 &  x122 &  x125 &  x131 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x161 &  x170 &  x173 &  x185 &  x188 &  x194 &  x200 &  x209 &  x212 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x251 &  x254 &  x257 &  x263 &  x266 &  x269 &  x272 &  x281 &  x284 &  x290 &  x296 &  x299 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x350 &  x353 &  x362 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x415 &  x419 &  x425 &  x428 &  x431 &  x434 &  x440 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x470 &  x473 &  x475 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x509 &  x512 &  x521 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x560 &  x563 &  x566 &  x569 &  x571 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x617 &  x620 &  x626 &  x629 &  x632 &  x635 &  x638 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x689 &  x698 &  x701 &  x710 &  x713 &  x716 &  x728 &  x731 &  x734 &  x737 &  x743 &  x746 &  x749 &  x755 &  x758 &  x764 &  x767 &  x770 &  x776 &  x779 &  x785 &  x788 &  x794 &  x797 &  x800 &  x809 &  x818 &  x821 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x851 &  x860 &  x863 &  x866 &  x875 &  x878 &  x887 &  x890 &  x893 &  x899 &  x905 &  x908 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x938 &  x941 &  x947 &  x950 &  x959 &  x962 &  x965 &  x968 &  x971 &  x977 &  x980 &  x983 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 & ~x201 & ~x390 & ~x429 & ~x468 & ~x507 & ~x846 & ~x891 & ~x912 & ~x933 & ~x1107;
assign c3154 =  x23 &  x26 &  x41 &  x53 &  x56 &  x62 &  x68 &  x71 &  x77 &  x80 &  x86 &  x92 &  x94 &  x110 &  x116 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x143 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x182 &  x188 &  x194 &  x197 &  x218 &  x227 &  x230 &  x242 &  x245 &  x263 &  x266 &  x278 &  x287 &  x290 &  x293 &  x299 &  x302 &  x308 &  x314 &  x323 &  x329 &  x335 &  x338 &  x341 &  x350 &  x356 &  x359 &  x368 &  x377 &  x383 &  x389 &  x398 &  x404 &  x407 &  x410 &  x419 &  x422 &  x431 &  x434 &  x446 &  x449 &  x452 &  x458 &  x461 &  x464 &  x470 &  x476 &  x482 &  x485 &  x488 &  x497 &  x500 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x536 &  x542 &  x545 &  x560 &  x563 &  x572 &  x575 &  x578 &  x581 &  x584 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x641 &  x644 &  x650 &  x653 &  x662 &  x665 &  x668 &  x671 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x713 &  x716 &  x728 &  x734 &  x737 &  x743 &  x752 &  x761 &  x767 &  x770 &  x776 &  x779 &  x785 &  x788 &  x791 &  x803 &  x812 &  x815 &  x827 &  x836 &  x839 &  x857 &  x866 &  x869 &  x872 &  x875 &  x878 &  x890 &  x896 &  x899 &  x902 &  x905 &  x923 &  x935 &  x941 &  x950 &  x959 &  x962 &  x965 &  x968 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1019 &  x1022 &  x1025 &  x1028 &  x1034 &  x1040 &  x1043 &  x1049 &  x1052 &  x1061 &  x1073 &  x1076 &  x1082 &  x1091 &  x1094 &  x1112 &  x1115 &  x1124 & ~x30 & ~x103 & ~x180 & ~x219 & ~x720 & ~x915 & ~x1026;
assign c3156 =  x5 &  x8 &  x11 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x44 &  x47 &  x53 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x121 &  x122 &  x128 &  x134 &  x137 &  x140 &  x143 &  x146 &  x152 &  x155 &  x158 &  x160 &  x161 &  x167 &  x170 &  x173 &  x179 &  x185 &  x194 &  x199 &  x203 &  x206 &  x212 &  x218 &  x227 &  x230 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x260 &  x263 &  x266 &  x269 &  x272 &  x277 &  x281 &  x284 &  x287 &  x293 &  x296 &  x305 &  x308 &  x311 &  x314 &  x316 &  x317 &  x320 &  x326 &  x332 &  x338 &  x341 &  x344 &  x350 &  x353 &  x356 &  x371 &  x380 &  x383 &  x389 &  x392 &  x394 &  x395 &  x404 &  x407 &  x410 &  x413 &  x419 &  x422 &  x428 &  x431 &  x433 &  x434 &  x437 &  x440 &  x443 &  x452 &  x455 &  x461 &  x470 &  x473 &  x476 &  x479 &  x482 &  x488 &  x491 &  x494 &  x497 &  x500 &  x509 &  x512 &  x518 &  x521 &  x524 &  x527 &  x533 &  x536 &  x542 &  x545 &  x548 &  x551 &  x553 &  x554 &  x557 &  x560 &  x566 &  x572 &  x575 &  x581 &  x584 &  x587 &  x590 &  x592 &  x596 &  x599 &  x602 &  x611 &  x617 &  x620 &  x626 &  x631 &  x635 &  x638 &  x641 &  x644 &  x653 &  x659 &  x668 &  x670 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x704 &  x707 &  x709 &  x710 &  x713 &  x716 &  x725 &  x728 &  x734 &  x737 &  x739 &  x740 &  x743 &  x746 &  x752 &  x755 &  x758 &  x761 &  x766 &  x767 &  x770 &  x778 &  x779 &  x785 &  x788 &  x791 &  x800 &  x805 &  x809 &  x812 &  x815 &  x817 &  x818 &  x824 &  x830 &  x836 &  x839 &  x845 &  x848 &  x854 &  x856 &  x857 &  x860 &  x863 &  x866 &  x875 &  x878 &  x881 &  x887 &  x890 &  x893 &  x896 &  x899 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x941 &  x944 &  x950 &  x953 &  x959 &  x965 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1052 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1088 &  x1094 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x105 & ~x144 & ~x366 & ~x405 & ~x444 & ~x546 & ~x585 & ~x624 & ~x702 & ~x741 & ~x742 & ~x780 & ~x781 & ~x819 & ~x822 & ~x858 & ~x861 & ~x897 & ~x900 & ~x936 & ~x1053;
assign c3158 =  x2 &  x5 &  x8 &  x11 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x265 &  x269 &  x272 &  x275 &  x278 &  x284 &  x287 &  x289 &  x290 &  x293 &  x296 &  x299 &  x302 &  x304 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x367 &  x368 &  x371 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x400 &  x401 &  x404 &  x406 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x439 &  x440 &  x443 &  x445 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x625 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x703 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x742 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x773 &  x776 &  x779 &  x781 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x893 &  x896 &  x899 &  x901 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x940 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x979 &  x980 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x570 & ~x1065 & ~x1104;
assign c3160 =  x1 &  x10 &  x11 &  x14 &  x17 &  x23 &  x32 &  x35 &  x38 &  x40 &  x41 &  x44 &  x49 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x71 &  x74 &  x79 &  x80 &  x83 &  x86 &  x89 &  x95 &  x98 &  x101 &  x104 &  x107 &  x113 &  x116 &  x119 &  x125 &  x128 &  x134 &  x137 &  x140 &  x146 &  x149 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x188 &  x194 &  x197 &  x200 &  x203 &  x209 &  x215 &  x224 &  x227 &  x230 &  x233 &  x236 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x346 &  x347 &  x350 &  x359 &  x362 &  x365 &  x368 &  x371 &  x377 &  x380 &  x382 &  x383 &  x386 &  x389 &  x395 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x425 &  x431 &  x434 &  x437 &  x440 &  x443 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x478 &  x479 &  x482 &  x485 &  x488 &  x494 &  x497 &  x500 &  x503 &  x506 &  x515 &  x517 &  x521 &  x524 &  x527 &  x530 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x559 &  x560 &  x563 &  x569 &  x572 &  x578 &  x584 &  x593 &  x596 &  x599 &  x605 &  x608 &  x614 &  x620 &  x623 &  x626 &  x632 &  x635 &  x641 &  x643 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x785 &  x788 &  x800 &  x806 &  x812 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x968 &  x971 &  x974 &  x977 &  x983 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1052 &  x1058 &  x1061 &  x1067 &  x1073 &  x1079 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x6 & ~x279 & ~x747;
assign c3162 =  x2 &  x11 &  x20 &  x23 &  x29 &  x32 &  x35 &  x41 &  x53 &  x56 &  x62 &  x65 &  x68 &  x71 &  x74 &  x82 &  x83 &  x86 &  x98 &  x101 &  x104 &  x110 &  x113 &  x121 &  x122 &  x125 &  x128 &  x137 &  x140 &  x143 &  x146 &  x158 &  x160 &  x170 &  x173 &  x176 &  x179 &  x182 &  x191 &  x194 &  x198 &  x199 &  x206 &  x212 &  x215 &  x218 &  x227 &  x251 &  x254 &  x257 &  x260 &  x266 &  x269 &  x277 &  x284 &  x287 &  x302 &  x305 &  x314 &  x323 &  x329 &  x332 &  x341 &  x353 &  x356 &  x359 &  x362 &  x368 &  x374 &  x380 &  x383 &  x386 &  x389 &  x394 &  x395 &  x398 &  x401 &  x404 &  x419 &  x422 &  x434 &  x449 &  x467 &  x473 &  x485 &  x491 &  x494 &  x500 &  x503 &  x506 &  x512 &  x530 &  x533 &  x548 &  x551 &  x557 &  x569 &  x575 &  x578 &  x581 &  x584 &  x587 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x631 &  x638 &  x653 &  x656 &  x665 &  x668 &  x670 &  x671 &  x674 &  x680 &  x695 &  x698 &  x704 &  x707 &  x713 &  x722 &  x727 &  x737 &  x740 &  x758 &  x761 &  x767 &  x773 &  x776 &  x782 &  x785 &  x806 &  x809 &  x812 &  x824 &  x827 &  x833 &  x844 &  x845 &  x854 &  x866 &  x875 &  x887 &  x890 &  x905 &  x914 &  x917 &  x929 &  x959 &  x962 &  x965 &  x989 &  x992 &  x995 &  x1001 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1034 &  x1037 &  x1049 &  x1052 &  x1061 &  x1070 &  x1079 &  x1091 &  x1094 &  x1103 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130 & ~x201 & ~x240 & ~x288 & ~x366 & ~x444 & ~x507 & ~x624 & ~x625 & ~x663 & ~x702 & ~x780 & ~x936 & ~x939 & ~x978 & ~x1014 & ~x1056;
assign c3164 =  x2 &  x8 &  x11 &  x14 &  x17 &  x23 &  x29 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x74 &  x77 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x110 &  x113 &  x116 &  x119 &  x125 &  x128 &  x131 &  x134 &  x143 &  x145 &  x149 &  x152 &  x155 &  x158 &  x161 &  x176 &  x179 &  x182 &  x188 &  x191 &  x194 &  x200 &  x203 &  x206 &  x209 &  x212 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x245 &  x248 &  x251 &  x254 &  x257 &  x266 &  x269 &  x272 &  x275 &  x281 &  x287 &  x290 &  x293 &  x296 &  x302 &  x308 &  x323 &  x326 &  x329 &  x335 &  x338 &  x343 &  x344 &  x347 &  x350 &  x353 &  x359 &  x362 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x389 &  x398 &  x400 &  x401 &  x404 &  x407 &  x413 &  x422 &  x425 &  x428 &  x431 &  x434 &  x439 &  x440 &  x443 &  x449 &  x452 &  x458 &  x461 &  x464 &  x467 &  x473 &  x479 &  x485 &  x488 &  x494 &  x497 &  x500 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x584 &  x586 &  x587 &  x590 &  x593 &  x596 &  x602 &  x608 &  x611 &  x625 &  x626 &  x629 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x659 &  x662 &  x664 &  x665 &  x668 &  x674 &  x677 &  x680 &  x683 &  x686 &  x695 &  x698 &  x701 &  x704 &  x716 &  x722 &  x731 &  x734 &  x737 &  x740 &  x742 &  x743 &  x746 &  x749 &  x752 &  x758 &  x761 &  x767 &  x773 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x815 &  x818 &  x821 &  x833 &  x836 &  x848 &  x851 &  x860 &  x862 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x901 &  x902 &  x905 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x943 &  x944 &  x947 &  x950 &  x953 &  x959 &  x962 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1046 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1085 &  x1088 &  x1091 &  x1094 &  x1100 &  x1106 &  x1109 &  x1111 &  x1112 &  x1115 &  x1118 &  x1124 &  x1130;
assign c3166 =  x2 &  x5 &  x8 &  x11 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x50 &  x52 &  x53 &  x56 &  x59 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x164 &  x167 &  x173 &  x176 &  x179 &  x185 &  x188 &  x194 &  x197 &  x200 &  x206 &  x212 &  x218 &  x221 &  x224 &  x227 &  x230 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x269 &  x272 &  x275 &  x277 &  x278 &  x281 &  x284 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x316 &  x317 &  x320 &  x323 &  x326 &  x329 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x355 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x389 &  x392 &  x394 &  x395 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x433 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x458 &  x464 &  x467 &  x470 &  x472 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x503 &  x506 &  x509 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x542 &  x545 &  x551 &  x554 &  x557 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x599 &  x602 &  x605 &  x608 &  x611 &  x620 &  x623 &  x626 &  x629 &  x632 &  x641 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x743 &  x746 &  x748 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x782 &  x785 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x875 &  x878 &  x881 &  x884 &  x887 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x944 &  x947 &  x950 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 & ~x300 & ~x339 & ~x378 & ~x379 & ~x417 & ~x423 & ~x858 & ~x897 & ~x936;
assign c3168 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x35 &  x38 &  x44 &  x50 &  x53 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x89 &  x92 &  x95 &  x98 &  x101 &  x103 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x125 &  x128 &  x131 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x181 &  x185 &  x188 &  x191 &  x193 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x242 &  x245 &  x248 &  x254 &  x257 &  x260 &  x263 &  x269 &  x272 &  x275 &  x278 &  x284 &  x287 &  x290 &  x292 &  x293 &  x296 &  x299 &  x301 &  x305 &  x308 &  x311 &  x317 &  x320 &  x323 &  x326 &  x329 &  x331 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x370 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x403 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x441 &  x442 &  x443 &  x446 &  x449 &  x452 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x478 &  x479 &  x481 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x554 &  x557 &  x569 &  x572 &  x575 &  x578 &  x581 &  x593 &  x596 &  x599 &  x602 &  x608 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x667 &  x668 &  x671 &  x677 &  x680 &  x683 &  x689 &  x692 &  x695 &  x698 &  x701 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x767 &  x770 &  x773 &  x776 &  x782 &  x785 &  x788 &  x791 &  x797 &  x800 &  x809 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x901 &  x902 &  x905 &  x908 &  x911 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x946 &  x947 &  x950 &  x953 &  x959 &  x962 &  x965 &  x968 &  x971 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1019 &  x1022 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1084 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130;
assign c3170 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x116 &  x119 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x322 &  x326 &  x329 &  x335 &  x341 &  x344 &  x347 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x419 &  x422 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x584 &  x587 &  x590 &  x593 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x707 &  x710 &  x712 &  x713 &  x716 &  x719 &  x722 &  x728 &  x731 &  x734 &  x737 &  x743 &  x746 &  x751 &  x752 &  x755 &  x758 &  x761 &  x767 &  x770 &  x773 &  x779 &  x782 &  x785 &  x788 &  x790 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x829 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x868 &  x869 &  x872 &  x875 &  x881 &  x884 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x907 &  x911 &  x914 &  x917 &  x920 &  x923 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x6 & ~x837 & ~x852 & ~x876 & ~x924 & ~x1089;
assign c3172 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x85 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x124 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x277 &  x278 &  x281 &  x284 &  x287 &  x289 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x316 &  x317 &  x320 &  x323 &  x326 &  x328 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x353 &  x355 &  x356 &  x359 &  x362 &  x365 &  x367 &  x368 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x394 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x419 &  x422 &  x425 &  x428 &  x430 &  x431 &  x433 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x508 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x548 &  x550 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x589 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x628 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x667 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x706 &  x707 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x826 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x901 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x940 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x968 &  x971 &  x974 &  x977 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1018 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130;
assign c3174 =  x5 &  x11 &  x14 &  x17 &  x20 &  x26 &  x29 &  x32 &  x38 &  x40 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x65 &  x71 &  x74 &  x77 &  x79 &  x80 &  x89 &  x92 &  x95 &  x98 &  x104 &  x107 &  x110 &  x113 &  x116 &  x118 &  x122 &  x134 &  x140 &  x143 &  x146 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x196 &  x200 &  x206 &  x209 &  x212 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x235 &  x239 &  x245 &  x248 &  x251 &  x257 &  x260 &  x263 &  x272 &  x274 &  x284 &  x287 &  x290 &  x296 &  x299 &  x305 &  x311 &  x313 &  x314 &  x317 &  x320 &  x323 &  x326 &  x332 &  x335 &  x338 &  x341 &  x344 &  x350 &  x353 &  x356 &  x359 &  x362 &  x368 &  x371 &  x374 &  x380 &  x386 &  x395 &  x398 &  x401 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x437 &  x440 &  x443 &  x446 &  x449 &  x455 &  x458 &  x464 &  x467 &  x470 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x509 &  x518 &  x521 &  x524 &  x527 &  x530 &  x539 &  x542 &  x545 &  x551 &  x554 &  x560 &  x566 &  x572 &  x575 &  x578 &  x581 &  x584 &  x596 &  x602 &  x605 &  x608 &  x611 &  x617 &  x623 &  x632 &  x638 &  x641 &  x647 &  x650 &  x656 &  x662 &  x665 &  x674 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x704 &  x710 &  x712 &  x713 &  x719 &  x722 &  x725 &  x728 &  x734 &  x737 &  x740 &  x749 &  x751 &  x752 &  x758 &  x761 &  x773 &  x776 &  x785 &  x788 &  x794 &  x797 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x827 &  x836 &  x839 &  x842 &  x848 &  x851 &  x854 &  x857 &  x866 &  x872 &  x875 &  x890 &  x893 &  x896 &  x902 &  x905 &  x908 &  x914 &  x917 &  x923 &  x929 &  x935 &  x938 &  x941 &  x944 &  x947 &  x953 &  x956 &  x965 &  x968 &  x971 &  x980 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 & ~x57 & ~x96 & ~x123 & ~x162 & ~x192 & ~x231 & ~x330 & ~x369 & ~x408 & ~x447 & ~x816 & ~x942 & ~x1098;
assign c3176 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x280 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x319 &  x320 &  x323 &  x325 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x363 &  x364 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x389 &  x392 &  x395 &  x398 &  x401 &  x403 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x442 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x745 &  x746 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x827 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x901 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x156 & ~x159 & ~x195 & ~x198 & ~x234 & ~x273 & ~x312 & ~x351 & ~x417 & ~x1107;
assign c3178 =  x5 &  x8 &  x11 &  x14 &  x17 &  x26 &  x41 &  x44 &  x47 &  x53 &  x56 &  x62 &  x71 &  x74 &  x83 &  x86 &  x104 &  x110 &  x116 &  x119 &  x134 &  x143 &  x146 &  x152 &  x155 &  x158 &  x167 &  x176 &  x179 &  x182 &  x191 &  x194 &  x206 &  x209 &  x212 &  x227 &  x233 &  x236 &  x239 &  x242 &  x260 &  x275 &  x290 &  x302 &  x314 &  x317 &  x320 &  x332 &  x335 &  x344 &  x347 &  x350 &  x356 &  x371 &  x389 &  x401 &  x410 &  x425 &  x428 &  x449 &  x452 &  x455 &  x458 &  x464 &  x467 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x503 &  x512 &  x521 &  x536 &  x539 &  x542 &  x557 &  x563 &  x566 &  x575 &  x578 &  x581 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x623 &  x629 &  x647 &  x650 &  x653 &  x662 &  x668 &  x674 &  x677 &  x689 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x725 &  x734 &  x745 &  x755 &  x761 &  x764 &  x767 &  x770 &  x784 &  x785 &  x788 &  x794 &  x800 &  x803 &  x809 &  x812 &  x818 &  x823 &  x827 &  x830 &  x833 &  x842 &  x848 &  x851 &  x854 &  x857 &  x860 &  x866 &  x878 &  x896 &  x899 &  x901 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x926 &  x932 &  x935 &  x938 &  x941 &  x943 &  x947 &  x953 &  x962 &  x968 &  x981 &  x982 &  x989 &  x995 &  x1013 &  x1021 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1064 &  x1070 &  x1073 &  x1082 &  x1085 &  x1094 &  x1100 &  x1103 &  x1124 &  x1130 & ~x156 & ~x234 & ~x273 & ~x351 & ~x831 & ~x912 & ~x957 & ~x996 & ~x1002;
assign c3180 =  x2 &  x5 &  x11 &  x14 &  x20 &  x26 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x80 &  x83 &  x89 &  x92 &  x98 &  x101 &  x107 &  x110 &  x116 &  x119 &  x121 &  x122 &  x128 &  x131 &  x134 &  x137 &  x140 &  x149 &  x155 &  x160 &  x161 &  x173 &  x179 &  x182 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x212 &  x221 &  x227 &  x233 &  x236 &  x238 &  x239 &  x245 &  x251 &  x254 &  x263 &  x266 &  x269 &  x272 &  x274 &  x277 &  x278 &  x287 &  x293 &  x296 &  x299 &  x302 &  x311 &  x313 &  x314 &  x316 &  x317 &  x320 &  x332 &  x341 &  x344 &  x347 &  x350 &  x353 &  x355 &  x356 &  x362 &  x365 &  x368 &  x380 &  x383 &  x386 &  x394 &  x395 &  x398 &  x401 &  x407 &  x410 &  x416 &  x419 &  x422 &  x425 &  x433 &  x434 &  x437 &  x440 &  x443 &  x446 &  x452 &  x455 &  x458 &  x461 &  x467 &  x470 &  x472 &  x476 &  x479 &  x482 &  x485 &  x488 &  x497 &  x500 &  x503 &  x509 &  x512 &  x515 &  x518 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x548 &  x553 &  x554 &  x557 &  x563 &  x566 &  x569 &  x572 &  x575 &  x584 &  x587 &  x590 &  x591 &  x592 &  x593 &  x596 &  x599 &  x605 &  x611 &  x617 &  x623 &  x626 &  x629 &  x638 &  x641 &  x650 &  x653 &  x656 &  x662 &  x670 &  x674 &  x677 &  x683 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x713 &  x716 &  x722 &  x725 &  x728 &  x737 &  x743 &  x746 &  x748 &  x755 &  x761 &  x764 &  x776 &  x782 &  x785 &  x788 &  x791 &  x794 &  x800 &  x803 &  x809 &  x811 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x844 &  x845 &  x848 &  x851 &  x854 &  x857 &  x865 &  x869 &  x872 &  x878 &  x881 &  x884 &  x889 &  x890 &  x899 &  x905 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x962 &  x965 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1021 &  x1022 &  x1028 &  x1034 &  x1046 &  x1049 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1106 &  x1112 & ~x327 & ~x483 & ~x663 & ~x702 & ~x703 & ~x741 & ~x742 & ~x781 & ~x819 & ~x822 & ~x858 & ~x900 & ~x936 & ~x975 & ~x978 & ~x1014 & ~x1017 & ~x1053 & ~x1056;
assign c3182 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x31 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x250 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x316 &  x317 &  x320 &  x323 &  x325 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x433 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x508 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x542 &  x545 &  x547 &  x548 &  x550 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x589 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x617 &  x623 &  x626 &  x628 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x667 &  x668 &  x671 &  x674 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x731 &  x734 &  x737 &  x740 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x815 &  x818 &  x821 &  x823 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x234 & ~x474 & ~x492 & ~x513;
assign c3184 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x68 &  x71 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x155 &  x161 &  x164 &  x167 &  x173 &  x179 &  x182 &  x188 &  x191 &  x194 &  x197 &  x203 &  x206 &  x215 &  x218 &  x221 &  x224 &  x226 &  x227 &  x230 &  x236 &  x239 &  x242 &  x245 &  x251 &  x254 &  x257 &  x260 &  x265 &  x266 &  x272 &  x275 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x304 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x332 &  x335 &  x338 &  x341 &  x344 &  x353 &  x356 &  x359 &  x365 &  x371 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x440 &  x443 &  x446 &  x448 &  x449 &  x452 &  x455 &  x458 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x497 &  x500 &  x503 &  x506 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x542 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x647 &  x650 &  x656 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x701 &  x707 &  x710 &  x713 &  x716 &  x719 &  x725 &  x728 &  x731 &  x743 &  x746 &  x749 &  x752 &  x755 &  x761 &  x764 &  x767 &  x770 &  x779 &  x781 &  x782 &  x784 &  x788 &  x791 &  x794 &  x797 &  x800 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x869 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x901 &  x902 &  x905 &  x907 &  x908 &  x914 &  x917 &  x923 &  x929 &  x938 &  x941 &  x944 &  x950 &  x953 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1100 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x951 & ~x990 & ~x993 & ~x1029 & ~x1032 & ~x1071 & ~x1110 & ~x1113;
assign c3186 =  x2 &  x5 &  x8 &  x11 &  x20 &  x23 &  x32 &  x41 &  x50 &  x56 &  x59 &  x62 &  x65 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x128 &  x131 &  x134 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x209 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x254 &  x257 &  x260 &  x266 &  x269 &  x278 &  x281 &  x284 &  x287 &  x290 &  x296 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x323 &  x326 &  x335 &  x338 &  x344 &  x347 &  x350 &  x353 &  x365 &  x371 &  x374 &  x383 &  x389 &  x392 &  x395 &  x401 &  x410 &  x416 &  x419 &  x425 &  x428 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x464 &  x470 &  x473 &  x476 &  x479 &  x482 &  x491 &  x494 &  x497 &  x500 &  x503 &  x515 &  x521 &  x533 &  x539 &  x542 &  x548 &  x551 &  x554 &  x557 &  x560 &  x566 &  x569 &  x572 &  x575 &  x581 &  x587 &  x590 &  x593 &  x596 &  x599 &  x605 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x659 &  x662 &  x665 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x734 &  x737 &  x746 &  x749 &  x764 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x794 &  x797 &  x800 &  x803 &  x806 &  x815 &  x818 &  x821 &  x824 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x857 &  x859 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x890 &  x896 &  x902 &  x911 &  x914 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x937 &  x940 &  x944 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x977 &  x979 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1018 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1052 &  x1054 &  x1055 &  x1058 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1093 &  x1094 &  x1096 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1130 & ~x882 & ~x960 & ~x988 & ~x999 & ~x1026 & ~x1065 & ~x1077 & ~x1078 & ~x1104 & ~x1116;
assign c3188 =  x1 &  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x40 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x65 &  x68 &  x71 &  x74 &  x77 &  x79 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x118 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x157 &  x158 &  x161 &  x164 &  x167 &  x170 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x196 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x449 &  x452 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x740 &  x743 &  x746 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x30 & ~x69 & ~x141 & ~x252 & ~x447 & ~x657 & ~x783 & ~x822 & ~x861 & ~x909 & ~x948 & ~x987 & ~x1026 & ~x1044 & ~x1065;
assign c3190 =  x2 &  x5 &  x11 &  x20 &  x26 &  x28 &  x29 &  x35 &  x38 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x71 &  x74 &  x77 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x131 &  x134 &  x140 &  x146 &  x149 &  x155 &  x158 &  x164 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x191 &  x200 &  x203 &  x209 &  x212 &  x215 &  x217 &  x218 &  x224 &  x245 &  x247 &  x248 &  x250 &  x251 &  x254 &  x257 &  x266 &  x269 &  x284 &  x289 &  x296 &  x299 &  x305 &  x308 &  x311 &  x314 &  x326 &  x332 &  x335 &  x341 &  x344 &  x347 &  x350 &  x353 &  x362 &  x368 &  x374 &  x380 &  x386 &  x389 &  x392 &  x398 &  x401 &  x407 &  x410 &  x425 &  x428 &  x433 &  x434 &  x440 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x476 &  x479 &  x482 &  x491 &  x494 &  x497 &  x503 &  x512 &  x515 &  x524 &  x527 &  x530 &  x533 &  x539 &  x545 &  x551 &  x557 &  x572 &  x590 &  x593 &  x599 &  x602 &  x605 &  x607 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x635 &  x638 &  x641 &  x644 &  x647 &  x653 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x698 &  x701 &  x707 &  x710 &  x713 &  x716 &  x719 &  x725 &  x731 &  x737 &  x746 &  x748 &  x752 &  x758 &  x770 &  x773 &  x782 &  x787 &  x797 &  x803 &  x809 &  x812 &  x821 &  x827 &  x830 &  x839 &  x842 &  x845 &  x854 &  x857 &  x860 &  x863 &  x865 &  x866 &  x869 &  x872 &  x875 &  x878 &  x887 &  x890 &  x893 &  x899 &  x904 &  x905 &  x911 &  x917 &  x920 &  x923 &  x929 &  x935 &  x938 &  x944 &  x947 &  x950 &  x953 &  x955 &  x956 &  x965 &  x968 &  x974 &  x977 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1025 &  x1028 &  x1034 &  x1037 &  x1039 &  x1040 &  x1043 &  x1046 &  x1052 &  x1058 &  x1061 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1088 &  x1094 &  x1097 &  x1100 &  x1109 &  x1115 &  x1118 &  x1124 &  x1127;
assign c3192 =  x2 &  x5 &  x8 &  x11 &  x23 &  x29 &  x32 &  x38 &  x41 &  x44 &  x56 &  x59 &  x62 &  x65 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x107 &  x110 &  x113 &  x122 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x155 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x200 &  x206 &  x209 &  x212 &  x218 &  x221 &  x224 &  x230 &  x236 &  x239 &  x242 &  x245 &  x248 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x278 &  x284 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x326 &  x329 &  x335 &  x338 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x380 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x419 &  x422 &  x428 &  x431 &  x434 &  x437 &  x443 &  x449 &  x458 &  x461 &  x464 &  x467 &  x470 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x508 &  x509 &  x512 &  x515 &  x518 &  x524 &  x527 &  x536 &  x539 &  x542 &  x551 &  x554 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x586 &  x587 &  x593 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x623 &  x625 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x659 &  x665 &  x668 &  x671 &  x674 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x707 &  x710 &  x713 &  x716 &  x722 &  x725 &  x734 &  x737 &  x740 &  x742 &  x743 &  x746 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x781 &  x782 &  x785 &  x788 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x818 &  x821 &  x824 &  x830 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x869 &  x875 &  x881 &  x884 &  x887 &  x893 &  x896 &  x901 &  x905 &  x908 &  x911 &  x914 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x950 &  x959 &  x962 &  x965 &  x971 &  x980 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1010 &  x1016 &  x1022 &  x1025 &  x1028 &  x1034 &  x1040 &  x1046 &  x1052 &  x1061 &  x1064 &  x1070 &  x1076 &  x1079 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1109 &  x1112 &  x1121 &  x1124 &  x1127 &  x1130 & ~x531 & ~x570 & ~x597 & ~x636 & ~x756 & ~x792 & ~x834 & ~x993 & ~x1026 & ~x1065 & ~x1104;
assign c3194 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x478 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x516 &  x517 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x556 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x595 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x901 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x940 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1018 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x312 & ~x348 & ~x351 & ~x387 & ~x816;
assign c3196 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x445 &  x446 &  x448 &  x449 &  x451 &  x452 &  x454 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x481 &  x482 &  x485 &  x488 &  x490 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x511 &  x512 &  x515 &  x518 &  x520 &  x521 &  x524 &  x527 &  x529 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x550 &  x551 &  x554 &  x557 &  x559 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x589 &  x590 &  x593 &  x596 &  x598 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x625 &  x626 &  x628 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x667 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x703 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x742 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x781 &  x782 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x820 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x859 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x893 &  x896 &  x899 &  x901 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x940 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130;
assign c3198 =  x23 &  x29 &  x35 &  x44 &  x56 &  x77 &  x85 &  x89 &  x101 &  x116 &  x122 &  x137 &  x143 &  x158 &  x164 &  x167 &  x206 &  x224 &  x260 &  x286 &  x314 &  x329 &  x347 &  x364 &  x389 &  x413 &  x437 &  x446 &  x455 &  x458 &  x473 &  x491 &  x500 &  x506 &  x515 &  x521 &  x533 &  x557 &  x563 &  x575 &  x608 &  x617 &  x656 &  x677 &  x695 &  x716 &  x731 &  x749 &  x758 &  x785 &  x788 &  x806 &  x812 &  x818 &  x821 &  x827 &  x839 &  x848 &  x854 &  x860 &  x911 &  x914 &  x920 &  x929 &  x950 &  x968 &  x971 &  x977 &  x980 &  x1010 &  x1016 &  x1022 &  x1034 &  x1037 &  x1040 &  x1049 &  x1109 &  x1121 & ~x118 & ~x196 & ~x228 & ~x274 & ~x313 & ~x417 & ~x969 & ~x1029;
assign c3200 =  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x101 &  x104 &  x107 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x134 &  x137 &  x143 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x206 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x448 &  x449 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x485 &  x488 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x722 &  x725 &  x728 &  x734 &  x737 &  x740 &  x743 &  x749 &  x755 &  x758 &  x764 &  x767 &  x770 &  x776 &  x779 &  x781 &  x782 &  x784 &  x785 &  x788 &  x794 &  x797 &  x800 &  x803 &  x809 &  x812 &  x815 &  x818 &  x820 &  x821 &  x823 &  x824 &  x827 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x866 &  x869 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x901 &  x902 &  x905 &  x908 &  x914 &  x917 &  x920 &  x929 &  x938 &  x940 &  x941 &  x944 &  x947 &  x950 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x976 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1018 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1057 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1085 &  x1088 &  x1091 &  x1093 &  x1094 &  x1096 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1118 &  x1124 &  x1127 &  x1130 & ~x699 & ~x738 & ~x804 & ~x843 & ~x882 & ~x921 & ~x951 & ~x960 & ~x990 & ~x993 & ~x1029 & ~x1032;
assign c3202 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x107 &  x113 &  x116 &  x119 &  x122 &  x125 &  x134 &  x137 &  x140 &  x149 &  x152 &  x155 &  x161 &  x164 &  x167 &  x170 &  x173 &  x179 &  x182 &  x185 &  x188 &  x194 &  x200 &  x203 &  x205 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x239 &  x242 &  x245 &  x248 &  x254 &  x257 &  x260 &  x263 &  x266 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x295 &  x296 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x334 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x361 &  x362 &  x368 &  x371 &  x373 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x395 &  x398 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x445 &  x449 &  x452 &  x455 &  x461 &  x467 &  x473 &  x476 &  x479 &  x481 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x506 &  x508 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x542 &  x545 &  x551 &  x554 &  x563 &  x578 &  x581 &  x586 &  x587 &  x590 &  x593 &  x596 &  x599 &  x605 &  x608 &  x611 &  x617 &  x623 &  x625 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x659 &  x662 &  x664 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x701 &  x703 &  x704 &  x713 &  x716 &  x719 &  x722 &  x725 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x764 &  x767 &  x770 &  x776 &  x781 &  x782 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x820 &  x821 &  x824 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x851 &  x854 &  x857 &  x863 &  x866 &  x869 &  x875 &  x878 &  x881 &  x890 &  x893 &  x896 &  x899 &  x901 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x938 &  x940 &  x941 &  x944 &  x950 &  x953 &  x956 &  x959 &  x968 &  x971 &  x974 &  x977 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1046 &  x1052 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x795 & ~x993;
assign c3204 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x38 &  x41 &  x44 &  x50 &  x56 &  x62 &  x65 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x134 &  x140 &  x143 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x280 &  x281 &  x290 &  x293 &  x296 &  x299 &  x305 &  x308 &  x311 &  x314 &  x317 &  x319 &  x320 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x403 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x464 &  x467 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x545 &  x548 &  x551 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x587 &  x590 &  x593 &  x596 &  x599 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x656 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x704 &  x707 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x845 &  x848 &  x851 &  x854 &  x857 &  x862 &  x863 &  x866 &  x869 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x901 &  x902 &  x905 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x940 &  x941 &  x944 &  x947 &  x953 &  x956 &  x959 &  x962 &  x965 &  x974 &  x977 &  x979 &  x980 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1018 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1055 &  x1057 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1096 &  x1097 &  x1100 &  x1103 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 & ~x159 & ~x195 & ~x234 & ~x273 & ~x312 & ~x417 & ~x456 & ~x921 & ~x960 & ~x972;
assign c3206 =  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x56 &  x68 &  x71 &  x80 &  x89 &  x92 &  x100 &  x104 &  x110 &  x112 &  x113 &  x125 &  x128 &  x131 &  x137 &  x143 &  x146 &  x151 &  x152 &  x158 &  x161 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x200 &  x209 &  x211 &  x212 &  x215 &  x239 &  x245 &  x248 &  x250 &  x256 &  x257 &  x263 &  x275 &  x284 &  x287 &  x295 &  x299 &  x305 &  x320 &  x335 &  x338 &  x341 &  x344 &  x353 &  x359 &  x362 &  x373 &  x374 &  x386 &  x389 &  x401 &  x403 &  x404 &  x409 &  x413 &  x416 &  x419 &  x422 &  x428 &  x431 &  x434 &  x440 &  x449 &  x451 &  x455 &  x458 &  x464 &  x473 &  x476 &  x481 &  x482 &  x491 &  x494 &  x509 &  x512 &  x524 &  x526 &  x530 &  x545 &  x548 &  x554 &  x556 &  x557 &  x560 &  x563 &  x566 &  x575 &  x578 &  x593 &  x596 &  x599 &  x605 &  x620 &  x623 &  x626 &  x629 &  x641 &  x644 &  x650 &  x659 &  x662 &  x665 &  x674 &  x682 &  x695 &  x701 &  x704 &  x707 &  x725 &  x731 &  x746 &  x749 &  x752 &  x755 &  x758 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x794 &  x797 &  x809 &  x818 &  x824 &  x830 &  x839 &  x842 &  x845 &  x854 &  x857 &  x859 &  x866 &  x868 &  x881 &  x887 &  x890 &  x896 &  x899 &  x929 &  x938 &  x947 &  x956 &  x964 &  x974 &  x977 &  x980 &  x992 &  x998 &  x1001 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1058 &  x1061 &  x1067 &  x1076 &  x1094 &  x1097 &  x1103 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127;
assign c3208 =  x1 &  x20 &  x23 &  x26 &  x32 &  x35 &  x41 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x74 &  x77 &  x83 &  x92 &  x95 &  x98 &  x101 &  x110 &  x113 &  x116 &  x118 &  x125 &  x128 &  x131 &  x137 &  x158 &  x161 &  x164 &  x173 &  x179 &  x182 &  x185 &  x188 &  x196 &  x206 &  x212 &  x221 &  x224 &  x233 &  x235 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x266 &  x269 &  x278 &  x281 &  x284 &  x287 &  x290 &  x296 &  x299 &  x305 &  x311 &  x313 &  x314 &  x316 &  x317 &  x320 &  x326 &  x344 &  x347 &  x350 &  x353 &  x355 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x386 &  x389 &  x392 &  x395 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x428 &  x434 &  x437 &  x440 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x467 &  x470 &  x473 &  x476 &  x482 &  x485 &  x491 &  x494 &  x500 &  x506 &  x509 &  x515 &  x521 &  x524 &  x527 &  x530 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x566 &  x569 &  x572 &  x587 &  x590 &  x593 &  x599 &  x605 &  x608 &  x620 &  x623 &  x632 &  x647 &  x650 &  x656 &  x659 &  x665 &  x668 &  x670 &  x671 &  x674 &  x680 &  x686 &  x689 &  x692 &  x698 &  x701 &  x704 &  x707 &  x712 &  x713 &  x716 &  x722 &  x725 &  x734 &  x740 &  x743 &  x748 &  x749 &  x751 &  x752 &  x755 &  x761 &  x764 &  x767 &  x770 &  x773 &  x782 &  x785 &  x788 &  x791 &  x797 &  x800 &  x803 &  x809 &  x812 &  x815 &  x824 &  x827 &  x842 &  x845 &  x848 &  x851 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x899 &  x902 &  x914 &  x917 &  x920 &  x923 &  x932 &  x944 &  x947 &  x950 &  x953 &  x956 &  x965 &  x971 &  x974 &  x980 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1016 &  x1019 &  x1022 &  x1028 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1088 &  x1091 &  x1097 &  x1106 &  x1109 &  x1115 &  x1118 &  x1124 &  x1127 &  x1130 & ~x663 & ~x702 & ~x741 & ~x780 & ~x837 & ~x1110;
assign c3210 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x298 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x337 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x364 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x403 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x442 &  x443 &  x446 &  x449 &  x452 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1060 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 &  x1130 & ~x3 & ~x42 & ~x81 & ~x82 & ~x120 & ~x121 & ~x159 & ~x160 & ~x198 & ~x237;
assign c3212 =  x2 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x29 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x77 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x140 &  x143 &  x148 &  x152 &  x155 &  x161 &  x164 &  x170 &  x176 &  x179 &  x182 &  x185 &  x191 &  x193 &  x194 &  x197 &  x203 &  x206 &  x209 &  x215 &  x224 &  x226 &  x227 &  x230 &  x232 &  x236 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x265 &  x266 &  x281 &  x284 &  x287 &  x290 &  x296 &  x299 &  x304 &  x305 &  x308 &  x314 &  x320 &  x323 &  x326 &  x329 &  x331 &  x332 &  x338 &  x347 &  x350 &  x353 &  x359 &  x362 &  x365 &  x370 &  x371 &  x374 &  x386 &  x389 &  x395 &  x403 &  x409 &  x410 &  x413 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x440 &  x442 &  x443 &  x446 &  x448 &  x455 &  x458 &  x461 &  x467 &  x470 &  x478 &  x479 &  x482 &  x485 &  x487 &  x491 &  x494 &  x497 &  x500 &  x506 &  x512 &  x515 &  x517 &  x518 &  x521 &  x527 &  x536 &  x539 &  x542 &  x545 &  x554 &  x557 &  x563 &  x566 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x629 &  x632 &  x638 &  x641 &  x643 &  x644 &  x650 &  x665 &  x674 &  x677 &  x680 &  x683 &  x689 &  x692 &  x695 &  x701 &  x704 &  x710 &  x716 &  x722 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x767 &  x770 &  x773 &  x776 &  x779 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x824 &  x833 &  x836 &  x842 &  x845 &  x848 &  x854 &  x857 &  x860 &  x866 &  x878 &  x884 &  x887 &  x893 &  x902 &  x905 &  x908 &  x914 &  x917 &  x920 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x956 &  x959 &  x965 &  x974 &  x977 &  x983 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1064 &  x1067 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130 & ~x312 & ~x390 & ~x834 & ~x873;
assign c3214 =  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x35 &  x41 &  x44 &  x47 &  x50 &  x56 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x95 &  x98 &  x107 &  x110 &  x113 &  x116 &  x122 &  x125 &  x128 &  x131 &  x134 &  x143 &  x146 &  x149 &  x155 &  x158 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x188 &  x191 &  x194 &  x203 &  x209 &  x212 &  x215 &  x218 &  x224 &  x230 &  x236 &  x239 &  x245 &  x248 &  x251 &  x254 &  x260 &  x263 &  x269 &  x272 &  x275 &  x281 &  x287 &  x290 &  x293 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x326 &  x329 &  x344 &  x347 &  x356 &  x359 &  x365 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x395 &  x398 &  x416 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x449 &  x455 &  x458 &  x461 &  x473 &  x476 &  x485 &  x488 &  x491 &  x494 &  x500 &  x512 &  x518 &  x521 &  x527 &  x533 &  x539 &  x542 &  x545 &  x548 &  x557 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x626 &  x632 &  x635 &  x638 &  x641 &  x647 &  x650 &  x653 &  x662 &  x665 &  x668 &  x671 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x704 &  x713 &  x716 &  x719 &  x725 &  x734 &  x737 &  x740 &  x749 &  x755 &  x767 &  x773 &  x776 &  x782 &  x784 &  x785 &  x791 &  x794 &  x797 &  x800 &  x803 &  x815 &  x818 &  x821 &  x827 &  x830 &  x833 &  x836 &  x839 &  x845 &  x851 &  x860 &  x862 &  x863 &  x872 &  x875 &  x881 &  x887 &  x890 &  x893 &  x896 &  x902 &  x914 &  x917 &  x926 &  x935 &  x941 &  x944 &  x947 &  x953 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x992 &  x995 &  x1007 &  x1013 &  x1019 &  x1025 &  x1028 &  x1040 &  x1043 &  x1046 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1118 &  x1124 &  x1130 & ~x27 & ~x66 & ~x105 & ~x183 & ~x234 & ~x261 & ~x300 & ~x339 & ~x378 & ~x840 & ~x918 & ~x1038 & ~x1074 & ~x1107 & ~x1128;
assign c3216 =  x8 &  x11 &  x17 &  x20 &  x26 &  x29 &  x32 &  x34 &  x35 &  x38 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x73 &  x77 &  x80 &  x83 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x116 &  x119 &  x122 &  x125 &  x128 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x263 &  x266 &  x269 &  x272 &  x281 &  x284 &  x287 &  x290 &  x299 &  x302 &  x305 &  x308 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x428 &  x431 &  x433 &  x434 &  x437 &  x443 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x479 &  x485 &  x488 &  x497 &  x506 &  x509 &  x515 &  x524 &  x527 &  x530 &  x536 &  x542 &  x545 &  x548 &  x554 &  x557 &  x563 &  x566 &  x569 &  x572 &  x578 &  x584 &  x586 &  x590 &  x596 &  x602 &  x605 &  x611 &  x617 &  x625 &  x626 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x674 &  x677 &  x686 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x737 &  x743 &  x746 &  x749 &  x752 &  x758 &  x761 &  x764 &  x767 &  x770 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x797 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x833 &  x836 &  x839 &  x842 &  x848 &  x851 &  x854 &  x857 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x901 &  x902 &  x905 &  x911 &  x914 &  x920 &  x923 &  x929 &  x935 &  x938 &  x941 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1016 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x609 & ~x648 & ~x675 & ~x687 & ~x726 & ~x792 & ~x795 & ~x834;
assign c3218 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x95 &  x98 &  x101 &  x107 &  x110 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x236 &  x239 &  x242 &  x244 &  x245 &  x248 &  x250 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x283 &  x284 &  x287 &  x289 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x316 &  x317 &  x320 &  x321 &  x322 &  x323 &  x326 &  x328 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x355 &  x356 &  x359 &  x361 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x391 &  x392 &  x394 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x430 &  x431 &  x433 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x469 &  x470 &  x472 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x508 &  x509 &  x511 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x547 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x589 &  x590 &  x593 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x628 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x667 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x869 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x905 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130;
assign c3220 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x41 &  x47 &  x50 &  x53 &  x56 &  x62 &  x65 &  x68 &  x77 &  x80 &  x89 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x131 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x356 &  x359 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x404 &  x407 &  x410 &  x413 &  x419 &  x425 &  x437 &  x440 &  x443 &  x446 &  x449 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x482 &  x484 &  x485 &  x488 &  x491 &  x494 &  x503 &  x506 &  x509 &  x527 &  x533 &  x536 &  x542 &  x545 &  x551 &  x560 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x590 &  x593 &  x596 &  x599 &  x602 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x656 &  x659 &  x662 &  x671 &  x672 &  x673 &  x674 &  x677 &  x680 &  x682 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x706 &  x707 &  x710 &  x712 &  x713 &  x716 &  x719 &  x722 &  x725 &  x731 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x773 &  x776 &  x779 &  x781 &  x782 &  x784 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x809 &  x812 &  x820 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x898 &  x901 &  x902 &  x905 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x937 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x977 &  x979 &  x980 &  x983 &  x986 &  x989 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1018 &  x1019 &  x1025 &  x1028 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1057 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130;
assign c3222 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x481 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x509 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x781 &  x782 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x820 &  x821 &  x823 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x859 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x901 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x273 & ~x312 & ~x351 & ~x612 & ~x651 & ~x993 & ~x1032 & ~x1044 & ~x1068 & ~x1083 & ~x1107 & ~x1122;
assign c3224 =  x13 &  x14 &  x41 &  x44 &  x77 &  x83 &  x92 &  x104 &  x122 &  x128 &  x149 &  x152 &  x155 &  x194 &  x203 &  x218 &  x227 &  x248 &  x272 &  x275 &  x284 &  x296 &  x308 &  x315 &  x392 &  x413 &  x428 &  x431 &  x443 &  x446 &  x475 &  x482 &  x491 &  x503 &  x521 &  x530 &  x554 &  x578 &  x581 &  x587 &  x602 &  x605 &  x608 &  x617 &  x620 &  x623 &  x659 &  x686 &  x694 &  x695 &  x722 &  x743 &  x755 &  x776 &  x779 &  x782 &  x788 &  x800 &  x830 &  x890 &  x893 &  x917 &  x920 &  x932 &  x950 &  x980 &  x992 &  x995 &  x998 &  x1013 &  x1019 &  x1025 &  x1058 &  x1061 &  x1073 &  x1100 &  x1115 & ~x225 & ~x405 & ~x406 & ~x444 & ~x702 & ~x819 & ~x936;
assign c3226 =  x2 &  x5 &  x8 &  x17 &  x20 &  x26 &  x35 &  x38 &  x41 &  x44 &  x50 &  x53 &  x59 &  x62 &  x68 &  x74 &  x80 &  x83 &  x86 &  x89 &  x95 &  x98 &  x104 &  x110 &  x113 &  x119 &  x122 &  x125 &  x128 &  x134 &  x137 &  x140 &  x146 &  x149 &  x152 &  x158 &  x164 &  x167 &  x170 &  x176 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x212 &  x224 &  x227 &  x230 &  x233 &  x239 &  x245 &  x248 &  x251 &  x260 &  x263 &  x266 &  x269 &  x272 &  x278 &  x281 &  x287 &  x293 &  x299 &  x302 &  x305 &  x311 &  x314 &  x317 &  x320 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x419 &  x425 &  x431 &  x437 &  x440 &  x446 &  x449 &  x455 &  x458 &  x461 &  x467 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x530 &  x533 &  x536 &  x538 &  x542 &  x545 &  x548 &  x551 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x577 &  x581 &  x584 &  x590 &  x593 &  x595 &  x599 &  x605 &  x608 &  x611 &  x614 &  x616 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x647 &  x650 &  x653 &  x655 &  x656 &  x659 &  x662 &  x665 &  x668 &  x677 &  x680 &  x683 &  x686 &  x692 &  x694 &  x695 &  x698 &  x701 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x743 &  x749 &  x755 &  x761 &  x767 &  x770 &  x776 &  x779 &  x785 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x845 &  x848 &  x851 &  x857 &  x860 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x926 &  x929 &  x932 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x977 &  x980 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1022 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x123 & ~x162 & ~x465 & ~x543 & ~x582 & ~x792 & ~x948 & ~x1065 & ~x1104;
assign c3228 =  x2 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x113 &  x116 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x322 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x360 &  x361 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x383 &  x386 &  x389 &  x400 &  x401 &  x403 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x434 &  x437 &  x440 &  x442 &  x443 &  x449 &  x452 &  x455 &  x461 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x494 &  x497 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x565 &  x566 &  x569 &  x572 &  x575 &  x578 &  x584 &  x593 &  x596 &  x599 &  x602 &  x604 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x626 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x656 &  x659 &  x671 &  x674 &  x677 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x707 &  x710 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x749 &  x752 &  x755 &  x761 &  x764 &  x767 &  x770 &  x773 &  x779 &  x782 &  x785 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x860 &  x863 &  x866 &  x872 &  x878 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x908 &  x911 &  x914 &  x917 &  x920 &  x922 &  x923 &  x926 &  x929 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1000 &  x1001 &  x1004 &  x1007 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1049 &  x1052 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x84;
assign c3230 =  x17 &  x44 &  x50 &  x56 &  x65 &  x68 &  x86 &  x92 &  x95 &  x107 &  x110 &  x113 &  x122 &  x128 &  x131 &  x134 &  x143 &  x155 &  x158 &  x166 &  x170 &  x172 &  x173 &  x188 &  x194 &  x205 &  x209 &  x211 &  x212 &  x215 &  x218 &  x221 &  x236 &  x245 &  x250 &  x254 &  x257 &  x275 &  x287 &  x296 &  x313 &  x314 &  x317 &  x320 &  x321 &  x323 &  x326 &  x332 &  x338 &  x341 &  x347 &  x352 &  x356 &  x361 &  x365 &  x377 &  x392 &  x398 &  x407 &  x416 &  x419 &  x428 &  x430 &  x440 &  x443 &  x452 &  x470 &  x479 &  x482 &  x494 &  x500 &  x508 &  x515 &  x518 &  x524 &  x530 &  x536 &  x542 &  x563 &  x569 &  x572 &  x602 &  x605 &  x608 &  x617 &  x620 &  x626 &  x659 &  x662 &  x683 &  x686 &  x692 &  x712 &  x716 &  x719 &  x722 &  x728 &  x734 &  x737 &  x740 &  x749 &  x764 &  x776 &  x779 &  x788 &  x790 &  x791 &  x800 &  x803 &  x812 &  x818 &  x821 &  x829 &  x830 &  x836 &  x848 &  x854 &  x866 &  x884 &  x890 &  x902 &  x905 &  x908 &  x926 &  x938 &  x956 &  x964 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1003 &  x1004 &  x1010 &  x1030 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1070 &  x1073 &  x1081 &  x1085 &  x1087 &  x1112;
assign c3232 =  x2 &  x5 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x131 &  x137 &  x143 &  x146 &  x151 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x197 &  x200 &  x203 &  x206 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x239 &  x242 &  x245 &  x248 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x283 &  x287 &  x290 &  x293 &  x296 &  x302 &  x311 &  x314 &  x316 &  x317 &  x320 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x356 &  x359 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x386 &  x392 &  x395 &  x398 &  x400 &  x401 &  x404 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x452 &  x455 &  x458 &  x464 &  x470 &  x476 &  x479 &  x482 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x530 &  x533 &  x536 &  x539 &  x542 &  x548 &  x551 &  x554 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x596 &  x602 &  x608 &  x611 &  x614 &  x620 &  x623 &  x626 &  x629 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x737 &  x740 &  x746 &  x749 &  x751 &  x752 &  x755 &  x761 &  x770 &  x773 &  x779 &  x782 &  x785 &  x787 &  x788 &  x791 &  x794 &  x803 &  x812 &  x815 &  x821 &  x826 &  x827 &  x833 &  x836 &  x839 &  x845 &  x848 &  x851 &  x854 &  x856 &  x857 &  x860 &  x866 &  x869 &  x872 &  x875 &  x878 &  x884 &  x890 &  x893 &  x895 &  x896 &  x902 &  x908 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x934 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x983 &  x986 &  x989 &  x995 &  x998 &  x1004 &  x1010 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1124 &  x1127 & ~x414 & ~x483;
assign c3234 =  x5 &  x11 &  x17 &  x23 &  x41 &  x44 &  x50 &  x59 &  x62 &  x71 &  x74 &  x80 &  x83 &  x107 &  x110 &  x113 &  x119 &  x131 &  x146 &  x149 &  x152 &  x161 &  x167 &  x170 &  x176 &  x185 &  x194 &  x197 &  x200 &  x203 &  x212 &  x218 &  x221 &  x223 &  x230 &  x236 &  x251 &  x257 &  x260 &  x263 &  x266 &  x272 &  x281 &  x284 &  x290 &  x299 &  x302 &  x341 &  x344 &  x356 &  x359 &  x365 &  x371 &  x374 &  x380 &  x386 &  x389 &  x392 &  x398 &  x407 &  x419 &  x422 &  x428 &  x431 &  x437 &  x440 &  x458 &  x467 &  x479 &  x490 &  x506 &  x509 &  x515 &  x524 &  x527 &  x528 &  x548 &  x551 &  x557 &  x563 &  x568 &  x569 &  x581 &  x590 &  x599 &  x607 &  x608 &  x611 &  x626 &  x629 &  x638 &  x641 &  x656 &  x662 &  x667 &  x668 &  x671 &  x680 &  x686 &  x689 &  x695 &  x701 &  x710 &  x719 &  x731 &  x734 &  x737 &  x749 &  x755 &  x758 &  x761 &  x767 &  x770 &  x776 &  x791 &  x800 &  x812 &  x827 &  x833 &  x851 &  x857 &  x863 &  x872 &  x875 &  x881 &  x884 &  x887 &  x893 &  x905 &  x914 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x941 &  x947 &  x974 &  x977 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1004 &  x1007 &  x1009 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1055 &  x1061 &  x1073 &  x1094 &  x1106 &  x1109 &  x1118 &  x1124 & ~x795 & ~x834;
assign c3236 =  x2 &  x8 &  x11 &  x13 &  x14 &  x17 &  x23 &  x29 &  x32 &  x38 &  x44 &  x47 &  x52 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x83 &  x86 &  x89 &  x92 &  x95 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x143 &  x149 &  x152 &  x155 &  x164 &  x167 &  x179 &  x182 &  x188 &  x191 &  x197 &  x200 &  x206 &  x209 &  x212 &  x218 &  x224 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x260 &  x263 &  x266 &  x269 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x308 &  x311 &  x316 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x353 &  x355 &  x356 &  x359 &  x362 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x395 &  x404 &  x407 &  x416 &  x419 &  x425 &  x433 &  x437 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x472 &  x475 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x503 &  x506 &  x509 &  x511 &  x513 &  x518 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x551 &  x553 &  x554 &  x557 &  x560 &  x569 &  x572 &  x575 &  x578 &  x584 &  x590 &  x592 &  x593 &  x596 &  x598 &  x599 &  x605 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x631 &  x637 &  x644 &  x647 &  x650 &  x652 &  x656 &  x659 &  x662 &  x665 &  x668 &  x670 &  x671 &  x674 &  x676 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x713 &  x715 &  x716 &  x728 &  x737 &  x743 &  x746 &  x749 &  x752 &  x754 &  x755 &  x758 &  x761 &  x764 &  x770 &  x773 &  x779 &  x782 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x827 &  x830 &  x839 &  x842 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x893 &  x899 &  x902 &  x905 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x944 &  x947 &  x950 &  x953 &  x956 &  x962 &  x965 &  x968 &  x974 &  x977 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1046 &  x1049 &  x1058 &  x1061 &  x1067 &  x1073 &  x1082 &  x1085 &  x1094 &  x1097 &  x1100 &  x1109 &  x1112 &  x1118 &  x1121 &  x1127 &  x1130 & ~x546 & ~x585 & ~x624 & ~x664 & ~x702 & ~x741 & ~x780 & ~x936 & ~x975 & ~x1014;
assign c3238 =  x2 &  x8 &  x10 &  x17 &  x20 &  x32 &  x35 &  x41 &  x77 &  x83 &  x89 &  x95 &  x98 &  x101 &  x104 &  x107 &  x116 &  x125 &  x128 &  x131 &  x140 &  x146 &  x149 &  x152 &  x158 &  x164 &  x170 &  x176 &  x179 &  x185 &  x191 &  x197 &  x200 &  x215 &  x218 &  x221 &  x227 &  x236 &  x239 &  x242 &  x248 &  x254 &  x260 &  x263 &  x269 &  x272 &  x278 &  x281 &  x284 &  x293 &  x299 &  x311 &  x314 &  x320 &  x322 &  x323 &  x329 &  x332 &  x341 &  x344 &  x347 &  x353 &  x355 &  x356 &  x361 &  x365 &  x374 &  x380 &  x383 &  x386 &  x389 &  x392 &  x394 &  x395 &  x398 &  x399 &  x401 &  x416 &  x422 &  x425 &  x431 &  x433 &  x434 &  x438 &  x439 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x472 &  x473 &  x494 &  x500 &  x509 &  x515 &  x517 &  x530 &  x533 &  x536 &  x542 &  x560 &  x569 &  x575 &  x578 &  x584 &  x587 &  x593 &  x596 &  x602 &  x608 &  x614 &  x617 &  x623 &  x626 &  x632 &  x638 &  x641 &  x647 &  x656 &  x665 &  x674 &  x680 &  x683 &  x704 &  x707 &  x716 &  x719 &  x722 &  x725 &  x737 &  x752 &  x758 &  x764 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x797 &  x800 &  x803 &  x809 &  x818 &  x821 &  x824 &  x833 &  x836 &  x842 &  x845 &  x848 &  x851 &  x854 &  x860 &  x863 &  x869 &  x887 &  x896 &  x920 &  x923 &  x929 &  x931 &  x944 &  x965 &  x971 &  x977 &  x980 &  x986 &  x989 &  x995 &  x1001 &  x1016 &  x1019 &  x1022 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1082 &  x1091 &  x1097 &  x1100 &  x1103 &  x1109 &  x1118 &  x1121 &  x1130 & ~x225;
assign c3240 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x23 &  x26 &  x32 &  x35 &  x38 &  x41 &  x44 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x101 &  x104 &  x107 &  x116 &  x119 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x146 &  x149 &  x155 &  x158 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x200 &  x206 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x269 &  x272 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x395 &  x398 &  x401 &  x407 &  x410 &  x416 &  x419 &  x425 &  x428 &  x434 &  x440 &  x442 &  x448 &  x449 &  x452 &  x455 &  x458 &  x461 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x494 &  x497 &  x500 &  x506 &  x509 &  x512 &  x515 &  x518 &  x520 &  x521 &  x524 &  x526 &  x527 &  x530 &  x533 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x559 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x587 &  x590 &  x596 &  x598 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x629 &  x635 &  x637 &  x638 &  x644 &  x650 &  x653 &  x656 &  x662 &  x671 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x706 &  x710 &  x713 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x745 &  x746 &  x749 &  x752 &  x758 &  x761 &  x764 &  x767 &  x776 &  x779 &  x782 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x815 &  x818 &  x823 &  x824 &  x827 &  x830 &  x839 &  x842 &  x848 &  x851 &  x854 &  x857 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x896 &  x899 &  x901 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x940 &  x944 &  x950 &  x959 &  x962 &  x971 &  x974 &  x977 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x1001 &  x1007 &  x1013 &  x1016 &  x1018 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1057 &  x1061 &  x1064 &  x1067 &  x1070 &  x1079 &  x1082 &  x1085 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1130 & ~x156 & ~x195 & ~x234 & ~x273 & ~x312 & ~x351 & ~x390 & ~x429 & ~x468 & ~x651 & ~x765 & ~x951 & ~x990 & ~x1029;
assign c3242 =  x2 &  x8 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x41 &  x50 &  x53 &  x74 &  x77 &  x83 &  x86 &  x95 &  x101 &  x104 &  x113 &  x116 &  x125 &  x128 &  x134 &  x152 &  x167 &  x173 &  x179 &  x182 &  x194 &  x197 &  x199 &  x200 &  x212 &  x215 &  x218 &  x224 &  x236 &  x238 &  x245 &  x251 &  x257 &  x269 &  x272 &  x277 &  x281 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x314 &  x320 &  x326 &  x350 &  x355 &  x356 &  x365 &  x380 &  x401 &  x413 &  x425 &  x433 &  x440 &  x443 &  x449 &  x452 &  x455 &  x458 &  x464 &  x479 &  x482 &  x497 &  x503 &  x509 &  x521 &  x524 &  x530 &  x539 &  x548 &  x551 &  x557 &  x566 &  x569 &  x572 &  x581 &  x584 &  x590 &  x592 &  x605 &  x611 &  x617 &  x620 &  x623 &  x631 &  x632 &  x635 &  x638 &  x644 &  x659 &  x668 &  x670 &  x674 &  x677 &  x683 &  x686 &  x689 &  x701 &  x704 &  x709 &  x725 &  x728 &  x746 &  x758 &  x764 &  x767 &  x773 &  x779 &  x785 &  x797 &  x800 &  x805 &  x806 &  x812 &  x824 &  x827 &  x830 &  x836 &  x848 &  x851 &  x854 &  x863 &  x872 &  x890 &  x893 &  x896 &  x902 &  x908 &  x911 &  x914 &  x929 &  x938 &  x941 &  x947 &  x959 &  x962 &  x977 &  x995 &  x1001 &  x1010 &  x1019 &  x1037 &  x1040 &  x1046 &  x1052 &  x1058 &  x1061 &  x1064 &  x1073 &  x1076 &  x1091 &  x1103 &  x1112 &  x1115 &  x1118 &  x1130 & ~x483 & ~x624 & ~x625 & ~x663 & ~x702 & ~x703 & ~x742 & ~x780 & ~x783 & ~x862 & ~x897 & ~x900 & ~x936 & ~x1014 & ~x1092;
assign c3244 =  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x89 &  x92 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x197 &  x203 &  x206 &  x209 &  x218 &  x221 &  x224 &  x227 &  x230 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x266 &  x272 &  x275 &  x281 &  x284 &  x287 &  x296 &  x299 &  x302 &  x308 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x350 &  x353 &  x355 &  x362 &  x374 &  x380 &  x386 &  x389 &  x392 &  x394 &  x398 &  x401 &  x404 &  x407 &  x410 &  x416 &  x419 &  x425 &  x428 &  x431 &  x433 &  x434 &  x437 &  x440 &  x443 &  x449 &  x452 &  x455 &  x458 &  x464 &  x467 &  x470 &  x472 &  x473 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x509 &  x511 &  x512 &  x515 &  x518 &  x521 &  x524 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x550 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x572 &  x575 &  x578 &  x581 &  x584 &  x589 &  x590 &  x596 &  x599 &  x605 &  x608 &  x611 &  x620 &  x623 &  x626 &  x629 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x709 &  x716 &  x719 &  x728 &  x737 &  x743 &  x748 &  x749 &  x752 &  x755 &  x761 &  x767 &  x770 &  x773 &  x776 &  x778 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x806 &  x812 &  x818 &  x833 &  x836 &  x839 &  x845 &  x848 &  x854 &  x856 &  x857 &  x860 &  x866 &  x875 &  x881 &  x887 &  x893 &  x895 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x929 &  x938 &  x941 &  x944 &  x956 &  x959 &  x962 &  x965 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1130 & ~x342 & ~x663 & ~x702 & ~x741 & ~x780 & ~x819 & ~x1104;
assign c3246 =  x2 &  x11 &  x14 &  x17 &  x20 &  x35 &  x41 &  x44 &  x47 &  x50 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x104 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x134 &  x137 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x212 &  x215 &  x218 &  x221 &  x227 &  x236 &  x239 &  x242 &  x248 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x277 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x316 &  x320 &  x323 &  x326 &  x329 &  x332 &  x338 &  x347 &  x350 &  x356 &  x359 &  x371 &  x374 &  x377 &  x380 &  x389 &  x392 &  x394 &  x395 &  x398 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x433 &  x434 &  x440 &  x443 &  x446 &  x449 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x482 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x509 &  x512 &  x517 &  x518 &  x524 &  x530 &  x536 &  x539 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x599 &  x602 &  x608 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x644 &  x647 &  x653 &  x656 &  x659 &  x665 &  x668 &  x670 &  x680 &  x686 &  x689 &  x692 &  x707 &  x709 &  x710 &  x716 &  x719 &  x722 &  x725 &  x731 &  x737 &  x739 &  x746 &  x749 &  x752 &  x758 &  x761 &  x764 &  x767 &  x773 &  x776 &  x782 &  x785 &  x787 &  x788 &  x797 &  x803 &  x815 &  x818 &  x821 &  x830 &  x833 &  x845 &  x848 &  x851 &  x854 &  x856 &  x857 &  x860 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x890 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x920 &  x926 &  x929 &  x932 &  x934 &  x935 &  x938 &  x947 &  x950 &  x956 &  x959 &  x965 &  x971 &  x974 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1016 &  x1019 &  x1022 &  x1031 &  x1034 &  x1040 &  x1043 &  x1049 &  x1052 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1127 &  x1130 & ~x150 & ~x600 & ~x663 & ~x702 & ~x717 & ~x741 & ~x819 & ~x858 & ~x891 & ~x936 & ~x951;
assign c3248 =  x8 &  x20 &  x23 &  x32 &  x38 &  x65 &  x68 &  x71 &  x74 &  x95 &  x101 &  x110 &  x116 &  x128 &  x131 &  x146 &  x149 &  x152 &  x191 &  x206 &  x215 &  x224 &  x245 &  x275 &  x281 &  x284 &  x287 &  x293 &  x296 &  x302 &  x314 &  x317 &  x322 &  x329 &  x347 &  x353 &  x356 &  x360 &  x383 &  x392 &  x400 &  x437 &  x452 &  x464 &  x494 &  x518 &  x524 &  x584 &  x611 &  x617 &  x623 &  x626 &  x632 &  x641 &  x665 &  x671 &  x677 &  x683 &  x689 &  x692 &  x695 &  x704 &  x716 &  x719 &  x737 &  x743 &  x752 &  x761 &  x770 &  x776 &  x779 &  x788 &  x797 &  x800 &  x812 &  x815 &  x823 &  x827 &  x830 &  x833 &  x836 &  x850 &  x857 &  x860 &  x867 &  x869 &  x878 &  x890 &  x896 &  x905 &  x908 &  x926 &  x935 &  x968 &  x971 &  x977 &  x980 &  x992 &  x998 &  x1019 &  x1025 &  x1028 &  x1037 &  x1049 &  x1052 &  x1064 &  x1070 &  x1076 &  x1094 &  x1097 &  x1112;
assign c3250 =  x2 &  x8 &  x11 &  x20 &  x23 &  x26 &  x35 &  x38 &  x41 &  x44 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x80 &  x83 &  x86 &  x107 &  x110 &  x113 &  x116 &  x122 &  x125 &  x128 &  x134 &  x140 &  x143 &  x146 &  x152 &  x155 &  x161 &  x173 &  x176 &  x179 &  x197 &  x203 &  x215 &  x224 &  x233 &  x236 &  x239 &  x248 &  x251 &  x254 &  x260 &  x263 &  x269 &  x272 &  x278 &  x281 &  x284 &  x293 &  x299 &  x305 &  x314 &  x317 &  x322 &  x323 &  x326 &  x335 &  x338 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x380 &  x383 &  x389 &  x398 &  x404 &  x407 &  x410 &  x413 &  x416 &  x425 &  x431 &  x440 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x478 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x512 &  x518 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x590 &  x596 &  x599 &  x605 &  x607 &  x608 &  x614 &  x617 &  x623 &  x629 &  x632 &  x635 &  x638 &  x644 &  x647 &  x653 &  x659 &  x665 &  x668 &  x671 &  x673 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x707 &  x710 &  x712 &  x713 &  x719 &  x722 &  x731 &  x734 &  x737 &  x746 &  x749 &  x755 &  x758 &  x764 &  x773 &  x776 &  x782 &  x788 &  x791 &  x794 &  x797 &  x803 &  x809 &  x812 &  x815 &  x818 &  x824 &  x830 &  x836 &  x839 &  x842 &  x848 &  x854 &  x857 &  x866 &  x868 &  x869 &  x875 &  x878 &  x887 &  x893 &  x907 &  x911 &  x917 &  x923 &  x938 &  x950 &  x956 &  x965 &  x968 &  x983 &  x986 &  x995 &  x998 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1064 &  x1076 &  x1079 &  x1082 &  x1088 &  x1100 &  x1106 &  x1109 &  x1118 &  x1124 &  x1127 &  x1130 & ~x84 & ~x387 & ~x471 & ~x552 & ~x591 & ~x630;
assign c3252 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x56 &  x62 &  x65 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x209 &  x212 &  x215 &  x218 &  x221 &  x227 &  x230 &  x236 &  x245 &  x248 &  x251 &  x254 &  x257 &  x263 &  x266 &  x269 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x302 &  x305 &  x308 &  x311 &  x314 &  x320 &  x326 &  x329 &  x331 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x359 &  x362 &  x368 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x401 &  x407 &  x410 &  x413 &  x416 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x452 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x482 &  x485 &  x488 &  x491 &  x497 &  x500 &  x503 &  x509 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x545 &  x548 &  x551 &  x560 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x593 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x662 &  x665 &  x668 &  x671 &  x674 &  x680 &  x686 &  x689 &  x692 &  x698 &  x701 &  x704 &  x707 &  x713 &  x716 &  x722 &  x725 &  x734 &  x740 &  x743 &  x746 &  x752 &  x755 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x784 &  x785 &  x788 &  x790 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x821 &  x823 &  x824 &  x827 &  x829 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x896 &  x899 &  x905 &  x908 &  x911 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x977 &  x980 &  x983 &  x986 &  x992 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x27 & ~x66 & ~x78 & ~x117 & ~x156 & ~x195 & ~x228 & ~x234 & ~x339 & ~x378 & ~x417 & ~x474 & ~x513;
assign c3254 =  x10 &  x11 &  x17 &  x20 &  x29 &  x44 &  x53 &  x56 &  x74 &  x80 &  x83 &  x95 &  x107 &  x116 &  x125 &  x131 &  x134 &  x158 &  x170 &  x179 &  x197 &  x212 &  x224 &  x239 &  x266 &  x274 &  x275 &  x281 &  x305 &  x313 &  x335 &  x350 &  x356 &  x365 &  x398 &  x413 &  x416 &  x422 &  x425 &  x491 &  x497 &  x512 &  x527 &  x533 &  x536 &  x575 &  x593 &  x596 &  x611 &  x629 &  x631 &  x635 &  x644 &  x647 &  x649 &  x670 &  x680 &  x686 &  x709 &  x710 &  x722 &  x725 &  x764 &  x766 &  x770 &  x797 &  x806 &  x818 &  x844 &  x848 &  x854 &  x869 &  x875 &  x878 &  x887 &  x890 &  x902 &  x905 &  x932 &  x938 &  x947 &  x950 &  x995 &  x1001 &  x1019 &  x1022 &  x1031 &  x1049 &  x1070 &  x1073 &  x1076 &  x1091 &  x1097 &  x1106 &  x1109 &  x1115 &  x1130 & ~x123 & ~x162 & ~x489 & ~x936 & ~x1053;
assign c3256 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x47 &  x50 &  x53 &  x56 &  x59 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x206 &  x209 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x317 &  x320 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x521 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x550 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x584 &  x587 &  x589 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x614 &  x617 &  x620 &  x623 &  x626 &  x628 &  x629 &  x632 &  x635 &  x638 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x667 &  x668 &  x671 &  x674 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x706 &  x707 &  x710 &  x713 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x743 &  x746 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x823 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x977 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x156 & ~x195 & ~x765 & ~x951 & ~x990 & ~x991 & ~x1029 & ~x1030 & ~x1035 & ~x1068 & ~x1074 & ~x1107 & ~x1113;
assign c3258 =  x2 &  x4 &  x11 &  x17 &  x23 &  x26 &  x32 &  x41 &  x43 &  x50 &  x53 &  x59 &  x62 &  x65 &  x68 &  x77 &  x80 &  x89 &  x92 &  x95 &  x98 &  x104 &  x113 &  x116 &  x119 &  x121 &  x125 &  x127 &  x128 &  x131 &  x134 &  x143 &  x146 &  x149 &  x161 &  x164 &  x166 &  x167 &  x170 &  x182 &  x185 &  x188 &  x191 &  x205 &  x209 &  x212 &  x215 &  x218 &  x221 &  x227 &  x230 &  x233 &  x238 &  x239 &  x242 &  x263 &  x272 &  x278 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x344 &  x347 &  x350 &  x353 &  x356 &  x362 &  x368 &  x371 &  x377 &  x380 &  x389 &  x392 &  x395 &  x401 &  x404 &  x410 &  x413 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x467 &  x470 &  x479 &  x482 &  x488 &  x491 &  x494 &  x497 &  x500 &  x506 &  x509 &  x511 &  x512 &  x518 &  x521 &  x527 &  x530 &  x539 &  x542 &  x545 &  x548 &  x551 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x581 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x656 &  x659 &  x662 &  x668 &  x677 &  x680 &  x686 &  x689 &  x692 &  x701 &  x704 &  x710 &  x716 &  x728 &  x734 &  x737 &  x746 &  x749 &  x752 &  x758 &  x761 &  x767 &  x770 &  x776 &  x782 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x821 &  x824 &  x836 &  x839 &  x842 &  x848 &  x854 &  x857 &  x860 &  x866 &  x875 &  x881 &  x884 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x959 &  x965 &  x968 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1043 &  x1049 &  x1058 &  x1061 &  x1067 &  x1070 &  x1076 &  x1079 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1124 &  x1127 & ~x36 & ~x37 & ~x927;
assign c3260 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x392 &  x395 &  x398 &  x401 &  x403 &  x404 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x442 &  x443 &  x446 &  x449 &  x452 &  x454 &  x455 &  x458 &  x460 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x481 &  x482 &  x484 &  x485 &  x488 &  x491 &  x493 &  x494 &  x497 &  x499 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x520 &  x521 &  x524 &  x527 &  x530 &  x532 &  x533 &  x536 &  x538 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x559 &  x560 &  x563 &  x566 &  x569 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x597 &  x598 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x637 &  x638 &  x641 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x731 &  x734 &  x737 &  x740 &  x743 &  x745 &  x746 &  x749 &  x752 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x901 &  x905 &  x908 &  x911 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x938 &  x940 &  x941 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x971 &  x974 &  x977 &  x979 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1018 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1057 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1096 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 & ~x990;
assign c3262 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x394 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x433 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x472 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x511 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x550 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x589 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x625 &  x626 &  x628 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x667 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x609 & ~x648 & ~x687 & ~x717 & ~x726 & ~x756 & ~x765 & ~x795 & ~x990 & ~x1029 & ~x1068;
assign c3264 =  x2 &  x23 &  x26 &  x29 &  x32 &  x44 &  x47 &  x50 &  x62 &  x65 &  x80 &  x86 &  x104 &  x110 &  x116 &  x119 &  x122 &  x125 &  x149 &  x155 &  x161 &  x164 &  x179 &  x182 &  x185 &  x188 &  x200 &  x206 &  x209 &  x226 &  x233 &  x239 &  x242 &  x245 &  x248 &  x254 &  x260 &  x263 &  x269 &  x287 &  x296 &  x305 &  x310 &  x311 &  x317 &  x326 &  x329 &  x331 &  x332 &  x335 &  x338 &  x344 &  x349 &  x353 &  x356 &  x359 &  x368 &  x371 &  x377 &  x380 &  x392 &  x398 &  x404 &  x413 &  x416 &  x422 &  x428 &  x434 &  x440 &  x441 &  x455 &  x461 &  x473 &  x476 &  x481 &  x511 &  x512 &  x520 &  x524 &  x530 &  x533 &  x542 &  x551 &  x554 &  x560 &  x563 &  x566 &  x572 &  x590 &  x596 &  x602 &  x608 &  x623 &  x625 &  x626 &  x629 &  x635 &  x638 &  x641 &  x644 &  x656 &  x664 &  x668 &  x671 &  x674 &  x686 &  x689 &  x692 &  x701 &  x703 &  x704 &  x706 &  x707 &  x710 &  x713 &  x725 &  x737 &  x740 &  x761 &  x770 &  x776 &  x779 &  x791 &  x797 &  x803 &  x815 &  x818 &  x823 &  x827 &  x842 &  x851 &  x860 &  x862 &  x866 &  x872 &  x884 &  x887 &  x902 &  x905 &  x914 &  x920 &  x923 &  x935 &  x947 &  x950 &  x956 &  x962 &  x965 &  x971 &  x977 &  x980 &  x983 &  x992 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1028 &  x1031 &  x1040 &  x1049 &  x1052 &  x1055 &  x1058 &  x1076 &  x1088 &  x1097 &  x1103 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 & ~x237 & ~x276;
assign c3266 =  x2 &  x5 &  x8 &  x11 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x44 &  x50 &  x53 &  x56 &  x62 &  x65 &  x68 &  x71 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x257 &  x259 &  x260 &  x263 &  x266 &  x269 &  x275 &  x284 &  x293 &  x298 &  x299 &  x302 &  x305 &  x308 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x364 &  x365 &  x368 &  x371 &  x374 &  x380 &  x386 &  x389 &  x392 &  x394 &  x395 &  x403 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x431 &  x433 &  x434 &  x437 &  x440 &  x443 &  x448 &  x452 &  x455 &  x458 &  x464 &  x467 &  x470 &  x472 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x508 &  x509 &  x511 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x547 &  x548 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x589 &  x590 &  x596 &  x599 &  x602 &  x605 &  x611 &  x614 &  x617 &  x620 &  x623 &  x625 &  x626 &  x628 &  x629 &  x632 &  x638 &  x644 &  x650 &  x653 &  x656 &  x659 &  x662 &  x667 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x722 &  x725 &  x728 &  x734 &  x737 &  x740 &  x743 &  x745 &  x746 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x812 &  x823 &  x824 &  x827 &  x830 &  x836 &  x839 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x878 &  x881 &  x884 &  x893 &  x899 &  x902 &  x905 &  x911 &  x914 &  x920 &  x923 &  x926 &  x929 &  x935 &  x938 &  x941 &  x944 &  x950 &  x959 &  x962 &  x968 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x1001 &  x1004 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x513 & ~x552 & ~x639 & ~x678;
assign c3268 =  x2 &  x5 &  x8 &  x11 &  x17 &  x26 &  x29 &  x32 &  x35 &  x53 &  x56 &  x62 &  x68 &  x80 &  x83 &  x86 &  x89 &  x92 &  x98 &  x104 &  x107 &  x110 &  x125 &  x128 &  x131 &  x149 &  x152 &  x155 &  x161 &  x164 &  x170 &  x179 &  x194 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x233 &  x239 &  x242 &  x248 &  x251 &  x254 &  x272 &  x275 &  x278 &  x281 &  x287 &  x305 &  x323 &  x329 &  x332 &  x341 &  x344 &  x347 &  x350 &  x353 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x404 &  x407 &  x410 &  x413 &  x422 &  x425 &  x428 &  x434 &  x446 &  x449 &  x455 &  x458 &  x467 &  x470 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x503 &  x506 &  x515 &  x521 &  x524 &  x527 &  x530 &  x533 &  x542 &  x548 &  x556 &  x557 &  x560 &  x566 &  x569 &  x581 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x617 &  x620 &  x629 &  x632 &  x635 &  x638 &  x641 &  x653 &  x656 &  x665 &  x677 &  x680 &  x683 &  x686 &  x695 &  x701 &  x710 &  x716 &  x719 &  x722 &  x725 &  x731 &  x734 &  x737 &  x740 &  x743 &  x749 &  x752 &  x764 &  x767 &  x770 &  x773 &  x779 &  x788 &  x797 &  x803 &  x806 &  x815 &  x824 &  x833 &  x842 &  x854 &  x857 &  x862 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x890 &  x899 &  x901 &  x905 &  x914 &  x920 &  x923 &  x926 &  x938 &  x941 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x986 &  x995 &  x1013 &  x1016 &  x1018 &  x1025 &  x1028 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1057 &  x1061 &  x1076 &  x1085 &  x1088 &  x1091 &  x1096 &  x1100 &  x1106 &  x1112 &  x1118 &  x1121 &  x1124 &  x1130 & ~x417 & ~x495 & ~x612 & ~x717 & ~x795 & ~x810 & ~x894;
assign c3270 =  x1 &  x2 &  x8 &  x11 &  x17 &  x20 &  x23 &  x32 &  x40 &  x41 &  x47 &  x50 &  x53 &  x56 &  x59 &  x61 &  x62 &  x65 &  x68 &  x74 &  x77 &  x86 &  x92 &  x95 &  x98 &  x100 &  x101 &  x107 &  x110 &  x131 &  x137 &  x138 &  x140 &  x143 &  x149 &  x158 &  x161 &  x167 &  x170 &  x173 &  x178 &  x179 &  x182 &  x185 &  x191 &  x194 &  x203 &  x206 &  x209 &  x215 &  x217 &  x218 &  x224 &  x230 &  x236 &  x242 &  x248 &  x251 &  x254 &  x260 &  x263 &  x266 &  x275 &  x278 &  x283 &  x284 &  x287 &  x299 &  x311 &  x313 &  x320 &  x326 &  x329 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x359 &  x362 &  x371 &  x383 &  x386 &  x389 &  x392 &  x401 &  x410 &  x413 &  x422 &  x431 &  x446 &  x458 &  x464 &  x470 &  x476 &  x479 &  x485 &  x488 &  x490 &  x491 &  x503 &  x509 &  x515 &  x518 &  x521 &  x524 &  x527 &  x529 &  x533 &  x536 &  x539 &  x542 &  x548 &  x557 &  x560 &  x563 &  x569 &  x572 &  x581 &  x584 &  x593 &  x602 &  x605 &  x607 &  x608 &  x620 &  x623 &  x626 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x665 &  x668 &  x671 &  x676 &  x677 &  x683 &  x692 &  x695 &  x698 &  x701 &  x715 &  x719 &  x728 &  x737 &  x740 &  x749 &  x761 &  x776 &  x779 &  x782 &  x785 &  x793 &  x803 &  x806 &  x815 &  x818 &  x827 &  x830 &  x839 &  x848 &  x854 &  x869 &  x881 &  x890 &  x893 &  x908 &  x911 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x941 &  x944 &  x950 &  x953 &  x965 &  x971 &  x974 &  x977 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1046 &  x1049 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1079 &  x1088 &  x1094 &  x1106 &  x1109 &  x1112 &  x1118 &  x1124 &  x1127 & ~x381;
assign c3272 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x209 &  x212 &  x214 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x239 &  x242 &  x245 &  x248 &  x251 &  x253 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x286 &  x287 &  x290 &  x292 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x325 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x364 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x403 &  x404 &  x407 &  x409 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x442 &  x443 &  x445 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x481 &  x482 &  x484 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x556 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x589 &  x590 &  x593 &  x595 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x628 &  x629 &  x632 &  x634 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x667 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x703 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x742 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x781 &  x782 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x820 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x859 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x898 &  x899 &  x901 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x937 &  x938 &  x940 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1018 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1057 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130;
assign c3274 =  x1 &  x2 &  x5 &  x8 &  x17 &  x20 &  x23 &  x29 &  x41 &  x47 &  x50 &  x53 &  x59 &  x62 &  x65 &  x71 &  x79 &  x80 &  x95 &  x101 &  x104 &  x110 &  x113 &  x116 &  x118 &  x122 &  x128 &  x134 &  x143 &  x152 &  x155 &  x157 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x191 &  x194 &  x196 &  x197 &  x200 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x235 &  x236 &  x239 &  x242 &  x245 &  x248 &  x260 &  x269 &  x272 &  x275 &  x278 &  x284 &  x287 &  x290 &  x296 &  x302 &  x305 &  x314 &  x320 &  x323 &  x329 &  x332 &  x335 &  x341 &  x347 &  x356 &  x359 &  x362 &  x368 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x398 &  x401 &  x404 &  x407 &  x410 &  x422 &  x425 &  x428 &  x434 &  x440 &  x443 &  x452 &  x458 &  x461 &  x464 &  x467 &  x470 &  x479 &  x482 &  x485 &  x488 &  x491 &  x500 &  x506 &  x515 &  x524 &  x530 &  x539 &  x541 &  x545 &  x551 &  x563 &  x572 &  x578 &  x587 &  x593 &  x596 &  x605 &  x614 &  x620 &  x623 &  x629 &  x632 &  x635 &  x641 &  x644 &  x647 &  x662 &  x665 &  x668 &  x671 &  x674 &  x680 &  x683 &  x692 &  x695 &  x710 &  x713 &  x731 &  x734 &  x737 &  x743 &  x746 &  x752 &  x758 &  x767 &  x776 &  x779 &  x797 &  x803 &  x806 &  x809 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x844 &  x845 &  x848 &  x851 &  x854 &  x860 &  x863 &  x866 &  x869 &  x875 &  x878 &  x881 &  x887 &  x902 &  x905 &  x908 &  x914 &  x917 &  x920 &  x923 &  x926 &  x935 &  x965 &  x968 &  x980 &  x983 &  x986 &  x989 &  x995 &  x1001 &  x1007 &  x1010 &  x1019 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1103 &  x1112 &  x1118 &  x1121 & ~x18 & ~x45 & ~x96 & ~x135 & ~x162 & ~x163 & ~x174 & ~x213 & ~x252;
assign c3276 =  x5 &  x8 &  x11 &  x17 &  x23 &  x26 &  x32 &  x41 &  x44 &  x50 &  x53 &  x59 &  x65 &  x71 &  x74 &  x80 &  x83 &  x86 &  x92 &  x101 &  x107 &  x110 &  x116 &  x119 &  x122 &  x125 &  x134 &  x137 &  x143 &  x146 &  x149 &  x152 &  x155 &  x161 &  x164 &  x167 &  x169 &  x170 &  x191 &  x200 &  x207 &  x208 &  x209 &  x218 &  x221 &  x227 &  x230 &  x236 &  x239 &  x248 &  x254 &  x257 &  x263 &  x272 &  x275 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x314 &  x329 &  x332 &  x335 &  x347 &  x356 &  x359 &  x362 &  x371 &  x380 &  x391 &  x392 &  x401 &  x404 &  x407 &  x419 &  x428 &  x430 &  x431 &  x434 &  x443 &  x452 &  x458 &  x464 &  x467 &  x469 &  x473 &  x494 &  x500 &  x503 &  x506 &  x518 &  x521 &  x524 &  x530 &  x533 &  x539 &  x542 &  x545 &  x550 &  x554 &  x569 &  x572 &  x587 &  x589 &  x590 &  x602 &  x605 &  x611 &  x614 &  x620 &  x623 &  x626 &  x628 &  x638 &  x644 &  x647 &  x650 &  x653 &  x656 &  x665 &  x667 &  x671 &  x674 &  x677 &  x680 &  x686 &  x692 &  x695 &  x704 &  x719 &  x722 &  x725 &  x728 &  x731 &  x740 &  x755 &  x758 &  x761 &  x770 &  x773 &  x782 &  x785 &  x787 &  x788 &  x797 &  x800 &  x809 &  x812 &  x821 &  x827 &  x830 &  x833 &  x839 &  x842 &  x848 &  x851 &  x854 &  x860 &  x869 &  x878 &  x884 &  x887 &  x904 &  x908 &  x911 &  x914 &  x923 &  x926 &  x929 &  x938 &  x943 &  x944 &  x947 &  x953 &  x956 &  x959 &  x965 &  x968 &  x980 &  x982 &  x983 &  x986 &  x992 &  x998 &  x1001 &  x1004 &  x1013 &  x1022 &  x1031 &  x1037 &  x1040 &  x1046 &  x1052 &  x1061 &  x1064 &  x1076 &  x1082 &  x1085 &  x1088 &  x1094 &  x1100 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x522 & ~x561 & ~x819 & ~x858 & ~x1053;
assign c3278 =  x14 &  x20 &  x23 &  x26 &  x35 &  x47 &  x50 &  x53 &  x59 &  x86 &  x92 &  x95 &  x101 &  x104 &  x116 &  x122 &  x134 &  x140 &  x149 &  x164 &  x170 &  x182 &  x185 &  x203 &  x206 &  x209 &  x212 &  x218 &  x221 &  x227 &  x230 &  x254 &  x269 &  x272 &  x275 &  x284 &  x287 &  x296 &  x299 &  x311 &  x320 &  x323 &  x326 &  x335 &  x341 &  x347 &  x353 &  x368 &  x374 &  x386 &  x404 &  x410 &  x413 &  x425 &  x428 &  x434 &  x449 &  x455 &  x464 &  x473 &  x476 &  x479 &  x494 &  x503 &  x518 &  x521 &  x527 &  x545 &  x554 &  x572 &  x575 &  x578 &  x581 &  x590 &  x596 &  x605 &  x608 &  x611 &  x614 &  x626 &  x629 &  x641 &  x647 &  x650 &  x659 &  x662 &  x665 &  x671 &  x674 &  x677 &  x680 &  x692 &  x695 &  x710 &  x719 &  x722 &  x734 &  x737 &  x740 &  x746 &  x752 &  x758 &  x764 &  x767 &  x770 &  x776 &  x782 &  x785 &  x806 &  x812 &  x818 &  x824 &  x827 &  x851 &  x857 &  x860 &  x872 &  x875 &  x881 &  x884 &  x911 &  x929 &  x935 &  x944 &  x947 &  x959 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1016 &  x1022 &  x1028 &  x1037 &  x1043 &  x1052 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1097 &  x1103 &  x1106 &  x1121 &  x1124 &  x1127 &  x1130 & ~x300 & ~x651 & ~x696 & ~x735 & ~x813 & ~x846 & ~x852 & ~x885 & ~x891 & ~x924 & ~x963 & ~x964 & ~x969 & ~x1002 & ~x1029 & ~x1068 & ~x1080 & ~x1108;
assign c3280 =  x2 &  x5 &  x11 &  x17 &  x23 &  x29 &  x32 &  x41 &  x44 &  x47 &  x50 &  x52 &  x53 &  x56 &  x59 &  x65 &  x68 &  x74 &  x77 &  x80 &  x98 &  x113 &  x121 &  x122 &  x125 &  x131 &  x137 &  x140 &  x152 &  x155 &  x158 &  x160 &  x161 &  x170 &  x176 &  x179 &  x182 &  x194 &  x197 &  x200 &  x212 &  x221 &  x230 &  x236 &  x242 &  x245 &  x248 &  x254 &  x257 &  x260 &  x269 &  x278 &  x281 &  x287 &  x305 &  x308 &  x313 &  x316 &  x317 &  x332 &  x335 &  x347 &  x352 &  x353 &  x354 &  x362 &  x383 &  x386 &  x392 &  x393 &  x394 &  x398 &  x401 &  x404 &  x407 &  x413 &  x422 &  x428 &  x433 &  x437 &  x440 &  x443 &  x449 &  x458 &  x464 &  x472 &  x476 &  x482 &  x494 &  x497 &  x503 &  x506 &  x509 &  x512 &  x515 &  x521 &  x527 &  x533 &  x536 &  x539 &  x551 &  x572 &  x578 &  x593 &  x596 &  x599 &  x602 &  x605 &  x611 &  x617 &  x623 &  x631 &  x635 &  x644 &  x647 &  x659 &  x662 &  x668 &  x671 &  x677 &  x683 &  x688 &  x689 &  x701 &  x704 &  x707 &  x709 &  x719 &  x725 &  x728 &  x737 &  x740 &  x746 &  x748 &  x749 &  x752 &  x764 &  x767 &  x773 &  x776 &  x779 &  x785 &  x787 &  x799 &  x803 &  x805 &  x806 &  x818 &  x821 &  x824 &  x830 &  x836 &  x839 &  x844 &  x845 &  x854 &  x860 &  x865 &  x866 &  x875 &  x881 &  x890 &  x896 &  x899 &  x908 &  x911 &  x929 &  x932 &  x938 &  x941 &  x944 &  x962 &  x968 &  x989 &  x992 &  x1004 &  x1007 &  x1010 &  x1025 &  x1028 &  x1043 &  x1049 &  x1058 &  x1061 &  x1067 &  x1076 &  x1082 &  x1088 &  x1091 &  x1100 &  x1103 &  x1109 &  x1112 &  x1118 &  x1127 &  x1130 & ~x663 & ~x702 & ~x780 & ~x897 & ~x936;
assign c3282 =  x2 &  x8 &  x11 &  x14 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x53 &  x59 &  x62 &  x65 &  x68 &  x74 &  x80 &  x86 &  x89 &  x92 &  x95 &  x98 &  x104 &  x110 &  x113 &  x122 &  x125 &  x137 &  x140 &  x143 &  x152 &  x158 &  x161 &  x164 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x203 &  x206 &  x215 &  x218 &  x224 &  x227 &  x230 &  x236 &  x245 &  x254 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x299 &  x305 &  x311 &  x317 &  x320 &  x323 &  x331 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x370 &  x374 &  x377 &  x380 &  x386 &  x389 &  x401 &  x404 &  x410 &  x413 &  x419 &  x425 &  x428 &  x431 &  x437 &  x440 &  x449 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x482 &  x485 &  x488 &  x491 &  x497 &  x506 &  x509 &  x511 &  x512 &  x515 &  x518 &  x527 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x563 &  x566 &  x572 &  x578 &  x587 &  x589 &  x593 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x628 &  x629 &  x632 &  x635 &  x641 &  x644 &  x647 &  x659 &  x662 &  x664 &  x665 &  x667 &  x668 &  x674 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x706 &  x707 &  x710 &  x716 &  x719 &  x722 &  x725 &  x734 &  x740 &  x742 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x781 &  x782 &  x785 &  x791 &  x794 &  x797 &  x800 &  x806 &  x809 &  x812 &  x815 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x842 &  x845 &  x848 &  x860 &  x862 &  x869 &  x872 &  x875 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x935 &  x938 &  x940 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1018 &  x1019 &  x1022 &  x1025 &  x1034 &  x1037 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x195 & ~x234 & ~x756 & ~x834 & ~x835 & ~x873 & ~x874 & ~x912 & ~x951 & ~x990;
assign c3284 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x242 &  x245 &  x251 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x451 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x481 &  x482 &  x485 &  x488 &  x490 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x519 &  x520 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x548 &  x551 &  x554 &  x556 &  x557 &  x559 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x589 &  x590 &  x593 &  x595 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x628 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x667 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x742 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x781 &  x782 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x820 &  x821 &  x823 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x859 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x898 &  x899 &  x901 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x937 &  x938 &  x940 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x976 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1091 &  x1094 &  x1096 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x429;
assign c3286 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x116 &  x119 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x146 &  x149 &  x152 &  x155 &  x158 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x191 &  x197 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x223 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x248 &  x254 &  x257 &  x262 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x356 &  x365 &  x371 &  x374 &  x377 &  x380 &  x383 &  x389 &  x392 &  x395 &  x398 &  x404 &  x407 &  x409 &  x410 &  x413 &  x416 &  x418 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x526 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x556 &  x557 &  x560 &  x566 &  x569 &  x578 &  x581 &  x584 &  x587 &  x590 &  x594 &  x595 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x703 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x742 &  x743 &  x746 &  x749 &  x752 &  x755 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x820 &  x821 &  x823 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x907 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x938 &  x940 &  x947 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x977 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1018 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130;
assign c3288 =  x2 &  x5 &  x8 &  x10 &  x14 &  x20 &  x32 &  x38 &  x41 &  x47 &  x49 &  x50 &  x53 &  x56 &  x65 &  x68 &  x71 &  x74 &  x88 &  x92 &  x95 &  x98 &  x107 &  x113 &  x116 &  x125 &  x128 &  x131 &  x137 &  x140 &  x143 &  x146 &  x155 &  x158 &  x164 &  x175 &  x179 &  x182 &  x185 &  x191 &  x197 &  x203 &  x209 &  x214 &  x215 &  x221 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x253 &  x257 &  x260 &  x263 &  x266 &  x272 &  x275 &  x287 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x322 &  x323 &  x326 &  x332 &  x335 &  x338 &  x350 &  x353 &  x359 &  x362 &  x368 &  x371 &  x377 &  x380 &  x383 &  x389 &  x404 &  x407 &  x425 &  x431 &  x434 &  x440 &  x446 &  x449 &  x452 &  x455 &  x461 &  x464 &  x470 &  x473 &  x476 &  x479 &  x485 &  x491 &  x494 &  x497 &  x500 &  x515 &  x524 &  x526 &  x527 &  x530 &  x533 &  x542 &  x545 &  x548 &  x551 &  x557 &  x563 &  x566 &  x578 &  x581 &  x590 &  x596 &  x599 &  x602 &  x605 &  x614 &  x617 &  x629 &  x650 &  x659 &  x665 &  x668 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x713 &  x716 &  x722 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x749 &  x752 &  x758 &  x761 &  x773 &  x776 &  x779 &  x785 &  x794 &  x800 &  x805 &  x806 &  x824 &  x830 &  x836 &  x842 &  x844 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x869 &  x875 &  x881 &  x883 &  x884 &  x886 &  x887 &  x890 &  x893 &  x899 &  x902 &  x905 &  x908 &  x911 &  x926 &  x929 &  x932 &  x935 &  x944 &  x947 &  x950 &  x959 &  x965 &  x968 &  x980 &  x989 &  x992 &  x995 &  x998 &  x1000 &  x1003 &  x1004 &  x1007 &  x1010 &  x1013 &  x1019 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1055 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1078 &  x1079 &  x1081 &  x1082 &  x1085 &  x1091 &  x1103 &  x1106 &  x1112 &  x1118 &  x1121 &  x1127;
assign c3290 =  x29 &  x32 &  x41 &  x44 &  x59 &  x65 &  x77 &  x83 &  x89 &  x92 &  x95 &  x119 &  x137 &  x167 &  x179 &  x185 &  x188 &  x209 &  x215 &  x218 &  x224 &  x227 &  x233 &  x248 &  x254 &  x260 &  x269 &  x272 &  x278 &  x281 &  x290 &  x296 &  x305 &  x314 &  x322 &  x332 &  x347 &  x353 &  x365 &  x386 &  x398 &  x407 &  x413 &  x419 &  x428 &  x482 &  x485 &  x488 &  x491 &  x494 &  x503 &  x509 &  x518 &  x521 &  x527 &  x536 &  x539 &  x542 &  x548 &  x550 &  x590 &  x599 &  x608 &  x628 &  x632 &  x638 &  x641 &  x647 &  x656 &  x662 &  x665 &  x674 &  x701 &  x710 &  x716 &  x719 &  x743 &  x746 &  x752 &  x770 &  x779 &  x782 &  x791 &  x803 &  x821 &  x830 &  x836 &  x860 &  x881 &  x884 &  x902 &  x905 &  x920 &  x935 &  x941 &  x950 &  x995 &  x1007 &  x1037 &  x1043 &  x1052 &  x1058 &  x1061 &  x1064 &  x1070 &  x1079 &  x1127 & ~x228 & ~x375 & ~x376 & ~x561 & ~x639 & ~x717 & ~x780 & ~x858;
assign c3292 =  x20 &  x23 &  x26 &  x32 &  x38 &  x41 &  x44 &  x62 &  x68 &  x71 &  x89 &  x92 &  x98 &  x101 &  x104 &  x107 &  x110 &  x116 &  x122 &  x128 &  x131 &  x137 &  x143 &  x146 &  x149 &  x152 &  x164 &  x167 &  x170 &  x179 &  x182 &  x185 &  x191 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x251 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x277 &  x278 &  x281 &  x284 &  x293 &  x296 &  x305 &  x320 &  x323 &  x329 &  x332 &  x335 &  x341 &  x362 &  x365 &  x368 &  x371 &  x377 &  x386 &  x389 &  x392 &  x398 &  x404 &  x410 &  x413 &  x431 &  x437 &  x440 &  x443 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x470 &  x473 &  x476 &  x488 &  x491 &  x494 &  x497 &  x512 &  x515 &  x524 &  x527 &  x530 &  x536 &  x542 &  x554 &  x556 &  x560 &  x563 &  x566 &  x569 &  x575 &  x584 &  x590 &  x593 &  x602 &  x608 &  x611 &  x617 &  x620 &  x623 &  x626 &  x632 &  x635 &  x638 &  x641 &  x647 &  x659 &  x665 &  x671 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x704 &  x707 &  x710 &  x713 &  x734 &  x737 &  x740 &  x752 &  x761 &  x764 &  x770 &  x782 &  x785 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x812 &  x815 &  x824 &  x833 &  x839 &  x842 &  x845 &  x851 &  x854 &  x857 &  x863 &  x872 &  x878 &  x881 &  x884 &  x890 &  x896 &  x899 &  x905 &  x908 &  x911 &  x914 &  x920 &  x923 &  x926 &  x932 &  x935 &  x941 &  x944 &  x947 &  x953 &  x956 &  x962 &  x971 &  x974 &  x977 &  x983 &  x992 &  x995 &  x998 &  x1007 &  x1010 &  x1013 &  x1025 &  x1028 &  x1034 &  x1037 &  x1043 &  x1046 &  x1052 &  x1055 &  x1064 &  x1076 &  x1079 &  x1082 &  x1091 &  x1097 &  x1100 &  x1109 &  x1112 &  x1115 &  x1118 &  x1130 & ~x27 & ~x297 & ~x336 & ~x337 & ~x375 & ~x1026;
assign c3294 =  x2 &  x5 &  x8 &  x10 &  x11 &  x14 &  x17 &  x23 &  x26 &  x35 &  x41 &  x43 &  x44 &  x47 &  x50 &  x53 &  x56 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x89 &  x95 &  x98 &  x101 &  x104 &  x107 &  x113 &  x116 &  x117 &  x118 &  x121 &  x122 &  x125 &  x128 &  x131 &  x143 &  x149 &  x152 &  x157 &  x158 &  x160 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x194 &  x197 &  x199 &  x203 &  x206 &  x209 &  x218 &  x221 &  x230 &  x233 &  x238 &  x239 &  x242 &  x245 &  x248 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x274 &  x275 &  x277 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x308 &  x311 &  x313 &  x316 &  x323 &  x326 &  x335 &  x338 &  x341 &  x344 &  x353 &  x359 &  x362 &  x365 &  x368 &  x371 &  x377 &  x383 &  x392 &  x394 &  x398 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x433 &  x437 &  x440 &  x443 &  x452 &  x455 &  x458 &  x461 &  x467 &  x479 &  x482 &  x485 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x524 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x556 &  x557 &  x560 &  x563 &  x569 &  x571 &  x572 &  x575 &  x578 &  x581 &  x587 &  x590 &  x592 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x610 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x631 &  x632 &  x635 &  x641 &  x649 &  x650 &  x653 &  x656 &  x662 &  x665 &  x668 &  x671 &  x680 &  x683 &  x686 &  x688 &  x692 &  x695 &  x698 &  x707 &  x713 &  x716 &  x719 &  x722 &  x727 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x754 &  x761 &  x764 &  x766 &  x770 &  x773 &  x776 &  x779 &  x785 &  x788 &  x794 &  x797 &  x800 &  x803 &  x805 &  x806 &  x809 &  x815 &  x818 &  x821 &  x830 &  x836 &  x842 &  x844 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x866 &  x869 &  x875 &  x878 &  x881 &  x883 &  x884 &  x887 &  x893 &  x896 &  x899 &  x905 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x959 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x705 & ~x744 & ~x783;
assign c3296 =  x5 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x41 &  x44 &  x47 &  x50 &  x59 &  x65 &  x68 &  x71 &  x74 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x137 &  x140 &  x143 &  x146 &  x152 &  x158 &  x161 &  x167 &  x173 &  x176 &  x179 &  x182 &  x191 &  x194 &  x203 &  x206 &  x209 &  x215 &  x221 &  x224 &  x230 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x293 &  x296 &  x299 &  x305 &  x308 &  x311 &  x314 &  x320 &  x326 &  x329 &  x332 &  x338 &  x341 &  x344 &  x350 &  x362 &  x364 &  x368 &  x371 &  x374 &  x380 &  x383 &  x386 &  x389 &  x392 &  x394 &  x395 &  x401 &  x403 &  x404 &  x407 &  x410 &  x416 &  x419 &  x425 &  x434 &  x440 &  x443 &  x446 &  x452 &  x461 &  x467 &  x476 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x506 &  x509 &  x511 &  x512 &  x515 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x548 &  x550 &  x551 &  x554 &  x557 &  x560 &  x563 &  x569 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x596 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x628 &  x632 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x665 &  x667 &  x668 &  x671 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x704 &  x706 &  x707 &  x710 &  x713 &  x719 &  x722 &  x728 &  x731 &  x734 &  x737 &  x743 &  x745 &  x746 &  x749 &  x752 &  x761 &  x764 &  x767 &  x770 &  x779 &  x782 &  x784 &  x791 &  x797 &  x800 &  x803 &  x815 &  x821 &  x823 &  x824 &  x827 &  x833 &  x836 &  x839 &  x845 &  x854 &  x857 &  x860 &  x862 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x901 &  x905 &  x908 &  x914 &  x917 &  x923 &  x929 &  x938 &  x941 &  x947 &  x950 &  x953 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x977 &  x983 &  x986 &  x989 &  x992 &  x1001 &  x1004 &  x1010 &  x1013 &  x1019 &  x1025 &  x1028 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x39 & ~x156 & ~x195 & ~x273 & ~x879 & ~x885 & ~x918 & ~x957 & ~x1092;
assign c3298 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x80 &  x83 &  x86 &  x89 &  x91 &  x95 &  x101 &  x107 &  x110 &  x113 &  x116 &  x122 &  x128 &  x131 &  x134 &  x137 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x167 &  x168 &  x169 &  x170 &  x173 &  x176 &  x182 &  x185 &  x188 &  x191 &  x197 &  x200 &  x203 &  x205 &  x206 &  x208 &  x209 &  x212 &  x215 &  x218 &  x221 &  x227 &  x230 &  x233 &  x236 &  x238 &  x239 &  x245 &  x248 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x277 &  x278 &  x281 &  x284 &  x290 &  x293 &  x296 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x329 &  x332 &  x335 &  x338 &  x344 &  x347 &  x350 &  x353 &  x355 &  x356 &  x362 &  x365 &  x368 &  x371 &  x377 &  x383 &  x386 &  x389 &  x391 &  x392 &  x394 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x433 &  x434 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x550 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x587 &  x589 &  x590 &  x596 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x734 &  x737 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x788 &  x791 &  x794 &  x797 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x896 &  x899 &  x902 &  x905 &  x908 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x117 & ~x405 & ~x444 & ~x483 & ~x522 & ~x741 & ~x780 & ~x819 & ~x858 & ~x897;
assign c31 =  x936 &  x991 &  x1068 & ~x1011;
assign c33 =  x70 &  x286 &  x475 &  x493 &  x553 & ~x675 & ~x792;
assign c35 =  x274 &  x993 & ~x207 & ~x435;
assign c37 =  x640 &  x991 &  x1062 &  x1092;
assign c39 =  x23 &  x44 &  x47 &  x83 &  x125 &  x128 &  x131 &  x137 &  x152 &  x176 &  x206 &  x212 &  x215 &  x241 &  x254 &  x269 &  x308 &  x344 &  x356 &  x374 &  x392 &  x410 &  x428 &  x449 &  x461 &  x469 &  x470 &  x500 &  x518 &  x566 &  x569 &  x605 &  x638 &  x656 &  x671 &  x683 &  x692 &  x722 &  x758 &  x785 &  x791 &  x803 &  x869 &  x893 &  x896 &  x917 &  x929 &  x950 &  x968 &  x995 &  x1004 &  x1019 &  x1043 &  x1049 &  x1061 &  x1067 &  x1073 &  x1079 &  x1094 &  x1097 &  x1121 & ~x324 & ~x363 & ~x489;
assign c311 =  x664 &  x834 &  x1068 & ~x732;
assign c313 =  x76 &  x127 &  x279 &  x357 & ~x681;
assign c315 =  x170 &  x470 &  x742 &  x838 &  x991 & ~x438;
assign c317 =  x912 & ~x844;
assign c319 =  x253 &  x410 &  x664 &  x863 &  x1088 & ~x276 & ~x942 & ~x943;
assign c321 =  x35 &  x521 &  x736 &  x763 &  x1128 & ~x51;
assign c323 =  x142 &  x152 &  x242 &  x279 &  x473 &  x488 &  x653 &  x689 &  x851 & ~x288 & ~x780;
assign c325 = ~x651 & ~x901;
assign c327 =  x482 &  x577 &  x857 &  x871 & ~x99 & ~x187 & ~x258;
assign c329 =  x11 &  x14 &  x17 &  x83 &  x104 &  x140 &  x182 &  x188 &  x224 &  x227 &  x290 &  x296 &  x320 &  x341 &  x347 &  x359 &  x374 &  x422 &  x434 &  x461 &  x467 &  x482 &  x518 &  x521 &  x524 &  x569 &  x581 &  x587 &  x611 &  x676 &  x686 &  x689 &  x713 &  x737 &  x758 &  x761 &  x770 &  x779 &  x782 &  x812 &  x842 &  x878 &  x890 &  x926 &  x986 &  x989 &  x1037 &  x1046 &  x1064 &  x1100 & ~x513 & ~x568 & ~x591;
assign c331 =  x71 &  x85 &  x161 &  x697 & ~x589;
assign c333 =  x397 &  x586 &  x666 & ~x402 & ~x480;
assign c335 =  x1117 & ~x48 & ~x364 & ~x441;
assign c337 =  x71 &  x169 &  x695 &  x819 &  x1092;
assign c339 =  x31 &  x70 &  x95 &  x128 &  x161 &  x197 &  x248 &  x370 &  x380 &  x449 &  x593 &  x614 &  x626 &  x674 &  x701 &  x703 &  x704 &  x731 &  x869 &  x950 &  x1076 & ~x756 & ~x786 & ~x942 & ~x954;
assign c341 =  x561 & ~x492 & ~x576;
assign c343 =  x10 &  x160 &  x445 &  x561 & ~x414;
assign c345 =  x1061 &  x1117 & ~x165 & ~x333 & ~x396 & ~x744;
assign c347 =  x38 &  x62 &  x74 &  x83 &  x101 &  x128 &  x287 &  x317 &  x323 &  x341 &  x350 &  x352 &  x362 &  x407 &  x410 &  x452 &  x521 &  x683 &  x710 &  x719 &  x743 &  x752 &  x764 &  x767 &  x773 &  x815 &  x908 &  x959 &  x980 &  x992 &  x1049 &  x1121 & ~x3 & ~x207 & ~x264 & ~x327;
assign c349 =  x838 &  x871 &  x910 &  x986 & ~x12 & ~x51 & ~x52 & ~x819;
assign c351 = ~x1127;
assign c353 =  x1117 & ~x75 & ~x546 & ~x550;
assign c355 =  x154 &  x586 &  x667 &  x1061 & ~x243 & ~x480 & ~x816;
assign c357 =  x146 &  x317 &  x347 &  x461 &  x470 &  x656 & ~x42 & ~x207 & ~x285 & ~x441 & ~x858 & ~x912;
assign c359 =  x56 &  x116 &  x140 &  x163 &  x470 &  x947 & ~x282 & ~x480 & ~x978;
assign c361 =  x316 &  x975 &  x1068;
assign c363 =  x17 &  x41 &  x77 &  x122 &  x137 &  x152 &  x181 &  x265 &  x266 &  x293 &  x296 &  x368 &  x404 &  x467 &  x494 &  x503 &  x505 &  x560 &  x635 &  x698 &  x704 &  x707 &  x746 &  x755 &  x767 &  x770 &  x785 &  x815 &  x884 &  x887 &  x968 &  x1028 &  x1034 &  x1064 &  x1070 &  x1112 & ~x237 & ~x558 & ~x708;
assign c365 =  x17 &  x35 &  x53 &  x80 &  x89 &  x119 &  x149 &  x152 &  x206 &  x215 &  x248 &  x341 &  x350 &  x383 &  x407 &  x416 &  x428 &  x449 &  x557 &  x566 &  x599 &  x623 &  x635 &  x680 &  x695 &  x701 &  x704 &  x716 &  x784 &  x806 &  x862 &  x875 &  x878 &  x890 &  x893 &  x901 &  x902 &  x905 &  x940 &  x950 &  x953 &  x989 &  x1049 &  x1067 &  x1076 &  x1103 &  x1127 & ~x351 & ~x354 & ~x402 & ~x441 & ~x597 & ~x636 & ~x753;
assign c367 =  x234 &  x837 & ~x168;
assign c369 =  x169 &  x494 &  x553 &  x719 & ~x321 & ~x516 & ~x555 & ~x672 & ~x831 & ~x1059;
assign c371 = ~x302;
assign c373 = ~x541 & ~x669 & ~x690 & ~x708;
assign c375 =  x567 &  x639 & ~x595;
assign c377 =  x658 & ~x675 & ~x904;
assign c379 =  x279 & ~x394 & ~x600;
assign c381 =  x553 & ~x433 & ~x636 & ~x714;
assign c383 =  x82 &  x113 &  x328 &  x785 &  x926 &  x991 &  x1125 &  x1126 & ~x927;
assign c385 =  x20 &  x35 &  x53 &  x158 &  x160 &  x197 &  x266 &  x302 &  x371 &  x443 &  x679 &  x797 &  x890 &  x986 &  x1066 & ~x210 & ~x249 & ~x531;
assign c387 =  x622 &  x1033 & ~x474 & ~x790 & ~x1119;
assign c389 =  x700 & ~x243 & ~x1021 & ~x1059 & ~x1119;
assign c391 =  x76 &  x784 &  x792 & ~x450;
assign c393 = ~x12 & ~x706;
assign c395 =  x70 &  x76 &  x115 &  x158 &  x497 &  x524 &  x695 &  x761 &  x953 &  x971 & ~x939 & ~x960 & ~x978;
assign c397 =  x835 & ~x475 & ~x514;
assign c399 =  x123 &  x730 &  x922 & ~x249;
assign c3101 =  x600 &  x639 & ~x615;
assign c3103 =  x200 &  x503 & ~x48 & ~x306 & ~x363 & ~x474 & ~x498;
assign c3105 = ~x318 & ~x550 & ~x1101;
assign c3107 =  x987 & ~x99 & ~x292;
assign c3109 = ~x899;
assign c3111 =  x17 &  x35 &  x53 &  x59 &  x68 &  x74 &  x98 &  x101 &  x104 &  x155 &  x188 &  x260 &  x269 &  x272 &  x275 &  x281 &  x293 &  x341 &  x356 &  x359 &  x401 &  x404 &  x431 &  x452 &  x458 &  x479 &  x488 &  x497 &  x509 &  x527 &  x530 &  x542 &  x545 &  x569 &  x581 &  x587 &  x590 &  x599 &  x608 &  x617 &  x632 &  x635 &  x650 &  x662 &  x664 &  x689 &  x704 &  x713 &  x728 &  x737 &  x749 &  x752 &  x779 &  x791 &  x809 &  x824 &  x833 &  x845 &  x854 &  x890 &  x905 &  x911 &  x926 &  x944 &  x971 &  x983 &  x989 &  x1007 &  x1031 &  x1040 &  x1064 &  x1067 &  x1076 &  x1103 &  x1115 &  x1124 & ~x288 & ~x555 & ~x786 & ~x846 & ~x963;
assign c3113 =  x223 &  x316 &  x332 &  x743 &  x749 &  x869 &  x1082 & ~x138 & ~x210 & ~x744;
assign c3115 =  x147;
assign c3117 =  x322 &  x538 &  x993 & ~x12;
assign c3119 =  x553 &  x823 & ~x433 & ~x636;
assign c3121 =  x5 &  x89 &  x119 &  x163 &  x202 &  x241 &  x284 &  x290 &  x293 &  x596 &  x623 &  x647 &  x734 &  x743 &  x935 & ~x321 & ~x399 & ~x756 & ~x1020 & ~x1059;
assign c3123 =  x248 &  x335 &  x467 &  x649 &  x805 &  x869 &  x881 &  x883 &  x971 &  x1001 &  x1079 & ~x9 & ~x207 & ~x459;
assign c3125 =  x589 & ~x277 & ~x523;
assign c3127 = ~x355 & ~x454;
assign c3129 =  x277 & ~x357 & ~x396 & ~x589;
assign c3131 =  x535 &  x736 &  x998 &  x1089;
assign c3133 =  x547 &  x932 &  x1037 & ~x321 & ~x327 & ~x441;
assign c3135 =  x34 &  x397 & ~x399 & ~x453 & ~x531;
assign c3137 = ~x472 & ~x597 & ~x792 & ~x870;
assign c3139 =  x20 &  x92 &  x143 &  x203 &  x257 &  x260 &  x305 &  x320 &  x323 &  x391 &  x527 &  x629 &  x653 &  x689 &  x725 &  x758 &  x773 &  x797 &  x863 &  x929 &  x986 &  x1004 &  x1019 &  x1061 &  x1066 &  x1091 &  x1103 &  x1109 & ~x12 & ~x51 & ~x129 & ~x285 & ~x741 & ~x897 & ~x936;
assign c3141 = ~x394 & ~x519 & ~x675;
assign c3143 =  x398 &  x845 &  x1055 &  x1105 & ~x474 & ~x513 & ~x705 & ~x744 & ~x936 & ~x1014;
assign c3145 =  x31 &  x46 & ~x126;
assign c3147 =  x813 &  x1047 & ~x498 & ~x786;
assign c3149 =  x208 &  x1092 & ~x276 & ~x1099;
assign c3151 =  x35 &  x68 &  x159 &  x160 &  x200 &  x257 &  x299 &  x328 &  x338 &  x389 &  x445 &  x452 &  x476 &  x527 &  x551 &  x566 &  x581 &  x638 &  x641 &  x725 &  x926 &  x1037 &  x1043 & ~x471 & ~x510;
assign c3153 = ~x433 & ~x790;
assign c3155 =  x601 &  x1105 & ~x15 & ~x537 & ~x628;
assign c3157 = ~x3 & ~x168 & ~x369 & ~x741 & ~x1107 & ~x1119;
assign c3159 =  x82 &  x279 &  x1003 & ~x288;
assign c3161 =  x549 & ~x81 & ~x324 & ~x523;
assign c3163 =  x2 &  x11 &  x17 &  x74 &  x86 &  x92 &  x98 &  x110 &  x113 &  x119 &  x122 &  x137 &  x143 &  x149 &  x158 &  x173 &  x194 &  x197 &  x200 &  x206 &  x215 &  x218 &  x221 &  x230 &  x242 &  x247 &  x257 &  x272 &  x278 &  x299 &  x311 &  x320 &  x332 &  x335 &  x338 &  x341 &  x356 &  x362 &  x371 &  x377 &  x380 &  x398 &  x410 &  x416 &  x419 &  x425 &  x434 &  x437 &  x449 &  x461 &  x464 &  x470 &  x479 &  x482 &  x518 &  x536 &  x569 &  x617 &  x626 &  x677 &  x680 &  x683 &  x689 &  x703 &  x704 &  x710 &  x716 &  x719 &  x728 &  x731 &  x742 &  x746 &  x749 &  x758 &  x788 &  x797 &  x809 &  x812 &  x815 &  x827 &  x857 &  x872 &  x884 &  x905 &  x908 &  x911 &  x929 &  x932 &  x941 &  x944 &  x959 &  x977 &  x989 &  x992 &  x998 &  x1022 &  x1031 &  x1043 &  x1055 &  x1094 &  x1097 &  x1103 &  x1115 & ~x276 & ~x438 & ~x477 & ~x708 & ~x756 & ~x759;
assign c3165 = ~x631 & ~x901;
assign c3167 = ~x953;
assign c3169 =  x553 &  x1035 & ~x798;
assign c3171 =  x561 &  x678 & ~x978;
assign c3173 = ~x550 & ~x1101;
assign c3175 =  x990 &  x1062 & ~x882 & ~x960;
assign c3177 = ~x3 & ~x51 & ~x168 & ~x369 & ~x624 & ~x858;
assign c3179 =  x274 &  x688 &  x749 &  x799 &  x967 & ~x3 & ~x324;
assign c3181 =  x430 &  x510 & ~x120;
assign c3183 =  x988 &  x1104 & ~x594 & ~x864;
assign c3185 =  x83 &  x443 & ~x15 & ~x51 & ~x54 & ~x285 & ~x780 & ~x897 & ~x1068;
assign c3187 = ~x805 & ~x862;
assign c3189 =  x104 &  x142 &  x163 &  x226 &  x227 &  x232 &  x563 & ~x117 & ~x441 & ~x669;
assign c3191 =  x190 &  x697 &  x1117 & ~x204 & ~x244 & ~x879;
assign c3193 =  x43 &  x82 &  x91 &  x95 &  x154 &  x190 &  x215 &  x229 &  x730 &  x764 &  x839 &  x965 & ~x1011;
assign c3195 =  x512 &  x737 &  x953 &  x1000 &  x1018 &  x1039 & ~x324 & ~x363 & ~x474 & ~x591;
assign c3197 =  x263 &  x379 &  x452 &  x971 &  x1010 &  x1049 & ~x315 & ~x429 & ~x654 & ~x786;
assign c3199 =  x547 &  x586 &  x799 & ~x789;
assign c3201 =  x316 &  x387 &  x950 &  x1036;
assign c3203 =  x10 &  x73 &  x82 &  x98 &  x163 &  x187 &  x265 &  x649 &  x1118 & ~x312;
assign c3205 = ~x790;
assign c3207 = ~x1010;
assign c3209 =  x601 &  x637 & ~x475;
assign c3211 =  x783 & ~x394 & ~x558 & ~x615;
assign c3213 = ~x9 & ~x403;
assign c3215 =  x993 & ~x177 & ~x214 & ~x1014;
assign c3217 =  x128 &  x212 &  x292 &  x425 &  x466 &  x577 &  x911 & ~x595 & ~x672 & ~x750;
assign c3219 = ~x188;
assign c3221 =  x600 & ~x297 & ~x531 & ~x549;
assign c3223 =  x611 &  x819 &  x1092 & ~x195 & ~x753;
assign c3225 =  x52 &  x115 &  x179 &  x571 &  x814 &  x1036 & ~x276;
assign c3227 =  x466 &  x922 &  x1033 & ~x148 & ~x216;
assign c3229 =  x325 & ~x472 & ~x546 & ~x720;
assign c3231 =  x742 & ~x54 & ~x901;
assign c3233 =  x163 &  x281 &  x371 &  x391 &  x641 &  x668 &  x926 &  x929 &  x1127 & ~x171 & ~x207 & ~x285 & ~x324;
assign c3235 =  x1032;
assign c3237 =  x423 & ~x825;
assign c3239 =  x835 & ~x693 & ~x805;
assign c3241 =  x122 &  x131 &  x155 &  x161 &  x179 &  x182 &  x224 &  x233 &  x338 &  x368 &  x398 &  x425 &  x446 &  x485 &  x527 &  x563 &  x587 &  x638 &  x641 &  x659 &  x668 &  x679 &  x683 &  x764 &  x779 &  x791 &  x796 &  x866 &  x887 &  x959 &  x1019 &  x1051 &  x1076 &  x1079 &  x1091 & ~x168 & ~x357;
assign c3243 =  x27 &  x39 &  x837;
assign c3245 =  x53 &  x104 &  x146 &  x194 &  x245 &  x269 &  x272 &  x365 &  x458 &  x503 &  x512 &  x551 &  x560 &  x569 &  x605 &  x650 &  x668 &  x719 &  x730 &  x761 &  x803 &  x911 &  x917 &  x968 &  x1004 &  x1034 &  x1043 &  x1067 &  x1085 &  x1091 &  x1106 & ~x90 & ~x451;
assign c3247 = ~x979;
assign c3249 =  x823 &  x1027 & ~x138 & ~x331;
assign c3251 = ~x610 & ~x784;
assign c3253 =  x553 &  x638 &  x722 &  x823 & ~x288 & ~x556 & ~x672 & ~x750;
assign c3255 =  x439 &  x819 & ~x753;
assign c3257 =  x974 &  x1027 &  x1037 & ~x399 & ~x567 & ~x708;
assign c3259 =  x852 &  x991 &  x1053;
assign c3261 =  x169 &  x819 & ~x546;
assign c3263 =  x236 &  x667 &  x701 &  x998 &  x1069 &  x1102 & ~x276 & ~x636 & ~x786;
assign c3265 =  x365 &  x374 &  x545 &  x587 &  x761 &  x832 &  x917 &  x983 &  x1025 &  x1088 &  x1124 & ~x276 & ~x312 & ~x603 & ~x642 & ~x786;
assign c3267 = ~x355 & ~x645 & ~x679;
assign c3269 = ~x866;
assign c3271 =  x200 &  x449 &  x665 &  x806 &  x1026 &  x1033 &  x1088 &  x1090 & ~x447 & ~x846;
assign c3273 =  x70 &  x544 &  x814 & ~x754;
assign c3275 =  x356 &  x560 &  x593 &  x757 & ~x288 & ~x475;
assign c3277 =  x70 & ~x354 & ~x438 & ~x679;
assign c3279 =  x23 &  x29 &  x32 &  x41 &  x47 &  x71 &  x119 &  x128 &  x146 &  x167 &  x169 &  x203 &  x208 &  x227 &  x236 &  x242 &  x251 &  x257 &  x269 &  x275 &  x278 &  x280 &  x296 &  x302 &  x308 &  x314 &  x319 &  x329 &  x332 &  x356 &  x358 &  x368 &  x371 &  x389 &  x392 &  x398 &  x404 &  x416 &  x419 &  x422 &  x436 &  x437 &  x461 &  x464 &  x476 &  x482 &  x503 &  x518 &  x530 &  x554 &  x572 &  x575 &  x587 &  x626 &  x632 &  x641 &  x650 &  x659 &  x662 &  x695 &  x704 &  x745 &  x749 &  x761 &  x776 &  x779 &  x794 &  x800 &  x803 &  x812 &  x815 &  x830 &  x839 &  x851 &  x857 &  x878 &  x884 &  x896 &  x914 &  x923 &  x941 &  x953 &  x989 &  x992 &  x1001 &  x1010 &  x1019 &  x1022 &  x1031 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1112 &  x1127 & ~x198 & ~x480;
assign c3281 =  x70 &  x214 &  x346 &  x350 & ~x276 & ~x438 & ~x1119;
assign c3283 =  x187 &  x226 &  x379 &  x547 & ~x156;
assign c3285 =  x156 & ~x12 & ~x13 & ~x327;
assign c3287 =  x551 &  x700 &  x905 & ~x754 & ~x1065;
assign c3289 =  x83 &  x110 &  x137 &  x190 &  x224 &  x248 &  x268 &  x305 &  x329 &  x407 &  x449 &  x536 &  x587 &  x767 &  x874 &  x1009 &  x1048 & ~x9 & ~x288;
assign c3291 =  x10 &  x76 &  x521 &  x755 &  x872 & ~x546 & ~x678 & ~x684;
assign c3293 =  x76 &  x397 &  x550 & ~x486 & ~x564;
assign c3295 =  x273 & ~x3 & ~x168 & ~x265;
assign c3297 =  x340 &  x510 &  x835 & ~x489;
assign c3299 = ~x78 & ~x117 & ~x285 & ~x324 & ~x375 & ~x459 & ~x741 & ~x1014;
assign c40 =  x2 &  x11 &  x14 &  x17 &  x20 &  x26 &  x29 &  x50 &  x59 &  x65 &  x74 &  x77 &  x80 &  x83 &  x86 &  x98 &  x101 &  x113 &  x119 &  x122 &  x125 &  x131 &  x134 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x164 &  x167 &  x170 &  x182 &  x188 &  x191 &  x197 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x233 &  x236 &  x239 &  x245 &  x254 &  x257 &  x263 &  x269 &  x272 &  x275 &  x281 &  x290 &  x293 &  x302 &  x308 &  x314 &  x317 &  x320 &  x332 &  x335 &  x338 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x364 &  x365 &  x374 &  x380 &  x383 &  x386 &  x389 &  x392 &  x398 &  x404 &  x407 &  x410 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x446 &  x449 &  x452 &  x455 &  x458 &  x464 &  x467 &  x473 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x518 &  x524 &  x530 &  x536 &  x539 &  x548 &  x554 &  x560 &  x563 &  x572 &  x575 &  x587 &  x593 &  x599 &  x601 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x695 &  x698 &  x701 &  x707 &  x710 &  x722 &  x728 &  x737 &  x752 &  x755 &  x758 &  x761 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x800 &  x803 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x835 &  x836 &  x842 &  x845 &  x851 &  x857 &  x860 &  x863 &  x878 &  x890 &  x896 &  x902 &  x908 &  x910 &  x911 &  x917 &  x923 &  x932 &  x938 &  x944 &  x947 &  x950 &  x956 &  x959 &  x962 &  x968 &  x977 &  x980 &  x983 &  x986 &  x992 &  x998 &  x1001 &  x1004 &  x1010 &  x1025 &  x1027 &  x1031 &  x1034 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1076 &  x1085 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1118 &  x1124 &  x1130 & ~x12 & ~x51 & ~x432 & ~x465 & ~x750;
assign c42 =  x2 &  x5 &  x8 &  x14 &  x17 &  x23 &  x29 &  x35 &  x38 &  x41 &  x44 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x152 &  x155 &  x158 &  x161 &  x167 &  x170 &  x173 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x206 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x269 &  x272 &  x277 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x316 &  x317 &  x323 &  x329 &  x332 &  x335 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x355 &  x356 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x394 &  x395 &  x398 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x484 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x508 &  x512 &  x515 &  x518 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x596 &  x598 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x707 &  x710 &  x713 &  x716 &  x718 &  x719 &  x722 &  x725 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x851 &  x854 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1027 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1066 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x513 & ~x552 & ~x666 & ~x705 & ~x783 & ~x822;
assign c44 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x503 &  x506 &  x509 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x542 &  x545 &  x548 &  x550 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x625 &  x626 &  x632 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x704 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x790 &  x791 &  x793 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x829 &  x830 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x941 &  x944 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x669 & ~x670 & ~x708 & ~x786 & ~x939 & ~x978;
assign c46 =  x5 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x44 &  x50 &  x53 &  x62 &  x83 &  x86 &  x89 &  x95 &  x98 &  x110 &  x113 &  x116 &  x122 &  x128 &  x137 &  x143 &  x149 &  x155 &  x164 &  x167 &  x170 &  x179 &  x185 &  x188 &  x191 &  x197 &  x206 &  x218 &  x230 &  x233 &  x236 &  x239 &  x242 &  x248 &  x251 &  x266 &  x269 &  x278 &  x284 &  x296 &  x308 &  x323 &  x326 &  x329 &  x338 &  x353 &  x356 &  x359 &  x380 &  x398 &  x404 &  x407 &  x413 &  x419 &  x425 &  x428 &  x434 &  x437 &  x440 &  x449 &  x455 &  x470 &  x473 &  x476 &  x479 &  x491 &  x494 &  x506 &  x512 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x581 &  x587 &  x590 &  x599 &  x602 &  x605 &  x608 &  x617 &  x620 &  x623 &  x629 &  x635 &  x641 &  x644 &  x650 &  x656 &  x665 &  x668 &  x677 &  x680 &  x686 &  x698 &  x704 &  x710 &  x713 &  x722 &  x743 &  x749 &  x758 &  x770 &  x776 &  x781 &  x785 &  x788 &  x797 &  x800 &  x803 &  x809 &  x812 &  x818 &  x827 &  x833 &  x839 &  x845 &  x848 &  x851 &  x854 &  x859 &  x863 &  x866 &  x869 &  x872 &  x875 &  x884 &  x902 &  x917 &  x926 &  x932 &  x941 &  x947 &  x953 &  x959 &  x962 &  x965 &  x971 &  x977 &  x980 &  x983 &  x986 &  x991 &  x995 &  x1007 &  x1022 &  x1025 &  x1028 &  x1030 &  x1040 &  x1046 &  x1049 &  x1052 &  x1064 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1112 &  x1121 & ~x321 & ~x849 & ~x888 & ~x903 & ~x928 & ~x960 & ~x966 & ~x1005 & ~x1011 & ~x1050 & ~x1089;
assign c48 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x109 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x355 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x394 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x433 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x472 &  x473 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x508 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x547 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x601 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x679 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x718 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x757 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x796 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x835 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x874 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x513 & ~x552 & ~x591 & ~x744 & ~x783 & ~x822 & ~x861;
assign c410 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x194 &  x196 &  x197 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x235 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x344 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x476 &  x479 &  x482 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x548 &  x551 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x889 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x917 &  x920 &  x923 &  x926 &  x928 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x953 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x66 & ~x357 & ~x396 & ~x420 & ~x435 & ~x474 & ~x501 & ~x549 & ~x588 & ~x627 & ~x666 & ~x705;
assign c412 =  x2 &  x8 &  x11 &  x20 &  x23 &  x26 &  x32 &  x41 &  x44 &  x53 &  x59 &  x62 &  x65 &  x68 &  x77 &  x83 &  x86 &  x89 &  x98 &  x101 &  x107 &  x110 &  x113 &  x116 &  x122 &  x131 &  x134 &  x137 &  x143 &  x146 &  x149 &  x155 &  x158 &  x164 &  x173 &  x176 &  x179 &  x182 &  x185 &  x191 &  x194 &  x200 &  x203 &  x206 &  x212 &  x218 &  x220 &  x221 &  x236 &  x239 &  x245 &  x257 &  x260 &  x263 &  x266 &  x272 &  x275 &  x281 &  x284 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x326 &  x329 &  x335 &  x341 &  x347 &  x350 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x380 &  x383 &  x389 &  x395 &  x404 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x464 &  x467 &  x470 &  x482 &  x488 &  x491 &  x497 &  x512 &  x515 &  x521 &  x524 &  x527 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x566 &  x569 &  x572 &  x575 &  x578 &  x587 &  x599 &  x602 &  x605 &  x617 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x659 &  x665 &  x668 &  x671 &  x677 &  x680 &  x683 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x719 &  x725 &  x731 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x767 &  x773 &  x776 &  x779 &  x782 &  x788 &  x794 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x820 &  x821 &  x830 &  x833 &  x836 &  x839 &  x845 &  x848 &  x860 &  x874 &  x875 &  x884 &  x890 &  x893 &  x899 &  x911 &  x914 &  x917 &  x926 &  x929 &  x935 &  x938 &  x947 &  x953 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x989 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1022 &  x1031 &  x1040 &  x1043 &  x1046 &  x1052 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1091 &  x1097 &  x1103 &  x1106 &  x1112 &  x1114 &  x1118 &  x1124 &  x1127 & ~x360 & ~x582 & ~x855 & ~x1017;
assign c414 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x92 &  x95 &  x98 &  x104 &  x107 &  x110 &  x116 &  x119 &  x122 &  x125 &  x131 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x155 &  x158 &  x160 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x188 &  x191 &  x194 &  x197 &  x199 &  x200 &  x206 &  x209 &  x212 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x235 &  x236 &  x238 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x260 &  x266 &  x272 &  x274 &  x275 &  x277 &  x278 &  x281 &  x284 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x316 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x391 &  x392 &  x395 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x517 &  x518 &  x521 &  x527 &  x530 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x555 &  x556 &  x557 &  x560 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x598 &  x599 &  x602 &  x608 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x707 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x821 &  x824 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x956 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 & ~x396 & ~x435 & ~x474 & ~x513 & ~x666 & ~x744;
assign c416 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x50 &  x53 &  x56 &  x59 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x113 &  x119 &  x122 &  x128 &  x131 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x254 &  x257 &  x263 &  x269 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x314 &  x320 &  x323 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x356 &  x362 &  x365 &  x368 &  x377 &  x380 &  x383 &  x386 &  x395 &  x398 &  x404 &  x407 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x443 &  x446 &  x449 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x479 &  x482 &  x485 &  x488 &  x491 &  x497 &  x500 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x584 &  x587 &  x589 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x617 &  x623 &  x626 &  x628 &  x632 &  x635 &  x638 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x668 &  x671 &  x674 &  x677 &  x683 &  x686 &  x692 &  x695 &  x701 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x728 &  x734 &  x737 &  x740 &  x743 &  x749 &  x752 &  x758 &  x761 &  x764 &  x767 &  x770 &  x776 &  x779 &  x781 &  x782 &  x785 &  x788 &  x791 &  x794 &  x806 &  x812 &  x815 &  x820 &  x821 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x859 &  x863 &  x867 &  x868 &  x869 &  x871 &  x872 &  x875 &  x878 &  x884 &  x887 &  x893 &  x899 &  x908 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1013 &  x1016 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x747 & ~x786 & ~x825 & ~x894;
assign c418 =  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x95 &  x97 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x131 &  x134 &  x136 &  x137 &  x140 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x173 &  x175 &  x176 &  x179 &  x185 &  x188 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x214 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x278 &  x284 &  x287 &  x290 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x320 &  x323 &  x326 &  x329 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x394 &  x398 &  x401 &  x407 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x433 &  x434 &  x437 &  x440 &  x443 &  x446 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x500 &  x506 &  x509 &  x511 &  x512 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x542 &  x548 &  x550 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x614 &  x617 &  x620 &  x626 &  x629 &  x632 &  x635 &  x641 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x725 &  x731 &  x734 &  x740 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x797 &  x800 &  x806 &  x809 &  x812 &  x815 &  x821 &  x824 &  x830 &  x836 &  x839 &  x842 &  x848 &  x851 &  x857 &  x860 &  x863 &  x875 &  x881 &  x884 &  x887 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x971 &  x977 &  x980 &  x986 &  x989 &  x992 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1034 &  x1037 &  x1046 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1130 & ~x117 & ~x156 & ~x444 & ~x615 & ~x654 & ~x693 & ~x975 & ~x1014 & ~x1053 & ~x1092;
assign c420 =  x2 &  x5 &  x8 &  x14 &  x20 &  x26 &  x32 &  x35 &  x41 &  x47 &  x62 &  x65 &  x68 &  x71 &  x80 &  x89 &  x101 &  x104 &  x107 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x140 &  x146 &  x149 &  x152 &  x155 &  x167 &  x170 &  x176 &  x179 &  x182 &  x197 &  x203 &  x212 &  x215 &  x223 &  x230 &  x233 &  x236 &  x242 &  x245 &  x251 &  x254 &  x257 &  x262 &  x272 &  x278 &  x284 &  x287 &  x293 &  x299 &  x302 &  x305 &  x314 &  x317 &  x326 &  x329 &  x335 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x368 &  x374 &  x377 &  x386 &  x389 &  x392 &  x398 &  x404 &  x410 &  x419 &  x425 &  x434 &  x437 &  x443 &  x446 &  x455 &  x458 &  x464 &  x470 &  x473 &  x482 &  x488 &  x491 &  x506 &  x512 &  x515 &  x521 &  x524 &  x527 &  x530 &  x539 &  x542 &  x545 &  x554 &  x557 &  x566 &  x569 &  x578 &  x584 &  x590 &  x599 &  x602 &  x605 &  x611 &  x617 &  x620 &  x626 &  x629 &  x632 &  x640 &  x641 &  x644 &  x647 &  x650 &  x656 &  x659 &  x662 &  x671 &  x677 &  x707 &  x710 &  x716 &  x719 &  x722 &  x725 &  x731 &  x737 &  x749 &  x764 &  x767 &  x773 &  x776 &  x782 &  x785 &  x794 &  x797 &  x800 &  x803 &  x809 &  x812 &  x818 &  x820 &  x821 &  x824 &  x830 &  x833 &  x836 &  x845 &  x848 &  x866 &  x869 &  x872 &  x890 &  x893 &  x896 &  x898 &  x899 &  x908 &  x914 &  x917 &  x920 &  x926 &  x929 &  x932 &  x937 &  x941 &  x944 &  x947 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x986 &  x992 &  x995 &  x1001 &  x1004 &  x1010 &  x1013 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1076 &  x1079 &  x1085 &  x1091 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 & ~x699 & ~x747 & ~x816 & ~x855 & ~x894 & ~x966 & ~x1017 & ~x1056;
assign c422 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x101 &  x104 &  x107 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x335 &  x338 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x469 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x494 &  x497 &  x500 &  x503 &  x506 &  x508 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x542 &  x545 &  x547 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x698 &  x701 &  x704 &  x707 &  x710 &  x716 &  x722 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x438 & ~x513 & ~x528 & ~x552 & ~x591 & ~x592 & ~x630 & ~x705 & ~x744 & ~x783 & ~x822 & ~x861;
assign c424 =  x11 &  x17 &  x26 &  x38 &  x41 &  x53 &  x62 &  x68 &  x71 &  x73 &  x74 &  x80 &  x89 &  x95 &  x101 &  x107 &  x110 &  x113 &  x116 &  x122 &  x125 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x164 &  x167 &  x170 &  x182 &  x185 &  x188 &  x194 &  x209 &  x212 &  x221 &  x230 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x269 &  x275 &  x278 &  x281 &  x287 &  x293 &  x296 &  x299 &  x305 &  x311 &  x314 &  x323 &  x335 &  x344 &  x350 &  x356 &  x365 &  x374 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x422 &  x431 &  x434 &  x437 &  x446 &  x452 &  x455 &  x461 &  x464 &  x470 &  x472 &  x476 &  x479 &  x485 &  x491 &  x494 &  x500 &  x506 &  x508 &  x509 &  x512 &  x515 &  x524 &  x530 &  x533 &  x536 &  x542 &  x550 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x575 &  x578 &  x581 &  x584 &  x590 &  x593 &  x596 &  x599 &  x608 &  x611 &  x614 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x640 &  x644 &  x647 &  x656 &  x668 &  x671 &  x677 &  x679 &  x680 &  x686 &  x689 &  x704 &  x707 &  x710 &  x713 &  x718 &  x719 &  x728 &  x731 &  x734 &  x740 &  x749 &  x752 &  x755 &  x757 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x779 &  x785 &  x788 &  x791 &  x806 &  x812 &  x821 &  x824 &  x827 &  x833 &  x836 &  x839 &  x848 &  x854 &  x857 &  x863 &  x872 &  x875 &  x881 &  x884 &  x890 &  x896 &  x914 &  x923 &  x929 &  x932 &  x938 &  x950 &  x953 &  x956 &  x959 &  x962 &  x968 &  x983 &  x986 &  x989 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1034 &  x1055 &  x1058 &  x1061 &  x1067 &  x1070 &  x1082 &  x1088 &  x1097 &  x1100 &  x1103 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x537 & ~x660;
assign c426 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x107 &  x110 &  x113 &  x116 &  x119 &  x121 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x160 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x196 &  x198 &  x199 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x227 &  x230 &  x233 &  x235 &  x236 &  x238 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x274 &  x277 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x401 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x442 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x464 &  x467 &  x470 &  x476 &  x479 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x632 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x679 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x710 &  x713 &  x716 &  x718 &  x725 &  x731 &  x734 &  x737 &  x740 &  x746 &  x749 &  x752 &  x755 &  x757 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x796 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x854 &  x857 &  x860 &  x866 &  x869 &  x872 &  x878 &  x881 &  x884 &  x887 &  x889 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x910 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x977 &  x980 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x318 & ~x333 & ~x357 & ~x588 & ~x627 & ~x666 & ~x705 & ~x744 & ~x783 & ~x858 & ~x897;
assign c428 =  x11 &  x14 &  x20 &  x26 &  x29 &  x35 &  x38 &  x56 &  x65 &  x71 &  x74 &  x80 &  x83 &  x92 &  x101 &  x104 &  x116 &  x122 &  x125 &  x137 &  x140 &  x146 &  x152 &  x155 &  x158 &  x164 &  x167 &  x176 &  x182 &  x191 &  x197 &  x200 &  x209 &  x212 &  x215 &  x224 &  x233 &  x235 &  x236 &  x239 &  x245 &  x248 &  x260 &  x263 &  x269 &  x274 &  x275 &  x284 &  x293 &  x296 &  x302 &  x308 &  x311 &  x320 &  x326 &  x329 &  x338 &  x341 &  x350 &  x352 &  x353 &  x356 &  x368 &  x371 &  x380 &  x382 &  x386 &  x389 &  x391 &  x398 &  x401 &  x404 &  x410 &  x419 &  x425 &  x431 &  x434 &  x437 &  x443 &  x455 &  x458 &  x461 &  x470 &  x473 &  x476 &  x479 &  x485 &  x497 &  x500 &  x512 &  x515 &  x518 &  x530 &  x533 &  x536 &  x539 &  x554 &  x557 &  x560 &  x563 &  x569 &  x578 &  x581 &  x584 &  x593 &  x596 &  x602 &  x608 &  x611 &  x617 &  x620 &  x626 &  x635 &  x638 &  x644 &  x650 &  x653 &  x662 &  x668 &  x671 &  x674 &  x683 &  x695 &  x710 &  x716 &  x718 &  x719 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x757 &  x761 &  x767 &  x773 &  x776 &  x779 &  x785 &  x788 &  x791 &  x794 &  x796 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x827 &  x830 &  x835 &  x839 &  x842 &  x854 &  x859 &  x863 &  x872 &  x874 &  x875 &  x878 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x905 &  x910 &  x911 &  x913 &  x926 &  x935 &  x937 &  x938 &  x944 &  x947 &  x953 &  x956 &  x959 &  x965 &  x968 &  x977 &  x992 &  x1004 &  x1007 &  x1010 &  x1013 &  x1019 &  x1028 &  x1034 &  x1037 &  x1040 &  x1049 &  x1058 &  x1067 &  x1073 &  x1082 &  x1085 &  x1088 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x1017 & ~x1095;
assign c430 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x122 &  x125 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x206 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x266 &  x269 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x332 &  x338 &  x341 &  x344 &  x347 &  x353 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x482 &  x485 &  x488 &  x494 &  x497 &  x500 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x550 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x703 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x742 &  x743 &  x746 &  x749 &  x751 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x789 &  x790 &  x791 &  x797 &  x800 &  x803 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x829 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x869 &  x872 &  x875 &  x881 &  x884 &  x887 &  x890 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x708 & ~x783 & ~x939 & ~x978 & ~x1017;
assign c432 =  x2 &  x11 &  x14 &  x17 &  x38 &  x50 &  x62 &  x68 &  x71 &  x74 &  x77 &  x89 &  x92 &  x101 &  x113 &  x116 &  x119 &  x122 &  x137 &  x146 &  x155 &  x158 &  x164 &  x185 &  x200 &  x203 &  x212 &  x221 &  x227 &  x236 &  x239 &  x257 &  x260 &  x263 &  x269 &  x272 &  x278 &  x284 &  x290 &  x304 &  x308 &  x338 &  x343 &  x344 &  x347 &  x356 &  x362 &  x365 &  x374 &  x382 &  x392 &  x404 &  x407 &  x410 &  x419 &  x421 &  x422 &  x428 &  x431 &  x434 &  x437 &  x440 &  x452 &  x455 &  x473 &  x476 &  x479 &  x497 &  x500 &  x515 &  x521 &  x533 &  x542 &  x548 &  x557 &  x569 &  x575 &  x578 &  x590 &  x605 &  x623 &  x626 &  x635 &  x638 &  x641 &  x644 &  x659 &  x668 &  x680 &  x705 &  x707 &  x725 &  x728 &  x737 &  x745 &  x752 &  x758 &  x761 &  x781 &  x783 &  x788 &  x797 &  x809 &  x821 &  x823 &  x824 &  x839 &  x862 &  x872 &  x881 &  x884 &  x905 &  x914 &  x926 &  x929 &  x932 &  x944 &  x953 &  x962 &  x968 &  x971 &  x974 &  x977 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1010 &  x1016 &  x1019 &  x1022 &  x1031 &  x1037 &  x1043 &  x1046 &  x1052 &  x1064 &  x1085 &  x1091 &  x1094 &  x1100 &  x1106 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x351 & ~x429 & ~x507 & ~x546 & ~x624 & ~x750 & ~x903;
assign c434 =  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x161 &  x164 &  x170 &  x173 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x251 &  x254 &  x260 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x314 &  x320 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x356 &  x362 &  x365 &  x368 &  x371 &  x380 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x476 &  x479 &  x482 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x508 &  x512 &  x515 &  x518 &  x524 &  x527 &  x530 &  x536 &  x542 &  x545 &  x547 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x620 &  x623 &  x626 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x695 &  x701 &  x704 &  x707 &  x713 &  x716 &  x722 &  x725 &  x728 &  x731 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x791 &  x794 &  x803 &  x806 &  x809 &  x812 &  x815 &  x821 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x863 &  x869 &  x872 &  x878 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x923 &  x929 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1034 &  x1037 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130 & ~x51 & ~x90 & ~x96 & ~x129 & ~x174 & ~x477 & ~x504 & ~x582 & ~x687 & ~x822 & ~x825 & ~x864 & ~x900;
assign c436 =  x5 &  x14 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x62 &  x68 &  x74 &  x77 &  x80 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x116 &  x119 &  x122 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x164 &  x167 &  x170 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x224 &  x230 &  x233 &  x236 &  x245 &  x248 &  x251 &  x254 &  x260 &  x263 &  x266 &  x269 &  x278 &  x281 &  x287 &  x296 &  x302 &  x305 &  x308 &  x311 &  x314 &  x323 &  x326 &  x329 &  x332 &  x335 &  x341 &  x344 &  x350 &  x356 &  x359 &  x365 &  x371 &  x377 &  x380 &  x383 &  x392 &  x395 &  x398 &  x401 &  x404 &  x419 &  x425 &  x431 &  x434 &  x437 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x473 &  x476 &  x479 &  x482 &  x488 &  x491 &  x497 &  x509 &  x512 &  x515 &  x521 &  x524 &  x527 &  x530 &  x536 &  x542 &  x548 &  x551 &  x554 &  x557 &  x560 &  x569 &  x572 &  x584 &  x593 &  x596 &  x605 &  x608 &  x611 &  x623 &  x626 &  x627 &  x629 &  x644 &  x647 &  x650 &  x653 &  x656 &  x668 &  x671 &  x674 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x728 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x758 &  x761 &  x767 &  x770 &  x773 &  x779 &  x781 &  x782 &  x785 &  x794 &  x803 &  x809 &  x812 &  x830 &  x836 &  x839 &  x842 &  x848 &  x851 &  x854 &  x863 &  x866 &  x869 &  x878 &  x884 &  x890 &  x893 &  x899 &  x902 &  x911 &  x917 &  x920 &  x923 &  x926 &  x932 &  x938 &  x947 &  x950 &  x953 &  x962 &  x965 &  x971 &  x974 &  x980 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1040 &  x1046 &  x1052 &  x1055 &  x1061 &  x1064 &  x1070 &  x1076 &  x1079 &  x1085 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1127 &  x1130 & ~x273 & ~x312 & ~x351 & ~x390 & ~x801 & ~x840 & ~x841 & ~x879 & ~x888 & ~x903 & ~x918 & ~x966;
assign c438 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x241 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x278 &  x280 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x319 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x419 &  x425 &  x428 &  x431 &  x432 &  x433 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x464 &  x467 &  x470 &  x472 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x506 &  x508 &  x509 &  x511 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x542 &  x545 &  x547 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x590 &  x593 &  x596 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x761 &  x764 &  x767 &  x770 &  x773 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x935 &  x938 &  x941 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1019 &  x1022 &  x1025 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1127 &  x1130 & ~x78 & ~x156 & ~x195 & ~x234 & ~x306 & ~x345 & ~x438;
assign c440 =  x2 &  x4 &  x5 &  x6 &  x7 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x43 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x80 &  x86 &  x89 &  x95 &  x98 &  x101 &  x107 &  x110 &  x116 &  x119 &  x121 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x159 &  x160 &  x161 &  x170 &  x173 &  x179 &  x182 &  x185 &  x191 &  x194 &  x196 &  x197 &  x198 &  x199 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x227 &  x233 &  x235 &  x236 &  x239 &  x248 &  x254 &  x257 &  x263 &  x266 &  x269 &  x272 &  x274 &  x275 &  x277 &  x278 &  x281 &  x284 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x404 &  x410 &  x413 &  x419 &  x422 &  x425 &  x428 &  x431 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x617 &  x620 &  x623 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x677 &  x680 &  x689 &  x692 &  x695 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x758 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x824 &  x830 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x896 &  x902 &  x905 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x935 &  x938 &  x944 &  x950 &  x953 &  x959 &  x962 &  x968 &  x971 &  x974 &  x977 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x168 & ~x663 & ~x702 & ~x780;
assign c442 =  x2 &  x5 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x35 &  x38 &  x41 &  x44 &  x47 &  x53 &  x59 &  x62 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x152 &  x161 &  x164 &  x170 &  x173 &  x176 &  x182 &  x185 &  x188 &  x191 &  x197 &  x200 &  x203 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x254 &  x257 &  x266 &  x269 &  x272 &  x275 &  x278 &  x284 &  x287 &  x290 &  x302 &  x305 &  x308 &  x311 &  x317 &  x320 &  x323 &  x329 &  x332 &  x335 &  x338 &  x347 &  x350 &  x353 &  x356 &  x362 &  x368 &  x371 &  x374 &  x377 &  x383 &  x386 &  x389 &  x392 &  x395 &  x397 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x446 &  x449 &  x452 &  x455 &  x458 &  x464 &  x476 &  x479 &  x482 &  x485 &  x491 &  x494 &  x500 &  x503 &  x506 &  x509 &  x511 &  x512 &  x515 &  x518 &  x521 &  x524 &  x530 &  x533 &  x536 &  x542 &  x550 &  x551 &  x554 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x586 &  x587 &  x593 &  x596 &  x599 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x625 &  x626 &  x632 &  x635 &  x638 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x668 &  x674 &  x677 &  x680 &  x683 &  x692 &  x695 &  x698 &  x701 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x761 &  x770 &  x773 &  x776 &  x779 &  x782 &  x793 &  x794 &  x797 &  x803 &  x806 &  x809 &  x812 &  x815 &  x821 &  x827 &  x836 &  x839 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x926 &  x929 &  x932 &  x935 &  x941 &  x944 &  x956 &  x959 &  x962 &  x965 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x555 & ~x630 & ~x669 & ~x670 & ~x708 & ~x747;
assign c444 =  x5 &  x8 &  x11 &  x14 &  x17 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x128 &  x134 &  x137 &  x140 &  x146 &  x149 &  x152 &  x161 &  x164 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x218 &  x221 &  x224 &  x230 &  x236 &  x239 &  x242 &  x251 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x308 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x353 &  x359 &  x362 &  x368 &  x371 &  x374 &  x377 &  x389 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x471 &  x472 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x506 &  x511 &  x512 &  x515 &  x518 &  x524 &  x527 &  x530 &  x536 &  x539 &  x542 &  x545 &  x547 &  x548 &  x550 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x584 &  x586 &  x587 &  x593 &  x596 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x704 &  x710 &  x713 &  x716 &  x719 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x749 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x785 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x821 &  x824 &  x827 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x860 &  x863 &  x872 &  x878 &  x884 &  x890 &  x896 &  x902 &  x905 &  x908 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x938 &  x947 &  x953 &  x956 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x992 &  x998 &  x1001 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x156 & ~x195 & ~x234 & ~x273 & ~x312 & ~x360 & ~x438 & ~x477 & ~x630;
assign c446 =  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x26 &  x32 &  x35 &  x38 &  x44 &  x50 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x77 &  x80 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x113 &  x116 &  x119 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x152 &  x158 &  x161 &  x164 &  x173 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x239 &  x245 &  x248 &  x251 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x287 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x317 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x362 &  x368 &  x371 &  x374 &  x377 &  x386 &  x389 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x431 &  x437 &  x440 &  x443 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x512 &  x518 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x550 &  x554 &  x557 &  x563 &  x566 &  x569 &  x575 &  x578 &  x581 &  x588 &  x589 &  x590 &  x593 &  x596 &  x599 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x647 &  x650 &  x653 &  x656 &  x662 &  x664 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x695 &  x698 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x773 &  x779 &  x788 &  x794 &  x797 &  x803 &  x806 &  x809 &  x812 &  x821 &  x824 &  x827 &  x836 &  x842 &  x845 &  x857 &  x860 &  x863 &  x869 &  x875 &  x878 &  x881 &  x887 &  x893 &  x896 &  x899 &  x905 &  x911 &  x914 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x968 &  x971 &  x974 &  x980 &  x983 &  x992 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1037 &  x1043 &  x1049 &  x1052 &  x1055 &  x1058 &  x1067 &  x1073 &  x1076 &  x1079 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x273 & ~x312 & ~x351 & ~x594 & ~x645 & ~x669 & ~x684 & ~x708 & ~x709 & ~x747;
assign c448 =  x2 &  x5 &  x11 &  x20 &  x35 &  x41 &  x47 &  x50 &  x59 &  x65 &  x80 &  x83 &  x89 &  x98 &  x101 &  x104 &  x116 &  x122 &  x125 &  x134 &  x137 &  x143 &  x146 &  x152 &  x176 &  x185 &  x191 &  x200 &  x206 &  x212 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x242 &  x245 &  x248 &  x251 &  x254 &  x263 &  x269 &  x275 &  x278 &  x290 &  x299 &  x305 &  x308 &  x311 &  x320 &  x326 &  x329 &  x335 &  x341 &  x350 &  x353 &  x365 &  x368 &  x371 &  x377 &  x380 &  x392 &  x398 &  x407 &  x410 &  x422 &  x425 &  x434 &  x440 &  x443 &  x452 &  x458 &  x461 &  x467 &  x471 &  x473 &  x479 &  x485 &  x500 &  x509 &  x511 &  x524 &  x533 &  x536 &  x539 &  x545 &  x548 &  x550 &  x557 &  x563 &  x566 &  x575 &  x578 &  x584 &  x587 &  x589 &  x596 &  x599 &  x602 &  x611 &  x620 &  x623 &  x629 &  x632 &  x635 &  x638 &  x650 &  x653 &  x662 &  x665 &  x668 &  x674 &  x677 &  x680 &  x683 &  x689 &  x695 &  x701 &  x703 &  x713 &  x725 &  x734 &  x737 &  x746 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x773 &  x776 &  x782 &  x788 &  x794 &  x797 &  x800 &  x803 &  x806 &  x827 &  x830 &  x833 &  x836 &  x842 &  x848 &  x854 &  x860 &  x863 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x893 &  x896 &  x899 &  x908 &  x917 &  x920 &  x929 &  x935 &  x941 &  x944 &  x956 &  x959 &  x974 &  x983 &  x986 &  x989 &  x992 &  x998 &  x1004 &  x1013 &  x1019 &  x1022 &  x1037 &  x1052 &  x1058 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1127 & ~x234 & ~x423 & ~x747 & ~x1056;
assign c450 =  x2 &  x11 &  x14 &  x20 &  x23 &  x32 &  x35 &  x44 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x83 &  x86 &  x95 &  x98 &  x101 &  x107 &  x131 &  x137 &  x143 &  x149 &  x155 &  x158 &  x161 &  x164 &  x179 &  x185 &  x197 &  x203 &  x209 &  x218 &  x221 &  x227 &  x230 &  x251 &  x254 &  x257 &  x260 &  x269 &  x275 &  x281 &  x296 &  x305 &  x308 &  x311 &  x314 &  x329 &  x332 &  x341 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x386 &  x392 &  x395 &  x398 &  x401 &  x404 &  x410 &  x413 &  x419 &  x428 &  x443 &  x449 &  x452 &  x458 &  x467 &  x479 &  x482 &  x485 &  x494 &  x500 &  x503 &  x506 &  x509 &  x521 &  x524 &  x532 &  x533 &  x542 &  x545 &  x551 &  x554 &  x563 &  x566 &  x569 &  x587 &  x590 &  x593 &  x596 &  x611 &  x620 &  x623 &  x629 &  x638 &  x641 &  x659 &  x662 &  x665 &  x668 &  x674 &  x680 &  x695 &  x698 &  x710 &  x713 &  x716 &  x719 &  x725 &  x728 &  x731 &  x737 &  x740 &  x746 &  x755 &  x761 &  x764 &  x767 &  x770 &  x779 &  x784 &  x785 &  x788 &  x791 &  x794 &  x803 &  x806 &  x809 &  x818 &  x827 &  x848 &  x851 &  x863 &  x869 &  x872 &  x875 &  x878 &  x887 &  x896 &  x898 &  x902 &  x911 &  x914 &  x920 &  x923 &  x932 &  x935 &  x937 &  x941 &  x947 &  x950 &  x953 &  x956 &  x962 &  x971 &  x974 &  x980 &  x989 &  x992 &  x995 &  x998 &  x1010 &  x1019 &  x1031 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1064 &  x1070 &  x1076 &  x1079 &  x1088 &  x1094 &  x1097 &  x1103 &  x1106 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x234 & ~x273 & ~x312 & ~x477 & ~x657 & ~x696 & ~x774 & ~x982 & ~x1020;
assign c452 =  x1 &  x4 &  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x29 &  x32 &  x35 &  x38 &  x41 &  x43 &  x44 &  x47 &  x50 &  x53 &  x56 &  x62 &  x65 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x118 &  x122 &  x125 &  x128 &  x131 &  x134 &  x140 &  x146 &  x152 &  x155 &  x157 &  x158 &  x161 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x196 &  x197 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x242 &  x245 &  x248 &  x251 &  x257 &  x260 &  x263 &  x266 &  x274 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x314 &  x317 &  x320 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x365 &  x368 &  x374 &  x377 &  x380 &  x383 &  x389 &  x392 &  x395 &  x398 &  x401 &  x407 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x440 &  x443 &  x445 &  x446 &  x449 &  x452 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x497 &  x500 &  x506 &  x509 &  x512 &  x515 &  x518 &  x530 &  x533 &  x539 &  x548 &  x554 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x587 &  x590 &  x593 &  x599 &  x602 &  x611 &  x614 &  x617 &  x620 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x761 &  x764 &  x767 &  x770 &  x773 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x800 &  x803 &  x806 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x832 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x860 &  x863 &  x866 &  x869 &  x871 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1130 & ~x30 & ~x63 & ~x102 & ~x141 & ~x153 & ~x192 & ~x270 & ~x309 & ~x336 & ~x381 & ~x504 & ~x543;
assign c454 =  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x35 &  x53 &  x59 &  x65 &  x80 &  x83 &  x92 &  x95 &  x98 &  x107 &  x110 &  x113 &  x122 &  x131 &  x140 &  x143 &  x149 &  x155 &  x179 &  x182 &  x194 &  x197 &  x200 &  x203 &  x209 &  x218 &  x220 &  x221 &  x233 &  x236 &  x239 &  x257 &  x266 &  x272 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x305 &  x308 &  x320 &  x335 &  x341 &  x350 &  x353 &  x359 &  x365 &  x368 &  x371 &  x374 &  x383 &  x389 &  x392 &  x395 &  x404 &  x407 &  x410 &  x422 &  x431 &  x434 &  x437 &  x440 &  x446 &  x455 &  x460 &  x464 &  x473 &  x479 &  x481 &  x488 &  x493 &  x494 &  x497 &  x499 &  x500 &  x503 &  x509 &  x514 &  x524 &  x532 &  x536 &  x548 &  x551 &  x553 &  x554 &  x560 &  x563 &  x566 &  x572 &  x578 &  x584 &  x587 &  x590 &  x596 &  x599 &  x602 &  x605 &  x608 &  x614 &  x617 &  x620 &  x623 &  x629 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x662 &  x665 &  x671 &  x674 &  x677 &  x680 &  x683 &  x695 &  x698 &  x704 &  x713 &  x716 &  x719 &  x722 &  x728 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x764 &  x779 &  x791 &  x794 &  x797 &  x800 &  x803 &  x812 &  x821 &  x824 &  x839 &  x842 &  x845 &  x848 &  x851 &  x857 &  x860 &  x863 &  x869 &  x875 &  x884 &  x887 &  x893 &  x901 &  x914 &  x929 &  x935 &  x938 &  x940 &  x953 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x998 &  x1001 &  x1004 &  x1007 &  x1016 &  x1019 &  x1022 &  x1031 &  x1067 &  x1070 &  x1073 &  x1091 &  x1094 &  x1103 &  x1115 &  x1124 &  x1127 &  x1130 & ~x117 & ~x273 & ~x312 & ~x429 & ~x468 & ~x507 & ~x585 & ~x618 & ~x624 & ~x750;
assign c456 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x265 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x304 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x343 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x472 &  x473 &  x476 &  x482 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x510 &  x511 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x549 &  x550 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x589 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130 & ~x156 & ~x195 & ~x234 & ~x273 & ~x312 & ~x351 & ~x390 & ~x429 & ~x708 & ~x747 & ~x786;
assign c458 =  x2 &  x8 &  x11 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x47 &  x50 &  x53 &  x59 &  x62 &  x65 &  x68 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x107 &  x110 &  x116 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x167 &  x170 &  x173 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x236 &  x237 &  x238 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x274 &  x275 &  x277 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x308 &  x311 &  x313 &  x314 &  x316 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x341 &  x344 &  x347 &  x350 &  x352 &  x355 &  x356 &  x359 &  x365 &  x368 &  x371 &  x374 &  x380 &  x383 &  x386 &  x392 &  x395 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x434 &  x440 &  x443 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x482 &  x491 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x517 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x545 &  x548 &  x554 &  x557 &  x560 &  x566 &  x569 &  x575 &  x578 &  x581 &  x584 &  x587 &  x593 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x623 &  x629 &  x632 &  x635 &  x638 &  x641 &  x647 &  x653 &  x656 &  x662 &  x665 &  x668 &  x671 &  x677 &  x683 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x710 &  x713 &  x719 &  x722 &  x725 &  x734 &  x737 &  x740 &  x743 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x842 &  x845 &  x851 &  x854 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1006 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x357 & ~x396 & ~x397 & ~x435 & ~x666 & ~x705 & ~x706 & ~x744 & ~x783 & ~x822 & ~x897 & ~x936 & ~x975 & ~x1014 & ~x1053 & ~x1092;
assign c460 =  x8 &  x11 &  x14 &  x17 &  x29 &  x32 &  x35 &  x41 &  x53 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x98 &  x101 &  x104 &  x110 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x173 &  x179 &  x182 &  x185 &  x188 &  x200 &  x203 &  x206 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x251 &  x254 &  x260 &  x263 &  x269 &  x275 &  x278 &  x281 &  x284 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x365 &  x374 &  x377 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x419 &  x421 &  x422 &  x425 &  x428 &  x431 &  x437 &  x443 &  x446 &  x452 &  x455 &  x458 &  x460 &  x461 &  x467 &  x479 &  x485 &  x488 &  x491 &  x497 &  x499 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x542 &  x545 &  x548 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x596 &  x599 &  x602 &  x605 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x680 &  x689 &  x701 &  x704 &  x707 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x742 &  x743 &  x746 &  x749 &  x752 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x779 &  x781 &  x782 &  x784 &  x785 &  x788 &  x791 &  x794 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x854 &  x859 &  x860 &  x863 &  x866 &  x869 &  x871 &  x872 &  x878 &  x881 &  x887 &  x893 &  x896 &  x905 &  x907 &  x908 &  x910 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x953 &  x956 &  x959 &  x962 &  x968 &  x974 &  x977 &  x980 &  x983 &  x989 &  x998 &  x1010 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1100 &  x1106 &  x1109 &  x1112 &  x1121 &  x1127 & ~x468 & ~x825;
assign c462 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x28 &  x29 &  x31 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x71 &  x77 &  x80 &  x86 &  x89 &  x92 &  x98 &  x101 &  x107 &  x110 &  x113 &  x116 &  x122 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x155 &  x158 &  x164 &  x167 &  x173 &  x176 &  x179 &  x182 &  x188 &  x191 &  x194 &  x197 &  x200 &  x212 &  x218 &  x221 &  x230 &  x233 &  x242 &  x245 &  x251 &  x254 &  x256 &  x257 &  x260 &  x262 &  x263 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x292 &  x293 &  x299 &  x301 &  x302 &  x305 &  x308 &  x311 &  x314 &  x320 &  x323 &  x326 &  x329 &  x332 &  x334 &  x337 &  x338 &  x344 &  x347 &  x350 &  x353 &  x358 &  x359 &  x368 &  x371 &  x374 &  x377 &  x386 &  x392 &  x395 &  x398 &  x401 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x467 &  x479 &  x485 &  x491 &  x494 &  x497 &  x503 &  x509 &  x512 &  x518 &  x524 &  x526 &  x527 &  x530 &  x533 &  x536 &  x542 &  x545 &  x548 &  x551 &  x560 &  x563 &  x569 &  x575 &  x578 &  x581 &  x584 &  x587 &  x589 &  x590 &  x593 &  x596 &  x599 &  x602 &  x604 &  x608 &  x617 &  x620 &  x623 &  x629 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x662 &  x665 &  x668 &  x680 &  x683 &  x686 &  x689 &  x692 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x722 &  x728 &  x734 &  x737 &  x743 &  x746 &  x749 &  x758 &  x761 &  x764 &  x770 &  x773 &  x782 &  x785 &  x788 &  x794 &  x800 &  x803 &  x806 &  x809 &  x812 &  x818 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x854 &  x857 &  x860 &  x866 &  x869 &  x872 &  x874 &  x875 &  x878 &  x881 &  x887 &  x890 &  x893 &  x899 &  x902 &  x905 &  x911 &  x913 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x938 &  x944 &  x947 &  x956 &  x962 &  x965 &  x968 &  x971 &  x974 &  x983 &  x986 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x234 & ~x273 & ~x312;
assign c464 =  x8 &  x26 &  x35 &  x40 &  x41 &  x47 &  x53 &  x56 &  x68 &  x86 &  x92 &  x116 &  x149 &  x161 &  x179 &  x182 &  x185 &  x194 &  x206 &  x209 &  x227 &  x287 &  x293 &  x308 &  x311 &  x314 &  x317 &  x320 &  x350 &  x359 &  x368 &  x374 &  x386 &  x389 &  x391 &  x392 &  x398 &  x413 &  x425 &  x430 &  x434 &  x443 &  x458 &  x464 &  x467 &  x482 &  x485 &  x488 &  x494 &  x524 &  x536 &  x539 &  x560 &  x563 &  x566 &  x569 &  x578 &  x620 &  x626 &  x641 &  x644 &  x647 &  x656 &  x677 &  x683 &  x686 &  x689 &  x692 &  x704 &  x718 &  x719 &  x725 &  x728 &  x731 &  x734 &  x743 &  x746 &  x749 &  x755 &  x770 &  x779 &  x785 &  x794 &  x809 &  x818 &  x821 &  x824 &  x827 &  x830 &  x835 &  x842 &  x875 &  x886 &  x902 &  x911 &  x920 &  x926 &  x932 &  x938 &  x941 &  x944 &  x950 &  x952 &  x953 &  x956 &  x965 &  x977 &  x980 &  x983 &  x992 &  x995 &  x1001 &  x1004 &  x1016 &  x1028 &  x1031 &  x1040 &  x1049 &  x1061 &  x1073 &  x1091 &  x1100 &  x1106 &  x1118 &  x1121 &  x1127 & ~x381 & ~x504 & ~x582 & ~x708;
assign c466 =  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x38 &  x41 &  x44 &  x47 &  x50 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x83 &  x86 &  x95 &  x98 &  x104 &  x107 &  x110 &  x119 &  x122 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x155 &  x158 &  x161 &  x164 &  x167 &  x173 &  x176 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x218 &  x224 &  x227 &  x230 &  x233 &  x242 &  x245 &  x251 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x311 &  x314 &  x317 &  x319 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x362 &  x371 &  x374 &  x377 &  x383 &  x386 &  x389 &  x392 &  x394 &  x398 &  x404 &  x407 &  x410 &  x413 &  x419 &  x422 &  x425 &  x432 &  x434 &  x440 &  x443 &  x449 &  x452 &  x455 &  x464 &  x467 &  x470 &  x472 &  x473 &  x479 &  x482 &  x485 &  x488 &  x494 &  x500 &  x503 &  x506 &  x508 &  x511 &  x512 &  x515 &  x518 &  x524 &  x533 &  x536 &  x542 &  x545 &  x547 &  x551 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x584 &  x586 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x625 &  x626 &  x629 &  x632 &  x635 &  x644 &  x647 &  x650 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x704 &  x707 &  x713 &  x716 &  x719 &  x725 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x752 &  x755 &  x758 &  x761 &  x767 &  x770 &  x773 &  x776 &  x782 &  x785 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x845 &  x848 &  x854 &  x857 &  x860 &  x866 &  x872 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x950 &  x953 &  x956 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x992 &  x998 &  x1001 &  x1007 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1097 &  x1103 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1130 & ~x591 & ~x592 & ~x630 & ~x631 & ~x669;
assign c468 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x238 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x277 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x316 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x352 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x391 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x430 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x467 &  x469 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x508 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x321 & ~x435 & ~x474 & ~x475 & ~x513 & ~x514 & ~x552 & ~x591 & ~x744 & ~x783 & ~x822 & ~x861 & ~x900 & ~x939 & ~x978 & ~x1017 & ~x1056;
assign c470 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x241 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x508 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x547 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x635 &  x638 &  x641 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x321 & ~x399 & ~x438 & ~x513 & ~x552 & ~x591 & ~x825 & ~x939 & ~x978;
assign c472 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x82 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x113 &  x116 &  x119 &  x120 &  x121 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x157 &  x158 &  x160 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x196 &  x197 &  x199 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x235 &  x236 &  x238 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x274 &  x275 &  x277 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x572 &  x575 &  x578 &  x581 &  x587 &  x590 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x93 & ~x165 & ~x216 & ~x264 & ~x303 & ~x342;
assign c474 =  x11 &  x20 &  x23 &  x26 &  x38 &  x41 &  x56 &  x59 &  x68 &  x71 &  x74 &  x80 &  x86 &  x95 &  x116 &  x119 &  x120 &  x121 &  x128 &  x137 &  x143 &  x155 &  x157 &  x158 &  x159 &  x164 &  x182 &  x196 &  x198 &  x200 &  x203 &  x212 &  x215 &  x218 &  x221 &  x224 &  x236 &  x245 &  x248 &  x263 &  x277 &  x287 &  x290 &  x302 &  x308 &  x314 &  x316 &  x317 &  x332 &  x338 &  x341 &  x353 &  x365 &  x377 &  x392 &  x398 &  x404 &  x416 &  x422 &  x428 &  x431 &  x434 &  x440 &  x442 &  x443 &  x449 &  x458 &  x461 &  x464 &  x479 &  x482 &  x485 &  x491 &  x494 &  x497 &  x500 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x542 &  x551 &  x554 &  x560 &  x566 &  x572 &  x575 &  x587 &  x590 &  x596 &  x601 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x641 &  x644 &  x650 &  x653 &  x659 &  x665 &  x668 &  x679 &  x686 &  x692 &  x698 &  x701 &  x707 &  x713 &  x716 &  x718 &  x719 &  x728 &  x731 &  x740 &  x752 &  x757 &  x758 &  x764 &  x776 &  x782 &  x794 &  x796 &  x800 &  x803 &  x815 &  x818 &  x824 &  x827 &  x833 &  x835 &  x854 &  x857 &  x869 &  x871 &  x875 &  x878 &  x887 &  x890 &  x893 &  x899 &  x916 &  x917 &  x926 &  x929 &  x941 &  x944 &  x971 &  x980 &  x983 &  x989 &  x995 &  x1016 &  x1025 &  x1034 &  x1046 &  x1052 &  x1070 &  x1073 &  x1079 &  x1088 &  x1091 &  x1097 &  x1100 &  x1109 &  x1115 &  x1118 & ~x240 & ~x280 & ~x318 & ~x357 & ~x819 & ~x858;
assign c476 =  x2 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x416 &  x419 &  x422 &  x425 &  x428 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x470 &  x473 &  x476 &  x482 &  x484 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x520 &  x521 &  x523 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x545 &  x548 &  x551 &  x554 &  x557 &  x559 &  x560 &  x563 &  x569 &  x572 &  x575 &  x577 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x601 &  x602 &  x605 &  x608 &  x610 &  x611 &  x614 &  x623 &  x626 &  x629 &  x631 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x781 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x820 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x859 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x898 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x937 &  x938 &  x941 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x976 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1015 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1054 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1093 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x657 & ~x750 & ~x903;
assign c478 =  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x40 &  x44 &  x47 &  x50 &  x53 &  x56 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x79 &  x80 &  x86 &  x89 &  x92 &  x95 &  x110 &  x118 &  x119 &  x122 &  x125 &  x128 &  x131 &  x137 &  x143 &  x146 &  x149 &  x155 &  x157 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x194 &  x196 &  x203 &  x206 &  x209 &  x212 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x235 &  x239 &  x242 &  x245 &  x248 &  x251 &  x260 &  x263 &  x266 &  x269 &  x272 &  x278 &  x281 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x323 &  x325 &  x326 &  x329 &  x335 &  x341 &  x344 &  x350 &  x356 &  x359 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x395 &  x398 &  x401 &  x407 &  x416 &  x419 &  x425 &  x431 &  x434 &  x437 &  x440 &  x446 &  x449 &  x452 &  x455 &  x464 &  x467 &  x476 &  x479 &  x482 &  x485 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x523 &  x524 &  x527 &  x530 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x562 &  x566 &  x572 &  x575 &  x577 &  x578 &  x581 &  x584 &  x587 &  x593 &  x596 &  x599 &  x601 &  x602 &  x605 &  x608 &  x611 &  x614 &  x616 &  x620 &  x623 &  x626 &  x629 &  x632 &  x640 &  x643 &  x644 &  x647 &  x650 &  x653 &  x659 &  x662 &  x665 &  x668 &  x671 &  x679 &  x680 &  x686 &  x692 &  x698 &  x701 &  x704 &  x707 &  x713 &  x716 &  x719 &  x721 &  x722 &  x725 &  x728 &  x734 &  x743 &  x746 &  x749 &  x752 &  x755 &  x760 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x796 &  x799 &  x800 &  x806 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x860 &  x866 &  x871 &  x872 &  x878 &  x881 &  x887 &  x890 &  x893 &  x896 &  x902 &  x908 &  x910 &  x917 &  x920 &  x935 &  x938 &  x949 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x971 &  x980 &  x983 &  x988 &  x992 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1039 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1130 & ~x240;
assign c480 =  x2 &  x5 &  x11 &  x29 &  x32 &  x44 &  x47 &  x50 &  x56 &  x83 &  x86 &  x98 &  x125 &  x128 &  x131 &  x146 &  x152 &  x173 &  x188 &  x194 &  x197 &  x200 &  x209 &  x218 &  x227 &  x248 &  x251 &  x257 &  x260 &  x287 &  x296 &  x299 &  x302 &  x317 &  x332 &  x344 &  x362 &  x365 &  x374 &  x389 &  x395 &  x398 &  x407 &  x410 &  x422 &  x431 &  x440 &  x446 &  x452 &  x458 &  x467 &  x473 &  x479 &  x482 &  x494 &  x497 &  x503 &  x511 &  x518 &  x527 &  x536 &  x539 &  x542 &  x545 &  x548 &  x550 &  x563 &  x578 &  x581 &  x584 &  x587 &  x590 &  x599 &  x602 &  x611 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x664 &  x674 &  x698 &  x704 &  x710 &  x722 &  x725 &  x728 &  x737 &  x740 &  x742 &  x743 &  x758 &  x764 &  x770 &  x803 &  x806 &  x809 &  x829 &  x839 &  x842 &  x857 &  x866 &  x884 &  x911 &  x920 &  x923 &  x935 &  x938 &  x941 &  x953 &  x968 &  x974 &  x986 &  x1001 &  x1031 &  x1034 &  x1037 &  x1046 &  x1052 &  x1061 &  x1064 &  x1067 &  x1076 &  x1088 &  x1091 &  x1124 & ~x390 & ~x555 & ~x709 & ~x748;
assign c482 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x251 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x278 &  x281 &  x284 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x325 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x436 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x475 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x512 &  x514 &  x515 &  x518 &  x521 &  x524 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x553 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x641 &  x647 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x692 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x890 &  x893 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x354 & ~x468 & ~x507 & ~x546 & ~x585 & ~x672 & ~x711 & ~x750 & ~x751 & ~x789 & ~x801 & ~x966;
assign c484 =  x8 &  x20 &  x26 &  x35 &  x38 &  x41 &  x59 &  x62 &  x68 &  x83 &  x86 &  x92 &  x95 &  x98 &  x113 &  x116 &  x128 &  x131 &  x134 &  x146 &  x149 &  x158 &  x164 &  x167 &  x170 &  x173 &  x179 &  x185 &  x200 &  x206 &  x209 &  x215 &  x218 &  x224 &  x227 &  x236 &  x239 &  x248 &  x251 &  x257 &  x269 &  x272 &  x275 &  x281 &  x293 &  x305 &  x314 &  x317 &  x323 &  x335 &  x338 &  x344 &  x347 &  x359 &  x362 &  x365 &  x371 &  x374 &  x377 &  x383 &  x386 &  x392 &  x395 &  x398 &  x401 &  x416 &  x422 &  x437 &  x455 &  x461 &  x470 &  x521 &  x542 &  x557 &  x581 &  x587 &  x599 &  x605 &  x616 &  x626 &  x629 &  x632 &  x635 &  x641 &  x647 &  x653 &  x662 &  x680 &  x689 &  x695 &  x701 &  x716 &  x734 &  x740 &  x746 &  x755 &  x767 &  x770 &  x779 &  x788 &  x809 &  x821 &  x823 &  x830 &  x833 &  x836 &  x842 &  x845 &  x851 &  x859 &  x887 &  x898 &  x899 &  x901 &  x908 &  x911 &  x914 &  x932 &  x935 &  x938 &  x940 &  x947 &  x968 &  x977 &  x980 &  x983 &  x995 &  x1001 &  x1004 &  x1013 &  x1016 &  x1022 &  x1025 &  x1031 &  x1037 &  x1052 &  x1058 &  x1067 &  x1068 &  x1073 &  x1076 &  x1079 &  x1085 &  x1097 &  x1103 &  x1107 &  x1109 &  x1115 & ~x273 & ~x390;
assign c486 =  x2 &  x5 &  x8 &  x11 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x157 &  x158 &  x159 &  x160 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x196 &  x197 &  x198 &  x199 &  x200 &  x203 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x235 &  x236 &  x237 &  x238 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x274 &  x275 &  x277 &  x278 &  x281 &  x284 &  x290 &  x293 &  x296 &  x299 &  x302 &  x308 &  x311 &  x313 &  x314 &  x316 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x391 &  x392 &  x395 &  x398 &  x401 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x442 &  x443 &  x449 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x481 &  x482 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x640 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x679 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x718 &  x719 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x757 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x800 &  x803 &  x806 &  x809 &  x812 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x835 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x980 &  x983 &  x986 &  x989 &  x992 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x318 & ~x357 & ~x358 & ~x396 & ~x397 & ~x435 & ~x897 & ~x936;
assign c488 =  x2 &  x14 &  x17 &  x23 &  x29 &  x41 &  x44 &  x47 &  x50 &  x53 &  x65 &  x71 &  x80 &  x86 &  x95 &  x101 &  x104 &  x113 &  x116 &  x128 &  x137 &  x140 &  x143 &  x149 &  x152 &  x158 &  x173 &  x179 &  x185 &  x194 &  x200 &  x203 &  x206 &  x215 &  x218 &  x224 &  x236 &  x239 &  x260 &  x275 &  x287 &  x293 &  x308 &  x311 &  x314 &  x317 &  x329 &  x332 &  x344 &  x350 &  x356 &  x370 &  x371 &  x374 &  x380 &  x383 &  x386 &  x392 &  x395 &  x401 &  x404 &  x413 &  x416 &  x428 &  x434 &  x440 &  x446 &  x449 &  x452 &  x461 &  x473 &  x479 &  x485 &  x493 &  x494 &  x496 &  x499 &  x503 &  x506 &  x512 &  x518 &  x521 &  x524 &  x527 &  x533 &  x538 &  x539 &  x545 &  x554 &  x563 &  x590 &  x593 &  x596 &  x611 &  x617 &  x620 &  x626 &  x638 &  x641 &  x644 &  x647 &  x656 &  x659 &  x662 &  x671 &  x677 &  x680 &  x683 &  x698 &  x701 &  x704 &  x725 &  x731 &  x734 &  x737 &  x743 &  x746 &  x749 &  x755 &  x761 &  x764 &  x776 &  x781 &  x785 &  x794 &  x803 &  x809 &  x812 &  x815 &  x820 &  x827 &  x830 &  x842 &  x845 &  x851 &  x863 &  x869 &  x875 &  x878 &  x884 &  x893 &  x896 &  x899 &  x905 &  x917 &  x923 &  x929 &  x935 &  x937 &  x947 &  x950 &  x953 &  x956 &  x959 &  x968 &  x971 &  x974 &  x992 &  x998 &  x1001 &  x1013 &  x1016 &  x1019 &  x1024 &  x1037 &  x1040 &  x1046 &  x1049 &  x1061 &  x1064 &  x1070 &  x1073 &  x1082 &  x1088 &  x1091 &  x1100 &  x1103 &  x1109 &  x1115 &  x1118 &  x1124 &  x1127 &  x1130 & ~x810 & ~x843 & ~x888 & ~x1059;
assign c490 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x32 &  x35 &  x38 &  x41 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x92 &  x95 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x143 &  x146 &  x149 &  x158 &  x161 &  x164 &  x167 &  x170 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x197 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x227 &  x230 &  x233 &  x236 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x358 &  x359 &  x362 &  x368 &  x371 &  x374 &  x377 &  x383 &  x386 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x455 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x506 &  x509 &  x512 &  x515 &  x518 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x581 &  x584 &  x587 &  x590 &  x599 &  x601 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x635 &  x638 &  x640 &  x647 &  x650 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x707 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x845 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x898 &  x899 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x120 & ~x159 & ~x696 & ~x855 & ~x933 & ~x1059 & ~x1098;
assign c492 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x703 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x742 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x781 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x871 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x910 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x946 &  x947 &  x949 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1030 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x723 & ~x747 & ~x762 & ~x786 & ~x801 & ~x840;
assign c494 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x23 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x227 &  x233 &  x239 &  x242 &  x245 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x464 &  x470 &  x473 &  x475 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x527 &  x530 &  x533 &  x539 &  x545 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x589 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x627 &  x628 &  x629 &  x632 &  x635 &  x638 &  x641 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x667 &  x668 &  x671 &  x674 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x703 &  x704 &  x706 &  x710 &  x716 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x785 &  x788 &  x791 &  x794 &  x809 &  x812 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1067 &  x1070 &  x1076 &  x1082 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x195 & ~x234 & ~x273 & ~x312 & ~x351 & ~x390 & ~x429 & ~x468 & ~x507 & ~x555 & ~x594 & ~x633 & ~x708 & ~x747;
assign c496 =  x5 &  x8 &  x20 &  x23 &  x26 &  x32 &  x35 &  x38 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x121 &  x122 &  x128 &  x131 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x157 &  x158 &  x160 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x196 &  x198 &  x199 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x227 &  x230 &  x233 &  x235 &  x236 &  x238 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x266 &  x269 &  x272 &  x274 &  x275 &  x276 &  x277 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x305 &  x311 &  x313 &  x314 &  x315 &  x317 &  x320 &  x323 &  x329 &  x332 &  x335 &  x341 &  x344 &  x350 &  x352 &  x353 &  x355 &  x356 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x386 &  x389 &  x392 &  x394 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x481 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x506 &  x509 &  x512 &  x517 &  x518 &  x521 &  x527 &  x530 &  x533 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x617 &  x620 &  x623 &  x626 &  x629 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x679 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x710 &  x713 &  x716 &  x718 &  x719 &  x722 &  x728 &  x734 &  x737 &  x740 &  x743 &  x749 &  x752 &  x755 &  x757 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x833 &  x836 &  x839 &  x842 &  x845 &  x863 &  x866 &  x869 &  x872 &  x875 &  x881 &  x887 &  x893 &  x896 &  x899 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x950 &  x953 &  x956 &  x962 &  x965 &  x971 &  x977 &  x983 &  x986 &  x989 &  x992 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x357 & ~x396 & ~x397;
assign c498 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x164 &  x170 &  x176 &  x179 &  x182 &  x188 &  x197 &  x200 &  x206 &  x212 &  x215 &  x218 &  x221 &  x227 &  x230 &  x233 &  x238 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x277 &  x278 &  x284 &  x287 &  x290 &  x293 &  x296 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x353 &  x356 &  x362 &  x365 &  x368 &  x374 &  x377 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x419 &  x422 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x452 &  x458 &  x464 &  x470 &  x473 &  x476 &  x479 &  x482 &  x488 &  x494 &  x500 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x575 &  x578 &  x581 &  x587 &  x590 &  x599 &  x602 &  x605 &  x608 &  x614 &  x617 &  x620 &  x626 &  x632 &  x638 &  x641 &  x644 &  x650 &  x653 &  x656 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x689 &  x692 &  x695 &  x701 &  x707 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x827 &  x833 &  x836 &  x839 &  x842 &  x848 &  x851 &  x854 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x905 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x968 &  x971 &  x974 &  x980 &  x986 &  x989 &  x992 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1022 &  x1025 &  x1028 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x54 & ~x55 & ~x72 & ~x93 & ~x126 & ~x588 & ~x744 & ~x783 & ~x822 & ~x861 & ~x900 & ~x936 & ~x939 & ~x975 & ~x1014 & ~x1053 & ~x1056 & ~x1092 & ~x1095 & ~x1107;
assign c4100 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x80 &  x89 &  x95 &  x101 &  x107 &  x110 &  x113 &  x116 &  x119 &  x121 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x146 &  x149 &  x152 &  x155 &  x159 &  x160 &  x161 &  x164 &  x170 &  x173 &  x179 &  x185 &  x188 &  x191 &  x194 &  x196 &  x198 &  x199 &  x200 &  x206 &  x209 &  x212 &  x215 &  x221 &  x227 &  x233 &  x235 &  x238 &  x239 &  x242 &  x245 &  x251 &  x257 &  x266 &  x269 &  x272 &  x274 &  x275 &  x278 &  x281 &  x284 &  x287 &  x299 &  x302 &  x308 &  x311 &  x317 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x352 &  x359 &  x362 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x419 &  x425 &  x428 &  x431 &  x437 &  x440 &  x452 &  x455 &  x458 &  x461 &  x467 &  x470 &  x476 &  x482 &  x485 &  x491 &  x494 &  x497 &  x503 &  x506 &  x509 &  x512 &  x518 &  x521 &  x523 &  x530 &  x536 &  x545 &  x548 &  x551 &  x554 &  x560 &  x566 &  x569 &  x575 &  x578 &  x581 &  x587 &  x590 &  x601 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x632 &  x635 &  x638 &  x644 &  x650 &  x656 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x704 &  x707 &  x710 &  x713 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x764 &  x767 &  x770 &  x776 &  x785 &  x788 &  x791 &  x794 &  x800 &  x812 &  x815 &  x821 &  x827 &  x833 &  x835 &  x836 &  x839 &  x842 &  x851 &  x854 &  x860 &  x863 &  x871 &  x872 &  x878 &  x887 &  x902 &  x905 &  x911 &  x914 &  x917 &  x920 &  x926 &  x935 &  x938 &  x941 &  x947 &  x950 &  x953 &  x956 &  x962 &  x968 &  x971 &  x974 &  x977 &  x980 &  x986 &  x992 &  x998 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1037 &  x1039 &  x1040 &  x1043 &  x1049 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1078 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x279 & ~x318 & ~x357 & ~x501 & ~x780 & ~x858 & ~x897 & ~x936 & ~x1014;
assign c4102 =  x2 &  x5 &  x8 &  x14 &  x20 &  x26 &  x32 &  x35 &  x38 &  x41 &  x50 &  x53 &  x56 &  x62 &  x68 &  x71 &  x80 &  x83 &  x86 &  x95 &  x107 &  x110 &  x116 &  x119 &  x122 &  x125 &  x128 &  x137 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x173 &  x182 &  x191 &  x215 &  x218 &  x221 &  x224 &  x233 &  x236 &  x242 &  x248 &  x254 &  x257 &  x263 &  x275 &  x281 &  x284 &  x287 &  x290 &  x296 &  x311 &  x317 &  x320 &  x323 &  x326 &  x332 &  x335 &  x338 &  x341 &  x344 &  x359 &  x365 &  x368 &  x374 &  x377 &  x383 &  x395 &  x398 &  x407 &  x410 &  x413 &  x416 &  x431 &  x433 &  x440 &  x449 &  x452 &  x455 &  x458 &  x461 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x494 &  x497 &  x500 &  x503 &  x506 &  x512 &  x515 &  x518 &  x524 &  x527 &  x530 &  x533 &  x539 &  x545 &  x547 &  x551 &  x557 &  x560 &  x575 &  x584 &  x590 &  x596 &  x599 &  x605 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x632 &  x635 &  x638 &  x647 &  x650 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x680 &  x689 &  x695 &  x704 &  x719 &  x725 &  x728 &  x734 &  x752 &  x755 &  x758 &  x761 &  x776 &  x779 &  x794 &  x797 &  x806 &  x809 &  x815 &  x827 &  x830 &  x833 &  x857 &  x860 &  x866 &  x869 &  x872 &  x878 &  x884 &  x899 &  x902 &  x905 &  x911 &  x914 &  x920 &  x929 &  x932 &  x935 &  x941 &  x953 &  x956 &  x965 &  x971 &  x974 &  x977 &  x983 &  x986 &  x989 &  x998 &  x1004 &  x1019 &  x1022 &  x1031 &  x1037 &  x1040 &  x1046 &  x1052 &  x1058 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1115 &  x1124 &  x1130 & ~x156 & ~x405 & ~x438 & ~x456 & ~x534 & ~x591 & ~x618 & ~x657 & ~x696;
assign c4104 =  x2 &  x5 &  x8 &  x11 &  x23 &  x26 &  x32 &  x38 &  x41 &  x44 &  x47 &  x53 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x95 &  x98 &  x104 &  x107 &  x110 &  x113 &  x116 &  x118 &  x119 &  x122 &  x128 &  x131 &  x140 &  x143 &  x146 &  x149 &  x155 &  x157 &  x158 &  x161 &  x170 &  x179 &  x185 &  x188 &  x191 &  x194 &  x196 &  x197 &  x200 &  x203 &  x209 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x242 &  x245 &  x251 &  x254 &  x263 &  x266 &  x269 &  x272 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x320 &  x323 &  x326 &  x329 &  x335 &  x341 &  x344 &  x347 &  x356 &  x359 &  x368 &  x374 &  x377 &  x383 &  x389 &  x392 &  x395 &  x401 &  x404 &  x406 &  x407 &  x410 &  x413 &  x419 &  x425 &  x434 &  x437 &  x440 &  x455 &  x461 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x491 &  x494 &  x497 &  x503 &  x506 &  x509 &  x515 &  x521 &  x530 &  x533 &  x539 &  x545 &  x548 &  x551 &  x554 &  x562 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x614 &  x617 &  x623 &  x626 &  x629 &  x635 &  x638 &  x644 &  x647 &  x650 &  x659 &  x662 &  x671 &  x677 &  x679 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x704 &  x707 &  x710 &  x716 &  x725 &  x728 &  x731 &  x734 &  x737 &  x743 &  x746 &  x749 &  x752 &  x758 &  x764 &  x770 &  x773 &  x776 &  x779 &  x782 &  x791 &  x794 &  x809 &  x812 &  x815 &  x824 &  x827 &  x830 &  x839 &  x842 &  x845 &  x851 &  x854 &  x857 &  x860 &  x869 &  x872 &  x875 &  x878 &  x884 &  x887 &  x890 &  x893 &  x902 &  x905 &  x908 &  x911 &  x917 &  x923 &  x926 &  x935 &  x938 &  x941 &  x944 &  x950 &  x956 &  x959 &  x962 &  x965 &  x977 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1013 &  x1016 &  x1028 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1082 &  x1085 &  x1088 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x264 & ~x336 & ~x348 & ~x423 & ~x588 & ~x627 & ~x774;
assign c4106 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x71 &  x74 &  x77 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x125 &  x131 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x155 &  x158 &  x161 &  x167 &  x170 &  x176 &  x179 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x218 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x323 &  x326 &  x332 &  x338 &  x341 &  x344 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x407 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x440 &  x443 &  x446 &  x449 &  x455 &  x461 &  x464 &  x467 &  x473 &  x479 &  x482 &  x485 &  x488 &  x494 &  x497 &  x500 &  x503 &  x506 &  x508 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x530 &  x533 &  x536 &  x539 &  x545 &  x547 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x677 &  x680 &  x683 &  x689 &  x695 &  x698 &  x701 &  x707 &  x710 &  x713 &  x715 &  x716 &  x719 &  x725 &  x728 &  x731 &  x737 &  x740 &  x743 &  x746 &  x752 &  x753 &  x754 &  x755 &  x761 &  x764 &  x767 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x793 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x815 &  x821 &  x824 &  x827 &  x830 &  x836 &  x842 &  x845 &  x848 &  x854 &  x857 &  x863 &  x869 &  x874 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x950 &  x952 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1079 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130 & ~x441 & ~x591 & ~x783 & ~x861;
assign c4108 =  x2 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x47 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x116 &  x128 &  x137 &  x140 &  x143 &  x149 &  x152 &  x161 &  x164 &  x167 &  x170 &  x185 &  x188 &  x194 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x230 &  x233 &  x236 &  x239 &  x242 &  x251 &  x254 &  x257 &  x260 &  x263 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x296 &  x299 &  x305 &  x308 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x341 &  x344 &  x350 &  x353 &  x359 &  x362 &  x365 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x398 &  x401 &  x404 &  x407 &  x413 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x472 &  x473 &  x476 &  x479 &  x488 &  x491 &  x494 &  x503 &  x506 &  x509 &  x511 &  x512 &  x515 &  x518 &  x521 &  x542 &  x548 &  x550 &  x554 &  x557 &  x563 &  x566 &  x569 &  x572 &  x575 &  x589 &  x590 &  x593 &  x599 &  x602 &  x605 &  x608 &  x611 &  x617 &  x620 &  x623 &  x626 &  x629 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x656 &  x662 &  x665 &  x671 &  x674 &  x683 &  x686 &  x692 &  x695 &  x698 &  x704 &  x716 &  x719 &  x722 &  x725 &  x728 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x767 &  x770 &  x776 &  x782 &  x785 &  x790 &  x791 &  x794 &  x797 &  x800 &  x806 &  x809 &  x812 &  x818 &  x821 &  x824 &  x827 &  x830 &  x839 &  x842 &  x845 &  x848 &  x857 &  x860 &  x866 &  x869 &  x872 &  x884 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x941 &  x950 &  x956 &  x959 &  x962 &  x968 &  x971 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1010 &  x1013 &  x1019 &  x1022 &  x1031 &  x1034 &  x1040 &  x1043 &  x1052 &  x1058 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1121 &  x1127 &  x1130 & ~x273 & ~x312 & ~x630 & ~x783 & ~x810 & ~x822 & ~x849 & ~x861;
assign c4110 =  x2 &  x5 &  x8 &  x11 &  x14 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x40 &  x44 &  x47 &  x56 &  x59 &  x65 &  x68 &  x71 &  x74 &  x77 &  x79 &  x80 &  x83 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x116 &  x118 &  x119 &  x122 &  x128 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x157 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x185 &  x191 &  x196 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x235 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x260 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x305 &  x308 &  x311 &  x313 &  x314 &  x317 &  x323 &  x329 &  x332 &  x335 &  x341 &  x347 &  x350 &  x353 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x407 &  x413 &  x422 &  x428 &  x431 &  x434 &  x437 &  x442 &  x443 &  x449 &  x455 &  x461 &  x464 &  x467 &  x473 &  x476 &  x479 &  x491 &  x494 &  x500 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x530 &  x548 &  x551 &  x554 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x596 &  x599 &  x601 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x623 &  x626 &  x632 &  x638 &  x640 &  x644 &  x647 &  x653 &  x656 &  x659 &  x665 &  x668 &  x674 &  x677 &  x679 &  x680 &  x686 &  x692 &  x695 &  x698 &  x704 &  x710 &  x713 &  x716 &  x718 &  x722 &  x728 &  x734 &  x743 &  x746 &  x757 &  x758 &  x761 &  x764 &  x767 &  x770 &  x776 &  x782 &  x788 &  x791 &  x797 &  x799 &  x800 &  x809 &  x815 &  x818 &  x821 &  x824 &  x827 &  x833 &  x836 &  x839 &  x842 &  x848 &  x854 &  x857 &  x863 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x899 &  x902 &  x905 &  x908 &  x911 &  x916 &  x920 &  x923 &  x932 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x989 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1097 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x279 & ~x396 & ~x435 & ~x471 & ~x588 & ~x627 & ~x666 & ~x705 & ~x744 & ~x783 & ~x822;
assign c4112 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x59 &  x62 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x155 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x209 &  x212 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x341 &  x347 &  x350 &  x353 &  x356 &  x362 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x542 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x668 &  x671 &  x674 &  x680 &  x683 &  x686 &  x692 &  x695 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x773 &  x776 &  x779 &  x782 &  x788 &  x791 &  x794 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x830 &  x836 &  x839 &  x842 &  x845 &  x848 &  x854 &  x857 &  x863 &  x869 &  x871 &  x872 &  x875 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x315 & ~x390 & ~x462 & ~x468 & ~x501 & ~x516 & ~x555 & ~x594 & ~x633 & ~x768;
assign c4114 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x59 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x272 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x302 &  x305 &  x308 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x394 &  x395 &  x398 &  x401 &  x404 &  x407 &  x413 &  x419 &  x425 &  x428 &  x431 &  x433 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x455 &  x458 &  x464 &  x467 &  x470 &  x476 &  x479 &  x482 &  x488 &  x491 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x545 &  x548 &  x551 &  x554 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x617 &  x620 &  x623 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x893 &  x896 &  x902 &  x905 &  x908 &  x911 &  x917 &  x920 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x971 &  x974 &  x977 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x0 & ~x39 & ~x78 & ~x117 & ~x267 & ~x321 & ~x552 & ~x591 & ~x630 & ~x783 & ~x822 & ~x861 & ~x900 & ~x939 & ~x1053 & ~x1092;
assign c4116 =  x22 &  x38 &  x41 &  x53 &  x71 &  x80 &  x86 &  x92 &  x104 &  x113 &  x119 &  x133 &  x137 &  x164 &  x167 &  x203 &  x206 &  x250 &  x260 &  x266 &  x272 &  x281 &  x290 &  x295 &  x296 &  x305 &  x307 &  x335 &  x341 &  x353 &  x368 &  x374 &  x392 &  x398 &  x407 &  x416 &  x440 &  x485 &  x488 &  x496 &  x515 &  x527 &  x560 &  x563 &  x569 &  x572 &  x575 &  x577 &  x590 &  x602 &  x626 &  x629 &  x632 &  x644 &  x653 &  x662 &  x668 &  x671 &  x698 &  x701 &  x728 &  x743 &  x752 &  x764 &  x767 &  x773 &  x781 &  x797 &  x800 &  x809 &  x812 &  x815 &  x820 &  x830 &  x839 &  x842 &  x845 &  x848 &  x851 &  x859 &  x869 &  x872 &  x881 &  x893 &  x896 &  x905 &  x917 &  x920 &  x926 &  x929 &  x944 &  x956 &  x971 &  x989 &  x1019 &  x1025 &  x1028 &  x1037 &  x1049 &  x1064 &  x1076 &  x1091 &  x1100 &  x1109 &  x1112 &  x1124 & ~x237 & ~x1056;
assign c4118 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x265 &  x266 &  x269 &  x272 &  x275 &  x278 &  x284 &  x287 &  x290 &  x293 &  x296 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x433 &  x434 &  x437 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x472 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x508 &  x509 &  x511 &  x512 &  x515 &  x518 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x550 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x830 &  x833 &  x836 &  x839 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x896 &  x899 &  x905 &  x908 &  x911 &  x917 &  x920 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x273 & ~x312 & ~x438 & ~x630 & ~x783;
assign c4120 =  x11 &  x14 &  x23 &  x35 &  x56 &  x67 &  x100 &  x116 &  x119 &  x122 &  x167 &  x191 &  x209 &  x223 &  x230 &  x245 &  x251 &  x287 &  x323 &  x371 &  x377 &  x416 &  x425 &  x443 &  x479 &  x485 &  x590 &  x602 &  x650 &  x662 &  x689 &  x692 &  x704 &  x818 &  x884 &  x899 &  x923 &  x941 &  x947 &  x952 &  x965 &  x1030 &  x1040 &  x1052 &  x1061 &  x1076 &  x1081 &  x1088 &  x1103 &  x1113 &  x1126 & ~x504 & ~x777;
assign c4122 =  x2 &  x5 &  x8 &  x17 &  x20 &  x29 &  x35 &  x38 &  x41 &  x44 &  x56 &  x65 &  x71 &  x92 &  x95 &  x101 &  x104 &  x116 &  x119 &  x128 &  x134 &  x137 &  x146 &  x149 &  x152 &  x155 &  x164 &  x167 &  x176 &  x179 &  x194 &  x206 &  x209 &  x212 &  x218 &  x230 &  x233 &  x236 &  x248 &  x260 &  x266 &  x272 &  x284 &  x287 &  x289 &  x290 &  x296 &  x299 &  x305 &  x308 &  x314 &  x320 &  x323 &  x326 &  x329 &  x338 &  x347 &  x359 &  x362 &  x365 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x392 &  x395 &  x398 &  x401 &  x416 &  x419 &  x422 &  x428 &  x437 &  x440 &  x449 &  x452 &  x455 &  x458 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x491 &  x494 &  x500 &  x506 &  x530 &  x533 &  x539 &  x563 &  x575 &  x581 &  x590 &  x602 &  x611 &  x620 &  x623 &  x626 &  x632 &  x635 &  x638 &  x647 &  x659 &  x665 &  x668 &  x671 &  x680 &  x683 &  x689 &  x692 &  x701 &  x703 &  x704 &  x707 &  x710 &  x713 &  x719 &  x722 &  x734 &  x743 &  x749 &  x755 &  x761 &  x767 &  x770 &  x773 &  x781 &  x785 &  x791 &  x800 &  x824 &  x827 &  x839 &  x845 &  x848 &  x851 &  x854 &  x857 &  x863 &  x869 &  x872 &  x875 &  x881 &  x893 &  x898 &  x908 &  x911 &  x914 &  x920 &  x923 &  x935 &  x937 &  x941 &  x947 &  x950 &  x952 &  x956 &  x962 &  x968 &  x977 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1019 &  x1022 &  x1031 &  x1037 &  x1049 &  x1055 &  x1069 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1094 &  x1097 &  x1100 &  x1106 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 &  x1130 & ~x438 & ~x804 & ~x816 & ~x849 & ~x855 & ~x903 & ~x942 & ~x1011 & ~x1050;
assign c4124 =  x2 &  x14 &  x21 &  x34 &  x110 &  x138 &  x176 &  x179 &  x188 &  x245 &  x256 &  x262 &  x272 &  x299 &  x302 &  x307 &  x311 &  x314 &  x317 &  x320 &  x323 &  x353 &  x359 &  x374 &  x440 &  x457 &  x461 &  x467 &  x470 &  x485 &  x488 &  x491 &  x497 &  x506 &  x533 &  x542 &  x566 &  x575 &  x578 &  x626 &  x665 &  x668 &  x704 &  x719 &  x764 &  x767 &  x773 &  x791 &  x806 &  x827 &  x845 &  x860 &  x898 &  x899 &  x902 &  x911 &  x920 &  x938 &  x947 &  x959 &  x1061 &  x1088 &  x1115 &  x1121;
assign c4126 =  x17 &  x20 &  x26 &  x62 &  x68 &  x71 &  x92 &  x98 &  x104 &  x107 &  x122 &  x134 &  x161 &  x164 &  x173 &  x198 &  x206 &  x239 &  x242 &  x248 &  x254 &  x260 &  x263 &  x272 &  x274 &  x278 &  x316 &  x332 &  x335 &  x344 &  x350 &  x365 &  x368 &  x383 &  x404 &  x410 &  x416 &  x419 &  x440 &  x446 &  x461 &  x512 &  x515 &  x521 &  x530 &  x545 &  x551 &  x560 &  x563 &  x581 &  x590 &  x593 &  x617 &  x629 &  x638 &  x644 &  x650 &  x653 &  x659 &  x665 &  x668 &  x671 &  x674 &  x677 &  x698 &  x731 &  x740 &  x746 &  x767 &  x776 &  x797 &  x818 &  x821 &  x824 &  x827 &  x866 &  x869 &  x887 &  x890 &  x908 &  x926 &  x932 &  x938 &  x947 &  x962 &  x983 &  x998 &  x1004 &  x1016 &  x1019 &  x1025 &  x1031 &  x1046 &  x1064 &  x1079 &  x1091 &  x1097 &  x1121 &  x1127 &  x1130 & ~x129 & ~x381 & ~x420 & ~x666 & ~x862;
assign c4128 =  x8 &  x11 &  x17 &  x20 &  x29 &  x35 &  x41 &  x44 &  x59 &  x62 &  x65 &  x71 &  x74 &  x83 &  x86 &  x89 &  x92 &  x95 &  x101 &  x107 &  x110 &  x122 &  x124 &  x128 &  x146 &  x160 &  x161 &  x164 &  x170 &  x173 &  x176 &  x179 &  x185 &  x194 &  x197 &  x198 &  x209 &  x218 &  x221 &  x227 &  x233 &  x238 &  x239 &  x245 &  x251 &  x254 &  x260 &  x266 &  x275 &  x278 &  x287 &  x290 &  x293 &  x305 &  x308 &  x314 &  x317 &  x320 &  x326 &  x332 &  x341 &  x344 &  x350 &  x362 &  x365 &  x371 &  x389 &  x392 &  x395 &  x401 &  x422 &  x425 &  x440 &  x446 &  x455 &  x458 &  x461 &  x470 &  x473 &  x476 &  x488 &  x491 &  x494 &  x506 &  x512 &  x518 &  x521 &  x527 &  x530 &  x548 &  x560 &  x575 &  x581 &  x587 &  x593 &  x596 &  x605 &  x614 &  x623 &  x629 &  x632 &  x638 &  x647 &  x650 &  x656 &  x662 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x713 &  x719 &  x725 &  x728 &  x737 &  x758 &  x764 &  x773 &  x782 &  x797 &  x803 &  x818 &  x824 &  x830 &  x833 &  x839 &  x848 &  x863 &  x866 &  x869 &  x875 &  x881 &  x884 &  x902 &  x905 &  x908 &  x914 &  x917 &  x926 &  x938 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x977 &  x980 &  x983 &  x986 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1022 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1052 &  x1055 &  x1061 &  x1064 &  x1073 &  x1082 &  x1094 &  x1100 &  x1106 &  x1109 &  x1112 &  x1124 &  x1130 & ~x192 & ~x210 & ~x783 & ~x822 & ~x900;
assign c4130 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x80 &  x89 &  x92 &  x98 &  x107 &  x110 &  x113 &  x116 &  x119 &  x120 &  x121 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x155 &  x157 &  x158 &  x159 &  x160 &  x161 &  x164 &  x167 &  x170 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x196 &  x197 &  x198 &  x199 &  x200 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x235 &  x236 &  x245 &  x248 &  x251 &  x260 &  x263 &  x266 &  x275 &  x277 &  x284 &  x290 &  x293 &  x296 &  x299 &  x305 &  x311 &  x313 &  x314 &  x316 &  x317 &  x320 &  x329 &  x332 &  x341 &  x344 &  x347 &  x350 &  x352 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x410 &  x413 &  x422 &  x428 &  x431 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x473 &  x476 &  x482 &  x491 &  x494 &  x497 &  x500 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x530 &  x539 &  x542 &  x545 &  x554 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x590 &  x593 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x632 &  x635 &  x638 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x779 &  x785 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x839 &  x842 &  x845 &  x848 &  x854 &  x860 &  x869 &  x872 &  x875 &  x878 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x920 &  x923 &  x926 &  x929 &  x932 &  x938 &  x941 &  x947 &  x950 &  x953 &  x956 &  x965 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1097 &  x1100 &  x1103 &  x1109 &  x1115 &  x1118 &  x1124 &  x1127 & ~x165 & ~x166 & ~x204 & ~x240 & ~x280 & ~x318 & ~x357 & ~x396 & ~x474;
assign c4132 =  x2 &  x8 &  x14 &  x20 &  x23 &  x29 &  x32 &  x35 &  x38 &  x44 &  x47 &  x50 &  x59 &  x62 &  x71 &  x74 &  x77 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x116 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x173 &  x179 &  x188 &  x194 &  x197 &  x200 &  x203 &  x205 &  x206 &  x209 &  x212 &  x218 &  x221 &  x224 &  x227 &  x233 &  x239 &  x244 &  x245 &  x248 &  x257 &  x263 &  x269 &  x272 &  x278 &  x287 &  x290 &  x293 &  x296 &  x302 &  x308 &  x311 &  x314 &  x317 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x386 &  x392 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x434 &  x443 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x476 &  x479 &  x482 &  x485 &  x487 &  x488 &  x494 &  x497 &  x499 &  x500 &  x503 &  x509 &  x512 &  x518 &  x524 &  x526 &  x527 &  x530 &  x533 &  x538 &  x539 &  x542 &  x545 &  x548 &  x551 &  x557 &  x560 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x608 &  x614 &  x617 &  x620 &  x626 &  x635 &  x638 &  x641 &  x647 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x674 &  x683 &  x686 &  x689 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x722 &  x725 &  x728 &  x731 &  x740 &  x743 &  x755 &  x758 &  x767 &  x773 &  x776 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x806 &  x809 &  x812 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x878 &  x884 &  x887 &  x893 &  x896 &  x901 &  x902 &  x908 &  x911 &  x917 &  x920 &  x923 &  x926 &  x932 &  x938 &  x944 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x974 &  x977 &  x983 &  x986 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1054 &  x1058 &  x1061 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1124 &  x1127 & ~x276 & ~x315 & ~x429 & ~x468 & ~x507 & ~x546 & ~x750;
assign c4134 =  x2 &  x8 &  x11 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x107 &  x110 &  x113 &  x116 &  x119 &  x125 &  x131 &  x134 &  x137 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x194 &  x197 &  x206 &  x209 &  x212 &  x218 &  x227 &  x233 &  x236 &  x238 &  x239 &  x245 &  x248 &  x254 &  x257 &  x260 &  x263 &  x269 &  x272 &  x277 &  x278 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x316 &  x317 &  x320 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x350 &  x353 &  x355 &  x356 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x404 &  x410 &  x416 &  x419 &  x425 &  x428 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x476 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x644 &  x647 &  x650 &  x653 &  x656 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x683 &  x686 &  x689 &  x695 &  x701 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x731 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x884 &  x887 &  x893 &  x896 &  x902 &  x905 &  x908 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x944 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x995 &  x998 &  x1007 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1100 &  x1103 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x15 & ~x435 & ~x474 & ~x475 & ~x513 & ~x528 & ~x591 & ~x606 & ~x744 & ~x783 & ~x822 & ~x1056;
assign c4136 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x364 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x832 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x870 &  x871 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x126 & ~x429 & ~x468 & ~x825 & ~x840 & ~x879;
assign c4138 =  x2 &  x11 &  x14 &  x17 &  x20 &  x23 &  x29 &  x38 &  x41 &  x47 &  x50 &  x53 &  x68 &  x71 &  x89 &  x92 &  x98 &  x104 &  x110 &  x116 &  x119 &  x125 &  x128 &  x131 &  x137 &  x140 &  x146 &  x155 &  x170 &  x176 &  x179 &  x182 &  x185 &  x191 &  x194 &  x197 &  x206 &  x215 &  x224 &  x227 &  x233 &  x245 &  x263 &  x266 &  x275 &  x278 &  x281 &  x284 &  x299 &  x308 &  x314 &  x320 &  x326 &  x329 &  x332 &  x344 &  x350 &  x356 &  x362 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x392 &  x401 &  x404 &  x406 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x445 &  x461 &  x470 &  x473 &  x479 &  x482 &  x488 &  x491 &  x497 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x554 &  x557 &  x560 &  x566 &  x569 &  x578 &  x581 &  x584 &  x590 &  x596 &  x599 &  x602 &  x605 &  x611 &  x614 &  x617 &  x620 &  x626 &  x629 &  x635 &  x641 &  x647 &  x650 &  x653 &  x659 &  x665 &  x668 &  x674 &  x677 &  x683 &  x689 &  x692 &  x695 &  x698 &  x701 &  x710 &  x722 &  x725 &  x728 &  x731 &  x740 &  x749 &  x755 &  x761 &  x767 &  x770 &  x776 &  x785 &  x788 &  x791 &  x797 &  x800 &  x803 &  x812 &  x815 &  x821 &  x824 &  x836 &  x842 &  x845 &  x851 &  x854 &  x857 &  x860 &  x866 &  x874 &  x875 &  x881 &  x890 &  x896 &  x898 &  x905 &  x908 &  x913 &  x914 &  x917 &  x923 &  x926 &  x935 &  x938 &  x947 &  x953 &  x956 &  x962 &  x965 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x1004 &  x1007 &  x1019 &  x1028 &  x1040 &  x1043 &  x1046 &  x1061 &  x1064 &  x1073 &  x1076 &  x1079 &  x1088 &  x1091 &  x1097 &  x1106 &  x1115 &  x1121 &  x1124 &  x1127 & ~x129 & ~x135 & ~x168 & ~x285 & ~x777 & ~x804;
assign c4140 =  x20 &  x32 &  x41 &  x47 &  x50 &  x68 &  x77 &  x92 &  x98 &  x104 &  x110 &  x122 &  x128 &  x131 &  x143 &  x161 &  x170 &  x173 &  x176 &  x179 &  x182 &  x188 &  x203 &  x209 &  x227 &  x245 &  x257 &  x266 &  x269 &  x275 &  x281 &  x284 &  x299 &  x314 &  x319 &  x332 &  x371 &  x401 &  x404 &  x413 &  x431 &  x432 &  x452 &  x479 &  x518 &  x530 &  x548 &  x550 &  x551 &  x554 &  x572 &  x587 &  x602 &  x625 &  x629 &  x632 &  x638 &  x671 &  x677 &  x680 &  x698 &  x710 &  x713 &  x770 &  x782 &  x788 &  x800 &  x824 &  x836 &  x851 &  x872 &  x875 &  x881 &  x893 &  x911 &  x926 &  x932 &  x935 &  x947 &  x950 &  x1007 &  x1025 &  x1037 &  x1073 &  x1094 &  x1100 &  x1103 &  x1115 & ~x438 & ~x504;
assign c4142 =  x2 &  x5 &  x8 &  x11 &  x32 &  x44 &  x47 &  x59 &  x62 &  x68 &  x74 &  x77 &  x83 &  x95 &  x98 &  x104 &  x110 &  x113 &  x116 &  x119 &  x125 &  x131 &  x134 &  x140 &  x143 &  x146 &  x149 &  x152 &  x176 &  x179 &  x182 &  x185 &  x197 &  x200 &  x203 &  x206 &  x209 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x242 &  x257 &  x260 &  x269 &  x278 &  x284 &  x287 &  x299 &  x302 &  x308 &  x314 &  x317 &  x326 &  x329 &  x335 &  x338 &  x344 &  x350 &  x358 &  x362 &  x365 &  x368 &  x371 &  x386 &  x392 &  x395 &  x401 &  x404 &  x407 &  x413 &  x416 &  x419 &  x422 &  x431 &  x434 &  x440 &  x449 &  x455 &  x458 &  x464 &  x467 &  x471 &  x472 &  x482 &  x485 &  x488 &  x491 &  x497 &  x500 &  x511 &  x512 &  x515 &  x521 &  x524 &  x527 &  x530 &  x536 &  x542 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x587 &  x590 &  x596 &  x602 &  x605 &  x608 &  x614 &  x632 &  x641 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x689 &  x698 &  x704 &  x710 &  x713 &  x719 &  x722 &  x725 &  x728 &  x731 &  x737 &  x740 &  x746 &  x749 &  x752 &  x758 &  x761 &  x764 &  x767 &  x770 &  x776 &  x782 &  x788 &  x791 &  x797 &  x815 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x845 &  x851 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x896 &  x920 &  x929 &  x935 &  x938 &  x941 &  x947 &  x953 &  x956 &  x965 &  x971 &  x974 &  x980 &  x983 &  x986 &  x995 &  x1004 &  x1010 &  x1016 &  x1022 &  x1025 &  x1031 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1064 &  x1076 &  x1094 &  x1100 &  x1103 &  x1109 &  x1115 &  x1118 &  x1121 &  x1130 & ~x234 & ~x273 & ~x438 & ~x478 & ~x516 & ~x591;
assign c4144 =  x2 &  x5 &  x8 &  x11 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x218 &  x224 &  x227 &  x230 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x394 &  x395 &  x398 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x428 &  x431 &  x433 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x470 &  x472 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x547 &  x548 &  x551 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x674 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x704 &  x707 &  x710 &  x713 &  x722 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x761 &  x764 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x806 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x860 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x890 &  x893 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x959 &  x962 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x156 & ~x195 & ~x234 & ~x273 & ~x360 & ~x363 & ~x477 & ~x591 & ~x618;
assign c4146 =  x2 &  x8 &  x11 &  x14 &  x17 &  x23 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x56 &  x59 &  x62 &  x65 &  x68 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x122 &  x128 &  x134 &  x137 &  x143 &  x146 &  x152 &  x155 &  x158 &  x164 &  x170 &  x176 &  x179 &  x188 &  x191 &  x194 &  x203 &  x206 &  x212 &  x215 &  x218 &  x224 &  x227 &  x233 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x263 &  x269 &  x281 &  x284 &  x287 &  x296 &  x305 &  x308 &  x311 &  x314 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x341 &  x344 &  x350 &  x353 &  x356 &  x359 &  x365 &  x368 &  x374 &  x377 &  x383 &  x389 &  x398 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x452 &  x455 &  x461 &  x470 &  x473 &  x476 &  x482 &  x491 &  x497 &  x500 &  x503 &  x506 &  x512 &  x518 &  x524 &  x527 &  x533 &  x536 &  x538 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x593 &  x599 &  x602 &  x608 &  x626 &  x629 &  x635 &  x638 &  x641 &  x647 &  x653 &  x656 &  x659 &  x662 &  x668 &  x671 &  x674 &  x680 &  x686 &  x689 &  x692 &  x695 &  x704 &  x707 &  x716 &  x725 &  x728 &  x734 &  x737 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x779 &  x782 &  x788 &  x791 &  x800 &  x803 &  x806 &  x809 &  x815 &  x821 &  x827 &  x833 &  x839 &  x842 &  x845 &  x869 &  x878 &  x884 &  x887 &  x893 &  x902 &  x908 &  x920 &  x929 &  x932 &  x935 &  x944 &  x947 &  x950 &  x953 &  x956 &  x968 &  x974 &  x986 &  x989 &  x992 &  x995 &  x1007 &  x1013 &  x1019 &  x1022 &  x1034 &  x1037 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 & ~x813 & ~x891 & ~x930 & ~x943 & ~x981 & ~x1008 & ~x1009 & ~x1098;
assign c4148 =  x17 &  x20 &  x47 &  x53 &  x62 &  x65 &  x74 &  x77 &  x80 &  x86 &  x101 &  x122 &  x125 &  x131 &  x146 &  x155 &  x158 &  x163 &  x173 &  x179 &  x185 &  x191 &  x194 &  x203 &  x221 &  x236 &  x241 &  x248 &  x251 &  x269 &  x272 &  x279 &  x280 &  x287 &  x293 &  x302 &  x323 &  x332 &  x341 &  x347 &  x353 &  x359 &  x362 &  x368 &  x374 &  x380 &  x386 &  x392 &  x410 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x446 &  x452 &  x455 &  x458 &  x461 &  x470 &  x476 &  x479 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x524 &  x533 &  x536 &  x542 &  x548 &  x557 &  x566 &  x569 &  x575 &  x596 &  x602 &  x605 &  x611 &  x626 &  x665 &  x668 &  x698 &  x701 &  x704 &  x707 &  x710 &  x722 &  x734 &  x740 &  x743 &  x746 &  x758 &  x761 &  x764 &  x767 &  x779 &  x785 &  x818 &  x821 &  x824 &  x830 &  x833 &  x836 &  x842 &  x851 &  x863 &  x878 &  x884 &  x887 &  x893 &  x896 &  x902 &  x907 &  x908 &  x938 &  x941 &  x947 &  x949 &  x956 &  x965 &  x971 &  x983 &  x998 &  x1001 &  x1004 &  x1019 &  x1025 &  x1028 &  x1049 &  x1061 &  x1073 &  x1076 &  x1079 &  x1091 &  x1094 &  x1106 &  x1121 &  x1124 &  x1127 &  x1130 & ~x1056 & ~x1095;
assign c4150 =  x2 &  x8 &  x11 &  x14 &  x26 &  x29 &  x32 &  x35 &  x38 &  x47 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x77 &  x86 &  x89 &  x95 &  x98 &  x101 &  x110 &  x116 &  x125 &  x131 &  x134 &  x140 &  x143 &  x152 &  x155 &  x158 &  x163 &  x167 &  x170 &  x173 &  x179 &  x181 &  x182 &  x185 &  x188 &  x191 &  x194 &  x200 &  x202 &  x203 &  x206 &  x212 &  x215 &  x218 &  x220 &  x221 &  x224 &  x230 &  x239 &  x241 &  x248 &  x251 &  x254 &  x260 &  x263 &  x275 &  x293 &  x296 &  x302 &  x311 &  x317 &  x320 &  x329 &  x332 &  x335 &  x344 &  x356 &  x362 &  x365 &  x371 &  x374 &  x389 &  x398 &  x401 &  x404 &  x407 &  x410 &  x416 &  x422 &  x428 &  x431 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x458 &  x461 &  x464 &  x467 &  x473 &  x476 &  x482 &  x485 &  x491 &  x494 &  x497 &  x506 &  x512 &  x518 &  x527 &  x530 &  x545 &  x557 &  x566 &  x569 &  x572 &  x578 &  x596 &  x599 &  x605 &  x608 &  x611 &  x614 &  x617 &  x623 &  x632 &  x635 &  x638 &  x644 &  x647 &  x656 &  x662 &  x668 &  x671 &  x686 &  x689 &  x692 &  x695 &  x701 &  x710 &  x713 &  x716 &  x719 &  x728 &  x743 &  x749 &  x755 &  x767 &  x773 &  x782 &  x785 &  x800 &  x803 &  x809 &  x812 &  x818 &  x827 &  x830 &  x833 &  x839 &  x842 &  x848 &  x854 &  x860 &  x869 &  x871 &  x875 &  x878 &  x881 &  x890 &  x896 &  x899 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x941 &  x944 &  x950 &  x953 &  x956 &  x959 &  x968 &  x971 &  x974 &  x977 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1052 &  x1055 &  x1058 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x360 & ~x399 & ~x450 & ~x528 & ~x567 & ~x1095;
assign c4152 =  x2 &  x8 &  x20 &  x23 &  x26 &  x32 &  x35 &  x47 &  x50 &  x53 &  x59 &  x62 &  x65 &  x71 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x98 &  x104 &  x107 &  x110 &  x116 &  x119 &  x125 &  x131 &  x134 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x218 &  x224 &  x227 &  x230 &  x236 &  x242 &  x245 &  x251 &  x254 &  x260 &  x263 &  x269 &  x272 &  x275 &  x278 &  x281 &  x287 &  x290 &  x293 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x329 &  x332 &  x334 &  x335 &  x338 &  x341 &  x344 &  x350 &  x353 &  x356 &  x358 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x392 &  x395 &  x401 &  x404 &  x407 &  x410 &  x413 &  x419 &  x422 &  x425 &  x428 &  x431 &  x436 &  x437 &  x440 &  x449 &  x455 &  x461 &  x467 &  x470 &  x475 &  x476 &  x482 &  x487 &  x490 &  x491 &  x500 &  x506 &  x509 &  x512 &  x518 &  x521 &  x524 &  x526 &  x527 &  x533 &  x536 &  x542 &  x548 &  x551 &  x553 &  x554 &  x557 &  x560 &  x563 &  x565 &  x569 &  x575 &  x578 &  x581 &  x587 &  x593 &  x599 &  x605 &  x608 &  x611 &  x617 &  x620 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x674 &  x689 &  x691 &  x692 &  x698 &  x701 &  x704 &  x706 &  x713 &  x716 &  x719 &  x722 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x745 &  x746 &  x749 &  x752 &  x761 &  x764 &  x767 &  x770 &  x776 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x821 &  x823 &  x827 &  x830 &  x836 &  x839 &  x842 &  x848 &  x851 &  x854 &  x860 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x890 &  x893 &  x899 &  x902 &  x905 &  x908 &  x914 &  x923 &  x929 &  x938 &  x941 &  x944 &  x947 &  x950 &  x956 &  x959 &  x968 &  x971 &  x974 &  x980 &  x983 &  x986 &  x989 &  x991 &  x992 &  x995 &  x998 &  x1001 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1058 &  x1061 &  x1064 &  x1076 &  x1082 &  x1088 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1118 &  x1124 &  x1130 & ~x843;
assign c4154 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x316 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x354 &  x355 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x391 &  x392 &  x394 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x430 &  x431 &  x433 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x469 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x508 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x547 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x952 &  x953 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x399 & ~x435 & ~x474 & ~x513 & ~x514 & ~x552 & ~x591;
assign c4156 =  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x32 &  x35 &  x38 &  x41 &  x44 &  x56 &  x65 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x110 &  x113 &  x116 &  x119 &  x125 &  x131 &  x134 &  x137 &  x140 &  x143 &  x149 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x179 &  x182 &  x185 &  x188 &  x194 &  x197 &  x203 &  x209 &  x215 &  x218 &  x224 &  x227 &  x233 &  x236 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x266 &  x272 &  x275 &  x278 &  x281 &  x284 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x335 &  x347 &  x356 &  x359 &  x362 &  x368 &  x374 &  x377 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x440 &  x443 &  x446 &  x449 &  x452 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x515 &  x524 &  x533 &  x536 &  x542 &  x545 &  x551 &  x557 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x593 &  x596 &  x602 &  x605 &  x608 &  x620 &  x623 &  x626 &  x629 &  x635 &  x638 &  x641 &  x656 &  x659 &  x662 &  x664 &  x668 &  x683 &  x689 &  x695 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x728 &  x731 &  x741 &  x742 &  x746 &  x749 &  x755 &  x758 &  x764 &  x767 &  x770 &  x773 &  x776 &  x781 &  x788 &  x791 &  x797 &  x800 &  x809 &  x815 &  x820 &  x824 &  x827 &  x829 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x860 &  x863 &  x868 &  x869 &  x872 &  x875 &  x881 &  x887 &  x890 &  x893 &  x899 &  x908 &  x911 &  x917 &  x923 &  x929 &  x938 &  x950 &  x953 &  x956 &  x965 &  x968 &  x971 &  x977 &  x980 &  x983 &  x986 &  x989 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1073 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1112 &  x1121 &  x1127 & ~x594 & ~x621 & ~x708 & ~x747 & ~x771 & ~x786 & ~x810 & ~x825 & ~x849 & ~x1038;
assign c4158 =  x2 &  x8 &  x11 &  x14 &  x17 &  x20 &  x29 &  x32 &  x35 &  x38 &  x41 &  x47 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x89 &  x92 &  x98 &  x101 &  x107 &  x110 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x143 &  x146 &  x149 &  x151 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x206 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x245 &  x251 &  x254 &  x257 &  x260 &  x266 &  x275 &  x281 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x323 &  x326 &  x335 &  x338 &  x344 &  x350 &  x353 &  x356 &  x359 &  x362 &  x368 &  x371 &  x374 &  x377 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x443 &  x446 &  x449 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x509 &  x512 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x557 &  x560 &  x566 &  x569 &  x572 &  x578 &  x581 &  x587 &  x590 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x698 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x743 &  x746 &  x749 &  x758 &  x770 &  x773 &  x779 &  x785 &  x788 &  x791 &  x793 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x854 &  x857 &  x863 &  x866 &  x875 &  x878 &  x881 &  x887 &  x890 &  x896 &  x899 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x926 &  x932 &  x938 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x983 &  x989 &  x991 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1121 &  x1124 &  x1127 &  x1130 & ~x351 & ~x390 & ~x429 & ~x516 & ~x555 & ~x556 & ~x594;
assign c4160 =  x2 &  x11 &  x17 &  x20 &  x29 &  x35 &  x38 &  x41 &  x44 &  x59 &  x71 &  x74 &  x80 &  x83 &  x92 &  x95 &  x98 &  x104 &  x110 &  x113 &  x125 &  x128 &  x134 &  x176 &  x179 &  x191 &  x194 &  x200 &  x209 &  x212 &  x218 &  x224 &  x230 &  x239 &  x245 &  x248 &  x260 &  x263 &  x284 &  x302 &  x308 &  x320 &  x323 &  x338 &  x341 &  x365 &  x368 &  x377 &  x383 &  x398 &  x407 &  x413 &  x416 &  x419 &  x437 &  x440 &  x446 &  x449 &  x458 &  x467 &  x479 &  x485 &  x491 &  x497 &  x506 &  x509 &  x512 &  x518 &  x521 &  x530 &  x536 &  x539 &  x542 &  x548 &  x551 &  x554 &  x557 &  x578 &  x590 &  x596 &  x602 &  x614 &  x620 &  x626 &  x635 &  x644 &  x656 &  x662 &  x665 &  x667 &  x668 &  x671 &  x674 &  x680 &  x706 &  x707 &  x710 &  x719 &  x725 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x767 &  x773 &  x776 &  x779 &  x781 &  x785 &  x788 &  x794 &  x800 &  x803 &  x812 &  x815 &  x820 &  x821 &  x839 &  x857 &  x860 &  x871 &  x884 &  x893 &  x899 &  x905 &  x914 &  x920 &  x935 &  x941 &  x953 &  x956 &  x968 &  x971 &  x992 &  x995 &  x1001 &  x1013 &  x1028 &  x1037 &  x1040 &  x1085 &  x1106 &  x1108 &  x1112 &  x1118 &  x1124 &  x1130 & ~x273 & ~x312 & ~x351 & ~x594 & ~x633 & ~x960 & ~x999;
assign c4162 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x382 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x482 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x698 &  x701 &  x703 &  x704 &  x707 &  x710 &  x713 &  x719 &  x722 &  x728 &  x731 &  x734 &  x737 &  x740 &  x742 &  x743 &  x746 &  x749 &  x752 &  x758 &  x761 &  x764 &  x767 &  x773 &  x776 &  x779 &  x781 &  x782 &  x785 &  x788 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x820 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x907 &  x908 &  x910 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x989 &  x992 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x351 & ~x747 & ~x786 & ~x787 & ~x825 & ~x826 & ~x864 & ~x865 & ~x903 & ~x904 & ~x942;
assign c4164 =  x2 &  x8 &  x11 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x44 &  x53 &  x62 &  x65 &  x68 &  x74 &  x80 &  x83 &  x89 &  x101 &  x104 &  x110 &  x116 &  x119 &  x125 &  x128 &  x134 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x173 &  x176 &  x179 &  x184 &  x188 &  x194 &  x200 &  x203 &  x212 &  x215 &  x218 &  x223 &  x236 &  x242 &  x245 &  x248 &  x251 &  x254 &  x266 &  x269 &  x275 &  x278 &  x281 &  x287 &  x290 &  x293 &  x302 &  x305 &  x308 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x335 &  x338 &  x341 &  x344 &  x350 &  x353 &  x362 &  x365 &  x368 &  x377 &  x380 &  x383 &  x386 &  x389 &  x407 &  x410 &  x413 &  x425 &  x428 &  x443 &  x449 &  x455 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x485 &  x497 &  x500 &  x503 &  x506 &  x515 &  x518 &  x521 &  x523 &  x524 &  x527 &  x533 &  x542 &  x548 &  x557 &  x560 &  x562 &  x566 &  x572 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x614 &  x617 &  x626 &  x635 &  x647 &  x650 &  x656 &  x665 &  x668 &  x677 &  x683 &  x689 &  x695 &  x698 &  x701 &  x707 &  x710 &  x716 &  x718 &  x719 &  x722 &  x731 &  x734 &  x737 &  x740 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x815 &  x818 &  x821 &  x824 &  x833 &  x835 &  x839 &  x842 &  x851 &  x854 &  x857 &  x863 &  x866 &  x871 &  x872 &  x874 &  x875 &  x878 &  x884 &  x893 &  x896 &  x902 &  x910 &  x911 &  x914 &  x919 &  x920 &  x932 &  x944 &  x950 &  x953 &  x956 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x983 &  x986 &  x992 &  x995 &  x1001 &  x1007 &  x1013 &  x1019 &  x1028 &  x1034 &  x1037 &  x1040 &  x1042 &  x1046 &  x1049 &  x1052 &  x1061 &  x1063 &  x1067 &  x1070 &  x1073 &  x1079 &  x1081 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1108 &  x1109 &  x1114 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x900 & ~x939 & ~x978 & ~x1017 & ~x1056;
assign c4166 =  x2 &  x5 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x41 &  x53 &  x59 &  x65 &  x71 &  x80 &  x92 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x128 &  x131 &  x134 &  x137 &  x152 &  x158 &  x161 &  x170 &  x173 &  x176 &  x182 &  x191 &  x197 &  x203 &  x206 &  x212 &  x215 &  x218 &  x221 &  x233 &  x236 &  x239 &  x248 &  x254 &  x257 &  x263 &  x269 &  x272 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x323 &  x326 &  x329 &  x335 &  x341 &  x344 &  x350 &  x356 &  x359 &  x362 &  x368 &  x371 &  x377 &  x380 &  x383 &  x389 &  x392 &  x398 &  x401 &  x404 &  x410 &  x416 &  x419 &  x425 &  x428 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x470 &  x473 &  x476 &  x479 &  x484 &  x488 &  x491 &  x503 &  x509 &  x515 &  x518 &  x521 &  x527 &  x530 &  x539 &  x542 &  x548 &  x554 &  x557 &  x560 &  x563 &  x566 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x601 &  x608 &  x611 &  x617 &  x620 &  x626 &  x629 &  x631 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x653 &  x656 &  x659 &  x665 &  x671 &  x674 &  x680 &  x683 &  x689 &  x701 &  x704 &  x707 &  x719 &  x722 &  x731 &  x734 &  x743 &  x746 &  x749 &  x752 &  x755 &  x764 &  x767 &  x770 &  x773 &  x776 &  x782 &  x788 &  x797 &  x803 &  x806 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x881 &  x884 &  x899 &  x908 &  x917 &  x923 &  x929 &  x932 &  x935 &  x936 &  x937 &  x938 &  x941 &  x947 &  x950 &  x953 &  x956 &  x959 &  x968 &  x971 &  x974 &  x977 &  x983 &  x989 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1015 &  x1016 &  x1028 &  x1031 &  x1040 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1073 &  x1076 &  x1079 &  x1085 &  x1091 &  x1093 &  x1097 &  x1100 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1130 & ~x996 & ~x1020 & ~x1059 & ~x1099;
assign c4168 =  x2 &  x14 &  x17 &  x20 &  x35 &  x47 &  x50 &  x53 &  x59 &  x62 &  x68 &  x80 &  x86 &  x92 &  x98 &  x107 &  x110 &  x113 &  x116 &  x119 &  x125 &  x131 &  x134 &  x137 &  x140 &  x149 &  x152 &  x157 &  x158 &  x159 &  x161 &  x167 &  x170 &  x176 &  x179 &  x188 &  x191 &  x200 &  x203 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x238 &  x245 &  x251 &  x254 &  x257 &  x263 &  x272 &  x275 &  x277 &  x281 &  x284 &  x293 &  x299 &  x302 &  x305 &  x326 &  x332 &  x335 &  x338 &  x344 &  x350 &  x362 &  x374 &  x377 &  x386 &  x389 &  x395 &  x404 &  x407 &  x410 &  x416 &  x422 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x455 &  x458 &  x470 &  x476 &  x479 &  x488 &  x494 &  x497 &  x500 &  x512 &  x515 &  x521 &  x530 &  x536 &  x539 &  x542 &  x545 &  x551 &  x554 &  x566 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x599 &  x602 &  x605 &  x611 &  x623 &  x635 &  x641 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x665 &  x677 &  x680 &  x683 &  x689 &  x695 &  x698 &  x701 &  x704 &  x716 &  x728 &  x731 &  x740 &  x746 &  x752 &  x758 &  x773 &  x776 &  x779 &  x785 &  x788 &  x791 &  x794 &  x803 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x836 &  x845 &  x851 &  x854 &  x857 &  x860 &  x869 &  x872 &  x878 &  x884 &  x887 &  x893 &  x896 &  x899 &  x902 &  x908 &  x911 &  x914 &  x920 &  x923 &  x926 &  x929 &  x938 &  x947 &  x950 &  x953 &  x956 &  x962 &  x968 &  x971 &  x974 &  x977 &  x980 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1034 &  x1037 &  x1040 &  x1049 &  x1052 &  x1085 &  x1088 &  x1097 &  x1103 &  x1109 &  x1115 &  x1124 &  x1127 &  x1130 & ~x165 & ~x294 & ~x333 & ~x342 & ~x357 & ~x420 & ~x744;
assign c4170 =  x2 &  x8 &  x32 &  x38 &  x41 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x86 &  x92 &  x95 &  x101 &  x104 &  x110 &  x116 &  x119 &  x131 &  x134 &  x137 &  x149 &  x158 &  x161 &  x164 &  x182 &  x188 &  x191 &  x194 &  x196 &  x200 &  x203 &  x206 &  x209 &  x221 &  x227 &  x233 &  x242 &  x248 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x299 &  x305 &  x311 &  x317 &  x326 &  x329 &  x332 &  x344 &  x347 &  x350 &  x356 &  x362 &  x365 &  x367 &  x368 &  x374 &  x377 &  x380 &  x383 &  x386 &  x395 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x445 &  x452 &  x455 &  x458 &  x464 &  x467 &  x482 &  x485 &  x491 &  x494 &  x500 &  x503 &  x506 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x542 &  x545 &  x551 &  x557 &  x562 &  x563 &  x566 &  x572 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x608 &  x614 &  x617 &  x623 &  x626 &  x629 &  x632 &  x635 &  x647 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x677 &  x689 &  x695 &  x698 &  x704 &  x707 &  x710 &  x713 &  x716 &  x718 &  x719 &  x722 &  x725 &  x731 &  x734 &  x740 &  x743 &  x746 &  x755 &  x758 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x796 &  x803 &  x806 &  x809 &  x821 &  x824 &  x833 &  x835 &  x845 &  x851 &  x857 &  x860 &  x874 &  x881 &  x890 &  x896 &  x902 &  x905 &  x911 &  x913 &  x914 &  x920 &  x929 &  x932 &  x937 &  x938 &  x941 &  x950 &  x952 &  x956 &  x962 &  x968 &  x980 &  x983 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1067 &  x1073 &  x1079 &  x1085 &  x1088 &  x1091 &  x1093 &  x1094 &  x1097 &  x1108 &  x1109 &  x1115 &  x1118 &  x1124 &  x1127 &  x1130 & ~x75 & ~x129 & ~x324 & ~x810 & ~x894;
assign c4172 =  x2 &  x5 &  x8 &  x11 &  x17 &  x19 &  x20 &  x23 &  x26 &  x35 &  x47 &  x59 &  x62 &  x65 &  x68 &  x74 &  x86 &  x92 &  x101 &  x104 &  x107 &  x110 &  x128 &  x131 &  x134 &  x140 &  x146 &  x149 &  x155 &  x158 &  x161 &  x179 &  x182 &  x185 &  x188 &  x197 &  x200 &  x209 &  x215 &  x221 &  x224 &  x226 &  x227 &  x233 &  x236 &  x239 &  x242 &  x260 &  x263 &  x265 &  x266 &  x269 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x299 &  x305 &  x314 &  x320 &  x329 &  x341 &  x350 &  x359 &  x362 &  x365 &  x371 &  x382 &  x383 &  x386 &  x392 &  x401 &  x404 &  x407 &  x431 &  x434 &  x437 &  x440 &  x442 &  x449 &  x461 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x487 &  x488 &  x491 &  x497 &  x500 &  x503 &  x506 &  x512 &  x520 &  x536 &  x548 &  x557 &  x563 &  x565 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x590 &  x596 &  x599 &  x602 &  x608 &  x620 &  x623 &  x638 &  x644 &  x649 &  x656 &  x659 &  x665 &  x668 &  x689 &  x707 &  x710 &  x725 &  x731 &  x746 &  x752 &  x755 &  x761 &  x767 &  x770 &  x773 &  x779 &  x791 &  x803 &  x806 &  x809 &  x821 &  x827 &  x848 &  x851 &  x863 &  x875 &  x878 &  x881 &  x911 &  x914 &  x920 &  x923 &  x926 &  x932 &  x938 &  x941 &  x950 &  x956 &  x959 &  x965 &  x971 &  x974 &  x977 &  x986 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1016 &  x1025 &  x1034 &  x1037 &  x1043 &  x1049 &  x1058 &  x1064 &  x1070 &  x1085 &  x1088 &  x1091 &  x1094 &  x1100 &  x1109 &  x1112 &  x1121 &  x1127 & ~x750 & ~x1008;
assign c4174 =  x5 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x41 &  x47 &  x50 &  x53 &  x56 &  x62 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x92 &  x95 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x152 &  x155 &  x158 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x191 &  x194 &  x197 &  x200 &  x203 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x287 &  x290 &  x299 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x377 &  x380 &  x383 &  x389 &  x392 &  x395 &  x398 &  x401 &  x407 &  x410 &  x413 &  x416 &  x425 &  x434 &  x455 &  x458 &  x461 &  x464 &  x467 &  x485 &  x488 &  x494 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x539 &  x545 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x632 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x674 &  x677 &  x680 &  x683 &  x689 &  x692 &  x698 &  x701 &  x710 &  x716 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x758 &  x764 &  x770 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x806 &  x809 &  x812 &  x815 &  x818 &  x820 &  x821 &  x824 &  x827 &  x830 &  x842 &  x845 &  x848 &  x851 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x884 &  x887 &  x890 &  x899 &  x905 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x941 &  x947 &  x950 &  x953 &  x959 &  x962 &  x965 &  x968 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x995 &  x1001 &  x1004 &  x1007 &  x1022 &  x1025 &  x1028 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1115 &  x1121 &  x1127 &  x1130 & ~x54 & ~x132 & ~x282 & ~x288 & ~x384 & ~x609 & ~x771 & ~x978;
assign c4176 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x23 &  x26 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x56 &  x59 &  x62 &  x68 &  x71 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x152 &  x158 &  x161 &  x164 &  x170 &  x173 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x254 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x596 &  x599 &  x602 &  x604 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x638 &  x641 &  x644 &  x647 &  x650 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x719 &  x722 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x752 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x781 &  x782 &  x785 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x941 &  x944 &  x947 &  x949 &  x950 &  x956 &  x959 &  x962 &  x965 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x405 & ~x444 & ~x540 & ~x579 & ~x1056;
assign c4178 =  x2 &  x8 &  x11 &  x14 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x41 &  x47 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x80 &  x86 &  x89 &  x92 &  x95 &  x98 &  x104 &  x107 &  x110 &  x113 &  x116 &  x122 &  x125 &  x131 &  x140 &  x143 &  x146 &  x149 &  x161 &  x170 &  x173 &  x176 &  x179 &  x188 &  x197 &  x203 &  x206 &  x209 &  x215 &  x218 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x326 &  x329 &  x332 &  x335 &  x341 &  x344 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x380 &  x383 &  x389 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x431 &  x434 &  x437 &  x440 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x485 &  x488 &  x491 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x563 &  x569 &  x578 &  x581 &  x587 &  x590 &  x593 &  x596 &  x602 &  x605 &  x617 &  x626 &  x629 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x659 &  x665 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x722 &  x725 &  x728 &  x731 &  x734 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x764 &  x767 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x794 &  x797 &  x800 &  x803 &  x809 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x839 &  x842 &  x845 &  x848 &  x854 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x896 &  x899 &  x902 &  x908 &  x911 &  x914 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1061 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x351 & ~x507 & ~x690 & ~x774 & ~x804 & ~x813 & ~x960 & ~x966 & ~x981 & ~x1005 & ~x1077;
assign c4180 =  x2 &  x5 &  x8 &  x11 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x50 &  x59 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x104 &  x110 &  x113 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x143 &  x146 &  x149 &  x152 &  x155 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x187 &  x188 &  x194 &  x197 &  x200 &  x206 &  x221 &  x224 &  x230 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x272 &  x278 &  x281 &  x284 &  x287 &  x293 &  x299 &  x302 &  x305 &  x314 &  x317 &  x320 &  x326 &  x329 &  x335 &  x338 &  x341 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x374 &  x383 &  x386 &  x389 &  x392 &  x394 &  x395 &  x398 &  x404 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x472 &  x473 &  x476 &  x479 &  x482 &  x485 &  x491 &  x494 &  x497 &  x500 &  x503 &  x509 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x548 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x584 &  x586 &  x587 &  x590 &  x596 &  x599 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x625 &  x629 &  x632 &  x635 &  x638 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x710 &  x713 &  x719 &  x722 &  x728 &  x731 &  x734 &  x737 &  x740 &  x746 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x788 &  x791 &  x793 &  x794 &  x797 &  x800 &  x803 &  x809 &  x815 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x854 &  x857 &  x863 &  x866 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x893 &  x896 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x968 &  x971 &  x974 &  x983 &  x989 &  x995 &  x998 &  x1004 &  x1007 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x708 & ~x709 & ~x747;
assign c4182 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x23 &  x29 &  x35 &  x38 &  x41 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x116 &  x119 &  x122 &  x125 &  x128 &  x134 &  x137 &  x140 &  x146 &  x152 &  x158 &  x161 &  x164 &  x170 &  x176 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x212 &  x215 &  x221 &  x224 &  x227 &  x233 &  x236 &  x242 &  x248 &  x254 &  x257 &  x260 &  x263 &  x266 &  x272 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x302 &  x308 &  x314 &  x317 &  x320 &  x323 &  x329 &  x332 &  x338 &  x341 &  x343 &  x344 &  x347 &  x350 &  x356 &  x359 &  x365 &  x368 &  x371 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x419 &  x422 &  x434 &  x443 &  x446 &  x449 &  x458 &  x461 &  x467 &  x476 &  x479 &  x482 &  x485 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x542 &  x545 &  x548 &  x550 &  x551 &  x554 &  x557 &  x563 &  x566 &  x575 &  x578 &  x581 &  x584 &  x587 &  x593 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x668 &  x671 &  x674 &  x680 &  x689 &  x692 &  x695 &  x701 &  x703 &  x707 &  x710 &  x716 &  x719 &  x725 &  x728 &  x731 &  x734 &  x737 &  x742 &  x743 &  x749 &  x752 &  x755 &  x764 &  x767 &  x770 &  x776 &  x779 &  x782 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x857 &  x860 &  x863 &  x866 &  x872 &  x875 &  x878 &  x887 &  x890 &  x893 &  x905 &  x911 &  x914 &  x917 &  x920 &  x926 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x953 &  x956 &  x959 &  x968 &  x974 &  x980 &  x983 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1022 &  x1028 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1112 &  x1124 &  x1127 & ~x195 & ~x234 & ~x273 & ~x312 & ~x351 & ~x390 & ~x483 & ~x594 & ~x708 & ~x807 & ~x846;
assign c4184 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x43 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x82 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x120 &  x121 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x157 &  x158 &  x159 &  x160 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x196 &  x199 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x235 &  x236 &  x237 &  x238 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x274 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x955 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x501 & ~x621 & ~x840;
assign c4186 =  x8 &  x11 &  x14 &  x17 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x53 &  x59 &  x62 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x194 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x278 &  x281 &  x284 &  x290 &  x293 &  x296 &  x299 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x368 &  x371 &  x374 &  x377 &  x380 &  x382 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x437 &  x440 &  x446 &  x449 &  x452 &  x455 &  x458 &  x460 &  x461 &  x464 &  x467 &  x470 &  x473 &  x479 &  x485 &  x488 &  x494 &  x497 &  x499 &  x500 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x560 &  x563 &  x566 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x593 &  x596 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x628 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x656 &  x659 &  x665 &  x667 &  x668 &  x671 &  x674 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x701 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x722 &  x725 &  x728 &  x731 &  x737 &  x740 &  x743 &  x745 &  x746 &  x749 &  x752 &  x758 &  x761 &  x767 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x815 &  x821 &  x823 &  x824 &  x827 &  x833 &  x836 &  x842 &  x845 &  x848 &  x851 &  x860 &  x862 &  x866 &  x869 &  x872 &  x875 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x901 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x949 &  x950 &  x953 &  x956 &  x962 &  x965 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 & ~x351 & ~x825 & ~x826 & ~x864 & ~x903;
assign c4188 =  x2 &  x5 &  x11 &  x14 &  x17 &  x20 &  x35 &  x44 &  x62 &  x77 &  x83 &  x89 &  x95 &  x113 &  x116 &  x122 &  x128 &  x134 &  x137 &  x143 &  x149 &  x176 &  x179 &  x182 &  x188 &  x197 &  x200 &  x206 &  x218 &  x227 &  x236 &  x239 &  x245 &  x251 &  x254 &  x257 &  x266 &  x287 &  x290 &  x296 &  x299 &  x305 &  x311 &  x317 &  x326 &  x332 &  x338 &  x344 &  x347 &  x350 &  x356 &  x362 &  x374 &  x380 &  x383 &  x386 &  x389 &  x395 &  x410 &  x416 &  x419 &  x422 &  x431 &  x440 &  x443 &  x452 &  x455 &  x473 &  x476 &  x479 &  x482 &  x506 &  x527 &  x542 &  x554 &  x557 &  x563 &  x572 &  x575 &  x584 &  x593 &  x596 &  x599 &  x611 &  x614 &  x617 &  x635 &  x638 &  x656 &  x659 &  x662 &  x671 &  x674 &  x680 &  x704 &  x728 &  x734 &  x740 &  x745 &  x755 &  x758 &  x764 &  x767 &  x779 &  x794 &  x797 &  x806 &  x809 &  x815 &  x820 &  x839 &  x881 &  x884 &  x893 &  x896 &  x898 &  x905 &  x914 &  x917 &  x920 &  x935 &  x941 &  x947 &  x956 &  x959 &  x965 &  x971 &  x977 &  x980 &  x983 &  x989 &  x992 &  x998 &  x1001 &  x1004 &  x1010 &  x1019 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1055 &  x1058 &  x1073 &  x1082 &  x1088 &  x1103 &  x1124 &  x1130 & ~x312 & ~x585 & ~x789 & ~x904 & ~x943 & ~x981;
assign c4190 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x22 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x61 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x137 &  x140 &  x146 &  x149 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x223 &  x224 &  x229 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x254 &  x257 &  x260 &  x263 &  x266 &  x268 &  x269 &  x271 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x301 &  x302 &  x308 &  x311 &  x314 &  x320 &  x323 &  x326 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x376 &  x377 &  x380 &  x383 &  x389 &  x392 &  x395 &  x398 &  x401 &  x403 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x431 &  x434 &  x437 &  x440 &  x442 &  x443 &  x446 &  x449 &  x452 &  x454 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x493 &  x494 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x643 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x722 &  x728 &  x731 &  x734 &  x737 &  x740 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x874 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x905 &  x908 &  x911 &  x913 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1108 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130;
assign c4192 =  x8 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x41 &  x47 &  x50 &  x56 &  x59 &  x65 &  x80 &  x86 &  x92 &  x104 &  x110 &  x113 &  x134 &  x137 &  x143 &  x152 &  x158 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x191 &  x194 &  x197 &  x203 &  x212 &  x218 &  x221 &  x233 &  x236 &  x239 &  x245 &  x248 &  x251 &  x260 &  x263 &  x266 &  x269 &  x272 &  x284 &  x287 &  x290 &  x302 &  x308 &  x314 &  x317 &  x329 &  x335 &  x338 &  x344 &  x350 &  x353 &  x356 &  x371 &  x374 &  x383 &  x386 &  x389 &  x398 &  x401 &  x407 &  x425 &  x428 &  x434 &  x437 &  x446 &  x449 &  x455 &  x458 &  x464 &  x467 &  x476 &  x479 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x539 &  x545 &  x551 &  x557 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x587 &  x590 &  x593 &  x599 &  x602 &  x608 &  x617 &  x620 &  x623 &  x626 &  x632 &  x635 &  x647 &  x650 &  x665 &  x671 &  x674 &  x680 &  x692 &  x698 &  x701 &  x704 &  x710 &  x713 &  x719 &  x725 &  x737 &  x740 &  x758 &  x761 &  x773 &  x779 &  x782 &  x785 &  x791 &  x794 &  x797 &  x800 &  x809 &  x812 &  x815 &  x818 &  x833 &  x839 &  x845 &  x851 &  x854 &  x857 &  x860 &  x871 &  x875 &  x878 &  x884 &  x887 &  x893 &  x896 &  x899 &  x902 &  x905 &  x914 &  x917 &  x920 &  x923 &  x929 &  x935 &  x938 &  x941 &  x950 &  x953 &  x959 &  x962 &  x965 &  x968 &  x983 &  x986 &  x995 &  x1007 &  x1016 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1049 &  x1055 &  x1058 &  x1061 &  x1064 &  x1070 &  x1076 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130 & ~x51 & ~x90 & ~x336 & ~x570 & ~x609 & ~x822 & ~x861 & ~x978 & ~x1056 & ~x1057 & ~x1095;
assign c4194 =  x2 &  x8 &  x11 &  x20 &  x23 &  x29 &  x32 &  x43 &  x44 &  x47 &  x50 &  x59 &  x65 &  x68 &  x77 &  x82 &  x89 &  x98 &  x104 &  x107 &  x119 &  x121 &  x122 &  x125 &  x134 &  x140 &  x143 &  x146 &  x149 &  x155 &  x157 &  x158 &  x160 &  x161 &  x164 &  x167 &  x170 &  x173 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x235 &  x236 &  x245 &  x254 &  x257 &  x266 &  x269 &  x272 &  x274 &  x275 &  x281 &  x284 &  x290 &  x293 &  x299 &  x305 &  x308 &  x311 &  x314 &  x317 &  x338 &  x341 &  x347 &  x359 &  x365 &  x368 &  x371 &  x374 &  x377 &  x389 &  x398 &  x401 &  x410 &  x413 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x445 &  x452 &  x455 &  x464 &  x470 &  x473 &  x479 &  x484 &  x488 &  x491 &  x494 &  x500 &  x503 &  x512 &  x518 &  x521 &  x530 &  x533 &  x536 &  x539 &  x545 &  x548 &  x551 &  x557 &  x560 &  x563 &  x566 &  x572 &  x575 &  x584 &  x587 &  x593 &  x596 &  x599 &  x601 &  x602 &  x605 &  x608 &  x617 &  x620 &  x623 &  x629 &  x635 &  x638 &  x640 &  x641 &  x644 &  x655 &  x656 &  x659 &  x662 &  x665 &  x674 &  x677 &  x679 &  x683 &  x686 &  x698 &  x704 &  x707 &  x710 &  x713 &  x718 &  x719 &  x728 &  x733 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x754 &  x758 &  x767 &  x773 &  x785 &  x797 &  x800 &  x809 &  x811 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x835 &  x836 &  x839 &  x845 &  x850 &  x851 &  x857 &  x860 &  x866 &  x869 &  x875 &  x878 &  x881 &  x884 &  x887 &  x893 &  x896 &  x899 &  x902 &  x910 &  x911 &  x914 &  x920 &  x929 &  x932 &  x935 &  x938 &  x941 &  x947 &  x955 &  x956 &  x959 &  x962 &  x965 &  x971 &  x974 &  x989 &  x992 &  x1001 &  x1007 &  x1010 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1039 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x705 & ~x741 & ~x780 & ~x783 & ~x1014;
assign c4196 =  x2 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x50 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x107 &  x110 &  x113 &  x119 &  x122 &  x134 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x298 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x326 &  x329 &  x332 &  x335 &  x337 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x407 &  x413 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x572 &  x578 &  x581 &  x584 &  x587 &  x593 &  x599 &  x602 &  x605 &  x608 &  x611 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x641 &  x644 &  x647 &  x653 &  x656 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1054 &  x1055 &  x1058 &  x1064 &  x1067 &  x1069 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1108 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 & ~x21 & ~x60 & ~x360 & ~x399 & ~x423 & ~x438 & ~x477;
assign c4198 =  x2 &  x5 &  x14 &  x17 &  x20 &  x26 &  x38 &  x41 &  x43 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x71 &  x74 &  x79 &  x80 &  x82 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x113 &  x116 &  x118 &  x119 &  x121 &  x122 &  x125 &  x128 &  x131 &  x134 &  x140 &  x143 &  x146 &  x149 &  x152 &  x160 &  x161 &  x164 &  x170 &  x173 &  x176 &  x182 &  x185 &  x191 &  x194 &  x199 &  x203 &  x206 &  x215 &  x218 &  x221 &  x227 &  x235 &  x236 &  x238 &  x239 &  x245 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x314 &  x317 &  x320 &  x323 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x368 &  x371 &  x374 &  x383 &  x386 &  x389 &  x395 &  x398 &  x401 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x434 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x473 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x503 &  x506 &  x515 &  x518 &  x521 &  x523 &  x527 &  x533 &  x536 &  x545 &  x548 &  x554 &  x560 &  x562 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x593 &  x596 &  x602 &  x605 &  x608 &  x614 &  x620 &  x626 &  x632 &  x635 &  x638 &  x640 &  x644 &  x647 &  x653 &  x659 &  x662 &  x665 &  x671 &  x677 &  x686 &  x689 &  x695 &  x698 &  x704 &  x710 &  x713 &  x716 &  x718 &  x719 &  x722 &  x725 &  x731 &  x734 &  x740 &  x743 &  x746 &  x749 &  x752 &  x757 &  x758 &  x761 &  x764 &  x770 &  x773 &  x776 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x863 &  x866 &  x872 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x920 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1051 &  x1052 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1082 &  x1088 &  x1091 &  x1094 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 &  x1130 & ~x90 & ~x387 & ~x426 & ~x465 & ~x549;
assign c4200 =  x2 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x35 &  x38 &  x44 &  x47 &  x50 &  x53 &  x65 &  x68 &  x71 &  x80 &  x86 &  x89 &  x92 &  x101 &  x104 &  x107 &  x116 &  x119 &  x122 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x161 &  x164 &  x173 &  x179 &  x188 &  x191 &  x197 &  x200 &  x206 &  x209 &  x212 &  x218 &  x224 &  x227 &  x230 &  x233 &  x239 &  x242 &  x245 &  x248 &  x254 &  x257 &  x260 &  x266 &  x269 &  x272 &  x275 &  x284 &  x287 &  x299 &  x308 &  x311 &  x320 &  x326 &  x329 &  x332 &  x335 &  x338 &  x350 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x410 &  x413 &  x416 &  x425 &  x437 &  x443 &  x452 &  x458 &  x467 &  x473 &  x479 &  x482 &  x488 &  x494 &  x497 &  x503 &  x506 &  x515 &  x518 &  x521 &  x524 &  x527 &  x536 &  x539 &  x542 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x593 &  x608 &  x611 &  x614 &  x629 &  x632 &  x635 &  x641 &  x644 &  x650 &  x656 &  x659 &  x665 &  x674 &  x677 &  x686 &  x692 &  x695 &  x698 &  x701 &  x704 &  x716 &  x719 &  x722 &  x728 &  x734 &  x746 &  x749 &  x752 &  x758 &  x761 &  x767 &  x779 &  x788 &  x791 &  x797 &  x806 &  x809 &  x812 &  x815 &  x824 &  x827 &  x833 &  x839 &  x842 &  x845 &  x848 &  x854 &  x860 &  x869 &  x881 &  x884 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x914 &  x920 &  x923 &  x932 &  x935 &  x944 &  x947 &  x950 &  x956 &  x959 &  x968 &  x977 &  x980 &  x983 &  x989 &  x992 &  x995 &  x1001 &  x1007 &  x1013 &  x1016 &  x1025 &  x1028 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1127 &  x1130 & ~x105 & ~x183 & ~x255 & ~x339 & ~x351 & ~x378 & ~x390 & ~x423 & ~x429 & ~x462 & ~x468 & ~x469 & ~x501 & ~x735 & ~x768 & ~x774 & ~x801 & ~x807 & ~x813 & ~x846 & ~x1002 & ~x1074 & ~x1113;
assign c4202 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x241 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x355 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x393 &  x394 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x430 &  x431 &  x433 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x469 &  x470 &  x472 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x508 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x637 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x675 &  x676 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x715 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x399 & ~x513 & ~x552 & ~x591;
assign c4204 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x62 &  x65 &  x68 &  x71 &  x77 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x119 &  x122 &  x125 &  x128 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x238 &  x239 &  x242 &  x245 &  x248 &  x254 &  x257 &  x263 &  x266 &  x269 &  x275 &  x277 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x315 &  x316 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x355 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x383 &  x386 &  x389 &  x392 &  x394 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x433 &  x434 &  x437 &  x440 &  x443 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x569 &  x575 &  x578 &  x581 &  x584 &  x590 &  x596 &  x599 &  x602 &  x608 &  x614 &  x620 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x716 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x845 &  x848 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x962 &  x965 &  x968 &  x971 &  x974 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x117 & ~x255 & ~x282 & ~x705 & ~x783 & ~x822 & ~x861;
assign c4206 =  x2 &  x11 &  x20 &  x23 &  x26 &  x32 &  x35 &  x38 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x122 &  x125 &  x128 &  x131 &  x140 &  x149 &  x152 &  x161 &  x167 &  x170 &  x173 &  x176 &  x182 &  x185 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x224 &  x227 &  x233 &  x239 &  x242 &  x245 &  x248 &  x254 &  x257 &  x263 &  x266 &  x269 &  x272 &  x278 &  x281 &  x284 &  x287 &  x290 &  x292 &  x293 &  x296 &  x299 &  x302 &  x305 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x331 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x359 &  x362 &  x365 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x398 &  x401 &  x404 &  x407 &  x410 &  x416 &  x422 &  x425 &  x434 &  x437 &  x440 &  x443 &  x449 &  x455 &  x458 &  x461 &  x470 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x506 &  x509 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x545 &  x551 &  x554 &  x557 &  x563 &  x569 &  x572 &  x578 &  x581 &  x584 &  x590 &  x593 &  x596 &  x608 &  x614 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x662 &  x665 &  x671 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x728 &  x731 &  x734 &  x740 &  x743 &  x752 &  x755 &  x758 &  x761 &  x770 &  x776 &  x779 &  x785 &  x791 &  x794 &  x797 &  x800 &  x809 &  x812 &  x815 &  x818 &  x821 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x857 &  x863 &  x866 &  x869 &  x872 &  x878 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x932 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1016 &  x1019 &  x1022 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1106 &  x1109 &  x1115 &  x1121 &  x1124 &  x1127 & ~x54 & ~x93 & ~x132 & ~x171 & ~x189 & ~x210 & ~x228 & ~x282 & ~x321 & ~x450 & ~x534 & ~x723 & ~x1008;
assign c4208 =  x44 &  x68 &  x170 &  x218 &  x266 &  x281 &  x353 &  x359 &  x413 &  x419 &  x455 &  x488 &  x491 &  x494 &  x521 &  x569 &  x578 &  x584 &  x716 &  x821 &  x823 &  x827 &  x833 &  x842 &  x851 &  x1067 &  x1073 &  x1079 &  x1103 & ~x864 & ~x889 & ~x918 & ~x981;
assign c4210 =  x5 &  x8 &  x14 &  x17 &  x20 &  x35 &  x44 &  x47 &  x50 &  x56 &  x59 &  x68 &  x74 &  x77 &  x80 &  x83 &  x92 &  x95 &  x98 &  x101 &  x110 &  x113 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x155 &  x167 &  x170 &  x173 &  x176 &  x179 &  x191 &  x206 &  x209 &  x221 &  x227 &  x230 &  x233 &  x236 &  x239 &  x251 &  x254 &  x260 &  x263 &  x272 &  x275 &  x278 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x316 &  x320 &  x323 &  x326 &  x329 &  x335 &  x341 &  x350 &  x352 &  x353 &  x355 &  x356 &  x359 &  x362 &  x365 &  x374 &  x377 &  x380 &  x383 &  x386 &  x391 &  x398 &  x401 &  x410 &  x425 &  x431 &  x440 &  x443 &  x446 &  x449 &  x452 &  x467 &  x470 &  x476 &  x479 &  x491 &  x494 &  x500 &  x503 &  x509 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x542 &  x545 &  x554 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x584 &  x587 &  x593 &  x595 &  x599 &  x602 &  x605 &  x614 &  x617 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x656 &  x659 &  x673 &  x674 &  x677 &  x679 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x712 &  x713 &  x716 &  x718 &  x722 &  x725 &  x746 &  x755 &  x758 &  x761 &  x764 &  x770 &  x773 &  x776 &  x785 &  x791 &  x794 &  x797 &  x800 &  x806 &  x812 &  x815 &  x821 &  x824 &  x830 &  x836 &  x839 &  x842 &  x848 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x881 &  x887 &  x890 &  x899 &  x902 &  x911 &  x914 &  x917 &  x926 &  x932 &  x938 &  x941 &  x950 &  x953 &  x965 &  x968 &  x971 &  x974 &  x980 &  x989 &  x995 &  x1004 &  x1013 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1061 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1103 &  x1109 &  x1112 &  x1124 &  x1130 & ~x93 & ~x165 & ~x435 & ~x705;
assign c4212 =  x5 &  x11 &  x14 &  x20 &  x23 &  x29 &  x32 &  x41 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x71 &  x74 &  x77 &  x83 &  x86 &  x92 &  x95 &  x101 &  x107 &  x110 &  x116 &  x119 &  x125 &  x128 &  x131 &  x134 &  x140 &  x143 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x242 &  x245 &  x251 &  x254 &  x260 &  x263 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x296 &  x302 &  x305 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x362 &  x371 &  x377 &  x383 &  x386 &  x392 &  x395 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x425 &  x431 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x458 &  x461 &  x464 &  x467 &  x473 &  x476 &  x482 &  x488 &  x491 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x542 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x605 &  x611 &  x614 &  x617 &  x620 &  x623 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x656 &  x659 &  x662 &  x665 &  x671 &  x674 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x704 &  x710 &  x713 &  x716 &  x719 &  x722 &  x728 &  x737 &  x743 &  x746 &  x749 &  x752 &  x758 &  x764 &  x770 &  x773 &  x776 &  x782 &  x785 &  x791 &  x794 &  x797 &  x800 &  x809 &  x815 &  x818 &  x821 &  x824 &  x827 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x893 &  x896 &  x902 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x977 &  x980 &  x989 &  x995 &  x1001 &  x1007 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1049 &  x1064 &  x1067 &  x1073 &  x1076 &  x1082 &  x1088 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1118 &  x1121 &  x1124 &  x1130 & ~x33 & ~x51 & ~x318 & ~x357 & ~x549 & ~x589 & ~x666 & ~x801 & ~x852 & ~x891 & ~x930 & ~x1002 & ~x1008;
assign c4214 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x50 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x164 &  x167 &  x170 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x263 &  x269 &  x280 &  x281 &  x284 &  x287 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x356 &  x359 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x419 &  x422 &  x425 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x472 &  x473 &  x476 &  x479 &  x485 &  x488 &  x491 &  x494 &  x497 &  x503 &  x506 &  x509 &  x511 &  x512 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x542 &  x548 &  x551 &  x554 &  x557 &  x566 &  x569 &  x575 &  x581 &  x584 &  x586 &  x587 &  x593 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x625 &  x632 &  x635 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x664 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x754 &  x755 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x815 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x854 &  x857 &  x860 &  x863 &  x866 &  x867 &  x869 &  x875 &  x878 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x929 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x989 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1061 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1130 & ~x786 & ~x825;
assign c4216 =  x4 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x53 &  x65 &  x80 &  x83 &  x92 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x122 &  x125 &  x128 &  x131 &  x134 &  x136 &  x137 &  x143 &  x146 &  x149 &  x161 &  x167 &  x170 &  x175 &  x179 &  x185 &  x191 &  x194 &  x206 &  x212 &  x221 &  x224 &  x227 &  x239 &  x242 &  x245 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x271 &  x278 &  x281 &  x284 &  x287 &  x299 &  x302 &  x317 &  x320 &  x326 &  x338 &  x341 &  x347 &  x350 &  x356 &  x362 &  x368 &  x371 &  x380 &  x392 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x431 &  x433 &  x434 &  x440 &  x443 &  x449 &  x452 &  x461 &  x467 &  x476 &  x479 &  x485 &  x494 &  x497 &  x500 &  x509 &  x511 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x548 &  x550 &  x560 &  x563 &  x575 &  x581 &  x584 &  x589 &  x596 &  x599 &  x602 &  x604 &  x605 &  x614 &  x617 &  x620 &  x626 &  x629 &  x632 &  x635 &  x641 &  x647 &  x650 &  x656 &  x659 &  x665 &  x668 &  x671 &  x680 &  x683 &  x695 &  x704 &  x707 &  x713 &  x716 &  x719 &  x725 &  x727 &  x728 &  x734 &  x740 &  x743 &  x746 &  x752 &  x755 &  x757 &  x758 &  x767 &  x770 &  x776 &  x788 &  x800 &  x812 &  x815 &  x818 &  x821 &  x827 &  x830 &  x833 &  x842 &  x845 &  x854 &  x863 &  x866 &  x874 &  x875 &  x884 &  x887 &  x896 &  x899 &  x902 &  x905 &  x908 &  x914 &  x917 &  x920 &  x929 &  x932 &  x938 &  x941 &  x944 &  x947 &  x955 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x986 &  x989 &  x998 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1040 &  x1052 &  x1058 &  x1064 &  x1067 &  x1070 &  x1085 &  x1094 &  x1097 &  x1100 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124;
assign c4218 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x238 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x276 &  x277 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x316 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x355 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x391 &  x392 &  x394 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x433 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x469 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x556 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x595 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x150 & ~x189 & ~x435 & ~x474 & ~x513 & ~x552 & ~x591 & ~x705 & ~x744 & ~x783 & ~x822;
assign c4220 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x194 &  x197 &  x199 &  x203 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x235 &  x236 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x274 &  x275 &  x277 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x314 &  x317 &  x320 &  x323 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x391 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x481 &  x482 &  x485 &  x488 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x718 &  x719 &  x722 &  x725 &  x728 &  x731 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x757 &  x758 &  x761 &  x764 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x796 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x959 &  x962 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x318 & ~x357 & ~x501 & ~x549 & ~x588 & ~x627 & ~x666 & ~x705 & ~x744 & ~x783 & ~x822 & ~x861 & ~x897 & ~x975 & ~x1014;
assign c4222 =  x2 &  x26 &  x38 &  x44 &  x50 &  x56 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x95 &  x98 &  x101 &  x122 &  x131 &  x134 &  x137 &  x140 &  x155 &  x158 &  x164 &  x170 &  x176 &  x179 &  x191 &  x194 &  x197 &  x200 &  x202 &  x203 &  x209 &  x218 &  x224 &  x227 &  x233 &  x239 &  x241 &  x242 &  x245 &  x251 &  x272 &  x275 &  x284 &  x293 &  x299 &  x302 &  x314 &  x317 &  x320 &  x323 &  x326 &  x338 &  x341 &  x347 &  x350 &  x353 &  x362 &  x368 &  x374 &  x383 &  x386 &  x389 &  x392 &  x395 &  x413 &  x419 &  x422 &  x443 &  x455 &  x458 &  x482 &  x485 &  x491 &  x500 &  x518 &  x521 &  x539 &  x542 &  x554 &  x563 &  x566 &  x575 &  x578 &  x587 &  x608 &  x611 &  x617 &  x620 &  x638 &  x641 &  x647 &  x664 &  x665 &  x674 &  x689 &  x692 &  x695 &  x716 &  x719 &  x722 &  x737 &  x746 &  x755 &  x758 &  x761 &  x764 &  x773 &  x782 &  x803 &  x815 &  x818 &  x821 &  x835 &  x842 &  x848 &  x857 &  x860 &  x863 &  x866 &  x869 &  x890 &  x893 &  x896 &  x905 &  x920 &  x926 &  x941 &  x944 &  x947 &  x950 &  x953 &  x959 &  x965 &  x968 &  x974 &  x977 &  x986 &  x995 &  x1013 &  x1019 &  x1022 &  x1037 &  x1049 &  x1052 &  x1058 &  x1064 &  x1067 &  x1082 &  x1091 &  x1097 &  x1100 &  x1115 &  x1130 & ~x669 & ~x894 & ~x978 & ~x1044 & ~x1056 & ~x1071;
assign c4224 =  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x121 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x146 &  x149 &  x152 &  x157 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x196 &  x197 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x227 &  x233 &  x235 &  x236 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x308 &  x311 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x523 &  x524 &  x527 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x566 &  x569 &  x572 &  x578 &  x584 &  x590 &  x593 &  x596 &  x601 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x626 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x656 &  x659 &  x662 &  x665 &  x668 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x757 &  x758 &  x761 &  x764 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x839 &  x845 &  x851 &  x854 &  x857 &  x863 &  x866 &  x869 &  x871 &  x872 &  x875 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x920 &  x923 &  x926 &  x932 &  x935 &  x941 &  x944 &  x950 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x995 &  x998 &  x1001 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 &  x1130 & ~x279 & ~x318 & ~x357 & ~x501 & ~x780 & ~x819 & ~x939 & ~x978 & ~x1014 & ~x1017 & ~x1053 & ~x1056;
assign c4226 =  x5 &  x41 &  x74 &  x86 &  x104 &  x107 &  x122 &  x128 &  x137 &  x164 &  x182 &  x194 &  x227 &  x239 &  x242 &  x245 &  x251 &  x269 &  x272 &  x278 &  x296 &  x308 &  x326 &  x329 &  x332 &  x335 &  x341 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x389 &  x401 &  x416 &  x428 &  x440 &  x452 &  x458 &  x464 &  x467 &  x473 &  x482 &  x488 &  x491 &  x494 &  x497 &  x512 &  x515 &  x548 &  x557 &  x563 &  x566 &  x575 &  x581 &  x584 &  x590 &  x593 &  x596 &  x611 &  x620 &  x641 &  x647 &  x665 &  x671 &  x677 &  x680 &  x689 &  x692 &  x728 &  x742 &  x743 &  x752 &  x764 &  x767 &  x773 &  x776 &  x782 &  x788 &  x797 &  x806 &  x812 &  x815 &  x818 &  x824 &  x830 &  x839 &  x845 &  x848 &  x851 &  x854 &  x866 &  x869 &  x887 &  x902 &  x905 &  x914 &  x917 &  x920 &  x935 &  x941 &  x944 &  x946 &  x947 &  x950 &  x998 &  x1004 &  x1025 &  x1028 &  x1030 &  x1046 &  x1049 &  x1055 &  x1067 &  x1070 &  x1073 &  x1097 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1130 & ~x81 & ~x399 & ~x894 & ~x933 & ~x966 & ~x972 & ~x1044 & ~x1056;
assign c4228 =  x2 &  x5 &  x8 &  x11 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x44 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x395 &  x398 &  x401 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x508 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x835 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x249 & ~x267 & ~x462 & ~x501 & ~x591 & ~x783 & ~x822 & ~x852 & ~x861;
assign c4230 =  x4 &  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x29 &  x32 &  x35 &  x41 &  x42 &  x43 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x79 &  x80 &  x81 &  x82 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x121 &  x122 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x157 &  x160 &  x161 &  x164 &  x167 &  x170 &  x173 &  x179 &  x185 &  x188 &  x191 &  x194 &  x196 &  x197 &  x199 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x281 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x323 &  x326 &  x329 &  x332 &  x338 &  x341 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x551 &  x554 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x605 &  x608 &  x611 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x665 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x718 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x743 &  x746 &  x749 &  x757 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x973 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1067 &  x1070 &  x1073 &  x1076 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x147 & ~x387 & ~x669;
assign c4232 =  x2 &  x5 &  x8 &  x11 &  x17 &  x29 &  x38 &  x41 &  x47 &  x53 &  x65 &  x68 &  x71 &  x77 &  x83 &  x89 &  x98 &  x110 &  x116 &  x119 &  x122 &  x125 &  x128 &  x137 &  x140 &  x146 &  x149 &  x155 &  x167 &  x173 &  x185 &  x188 &  x197 &  x203 &  x206 &  x209 &  x224 &  x233 &  x239 &  x245 &  x248 &  x251 &  x254 &  x257 &  x269 &  x272 &  x275 &  x281 &  x284 &  x287 &  x290 &  x305 &  x308 &  x311 &  x314 &  x317 &  x323 &  x338 &  x344 &  x347 &  x350 &  x357 &  x362 &  x368 &  x371 &  x377 &  x383 &  x389 &  x392 &  x401 &  x404 &  x413 &  x422 &  x437 &  x443 &  x449 &  x458 &  x461 &  x464 &  x467 &  x470 &  x471 &  x472 &  x473 &  x476 &  x479 &  x482 &  x485 &  x494 &  x510 &  x512 &  x515 &  x521 &  x524 &  x527 &  x536 &  x550 &  x557 &  x560 &  x563 &  x566 &  x569 &  x578 &  x581 &  x584 &  x587 &  x589 &  x599 &  x608 &  x614 &  x617 &  x623 &  x629 &  x638 &  x647 &  x659 &  x662 &  x665 &  x671 &  x674 &  x677 &  x680 &  x689 &  x698 &  x707 &  x722 &  x725 &  x731 &  x734 &  x740 &  x746 &  x758 &  x764 &  x767 &  x770 &  x773 &  x797 &  x800 &  x809 &  x818 &  x821 &  x827 &  x830 &  x836 &  x839 &  x845 &  x848 &  x854 &  x860 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x899 &  x905 &  x917 &  x929 &  x932 &  x947 &  x950 &  x953 &  x956 &  x962 &  x965 &  x977 &  x983 &  x986 &  x998 &  x1001 &  x1004 &  x1010 &  x1022 &  x1025 &  x1034 &  x1037 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1082 &  x1091 &  x1094 &  x1097 &  x1100 &  x1109 &  x1112 &  x1118 &  x1124 &  x1130 & ~x273 & ~x312 & ~x477;
assign c4234 =  x2 &  x5 &  x14 &  x20 &  x26 &  x32 &  x38 &  x47 &  x56 &  x59 &  x62 &  x65 &  x80 &  x83 &  x86 &  x89 &  x92 &  x101 &  x107 &  x119 &  x128 &  x137 &  x140 &  x146 &  x149 &  x152 &  x155 &  x158 &  x164 &  x167 &  x173 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x212 &  x215 &  x224 &  x227 &  x230 &  x236 &  x245 &  x254 &  x257 &  x263 &  x266 &  x269 &  x275 &  x278 &  x281 &  x287 &  x293 &  x298 &  x302 &  x305 &  x308 &  x311 &  x317 &  x320 &  x323 &  x329 &  x332 &  x341 &  x344 &  x350 &  x353 &  x356 &  x359 &  x368 &  x380 &  x383 &  x395 &  x401 &  x404 &  x407 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x446 &  x452 &  x455 &  x461 &  x473 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x503 &  x509 &  x515 &  x518 &  x521 &  x527 &  x530 &  x539 &  x542 &  x548 &  x554 &  x560 &  x563 &  x569 &  x572 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x620 &  x623 &  x638 &  x641 &  x647 &  x653 &  x656 &  x659 &  x664 &  x665 &  x674 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x703 &  x704 &  x719 &  x722 &  x725 &  x731 &  x737 &  x740 &  x743 &  x749 &  x752 &  x755 &  x761 &  x767 &  x782 &  x788 &  x794 &  x797 &  x806 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x848 &  x851 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x890 &  x899 &  x911 &  x914 &  x917 &  x920 &  x926 &  x932 &  x938 &  x947 &  x950 &  x953 &  x956 &  x959 &  x965 &  x968 &  x971 &  x977 &  x980 &  x989 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1040 &  x1049 &  x1055 &  x1061 &  x1064 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x273 & ~x312 & ~x351 & ~x429 & ~x468 & ~x507 & ~x594 & ~x633 & ~x747 & ~x1017;
assign c4236 =  x20 &  x47 &  x65 &  x79 &  x92 &  x101 &  x134 &  x152 &  x164 &  x182 &  x194 &  x197 &  x218 &  x236 &  x242 &  x269 &  x289 &  x290 &  x311 &  x320 &  x335 &  x350 &  x367 &  x371 &  x383 &  x401 &  x419 &  x424 &  x428 &  x431 &  x448 &  x455 &  x458 &  x461 &  x473 &  x494 &  x530 &  x533 &  x545 &  x554 &  x560 &  x566 &  x593 &  x656 &  x677 &  x716 &  x725 &  x749 &  x791 &  x818 &  x820 &  x824 &  x830 &  x833 &  x860 &  x866 &  x881 &  x898 &  x902 &  x917 &  x920 &  x953 &  x959 &  x962 &  x986 &  x1001 &  x1010 &  x1034 &  x1037 &  x1054 &  x1061 &  x1079 &  x1094 &  x1097 &  x1106 &  x1108 & ~x1059 & ~x1071 & ~x1110;
assign c4238 =  x2 &  x11 &  x14 &  x17 &  x20 &  x23 &  x29 &  x38 &  x41 &  x44 &  x59 &  x62 &  x71 &  x74 &  x83 &  x86 &  x92 &  x101 &  x107 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x146 &  x152 &  x158 &  x170 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x251 &  x254 &  x257 &  x263 &  x266 &  x269 &  x272 &  x278 &  x281 &  x284 &  x290 &  x293 &  x296 &  x304 &  x308 &  x311 &  x314 &  x320 &  x323 &  x326 &  x329 &  x332 &  x337 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x371 &  x374 &  x377 &  x383 &  x386 &  x389 &  x392 &  x395 &  x404 &  x407 &  x410 &  x419 &  x422 &  x428 &  x431 &  x434 &  x437 &  x440 &  x446 &  x449 &  x455 &  x461 &  x464 &  x467 &  x473 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x503 &  x509 &  x518 &  x527 &  x530 &  x536 &  x538 &  x539 &  x545 &  x551 &  x554 &  x560 &  x575 &  x578 &  x581 &  x587 &  x590 &  x593 &  x599 &  x602 &  x605 &  x608 &  x611 &  x617 &  x620 &  x635 &  x638 &  x644 &  x647 &  x650 &  x653 &  x664 &  x665 &  x668 &  x671 &  x674 &  x683 &  x686 &  x692 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x731 &  x737 &  x743 &  x746 &  x752 &  x755 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x860 &  x863 &  x866 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x896 &  x905 &  x907 &  x908 &  x910 &  x911 &  x914 &  x917 &  x920 &  x926 &  x935 &  x941 &  x944 &  x947 &  x949 &  x952 &  x953 &  x959 &  x962 &  x965 &  x974 &  x977 &  x983 &  x986 &  x992 &  x995 &  x1004 &  x1016 &  x1025 &  x1028 &  x1031 &  x1040 &  x1043 &  x1046 &  x1055 &  x1058 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x1056 & ~x1095;
assign c4240 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x280 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x316 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x355 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x433 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x506 &  x508 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x547 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x611 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x363 & ~x399 & ~x402 & ~x438 & ~x576 & ~x615;
assign c4242 =  x2 &  x5 &  x11 &  x17 &  x20 &  x23 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x89 &  x92 &  x95 &  x104 &  x110 &  x113 &  x122 &  x128 &  x137 &  x140 &  x143 &  x164 &  x167 &  x170 &  x185 &  x194 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x227 &  x233 &  x236 &  x242 &  x245 &  x248 &  x254 &  x257 &  x260 &  x263 &  x269 &  x272 &  x275 &  x281 &  x284 &  x290 &  x293 &  x299 &  x305 &  x314 &  x323 &  x326 &  x332 &  x338 &  x344 &  x353 &  x359 &  x362 &  x365 &  x371 &  x374 &  x383 &  x386 &  x389 &  x392 &  x398 &  x401 &  x407 &  x410 &  x416 &  x422 &  x425 &  x428 &  x431 &  x437 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x470 &  x473 &  x482 &  x494 &  x506 &  x515 &  x521 &  x524 &  x533 &  x557 &  x563 &  x572 &  x578 &  x581 &  x587 &  x590 &  x593 &  x596 &  x602 &  x608 &  x611 &  x623 &  x626 &  x629 &  x647 &  x653 &  x656 &  x659 &  x665 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x704 &  x707 &  x710 &  x719 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x776 &  x782 &  x785 &  x791 &  x794 &  x797 &  x800 &  x803 &  x809 &  x812 &  x818 &  x821 &  x824 &  x830 &  x833 &  x836 &  x845 &  x848 &  x854 &  x860 &  x866 &  x875 &  x881 &  x884 &  x896 &  x902 &  x911 &  x917 &  x923 &  x926 &  x932 &  x944 &  x947 &  x950 &  x956 &  x959 &  x962 &  x980 &  x983 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1013 &  x1016 &  x1019 &  x1028 &  x1034 &  x1040 &  x1043 &  x1046 &  x1055 &  x1058 &  x1067 &  x1070 &  x1076 &  x1085 &  x1091 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x273 & ~x288 & ~x327 & ~x528 & ~x546 & ~x735 & ~x736 & ~x774 & ~x807 & ~x963 & ~x966 & ~x1005;
assign c4244 =  x2 &  x8 &  x17 &  x20 &  x23 &  x29 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x59 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x89 &  x95 &  x107 &  x110 &  x113 &  x116 &  x122 &  x128 &  x131 &  x134 &  x137 &  x143 &  x149 &  x152 &  x158 &  x167 &  x170 &  x173 &  x176 &  x182 &  x185 &  x188 &  x194 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x227 &  x233 &  x236 &  x242 &  x245 &  x254 &  x263 &  x278 &  x284 &  x293 &  x296 &  x302 &  x311 &  x314 &  x320 &  x323 &  x326 &  x329 &  x335 &  x338 &  x344 &  x356 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x404 &  x407 &  x410 &  x416 &  x422 &  x425 &  x428 &  x431 &  x433 &  x434 &  x437 &  x440 &  x443 &  x452 &  x458 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x494 &  x500 &  x503 &  x506 &  x509 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x542 &  x545 &  x547 &  x548 &  x551 &  x557 &  x560 &  x575 &  x584 &  x590 &  x593 &  x599 &  x602 &  x605 &  x608 &  x614 &  x620 &  x623 &  x626 &  x629 &  x634 &  x635 &  x637 &  x638 &  x647 &  x656 &  x662 &  x665 &  x668 &  x671 &  x674 &  x676 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x722 &  x728 &  x731 &  x734 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x761 &  x779 &  x782 &  x785 &  x791 &  x797 &  x800 &  x806 &  x812 &  x830 &  x833 &  x839 &  x845 &  x851 &  x857 &  x860 &  x863 &  x866 &  x869 &  x875 &  x878 &  x881 &  x884 &  x887 &  x893 &  x902 &  x908 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x962 &  x965 &  x968 &  x974 &  x980 &  x986 &  x989 &  x992 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1019 &  x1025 &  x1028 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1070 &  x1082 &  x1088 &  x1091 &  x1094 &  x1100 &  x1103 &  x1121 &  x1124 &  x1130 & ~x399 & ~x513 & ~x552 & ~x553 & ~x591 & ~x630 & ~x822;
assign c4246 =  x11 &  x17 &  x23 &  x38 &  x41 &  x44 &  x62 &  x65 &  x68 &  x74 &  x77 &  x80 &  x89 &  x95 &  x110 &  x116 &  x134 &  x140 &  x152 &  x155 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x188 &  x194 &  x199 &  x209 &  x215 &  x218 &  x221 &  x224 &  x233 &  x236 &  x238 &  x239 &  x242 &  x245 &  x251 &  x257 &  x269 &  x272 &  x275 &  x278 &  x284 &  x290 &  x293 &  x296 &  x302 &  x305 &  x308 &  x311 &  x314 &  x320 &  x323 &  x338 &  x347 &  x350 &  x356 &  x359 &  x362 &  x368 &  x371 &  x377 &  x383 &  x386 &  x389 &  x398 &  x410 &  x419 &  x428 &  x434 &  x437 &  x443 &  x446 &  x455 &  x470 &  x473 &  x485 &  x488 &  x494 &  x497 &  x500 &  x503 &  x512 &  x515 &  x523 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x548 &  x554 &  x557 &  x560 &  x563 &  x569 &  x575 &  x578 &  x581 &  x587 &  x595 &  x596 &  x599 &  x601 &  x605 &  x611 &  x617 &  x623 &  x626 &  x632 &  x641 &  x656 &  x659 &  x662 &  x668 &  x671 &  x677 &  x679 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x704 &  x707 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x755 &  x758 &  x761 &  x764 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x794 &  x800 &  x803 &  x809 &  x812 &  x818 &  x827 &  x830 &  x835 &  x838 &  x848 &  x851 &  x854 &  x857 &  x863 &  x866 &  x869 &  x875 &  x877 &  x878 &  x884 &  x893 &  x902 &  x905 &  x911 &  x914 &  x916 &  x917 &  x920 &  x923 &  x941 &  x947 &  x950 &  x959 &  x965 &  x968 &  x974 &  x980 &  x986 &  x989 &  x992 &  x998 &  x1000 &  x1004 &  x1012 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1039 &  x1046 &  x1052 &  x1058 &  x1064 &  x1076 &  x1078 &  x1082 &  x1085 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x210 & ~x357 & ~x396;
assign c4248 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x511 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x550 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x589 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x686 &  x689 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x718 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x399 & ~x438 & ~x477 & ~x708 & ~x723;
assign c4250 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x125 &  x128 &  x134 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x251 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x308 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x338 &  x341 &  x344 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x536 &  x542 &  x545 &  x554 &  x569 &  x572 &  x575 &  x578 &  x581 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x770 &  x773 &  x776 &  x779 &  x785 &  x788 &  x791 &  x794 &  x796 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x835 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 &  x1130 & ~x630 & ~x645 & ~x657 & ~x669 & ~x684 & ~x723 & ~x921 & ~x1056;
assign c4252 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x83 &  x86 &  x89 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x198 &  x199 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x235 &  x236 &  x237 &  x238 &  x239 &  x242 &  x245 &  x248 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x274 &  x275 &  x277 &  x278 &  x281 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x308 &  x311 &  x314 &  x316 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x391 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x455 &  x464 &  x467 &  x470 &  x473 &  x476 &  x478 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x503 &  x506 &  x512 &  x515 &  x518 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x204 & ~x318 & ~x319 & ~x357 & ~x358 & ~x396 & ~x435 & ~x436;
assign c4254 =  x2 &  x11 &  x14 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x44 &  x47 &  x50 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x92 &  x95 &  x98 &  x104 &  x107 &  x113 &  x119 &  x122 &  x125 &  x131 &  x140 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x185 &  x191 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x239 &  x241 &  x242 &  x245 &  x248 &  x251 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x299 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x433 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x508 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x542 &  x547 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x617 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x676 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x715 &  x716 &  x719 &  x722 &  x731 &  x737 &  x740 &  x743 &  x749 &  x752 &  x754 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x788 &  x791 &  x794 &  x797 &  x800 &  x806 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x833 &  x836 &  x842 &  x845 &  x848 &  x851 &  x857 &  x860 &  x863 &  x866 &  x869 &  x875 &  x878 &  x887 &  x890 &  x893 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1085 &  x1088 &  x1091 &  x1094 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x117 & ~x195 & ~x234 & ~x360 & ~x399 & ~x552 & ~x591 & ~x783 & ~x861;
assign c4256 =  x2 &  x11 &  x14 &  x17 &  x20 &  x23 &  x29 &  x35 &  x41 &  x44 &  x53 &  x56 &  x59 &  x62 &  x65 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x95 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x140 &  x143 &  x149 &  x152 &  x155 &  x158 &  x164 &  x167 &  x173 &  x176 &  x179 &  x182 &  x191 &  x194 &  x197 &  x199 &  x200 &  x209 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x237 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x260 &  x263 &  x269 &  x272 &  x275 &  x276 &  x277 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x314 &  x316 &  x317 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x352 &  x353 &  x355 &  x356 &  x359 &  x362 &  x368 &  x371 &  x374 &  x380 &  x383 &  x386 &  x389 &  x391 &  x392 &  x398 &  x401 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x446 &  x452 &  x458 &  x461 &  x464 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x556 &  x557 &  x560 &  x566 &  x569 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x595 &  x596 &  x601 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x634 &  x635 &  x638 &  x640 &  x641 &  x647 &  x650 &  x656 &  x659 &  x662 &  x665 &  x671 &  x674 &  x676 &  x679 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x718 &  x722 &  x725 &  x728 &  x731 &  x740 &  x743 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x782 &  x785 &  x788 &  x793 &  x794 &  x796 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x827 &  x830 &  x833 &  x835 &  x836 &  x839 &  x842 &  x848 &  x851 &  x854 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x941 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x992 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1067 &  x1073 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x396 & ~x435;
assign c4258 =  x2 &  x5 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x35 &  x38 &  x41 &  x47 &  x50 &  x53 &  x56 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x89 &  x92 &  x98 &  x104 &  x107 &  x110 &  x113 &  x116 &  x123 &  x124 &  x125 &  x128 &  x131 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x170 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x199 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x237 &  x248 &  x251 &  x254 &  x263 &  x266 &  x269 &  x272 &  x275 &  x276 &  x278 &  x287 &  x290 &  x302 &  x305 &  x308 &  x311 &  x314 &  x315 &  x316 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x347 &  x353 &  x355 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x383 &  x386 &  x389 &  x394 &  x395 &  x398 &  x401 &  x404 &  x407 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x479 &  x482 &  x485 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x530 &  x533 &  x536 &  x542 &  x548 &  x551 &  x554 &  x557 &  x560 &  x572 &  x578 &  x581 &  x584 &  x587 &  x590 &  x596 &  x599 &  x602 &  x605 &  x614 &  x617 &  x620 &  x623 &  x629 &  x632 &  x638 &  x641 &  x644 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x764 &  x767 &  x773 &  x779 &  x782 &  x785 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x845 &  x848 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x887 &  x890 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x962 &  x965 &  x968 &  x971 &  x977 &  x980 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1100 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x228 & ~x243 & ~x282;
assign c4260 =  x2 &  x5 &  x11 &  x14 &  x17 &  x23 &  x29 &  x32 &  x35 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x365 &  x368 &  x371 &  x374 &  x380 &  x383 &  x386 &  x389 &  x391 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x430 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x512 &  x515 &  x518 &  x521 &  x523 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x578 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x623 &  x626 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x715 &  x716 &  x718 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x757 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x796 &  x797 &  x800 &  x803 &  x806 &  x809 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x835 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x874 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1084 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1123 &  x1127 &  x1130 & ~x231 & ~x435 & ~x474 & ~x513 & ~x552 & ~x822 & ~x900;
assign c4262 =  x20 &  x23 &  x35 &  x41 &  x53 &  x62 &  x68 &  x92 &  x113 &  x119 &  x122 &  x137 &  x146 &  x167 &  x170 &  x173 &  x197 &  x203 &  x212 &  x251 &  x254 &  x260 &  x269 &  x278 &  x293 &  x308 &  x311 &  x317 &  x323 &  x353 &  x362 &  x386 &  x401 &  x404 &  x425 &  x434 &  x512 &  x524 &  x526 &  x530 &  x539 &  x545 &  x551 &  x554 &  x565 &  x572 &  x577 &  x584 &  x602 &  x611 &  x641 &  x647 &  x653 &  x683 &  x698 &  x701 &  x705 &  x706 &  x728 &  x734 &  x743 &  x749 &  x755 &  x761 &  x764 &  x788 &  x797 &  x800 &  x809 &  x812 &  x869 &  x890 &  x901 &  x905 &  x920 &  x947 &  x974 &  x983 &  x1046 &  x1055 &  x1061 &  x1073 &  x1076 &  x1085 &  x1127 &  x1130 & ~x312 & ~x429 & ~x468 & ~x507 & ~x585 & ~x942 & ~x943 & ~x981;
assign c4264 =  x2 &  x8 &  x14 &  x17 &  x20 &  x26 &  x29 &  x32 &  x41 &  x44 &  x53 &  x56 &  x59 &  x68 &  x71 &  x77 &  x80 &  x89 &  x92 &  x101 &  x104 &  x110 &  x113 &  x116 &  x122 &  x125 &  x131 &  x137 &  x140 &  x146 &  x149 &  x161 &  x164 &  x179 &  x182 &  x185 &  x188 &  x194 &  x200 &  x212 &  x215 &  x218 &  x227 &  x230 &  x248 &  x251 &  x254 &  x260 &  x266 &  x269 &  x272 &  x278 &  x284 &  x287 &  x296 &  x305 &  x311 &  x314 &  x317 &  x320 &  x326 &  x329 &  x335 &  x344 &  x353 &  x356 &  x362 &  x374 &  x380 &  x383 &  x386 &  x392 &  x395 &  x401 &  x413 &  x416 &  x425 &  x428 &  x434 &  x437 &  x443 &  x449 &  x452 &  x455 &  x464 &  x467 &  x473 &  x476 &  x479 &  x485 &  x488 &  x494 &  x497 &  x521 &  x524 &  x527 &  x530 &  x536 &  x545 &  x553 &  x554 &  x566 &  x590 &  x593 &  x599 &  x611 &  x614 &  x617 &  x620 &  x638 &  x641 &  x644 &  x662 &  x665 &  x668 &  x671 &  x674 &  x686 &  x706 &  x707 &  x710 &  x713 &  x719 &  x725 &  x728 &  x734 &  x737 &  x746 &  x749 &  x755 &  x758 &  x761 &  x767 &  x776 &  x785 &  x794 &  x800 &  x803 &  x806 &  x818 &  x820 &  x821 &  x823 &  x827 &  x833 &  x839 &  x848 &  x851 &  x854 &  x860 &  x862 &  x866 &  x869 &  x872 &  x875 &  x893 &  x896 &  x899 &  x901 &  x902 &  x905 &  x911 &  x917 &  x920 &  x929 &  x935 &  x938 &  x941 &  x950 &  x953 &  x956 &  x959 &  x971 &  x974 &  x980 &  x983 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1016 &  x1019 &  x1022 &  x1031 &  x1034 &  x1040 &  x1046 &  x1055 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1085 &  x1091 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 & ~x390 & ~x468 & ~x546 & ~x585 & ~x636 & ~x903 & ~x924;
assign c4266 =  x14 &  x17 &  x23 &  x26 &  x41 &  x44 &  x47 &  x53 &  x56 &  x65 &  x77 &  x80 &  x83 &  x95 &  x101 &  x107 &  x110 &  x113 &  x128 &  x131 &  x134 &  x140 &  x146 &  x155 &  x158 &  x167 &  x170 &  x173 &  x185 &  x206 &  x209 &  x212 &  x224 &  x236 &  x242 &  x254 &  x257 &  x260 &  x263 &  x266 &  x275 &  x287 &  x296 &  x302 &  x316 &  x320 &  x323 &  x326 &  x338 &  x341 &  x350 &  x359 &  x362 &  x368 &  x374 &  x377 &  x383 &  x386 &  x395 &  x398 &  x401 &  x407 &  x410 &  x428 &  x431 &  x433 &  x434 &  x437 &  x446 &  x449 &  x452 &  x455 &  x464 &  x467 &  x473 &  x494 &  x503 &  x508 &  x518 &  x530 &  x536 &  x545 &  x548 &  x554 &  x557 &  x560 &  x563 &  x569 &  x584 &  x587 &  x590 &  x593 &  x602 &  x617 &  x620 &  x623 &  x629 &  x635 &  x637 &  x644 &  x647 &  x671 &  x672 &  x674 &  x677 &  x707 &  x713 &  x722 &  x725 &  x731 &  x743 &  x749 &  x755 &  x758 &  x764 &  x767 &  x788 &  x791 &  x797 &  x800 &  x806 &  x824 &  x827 &  x833 &  x836 &  x839 &  x848 &  x851 &  x866 &  x869 &  x874 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x941 &  x947 &  x959 &  x965 &  x974 &  x977 &  x980 &  x986 &  x989 &  x1004 &  x1007 &  x1019 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1064 &  x1079 &  x1082 &  x1085 &  x1088 &  x1103 &  x1106 &  x1112 & ~x474 & ~x552 & ~x705 & ~x744 & ~x783;
assign c4268 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x50 &  x53 &  x56 &  x59 &  x62 &  x64 &  x65 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x194 &  x197 &  x200 &  x202 &  x203 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x245 &  x248 &  x251 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x377 &  x383 &  x389 &  x392 &  x394 &  x395 &  x398 &  x401 &  x404 &  x407 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x433 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x464 &  x467 &  x470 &  x472 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x511 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x581 &  x584 &  x587 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x725 &  x728 &  x731 &  x737 &  x743 &  x746 &  x749 &  x752 &  x758 &  x761 &  x764 &  x767 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x830 &  x833 &  x836 &  x839 &  x845 &  x848 &  x851 &  x854 &  x857 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x926 &  x929 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x952 &  x953 &  x959 &  x962 &  x965 &  x968 &  x974 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x39 & ~x78 & ~x117 & ~x156 & ~x195 & ~x360 & ~x399 & ~x438 & ~x699;
assign c4270 =  x5 &  x11 &  x14 &  x17 &  x20 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x53 &  x59 &  x62 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x149 &  x152 &  x155 &  x158 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x194 &  x197 &  x199 &  x200 &  x203 &  x206 &  x212 &  x215 &  x218 &  x221 &  x224 &  x230 &  x233 &  x238 &  x239 &  x248 &  x254 &  x260 &  x263 &  x269 &  x276 &  x277 &  x278 &  x281 &  x290 &  x296 &  x305 &  x308 &  x311 &  x313 &  x316 &  x320 &  x323 &  x326 &  x332 &  x338 &  x341 &  x347 &  x350 &  x353 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x386 &  x389 &  x394 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x425 &  x431 &  x440 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x473 &  x476 &  x485 &  x491 &  x494 &  x497 &  x500 &  x506 &  x509 &  x515 &  x518 &  x521 &  x530 &  x542 &  x545 &  x548 &  x551 &  x556 &  x560 &  x566 &  x569 &  x572 &  x578 &  x581 &  x590 &  x596 &  x599 &  x608 &  x611 &  x617 &  x623 &  x632 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x668 &  x671 &  x677 &  x679 &  x683 &  x686 &  x689 &  x692 &  x695 &  x704 &  x707 &  x713 &  x716 &  x719 &  x725 &  x734 &  x737 &  x743 &  x746 &  x749 &  x752 &  x755 &  x761 &  x764 &  x773 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x818 &  x821 &  x833 &  x835 &  x839 &  x842 &  x845 &  x848 &  x851 &  x857 &  x860 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x902 &  x905 &  x908 &  x910 &  x911 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x953 &  x956 &  x959 &  x962 &  x965 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x995 &  x998 &  x1007 &  x1010 &  x1013 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1073 &  x1076 &  x1085 &  x1091 &  x1097 &  x1106 &  x1109 &  x1112 &  x1121 &  x1127 &  x1130 & ~x318 & ~x357 & ~x358 & ~x396 & ~x435 & ~x588 & ~x783 & ~x822;
assign c4272 =  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x32 &  x35 &  x38 &  x41 &  x43 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x79 &  x80 &  x82 &  x89 &  x101 &  x104 &  x107 &  x116 &  x125 &  x128 &  x131 &  x137 &  x143 &  x146 &  x149 &  x152 &  x157 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x191 &  x194 &  x196 &  x200 &  x203 &  x209 &  x218 &  x221 &  x224 &  x235 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x274 &  x275 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x313 &  x314 &  x317 &  x326 &  x332 &  x341 &  x347 &  x350 &  x352 &  x353 &  x356 &  x362 &  x365 &  x371 &  x380 &  x392 &  x401 &  x404 &  x407 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x437 &  x446 &  x455 &  x461 &  x467 &  x470 &  x473 &  x479 &  x481 &  x482 &  x485 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x517 &  x520 &  x521 &  x523 &  x524 &  x530 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x560 &  x563 &  x566 &  x569 &  x572 &  x584 &  x587 &  x590 &  x595 &  x596 &  x599 &  x602 &  x608 &  x614 &  x617 &  x620 &  x623 &  x629 &  x634 &  x635 &  x638 &  x640 &  x644 &  x647 &  x649 &  x650 &  x653 &  x668 &  x674 &  x677 &  x679 &  x680 &  x683 &  x686 &  x688 &  x689 &  x691 &  x695 &  x698 &  x701 &  x704 &  x710 &  x716 &  x722 &  x725 &  x727 &  x728 &  x730 &  x731 &  x743 &  x749 &  x752 &  x754 &  x755 &  x758 &  x761 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x815 &  x821 &  x824 &  x827 &  x830 &  x833 &  x838 &  x842 &  x845 &  x848 &  x851 &  x856 &  x857 &  x860 &  x863 &  x866 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x905 &  x908 &  x911 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x944 &  x947 &  x959 &  x962 &  x965 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1022 &  x1025 &  x1034 &  x1040 &  x1043 &  x1052 &  x1064 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1097 &  x1106 &  x1115 &  x1118 &  x1127 &  x1130;
assign c4274 =  x2 &  x5 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x41 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x95 &  x98 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x128 &  x134 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x175 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x206 &  x212 &  x215 &  x218 &  x221 &  x227 &  x230 &  x233 &  x236 &  x239 &  x251 &  x254 &  x257 &  x260 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x362 &  x365 &  x368 &  x374 &  x377 &  x383 &  x386 &  x392 &  x395 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x434 &  x440 &  x443 &  x449 &  x452 &  x455 &  x458 &  x460 &  x461 &  x464 &  x476 &  x479 &  x482 &  x488 &  x491 &  x493 &  x494 &  x496 &  x497 &  x499 &  x500 &  x506 &  x509 &  x512 &  x514 &  x515 &  x521 &  x526 &  x527 &  x530 &  x533 &  x535 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x565 &  x566 &  x569 &  x572 &  x575 &  x577 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x659 &  x665 &  x667 &  x668 &  x671 &  x677 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x728 &  x731 &  x737 &  x745 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x779 &  x782 &  x785 &  x788 &  x794 &  x797 &  x800 &  x806 &  x809 &  x815 &  x818 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x866 &  x869 &  x872 &  x878 &  x884 &  x887 &  x890 &  x899 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x983 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x429 & ~x852;
assign c4276 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x197 &  x199 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x238 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x277 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x314 &  x315 &  x316 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x355 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x433 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x520 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x562 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x623 &  x626 &  x629 &  x632 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x679 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x869 &  x872 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x396 & ~x435 & ~x436 & ~x474 & ~x475 & ~x513;
assign c4278 =  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x41 &  x44 &  x47 &  x50 &  x59 &  x62 &  x68 &  x71 &  x74 &  x77 &  x86 &  x92 &  x95 &  x101 &  x104 &  x107 &  x110 &  x113 &  x128 &  x131 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x167 &  x170 &  x173 &  x176 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x206 &  x212 &  x215 &  x221 &  x224 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x254 &  x257 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x317 &  x320 &  x323 &  x326 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x359 &  x362 &  x368 &  x371 &  x374 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x410 &  x416 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x446 &  x452 &  x455 &  x461 &  x464 &  x467 &  x470 &  x473 &  x482 &  x488 &  x491 &  x494 &  x497 &  x500 &  x509 &  x512 &  x515 &  x518 &  x524 &  x530 &  x536 &  x539 &  x544 &  x545 &  x548 &  x551 &  x554 &  x557 &  x563 &  x566 &  x569 &  x572 &  x575 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x626 &  x629 &  x638 &  x641 &  x644 &  x647 &  x653 &  x659 &  x665 &  x668 &  x671 &  x677 &  x683 &  x686 &  x689 &  x692 &  x698 &  x701 &  x707 &  x722 &  x725 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x764 &  x770 &  x776 &  x779 &  x781 &  x794 &  x797 &  x800 &  x809 &  x812 &  x818 &  x821 &  x824 &  x830 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x859 &  x860 &  x866 &  x875 &  x878 &  x881 &  x887 &  x893 &  x896 &  x902 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x944 &  x947 &  x949 &  x950 &  x956 &  x962 &  x965 &  x968 &  x971 &  x977 &  x980 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1040 &  x1049 &  x1055 &  x1058 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1091 &  x1097 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1130 & ~x594 & ~x687 & ~x726 & ~x747 & ~x765 & ~x786 & ~x882 & ~x960 & ~x1044;
assign c4280 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x82 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x107 &  x110 &  x113 &  x116 &  x119 &  x121 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x157 &  x158 &  x159 &  x160 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x196 &  x197 &  x198 &  x199 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x235 &  x236 &  x238 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x274 &  x275 &  x277 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x314 &  x316 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x356 &  x359 &  x362 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x391 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x442 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x481 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x671 &  x674 &  x677 &  x679 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x752 &  x755 &  x757 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x165 & ~x279 & ~x318 & ~x357 & ~x588 & ~x627 & ~x666 & ~x705;
assign c4282 =  x2 &  x5 &  x11 &  x17 &  x28 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x71 &  x74 &  x80 &  x82 &  x83 &  x95 &  x98 &  x101 &  x107 &  x110 &  x116 &  x118 &  x119 &  x121 &  x122 &  x125 &  x137 &  x149 &  x152 &  x155 &  x157 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x196 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x221 &  x227 &  x230 &  x233 &  x245 &  x251 &  x257 &  x260 &  x263 &  x272 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x326 &  x329 &  x332 &  x335 &  x341 &  x344 &  x350 &  x352 &  x353 &  x356 &  x362 &  x368 &  x377 &  x380 &  x383 &  x386 &  x392 &  x395 &  x401 &  x404 &  x413 &  x416 &  x425 &  x428 &  x431 &  x437 &  x440 &  x443 &  x446 &  x449 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x503 &  x506 &  x512 &  x515 &  x518 &  x520 &  x523 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x551 &  x554 &  x560 &  x563 &  x566 &  x569 &  x578 &  x590 &  x593 &  x596 &  x599 &  x601 &  x602 &  x605 &  x608 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x640 &  x644 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x674 &  x677 &  x679 &  x683 &  x686 &  x698 &  x701 &  x707 &  x710 &  x713 &  x718 &  x719 &  x722 &  x728 &  x737 &  x740 &  x743 &  x746 &  x752 &  x755 &  x757 &  x758 &  x760 &  x761 &  x764 &  x767 &  x770 &  x782 &  x785 &  x788 &  x791 &  x794 &  x796 &  x797 &  x799 &  x800 &  x803 &  x809 &  x818 &  x821 &  x824 &  x827 &  x830 &  x835 &  x836 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x863 &  x869 &  x872 &  x874 &  x875 &  x881 &  x893 &  x896 &  x898 &  x899 &  x905 &  x908 &  x911 &  x913 &  x914 &  x920 &  x923 &  x929 &  x932 &  x937 &  x938 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x977 &  x980 &  x989 &  x1001 &  x1004 &  x1010 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1054 &  x1055 &  x1058 &  x1064 &  x1069 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1091 &  x1093 &  x1094 &  x1097 &  x1100 &  x1109 &  x1112 &  x1118 &  x1124 &  x1127;
assign c4284 =  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x47 &  x50 &  x59 &  x62 &  x65 &  x71 &  x77 &  x80 &  x83 &  x89 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x121 &  x128 &  x134 &  x137 &  x143 &  x146 &  x152 &  x155 &  x158 &  x160 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x188 &  x191 &  x194 &  x196 &  x197 &  x203 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x248 &  x251 &  x257 &  x263 &  x266 &  x272 &  x275 &  x278 &  x281 &  x287 &  x290 &  x296 &  x299 &  x302 &  x311 &  x314 &  x317 &  x320 &  x323 &  x329 &  x332 &  x338 &  x341 &  x344 &  x356 &  x362 &  x365 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x395 &  x401 &  x404 &  x407 &  x410 &  x419 &  x422 &  x425 &  x431 &  x434 &  x437 &  x440 &  x443 &  x449 &  x452 &  x455 &  x461 &  x467 &  x473 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x542 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x584 &  x587 &  x590 &  x602 &  x611 &  x620 &  x623 &  x626 &  x632 &  x635 &  x638 &  x641 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x698 &  x701 &  x707 &  x710 &  x713 &  x719 &  x722 &  x728 &  x731 &  x734 &  x737 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x773 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x830 &  x833 &  x848 &  x854 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x893 &  x899 &  x905 &  x908 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x938 &  x941 &  x947 &  x950 &  x959 &  x965 &  x968 &  x974 &  x977 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1019 &  x1028 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1073 &  x1082 &  x1085 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1115 &  x1121 &  x1124 &  x1127 & ~x9 & ~x33 & ~x48 & ~x51 & ~x99 & ~x270 & ~x309 & ~x504;
assign c4286 =  x5 &  x20 &  x26 &  x32 &  x38 &  x44 &  x53 &  x56 &  x59 &  x62 &  x68 &  x74 &  x77 &  x83 &  x89 &  x92 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x125 &  x131 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x167 &  x170 &  x173 &  x176 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x215 &  x221 &  x230 &  x242 &  x245 &  x251 &  x257 &  x263 &  x266 &  x269 &  x272 &  x278 &  x281 &  x287 &  x290 &  x293 &  x302 &  x308 &  x323 &  x326 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x377 &  x383 &  x386 &  x389 &  x395 &  x398 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x437 &  x443 &  x446 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x479 &  x484 &  x485 &  x488 &  x491 &  x497 &  x500 &  x506 &  x509 &  x512 &  x515 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x545 &  x551 &  x557 &  x560 &  x569 &  x572 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x601 &  x602 &  x605 &  x611 &  x614 &  x620 &  x623 &  x626 &  x632 &  x638 &  x641 &  x644 &  x647 &  x653 &  x656 &  x662 &  x665 &  x671 &  x674 &  x677 &  x683 &  x692 &  x704 &  x707 &  x713 &  x716 &  x719 &  x722 &  x728 &  x731 &  x734 &  x740 &  x743 &  x752 &  x755 &  x758 &  x764 &  x770 &  x773 &  x776 &  x779 &  x782 &  x788 &  x791 &  x794 &  x797 &  x800 &  x824 &  x827 &  x830 &  x833 &  x836 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x863 &  x866 &  x869 &  x875 &  x881 &  x887 &  x890 &  x899 &  x902 &  x914 &  x917 &  x923 &  x929 &  x938 &  x941 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x980 &  x983 &  x986 &  x989 &  x990 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1015 &  x1016 &  x1019 &  x1022 &  x1025 &  x1030 &  x1031 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1070 &  x1076 &  x1079 &  x1093 &  x1094 &  x1097 &  x1103 &  x1109 &  x1115 &  x1118 &  x1127 & ~x393 & ~x585 & ~x930 & ~x1020;
assign c4288 =  x8 &  x26 &  x35 &  x38 &  x44 &  x50 &  x53 &  x62 &  x71 &  x83 &  x89 &  x98 &  x110 &  x143 &  x170 &  x185 &  x191 &  x197 &  x200 &  x224 &  x227 &  x236 &  x251 &  x263 &  x272 &  x278 &  x287 &  x293 &  x296 &  x308 &  x314 &  x323 &  x326 &  x329 &  x332 &  x350 &  x353 &  x362 &  x365 &  x395 &  x419 &  x434 &  x440 &  x446 &  x452 &  x467 &  x479 &  x481 &  x482 &  x485 &  x494 &  x506 &  x515 &  x554 &  x563 &  x569 &  x572 &  x578 &  x599 &  x602 &  x617 &  x632 &  x635 &  x641 &  x647 &  x653 &  x659 &  x665 &  x671 &  x674 &  x683 &  x692 &  x698 &  x704 &  x707 &  x716 &  x719 &  x728 &  x734 &  x752 &  x764 &  x773 &  x779 &  x788 &  x797 &  x806 &  x830 &  x832 &  x836 &  x839 &  x871 &  x893 &  x905 &  x911 &  x920 &  x926 &  x941 &  x947 &  x950 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x1007 &  x1031 &  x1043 &  x1049 &  x1073 &  x1097 &  x1100 &  x1109 & ~x204 & ~x633 & ~x786 & ~x1095;
assign c4290 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x113 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x191 &  x194 &  x197 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x238 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x276 &  x277 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x315 &  x316 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x355 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x391 &  x392 &  x394 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x433 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x497 &  x500 &  x503 &  x506 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x556 &  x557 &  x560 &  x563 &  x566 &  x569 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x595 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x634 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x396 & ~x435 & ~x513 & ~x588 & ~x705 & ~x744 & ~x783 & ~x822 & ~x861 & ~x1053 & ~x1092;
assign c4292 =  x59 &  x89 &  x128 &  x143 &  x185 &  x200 &  x203 &  x209 &  x224 &  x230 &  x305 &  x344 &  x373 &  x398 &  x401 &  x449 &  x479 &  x488 &  x491 &  x500 &  x524 &  x547 &  x557 &  x602 &  x608 &  x625 &  x626 &  x629 &  x638 &  x647 &  x656 &  x664 &  x665 &  x707 &  x719 &  x722 &  x737 &  x754 &  x776 &  x781 &  x791 &  x797 &  x806 &  x866 &  x868 &  x887 &  x899 &  x902 &  x971 &  x986 &  x992 &  x995 &  x1049 &  x1070 &  x1073 &  x1082 &  x1097 &  x1103 & ~x504 & ~x555 & ~x978 & ~x1017;
assign c4294 =  x2 &  x5 &  x11 &  x14 &  x20 &  x26 &  x32 &  x41 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x74 &  x80 &  x86 &  x92 &  x95 &  x98 &  x101 &  x107 &  x113 &  x119 &  x122 &  x125 &  x128 &  x134 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x170 &  x173 &  x179 &  x182 &  x191 &  x194 &  x197 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x248 &  x251 &  x263 &  x269 &  x278 &  x284 &  x287 &  x293 &  x296 &  x302 &  x305 &  x308 &  x311 &  x314 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x350 &  x353 &  x356 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x389 &  x392 &  x395 &  x398 &  x404 &  x407 &  x416 &  x422 &  x425 &  x428 &  x431 &  x434 &  x440 &  x443 &  x449 &  x452 &  x458 &  x461 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x494 &  x500 &  x506 &  x509 &  x512 &  x515 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x590 &  x599 &  x605 &  x608 &  x614 &  x617 &  x620 &  x623 &  x629 &  x632 &  x635 &  x638 &  x641 &  x647 &  x650 &  x656 &  x665 &  x668 &  x674 &  x680 &  x683 &  x689 &  x692 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x718 &  x719 &  x722 &  x725 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x757 &  x758 &  x761 &  x764 &  x767 &  x770 &  x776 &  x779 &  x782 &  x788 &  x791 &  x796 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x824 &  x827 &  x833 &  x835 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x863 &  x866 &  x869 &  x874 &  x875 &  x878 &  x881 &  x884 &  x887 &  x893 &  x896 &  x899 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x941 &  x944 &  x950 &  x953 &  x959 &  x965 &  x971 &  x974 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1058 &  x1064 &  x1067 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1130 & ~x348 & ~x459 & ~x525 & ~x564 & ~x777 & ~x778 & ~x1038;
assign c4296 =  x5 &  x14 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x59 &  x65 &  x68 &  x80 &  x82 &  x86 &  x89 &  x98 &  x101 &  x107 &  x110 &  x116 &  x119 &  x120 &  x121 &  x122 &  x125 &  x131 &  x134 &  x137 &  x140 &  x149 &  x152 &  x157 &  x158 &  x170 &  x176 &  x179 &  x185 &  x191 &  x194 &  x199 &  x200 &  x206 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x254 &  x269 &  x274 &  x278 &  x284 &  x287 &  x293 &  x296 &  x305 &  x311 &  x317 &  x320 &  x323 &  x332 &  x338 &  x341 &  x344 &  x350 &  x371 &  x374 &  x377 &  x383 &  x386 &  x401 &  x404 &  x416 &  x419 &  x428 &  x431 &  x440 &  x443 &  x446 &  x449 &  x458 &  x461 &  x464 &  x467 &  x473 &  x476 &  x479 &  x485 &  x494 &  x503 &  x509 &  x518 &  x521 &  x523 &  x524 &  x530 &  x539 &  x545 &  x551 &  x554 &  x557 &  x560 &  x566 &  x569 &  x584 &  x593 &  x596 &  x605 &  x611 &  x620 &  x626 &  x629 &  x632 &  x635 &  x641 &  x644 &  x650 &  x656 &  x665 &  x679 &  x680 &  x692 &  x698 &  x710 &  x713 &  x716 &  x718 &  x725 &  x728 &  x731 &  x737 &  x740 &  x755 &  x767 &  x770 &  x773 &  x776 &  x779 &  x785 &  x788 &  x791 &  x794 &  x800 &  x803 &  x815 &  x821 &  x824 &  x827 &  x833 &  x835 &  x839 &  x842 &  x848 &  x851 &  x854 &  x863 &  x866 &  x893 &  x899 &  x902 &  x911 &  x914 &  x920 &  x929 &  x932 &  x938 &  x947 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x995 &  x1004 &  x1007 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1067 &  x1070 &  x1076 &  x1085 &  x1091 &  x1097 &  x1103 &  x1106 &  x1112 &  x1115 &  x1117 &  x1118 &  x1121 &  x1124 &  x1130 & ~x105 & ~x357 & ~x501;
assign c4298 =  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x29 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x194 &  x197 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x230 &  x233 &  x238 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x277 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x316 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x398 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x434 &  x440 &  x443 &  x449 &  x452 &  x458 &  x464 &  x467 &  x470 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x542 &  x545 &  x548 &  x554 &  x557 &  x560 &  x563 &  x566 &  x572 &  x575 &  x578 &  x587 &  x590 &  x593 &  x596 &  x599 &  x605 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x671 &  x674 &  x680 &  x683 &  x686 &  x692 &  x695 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x725 &  x728 &  x731 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x824 &  x830 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x857 &  x869 &  x872 &  x878 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x947 &  x953 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x980 &  x983 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1025 &  x1031 &  x1034 &  x1040 &  x1043 &  x1045 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1084 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x15 & ~x54 & ~x138 & ~x465 & ~x744 & ~x783 & ~x822 & ~x861 & ~x900 & ~x939 & ~x978 & ~x1014 & ~x1092;
assign c41 =  x5 &  x14 &  x20 &  x23 &  x29 &  x44 &  x56 &  x59 &  x65 &  x77 &  x98 &  x107 &  x122 &  x137 &  x140 &  x185 &  x197 &  x215 &  x218 &  x224 &  x230 &  x239 &  x242 &  x245 &  x284 &  x296 &  x299 &  x311 &  x323 &  x329 &  x338 &  x352 &  x355 &  x391 &  x398 &  x401 &  x407 &  x413 &  x422 &  x431 &  x458 &  x464 &  x467 &  x479 &  x491 &  x497 &  x506 &  x512 &  x542 &  x551 &  x563 &  x578 &  x596 &  x602 &  x608 &  x611 &  x623 &  x650 &  x659 &  x695 &  x740 &  x773 &  x788 &  x806 &  x818 &  x827 &  x836 &  x839 &  x851 &  x860 &  x863 &  x872 &  x875 &  x896 &  x938 &  x941 &  x944 &  x953 &  x1004 &  x1025 &  x1028 &  x1055 &  x1064 &  x1097 &  x1103 &  x1106 &  x1127 & ~x363 & ~x402 & ~x480 & ~x585 & ~x597 & ~x780;
assign c43 =  x38 &  x101 &  x191 &  x293 &  x302 &  x335 &  x359 &  x380 &  x392 &  x398 &  x443 &  x449 &  x472 &  x473 &  x494 &  x503 &  x515 &  x524 &  x553 &  x574 &  x605 &  x608 &  x631 &  x649 &  x653 &  x671 &  x688 &  x731 &  x754 &  x803 &  x832 &  x881 &  x923 &  x949 &  x983 &  x988 & ~x663;
assign c45 =  x399 &  x468 & ~x198;
assign c47 =  x131 &  x251 &  x377 &  x398 &  x434 &  x440 &  x491 &  x494 &  x505 &  x530 &  x605 &  x659 &  x749 &  x815 &  x854 &  x875 &  x896 &  x938 &  x1034 &  x1097 &  x1121 & ~x468 & ~x585 & ~x669 & ~x708 & ~x870 & ~x909;
assign c49 =  x35 &  x74 &  x188 &  x194 &  x248 &  x343 &  x395 &  x485 &  x692 &  x719 &  x776 &  x800 &  x898 &  x989 &  x1056 &  x1095 & ~x954 & ~x1104;
assign c411 =  x5 &  x14 &  x113 &  x128 &  x149 &  x173 &  x194 &  x209 &  x218 &  x233 &  x272 &  x436 &  x440 &  x443 &  x458 &  x473 &  x485 &  x514 &  x524 &  x563 &  x599 &  x629 &  x668 &  x824 &  x875 &  x911 &  x937 &  x944 &  x986 &  x1001 &  x1094 &  x1118 &  x1127 & ~x588 & ~x909 & ~x1026 & ~x1105;
assign c413 =  x17 &  x200 &  x245 &  x317 &  x344 &  x509 &  x814 &  x917 &  x962 &  x1109 & ~x87 & ~x126 & ~x273 & ~x354 & ~x843;
assign c415 =  x143 &  x152 &  x167 &  x320 &  x341 &  x343 &  x481 &  x509 &  x559 &  x566 &  x665 &  x668 &  x749 &  x755 &  x1037 &  x1073 &  x1127 & ~x393 & ~x726 & ~x909 & ~x987;
assign c417 =  x10 &  x14 &  x17 &  x20 &  x23 &  x29 &  x32 &  x35 &  x38 &  x50 &  x53 &  x56 &  x62 &  x71 &  x77 &  x83 &  x86 &  x101 &  x104 &  x146 &  x158 &  x167 &  x173 &  x185 &  x197 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x230 &  x257 &  x278 &  x287 &  x290 &  x296 &  x299 &  x302 &  x323 &  x332 &  x335 &  x350 &  x368 &  x371 &  x374 &  x380 &  x386 &  x389 &  x392 &  x404 &  x407 &  x410 &  x419 &  x434 &  x449 &  x461 &  x470 &  x473 &  x491 &  x503 &  x506 &  x512 &  x518 &  x524 &  x530 &  x536 &  x542 &  x548 &  x551 &  x554 &  x557 &  x566 &  x578 &  x581 &  x584 &  x602 &  x608 &  x614 &  x617 &  x626 &  x635 &  x638 &  x641 &  x647 &  x659 &  x677 &  x689 &  x695 &  x710 &  x713 &  x716 &  x719 &  x722 &  x746 &  x755 &  x758 &  x760 &  x770 &  x773 &  x779 &  x782 &  x788 &  x791 &  x800 &  x815 &  x818 &  x821 &  x836 &  x839 &  x842 &  x848 &  x860 &  x863 &  x872 &  x877 &  x890 &  x905 &  x908 &  x917 &  x920 &  x923 &  x926 &  x962 &  x1001 &  x1004 &  x1022 &  x1031 &  x1058 &  x1061 &  x1073 &  x1085 &  x1103 &  x1109 &  x1124 & ~x441 & ~x585 & ~x741 & ~x780 & ~x783;
assign c419 =  x239 &  x322 &  x326 &  x329 &  x361 & ~x117 & ~x195 & ~x396 & ~x531;
assign c421 =  x335 &  x446 &  x533 &  x706 &  x863 &  x959 & ~x354 & ~x393 & ~x432 & ~x513 & ~x592;
assign c423 =  x10 &  x23 &  x38 &  x161 &  x179 &  x260 &  x263 &  x356 &  x374 &  x389 &  x437 &  x521 &  x548 &  x551 &  x560 &  x584 &  x592 &  x623 &  x632 &  x656 &  x698 &  x719 &  x737 &  x767 &  x806 &  x833 &  x884 &  x890 &  x920 &  x995 &  x1009 &  x1022 &  x1043 &  x1061 &  x1085 &  x1097 & ~x831 & ~x870 & ~x909 & ~x1065;
assign c425 =  x71 &  x194 &  x215 &  x248 &  x283 &  x293 &  x361 &  x469 &  x470 &  x527 &  x608 &  x689 &  x812 &  x833 &  x1004 &  x1091 &  x1106 & ~x195 & ~x435 & ~x672;
assign c427 =  x236 &  x248 &  x323 &  x356 &  x395 &  x397 &  x410 &  x485 &  x488 &  x524 &  x566 &  x592 &  x740 &  x764 &  x815 &  x844 &  x887 &  x950 &  x965 &  x977 &  x1007 &  x1060 & ~x363 & ~x906;
assign c429 =  x80 &  x83 &  x104 &  x131 &  x179 &  x200 &  x212 &  x283 &  x287 &  x296 &  x321 &  x371 &  x377 &  x389 &  x395 &  x400 &  x542 &  x566 &  x614 &  x674 &  x725 &  x746 &  x914 &  x923 &  x929 &  x938 &  x1007 & ~x48 & ~x156;
assign c431 =  x23 &  x59 &  x71 &  x98 &  x164 &  x188 &  x212 &  x245 &  x410 &  x413 &  x437 &  x521 &  x529 &  x533 &  x602 &  x614 &  x650 &  x653 &  x680 &  x692 &  x701 &  x728 &  x764 &  x785 &  x815 &  x842 &  x848 &  x850 &  x980 &  x1006 &  x1016 &  x1028 &  x1040 & ~x3 & ~x42;
assign c433 =  x11 &  x14 &  x23 &  x47 &  x59 &  x86 &  x152 &  x185 &  x188 &  x278 &  x347 &  x383 &  x506 &  x509 &  x539 &  x572 &  x578 &  x581 &  x590 &  x647 &  x650 &  x662 &  x722 &  x737 &  x743 &  x746 &  x752 &  x758 &  x788 &  x827 &  x851 &  x863 &  x866 &  x881 &  x893 &  x911 &  x998 &  x1016 &  x1031 &  x1046 &  x1057 & ~x726 & ~x972 & ~x987 & ~x990;
assign c435 =  x358 &  x943 & ~x393 & ~x510 & ~x876;
assign c437 =  x53 &  x88 &  x125 &  x127 &  x134 &  x166 &  x230 &  x234 &  x269 &  x290 &  x329 &  x386 &  x497 &  x532 &  x596 &  x626 &  x677 &  x704 &  x794 &  x806 &  x830 &  x854 &  x875 &  x881 &  x944 &  x1028 &  x1100 & ~x585 & ~x702;
assign c439 =  x256 &  x326 &  x451 &  x482 &  x544 &  x676 &  x716 &  x727 &  x911 &  x914 &  x956 &  x1060 & ~x906;
assign c441 =  x191 &  x248 &  x352 &  x385 &  x391 &  x463 &  x502 &  x656 &  x734 &  x896 & ~x376 & ~x477 & ~x516 & ~x555;
assign c443 =  x8 &  x29 &  x32 &  x50 &  x83 &  x95 &  x107 &  x143 &  x164 &  x173 &  x179 &  x206 &  x227 &  x230 &  x239 &  x245 &  x254 &  x263 &  x266 &  x281 &  x293 &  x305 &  x314 &  x332 &  x340 &  x341 &  x347 &  x350 &  x362 &  x368 &  x377 &  x379 &  x383 &  x386 &  x403 &  x409 &  x418 &  x428 &  x437 &  x442 &  x460 &  x461 &  x476 &  x485 &  x487 &  x500 &  x515 &  x530 &  x560 &  x569 &  x572 &  x581 &  x593 &  x611 &  x614 &  x626 &  x634 &  x638 &  x650 &  x674 &  x695 &  x698 &  x710 &  x716 &  x728 &  x737 &  x740 &  x746 &  x751 &  x752 &  x791 &  x794 &  x821 &  x833 &  x836 &  x857 &  x881 &  x896 &  x905 &  x908 &  x944 &  x959 &  x974 &  x977 &  x998 &  x1001 &  x1022 &  x1070 &  x1076 &  x1085 &  x1091 &  x1094 &  x1112 &  x1127 & ~x351 & ~x390 & ~x429 & ~x432;
assign c445 =  x502 &  x981 & ~x282;
assign c447 =  x35 &  x59 &  x62 &  x77 &  x95 &  x140 &  x217 &  x322 &  x368 &  x407 &  x439 &  x488 &  x587 &  x713 &  x725 &  x740 &  x746 &  x752 &  x764 &  x806 &  x824 &  x842 &  x860 &  x935 &  x989 &  x1010 &  x1073 & ~x123 & ~x876 & ~x939 & ~x1005;
assign c449 =  x704 &  x751 & ~x579 & ~x954;
assign c451 =  x2 &  x14 &  x20 &  x23 &  x29 &  x32 &  x38 &  x44 &  x47 &  x50 &  x53 &  x59 &  x62 &  x68 &  x74 &  x83 &  x86 &  x98 &  x107 &  x110 &  x116 &  x119 &  x134 &  x146 &  x152 &  x155 &  x158 &  x161 &  x170 &  x173 &  x179 &  x185 &  x188 &  x191 &  x197 &  x200 &  x203 &  x206 &  x212 &  x218 &  x221 &  x236 &  x239 &  x242 &  x248 &  x251 &  x260 &  x263 &  x269 &  x272 &  x275 &  x281 &  x284 &  x287 &  x293 &  x302 &  x314 &  x320 &  x323 &  x332 &  x335 &  x338 &  x347 &  x359 &  x362 &  x365 &  x371 &  x374 &  x380 &  x383 &  x389 &  x392 &  x395 &  x401 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x434 &  x440 &  x443 &  x446 &  x452 &  x455 &  x464 &  x467 &  x470 &  x473 &  x476 &  x482 &  x485 &  x488 &  x494 &  x500 &  x509 &  x512 &  x527 &  x530 &  x533 &  x539 &  x542 &  x548 &  x551 &  x554 &  x557 &  x560 &  x572 &  x575 &  x578 &  x581 &  x590 &  x602 &  x611 &  x614 &  x620 &  x623 &  x629 &  x635 &  x638 &  x641 &  x653 &  x659 &  x665 &  x668 &  x671 &  x673 &  x674 &  x689 &  x692 &  x698 &  x704 &  x710 &  x725 &  x728 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x773 &  x776 &  x779 &  x782 &  x785 &  x790 &  x797 &  x800 &  x803 &  x815 &  x818 &  x827 &  x833 &  x836 &  x839 &  x842 &  x845 &  x851 &  x854 &  x857 &  x863 &  x872 &  x875 &  x881 &  x887 &  x893 &  x902 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x941 &  x947 &  x953 &  x962 &  x965 &  x968 &  x971 &  x974 &  x980 &  x986 &  x989 &  x992 &  x1004 &  x1007 &  x1013 &  x1019 &  x1022 &  x1034 &  x1037 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1076 &  x1079 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1112 &  x1115 &  x1130 & ~x48 & ~x165 & ~x234 & ~x354 & ~x432;
assign c453 =  x5 &  x17 &  x29 &  x38 &  x53 &  x68 &  x77 &  x104 &  x128 &  x152 &  x155 &  x161 &  x170 &  x239 &  x245 &  x269 &  x272 &  x290 &  x299 &  x331 &  x335 &  x353 &  x368 &  x401 &  x449 &  x452 &  x455 &  x509 &  x521 &  x584 &  x623 &  x629 &  x644 &  x664 &  x728 &  x782 &  x797 &  x815 &  x818 &  x824 &  x827 &  x836 &  x902 &  x923 &  x937 &  x956 &  x974 &  x998 &  x1019 &  x1025 &  x1040 &  x1073 &  x1085 &  x1091 & ~x687 & ~x792 & ~x948 & ~x987 & ~x1027;
assign c455 =  x547 &  x625 &  x629 &  x908 & ~x234 & ~x354 & ~x492 & ~x513;
assign c457 =  x801 & ~x160;
assign c459 =  x2 &  x11 &  x23 &  x32 &  x35 &  x41 &  x53 &  x56 &  x59 &  x62 &  x68 &  x74 &  x77 &  x80 &  x83 &  x92 &  x101 &  x104 &  x122 &  x128 &  x134 &  x137 &  x140 &  x143 &  x152 &  x155 &  x161 &  x167 &  x170 &  x173 &  x178 &  x179 &  x188 &  x191 &  x194 &  x203 &  x209 &  x215 &  x218 &  x221 &  x239 &  x251 &  x254 &  x256 &  x263 &  x266 &  x269 &  x275 &  x278 &  x287 &  x290 &  x293 &  x296 &  x299 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x338 &  x341 &  x350 &  x359 &  x362 &  x374 &  x380 &  x386 &  x395 &  x407 &  x410 &  x413 &  x434 &  x439 &  x446 &  x449 &  x455 &  x458 &  x476 &  x478 &  x482 &  x488 &  x491 &  x494 &  x506 &  x509 &  x512 &  x521 &  x530 &  x536 &  x547 &  x554 &  x557 &  x563 &  x566 &  x581 &  x584 &  x586 &  x590 &  x596 &  x599 &  x605 &  x611 &  x617 &  x620 &  x623 &  x632 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x662 &  x664 &  x671 &  x680 &  x683 &  x686 &  x689 &  x695 &  x698 &  x701 &  x703 &  x707 &  x716 &  x725 &  x734 &  x740 &  x746 &  x749 &  x755 &  x758 &  x788 &  x791 &  x797 &  x806 &  x809 &  x815 &  x818 &  x821 &  x830 &  x833 &  x836 &  x839 &  x842 &  x854 &  x857 &  x859 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x887 &  x893 &  x896 &  x898 &  x902 &  x905 &  x908 &  x917 &  x919 &  x926 &  x929 &  x937 &  x944 &  x950 &  x953 &  x956 &  x958 &  x965 &  x971 &  x976 &  x977 &  x983 &  x989 &  x992 &  x1004 &  x1019 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1058 &  x1067 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1100 &  x1103 &  x1106 &  x1118 &  x1121 & ~x513 & ~x591;
assign c461 =  x442 &  x546 &  x586 &  x893 &  x968 & ~x393 & ~x792;
assign c463 =  x438 &  x449 &  x673 &  x841 & ~x120;
assign c465 =  x89 &  x1111 & ~x675 & ~x756 & ~x757;
assign c467 =  x71 &  x92 &  x98 &  x125 &  x227 &  x263 &  x299 &  x308 &  x343 &  x380 &  x403 &  x442 &  x449 &  x476 &  x479 &  x500 &  x506 &  x523 &  x539 &  x614 &  x647 &  x665 &  x668 &  x686 &  x695 &  x728 &  x742 &  x809 &  x821 &  x839 &  x872 &  x929 &  x938 &  x950 &  x953 &  x998 &  x1058 &  x1067 &  x1079 &  x1106 & ~x792 & ~x831 & ~x870 & ~x909 & ~x987 & ~x1065;
assign c469 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x23 &  x29 &  x32 &  x38 &  x41 &  x47 &  x50 &  x53 &  x62 &  x68 &  x71 &  x74 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x107 &  x110 &  x122 &  x125 &  x134 &  x137 &  x143 &  x149 &  x152 &  x155 &  x158 &  x164 &  x167 &  x170 &  x173 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x212 &  x224 &  x227 &  x233 &  x236 &  x245 &  x248 &  x263 &  x266 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x323 &  x326 &  x329 &  x332 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x359 &  x365 &  x368 &  x371 &  x386 &  x391 &  x392 &  x401 &  x407 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x470 &  x476 &  x479 &  x482 &  x485 &  x488 &  x500 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x533 &  x536 &  x542 &  x545 &  x548 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x584 &  x587 &  x590 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x635 &  x638 &  x641 &  x644 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x704 &  x707 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x740 &  x743 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x773 &  x776 &  x779 &  x782 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x809 &  x812 &  x815 &  x821 &  x827 &  x833 &  x839 &  x842 &  x845 &  x848 &  x857 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1010 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1094 &  x1103 &  x1106 &  x1109 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x402 & ~x441 & ~x480 & ~x585 & ~x597 & ~x663 & ~x705 & ~x744 & ~x783 & ~x822 & ~x861;
assign c471 =  x5 &  x11 &  x17 &  x20 &  x23 &  x26 &  x29 &  x38 &  x44 &  x47 &  x50 &  x53 &  x59 &  x62 &  x68 &  x71 &  x77 &  x80 &  x83 &  x89 &  x95 &  x101 &  x116 &  x122 &  x125 &  x128 &  x131 &  x140 &  x149 &  x155 &  x158 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x224 &  x227 &  x230 &  x233 &  x239 &  x242 &  x245 &  x248 &  x251 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x401 &  x407 &  x410 &  x419 &  x434 &  x440 &  x443 &  x446 &  x449 &  x452 &  x458 &  x461 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x488 &  x491 &  x500 &  x509 &  x512 &  x515 &  x518 &  x521 &  x526 &  x527 &  x529 &  x530 &  x533 &  x536 &  x539 &  x551 &  x554 &  x560 &  x563 &  x565 &  x566 &  x569 &  x572 &  x575 &  x581 &  x587 &  x590 &  x593 &  x599 &  x605 &  x614 &  x617 &  x620 &  x623 &  x629 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x665 &  x668 &  x671 &  x674 &  x683 &  x686 &  x689 &  x692 &  x695 &  x704 &  x707 &  x710 &  x712 &  x722 &  x734 &  x743 &  x746 &  x749 &  x751 &  x752 &  x755 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x794 &  x797 &  x800 &  x806 &  x809 &  x812 &  x821 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x851 &  x854 &  x857 &  x860 &  x866 &  x869 &  x872 &  x878 &  x881 &  x884 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x929 &  x938 &  x941 &  x944 &  x947 &  x950 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x989 &  x992 &  x998 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1100 &  x1103 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 & ~x432 & ~x471 & ~x837 & ~x876 & ~x954;
assign c473 =  x8 &  x29 &  x32 &  x41 &  x56 &  x65 &  x68 &  x92 &  x104 &  x110 &  x122 &  x137 &  x152 &  x176 &  x182 &  x185 &  x191 &  x194 &  x209 &  x218 &  x221 &  x227 &  x239 &  x245 &  x254 &  x257 &  x278 &  x287 &  x293 &  x296 &  x314 &  x320 &  x329 &  x338 &  x341 &  x353 &  x356 &  x359 &  x362 &  x383 &  x392 &  x401 &  x410 &  x416 &  x428 &  x431 &  x437 &  x443 &  x470 &  x473 &  x479 &  x485 &  x497 &  x503 &  x533 &  x542 &  x548 &  x557 &  x563 &  x578 &  x626 &  x632 &  x635 &  x638 &  x650 &  x653 &  x674 &  x680 &  x689 &  x698 &  x710 &  x713 &  x719 &  x722 &  x728 &  x734 &  x737 &  x743 &  x749 &  x752 &  x755 &  x770 &  x776 &  x785 &  x788 &  x818 &  x881 &  x899 &  x932 &  x941 &  x950 &  x959 &  x962 &  x977 &  x1001 &  x1010 &  x1016 &  x1022 &  x1028 &  x1037 &  x1052 &  x1064 &  x1070 &  x1076 &  x1082 &  x1121 &  x1124 &  x1127 &  x1130 & ~x78 & ~x237 & ~x276 & ~x792 & ~x897 & ~x936;
assign c475 =  x62 &  x98 &  x119 &  x179 &  x191 &  x218 &  x248 &  x254 &  x299 &  x401 &  x410 &  x416 &  x419 &  x452 &  x469 &  x479 &  x509 &  x515 &  x557 &  x575 &  x578 &  x584 &  x596 &  x608 &  x620 &  x628 &  x629 &  x641 &  x710 &  x713 &  x737 &  x761 &  x773 &  x794 &  x806 &  x809 &  x818 &  x833 &  x863 &  x875 &  x881 &  x884 &  x887 &  x905 &  x908 &  x914 &  x965 &  x983 &  x1067 &  x1106 &  x1115 &  x1121 &  x1127 & ~x531 & ~x636 & ~x675 & ~x741;
assign c477 =  x321 &  x361 &  x626 & ~x120 & ~x397;
assign c479 =  x205 &  x657 &  x769 &  x782 & ~x3;
assign c481 =  x17 &  x26 &  x80 &  x92 &  x134 &  x137 &  x197 &  x209 &  x218 &  x248 &  x266 &  x272 &  x278 &  x302 &  x314 &  x335 &  x347 &  x353 &  x383 &  x389 &  x455 &  x464 &  x470 &  x476 &  x485 &  x593 &  x595 &  x602 &  x635 &  x662 &  x664 &  x710 &  x725 &  x740 &  x806 &  x854 &  x863 &  x875 &  x881 &  x890 &  x932 &  x956 &  x1001 &  x1025 &  x1040 & ~x156 & ~x195 & ~x315 & ~x354 & ~x432;
assign c483 = ~x1091;
assign c485 =  x475 &  x532 &  x558 &  x636 &  x1098 & ~x546;
assign c487 =  x206 &  x299 &  x332 &  x404 &  x461 &  x479 &  x497 &  x881 &  x1001 &  x1031 &  x1070 &  x1094 & ~x339 & ~x364 & ~x402 & ~x480 & ~x519 & ~x663 & ~x672;
assign c489 =  x32 &  x65 &  x83 &  x86 &  x107 &  x122 &  x128 &  x137 &  x170 &  x185 &  x188 &  x206 &  x209 &  x233 &  x239 &  x242 &  x245 &  x260 &  x263 &  x278 &  x311 &  x479 &  x512 &  x524 &  x587 &  x617 &  x623 &  x656 &  x683 &  x709 &  x710 &  x737 &  x747 &  x749 &  x770 &  x776 &  x779 &  x787 &  x788 &  x791 &  x793 &  x809 &  x821 &  x825 &  x845 &  x857 &  x866 &  x870 &  x908 &  x917 &  x923 &  x929 &  x944 &  x947 &  x949 &  x956 &  x959 &  x965 &  x980 &  x988 &  x989 &  x995 &  x1064 &  x1088 &  x1097 &  x1100 &  x1103 &  x1112 &  x1115 &  x1121;
assign c491 =  x5 &  x11 &  x17 &  x23 &  x26 &  x44 &  x47 &  x53 &  x56 &  x80 &  x86 &  x89 &  x98 &  x101 &  x104 &  x113 &  x119 &  x122 &  x125 &  x131 &  x143 &  x152 &  x158 &  x179 &  x185 &  x188 &  x191 &  x206 &  x218 &  x224 &  x230 &  x236 &  x251 &  x269 &  x287 &  x293 &  x311 &  x320 &  x332 &  x341 &  x353 &  x359 &  x374 &  x386 &  x388 &  x392 &  x395 &  x422 &  x434 &  x443 &  x451 &  x452 &  x455 &  x466 &  x476 &  x494 &  x497 &  x503 &  x509 &  x521 &  x524 &  x542 &  x545 &  x548 &  x551 &  x554 &  x569 &  x572 &  x575 &  x581 &  x590 &  x632 &  x641 &  x644 &  x650 &  x665 &  x677 &  x692 &  x712 &  x713 &  x716 &  x722 &  x725 &  x731 &  x734 &  x740 &  x743 &  x746 &  x767 &  x770 &  x776 &  x779 &  x791 &  x797 &  x800 &  x833 &  x842 &  x851 &  x863 &  x878 &  x896 &  x905 &  x908 &  x920 &  x938 &  x941 &  x950 &  x956 &  x959 &  x962 &  x968 &  x1004 &  x1010 &  x1016 &  x1037 &  x1049 &  x1052 &  x1058 &  x1061 &  x1070 &  x1079 &  x1088 &  x1103 &  x1115 &  x1118 &  x1124 & ~x912 & ~x990;
assign c493 =  x49 &  x50 &  x91 &  x119 &  x155 &  x158 &  x164 &  x166 &  x209 &  x233 &  x242 &  x244 &  x284 &  x377 &  x413 &  x422 &  x524 &  x539 &  x542 &  x551 &  x554 &  x557 &  x581 &  x587 &  x731 &  x752 &  x773 &  x802 &  x914 &  x947 &  x959 &  x989 &  x1076 & ~x279 & ~x336 & ~x375 & ~x414;
assign c495 =  x5 &  x11 &  x13 &  x20 &  x23 &  x56 &  x74 &  x77 &  x83 &  x88 &  x89 &  x116 &  x119 &  x127 &  x146 &  x164 &  x166 &  x185 &  x188 &  x236 &  x254 &  x281 &  x284 &  x296 &  x314 &  x320 &  x323 &  x338 &  x341 &  x362 &  x365 &  x380 &  x410 &  x425 &  x428 &  x485 &  x497 &  x503 &  x506 &  x515 &  x548 &  x584 &  x596 &  x605 &  x608 &  x611 &  x653 &  x716 &  x749 &  x773 &  x782 &  x794 &  x815 &  x821 &  x848 &  x851 &  x854 &  x860 &  x866 &  x884 &  x887 &  x956 &  x959 &  x977 &  x980 &  x1007 &  x1010 &  x1016 &  x1031 &  x1040 &  x1058 &  x1094 & ~x594 & ~x633 & ~x663 & ~x705 & ~x744 & ~x783;
assign c497 =  x254 &  x347 &  x467 &  x530 &  x635 &  x749 &  x791 &  x947 &  x953 & ~x354 & ~x393 & ~x432 & ~x588 & ~x627 & ~x759 & ~x990;
assign c499 =  x23 &  x68 &  x74 &  x233 &  x322 &  x536 &  x550 &  x932 &  x1085 & ~x600 & ~x678 & ~x780 & ~x789 & ~x897;
assign c4101 =  x422 &  x432 &  x553 &  x877 &  x911 & ~x522;
assign c4103 =  x11 &  x38 &  x65 &  x86 &  x89 &  x95 &  x140 &  x152 &  x164 &  x166 &  x221 &  x235 &  x254 &  x284 &  x296 &  x313 &  x368 &  x479 &  x491 &  x500 &  x506 &  x566 &  x635 &  x731 &  x839 &  x872 &  x878 &  x908 &  x989 &  x1007 &  x1130 & ~x201 & ~x363 & ~x585 & ~x705 & ~x741;
assign c4105 =  x29 &  x74 &  x95 &  x116 &  x248 &  x260 &  x266 &  x329 &  x344 &  x371 &  x431 &  x436 &  x467 &  x470 &  x475 &  x476 &  x485 &  x553 &  x578 &  x649 &  x673 &  x692 &  x751 &  x755 &  x790 &  x908 &  x983 &  x992 &  x998 &  x1004 &  x1022 &  x1045 &  x1106 &  x1109 &  x1127 & ~x585;
assign c4107 =  x41 &  x107 &  x146 &  x152 &  x197 &  x218 &  x260 &  x287 &  x314 &  x347 &  x380 &  x383 &  x386 &  x434 &  x449 &  x469 &  x485 &  x506 &  x515 &  x563 &  x587 &  x611 &  x617 &  x638 &  x668 &  x713 &  x773 &  x800 &  x818 &  x893 &  x965 &  x977 &  x1121 & ~x81 & ~x597 & ~x636 & ~x675 & ~x702;
assign c4109 =  x589 &  x613 & ~x382 & ~x600;
assign c4111 =  x2 &  x56 &  x71 &  x119 &  x137 &  x143 &  x227 &  x248 &  x263 &  x278 &  x301 &  x311 &  x317 &  x416 &  x482 &  x506 &  x512 &  x665 &  x731 &  x815 &  x884 &  x923 &  x935 &  x941 &  x995 &  x1031 &  x1064 &  x1130 & ~x351 & ~x471 & ~x588 & ~x708 & ~x1026;
assign c4113 =  x5 &  x8 &  x11 &  x14 &  x20 &  x26 &  x32 &  x35 &  x38 &  x44 &  x50 &  x62 &  x68 &  x71 &  x74 &  x80 &  x83 &  x92 &  x101 &  x104 &  x107 &  x110 &  x116 &  x122 &  x125 &  x131 &  x140 &  x146 &  x149 &  x158 &  x164 &  x167 &  x173 &  x191 &  x200 &  x203 &  x209 &  x215 &  x218 &  x227 &  x230 &  x233 &  x239 &  x251 &  x254 &  x257 &  x260 &  x266 &  x284 &  x293 &  x299 &  x302 &  x308 &  x314 &  x316 &  x317 &  x320 &  x323 &  x332 &  x338 &  x353 &  x362 &  x368 &  x374 &  x377 &  x383 &  x386 &  x389 &  x392 &  x398 &  x401 &  x407 &  x416 &  x419 &  x422 &  x425 &  x440 &  x443 &  x446 &  x449 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x476 &  x482 &  x485 &  x491 &  x506 &  x512 &  x515 &  x518 &  x524 &  x527 &  x533 &  x536 &  x539 &  x545 &  x548 &  x551 &  x553 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x592 &  x593 &  x599 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x629 &  x632 &  x647 &  x650 &  x656 &  x659 &  x665 &  x670 &  x677 &  x686 &  x695 &  x704 &  x710 &  x716 &  x719 &  x737 &  x743 &  x746 &  x752 &  x755 &  x761 &  x773 &  x776 &  x782 &  x785 &  x794 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x824 &  x827 &  x830 &  x848 &  x854 &  x857 &  x860 &  x869 &  x872 &  x875 &  x877 &  x881 &  x887 &  x896 &  x902 &  x905 &  x908 &  x911 &  x914 &  x920 &  x929 &  x932 &  x935 &  x938 &  x941 &  x947 &  x949 &  x953 &  x959 &  x968 &  x974 &  x977 &  x980 &  x986 &  x989 &  x1013 &  x1016 &  x1022 &  x1028 &  x1034 &  x1037 &  x1040 &  x1073 &  x1076 &  x1079 &  x1082 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1130 & ~x522 & ~x663 & ~x702 & ~x741 & ~x780 & ~x858;
assign c4115 =  x272 &  x667 &  x705 &  x826 &  x1027 & ~x1053;
assign c4117 =  x712 &  x783 &  x836 &  x941 &  x982 &  x1021 &  x1064;
assign c4119 =  x169 &  x656 &  x745 & ~x835 & ~x1092;
assign c4121 =  x20 &  x35 &  x38 &  x41 &  x68 &  x143 &  x146 &  x158 &  x203 &  x215 &  x221 &  x236 &  x251 &  x257 &  x266 &  x287 &  x305 &  x320 &  x329 &  x335 &  x359 &  x374 &  x379 &  x380 &  x407 &  x436 &  x440 &  x458 &  x475 &  x514 &  x521 &  x566 &  x602 &  x605 &  x635 &  x650 &  x662 &  x664 &  x677 &  x680 &  x701 &  x725 &  x797 &  x803 &  x806 &  x821 &  x851 &  x860 &  x869 &  x878 &  x884 &  x929 &  x938 &  x968 &  x977 &  x1028 &  x1037 &  x1046 &  x1055 &  x1124 & ~x510 & ~x549 & ~x591 & ~x630;
assign c4123 =  x348 &  x368 &  x443 &  x839 &  x953 &  x1021 &  x1082 & ~x393 & ~x432;
assign c4125 =  x2 &  x10 &  x53 &  x74 &  x86 &  x88 &  x92 &  x127 &  x134 &  x137 &  x167 &  x173 &  x176 &  x188 &  x191 &  x194 &  x196 &  x203 &  x209 &  x266 &  x278 &  x284 &  x287 &  x296 &  x323 &  x326 &  x335 &  x350 &  x356 &  x380 &  x395 &  x398 &  x404 &  x461 &  x482 &  x502 &  x509 &  x527 &  x545 &  x557 &  x572 &  x575 &  x578 &  x581 &  x583 &  x584 &  x587 &  x599 &  x605 &  x614 &  x623 &  x635 &  x665 &  x716 &  x725 &  x734 &  x787 &  x788 &  x797 &  x806 &  x839 &  x845 &  x848 &  x851 &  x863 &  x872 &  x890 &  x893 &  x905 &  x917 &  x935 &  x959 &  x962 &  x965 &  x1001 &  x1007 &  x1037 &  x1052 &  x1061 &  x1085 &  x1091 &  x1129;
assign c4127 =  x891 &  x1008;
assign c4129 =  x5 &  x13 &  x17 &  x20 &  x23 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x59 &  x62 &  x71 &  x86 &  x91 &  x119 &  x128 &  x130 &  x131 &  x134 &  x149 &  x164 &  x169 &  x170 &  x194 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x227 &  x230 &  x242 &  x248 &  x254 &  x266 &  x275 &  x278 &  x281 &  x290 &  x293 &  x314 &  x317 &  x323 &  x326 &  x329 &  x332 &  x335 &  x347 &  x350 &  x365 &  x371 &  x377 &  x380 &  x383 &  x398 &  x401 &  x407 &  x422 &  x425 &  x428 &  x431 &  x437 &  x440 &  x451 &  x464 &  x467 &  x476 &  x479 &  x485 &  x491 &  x494 &  x506 &  x515 &  x518 &  x521 &  x527 &  x533 &  x554 &  x563 &  x566 &  x568 &  x575 &  x578 &  x607 &  x608 &  x611 &  x614 &  x629 &  x635 &  x644 &  x656 &  x659 &  x671 &  x683 &  x686 &  x707 &  x710 &  x713 &  x716 &  x722 &  x734 &  x737 &  x743 &  x752 &  x782 &  x785 &  x800 &  x806 &  x814 &  x815 &  x824 &  x839 &  x842 &  x845 &  x851 &  x853 &  x884 &  x887 &  x899 &  x902 &  x905 &  x919 &  x923 &  x929 &  x931 &  x932 &  x935 &  x938 &  x947 &  x956 &  x959 &  x965 &  x998 &  x1004 &  x1010 &  x1019 &  x1043 &  x1055 &  x1067 &  x1076 &  x1079 &  x1085 &  x1103 &  x1106 &  x1115 &  x1121 &  x1127 &  x1130;
assign c4131 =  x47 &  x188 &  x317 &  x355 &  x709 &  x824 &  x850 &  x908 &  x916 &  x955 &  x1052 &  x1123 & ~x561 & ~x717;
assign c4133 =  x17 &  x241 &  x479 &  x747 &  x786 &  x903 &  x1097;
assign c4135 =  x478 &  x559 &  x663 & ~x237 & ~x591;
assign c4137 =  x688 &  x694 & ~x405 & ~x445 & ~x780 & ~x819;
assign c4139 =  x204 &  x244 &  x352 &  x383 &  x479 &  x544 &  x785 &  x953 &  x1121 & ~x1107;
assign c4141 =  x478 &  x585 &  x703 &  x742 &  x898 &  x956 & ~x513 & ~x711 & ~x750;
assign c4143 =  x775 &  x817 & ~x522 & ~x562;
assign c4145 =  x2 &  x8 &  x11 &  x14 &  x20 &  x26 &  x29 &  x32 &  x35 &  x41 &  x47 &  x59 &  x62 &  x65 &  x68 &  x74 &  x77 &  x83 &  x86 &  x89 &  x110 &  x113 &  x116 &  x125 &  x137 &  x140 &  x143 &  x146 &  x152 &  x158 &  x164 &  x167 &  x182 &  x188 &  x200 &  x203 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x296 &  x305 &  x311 &  x317 &  x322 &  x335 &  x341 &  x344 &  x347 &  x353 &  x365 &  x368 &  x383 &  x386 &  x392 &  x395 &  x410 &  x413 &  x428 &  x431 &  x433 &  x434 &  x440 &  x443 &  x449 &  x452 &  x455 &  x458 &  x461 &  x467 &  x470 &  x472 &  x479 &  x482 &  x485 &  x488 &  x494 &  x497 &  x500 &  x503 &  x509 &  x511 &  x512 &  x521 &  x527 &  x533 &  x536 &  x539 &  x545 &  x548 &  x550 &  x557 &  x560 &  x563 &  x575 &  x581 &  x584 &  x587 &  x590 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x632 &  x638 &  x641 &  x647 &  x653 &  x662 &  x665 &  x668 &  x674 &  x677 &  x689 &  x701 &  x710 &  x713 &  x716 &  x719 &  x728 &  x731 &  x734 &  x740 &  x746 &  x758 &  x770 &  x773 &  x779 &  x791 &  x794 &  x803 &  x806 &  x812 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x845 &  x848 &  x851 &  x854 &  x857 &  x863 &  x872 &  x884 &  x890 &  x893 &  x896 &  x899 &  x902 &  x908 &  x914 &  x920 &  x923 &  x941 &  x947 &  x950 &  x956 &  x959 &  x965 &  x971 &  x983 &  x986 &  x995 &  x998 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1028 &  x1031 &  x1040 &  x1043 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1106 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x303 & ~x672 & ~x741 & ~x780;
assign c4147 =  x5 &  x11 &  x17 &  x20 &  x29 &  x32 &  x56 &  x71 &  x74 &  x80 &  x86 &  x98 &  x101 &  x107 &  x110 &  x131 &  x146 &  x158 &  x164 &  x188 &  x194 &  x206 &  x236 &  x239 &  x245 &  x269 &  x287 &  x329 &  x344 &  x347 &  x365 &  x368 &  x371 &  x380 &  x437 &  x446 &  x485 &  x491 &  x497 &  x524 &  x551 &  x554 &  x563 &  x572 &  x575 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x620 &  x628 &  x635 &  x644 &  x647 &  x665 &  x695 &  x701 &  x716 &  x779 &  x785 &  x791 &  x797 &  x800 &  x806 &  x809 &  x815 &  x857 &  x881 &  x902 &  x905 &  x911 &  x920 &  x980 &  x986 &  x1010 &  x1043 &  x1046 &  x1061 &  x1082 &  x1088 &  x1100 &  x1106 &  x1121 &  x1127 & ~x630 & ~x648 & ~x669 & ~x747 & ~x792 & ~x831 & ~x834;
assign c4149 =  x10 &  x29 &  x53 &  x59 &  x77 &  x88 &  x101 &  x118 &  x146 &  x236 &  x248 &  x257 &  x263 &  x266 &  x281 &  x296 &  x314 &  x353 &  x374 &  x377 &  x440 &  x455 &  x506 &  x527 &  x530 &  x557 &  x592 &  x602 &  x622 &  x626 &  x638 &  x653 &  x656 &  x665 &  x668 &  x725 &  x787 &  x826 &  x836 &  x845 &  x941 &  x989 &  x1019 &  x1070 &  x1082 &  x1088 &  x1094 &  x1121 &  x1129;
assign c4151 =  x2 &  x5 &  x11 &  x23 &  x26 &  x29 &  x32 &  x41 &  x44 &  x53 &  x59 &  x62 &  x65 &  x80 &  x83 &  x86 &  x95 &  x104 &  x116 &  x119 &  x125 &  x137 &  x140 &  x143 &  x146 &  x152 &  x158 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x197 &  x212 &  x221 &  x224 &  x233 &  x242 &  x251 &  x260 &  x269 &  x275 &  x281 &  x284 &  x290 &  x293 &  x296 &  x299 &  x301 &  x308 &  x311 &  x317 &  x320 &  x323 &  x338 &  x341 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x410 &  x413 &  x416 &  x434 &  x440 &  x443 &  x452 &  x461 &  x464 &  x467 &  x470 &  x473 &  x479 &  x482 &  x491 &  x494 &  x497 &  x506 &  x512 &  x521 &  x524 &  x527 &  x530 &  x542 &  x548 &  x551 &  x554 &  x560 &  x563 &  x566 &  x572 &  x575 &  x578 &  x584 &  x590 &  x602 &  x614 &  x623 &  x626 &  x632 &  x635 &  x641 &  x644 &  x647 &  x650 &  x665 &  x668 &  x674 &  x677 &  x692 &  x707 &  x710 &  x713 &  x719 &  x722 &  x734 &  x737 &  x740 &  x746 &  x749 &  x752 &  x755 &  x758 &  x764 &  x767 &  x779 &  x782 &  x785 &  x788 &  x800 &  x806 &  x809 &  x812 &  x814 &  x818 &  x830 &  x836 &  x839 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x893 &  x896 &  x899 &  x908 &  x914 &  x917 &  x923 &  x935 &  x941 &  x947 &  x959 &  x962 &  x965 &  x968 &  x971 &  x983 &  x986 &  x992 &  x998 &  x1034 &  x1037 &  x1040 &  x1046 &  x1052 &  x1055 &  x1058 &  x1064 &  x1067 &  x1070 &  x1079 &  x1082 &  x1085 &  x1091 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1130 & ~x354 & ~x393 & ~x630 & ~x669 & ~x831;
assign c4153 =  x29 &  x41 &  x50 &  x59 &  x74 &  x80 &  x83 &  x89 &  x104 &  x107 &  x113 &  x119 &  x152 &  x155 &  x170 &  x188 &  x197 &  x200 &  x215 &  x221 &  x227 &  x245 &  x260 &  x296 &  x317 &  x338 &  x344 &  x362 &  x368 &  x386 &  x395 &  x398 &  x410 &  x416 &  x440 &  x443 &  x446 &  x449 &  x458 &  x470 &  x473 &  x482 &  x485 &  x494 &  x512 &  x545 &  x572 &  x575 &  x587 &  x596 &  x623 &  x626 &  x632 &  x641 &  x649 &  x650 &  x656 &  x688 &  x689 &  x722 &  x727 &  x731 &  x737 &  x779 &  x791 &  x794 &  x803 &  x805 &  x812 &  x821 &  x833 &  x845 &  x857 &  x893 &  x895 &  x899 &  x902 &  x911 &  x914 &  x920 &  x923 &  x926 &  x929 &  x934 &  x941 &  x944 &  x947 &  x956 &  x983 &  x986 &  x1055 &  x1058 &  x1067 &  x1076 &  x1118 & ~x396 & ~x402 & ~x480 & ~x519 & ~x558;
assign c4155 =  x248 &  x544 &  x623 &  x635 &  x979 &  x1079 &  x1085 & ~x804 & ~x825 & ~x882 & ~x948 & ~x951 & ~x987;
assign c4157 =  x8 &  x41 &  x47 &  x59 &  x83 &  x119 &  x155 &  x179 &  x185 &  x212 &  x227 &  x248 &  x260 &  x284 &  x440 &  x467 &  x494 &  x497 &  x545 &  x599 &  x611 &  x623 &  x632 &  x677 &  x680 &  x698 &  x749 &  x785 &  x839 &  x845 &  x875 &  x898 &  x923 &  x944 &  x1004 &  x1015 &  x1037 &  x1073 &  x1100 &  x1124 & ~x276 & ~x909 & ~x954 & ~x987 & ~x990;
assign c4159 =  x11 &  x23 &  x32 &  x35 &  x41 &  x62 &  x74 &  x92 &  x104 &  x113 &  x119 &  x125 &  x131 &  x140 &  x149 &  x173 &  x182 &  x206 &  x260 &  x266 &  x269 &  x290 &  x302 &  x311 &  x316 &  x323 &  x344 &  x352 &  x359 &  x377 &  x380 &  x391 &  x398 &  x401 &  x404 &  x410 &  x422 &  x440 &  x446 &  x455 &  x458 &  x467 &  x470 &  x479 &  x485 &  x512 &  x527 &  x533 &  x548 &  x551 &  x566 &  x578 &  x581 &  x584 &  x587 &  x599 &  x611 &  x626 &  x650 &  x656 &  x665 &  x674 &  x689 &  x701 &  x707 &  x737 &  x746 &  x752 &  x755 &  x776 &  x779 &  x788 &  x818 &  x872 &  x875 &  x881 &  x911 &  x920 &  x926 &  x950 &  x1001 &  x1004 &  x1007 &  x1019 &  x1070 &  x1085 &  x1088 &  x1091 &  x1100 &  x1109 &  x1124 &  x1127 & ~x480 & ~x519 & ~x594 & ~x675 & ~x702;
assign c4161 =  x14 &  x17 &  x20 &  x32 &  x65 &  x71 &  x86 &  x113 &  x122 &  x134 &  x143 &  x146 &  x152 &  x158 &  x179 &  x188 &  x197 &  x203 &  x221 &  x230 &  x236 &  x239 &  x269 &  x290 &  x299 &  x314 &  x326 &  x329 &  x335 &  x344 &  x362 &  x368 &  x395 &  x413 &  x416 &  x425 &  x437 &  x443 &  x449 &  x458 &  x464 &  x473 &  x482 &  x497 &  x500 &  x512 &  x515 &  x530 &  x533 &  x536 &  x554 &  x557 &  x566 &  x572 &  x584 &  x608 &  x611 &  x614 &  x629 &  x632 &  x653 &  x674 &  x677 &  x686 &  x689 &  x692 &  x698 &  x701 &  x707 &  x713 &  x734 &  x740 &  x752 &  x755 &  x764 &  x770 &  x773 &  x776 &  x791 &  x794 &  x809 &  x827 &  x830 &  x833 &  x836 &  x845 &  x848 &  x890 &  x893 &  x896 &  x905 &  x914 &  x920 &  x923 &  x926 &  x935 &  x941 &  x944 &  x950 &  x953 &  x959 &  x968 &  x974 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1031 &  x1034 &  x1067 &  x1073 &  x1097 &  x1099 & ~x3 & ~x42 & ~x354 & ~x393 & ~x432 & ~x588 & ~x627;
assign c4163 =  x23 &  x26 &  x41 &  x50 &  x134 &  x187 &  x227 &  x286 &  x299 &  x395 &  x494 &  x539 &  x638 &  x662 &  x664 &  x674 &  x728 &  x731 &  x836 &  x839 &  x872 &  x886 &  x1019 &  x1049 & ~x831;
assign c4165 =  x131 &  x170 &  x365 &  x602 &  x628 &  x703 &  x706 &  x745 &  x781 &  x823 &  x901 &  x1018 & ~x513;
assign c4167 = ~x156 & ~x276 & ~x687 & ~x753 & ~x831 & ~x909 & ~x1026;
assign c4169 =  x20 &  x47 &  x56 &  x59 &  x80 &  x95 &  x98 &  x107 &  x116 &  x122 &  x125 &  x131 &  x152 &  x164 &  x191 &  x209 &  x227 &  x248 &  x254 &  x263 &  x269 &  x278 &  x290 &  x314 &  x329 &  x341 &  x350 &  x368 &  x374 &  x404 &  x406 &  x413 &  x416 &  x428 &  x446 &  x458 &  x467 &  x470 &  x497 &  x503 &  x512 &  x527 &  x530 &  x536 &  x545 &  x551 &  x590 &  x602 &  x635 &  x638 &  x662 &  x664 &  x665 &  x674 &  x683 &  x698 &  x707 &  x716 &  x737 &  x740 &  x749 &  x764 &  x773 &  x779 &  x782 &  x788 &  x803 &  x809 &  x818 &  x827 &  x839 &  x854 &  x872 &  x875 &  x878 &  x902 &  x908 &  x920 &  x950 &  x953 &  x959 &  x968 &  x974 &  x986 &  x995 &  x1019 &  x1052 &  x1061 &  x1073 &  x1082 &  x1091 &  x1103 & ~x315 & ~x351 & ~x630 & ~x792;
assign c4171 =  x13 &  x38 &  x50 &  x65 &  x91 &  x110 &  x130 &  x149 &  x299 &  x341 &  x365 &  x383 &  x461 &  x494 &  x524 &  x533 &  x545 &  x575 &  x605 &  x614 &  x623 &  x626 &  x635 &  x641 &  x695 &  x755 &  x773 &  x775 &  x791 &  x806 &  x841 &  x842 &  x860 &  x880 &  x935 &  x971 &  x980 &  x1028 &  x1055 &  x1061 &  x1100 &  x1127 & ~x594 & ~x828;
assign c4173 =  x101 &  x125 &  x149 &  x257 &  x428 &  x506 &  x542 &  x554 &  x623 &  x626 &  x674 &  x698 &  x710 &  x761 &  x842 &  x848 &  x860 &  x916 &  x938 &  x1001 &  x1019 & ~x402 & ~x441 & ~x480 & ~x519 & ~x636 & ~x702 & ~x822;
assign c4175 =  x2 &  x14 &  x17 &  x20 &  x29 &  x35 &  x38 &  x44 &  x47 &  x50 &  x53 &  x62 &  x65 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x107 &  x110 &  x122 &  x131 &  x143 &  x146 &  x170 &  x176 &  x191 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x233 &  x236 &  x242 &  x248 &  x251 &  x254 &  x260 &  x266 &  x272 &  x278 &  x284 &  x287 &  x302 &  x305 &  x308 &  x311 &  x317 &  x332 &  x335 &  x343 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x374 &  x389 &  x392 &  x398 &  x401 &  x410 &  x419 &  x422 &  x425 &  x431 &  x434 &  x437 &  x440 &  x443 &  x449 &  x461 &  x464 &  x467 &  x470 &  x482 &  x485 &  x497 &  x500 &  x503 &  x509 &  x521 &  x524 &  x530 &  x533 &  x539 &  x542 &  x545 &  x551 &  x554 &  x563 &  x569 &  x575 &  x578 &  x581 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x623 &  x626 &  x632 &  x635 &  x638 &  x644 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x689 &  x692 &  x698 &  x707 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x743 &  x746 &  x749 &  x752 &  x758 &  x767 &  x770 &  x776 &  x779 &  x785 &  x791 &  x794 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x824 &  x827 &  x833 &  x836 &  x839 &  x842 &  x851 &  x860 &  x863 &  x875 &  x878 &  x881 &  x884 &  x893 &  x902 &  x920 &  x923 &  x929 &  x932 &  x938 &  x941 &  x944 &  x953 &  x956 &  x962 &  x965 &  x980 &  x986 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1046 &  x1049 &  x1052 &  x1079 &  x1088 &  x1091 &  x1097 &  x1100 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x42 & ~x315 & ~x354 & ~x393 & ~x471 & ~x588 & ~x627 & ~x705 & ~x765;
assign c4177 =  x116 &  x155 &  x182 &  x302 &  x320 &  x377 &  x394 &  x404 &  x431 &  x461 &  x509 &  x512 &  x515 &  x539 &  x557 &  x571 &  x584 &  x638 &  x680 &  x728 &  x743 &  x800 &  x812 &  x850 &  x863 &  x884 &  x950 &  x961 &  x977 &  x980 &  x1000 &  x1022 &  x1028 &  x1031 &  x1058 &  x1085 & ~x561 & ~x600 & ~x639 & ~x663 & ~x780;
assign c4179 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x35 &  x41 &  x44 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x137 &  x140 &  x143 &  x146 &  x152 &  x155 &  x161 &  x166 &  x170 &  x173 &  x176 &  x179 &  x182 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x205 &  x206 &  x212 &  x215 &  x218 &  x221 &  x227 &  x233 &  x236 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x274 &  x275 &  x278 &  x283 &  x284 &  x287 &  x290 &  x293 &  x296 &  x302 &  x305 &  x308 &  x311 &  x313 &  x314 &  x317 &  x320 &  x322 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x356 &  x362 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x389 &  x391 &  x392 &  x395 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x422 &  x425 &  x430 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x469 &  x470 &  x473 &  x476 &  x479 &  x482 &  x488 &  x491 &  x494 &  x497 &  x500 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x545 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x608 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x680 &  x683 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x850 &  x851 &  x854 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x889 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x922 &  x923 &  x926 &  x928 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 &  x1130 & ~x318;
assign c4181 =  x17 &  x23 &  x35 &  x44 &  x53 &  x71 &  x80 &  x92 &  x95 &  x113 &  x122 &  x128 &  x176 &  x212 &  x224 &  x230 &  x233 &  x236 &  x263 &  x293 &  x359 &  x401 &  x413 &  x425 &  x488 &  x509 &  x548 &  x563 &  x593 &  x611 &  x632 &  x641 &  x706 &  x731 &  x745 &  x755 &  x800 &  x803 &  x806 &  x812 &  x815 &  x836 &  x839 &  x878 &  x914 &  x917 &  x923 &  x926 &  x929 &  x962 &  x989 &  x1001 &  x1019 &  x1027 &  x1043 &  x1067 &  x1073 &  x1079 &  x1085 &  x1094 &  x1124 & ~x639 & ~x678 & ~x897 & ~x936;
assign c4183 =  x5 &  x8 &  x11 &  x20 &  x29 &  x41 &  x68 &  x80 &  x89 &  x143 &  x164 &  x188 &  x203 &  x251 &  x254 &  x287 &  x320 &  x355 &  x383 &  x391 &  x410 &  x422 &  x425 &  x437 &  x449 &  x452 &  x473 &  x488 &  x533 &  x545 &  x554 &  x602 &  x605 &  x623 &  x641 &  x698 &  x713 &  x719 &  x749 &  x800 &  x824 &  x827 &  x854 &  x857 &  x866 &  x875 &  x887 &  x893 &  x899 &  x902 &  x908 &  x911 &  x971 &  x998 &  x1004 &  x1019 &  x1049 &  x1052 &  x1112 &  x1121 & ~x441 & ~x480 & ~x519 & ~x558 & ~x585 & ~x624 & ~x741 & ~x780 & ~x819 & ~x858;
assign c4185 =  x20 &  x44 &  x50 &  x119 &  x152 &  x167 &  x194 &  x209 &  x233 &  x242 &  x281 &  x305 &  x362 &  x365 &  x371 &  x374 &  x386 &  x401 &  x416 &  x428 &  x437 &  x472 &  x488 &  x491 &  x503 &  x515 &  x539 &  x548 &  x553 &  x578 &  x584 &  x596 &  x608 &  x626 &  x631 &  x650 &  x656 &  x665 &  x668 &  x688 &  x716 &  x767 &  x779 &  x827 &  x830 &  x854 &  x944 &  x968 &  x971 &  x974 &  x983 &  x998 &  x1031 &  x1046 &  x1058 &  x1085 &  x1106 &  x1121 & ~x522 & ~x663 & ~x741 & ~x936;
assign c4187 =  x812 &  x822 &  x982;
assign c4189 =  x14 &  x17 &  x41 &  x68 &  x77 &  x104 &  x134 &  x167 &  x226 &  x233 &  x260 &  x266 &  x275 &  x278 &  x304 &  x323 &  x455 &  x458 &  x461 &  x506 &  x533 &  x554 &  x599 &  x611 &  x614 &  x680 &  x683 &  x703 &  x737 &  x742 &  x755 &  x803 &  x820 &  x827 &  x836 &  x854 &  x902 &  x926 &  x962 &  x977 &  x1007 &  x1010 &  x1013 &  x1049 &  x1061 &  x1070 & ~x432 & ~x471 & ~x870 & ~x948 & ~x1026 & ~x1065;
assign c4191 =  x44 &  x77 &  x161 &  x188 &  x284 &  x374 &  x521 &  x566 &  x608 &  x617 &  x691 &  x701 &  x782 &  x806 &  x818 &  x827 &  x890 &  x917 &  x971 &  x989 &  x1027 &  x1037 &  x1049 & ~x477 & ~x522 & ~x594 & ~x600 & ~x702 & ~x897;
assign c4193 =  x26 &  x35 &  x71 &  x80 &  x86 &  x89 &  x91 &  x113 &  x128 &  x158 &  x161 &  x167 &  x209 &  x269 &  x322 &  x323 &  x329 &  x344 &  x347 &  x350 &  x440 &  x446 &  x452 &  x455 &  x461 &  x473 &  x488 &  x491 &  x494 &  x506 &  x536 &  x539 &  x548 &  x584 &  x593 &  x650 &  x671 &  x689 &  x698 &  x719 &  x728 &  x773 &  x776 &  x779 &  x794 &  x830 &  x833 &  x854 &  x878 &  x887 &  x899 &  x923 &  x947 &  x950 &  x995 &  x1001 &  x1022 &  x1028 &  x1034 &  x1046 &  x1061 &  x1073 &  x1076 &  x1079 &  x1127 & ~x264 & ~x624 & ~x702 & ~x819 & ~x858 & ~x1047;
assign c4195 =  x53 &  x71 &  x197 &  x200 &  x338 &  x353 &  x438 &  x478 &  x508 &  x704 &  x860 &  x875 & ~x237 & ~x513;
assign c4197 =  x217 &  x322 &  x852 &  x1048 & ~x906;
assign c4199 =  x8 &  x26 &  x38 &  x41 &  x62 &  x65 &  x68 &  x89 &  x95 &  x101 &  x110 &  x128 &  x152 &  x155 &  x167 &  x197 &  x212 &  x224 &  x242 &  x245 &  x248 &  x260 &  x263 &  x269 &  x278 &  x293 &  x296 &  x305 &  x317 &  x323 &  x326 &  x337 &  x338 &  x350 &  x356 &  x437 &  x455 &  x458 &  x461 &  x467 &  x473 &  x509 &  x521 &  x545 &  x554 &  x559 &  x560 &  x563 &  x565 &  x581 &  x584 &  x598 &  x608 &  x620 &  x632 &  x635 &  x637 &  x671 &  x712 &  x737 &  x740 &  x751 &  x767 &  x794 &  x800 &  x830 &  x833 &  x848 &  x854 &  x857 &  x863 &  x887 &  x908 &  x941 &  x950 &  x959 &  x962 &  x968 &  x974 &  x998 &  x1001 &  x1019 &  x1028 &  x1040 &  x1046 &  x1064 &  x1073 &  x1082 &  x1097 &  x1112 & ~x354 & ~x837;
assign c4201 =  x371 &  x743 &  x998 &  x1018 &  x1052 & ~x390 & ~x669 & ~x831 & ~x951;
assign c4203 =  x116 &  x233 &  x338 &  x413 & ~x3 & ~x174 & ~x516 & ~x633 & ~x750 & ~x780 & ~x897;
assign c4205 =  x661 &  x816 &  x877 & ~x441;
assign c4207 =  x29 &  x77 &  x83 &  x98 &  x101 &  x113 &  x122 &  x149 &  x164 &  x176 &  x215 &  x218 &  x290 &  x320 &  x365 &  x410 &  x416 &  x443 &  x476 &  x482 &  x518 &  x587 &  x710 &  x742 &  x761 &  x767 &  x800 &  x857 &  x863 &  x950 &  x974 &  x980 &  x1019 &  x1028 &  x1058 &  x1115 &  x1121 & ~x351 & ~x432 & ~x792 & ~x870 & ~x948 & ~x1065;
assign c4209 =  x2 &  x44 &  x83 &  x95 &  x101 &  x110 &  x119 &  x131 &  x169 &  x173 &  x179 &  x197 &  x209 &  x263 &  x266 &  x269 &  x272 &  x286 &  x296 &  x305 &  x335 &  x362 &  x374 &  x383 &  x404 &  x419 &  x467 &  x500 &  x506 &  x509 &  x521 &  x530 &  x542 &  x554 &  x578 &  x584 &  x586 &  x617 &  x620 &  x623 &  x625 &  x629 &  x647 &  x680 &  x701 &  x716 &  x719 &  x722 &  x737 &  x743 &  x779 &  x785 &  x818 &  x848 &  x854 &  x857 &  x863 &  x878 &  x890 &  x905 &  x908 &  x965 &  x974 &  x1013 &  x1022 &  x1043 &  x1061 &  x1085 &  x1097 &  x1100 &  x1124 &  x1127 & ~x636 & ~x714 & ~x831 & ~x870 & ~x909;
assign c4211 = ~x679;
assign c4213 =  x77 &  x113 &  x703 &  x1085 & ~x471 & ~x871 & ~x910 & ~x1065;
assign c4215 =  x17 &  x29 &  x32 &  x44 &  x74 &  x77 &  x80 &  x86 &  x122 &  x131 &  x140 &  x143 &  x167 &  x176 &  x212 &  x215 &  x242 &  x245 &  x254 &  x257 &  x266 &  x308 &  x353 &  x362 &  x365 &  x368 &  x392 &  x398 &  x422 &  x430 &  x434 &  x458 &  x464 &  x469 &  x488 &  x508 &  x511 &  x518 &  x539 &  x550 &  x560 &  x566 &  x569 &  x572 &  x587 &  x589 &  x599 &  x602 &  x608 &  x650 &  x653 &  x695 &  x709 &  x716 &  x758 &  x779 &  x800 &  x806 &  x818 &  x851 &  x854 &  x884 &  x893 &  x917 &  x956 &  x965 &  x971 &  x1001 &  x1004 &  x1037 &  x1040 &  x1049 &  x1058 &  x1064 &  x1082 &  x1091 &  x1100 &  x1103 &  x1118 &  x1124 &  x1130 & ~x597 & ~x675;
assign c4217 =  x92 &  x104 &  x188 &  x311 &  x356 &  x374 &  x416 &  x527 &  x557 &  x560 &  x566 &  x605 &  x641 &  x665 &  x683 &  x703 &  x713 &  x752 &  x776 &  x809 &  x815 &  x863 &  x896 &  x902 &  x944 &  x986 &  x1001 &  x1031 &  x1076 &  x1100 & ~x39 & ~x156 & ~x195 & ~x354 & ~x432 & ~x510 & ~x588;
assign c4219 =  x451 &  x502 &  x856 & ~x651;
assign c4221 =  x59 &  x490 &  x748 &  x869 &  x884 &  x892 &  x895 &  x1076 &  x1088 &  x1103 &  x1115 & ~x675;
assign c4223 =  x149 &  x164 &  x230 &  x281 &  x497 &  x653 &  x742 &  x797 &  x848 &  x896 &  x950 & ~x243 & ~x351 & ~x390 & ~x432 & ~x588 & ~x708;
assign c4225 =  x284 &  x625 &  x629 &  x734 &  x752 & ~x237 & ~x276 & ~x315 & ~x393 & ~x552;
assign c4227 =  x8 &  x257 &  x311 &  x485 &  x797 &  x806 & ~x246 & ~x402 & ~x480 & ~x519 & ~x585 & ~x873 & ~x951 & ~x1062;
assign c4229 =  x218 &  x310 &  x389 &  x695 &  x748 &  x806 &  x992 &  x1027 & ~x639 & ~x858 & ~x936;
assign c4231 = ~x221;
assign c4233 =  x2 &  x5 &  x11 &  x17 &  x20 &  x29 &  x35 &  x38 &  x44 &  x47 &  x50 &  x53 &  x62 &  x68 &  x71 &  x74 &  x77 &  x86 &  x89 &  x92 &  x95 &  x101 &  x113 &  x116 &  x122 &  x125 &  x131 &  x134 &  x137 &  x140 &  x143 &  x158 &  x164 &  x170 &  x176 &  x182 &  x185 &  x188 &  x194 &  x203 &  x209 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x242 &  x245 &  x251 &  x257 &  x263 &  x266 &  x269 &  x271 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x299 &  x302 &  x308 &  x310 &  x311 &  x320 &  x326 &  x329 &  x332 &  x338 &  x341 &  x344 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x377 &  x379 &  x380 &  x383 &  x386 &  x395 &  x398 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x437 &  x440 &  x449 &  x452 &  x455 &  x464 &  x473 &  x476 &  x488 &  x491 &  x494 &  x497 &  x506 &  x512 &  x518 &  x527 &  x533 &  x536 &  x545 &  x548 &  x554 &  x560 &  x566 &  x569 &  x575 &  x578 &  x584 &  x590 &  x596 &  x611 &  x614 &  x617 &  x620 &  x641 &  x644 &  x647 &  x650 &  x659 &  x665 &  x668 &  x671 &  x674 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x710 &  x713 &  x719 &  x722 &  x728 &  x731 &  x737 &  x746 &  x755 &  x758 &  x764 &  x770 &  x776 &  x779 &  x782 &  x785 &  x791 &  x794 &  x797 &  x800 &  x809 &  x812 &  x815 &  x821 &  x827 &  x830 &  x839 &  x848 &  x851 &  x854 &  x857 &  x860 &  x869 &  x872 &  x878 &  x887 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x917 &  x920 &  x929 &  x935 &  x938 &  x941 &  x944 &  x953 &  x956 &  x977 &  x986 &  x989 &  x992 &  x995 &  x1004 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1061 &  x1067 &  x1076 &  x1079 &  x1082 &  x1085 &  x1094 &  x1097 &  x1100 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x393 & ~x471 & ~x510 & ~x909 & ~x948 & ~x1026 & ~x1065 & ~x1104;
assign c4235 =  x2 &  x41 &  x71 &  x77 &  x92 &  x125 &  x166 &  x205 &  x221 &  x244 &  x313 &  x316 &  x335 &  x509 &  x548 &  x626 &  x644 &  x683 &  x698 &  x704 &  x761 &  x824 &  x857 &  x866 &  x872 &  x947 &  x986 &  x1064 & ~x483 & ~x585 & ~x702 & ~x780 & ~x819;
assign c4237 =  x11 &  x47 &  x137 &  x329 &  x422 &  x434 &  x533 &  x571 &  x740 &  x817 &  x856 & ~x148 & ~x246;
assign c4239 =  x648 & ~x976;
assign c4241 =  x8 &  x20 &  x35 &  x44 &  x68 &  x80 &  x89 &  x116 &  x122 &  x146 &  x200 &  x212 &  x227 &  x233 &  x260 &  x317 &  x374 &  x431 &  x599 &  x635 &  x641 &  x722 &  x728 &  x761 &  x779 &  x803 &  x818 &  x887 &  x914 &  x950 &  x953 &  x962 &  x977 &  x1042 &  x1055 &  x1073 &  x1088 &  x1100 &  x1127 & ~x276 & ~x591 & ~x753 & ~x792;
assign c4243 =  x502 & ~x597 & ~x793;
assign c4245 =  x508 &  x589 &  x685 &  x763 &  x1111 & ~x675;
assign c4247 =  x2 &  x5 &  x8 &  x14 &  x23 &  x29 &  x32 &  x44 &  x62 &  x74 &  x80 &  x83 &  x89 &  x101 &  x131 &  x137 &  x149 &  x152 &  x158 &  x161 &  x170 &  x173 &  x176 &  x179 &  x182 &  x191 &  x194 &  x200 &  x203 &  x206 &  x209 &  x218 &  x224 &  x227 &  x254 &  x266 &  x269 &  x272 &  x284 &  x287 &  x293 &  x308 &  x320 &  x323 &  x332 &  x341 &  x344 &  x353 &  x359 &  x365 &  x377 &  x395 &  x398 &  x407 &  x413 &  x416 &  x440 &  x461 &  x464 &  x473 &  x479 &  x485 &  x497 &  x515 &  x518 &  x521 &  x524 &  x530 &  x542 &  x548 &  x551 &  x557 &  x578 &  x587 &  x595 &  x596 &  x617 &  x623 &  x634 &  x644 &  x656 &  x665 &  x668 &  x673 &  x674 &  x686 &  x692 &  x703 &  x704 &  x719 &  x737 &  x740 &  x742 &  x746 &  x751 &  x755 &  x758 &  x764 &  x776 &  x779 &  x785 &  x800 &  x815 &  x818 &  x821 &  x824 &  x830 &  x833 &  x839 &  x842 &  x845 &  x851 &  x854 &  x860 &  x872 &  x881 &  x902 &  x905 &  x908 &  x911 &  x914 &  x929 &  x944 &  x950 &  x953 &  x959 &  x974 &  x977 &  x986 &  x992 &  x995 &  x1007 &  x1010 &  x1013 &  x1016 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1046 &  x1049 &  x1058 &  x1061 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1100 &  x1106 &  x1112 &  x1118 &  x1121 &  x1127 &  x1130 & ~x432 & ~x471 & ~x732 & ~x771;
assign c4249 = ~x549 & ~x871 & ~x912 & ~x1068;
assign c4251 =  x35 &  x71 &  x116 &  x137 &  x152 &  x182 &  x251 &  x272 &  x281 &  x329 &  x380 &  x443 &  x512 &  x515 &  x554 &  x563 &  x626 &  x629 &  x722 &  x800 &  x806 &  x815 &  x902 &  x917 &  x965 & ~x234 & ~x276 & ~x471 & ~x909 & ~x954 & ~x987 & ~x1065 & ~x1104;
assign c4253 =  x8 &  x14 &  x17 &  x23 &  x32 &  x41 &  x50 &  x53 &  x74 &  x86 &  x92 &  x95 &  x98 &  x107 &  x110 &  x116 &  x122 &  x140 &  x146 &  x155 &  x164 &  x182 &  x197 &  x206 &  x215 &  x224 &  x230 &  x233 &  x236 &  x239 &  x242 &  x248 &  x281 &  x284 &  x290 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x323 &  x326 &  x332 &  x335 &  x355 &  x356 &  x362 &  x386 &  x401 &  x413 &  x422 &  x428 &  x436 &  x440 &  x443 &  x446 &  x461 &  x464 &  x467 &  x473 &  x475 &  x476 &  x479 &  x488 &  x494 &  x521 &  x527 &  x536 &  x545 &  x548 &  x553 &  x560 &  x569 &  x578 &  x581 &  x584 &  x602 &  x605 &  x611 &  x614 &  x617 &  x632 &  x635 &  x637 &  x638 &  x641 &  x656 &  x662 &  x670 &  x676 &  x680 &  x683 &  x686 &  x695 &  x698 &  x704 &  x709 &  x710 &  x713 &  x715 &  x725 &  x731 &  x740 &  x746 &  x752 &  x758 &  x770 &  x773 &  x785 &  x803 &  x812 &  x818 &  x821 &  x830 &  x839 &  x857 &  x863 &  x890 &  x899 &  x905 &  x911 &  x932 &  x938 &  x941 &  x950 &  x971 &  x977 &  x980 &  x1004 &  x1010 &  x1019 &  x1028 &  x1040 &  x1052 &  x1058 &  x1067 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1100 &  x1103 &  x1109 &  x1112 &  x1124 &  x1130 & ~x405 & ~x585 & ~x624 & ~x702 & ~x744 & ~x822;
assign c4255 =  x1012 & ~x81 & ~x198 & ~x315 & ~x432 & ~x642;
assign c4257 =  x8 &  x59 &  x209 &  x224 &  x290 &  x329 &  x419 &  x431 &  x503 &  x506 &  x557 &  x608 &  x659 &  x695 &  x709 &  x776 &  x797 &  x890 &  x902 &  x911 &  x938 &  x944 &  x1070 &  x1117 & ~x522 & ~x562 & ~x678;
assign c4259 =  x38 &  x62 &  x68 &  x149 &  x166 &  x173 &  x185 &  x248 &  x251 &  x413 &  x462 &  x463 &  x540 &  x602 &  x605 &  x617 &  x707 &  x776 &  x818 &  x881 &  x917 &  x944 &  x989 &  x1016 &  x1106 & ~x318 & ~x744;
assign c4261 =  x8 &  x14 &  x26 &  x44 &  x53 &  x62 &  x65 &  x68 &  x86 &  x92 &  x101 &  x104 &  x125 &  x134 &  x137 &  x143 &  x146 &  x161 &  x170 &  x179 &  x182 &  x185 &  x188 &  x191 &  x197 &  x206 &  x221 &  x233 &  x242 &  x245 &  x248 &  x257 &  x260 &  x266 &  x296 &  x299 &  x305 &  x308 &  x323 &  x326 &  x329 &  x341 &  x353 &  x368 &  x371 &  x374 &  x380 &  x386 &  x389 &  x398 &  x407 &  x425 &  x437 &  x440 &  x443 &  x452 &  x458 &  x467 &  x470 &  x476 &  x479 &  x509 &  x518 &  x527 &  x539 &  x548 &  x572 &  x578 &  x584 &  x593 &  x596 &  x611 &  x619 &  x620 &  x629 &  x638 &  x647 &  x650 &  x659 &  x665 &  x674 &  x680 &  x686 &  x697 &  x698 &  x701 &  x704 &  x707 &  x710 &  x716 &  x725 &  x731 &  x734 &  x736 &  x737 &  x743 &  x749 &  x755 &  x764 &  x767 &  x773 &  x775 &  x776 &  x800 &  x803 &  x809 &  x812 &  x821 &  x836 &  x842 &  x845 &  x848 &  x851 &  x857 &  x863 &  x872 &  x878 &  x881 &  x884 &  x887 &  x898 &  x902 &  x905 &  x914 &  x926 &  x929 &  x937 &  x944 &  x947 &  x962 &  x980 &  x983 &  x989 &  x1001 &  x1004 &  x1013 &  x1016 &  x1034 &  x1037 &  x1040 &  x1043 &  x1052 &  x1064 &  x1070 &  x1088 &  x1091 &  x1097 &  x1106 &  x1115 &  x1127 &  x1130 & ~x597 & ~x675 & ~x792 & ~x909 & ~x948;
assign c4263 =  x83 &  x131 &  x191 &  x203 &  x245 &  x302 &  x344 &  x377 &  x380 &  x404 &  x470 &  x473 &  x521 &  x547 &  x746 &  x791 &  x800 &  x884 &  x971 &  x1007 &  x1018 &  x1097 & ~x636 & ~x675 & ~x714 & ~x756 & ~x792;
assign c4265 = ~x258 & ~x714 & ~x871 & ~x948;
assign c4267 =  x113 &  x212 &  x422 &  x586 &  x625 &  x731 &  x761 &  x929 &  x998 &  x1001 &  x1124 & ~x39 & ~x315 & ~x432 & ~x792 & ~x831;
assign c4269 =  x745 & ~x718 & ~x897;
assign c4271 =  x5 &  x14 &  x20 &  x23 &  x35 &  x44 &  x59 &  x62 &  x86 &  x89 &  x92 &  x113 &  x122 &  x146 &  x167 &  x173 &  x182 &  x185 &  x194 &  x200 &  x203 &  x209 &  x212 &  x238 &  x239 &  x272 &  x274 &  x278 &  x313 &  x316 &  x341 &  x419 &  x434 &  x440 &  x475 &  x482 &  x488 &  x514 &  x515 &  x521 &  x533 &  x542 &  x548 &  x560 &  x563 &  x569 &  x575 &  x587 &  x593 &  x596 &  x608 &  x614 &  x620 &  x631 &  x635 &  x637 &  x641 &  x676 &  x677 &  x683 &  x692 &  x704 &  x719 &  x749 &  x767 &  x779 &  x782 &  x791 &  x806 &  x809 &  x812 &  x836 &  x860 &  x863 &  x869 &  x881 &  x896 &  x917 &  x938 &  x959 &  x971 &  x974 &  x983 &  x989 &  x995 &  x1004 &  x1013 &  x1046 &  x1049 &  x1061 &  x1070 &  x1076 &  x1097 &  x1103 &  x1121 & ~x366 & ~x585 & ~x861;
assign c4273 =  x2 &  x14 &  x35 &  x47 &  x56 &  x59 &  x62 &  x71 &  x83 &  x86 &  x95 &  x98 &  x110 &  x113 &  x116 &  x164 &  x182 &  x185 &  x188 &  x194 &  x197 &  x206 &  x215 &  x224 &  x275 &  x290 &  x302 &  x305 &  x311 &  x314 &  x335 &  x350 &  x362 &  x383 &  x392 &  x401 &  x416 &  x431 &  x449 &  x452 &  x458 &  x467 &  x470 &  x476 &  x482 &  x500 &  x518 &  x524 &  x542 &  x545 &  x551 &  x560 &  x569 &  x572 &  x581 &  x587 &  x590 &  x593 &  x620 &  x626 &  x635 &  x638 &  x641 &  x656 &  x662 &  x667 &  x671 &  x677 &  x686 &  x698 &  x701 &  x704 &  x716 &  x719 &  x725 &  x740 &  x746 &  x752 &  x767 &  x770 &  x773 &  x784 &  x785 &  x788 &  x791 &  x800 &  x803 &  x812 &  x818 &  x821 &  x833 &  x836 &  x845 &  x851 &  x854 &  x857 &  x860 &  x863 &  x865 &  x872 &  x881 &  x884 &  x887 &  x899 &  x905 &  x908 &  x911 &  x932 &  x938 &  x941 &  x950 &  x953 &  x959 &  x968 &  x971 &  x974 &  x989 &  x992 &  x998 &  x1007 &  x1016 &  x1019 &  x1022 &  x1025 &  x1037 &  x1040 &  x1055 &  x1058 &  x1076 &  x1079 &  x1085 &  x1115 &  x1121 & ~x756 & ~x795 & ~x798;
assign c4275 =  x5 &  x13 &  x51 &  x113 &  x149 &  x173 &  x179 &  x281 &  x410 &  x467 &  x482 &  x491 &  x524 &  x812 &  x857 &  x872 &  x923 &  x959 &  x1027 & ~x702 & ~x780 & ~x819 & ~x858;
assign c4277 =  x2 &  x8 &  x11 &  x23 &  x26 &  x29 &  x32 &  x38 &  x44 &  x47 &  x50 &  x53 &  x56 &  x77 &  x83 &  x86 &  x104 &  x110 &  x116 &  x119 &  x122 &  x125 &  x128 &  x137 &  x140 &  x143 &  x152 &  x161 &  x164 &  x166 &  x167 &  x170 &  x194 &  x197 &  x200 &  x203 &  x209 &  x212 &  x221 &  x230 &  x242 &  x248 &  x251 &  x266 &  x275 &  x281 &  x302 &  x305 &  x314 &  x320 &  x323 &  x329 &  x332 &  x341 &  x350 &  x352 &  x365 &  x368 &  x371 &  x377 &  x383 &  x389 &  x391 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x431 &  x440 &  x449 &  x476 &  x479 &  x500 &  x506 &  x524 &  x533 &  x536 &  x542 &  x545 &  x554 &  x560 &  x563 &  x569 &  x575 &  x578 &  x581 &  x599 &  x605 &  x617 &  x620 &  x623 &  x626 &  x635 &  x644 &  x650 &  x653 &  x659 &  x683 &  x692 &  x701 &  x707 &  x716 &  x722 &  x731 &  x734 &  x737 &  x743 &  x749 &  x758 &  x761 &  x764 &  x770 &  x773 &  x779 &  x782 &  x788 &  x794 &  x797 &  x806 &  x818 &  x827 &  x830 &  x836 &  x842 &  x845 &  x848 &  x851 &  x854 &  x860 &  x869 &  x872 &  x878 &  x887 &  x902 &  x905 &  x923 &  x941 &  x944 &  x947 &  x962 &  x965 &  x968 &  x974 &  x980 &  x983 &  x989 &  x995 &  x998 &  x1007 &  x1016 &  x1022 &  x1025 &  x1034 &  x1040 &  x1046 &  x1052 &  x1058 &  x1070 &  x1073 &  x1088 &  x1100 &  x1103 &  x1109 &  x1112 &  x1118 &  x1121 &  x1130 & ~x330 & ~x477 & ~x516 & ~x555 & ~x633 & ~x672 & ~x702;
assign c4279 =  x2 &  x5 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x50 &  x53 &  x56 &  x59 &  x65 &  x71 &  x77 &  x80 &  x86 &  x89 &  x92 &  x101 &  x113 &  x116 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x143 &  x146 &  x149 &  x158 &  x161 &  x164 &  x170 &  x179 &  x191 &  x197 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x230 &  x233 &  x239 &  x242 &  x248 &  x251 &  x257 &  x263 &  x266 &  x269 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x299 &  x302 &  x305 &  x308 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x365 &  x371 &  x380 &  x383 &  x389 &  x392 &  x395 &  x398 &  x404 &  x407 &  x410 &  x413 &  x428 &  x434 &  x437 &  x440 &  x443 &  x446 &  x455 &  x458 &  x461 &  x467 &  x479 &  x482 &  x485 &  x491 &  x494 &  x497 &  x500 &  x512 &  x514 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x554 &  x560 &  x563 &  x572 &  x575 &  x584 &  x590 &  x596 &  x599 &  x608 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x656 &  x659 &  x665 &  x668 &  x674 &  x680 &  x683 &  x686 &  x695 &  x698 &  x707 &  x710 &  x716 &  x722 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x779 &  x782 &  x785 &  x788 &  x791 &  x797 &  x800 &  x806 &  x809 &  x818 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x845 &  x848 &  x854 &  x857 &  x863 &  x875 &  x878 &  x884 &  x887 &  x890 &  x896 &  x899 &  x905 &  x908 &  x911 &  x920 &  x923 &  x926 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x968 &  x971 &  x974 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1013 &  x1019 &  x1022 &  x1025 &  x1028 &  x1034 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1058 &  x1060 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1082 &  x1085 &  x1091 &  x1094 &  x1097 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x3 & ~x42 & ~x81 & ~x588 & ~x627;
assign c4281 =  x8 &  x11 &  x14 &  x17 &  x23 &  x32 &  x38 &  x41 &  x47 &  x50 &  x56 &  x59 &  x62 &  x80 &  x83 &  x86 &  x89 &  x98 &  x104 &  x107 &  x116 &  x122 &  x137 &  x143 &  x146 &  x149 &  x158 &  x164 &  x170 &  x179 &  x182 &  x185 &  x188 &  x191 &  x197 &  x209 &  x212 &  x214 &  x221 &  x224 &  x239 &  x242 &  x245 &  x248 &  x251 &  x253 &  x254 &  x257 &  x263 &  x266 &  x269 &  x275 &  x281 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x311 &  x317 &  x320 &  x323 &  x326 &  x329 &  x335 &  x341 &  x344 &  x353 &  x365 &  x368 &  x380 &  x389 &  x392 &  x398 &  x401 &  x404 &  x407 &  x409 &  x410 &  x416 &  x419 &  x422 &  x437 &  x443 &  x446 &  x448 &  x449 &  x458 &  x461 &  x464 &  x467 &  x470 &  x479 &  x482 &  x485 &  x494 &  x503 &  x506 &  x509 &  x524 &  x527 &  x542 &  x551 &  x554 &  x557 &  x563 &  x566 &  x569 &  x575 &  x584 &  x587 &  x593 &  x599 &  x605 &  x608 &  x611 &  x623 &  x626 &  x629 &  x632 &  x635 &  x650 &  x653 &  x656 &  x662 &  x671 &  x677 &  x680 &  x695 &  x698 &  x703 &  x710 &  x713 &  x716 &  x719 &  x728 &  x731 &  x734 &  x737 &  x740 &  x742 &  x743 &  x749 &  x752 &  x773 &  x776 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x803 &  x809 &  x812 &  x818 &  x830 &  x836 &  x842 &  x845 &  x848 &  x854 &  x863 &  x869 &  x878 &  x884 &  x890 &  x896 &  x899 &  x902 &  x904 &  x905 &  x908 &  x911 &  x920 &  x926 &  x929 &  x935 &  x938 &  x947 &  x950 &  x953 &  x956 &  x962 &  x965 &  x968 &  x971 &  x977 &  x983 &  x986 &  x995 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1037 &  x1043 &  x1046 &  x1049 &  x1055 &  x1073 &  x1085 &  x1088 &  x1091 &  x1094 &  x1112 &  x1127 & ~x471;
assign c4283 =  x354 &  x475 &  x592 & ~x522;
assign c4285 =  x38 &  x362 &  x551 &  x584 &  x833 &  x859 &  x940 &  x1018 & ~x870 & ~x1065;
assign c4287 =  x373 &  x383 &  x477 &  x547 &  x548 &  x556 &  x625 &  x1037 & ~x219;
assign c4289 =  x2 &  x5 &  x11 &  x17 &  x23 &  x29 &  x32 &  x35 &  x38 &  x44 &  x50 &  x56 &  x62 &  x71 &  x74 &  x80 &  x83 &  x86 &  x89 &  x95 &  x107 &  x110 &  x113 &  x116 &  x122 &  x125 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x188 &  x191 &  x194 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x227 &  x233 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x266 &  x272 &  x278 &  x281 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x308 &  x317 &  x320 &  x323 &  x329 &  x332 &  x341 &  x344 &  x350 &  x353 &  x362 &  x371 &  x374 &  x377 &  x391 &  x392 &  x401 &  x404 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x431 &  x434 &  x437 &  x440 &  x449 &  x452 &  x455 &  x458 &  x461 &  x470 &  x473 &  x476 &  x479 &  x482 &  x488 &  x491 &  x497 &  x503 &  x506 &  x509 &  x515 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x545 &  x548 &  x554 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x581 &  x587 &  x590 &  x596 &  x599 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x644 &  x647 &  x650 &  x653 &  x656 &  x662 &  x668 &  x671 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x713 &  x716 &  x722 &  x731 &  x734 &  x737 &  x740 &  x743 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x779 &  x785 &  x791 &  x794 &  x797 &  x800 &  x812 &  x815 &  x818 &  x821 &  x824 &  x836 &  x839 &  x845 &  x851 &  x860 &  x869 &  x872 &  x875 &  x878 &  x881 &  x890 &  x896 &  x902 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x935 &  x944 &  x947 &  x950 &  x953 &  x962 &  x965 &  x968 &  x971 &  x974 &  x980 &  x983 &  x986 &  x992 &  x995 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1052 &  x1055 &  x1058 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x441 & ~x453 & ~x480 & ~x519 & ~x558 & ~x675 & ~x714 & ~x780 & ~x819;
assign c4291 =  x379 &  x436 &  x478 &  x555;
assign c4293 =  x2 &  x14 &  x20 &  x50 &  x59 &  x92 &  x104 &  x125 &  x149 &  x176 &  x197 &  x200 &  x230 &  x260 &  x293 &  x314 &  x320 &  x335 &  x389 &  x410 &  x413 &  x431 &  x476 &  x485 &  x494 &  x500 &  x511 &  x535 &  x632 &  x647 &  x650 &  x653 &  x659 &  x677 &  x683 &  x695 &  x709 &  x713 &  x716 &  x722 &  x767 &  x770 &  x826 &  x848 &  x866 &  x878 &  x883 &  x887 &  x890 &  x893 &  x902 &  x908 &  x929 &  x947 &  x949 &  x959 &  x968 &  x971 &  x980 &  x992 &  x1007 &  x1016 &  x1037 &  x1043 &  x1070 &  x1082 &  x1085 &  x1109 &  x1112 &  x1115 & ~x444 & ~x702 & ~x741 & ~x819;
assign c4295 =  x47 &  x50 &  x77 &  x83 &  x140 &  x197 &  x218 &  x224 &  x269 &  x281 &  x425 &  x629 &  x737 &  x884 &  x899 &  x977 &  x994 &  x1013 &  x1016 &  x1031 &  x1097 & ~x246 & ~x324 & ~x441 & ~x480 & ~x507 & ~x585 & ~x741 & ~x780 & ~x819 & ~x897 & ~x975;
assign c4297 =  x152 &  x482 &  x533 &  x632 &  x638 &  x744 &  x887 &  x904 &  x932 &  x1007 &  x1010 &  x1088 &  x1105;
assign c4299 =  x1018 & ~x474 & ~x640;
assign c50 =  x2 &  x8 &  x11 &  x14 &  x20 &  x23 &  x32 &  x38 &  x44 &  x47 &  x53 &  x59 &  x62 &  x68 &  x77 &  x80 &  x83 &  x95 &  x98 &  x101 &  x107 &  x110 &  x113 &  x119 &  x125 &  x128 &  x131 &  x137 &  x140 &  x146 &  x149 &  x152 &  x158 &  x161 &  x170 &  x173 &  x176 &  x185 &  x191 &  x203 &  x206 &  x209 &  x224 &  x227 &  x242 &  x251 &  x254 &  x269 &  x302 &  x314 &  x317 &  x329 &  x356 &  x365 &  x368 &  x371 &  x380 &  x383 &  x392 &  x395 &  x397 &  x401 &  x410 &  x431 &  x436 &  x440 &  x452 &  x455 &  x461 &  x464 &  x467 &  x470 &  x476 &  x482 &  x488 &  x491 &  x494 &  x509 &  x512 &  x515 &  x518 &  x521 &  x530 &  x533 &  x542 &  x545 &  x548 &  x551 &  x557 &  x566 &  x569 &  x578 &  x580 &  x581 &  x587 &  x590 &  x596 &  x605 &  x608 &  x611 &  x617 &  x623 &  x629 &  x632 &  x635 &  x641 &  x644 &  x650 &  x653 &  x656 &  x659 &  x668 &  x674 &  x677 &  x680 &  x689 &  x692 &  x695 &  x719 &  x740 &  x743 &  x746 &  x755 &  x767 &  x770 &  x781 &  x785 &  x788 &  x791 &  x806 &  x821 &  x827 &  x842 &  x848 &  x869 &  x872 &  x875 &  x890 &  x896 &  x902 &  x905 &  x908 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x938 &  x940 &  x941 &  x959 &  x965 &  x971 &  x974 &  x983 &  x986 &  x998 &  x1004 &  x1010 &  x1022 &  x1025 &  x1028 &  x1034 &  x1043 &  x1046 &  x1055 &  x1058 &  x1070 &  x1073 &  x1076 &  x1088 &  x1091 &  x1097 &  x1115 &  x1127 &  x1130 & ~x9 & ~x48 & ~x87 & ~x315 & ~x558 & ~x597 & ~x636 & ~x675 & ~x714 & ~x870 & ~x909;
assign c52 =  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x29 &  x32 &  x38 &  x40 &  x47 &  x50 &  x53 &  x59 &  x68 &  x71 &  x79 &  x86 &  x92 &  x98 &  x101 &  x116 &  x118 &  x119 &  x131 &  x134 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x167 &  x170 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x206 &  x215 &  x221 &  x230 &  x235 &  x236 &  x242 &  x245 &  x248 &  x254 &  x257 &  x266 &  x269 &  x272 &  x275 &  x278 &  x284 &  x287 &  x290 &  x293 &  x299 &  x308 &  x311 &  x313 &  x314 &  x317 &  x326 &  x332 &  x335 &  x338 &  x347 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x377 &  x383 &  x386 &  x389 &  x392 &  x394 &  x398 &  x401 &  x407 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x446 &  x452 &  x461 &  x464 &  x473 &  x479 &  x482 &  x488 &  x494 &  x497 &  x503 &  x506 &  x512 &  x524 &  x527 &  x533 &  x542 &  x548 &  x551 &  x563 &  x569 &  x571 &  x581 &  x584 &  x590 &  x593 &  x596 &  x602 &  x605 &  x611 &  x623 &  x629 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x659 &  x665 &  x668 &  x677 &  x680 &  x686 &  x689 &  x695 &  x716 &  x728 &  x731 &  x734 &  x737 &  x740 &  x749 &  x755 &  x770 &  x773 &  x782 &  x791 &  x794 &  x797 &  x803 &  x809 &  x815 &  x824 &  x830 &  x836 &  x839 &  x844 &  x848 &  x854 &  x857 &  x881 &  x884 &  x890 &  x893 &  x896 &  x899 &  x902 &  x908 &  x911 &  x917 &  x920 &  x923 &  x929 &  x935 &  x938 &  x941 &  x953 &  x968 &  x971 &  x974 &  x986 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1055 &  x1061 &  x1064 &  x1070 &  x1073 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1103 &  x1109 &  x1112 &  x1121 &  x1124 &  x1127 & ~x4 & ~x42 & ~x213 & ~x252 & ~x291 & ~x405 & ~x444 & ~x585 & ~x624 & ~x663 & ~x702 & ~x741 & ~x744 & ~x780 & ~x819 & ~x822 & ~x858 & ~x897;
assign c54 =  x11 &  x17 &  x20 &  x26 &  x35 &  x47 &  x53 &  x80 &  x89 &  x92 &  x95 &  x101 &  x155 &  x173 &  x179 &  x197 &  x206 &  x239 &  x242 &  x266 &  x293 &  x314 &  x335 &  x338 &  x362 &  x368 &  x380 &  x386 &  x395 &  x440 &  x452 &  x464 &  x482 &  x494 &  x521 &  x524 &  x533 &  x548 &  x551 &  x590 &  x593 &  x599 &  x602 &  x620 &  x623 &  x659 &  x662 &  x671 &  x680 &  x686 &  x688 &  x689 &  x707 &  x722 &  x725 &  x728 &  x731 &  x734 &  x746 &  x764 &  x794 &  x812 &  x851 &  x866 &  x869 &  x878 &  x884 &  x953 &  x956 &  x962 &  x986 &  x1001 &  x1004 &  x1010 &  x1028 &  x1040 &  x1061 &  x1085 &  x1103 &  x1124 & ~x42 & ~x81 & ~x120 & ~x159 & ~x160 & ~x198 & ~x238 & ~x276 & ~x375 & ~x453 & ~x561 & ~x600 & ~x897 & ~x936;
assign c56 =  x8 &  x14 &  x29 &  x35 &  x44 &  x50 &  x56 &  x62 &  x68 &  x71 &  x79 &  x95 &  x98 &  x104 &  x107 &  x110 &  x118 &  x119 &  x122 &  x134 &  x137 &  x143 &  x157 &  x170 &  x179 &  x185 &  x191 &  x196 &  x197 &  x203 &  x212 &  x215 &  x218 &  x221 &  x224 &  x233 &  x235 &  x242 &  x245 &  x248 &  x260 &  x272 &  x274 &  x281 &  x284 &  x293 &  x296 &  x311 &  x317 &  x332 &  x341 &  x344 &  x352 &  x353 &  x355 &  x356 &  x359 &  x362 &  x368 &  x374 &  x377 &  x386 &  x394 &  x395 &  x401 &  x410 &  x422 &  x425 &  x437 &  x446 &  x449 &  x452 &  x479 &  x482 &  x491 &  x503 &  x515 &  x518 &  x530 &  x533 &  x539 &  x554 &  x581 &  x584 &  x587 &  x590 &  x596 &  x602 &  x605 &  x611 &  x614 &  x626 &  x638 &  x653 &  x674 &  x692 &  x695 &  x716 &  x722 &  x725 &  x728 &  x731 &  x740 &  x743 &  x746 &  x752 &  x755 &  x767 &  x773 &  x794 &  x803 &  x815 &  x818 &  x833 &  x842 &  x845 &  x863 &  x869 &  x878 &  x881 &  x893 &  x896 &  x905 &  x938 &  x950 &  x962 &  x971 &  x974 &  x977 &  x980 &  x992 &  x1001 &  x1010 &  x1013 &  x1022 &  x1034 &  x1064 &  x1067 &  x1070 &  x1076 &  x1085 &  x1094 &  x1097 &  x1100 &  x1106 &  x1130 & ~x3 & ~x4 & ~x108 & ~x129 & ~x148 & ~x168 & ~x186 & ~x207 & ~x252 & ~x405 & ~x444 & ~x741 & ~x780 & ~x936;
assign c58 =  x2 &  x14 &  x26 &  x29 &  x47 &  x50 &  x56 &  x71 &  x74 &  x80 &  x86 &  x104 &  x107 &  x119 &  x125 &  x149 &  x152 &  x161 &  x164 &  x167 &  x170 &  x173 &  x182 &  x185 &  x188 &  x191 &  x200 &  x203 &  x212 &  x215 &  x224 &  x227 &  x242 &  x245 &  x248 &  x263 &  x269 &  x281 &  x284 &  x302 &  x305 &  x308 &  x311 &  x332 &  x335 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x398 &  x413 &  x419 &  x425 &  x434 &  x440 &  x446 &  x455 &  x458 &  x464 &  x479 &  x482 &  x485 &  x488 &  x497 &  x500 &  x509 &  x512 &  x515 &  x518 &  x533 &  x536 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x566 &  x569 &  x578 &  x587 &  x602 &  x605 &  x608 &  x614 &  x617 &  x632 &  x638 &  x644 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x671 &  x680 &  x683 &  x689 &  x692 &  x695 &  x701 &  x703 &  x707 &  x713 &  x716 &  x728 &  x731 &  x734 &  x746 &  x749 &  x752 &  x761 &  x788 &  x791 &  x794 &  x809 &  x821 &  x833 &  x845 &  x848 &  x857 &  x861 &  x869 &  x878 &  x887 &  x890 &  x900 &  x901 &  x920 &  x926 &  x935 &  x940 &  x941 &  x944 &  x950 &  x959 &  x983 &  x992 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1031 &  x1034 &  x1037 &  x1055 &  x1073 &  x1082 &  x1085 &  x1094 &  x1097 &  x1100 &  x1115 &  x1121 & ~x273 & ~x511 & ~x558 & ~x636 & ~x714;
assign c510 =  x2 &  x5 &  x17 &  x20 &  x35 &  x38 &  x41 &  x47 &  x56 &  x65 &  x74 &  x77 &  x101 &  x104 &  x113 &  x128 &  x143 &  x146 &  x164 &  x179 &  x194 &  x200 &  x203 &  x209 &  x224 &  x233 &  x245 &  x251 &  x260 &  x269 &  x272 &  x287 &  x305 &  x308 &  x314 &  x319 &  x320 &  x323 &  x341 &  x368 &  x371 &  x374 &  x377 &  x410 &  x413 &  x431 &  x443 &  x452 &  x464 &  x475 &  x494 &  x506 &  x521 &  x523 &  x530 &  x533 &  x563 &  x581 &  x593 &  x605 &  x614 &  x620 &  x623 &  x641 &  x659 &  x671 &  x680 &  x692 &  x698 &  x701 &  x716 &  x719 &  x731 &  x746 &  x761 &  x782 &  x788 &  x806 &  x820 &  x836 &  x839 &  x857 &  x860 &  x872 &  x890 &  x898 &  x902 &  x905 &  x923 &  x929 &  x935 &  x937 &  x941 &  x953 &  x962 &  x965 &  x968 &  x974 &  x989 &  x998 &  x1004 &  x1034 &  x1037 &  x1040 &  x1043 &  x1058 &  x1061 &  x1064 &  x1079 &  x1088 &  x1091 &  x1103 &  x1106 &  x1109 &  x1115 &  x1130 & ~x237 & ~x597 & ~x903 & ~x948 & ~x951;
assign c512 =  x92 &  x227 &  x457 &  x579 &  x725 &  x884 & ~x504 & ~x909;
assign c514 =  x11 &  x26 &  x44 &  x47 &  x65 &  x83 &  x104 &  x107 &  x110 &  x143 &  x155 &  x167 &  x176 &  x179 &  x185 &  x188 &  x224 &  x230 &  x233 &  x242 &  x251 &  x260 &  x272 &  x284 &  x287 &  x293 &  x296 &  x299 &  x329 &  x338 &  x341 &  x356 &  x374 &  x413 &  x416 &  x428 &  x437 &  x461 &  x470 &  x476 &  x491 &  x530 &  x533 &  x548 &  x551 &  x560 &  x590 &  x599 &  x605 &  x617 &  x629 &  x632 &  x638 &  x644 &  x662 &  x665 &  x674 &  x683 &  x695 &  x707 &  x719 &  x731 &  x782 &  x794 &  x800 &  x806 &  x809 &  x812 &  x818 &  x836 &  x839 &  x845 &  x848 &  x851 &  x857 &  x872 &  x881 &  x899 &  x908 &  x911 &  x917 &  x920 &  x923 &  x941 &  x962 &  x968 &  x977 &  x992 &  x1022 &  x1043 &  x1046 &  x1049 &  x1061 &  x1064 &  x1070 &  x1091 &  x1094 &  x1103 &  x1115 &  x1127 & ~x9 & ~x48 & ~x87 & ~x282 & ~x361 & ~x400 & ~x595 & ~x672 & ~x750 & ~x864 & ~x942 & ~x1068;
assign c516 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x95 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x125 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x239 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x341 &  x344 &  x347 &  x350 &  x353 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x380 &  x383 &  x386 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x560 &  x563 &  x566 &  x569 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x704 &  x710 &  x716 &  x719 &  x722 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x974 &  x977 &  x980 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 & ~x159 & ~x160 & ~x198 & ~x207 & ~x237 & ~x246 & ~x363 & ~x444 & ~x522 & ~x561 & ~x600 & ~x678 & ~x717 & ~x846 & ~x885 & ~x984 & ~x1029 & ~x1086;
assign c518 =  x5 &  x8 &  x11 &  x20 &  x23 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x62 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x98 &  x101 &  x107 &  x113 &  x116 &  x122 &  x125 &  x128 &  x131 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x170 &  x173 &  x176 &  x179 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x290 &  x293 &  x299 &  x305 &  x308 &  x314 &  x317 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x380 &  x383 &  x392 &  x395 &  x398 &  x401 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x446 &  x449 &  x452 &  x455 &  x467 &  x470 &  x473 &  x476 &  x479 &  x485 &  x488 &  x494 &  x500 &  x503 &  x509 &  x515 &  x518 &  x524 &  x527 &  x530 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x563 &  x566 &  x572 &  x581 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x629 &  x632 &  x635 &  x638 &  x644 &  x647 &  x650 &  x653 &  x659 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x704 &  x707 &  x710 &  x713 &  x719 &  x722 &  x725 &  x728 &  x734 &  x743 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x779 &  x782 &  x785 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x893 &  x896 &  x899 &  x902 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x932 &  x935 &  x938 &  x944 &  x947 &  x950 &  x953 &  x956 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1118 &  x1127 &  x1130 & ~x159 & ~x160 & ~x199 & ~x207 & ~x237 & ~x246 & ~x276 & ~x363 & ~x364 & ~x402 & ~x441 & ~x480 & ~x717 & ~x756 & ~x951;
assign c520 =  x53 &  x191 &  x226 &  x440 &  x457 &  x461 &  x803 &  x905 &  x947 &  x998 & ~x223 & ~x798 & ~x837;
assign c522 =  x14 &  x17 &  x23 &  x35 &  x44 &  x53 &  x68 &  x80 &  x83 &  x89 &  x101 &  x104 &  x107 &  x113 &  x122 &  x128 &  x134 &  x137 &  x146 &  x152 &  x158 &  x167 &  x170 &  x182 &  x185 &  x197 &  x209 &  x221 &  x227 &  x242 &  x245 &  x254 &  x260 &  x281 &  x284 &  x293 &  x302 &  x314 &  x323 &  x338 &  x344 &  x347 &  x368 &  x383 &  x392 &  x395 &  x407 &  x425 &  x431 &  x440 &  x452 &  x455 &  x461 &  x467 &  x470 &  x473 &  x479 &  x488 &  x491 &  x500 &  x503 &  x506 &  x509 &  x512 &  x518 &  x521 &  x533 &  x551 &  x557 &  x560 &  x563 &  x581 &  x584 &  x605 &  x611 &  x629 &  x632 &  x635 &  x644 &  x647 &  x662 &  x665 &  x668 &  x674 &  x677 &  x683 &  x695 &  x698 &  x704 &  x710 &  x713 &  x719 &  x722 &  x728 &  x737 &  x743 &  x746 &  x749 &  x758 &  x776 &  x809 &  x815 &  x833 &  x839 &  x845 &  x851 &  x866 &  x869 &  x887 &  x893 &  x899 &  x902 &  x935 &  x941 &  x944 &  x962 &  x977 &  x992 &  x1007 &  x1025 &  x1046 &  x1049 &  x1052 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1088 &  x1127 &  x1130 & ~x550 & ~x589 & ~x621 & ~x675 & ~x699 & ~x738 & ~x834 & ~x912 & ~x952 & ~x1068;
assign c524 =  x20 &  x26 &  x40 &  x41 &  x44 &  x79 &  x86 &  x152 &  x158 &  x182 &  x188 &  x191 &  x203 &  x217 &  x242 &  x287 &  x302 &  x320 &  x326 &  x335 &  x350 &  x356 &  x368 &  x379 &  x386 &  x392 &  x398 &  x404 &  x410 &  x418 &  x457 &  x461 &  x470 &  x509 &  x515 &  x530 &  x554 &  x563 &  x578 &  x587 &  x611 &  x632 &  x635 &  x653 &  x677 &  x700 &  x713 &  x770 &  x773 &  x808 &  x818 &  x848 &  x893 &  x911 &  x932 &  x935 &  x944 &  x956 &  x965 &  x973 &  x977 &  x1001 &  x1004 &  x1013 &  x1028 &  x1040 &  x1055 &  x1064 &  x1070 &  x1073 &  x1075 &  x1076 &  x1106 &  x1109 & ~x516 & ~x828;
assign c526 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x77 &  x86 &  x92 &  x95 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x196 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x235 &  x242 &  x245 &  x248 &  x251 &  x254 &  x260 &  x263 &  x269 &  x272 &  x274 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x391 &  x395 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x430 &  x431 &  x434 &  x437 &  x440 &  x443 &  x449 &  x452 &  x458 &  x464 &  x467 &  x469 &  x470 &  x473 &  x476 &  x479 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x511 &  x512 &  x518 &  x521 &  x524 &  x527 &  x533 &  x536 &  x545 &  x548 &  x557 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x695 &  x698 &  x701 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x767 &  x770 &  x773 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x869 &  x875 &  x877 &  x878 &  x881 &  x884 &  x893 &  x896 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x971 &  x974 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1070 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x159 & ~x198 & ~x199 & ~x237 & ~x402 & ~x519 & ~x561 & ~x600 & ~x639 & ~x789;
assign c528 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x29 &  x32 &  x35 &  x38 &  x44 &  x50 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x79 &  x80 &  x83 &  x86 &  x92 &  x95 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x118 &  x119 &  x122 &  x131 &  x137 &  x143 &  x146 &  x152 &  x155 &  x157 &  x164 &  x167 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x194 &  x197 &  x200 &  x203 &  x206 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x235 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x260 &  x263 &  x269 &  x272 &  x276 &  x277 &  x278 &  x281 &  x287 &  x296 &  x299 &  x302 &  x308 &  x311 &  x313 &  x314 &  x316 &  x323 &  x326 &  x332 &  x335 &  x341 &  x347 &  x350 &  x353 &  x355 &  x356 &  x359 &  x362 &  x368 &  x374 &  x377 &  x383 &  x386 &  x389 &  x394 &  x395 &  x401 &  x404 &  x413 &  x416 &  x431 &  x434 &  x437 &  x443 &  x446 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x473 &  x476 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x506 &  x509 &  x515 &  x518 &  x521 &  x524 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x551 &  x554 &  x557 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x629 &  x635 &  x641 &  x647 &  x650 &  x653 &  x656 &  x671 &  x674 &  x677 &  x680 &  x686 &  x689 &  x695 &  x698 &  x701 &  x707 &  x710 &  x716 &  x719 &  x725 &  x728 &  x731 &  x734 &  x737 &  x743 &  x746 &  x752 &  x758 &  x770 &  x773 &  x776 &  x788 &  x791 &  x793 &  x794 &  x803 &  x806 &  x809 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x832 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x866 &  x869 &  x871 &  x875 &  x878 &  x881 &  x884 &  x890 &  x893 &  x896 &  x905 &  x910 &  x911 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x956 &  x959 &  x968 &  x971 &  x977 &  x980 &  x983 &  x986 &  x988 &  x989 &  x992 &  x998 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x24 & ~x63 & ~x102 & ~x174 & ~x213 & ~x288 & ~x327 & ~x444 & ~x546 & ~x585 & ~x663 & ~x897 & ~x936;
assign c530 =  x2 &  x5 &  x11 &  x17 &  x20 &  x23 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x59 &  x62 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x122 &  x125 &  x128 &  x137 &  x140 &  x143 &  x146 &  x152 &  x158 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x469 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x524 &  x533 &  x536 &  x539 &  x542 &  x545 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x584 &  x587 &  x590 &  x593 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x653 &  x656 &  x662 &  x668 &  x671 &  x674 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x773 &  x776 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x818 &  x821 &  x827 &  x833 &  x836 &  x839 &  x842 &  x848 &  x857 &  x860 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x905 &  x908 &  x911 &  x917 &  x920 &  x926 &  x929 &  x932 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x81 & ~x82 & ~x90 & ~x120 & ~x246 & ~x363 & ~x402 & ~x462 & ~x501 & ~x540 & ~x780 & ~x1014 & ~x1047 & ~x1053 & ~x1086 & ~x1092;
assign c532 =  x2 &  x5 &  x14 &  x29 &  x38 &  x44 &  x46 &  x71 &  x79 &  x85 &  x86 &  x98 &  x110 &  x116 &  x118 &  x119 &  x124 &  x125 &  x146 &  x152 &  x161 &  x164 &  x185 &  x188 &  x200 &  x203 &  x221 &  x224 &  x242 &  x254 &  x260 &  x281 &  x293 &  x302 &  x308 &  x313 &  x314 &  x323 &  x326 &  x329 &  x332 &  x347 &  x352 &  x359 &  x365 &  x368 &  x374 &  x380 &  x386 &  x391 &  x398 &  x404 &  x425 &  x440 &  x461 &  x467 &  x472 &  x476 &  x485 &  x497 &  x511 &  x530 &  x542 &  x545 &  x557 &  x560 &  x569 &  x581 &  x590 &  x605 &  x608 &  x617 &  x623 &  x632 &  x635 &  x641 &  x644 &  x659 &  x668 &  x683 &  x686 &  x689 &  x701 &  x716 &  x728 &  x737 &  x755 &  x761 &  x770 &  x794 &  x809 &  x812 &  x830 &  x836 &  x842 &  x863 &  x866 &  x869 &  x871 &  x872 &  x877 &  x881 &  x896 &  x899 &  x908 &  x910 &  x917 &  x920 &  x935 &  x938 &  x949 &  x953 &  x959 &  x965 &  x968 &  x983 &  x989 &  x992 &  x995 &  x1004 &  x1022 &  x1025 &  x1037 &  x1055 &  x1064 &  x1066 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1105 &  x1115 &  x1121 & ~x741 & ~x1068;
assign c534 =  x2 &  x8 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x56 &  x59 &  x62 &  x65 &  x71 &  x74 &  x80 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x119 &  x122 &  x125 &  x128 &  x131 &  x140 &  x152 &  x155 &  x158 &  x161 &  x167 &  x170 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x206 &  x209 &  x212 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x245 &  x251 &  x254 &  x257 &  x260 &  x263 &  x269 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x317 &  x323 &  x326 &  x329 &  x338 &  x347 &  x350 &  x353 &  x359 &  x362 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x443 &  x449 &  x464 &  x467 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x506 &  x509 &  x512 &  x518 &  x521 &  x524 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x589 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x614 &  x623 &  x626 &  x628 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x646 &  x647 &  x650 &  x653 &  x656 &  x659 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x725 &  x727 &  x734 &  x737 &  x740 &  x746 &  x761 &  x766 &  x767 &  x773 &  x782 &  x784 &  x785 &  x791 &  x797 &  x803 &  x805 &  x809 &  x812 &  x815 &  x824 &  x830 &  x833 &  x842 &  x844 &  x854 &  x863 &  x869 &  x872 &  x875 &  x878 &  x880 &  x884 &  x889 &  x896 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x935 &  x944 &  x959 &  x965 &  x968 &  x974 &  x980 &  x989 &  x1001 &  x1010 &  x1013 &  x1016 &  x1022 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1057 &  x1058 &  x1061 &  x1067 &  x1070 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1096 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 & ~x42;
assign c536 =  x2 &  x5 &  x8 &  x11 &  x17 &  x20 &  x26 &  x29 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x230 &  x233 &  x236 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x392 &  x395 &  x397 &  x398 &  x401 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x436 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x464 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x617 &  x620 &  x623 &  x626 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x800 &  x803 &  x806 &  x809 &  x812 &  x818 &  x821 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x977 &  x980 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x120 & ~x159 & ~x198 & ~x231 & ~x237 & ~x270 & ~x309 & ~x330 & ~x348 & ~x369 & ~x639 & ~x828 & ~x906 & ~x984;
assign c538 =  x8 &  x11 &  x14 &  x29 &  x32 &  x35 &  x44 &  x50 &  x62 &  x98 &  x104 &  x110 &  x116 &  x125 &  x131 &  x152 &  x158 &  x167 &  x170 &  x179 &  x182 &  x191 &  x206 &  x215 &  x218 &  x227 &  x239 &  x245 &  x251 &  x260 &  x263 &  x266 &  x275 &  x278 &  x284 &  x287 &  x296 &  x299 &  x308 &  x326 &  x347 &  x353 &  x359 &  x374 &  x395 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x428 &  x431 &  x434 &  x436 &  x437 &  x440 &  x449 &  x464 &  x470 &  x476 &  x479 &  x482 &  x488 &  x497 &  x512 &  x524 &  x527 &  x536 &  x539 &  x542 &  x545 &  x547 &  x548 &  x554 &  x572 &  x575 &  x590 &  x593 &  x602 &  x617 &  x623 &  x635 &  x638 &  x659 &  x665 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x701 &  x704 &  x710 &  x722 &  x725 &  x731 &  x740 &  x745 &  x749 &  x755 &  x761 &  x764 &  x770 &  x773 &  x784 &  x788 &  x791 &  x794 &  x797 &  x803 &  x806 &  x818 &  x824 &  x836 &  x844 &  x851 &  x854 &  x860 &  x863 &  x872 &  x875 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x926 &  x929 &  x947 &  x950 &  x968 &  x980 &  x983 &  x995 &  x1001 &  x1010 &  x1013 &  x1019 &  x1022 &  x1034 &  x1040 &  x1049 &  x1070 &  x1091 &  x1094 &  x1100 &  x1106 &  x1121 & ~x393 & ~x759 & ~x795 & ~x798 & ~x835 & ~x873;
assign c540 =  x14 &  x23 &  x110 &  x122 &  x125 &  x158 &  x172 &  x173 &  x290 &  x296 &  x329 &  x368 &  x373 &  x383 &  x406 &  x434 &  x449 &  x479 &  x529 &  x542 &  x553 &  x557 &  x632 &  x680 &  x685 &  x725 &  x731 &  x742 &  x780 &  x781 &  x803 &  x806 &  x819 &  x863 &  x878 &  x893 &  x896 &  x920 &  x1007 &  x1022 &  x1052 &  x1057 &  x1096 &  x1112 & ~x636 & ~x753 & ~x909 & ~x987;
assign c542 =  x8 &  x11 &  x20 &  x29 &  x53 &  x56 &  x62 &  x71 &  x83 &  x89 &  x95 &  x100 &  x104 &  x110 &  x112 &  x113 &  x119 &  x122 &  x137 &  x143 &  x149 &  x173 &  x176 &  x178 &  x188 &  x194 &  x242 &  x248 &  x254 &  x266 &  x269 &  x281 &  x284 &  x290 &  x305 &  x314 &  x317 &  x334 &  x341 &  x353 &  x356 &  x359 &  x362 &  x371 &  x373 &  x374 &  x377 &  x380 &  x392 &  x413 &  x416 &  x419 &  x424 &  x449 &  x461 &  x464 &  x467 &  x470 &  x485 &  x502 &  x506 &  x509 &  x512 &  x521 &  x527 &  x545 &  x557 &  x563 &  x578 &  x587 &  x593 &  x596 &  x611 &  x617 &  x626 &  x644 &  x653 &  x662 &  x668 &  x677 &  x683 &  x686 &  x695 &  x698 &  x710 &  x716 &  x731 &  x734 &  x737 &  x740 &  x749 &  x752 &  x764 &  x767 &  x773 &  x782 &  x785 &  x791 &  x806 &  x815 &  x818 &  x823 &  x833 &  x836 &  x848 &  x854 &  x857 &  x863 &  x875 &  x878 &  x884 &  x895 &  x896 &  x902 &  x920 &  x923 &  x926 &  x928 &  x929 &  x934 &  x941 &  x944 &  x965 &  x968 &  x989 &  x995 &  x998 &  x1001 &  x1031 &  x1034 &  x1043 &  x1055 &  x1061 &  x1072 &  x1073 &  x1076 &  x1079 &  x1084 &  x1088 &  x1097 &  x1100 &  x1111 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130;
assign c544 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x35 &  x38 &  x41 &  x44 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x146 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x280 &  x281 &  x284 &  x287 &  x290 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x319 &  x320 &  x323 &  x326 &  x329 &  x332 &  x341 &  x344 &  x347 &  x350 &  x353 &  x362 &  x365 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x395 &  x397 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x458 &  x461 &  x464 &  x467 &  x473 &  x476 &  x479 &  x482 &  x488 &  x491 &  x494 &  x497 &  x500 &  x506 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x611 &  x614 &  x617 &  x620 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x674 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x719 &  x722 &  x728 &  x731 &  x734 &  x737 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x803 &  x806 &  x809 &  x812 &  x818 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x889 &  x890 &  x893 &  x896 &  x905 &  x908 &  x911 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x950 &  x953 &  x956 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1070 &  x1072 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1099 &  x1100 &  x1103 &  x1109 &  x1111 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x42 & ~x291 & ~x858;
assign c546 =  x29 &  x38 &  x80 &  x86 &  x89 &  x107 &  x116 &  x125 &  x134 &  x179 &  x236 &  x239 &  x242 &  x254 &  x284 &  x308 &  x335 &  x338 &  x346 &  x371 &  x386 &  x392 &  x398 &  x419 &  x436 &  x437 &  x467 &  x475 &  x508 &  x524 &  x547 &  x575 &  x581 &  x605 &  x608 &  x635 &  x647 &  x683 &  x706 &  x731 &  x737 &  x749 &  x755 &  x764 &  x788 &  x803 &  x806 &  x809 &  x823 &  x857 &  x881 &  x884 &  x893 &  x896 &  x905 &  x908 &  x920 &  x932 &  x935 &  x938 &  x950 &  x959 &  x965 &  x974 &  x992 &  x1007 &  x1013 &  x1016 &  x1022 &  x1028 &  x1058 &  x1064 &  x1076 &  x1085 &  x1091 &  x1100 &  x1106 &  x1112 &  x1118 & ~x394 & ~x432 & ~x870;
assign c548 =  x2 &  x5 &  x11 &  x23 &  x29 &  x32 &  x38 &  x44 &  x47 &  x65 &  x71 &  x74 &  x79 &  x80 &  x86 &  x101 &  x104 &  x110 &  x116 &  x118 &  x122 &  x128 &  x131 &  x137 &  x140 &  x149 &  x155 &  x158 &  x161 &  x164 &  x167 &  x185 &  x196 &  x200 &  x203 &  x209 &  x218 &  x221 &  x224 &  x230 &  x233 &  x235 &  x239 &  x242 &  x248 &  x251 &  x260 &  x263 &  x266 &  x272 &  x275 &  x278 &  x290 &  x296 &  x305 &  x308 &  x314 &  x317 &  x329 &  x332 &  x335 &  x347 &  x353 &  x356 &  x362 &  x365 &  x371 &  x377 &  x383 &  x386 &  x389 &  x392 &  x394 &  x398 &  x401 &  x404 &  x407 &  x413 &  x419 &  x422 &  x425 &  x428 &  x437 &  x440 &  x446 &  x452 &  x455 &  x458 &  x470 &  x473 &  x476 &  x485 &  x488 &  x494 &  x497 &  x500 &  x506 &  x509 &  x512 &  x515 &  x521 &  x524 &  x527 &  x530 &  x539 &  x542 &  x545 &  x548 &  x551 &  x560 &  x575 &  x578 &  x584 &  x593 &  x602 &  x608 &  x617 &  x620 &  x626 &  x629 &  x635 &  x653 &  x659 &  x662 &  x677 &  x683 &  x689 &  x692 &  x695 &  x701 &  x704 &  x707 &  x710 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x749 &  x758 &  x761 &  x770 &  x788 &  x794 &  x803 &  x809 &  x812 &  x815 &  x818 &  x830 &  x833 &  x839 &  x845 &  x851 &  x857 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x884 &  x893 &  x905 &  x911 &  x914 &  x920 &  x923 &  x926 &  x935 &  x938 &  x947 &  x956 &  x959 &  x962 &  x965 &  x971 &  x977 &  x986 &  x992 &  x998 &  x1001 &  x1010 &  x1016 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1043 &  x1046 &  x1055 &  x1058 &  x1064 &  x1070 &  x1073 &  x1076 &  x1088 &  x1100 &  x1103 &  x1112 &  x1118 &  x1124 &  x1127 & ~x12 & ~x52 & ~x114 & ~x153 & ~x154 & ~x192 & ~x207 & ~x231 & ~x246 & ~x288 & ~x327 & ~x328 & ~x366 & ~x405 & ~x444 & ~x624 & ~x663;
assign c550 =  x8 &  x26 &  x59 &  x86 &  x89 &  x95 &  x134 &  x140 &  x155 &  x164 &  x167 &  x173 &  x179 &  x182 &  x191 &  x212 &  x236 &  x320 &  x335 &  x344 &  x383 &  x404 &  x416 &  x434 &  x440 &  x473 &  x494 &  x506 &  x521 &  x545 &  x563 &  x569 &  x584 &  x593 &  x605 &  x626 &  x635 &  x650 &  x665 &  x683 &  x692 &  x734 &  x742 &  x761 &  x770 &  x781 &  x803 &  x830 &  x842 &  x866 &  x878 &  x887 &  x890 &  x893 &  x896 &  x905 &  x911 &  x914 &  x917 &  x926 &  x950 &  x953 &  x1004 &  x1007 &  x1028 &  x1043 &  x1049 &  x1096 &  x1109 &  x1112 &  x1130 & ~x468 & ~x667 & ~x675;
assign c552 =  x20 &  x26 &  x32 &  x35 &  x38 &  x44 &  x47 &  x56 &  x59 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x101 &  x104 &  x110 &  x116 &  x119 &  x122 &  x125 &  x131 &  x134 &  x137 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x191 &  x194 &  x197 &  x200 &  x209 &  x212 &  x215 &  x227 &  x230 &  x233 &  x239 &  x242 &  x248 &  x251 &  x257 &  x260 &  x269 &  x272 &  x278 &  x287 &  x293 &  x296 &  x308 &  x317 &  x320 &  x326 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x352 &  x353 &  x356 &  x359 &  x365 &  x371 &  x374 &  x380 &  x383 &  x386 &  x389 &  x395 &  x398 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x428 &  x443 &  x446 &  x449 &  x458 &  x461 &  x470 &  x479 &  x482 &  x488 &  x491 &  x494 &  x497 &  x500 &  x509 &  x512 &  x515 &  x518 &  x521 &  x527 &  x533 &  x536 &  x539 &  x542 &  x548 &  x554 &  x566 &  x569 &  x575 &  x581 &  x584 &  x593 &  x602 &  x608 &  x610 &  x611 &  x614 &  x623 &  x626 &  x629 &  x638 &  x641 &  x647 &  x649 &  x656 &  x671 &  x674 &  x688 &  x689 &  x691 &  x692 &  x695 &  x707 &  x719 &  x725 &  x728 &  x731 &  x734 &  x740 &  x749 &  x752 &  x755 &  x758 &  x767 &  x770 &  x779 &  x782 &  x791 &  x794 &  x797 &  x800 &  x806 &  x815 &  x821 &  x827 &  x830 &  x833 &  x836 &  x842 &  x848 &  x851 &  x857 &  x866 &  x875 &  x884 &  x890 &  x902 &  x905 &  x908 &  x914 &  x920 &  x923 &  x926 &  x929 &  x935 &  x938 &  x950 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x977 &  x995 &  x1001 &  x1007 &  x1010 &  x1016 &  x1025 &  x1055 &  x1058 &  x1061 &  x1064 &  x1088 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1115 &  x1124 &  x1127 & ~x3 & ~x12 & ~x51 & ~x82 & ~x90 & ~x291 & ~x292 & ~x330 & ~x370 & ~x408;
assign c554 =  x38 &  x101 &  x191 &  x200 &  x290 &  x335 &  x344 &  x434 &  x436 &  x440 &  x491 &  x551 &  x620 &  x653 &  x680 &  x713 &  x731 &  x781 &  x803 &  x820 &  x917 &  x938 &  x1095 &  x1096 &  x1121 &  x1127 &  x1130 & ~x510 & ~x627 & ~x705 & ~x706;
assign c556 =  x1 &  x2 &  x5 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x40 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x65 &  x68 &  x71 &  x74 &  x77 &  x79 &  x80 &  x83 &  x89 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x157 &  x158 &  x161 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x323 &  x326 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x353 &  x356 &  x362 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x544 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x716 &  x719 &  x722 &  x725 &  x728 &  x734 &  x737 &  x740 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x12 & ~x13 & ~x51 & ~x52 & ~x90 & ~x129 & ~x168 & ~x186 & ~x246 & ~x285 & ~x328 & ~x366 & ~x405 & ~x444 & ~x546 & ~x585 & ~x633;
assign c558 =  x5 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x107 &  x113 &  x119 &  x128 &  x131 &  x146 &  x170 &  x176 &  x182 &  x197 &  x211 &  x212 &  x224 &  x227 &  x230 &  x235 &  x236 &  x251 &  x254 &  x257 &  x260 &  x266 &  x269 &  x274 &  x275 &  x281 &  x284 &  x290 &  x293 &  x311 &  x317 &  x329 &  x350 &  x352 &  x359 &  x362 &  x365 &  x374 &  x377 &  x389 &  x391 &  x395 &  x404 &  x410 &  x419 &  x422 &  x430 &  x431 &  x443 &  x446 &  x449 &  x452 &  x464 &  x467 &  x485 &  x497 &  x500 &  x503 &  x506 &  x509 &  x511 &  x512 &  x515 &  x521 &  x536 &  x539 &  x545 &  x548 &  x550 &  x566 &  x569 &  x599 &  x602 &  x608 &  x620 &  x623 &  x629 &  x632 &  x635 &  x641 &  x644 &  x650 &  x662 &  x665 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x701 &  x704 &  x707 &  x719 &  x728 &  x734 &  x737 &  x740 &  x743 &  x758 &  x764 &  x770 &  x776 &  x779 &  x782 &  x788 &  x791 &  x794 &  x797 &  x806 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x839 &  x845 &  x860 &  x875 &  x881 &  x887 &  x890 &  x896 &  x911 &  x920 &  x929 &  x935 &  x944 &  x947 &  x953 &  x959 &  x968 &  x971 &  x974 &  x986 &  x989 &  x998 &  x1001 &  x1007 &  x1013 &  x1016 &  x1019 &  x1025 &  x1034 &  x1043 &  x1055 &  x1067 &  x1073 &  x1079 &  x1085 &  x1100 &  x1112 &  x1124 &  x1127 &  x1130 & ~x199 & ~x237 & ~x324 & ~x336 & ~x441 & ~x600;
assign c560 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x79 &  x83 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x152 &  x155 &  x157 &  x158 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x188 &  x191 &  x194 &  x195 &  x196 &  x203 &  x206 &  x212 &  x215 &  x218 &  x221 &  x230 &  x233 &  x235 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x266 &  x269 &  x274 &  x281 &  x284 &  x287 &  x290 &  x302 &  x305 &  x308 &  x311 &  x323 &  x326 &  x332 &  x335 &  x338 &  x344 &  x347 &  x352 &  x353 &  x355 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x394 &  x395 &  x404 &  x413 &  x416 &  x419 &  x422 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x458 &  x461 &  x464 &  x470 &  x472 &  x473 &  x476 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x524 &  x530 &  x533 &  x539 &  x542 &  x548 &  x554 &  x557 &  x560 &  x563 &  x569 &  x572 &  x578 &  x581 &  x583 &  x584 &  x587 &  x590 &  x596 &  x602 &  x605 &  x608 &  x614 &  x620 &  x622 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x665 &  x671 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x701 &  x710 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x761 &  x767 &  x776 &  x779 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x821 &  x824 &  x830 &  x833 &  x836 &  x838 &  x839 &  x842 &  x845 &  x848 &  x851 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x877 &  x881 &  x884 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x914 &  x916 &  x920 &  x926 &  x935 &  x938 &  x941 &  x947 &  x950 &  x953 &  x956 &  x959 &  x968 &  x971 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1073 &  x1076 &  x1085 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1130 & ~x42 & ~x81 & ~x82;
assign c562 =  x8 &  x17 &  x20 &  x29 &  x32 &  x41 &  x47 &  x50 &  x56 &  x59 &  x62 &  x68 &  x74 &  x77 &  x86 &  x89 &  x95 &  x98 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x158 &  x161 &  x164 &  x167 &  x173 &  x176 &  x188 &  x191 &  x197 &  x200 &  x206 &  x209 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x290 &  x293 &  x299 &  x305 &  x308 &  x314 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x353 &  x359 &  x362 &  x365 &  x377 &  x383 &  x386 &  x389 &  x397 &  x401 &  x404 &  x413 &  x416 &  x422 &  x425 &  x428 &  x436 &  x437 &  x443 &  x446 &  x452 &  x458 &  x464 &  x485 &  x491 &  x497 &  x500 &  x503 &  x509 &  x518 &  x521 &  x527 &  x533 &  x539 &  x542 &  x545 &  x548 &  x563 &  x569 &  x572 &  x578 &  x581 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x608 &  x611 &  x617 &  x620 &  x626 &  x629 &  x632 &  x638 &  x647 &  x656 &  x662 &  x668 &  x671 &  x683 &  x686 &  x695 &  x704 &  x710 &  x713 &  x716 &  x719 &  x722 &  x731 &  x740 &  x743 &  x752 &  x755 &  x764 &  x767 &  x776 &  x779 &  x782 &  x785 &  x791 &  x794 &  x797 &  x803 &  x809 &  x815 &  x827 &  x836 &  x839 &  x842 &  x845 &  x857 &  x860 &  x863 &  x884 &  x887 &  x890 &  x896 &  x899 &  x905 &  x911 &  x914 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x959 &  x965 &  x968 &  x971 &  x974 &  x983 &  x986 &  x989 &  x998 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1049 &  x1052 &  x1058 &  x1061 &  x1073 &  x1076 &  x1079 &  x1088 &  x1091 &  x1094 &  x1097 &  x1112 &  x1115 &  x1121 &  x1124 & ~x159 & ~x198 & ~x237 & ~x315 & ~x354 & ~x441 & ~x519 & ~x558 & ~x559 & ~x597 & ~x636 & ~x675 & ~x714 & ~x735 & ~x753 & ~x831;
assign c564 =  x11 &  x35 &  x38 &  x41 &  x47 &  x95 &  x110 &  x113 &  x137 &  x140 &  x149 &  x167 &  x170 &  x185 &  x194 &  x209 &  x212 &  x230 &  x233 &  x245 &  x254 &  x263 &  x272 &  x281 &  x290 &  x299 &  x314 &  x323 &  x337 &  x341 &  x344 &  x365 &  x374 &  x383 &  x386 &  x389 &  x395 &  x413 &  x419 &  x425 &  x437 &  x446 &  x449 &  x458 &  x482 &  x491 &  x494 &  x509 &  x514 &  x521 &  x527 &  x533 &  x548 &  x569 &  x599 &  x601 &  x608 &  x613 &  x626 &  x632 &  x635 &  x652 &  x677 &  x709 &  x710 &  x713 &  x734 &  x740 &  x749 &  x752 &  x764 &  x767 &  x776 &  x797 &  x800 &  x809 &  x818 &  x827 &  x836 &  x857 &  x866 &  x878 &  x893 &  x898 &  x920 &  x923 &  x926 &  x932 &  x968 &  x976 &  x989 &  x992 &  x998 &  x1015 &  x1016 &  x1022 &  x1025 &  x1031 &  x1037 &  x1046 &  x1073 &  x1076 &  x1079 &  x1085 &  x1097 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1130 & ~x627 & ~x628 & ~x870 & ~x915 & ~x1065;
assign c566 =  x2 &  x5 &  x14 &  x35 &  x53 &  x56 &  x80 &  x83 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x137 &  x143 &  x146 &  x152 &  x173 &  x176 &  x179 &  x188 &  x191 &  x194 &  x197 &  x200 &  x206 &  x212 &  x221 &  x230 &  x233 &  x263 &  x269 &  x272 &  x278 &  x296 &  x314 &  x323 &  x326 &  x332 &  x338 &  x347 &  x353 &  x362 &  x365 &  x374 &  x392 &  x404 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x449 &  x455 &  x464 &  x467 &  x473 &  x476 &  x494 &  x500 &  x512 &  x527 &  x536 &  x542 &  x548 &  x551 &  x563 &  x566 &  x569 &  x581 &  x590 &  x608 &  x635 &  x638 &  x644 &  x647 &  x650 &  x659 &  x665 &  x667 &  x677 &  x689 &  x698 &  x706 &  x719 &  x722 &  x737 &  x740 &  x745 &  x749 &  x761 &  x767 &  x770 &  x779 &  x785 &  x800 &  x821 &  x833 &  x848 &  x860 &  x875 &  x890 &  x902 &  x905 &  x926 &  x929 &  x935 &  x941 &  x950 &  x962 &  x974 &  x980 &  x986 &  x998 &  x1001 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1037 &  x1040 &  x1058 &  x1061 &  x1070 &  x1079 &  x1082 &  x1088 &  x1091 &  x1103 &  x1109 &  x1112 &  x1121 &  x1124 &  x1130 & ~x324 & ~x348 & ~x558 & ~x564 & ~x600 & ~x678 & ~x717 & ~x819 & ~x1014 & ~x1125;
assign c568 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x29 &  x32 &  x35 &  x38 &  x40 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x79 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x112 &  x113 &  x116 &  x118 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x151 &  x152 &  x155 &  x157 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x178 &  x179 &  x182 &  x185 &  x188 &  x190 &  x191 &  x194 &  x196 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x229 &  x230 &  x233 &  x235 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x274 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x493 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x583 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x622 &  x623 &  x626 &  x629 &  x632 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x694 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x733 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x928 &  x929 &  x932 &  x934 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x967 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x997 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x36;
assign c570 =  x20 &  x35 &  x59 &  x101 &  x113 &  x170 &  x176 &  x179 &  x188 &  x203 &  x212 &  x236 &  x274 &  x287 &  x302 &  x317 &  x335 &  x341 &  x344 &  x353 &  x356 &  x358 &  x359 &  x374 &  x431 &  x469 &  x470 &  x503 &  x512 &  x548 &  x551 &  x588 &  x589 &  x596 &  x638 &  x659 &  x668 &  x671 &  x688 &  x722 &  x727 &  x734 &  x740 &  x755 &  x766 &  x770 &  x785 &  x812 &  x821 &  x848 &  x851 &  x866 &  x872 &  x875 &  x896 &  x926 &  x947 &  x977 &  x986 &  x989 &  x1004 &  x1016 &  x1067 &  x1088 &  x1100 &  x1124 &  x1127 &  x1130 & ~x558;
assign c572 =  x8 &  x20 &  x32 &  x35 &  x41 &  x65 &  x68 &  x110 &  x116 &  x122 &  x167 &  x173 &  x221 &  x248 &  x257 &  x272 &  x293 &  x305 &  x314 &  x350 &  x362 &  x416 &  x467 &  x506 &  x529 &  x551 &  x554 &  x557 &  x578 &  x593 &  x614 &  x623 &  x646 &  x647 &  x686 &  x724 &  x740 &  x746 &  x764 &  x767 &  x812 &  x819 &  x830 &  x833 &  x872 &  x890 &  x893 &  x897 &  x899 &  x986 &  x989 &  x998 &  x1037 &  x1079 &  x1085 &  x1100 &  x1112 &  x1127 & ~x589 & ~x714;
assign c574 =  x5 &  x8 &  x23 &  x41 &  x89 &  x98 &  x113 &  x155 &  x197 &  x206 &  x218 &  x224 &  x235 &  x242 &  x257 &  x260 &  x287 &  x299 &  x313 &  x317 &  x332 &  x350 &  x377 &  x395 &  x401 &  x410 &  x416 &  x430 &  x440 &  x458 &  x469 &  x506 &  x509 &  x515 &  x518 &  x539 &  x569 &  x572 &  x581 &  x599 &  x602 &  x608 &  x617 &  x629 &  x698 &  x704 &  x707 &  x716 &  x746 &  x767 &  x794 &  x833 &  x839 &  x848 &  x869 &  x899 &  x905 &  x908 &  x911 &  x926 &  x929 &  x944 &  x947 &  x962 &  x965 &  x986 &  x1001 &  x1019 &  x1025 &  x1028 &  x1031 &  x1046 &  x1085 &  x1091 &  x1109 &  x1121 & ~x277 & ~x441 & ~x519 & ~x558 & ~x561 & ~x600 & ~x828;
assign c576 =  x2 &  x5 &  x17 &  x32 &  x35 &  x44 &  x58 &  x59 &  x71 &  x74 &  x77 &  x83 &  x86 &  x89 &  x98 &  x109 &  x110 &  x122 &  x128 &  x134 &  x148 &  x149 &  x155 &  x161 &  x164 &  x167 &  x179 &  x182 &  x188 &  x191 &  x200 &  x208 &  x212 &  x218 &  x236 &  x239 &  x245 &  x251 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x281 &  x287 &  x299 &  x302 &  x305 &  x308 &  x311 &  x317 &  x320 &  x326 &  x332 &  x335 &  x338 &  x347 &  x353 &  x368 &  x374 &  x383 &  x386 &  x392 &  x398 &  x404 &  x410 &  x413 &  x422 &  x425 &  x428 &  x431 &  x452 &  x457 &  x458 &  x461 &  x467 &  x473 &  x476 &  x479 &  x482 &  x497 &  x503 &  x506 &  x509 &  x518 &  x523 &  x524 &  x527 &  x530 &  x536 &  x545 &  x554 &  x560 &  x563 &  x566 &  x568 &  x581 &  x587 &  x599 &  x602 &  x611 &  x614 &  x635 &  x644 &  x646 &  x653 &  x656 &  x662 &  x665 &  x671 &  x674 &  x680 &  x683 &  x685 &  x686 &  x689 &  x695 &  x698 &  x713 &  x716 &  x719 &  x725 &  x737 &  x755 &  x763 &  x764 &  x779 &  x782 &  x794 &  x800 &  x803 &  x818 &  x820 &  x830 &  x833 &  x839 &  x854 &  x860 &  x866 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x911 &  x917 &  x929 &  x941 &  x947 &  x962 &  x965 &  x968 &  x977 &  x986 &  x995 &  x998 &  x1001 &  x1007 &  x1013 &  x1016 &  x1019 &  x1025 &  x1034 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1064 &  x1070 &  x1079 &  x1085 &  x1094 &  x1097 &  x1109 &  x1112 &  x1115 &  x1118 & ~x360;
assign c578 =  x26 &  x221 &  x290 &  x338 &  x464 &  x515 &  x529 &  x579 &  x584 &  x641 &  x644 &  x665 &  x713 &  x724 &  x1043 &  x1097 & ~x1027;
assign c580 =  x5 &  x17 &  x23 &  x35 &  x41 &  x46 &  x50 &  x53 &  x56 &  x59 &  x74 &  x77 &  x89 &  x92 &  x95 &  x107 &  x112 &  x116 &  x122 &  x143 &  x161 &  x163 &  x167 &  x184 &  x188 &  x191 &  x194 &  x215 &  x223 &  x224 &  x235 &  x239 &  x241 &  x242 &  x263 &  x266 &  x269 &  x272 &  x275 &  x284 &  x287 &  x290 &  x293 &  x299 &  x319 &  x332 &  x338 &  x340 &  x341 &  x347 &  x352 &  x368 &  x377 &  x380 &  x383 &  x391 &  x397 &  x398 &  x410 &  x425 &  x428 &  x431 &  x434 &  x443 &  x446 &  x452 &  x457 &  x461 &  x464 &  x473 &  x479 &  x506 &  x515 &  x518 &  x524 &  x533 &  x542 &  x551 &  x557 &  x563 &  x566 &  x572 &  x575 &  x587 &  x599 &  x605 &  x608 &  x611 &  x623 &  x629 &  x632 &  x647 &  x650 &  x653 &  x659 &  x662 &  x668 &  x674 &  x677 &  x680 &  x683 &  x689 &  x692 &  x695 &  x701 &  x704 &  x707 &  x713 &  x725 &  x728 &  x731 &  x737 &  x740 &  x752 &  x763 &  x764 &  x767 &  x770 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x802 &  x818 &  x824 &  x830 &  x841 &  x842 &  x845 &  x851 &  x854 &  x866 &  x878 &  x902 &  x908 &  x916 &  x920 &  x923 &  x929 &  x947 &  x950 &  x956 &  x962 &  x965 &  x974 &  x994 &  x995 &  x998 &  x1001 &  x1004 &  x1013 &  x1022 &  x1028 &  x1034 &  x1043 &  x1049 &  x1058 &  x1073 &  x1076 &  x1079 &  x1085 &  x1091 &  x1097 &  x1103 &  x1112 &  x1118 &  x1121 &  x1127 &  x1130;
assign c582 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x26 &  x29 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x107 &  x110 &  x113 &  x116 &  x122 &  x128 &  x131 &  x137 &  x140 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x172 &  x173 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x211 &  x212 &  x215 &  x218 &  x230 &  x233 &  x235 &  x236 &  x239 &  x245 &  x250 &  x251 &  x257 &  x263 &  x266 &  x274 &  x275 &  x281 &  x284 &  x289 &  x290 &  x293 &  x296 &  x299 &  x305 &  x308 &  x311 &  x313 &  x314 &  x317 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x352 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x380 &  x389 &  x391 &  x395 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x425 &  x430 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x469 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x491 &  x500 &  x503 &  x506 &  x508 &  x509 &  x512 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x542 &  x545 &  x547 &  x548 &  x551 &  x554 &  x557 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x625 &  x626 &  x629 &  x635 &  x644 &  x647 &  x650 &  x656 &  x659 &  x662 &  x665 &  x668 &  x674 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x758 &  x761 &  x767 &  x776 &  x779 &  x785 &  x788 &  x791 &  x794 &  x797 &  x803 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x905 &  x908 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x934 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x959 &  x962 &  x965 &  x971 &  x974 &  x977 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1130 & ~x237 & ~x276 & ~x277 & ~x315 & ~x597;
assign c584 =  x2 &  x5 &  x20 &  x26 &  x35 &  x38 &  x47 &  x52 &  x62 &  x65 &  x86 &  x92 &  x128 &  x134 &  x155 &  x169 &  x176 &  x182 &  x191 &  x200 &  x206 &  x212 &  x230 &  x242 &  x257 &  x278 &  x281 &  x296 &  x314 &  x329 &  x380 &  x392 &  x404 &  x416 &  x419 &  x425 &  x437 &  x440 &  x446 &  x449 &  x452 &  x455 &  x461 &  x467 &  x473 &  x476 &  x479 &  x491 &  x497 &  x500 &  x512 &  x521 &  x530 &  x533 &  x566 &  x569 &  x578 &  x580 &  x590 &  x596 &  x617 &  x626 &  x650 &  x653 &  x656 &  x659 &  x665 &  x680 &  x683 &  x686 &  x695 &  x713 &  x719 &  x724 &  x728 &  x737 &  x746 &  x755 &  x761 &  x776 &  x779 &  x781 &  x791 &  x797 &  x815 &  x820 &  x833 &  x845 &  x851 &  x857 &  x869 &  x881 &  x890 &  x893 &  x896 &  x923 &  x938 &  x940 &  x944 &  x953 &  x970 &  x998 &  x1001 &  x1013 &  x1019 &  x1031 &  x1040 &  x1043 &  x1048 &  x1055 &  x1057 &  x1061 &  x1064 &  x1088 &  x1103 &  x1106 &  x1118 &  x1121 &  x1127 & ~x315 & ~x798;
assign c586 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x26 &  x29 &  x35 &  x38 &  x44 &  x47 &  x50 &  x53 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x89 &  x92 &  x95 &  x110 &  x116 &  x119 &  x122 &  x125 &  x131 &  x140 &  x143 &  x149 &  x152 &  x158 &  x161 &  x164 &  x170 &  x173 &  x179 &  x182 &  x188 &  x191 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x254 &  x257 &  x260 &  x263 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x293 &  x296 &  x302 &  x308 &  x311 &  x314 &  x317 &  x320 &  x326 &  x329 &  x335 &  x338 &  x341 &  x347 &  x350 &  x356 &  x359 &  x362 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x398 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x467 &  x470 &  x476 &  x479 &  x482 &  x488 &  x491 &  x494 &  x497 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x547 &  x548 &  x551 &  x560 &  x563 &  x566 &  x572 &  x575 &  x578 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x617 &  x620 &  x623 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x662 &  x665 &  x667 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x698 &  x701 &  x704 &  x706 &  x707 &  x710 &  x722 &  x728 &  x731 &  x734 &  x737 &  x740 &  x745 &  x746 &  x749 &  x752 &  x758 &  x761 &  x764 &  x767 &  x773 &  x776 &  x779 &  x782 &  x784 &  x788 &  x791 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x869 &  x875 &  x881 &  x893 &  x896 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x929 &  x938 &  x941 &  x944 &  x947 &  x953 &  x962 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x237 & ~x276 & ~x315 & ~x316 & ~x354 & ~x355 & ~x375 & ~x414 & ~x453 & ~x678;
assign c588 =  x5 &  x8 &  x11 &  x17 &  x20 &  x23 &  x29 &  x32 &  x38 &  x44 &  x47 &  x53 &  x59 &  x68 &  x71 &  x74 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x110 &  x116 &  x119 &  x122 &  x123 &  x124 &  x131 &  x134 &  x149 &  x152 &  x158 &  x161 &  x163 &  x167 &  x173 &  x176 &  x200 &  x202 &  x203 &  x209 &  x212 &  x233 &  x239 &  x242 &  x245 &  x248 &  x263 &  x266 &  x269 &  x275 &  x278 &  x280 &  x284 &  x287 &  x290 &  x296 &  x299 &  x302 &  x308 &  x311 &  x319 &  x320 &  x326 &  x338 &  x341 &  x344 &  x350 &  x356 &  x358 &  x368 &  x371 &  x374 &  x389 &  x410 &  x416 &  x419 &  x434 &  x440 &  x443 &  x446 &  x449 &  x458 &  x461 &  x467 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x527 &  x530 &  x536 &  x548 &  x563 &  x569 &  x572 &  x584 &  x614 &  x617 &  x623 &  x626 &  x638 &  x641 &  x659 &  x662 &  x668 &  x674 &  x677 &  x686 &  x689 &  x692 &  x698 &  x701 &  x713 &  x719 &  x725 &  x737 &  x746 &  x749 &  x752 &  x758 &  x766 &  x770 &  x776 &  x782 &  x794 &  x803 &  x805 &  x806 &  x815 &  x818 &  x824 &  x827 &  x830 &  x833 &  x842 &  x844 &  x845 &  x854 &  x860 &  x875 &  x878 &  x881 &  x883 &  x887 &  x893 &  x908 &  x922 &  x929 &  x935 &  x941 &  x947 &  x953 &  x965 &  x971 &  x980 &  x986 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1013 &  x1037 &  x1039 &  x1043 &  x1045 &  x1055 &  x1079 &  x1088 &  x1100 &  x1112 &  x1115 &  x1118 &  x1121;
assign c590 =  x2 &  x7 &  x8 &  x16 &  x20 &  x41 &  x47 &  x62 &  x65 &  x74 &  x80 &  x83 &  x86 &  x92 &  x98 &  x101 &  x107 &  x113 &  x119 &  x125 &  x134 &  x139 &  x140 &  x146 &  x152 &  x155 &  x158 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x212 &  x218 &  x221 &  x235 &  x239 &  x242 &  x251 &  x257 &  x260 &  x263 &  x269 &  x274 &  x278 &  x287 &  x293 &  x308 &  x313 &  x323 &  x326 &  x329 &  x374 &  x377 &  x386 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x440 &  x446 &  x452 &  x457 &  x458 &  x467 &  x473 &  x488 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x527 &  x536 &  x545 &  x548 &  x560 &  x563 &  x569 &  x572 &  x574 &  x581 &  x587 &  x605 &  x620 &  x649 &  x655 &  x656 &  x659 &  x677 &  x692 &  x694 &  x704 &  x716 &  x724 &  x725 &  x728 &  x761 &  x763 &  x767 &  x776 &  x815 &  x818 &  x827 &  x830 &  x842 &  x850 &  x851 &  x854 &  x869 &  x872 &  x881 &  x884 &  x887 &  x890 &  x893 &  x902 &  x914 &  x950 &  x962 &  x977 &  x983 &  x998 &  x1007 &  x1010 &  x1013 &  x1016 &  x1034 &  x1040 &  x1046 &  x1049 &  x1058 &  x1067 &  x1070 &  x1088 &  x1091 &  x1097 &  x1103 &  x1109 &  x1115 & ~x207;
assign c592 =  x53 &  x71 &  x74 &  x80 &  x86 &  x89 &  x116 &  x155 &  x179 &  x182 &  x194 &  x203 &  x224 &  x236 &  x254 &  x272 &  x314 &  x320 &  x329 &  x332 &  x347 &  x356 &  x371 &  x383 &  x386 &  x413 &  x416 &  x422 &  x464 &  x470 &  x479 &  x491 &  x509 &  x518 &  x557 &  x602 &  x620 &  x632 &  x656 &  x683 &  x689 &  x695 &  x698 &  x725 &  x740 &  x770 &  x791 &  x797 &  x806 &  x809 &  x833 &  x848 &  x863 &  x884 &  x896 &  x905 &  x923 &  x929 &  x947 &  x968 &  x977 &  x1017 &  x1049 &  x1093 &  x1096 &  x1097 &  x1100 &  x1118 &  x1121 &  x1124 & ~x312 & ~x468 & ~x549 & ~x628 & ~x777 & ~x849 & ~x870 & ~x909 & ~x948;
assign c594 =  x23 &  x26 &  x140 &  x251 &  x311 &  x332 &  x395 &  x575 &  x611 &  x683 &  x709 &  x719 &  x858 &  x986 &  x1057 & ~x438 & ~x706;
assign c596 =  x16 &  x17 &  x26 &  x28 &  x34 &  x53 &  x68 &  x71 &  x72 &  x83 &  x101 &  x107 &  x110 &  x122 &  x128 &  x149 &  x161 &  x173 &  x176 &  x178 &  x182 &  x191 &  x227 &  x248 &  x263 &  x266 &  x284 &  x290 &  x301 &  x305 &  x308 &  x311 &  x317 &  x323 &  x338 &  x356 &  x359 &  x380 &  x385 &  x449 &  x458 &  x461 &  x476 &  x554 &  x557 &  x562 &  x568 &  x584 &  x593 &  x607 &  x614 &  x617 &  x632 &  x635 &  x652 &  x653 &  x656 &  x657 &  x659 &  x674 &  x686 &  x695 &  x710 &  x728 &  x734 &  x749 &  x758 &  x763 &  x764 &  x785 &  x791 &  x797 &  x824 &  x830 &  x836 &  x842 &  x863 &  x872 &  x892 &  x935 &  x938 &  x944 &  x959 &  x974 &  x998 &  x1001 &  x1010 &  x1016 &  x1019 &  x1031 &  x1034 &  x1046 &  x1055 &  x1070 &  x1073 &  x1076 &  x1079 &  x1088 &  x1097 &  x1103 &  x1109 &  x1118 &  x1120 &  x1121;
assign c598 =  x5 &  x8 &  x14 &  x17 &  x20 &  x26 &  x29 &  x38 &  x44 &  x50 &  x53 &  x56 &  x65 &  x68 &  x74 &  x77 &  x80 &  x86 &  x92 &  x98 &  x104 &  x107 &  x110 &  x119 &  x122 &  x128 &  x131 &  x134 &  x140 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x185 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x218 &  x221 &  x227 &  x230 &  x233 &  x239 &  x242 &  x245 &  x251 &  x254 &  x260 &  x263 &  x266 &  x272 &  x275 &  x278 &  x281 &  x284 &  x299 &  x305 &  x308 &  x311 &  x314 &  x317 &  x323 &  x326 &  x329 &  x341 &  x347 &  x350 &  x356 &  x359 &  x362 &  x374 &  x377 &  x383 &  x389 &  x392 &  x395 &  x398 &  x401 &  x407 &  x410 &  x422 &  x428 &  x434 &  x452 &  x455 &  x458 &  x461 &  x464 &  x470 &  x473 &  x479 &  x482 &  x485 &  x488 &  x491 &  x497 &  x506 &  x515 &  x518 &  x521 &  x530 &  x533 &  x536 &  x539 &  x542 &  x548 &  x551 &  x554 &  x560 &  x563 &  x566 &  x569 &  x578 &  x587 &  x590 &  x599 &  x611 &  x613 &  x617 &  x620 &  x626 &  x632 &  x635 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x680 &  x686 &  x701 &  x713 &  x716 &  x722 &  x731 &  x734 &  x740 &  x743 &  x746 &  x752 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x781 &  x782 &  x785 &  x788 &  x791 &  x794 &  x803 &  x806 &  x812 &  x815 &  x818 &  x819 &  x820 &  x821 &  x827 &  x830 &  x833 &  x839 &  x842 &  x845 &  x857 &  x859 &  x860 &  x863 &  x866 &  x869 &  x872 &  x878 &  x884 &  x890 &  x896 &  x899 &  x902 &  x905 &  x911 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x937 &  x938 &  x941 &  x947 &  x950 &  x953 &  x962 &  x965 &  x968 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1013 &  x1019 &  x1022 &  x1028 &  x1031 &  x1037 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1070 &  x1076 &  x1082 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1118 &  x1124 &  x1127 & ~x549 & ~x588 & ~x589 & ~x621 & ~x627 & ~x660 & ~x699 & ~x837 & ~x876 & ~x915 & ~x948 & ~x1029 & ~x1068;
assign c5100 =  x8 &  x26 &  x32 &  x35 &  x47 &  x53 &  x59 &  x62 &  x68 &  x86 &  x89 &  x101 &  x104 &  x113 &  x116 &  x119 &  x128 &  x134 &  x140 &  x143 &  x146 &  x152 &  x155 &  x158 &  x161 &  x164 &  x173 &  x176 &  x182 &  x194 &  x197 &  x206 &  x209 &  x212 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x239 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x266 &  x272 &  x275 &  x278 &  x281 &  x287 &  x290 &  x293 &  x299 &  x317 &  x338 &  x346 &  x347 &  x359 &  x362 &  x365 &  x371 &  x377 &  x380 &  x385 &  x389 &  x392 &  x395 &  x413 &  x416 &  x419 &  x431 &  x434 &  x440 &  x443 &  x446 &  x458 &  x461 &  x464 &  x469 &  x470 &  x476 &  x485 &  x494 &  x500 &  x508 &  x509 &  x515 &  x518 &  x527 &  x530 &  x533 &  x536 &  x539 &  x545 &  x551 &  x557 &  x566 &  x575 &  x581 &  x584 &  x590 &  x599 &  x602 &  x611 &  x614 &  x626 &  x629 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x689 &  x692 &  x701 &  x704 &  x710 &  x719 &  x725 &  x728 &  x731 &  x734 &  x740 &  x749 &  x752 &  x755 &  x761 &  x764 &  x767 &  x770 &  x776 &  x779 &  x782 &  x785 &  x788 &  x794 &  x809 &  x812 &  x821 &  x824 &  x827 &  x833 &  x839 &  x842 &  x848 &  x851 &  x854 &  x857 &  x863 &  x869 &  x872 &  x875 &  x884 &  x890 &  x896 &  x905 &  x911 &  x914 &  x920 &  x929 &  x932 &  x947 &  x950 &  x962 &  x983 &  x986 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1022 &  x1031 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1067 &  x1070 &  x1076 &  x1079 &  x1088 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1124 &  x1127 &  x1130 & ~x237 & ~x277 & ~x315 & ~x426 & ~x427 & ~x465 & ~x564;
assign c5102 =  x5 &  x35 &  x38 &  x47 &  x53 &  x59 &  x65 &  x74 &  x83 &  x86 &  x98 &  x101 &  x107 &  x137 &  x143 &  x149 &  x155 &  x161 &  x179 &  x185 &  x197 &  x200 &  x212 &  x215 &  x221 &  x230 &  x236 &  x248 &  x254 &  x257 &  x260 &  x269 &  x272 &  x275 &  x281 &  x287 &  x308 &  x314 &  x320 &  x323 &  x332 &  x335 &  x338 &  x341 &  x365 &  x392 &  x407 &  x410 &  x425 &  x434 &  x446 &  x467 &  x476 &  x479 &  x485 &  x491 &  x500 &  x509 &  x515 &  x518 &  x523 &  x527 &  x530 &  x539 &  x545 &  x561 &  x566 &  x569 &  x572 &  x590 &  x599 &  x605 &  x608 &  x611 &  x617 &  x629 &  x635 &  x647 &  x656 &  x665 &  x668 &  x671 &  x692 &  x695 &  x701 &  x704 &  x713 &  x722 &  x725 &  x728 &  x734 &  x737 &  x761 &  x764 &  x770 &  x776 &  x779 &  x781 &  x782 &  x788 &  x791 &  x797 &  x806 &  x820 &  x824 &  x845 &  x851 &  x857 &  x859 &  x872 &  x878 &  x893 &  x899 &  x902 &  x911 &  x932 &  x941 &  x947 &  x965 &  x980 &  x989 &  x992 &  x1007 &  x1010 &  x1019 &  x1025 &  x1034 &  x1046 &  x1049 &  x1055 &  x1064 &  x1070 &  x1073 &  x1076 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1112 &  x1115 &  x1121 & ~x273 & ~x351 & ~x471 & ~x510 & ~x550 & ~x675 & ~x714 & ~x792;
assign c5104 =  x5 &  x8 &  x11 &  x14 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x40 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x77 &  x80 &  x83 &  x98 &  x101 &  x107 &  x110 &  x113 &  x116 &  x118 &  x119 &  x125 &  x128 &  x131 &  x137 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x176 &  x179 &  x182 &  x188 &  x191 &  x194 &  x196 &  x197 &  x200 &  x206 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x235 &  x236 &  x242 &  x248 &  x251 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x320 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x380 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x455 &  x458 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x491 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x572 &  x575 &  x578 &  x581 &  x584 &  x590 &  x599 &  x605 &  x608 &  x610 &  x611 &  x614 &  x617 &  x623 &  x626 &  x632 &  x635 &  x644 &  x647 &  x649 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x674 &  x677 &  x680 &  x683 &  x686 &  x688 &  x689 &  x695 &  x698 &  x704 &  x707 &  x713 &  x716 &  x719 &  x722 &  x725 &  x727 &  x728 &  x731 &  x734 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x764 &  x770 &  x773 &  x776 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x812 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x850 &  x851 &  x854 &  x860 &  x863 &  x866 &  x869 &  x875 &  x878 &  x881 &  x887 &  x890 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x950 &  x953 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 & ~x42 & ~x81 & ~x225 & ~x252 & ~x291 & ~x324 & ~x330 & ~x369 & ~x444 & ~x483 & ~x522 & ~x600 & ~x633 & ~x711;
assign c5106 =  x122 &  x173 &  x194 &  x248 &  x260 &  x284 &  x302 &  x359 &  x365 &  x380 &  x474 &  x506 &  x553 &  x632 &  x641 &  x703 &  x788 &  x830 &  x863 &  x901 &  x929 &  x938 &  x1043 &  x1097 & ~x511;
assign c5108 =  x269 &  x337 &  x386 &  x618 &  x670 &  x671 &  x722 &  x724 &  x757 &  x775 &  x853 &  x887 &  x892 &  x969 &  x998 &  x1073 &  x1085 &  x1093;
assign c5110 =  x2 &  x5 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x128 &  x131 &  x134 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x479 &  x482 &  x485 &  x491 &  x494 &  x497 &  x500 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x571 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x602 &  x605 &  x608 &  x610 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x644 &  x649 &  x650 &  x653 &  x656 &  x659 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x688 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x725 &  x728 &  x731 &  x734 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x788 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x821 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x911 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x961 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1000 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x42 & ~x51 & ~x81 & ~x82 & ~x291 & ~x292 & ~x324 & ~x330 & ~x370 & ~x408;
assign c5112 =  x26 &  x35 &  x97 &  x98 &  x101 &  x107 &  x110 &  x119 &  x125 &  x137 &  x140 &  x143 &  x146 &  x152 &  x164 &  x167 &  x185 &  x191 &  x203 &  x215 &  x224 &  x230 &  x251 &  x278 &  x281 &  x290 &  x296 &  x302 &  x305 &  x311 &  x332 &  x335 &  x380 &  x383 &  x407 &  x413 &  x422 &  x440 &  x449 &  x473 &  x488 &  x491 &  x494 &  x500 &  x572 &  x575 &  x602 &  x605 &  x608 &  x620 &  x623 &  x626 &  x629 &  x632 &  x653 &  x656 &  x662 &  x665 &  x668 &  x698 &  x713 &  x722 &  x725 &  x731 &  x737 &  x749 &  x770 &  x773 &  x791 &  x797 &  x803 &  x809 &  x821 &  x830 &  x836 &  x861 &  x875 &  x878 &  x890 &  x901 &  x902 &  x905 &  x911 &  x917 &  x923 &  x932 &  x941 &  x950 &  x956 &  x959 &  x962 &  x965 &  x986 &  x995 &  x998 &  x1004 &  x1007 &  x1025 &  x1028 &  x1046 &  x1055 &  x1058 &  x1070 &  x1073 &  x1097 &  x1100 &  x1109 &  x1112 &  x1115 & ~x312 & ~x480 & ~x675 & ~x720 & ~x798 & ~x1068;
assign c5114 =  x1 &  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x29 &  x32 &  x35 &  x41 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x77 &  x79 &  x80 &  x83 &  x86 &  x89 &  x92 &  x98 &  x101 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x155 &  x157 &  x158 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x235 &  x236 &  x239 &  x245 &  x248 &  x251 &  x254 &  x257 &  x263 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x311 &  x313 &  x314 &  x317 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x344 &  x347 &  x350 &  x353 &  x359 &  x362 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x389 &  x394 &  x395 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x432 &  x433 &  x434 &  x437 &  x443 &  x446 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x472 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x506 &  x511 &  x512 &  x515 &  x521 &  x524 &  x527 &  x533 &  x536 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x626 &  x629 &  x632 &  x638 &  x641 &  x644 &  x647 &  x653 &  x662 &  x665 &  x671 &  x674 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x701 &  x707 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x734 &  x737 &  x743 &  x746 &  x752 &  x755 &  x758 &  x764 &  x767 &  x770 &  x776 &  x779 &  x785 &  x791 &  x794 &  x797 &  x800 &  x806 &  x821 &  x827 &  x830 &  x836 &  x848 &  x851 &  x854 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x905 &  x908 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x938 &  x944 &  x947 &  x950 &  x953 &  x959 &  x962 &  x971 &  x974 &  x977 &  x980 &  x983 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x207 & ~x264 & ~x303 & ~x546 & ~x585 & ~x633 & ~x672 & ~x789 & ~x828;
assign c5116 =  x2 &  x17 &  x23 &  x26 &  x89 &  x101 &  x107 &  x110 &  x116 &  x122 &  x134 &  x146 &  x158 &  x197 &  x206 &  x209 &  x215 &  x242 &  x248 &  x254 &  x293 &  x299 &  x311 &  x317 &  x320 &  x338 &  x341 &  x359 &  x362 &  x374 &  x380 &  x389 &  x401 &  x422 &  x431 &  x440 &  x446 &  x449 &  x455 &  x467 &  x473 &  x476 &  x479 &  x491 &  x497 &  x503 &  x512 &  x514 &  x518 &  x527 &  x539 &  x545 &  x548 &  x572 &  x578 &  x584 &  x590 &  x617 &  x620 &  x635 &  x644 &  x656 &  x671 &  x683 &  x719 &  x728 &  x749 &  x755 &  x767 &  x773 &  x779 &  x782 &  x785 &  x788 &  x791 &  x797 &  x800 &  x818 &  x836 &  x881 &  x898 &  x917 &  x935 &  x940 &  x947 &  x950 &  x962 &  x965 &  x971 &  x995 &  x1034 &  x1052 &  x1058 &  x1067 &  x1073 &  x1085 &  x1096 &  x1112 &  x1118 &  x1121 & ~x312 & ~x510 & ~x588 & ~x628 & ~x675 & ~x831 & ~x954;
assign c5118 =  x8 &  x44 &  x50 &  x56 &  x61 &  x110 &  x134 &  x175 &  x185 &  x230 &  x233 &  x239 &  x242 &  x326 &  x344 &  x410 &  x443 &  x494 &  x503 &  x506 &  x529 &  x539 &  x545 &  x566 &  x569 &  x616 &  x620 &  x647 &  x695 &  x698 &  x728 &  x731 &  x836 &  x854 &  x884 &  x887 &  x892 &  x893 &  x938 &  x956 &  x983 &  x995 &  x998 &  x1010 &  x1018 &  x1040 &  x1097 & ~x276 & ~x906;
assign c5120 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x23 &  x29 &  x32 &  x35 &  x38 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x119 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x230 &  x233 &  x235 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x274 &  x275 &  x278 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x314 &  x317 &  x320 &  x326 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x352 &  x356 &  x365 &  x368 &  x377 &  x380 &  x383 &  x386 &  x391 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x428 &  x431 &  x434 &  x437 &  x440 &  x449 &  x452 &  x458 &  x461 &  x467 &  x469 &  x470 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x508 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x584 &  x587 &  x589 &  x590 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x628 &  x629 &  x632 &  x635 &  x641 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x818 &  x821 &  x824 &  x827 &  x833 &  x842 &  x845 &  x848 &  x851 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x893 &  x896 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x932 &  x935 &  x941 &  x944 &  x947 &  x950 &  x953 &  x959 &  x962 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1037 &  x1040 &  x1043 &  x1046 &  x1055 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1097 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x238 & ~x483 & ~x522 & ~x523 & ~x561 & ~x562 & ~x600 & ~x639;
assign c5122 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x83 &  x86 &  x89 &  x92 &  x95 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x157 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x308 &  x311 &  x313 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x394 &  x395 &  x398 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x440 &  x443 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x512 &  x515 &  x518 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x587 &  x593 &  x596 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x830 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x971 &  x977 &  x980 &  x983 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130 & ~x3 & ~x12 & ~x42 & ~x43 & ~x51 & ~x81 & ~x90 & ~x91 & ~x129 & ~x168 & ~x169 & ~x246 & ~x285 & ~x324 & ~x363 & ~x585 & ~x663 & ~x702 & ~x741 & ~x780 & ~x819 & ~x858 & ~x897 & ~x936 & ~x975 & ~x1014 & ~x1053 & ~x1092;
assign c5124 =  x5 &  x8 &  x11 &  x20 &  x26 &  x32 &  x62 &  x83 &  x86 &  x92 &  x95 &  x98 &  x125 &  x137 &  x140 &  x143 &  x149 &  x158 &  x161 &  x164 &  x170 &  x173 &  x176 &  x179 &  x185 &  x188 &  x194 &  x197 &  x200 &  x206 &  x209 &  x218 &  x221 &  x227 &  x230 &  x233 &  x239 &  x245 &  x248 &  x254 &  x263 &  x275 &  x281 &  x284 &  x296 &  x311 &  x314 &  x350 &  x353 &  x356 &  x368 &  x377 &  x380 &  x401 &  x404 &  x407 &  x410 &  x419 &  x425 &  x428 &  x437 &  x443 &  x445 &  x455 &  x458 &  x464 &  x482 &  x485 &  x497 &  x500 &  x503 &  x514 &  x523 &  x530 &  x533 &  x539 &  x542 &  x548 &  x553 &  x554 &  x560 &  x563 &  x566 &  x575 &  x587 &  x593 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x629 &  x638 &  x641 &  x662 &  x665 &  x668 &  x671 &  x686 &  x695 &  x707 &  x713 &  x716 &  x725 &  x734 &  x737 &  x740 &  x742 &  x746 &  x752 &  x761 &  x779 &  x781 &  x782 &  x785 &  x788 &  x806 &  x812 &  x820 &  x821 &  x824 &  x836 &  x839 &  x842 &  x845 &  x854 &  x859 &  x863 &  x875 &  x878 &  x884 &  x887 &  x893 &  x911 &  x914 &  x920 &  x932 &  x938 &  x941 &  x944 &  x950 &  x953 &  x956 &  x959 &  x968 &  x983 &  x989 &  x992 &  x998 &  x1007 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1054 &  x1055 &  x1076 &  x1079 &  x1082 &  x1103 &  x1118 &  x1127 &  x1130 & ~x315 & ~x393 & ~x471 & ~x486 & ~x549 & ~x687 & ~x714 & ~x831;
assign c5126 =  x20 &  x26 &  x29 &  x32 &  x41 &  x56 &  x65 &  x68 &  x77 &  x80 &  x83 &  x86 &  x92 &  x110 &  x113 &  x125 &  x128 &  x140 &  x155 &  x167 &  x173 &  x188 &  x194 &  x206 &  x209 &  x233 &  x239 &  x242 &  x254 &  x257 &  x269 &  x278 &  x280 &  x293 &  x296 &  x302 &  x305 &  x323 &  x335 &  x345 &  x359 &  x368 &  x371 &  x380 &  x389 &  x398 &  x401 &  x410 &  x419 &  x425 &  x431 &  x434 &  x443 &  x482 &  x485 &  x491 &  x506 &  x509 &  x512 &  x521 &  x533 &  x551 &  x560 &  x572 &  x578 &  x590 &  x608 &  x614 &  x626 &  x635 &  x644 &  x647 &  x659 &  x665 &  x671 &  x674 &  x689 &  x692 &  x728 &  x731 &  x737 &  x764 &  x779 &  x782 &  x809 &  x812 &  x833 &  x842 &  x860 &  x863 &  x866 &  x869 &  x884 &  x887 &  x893 &  x896 &  x905 &  x917 &  x926 &  x947 &  x983 &  x992 &  x1034 &  x1052 &  x1055 &  x1061 &  x1067 &  x1076 &  x1085 &  x1094 &  x1115 & ~x237 & ~x354 & ~x375 & ~x519 & ~x558 & ~x714;
assign c5128 =  x8 &  x110 &  x233 &  x323 &  x419 &  x581 &  x617 &  x743 &  x797 &  x830 &  x863 & ~x355 & ~x427;
assign c5130 =  x2 &  x5 &  x11 &  x14 &  x20 &  x26 &  x29 &  x32 &  x35 &  x41 &  x44 &  x47 &  x50 &  x53 &  x59 &  x62 &  x65 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x101 &  x104 &  x107 &  x110 &  x116 &  x118 &  x119 &  x125 &  x128 &  x131 &  x137 &  x143 &  x146 &  x149 &  x164 &  x167 &  x170 &  x176 &  x185 &  x188 &  x191 &  x194 &  x196 &  x197 &  x200 &  x209 &  x212 &  x215 &  x218 &  x221 &  x227 &  x230 &  x233 &  x235 &  x236 &  x239 &  x242 &  x245 &  x248 &  x254 &  x257 &  x263 &  x266 &  x269 &  x272 &  x274 &  x275 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x311 &  x312 &  x313 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x347 &  x350 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x391 &  x392 &  x395 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x437 &  x443 &  x449 &  x452 &  x458 &  x461 &  x467 &  x470 &  x472 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x500 &  x503 &  x512 &  x515 &  x518 &  x521 &  x524 &  x530 &  x533 &  x536 &  x542 &  x545 &  x548 &  x550 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x587 &  x590 &  x593 &  x596 &  x602 &  x605 &  x608 &  x614 &  x617 &  x620 &  x623 &  x629 &  x635 &  x638 &  x641 &  x650 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x688 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x713 &  x719 &  x722 &  x725 &  x727 &  x728 &  x734 &  x737 &  x740 &  x749 &  x755 &  x758 &  x761 &  x764 &  x766 &  x770 &  x773 &  x776 &  x779 &  x782 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x812 &  x821 &  x824 &  x830 &  x836 &  x839 &  x842 &  x848 &  x851 &  x857 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x890 &  x896 &  x902 &  x911 &  x914 &  x917 &  x920 &  x923 &  x935 &  x938 &  x941 &  x944 &  x953 &  x956 &  x959 &  x962 &  x965 &  x974 &  x977 &  x980 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1034 &  x1037 &  x1043 &  x1052 &  x1055 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x42 & ~x81 & ~x120 & ~x121 & ~x159 & ~x246 & ~x303 & ~x363;
assign c5132 =  x11 &  x13 &  x17 &  x20 &  x34 &  x52 &  x53 &  x61 &  x73 &  x92 &  x98 &  x100 &  x101 &  x104 &  x116 &  x119 &  x128 &  x131 &  x137 &  x143 &  x152 &  x155 &  x170 &  x178 &  x179 &  x182 &  x190 &  x206 &  x212 &  x230 &  x245 &  x263 &  x268 &  x281 &  x284 &  x287 &  x293 &  x305 &  x307 &  x317 &  x323 &  x335 &  x344 &  x356 &  x368 &  x374 &  x383 &  x385 &  x386 &  x392 &  x398 &  x416 &  x425 &  x431 &  x434 &  x440 &  x446 &  x449 &  x458 &  x467 &  x485 &  x488 &  x491 &  x497 &  x500 &  x506 &  x512 &  x521 &  x524 &  x533 &  x542 &  x560 &  x602 &  x608 &  x614 &  x620 &  x632 &  x638 &  x641 &  x650 &  x662 &  x671 &  x677 &  x683 &  x695 &  x701 &  x704 &  x713 &  x719 &  x739 &  x743 &  x749 &  x764 &  x776 &  x779 &  x800 &  x803 &  x815 &  x827 &  x836 &  x857 &  x862 &  x863 &  x866 &  x872 &  x875 &  x887 &  x901 &  x902 &  x914 &  x920 &  x929 &  x932 &  x934 &  x941 &  x953 &  x959 &  x965 &  x992 &  x1001 &  x1013 &  x1031 &  x1036 &  x1043 &  x1046 &  x1061 &  x1067 &  x1094 &  x1097 &  x1109 &  x1112 &  x1115 &  x1124;
assign c5134 =  x2 &  x5 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x476 &  x479 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x626 &  x632 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x701 &  x704 &  x707 &  x710 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x794 &  x800 &  x803 &  x806 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x857 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x159 & ~x198 & ~x199 & ~x237 & ~x276 & ~x369 & ~x402 & ~x441 & ~x486 & ~x519 & ~x525 & ~x1053 & ~x1068 & ~x1107;
assign c5136 =  x2 &  x14 &  x17 &  x23 &  x35 &  x38 &  x47 &  x50 &  x53 &  x56 &  x62 &  x68 &  x71 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x122 &  x134 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x167 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x242 &  x245 &  x254 &  x257 &  x260 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x293 &  x296 &  x299 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x332 &  x335 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x437 &  x443 &  x446 &  x449 &  x455 &  x461 &  x464 &  x467 &  x473 &  x479 &  x482 &  x485 &  x488 &  x494 &  x497 &  x500 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x587 &  x590 &  x593 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x628 &  x629 &  x632 &  x635 &  x638 &  x641 &  x647 &  x650 &  x653 &  x656 &  x665 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x692 &  x701 &  x704 &  x707 &  x713 &  x716 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x743 &  x746 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x782 &  x785 &  x794 &  x797 &  x800 &  x803 &  x809 &  x812 &  x815 &  x818 &  x824 &  x827 &  x830 &  x839 &  x842 &  x845 &  x848 &  x851 &  x857 &  x863 &  x866 &  x869 &  x872 &  x878 &  x881 &  x884 &  x887 &  x893 &  x896 &  x899 &  x905 &  x908 &  x911 &  x920 &  x929 &  x932 &  x938 &  x947 &  x950 &  x953 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x983 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1028 &  x1033 &  x1034 &  x1043 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1072 &  x1073 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 & ~x0 & ~x120 & ~x160 & ~x199 & ~x246 & ~x285 & ~x324 & ~x363 & ~x402 & ~x600 & ~x639 & ~x819 & ~x897 & ~x975 & ~x1014;
assign c5138 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x59 &  x62 &  x65 &  x71 &  x77 &  x79 &  x80 &  x86 &  x92 &  x95 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x118 &  x119 &  x122 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x206 &  x209 &  x212 &  x215 &  x227 &  x230 &  x233 &  x235 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x266 &  x269 &  x272 &  x274 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x312 &  x313 &  x314 &  x317 &  x320 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x352 &  x355 &  x356 &  x359 &  x365 &  x368 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x391 &  x392 &  x394 &  x395 &  x398 &  x404 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x467 &  x470 &  x472 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x521 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x566 &  x569 &  x575 &  x578 &  x581 &  x583 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x680 &  x683 &  x686 &  x688 &  x689 &  x692 &  x695 &  x698 &  x701 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x743 &  x746 &  x749 &  x752 &  x758 &  x761 &  x764 &  x767 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1058 &  x1064 &  x1067 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x81 & ~x82 & ~x120 & ~x121 & ~x363 & ~x585 & ~x624 & ~x663 & ~x702;
assign c5140 =  x2 &  x5 &  x11 &  x14 &  x23 &  x35 &  x40 &  x50 &  x62 &  x68 &  x71 &  x74 &  x77 &  x79 &  x80 &  x83 &  x92 &  x95 &  x104 &  x107 &  x110 &  x112 &  x113 &  x116 &  x118 &  x131 &  x140 &  x146 &  x152 &  x155 &  x161 &  x164 &  x167 &  x173 &  x178 &  x179 &  x182 &  x188 &  x197 &  x209 &  x212 &  x218 &  x224 &  x230 &  x233 &  x235 &  x236 &  x242 &  x248 &  x251 &  x256 &  x260 &  x272 &  x274 &  x278 &  x284 &  x287 &  x290 &  x299 &  x302 &  x311 &  x314 &  x323 &  x332 &  x338 &  x347 &  x359 &  x362 &  x383 &  x386 &  x389 &  x395 &  x404 &  x407 &  x413 &  x416 &  x419 &  x422 &  x425 &  x434 &  x443 &  x449 &  x452 &  x455 &  x461 &  x467 &  x473 &  x485 &  x491 &  x500 &  x505 &  x515 &  x524 &  x527 &  x530 &  x548 &  x551 &  x554 &  x560 &  x563 &  x566 &  x575 &  x581 &  x583 &  x584 &  x587 &  x590 &  x599 &  x602 &  x608 &  x617 &  x620 &  x622 &  x629 &  x638 &  x641 &  x644 &  x647 &  x649 &  x650 &  x653 &  x656 &  x665 &  x668 &  x674 &  x680 &  x683 &  x695 &  x731 &  x734 &  x740 &  x749 &  x752 &  x761 &  x767 &  x776 &  x779 &  x782 &  x784 &  x785 &  x788 &  x791 &  x794 &  x800 &  x803 &  x806 &  x812 &  x815 &  x818 &  x821 &  x823 &  x827 &  x833 &  x839 &  x848 &  x850 &  x851 &  x854 &  x860 &  x869 &  x875 &  x881 &  x890 &  x893 &  x899 &  x905 &  x916 &  x917 &  x919 &  x920 &  x923 &  x932 &  x938 &  x947 &  x953 &  x955 &  x956 &  x965 &  x968 &  x971 &  x974 &  x980 &  x989 &  x994 &  x995 &  x1004 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1040 &  x1043 &  x1046 &  x1055 &  x1067 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1100 &  x1115 &  x1121 &  x1124;
assign c5142 =  x2 &  x5 &  x8 &  x11 &  x14 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x74 &  x77 &  x80 &  x83 &  x85 &  x86 &  x89 &  x92 &  x95 &  x98 &  x104 &  x107 &  x110 &  x113 &  x116 &  x122 &  x124 &  x125 &  x134 &  x143 &  x146 &  x152 &  x158 &  x161 &  x167 &  x170 &  x176 &  x185 &  x191 &  x197 &  x203 &  x212 &  x215 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x241 &  x251 &  x257 &  x260 &  x266 &  x269 &  x278 &  x280 &  x281 &  x284 &  x287 &  x290 &  x293 &  x299 &  x305 &  x314 &  x317 &  x319 &  x323 &  x326 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x362 &  x368 &  x371 &  x374 &  x377 &  x383 &  x386 &  x398 &  x404 &  x407 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x467 &  x470 &  x473 &  x476 &  x482 &  x485 &  x488 &  x500 &  x503 &  x512 &  x515 &  x518 &  x527 &  x530 &  x533 &  x539 &  x545 &  x557 &  x560 &  x563 &  x569 &  x575 &  x581 &  x584 &  x587 &  x593 &  x596 &  x599 &  x602 &  x608 &  x611 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x647 &  x650 &  x653 &  x662 &  x665 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x701 &  x704 &  x707 &  x710 &  x716 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x746 &  x752 &  x761 &  x764 &  x767 &  x772 &  x776 &  x779 &  x788 &  x797 &  x800 &  x809 &  x812 &  x815 &  x827 &  x836 &  x839 &  x842 &  x845 &  x854 &  x857 &  x863 &  x878 &  x884 &  x890 &  x893 &  x902 &  x905 &  x908 &  x911 &  x914 &  x923 &  x926 &  x929 &  x935 &  x938 &  x941 &  x944 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x977 &  x980 &  x983 &  x989 &  x992 &  x1004 &  x1007 &  x1010 &  x1028 &  x1034 &  x1043 &  x1046 &  x1049 &  x1055 &  x1061 &  x1064 &  x1067 &  x1076 &  x1079 &  x1085 &  x1088 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1127 & ~x198 & ~x237 & ~x555 & ~x633 & ~x672 & ~x711 & ~x750 & ~x828 & ~x867 & ~x1062 & ~x1101;
assign c5144 =  x2 &  x8 &  x11 &  x17 &  x32 &  x35 &  x47 &  x50 &  x65 &  x71 &  x74 &  x77 &  x83 &  x86 &  x89 &  x95 &  x101 &  x104 &  x116 &  x119 &  x122 &  x125 &  x131 &  x134 &  x143 &  x149 &  x164 &  x179 &  x200 &  x209 &  x218 &  x221 &  x224 &  x233 &  x239 &  x242 &  x245 &  x254 &  x257 &  x269 &  x275 &  x281 &  x290 &  x293 &  x302 &  x308 &  x311 &  x317 &  x326 &  x329 &  x335 &  x347 &  x353 &  x359 &  x374 &  x377 &  x380 &  x383 &  x392 &  x416 &  x419 &  x428 &  x431 &  x434 &  x449 &  x476 &  x479 &  x482 &  x488 &  x500 &  x512 &  x530 &  x533 &  x539 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x584 &  x587 &  x593 &  x605 &  x608 &  x611 &  x614 &  x623 &  x626 &  x632 &  x635 &  x638 &  x641 &  x644 &  x659 &  x671 &  x677 &  x710 &  x719 &  x725 &  x731 &  x737 &  x740 &  x743 &  x746 &  x752 &  x761 &  x767 &  x776 &  x779 &  x785 &  x791 &  x809 &  x812 &  x821 &  x824 &  x830 &  x836 &  x842 &  x848 &  x851 &  x872 &  x875 &  x890 &  x901 &  x902 &  x905 &  x908 &  x920 &  x929 &  x941 &  x962 &  x971 &  x977 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1046 &  x1049 &  x1052 &  x1058 &  x1067 &  x1070 &  x1073 &  x1076 &  x1085 &  x1088 &  x1091 &  x1094 &  x1100 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 & ~x120 & ~x159 & ~x198 & ~x276 & ~x316 & ~x375 & ~x453 & ~x492 & ~x531 & ~x678 & ~x681 & ~x720;
assign c5146 =  x2 &  x25 &  x26 &  x35 &  x53 &  x59 &  x65 &  x86 &  x119 &  x125 &  x143 &  x155 &  x167 &  x173 &  x194 &  x209 &  x212 &  x233 &  x236 &  x239 &  x248 &  x251 &  x269 &  x272 &  x284 &  x287 &  x311 &  x320 &  x338 &  x341 &  x344 &  x362 &  x365 &  x377 &  x383 &  x395 &  x422 &  x428 &  x455 &  x479 &  x491 &  x506 &  x509 &  x524 &  x530 &  x566 &  x596 &  x608 &  x632 &  x644 &  x647 &  x662 &  x674 &  x680 &  x686 &  x689 &  x713 &  x749 &  x755 &  x758 &  x764 &  x767 &  x776 &  x827 &  x848 &  x860 &  x862 &  x869 &  x872 &  x875 &  x884 &  x887 &  x890 &  x901 &  x908 &  x923 &  x962 &  x965 &  x979 &  x983 &  x989 &  x1001 &  x1004 &  x1007 &  x1010 &  x1019 &  x1022 &  x1037 &  x1070 &  x1088 &  x1094 &  x1097 &  x1103 &  x1112 &  x1121 &  x1130 & ~x87 & ~x126 & ~x165 & ~x283 & ~x390 & ~x549;
assign c5148 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x32 &  x41 &  x44 &  x53 &  x56 &  x59 &  x65 &  x68 &  x74 &  x77 &  x80 &  x89 &  x92 &  x101 &  x104 &  x107 &  x113 &  x116 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x191 &  x194 &  x197 &  x203 &  x206 &  x209 &  x218 &  x221 &  x224 &  x227 &  x230 &  x242 &  x248 &  x251 &  x254 &  x257 &  x263 &  x266 &  x269 &  x278 &  x281 &  x284 &  x293 &  x302 &  x311 &  x314 &  x317 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x350 &  x353 &  x359 &  x362 &  x365 &  x380 &  x383 &  x386 &  x389 &  x392 &  x398 &  x401 &  x404 &  x407 &  x410 &  x428 &  x434 &  x443 &  x446 &  x452 &  x454 &  x458 &  x461 &  x464 &  x476 &  x479 &  x482 &  x485 &  x491 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x521 &  x527 &  x533 &  x536 &  x542 &  x545 &  x548 &  x554 &  x557 &  x560 &  x566 &  x569 &  x575 &  x578 &  x581 &  x583 &  x584 &  x587 &  x590 &  x593 &  x599 &  x608 &  x611 &  x614 &  x617 &  x620 &  x622 &  x626 &  x629 &  x635 &  x641 &  x644 &  x647 &  x649 &  x650 &  x653 &  x659 &  x665 &  x668 &  x671 &  x674 &  x680 &  x688 &  x689 &  x692 &  x695 &  x698 &  x701 &  x707 &  x713 &  x722 &  x725 &  x727 &  x734 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x815 &  x818 &  x824 &  x830 &  x836 &  x839 &  x845 &  x848 &  x851 &  x854 &  x860 &  x863 &  x866 &  x869 &  x875 &  x878 &  x881 &  x889 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x916 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x953 &  x959 &  x965 &  x968 &  x974 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1060 &  x1061 &  x1064 &  x1067 &  x1078 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1099 &  x1103 &  x1106 &  x1109 &  x1112 &  x1117 &  x1118 &  x1121 &  x1127 & ~x42 & ~x81 & ~x102 & ~x789 & ~x858;
assign c5150 =  x2 &  x5 &  x11 &  x14 &  x17 &  x23 &  x26 &  x29 &  x32 &  x41 &  x53 &  x56 &  x59 &  x61 &  x71 &  x74 &  x77 &  x83 &  x89 &  x101 &  x107 &  x113 &  x128 &  x131 &  x137 &  x140 &  x146 &  x149 &  x152 &  x155 &  x161 &  x164 &  x167 &  x170 &  x173 &  x182 &  x185 &  x188 &  x191 &  x194 &  x203 &  x206 &  x209 &  x215 &  x221 &  x224 &  x227 &  x230 &  x236 &  x239 &  x242 &  x263 &  x269 &  x274 &  x275 &  x281 &  x284 &  x287 &  x290 &  x296 &  x302 &  x305 &  x308 &  x311 &  x317 &  x323 &  x329 &  x332 &  x335 &  x338 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x395 &  x401 &  x404 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x437 &  x440 &  x446 &  x449 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x488 &  x491 &  x503 &  x506 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x545 &  x551 &  x557 &  x563 &  x575 &  x578 &  x587 &  x590 &  x596 &  x605 &  x608 &  x611 &  x620 &  x623 &  x626 &  x638 &  x650 &  x653 &  x659 &  x665 &  x668 &  x671 &  x674 &  x677 &  x683 &  x686 &  x689 &  x707 &  x710 &  x716 &  x722 &  x725 &  x731 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x758 &  x761 &  x764 &  x773 &  x776 &  x779 &  x791 &  x797 &  x803 &  x806 &  x815 &  x818 &  x821 &  x830 &  x833 &  x836 &  x842 &  x848 &  x854 &  x866 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x896 &  x902 &  x908 &  x917 &  x920 &  x926 &  x929 &  x935 &  x941 &  x947 &  x953 &  x959 &  x965 &  x968 &  x977 &  x980 &  x986 &  x995 &  x998 &  x1004 &  x1010 &  x1019 &  x1022 &  x1028 &  x1037 &  x1046 &  x1049 &  x1052 &  x1055 &  x1067 &  x1070 &  x1073 &  x1082 &  x1088 &  x1091 &  x1097 &  x1100 &  x1106 &  x1121 &  x1124 &  x1130 & ~x3 & ~x4 & ~x42 & ~x135 & ~x174 & ~x175 & ~x207 & ~x213 & ~x291 & ~x741 & ~x780 & ~x858 & ~x897;
assign c5152 =  x8 &  x11 &  x29 &  x41 &  x53 &  x56 &  x77 &  x119 &  x131 &  x146 &  x170 &  x191 &  x212 &  x215 &  x221 &  x236 &  x257 &  x272 &  x278 &  x296 &  x308 &  x326 &  x335 &  x356 &  x368 &  x371 &  x374 &  x377 &  x380 &  x422 &  x467 &  x469 &  x485 &  x518 &  x530 &  x548 &  x584 &  x596 &  x599 &  x626 &  x632 &  x641 &  x665 &  x674 &  x683 &  x698 &  x737 &  x743 &  x749 &  x755 &  x761 &  x764 &  x788 &  x806 &  x809 &  x812 &  x821 &  x823 &  x824 &  x848 &  x863 &  x887 &  x893 &  x901 &  x908 &  x911 &  x929 &  x938 &  x953 &  x965 &  x992 &  x998 &  x1007 &  x1025 &  x1040 &  x1049 &  x1088 &  x1100 &  x1118 &  x1130 & ~x198 & ~x276 & ~x316 & ~x642 & ~x678;
assign c5154 =  x5 &  x14 &  x17 &  x20 &  x26 &  x32 &  x40 &  x44 &  x50 &  x56 &  x59 &  x65 &  x68 &  x79 &  x80 &  x86 &  x92 &  x107 &  x110 &  x113 &  x116 &  x118 &  x122 &  x128 &  x131 &  x134 &  x137 &  x140 &  x146 &  x155 &  x157 &  x158 &  x167 &  x191 &  x196 &  x215 &  x224 &  x233 &  x234 &  x235 &  x248 &  x251 &  x263 &  x266 &  x275 &  x281 &  x287 &  x293 &  x308 &  x311 &  x313 &  x314 &  x326 &  x338 &  x344 &  x347 &  x352 &  x353 &  x365 &  x368 &  x371 &  x377 &  x386 &  x394 &  x401 &  x404 &  x407 &  x410 &  x419 &  x428 &  x434 &  x449 &  x452 &  x458 &  x464 &  x467 &  x479 &  x485 &  x488 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x524 &  x527 &  x533 &  x548 &  x551 &  x572 &  x578 &  x599 &  x614 &  x620 &  x623 &  x626 &  x647 &  x653 &  x656 &  x665 &  x671 &  x674 &  x683 &  x689 &  x698 &  x701 &  x719 &  x722 &  x725 &  x728 &  x743 &  x746 &  x749 &  x755 &  x767 &  x770 &  x773 &  x779 &  x803 &  x812 &  x818 &  x833 &  x839 &  x842 &  x845 &  x848 &  x854 &  x857 &  x863 &  x869 &  x872 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x920 &  x932 &  x941 &  x944 &  x947 &  x962 &  x968 &  x983 &  x992 &  x995 &  x1010 &  x1013 &  x1016 &  x1022 &  x1028 &  x1034 &  x1043 &  x1058 &  x1064 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1097 &  x1103 &  x1109 &  x1112 &  x1130 & ~x3 & ~x4 & ~x42 & ~x90 & ~x129 & ~x148 & ~x180 & ~x405 & ~x444 & ~x663 & ~x780 & ~x819 & ~x897;
assign c5156 =  x20 &  x44 &  x50 &  x58 &  x71 &  x80 &  x92 &  x95 &  x103 &  x119 &  x131 &  x134 &  x140 &  x143 &  x149 &  x161 &  x167 &  x176 &  x203 &  x206 &  x212 &  x227 &  x245 &  x254 &  x260 &  x263 &  x278 &  x281 &  x302 &  x311 &  x320 &  x329 &  x350 &  x353 &  x368 &  x392 &  x431 &  x437 &  x446 &  x470 &  x473 &  x485 &  x497 &  x503 &  x509 &  x518 &  x524 &  x527 &  x536 &  x542 &  x547 &  x554 &  x563 &  x572 &  x581 &  x587 &  x596 &  x599 &  x608 &  x617 &  x626 &  x632 &  x638 &  x647 &  x650 &  x659 &  x662 &  x680 &  x686 &  x701 &  x710 &  x716 &  x728 &  x740 &  x758 &  x764 &  x767 &  x770 &  x776 &  x779 &  x794 &  x800 &  x803 &  x815 &  x823 &  x824 &  x833 &  x836 &  x854 &  x860 &  x869 &  x872 &  x875 &  x878 &  x908 &  x914 &  x923 &  x926 &  x938 &  x941 &  x947 &  x962 &  x974 &  x998 &  x1001 &  x1028 &  x1049 &  x1061 &  x1070 &  x1076 &  x1094 &  x1106 &  x1112 & ~x394 & ~x432 & ~x537 & ~x558;
assign c5158 =  x2 &  x5 &  x14 &  x17 &  x26 &  x32 &  x35 &  x44 &  x47 &  x53 &  x59 &  x62 &  x68 &  x83 &  x86 &  x101 &  x104 &  x107 &  x110 &  x116 &  x122 &  x125 &  x131 &  x134 &  x140 &  x143 &  x155 &  x158 &  x161 &  x164 &  x173 &  x182 &  x185 &  x191 &  x194 &  x197 &  x200 &  x206 &  x209 &  x212 &  x221 &  x224 &  x233 &  x236 &  x242 &  x245 &  x248 &  x251 &  x260 &  x266 &  x269 &  x272 &  x275 &  x284 &  x293 &  x296 &  x308 &  x314 &  x317 &  x326 &  x329 &  x332 &  x338 &  x341 &  x347 &  x350 &  x353 &  x356 &  x359 &  x365 &  x371 &  x380 &  x383 &  x389 &  x395 &  x398 &  x404 &  x416 &  x425 &  x428 &  x431 &  x434 &  x437 &  x446 &  x449 &  x467 &  x470 &  x476 &  x485 &  x488 &  x491 &  x506 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x539 &  x545 &  x548 &  x551 &  x554 &  x560 &  x563 &  x566 &  x569 &  x571 &  x572 &  x581 &  x584 &  x587 &  x593 &  x611 &  x614 &  x617 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x649 &  x650 &  x653 &  x656 &  x665 &  x671 &  x683 &  x689 &  x695 &  x698 &  x701 &  x707 &  x710 &  x719 &  x722 &  x725 &  x727 &  x731 &  x734 &  x740 &  x752 &  x761 &  x769 &  x770 &  x773 &  x776 &  x779 &  x791 &  x794 &  x809 &  x815 &  x821 &  x824 &  x833 &  x839 &  x842 &  x845 &  x848 &  x854 &  x860 &  x872 &  x881 &  x887 &  x896 &  x905 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x947 &  x950 &  x956 &  x959 &  x962 &  x971 &  x980 &  x983 &  x986 &  x989 &  x995 &  x998 &  x1004 &  x1007 &  x1013 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1088 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1115 &  x1121 & ~x120 & ~x213 & ~x214 & ~x253 & ~x292 & ~x331 & ~x408 & ~x558;
assign c5160 =  x2 &  x5 &  x11 &  x20 &  x29 &  x50 &  x56 &  x58 &  x62 &  x80 &  x86 &  x116 &  x125 &  x146 &  x149 &  x158 &  x161 &  x167 &  x176 &  x179 &  x182 &  x191 &  x194 &  x200 &  x203 &  x206 &  x212 &  x214 &  x221 &  x236 &  x239 &  x248 &  x254 &  x257 &  x269 &  x272 &  x275 &  x278 &  x299 &  x314 &  x317 &  x335 &  x344 &  x362 &  x368 &  x371 &  x380 &  x386 &  x392 &  x401 &  x410 &  x418 &  x419 &  x425 &  x428 &  x437 &  x446 &  x464 &  x473 &  x485 &  x497 &  x506 &  x514 &  x515 &  x524 &  x536 &  x542 &  x545 &  x547 &  x557 &  x560 &  x563 &  x575 &  x584 &  x587 &  x590 &  x605 &  x611 &  x614 &  x620 &  x623 &  x659 &  x662 &  x671 &  x683 &  x701 &  x704 &  x713 &  x722 &  x725 &  x728 &  x734 &  x755 &  x758 &  x761 &  x767 &  x773 &  x779 &  x788 &  x818 &  x830 &  x839 &  x860 &  x862 &  x863 &  x872 &  x881 &  x908 &  x914 &  x923 &  x953 &  x959 &  x965 &  x967 &  x971 &  x974 &  x980 &  x989 &  x995 &  x1010 &  x1052 &  x1061 &  x1088 &  x1091 &  x1097 &  x1103 &  x1112 &  x1124 & ~x597;
assign c5162 =  x2 &  x8 &  x11 &  x14 &  x29 &  x32 &  x35 &  x47 &  x50 &  x59 &  x65 &  x71 &  x83 &  x95 &  x98 &  x101 &  x104 &  x107 &  x119 &  x122 &  x125 &  x128 &  x137 &  x140 &  x158 &  x188 &  x194 &  x200 &  x203 &  x212 &  x221 &  x239 &  x242 &  x245 &  x269 &  x275 &  x284 &  x293 &  x299 &  x302 &  x305 &  x308 &  x314 &  x320 &  x329 &  x332 &  x338 &  x344 &  x347 &  x350 &  x374 &  x380 &  x395 &  x401 &  x410 &  x413 &  x440 &  x443 &  x452 &  x455 &  x458 &  x461 &  x470 &  x473 &  x482 &  x488 &  x491 &  x509 &  x512 &  x539 &  x547 &  x551 &  x566 &  x569 &  x575 &  x587 &  x599 &  x605 &  x620 &  x629 &  x641 &  x647 &  x650 &  x653 &  x656 &  x659 &  x671 &  x674 &  x692 &  x701 &  x704 &  x707 &  x728 &  x743 &  x746 &  x761 &  x764 &  x767 &  x785 &  x794 &  x818 &  x822 &  x833 &  x842 &  x857 &  x872 &  x878 &  x881 &  x884 &  x887 &  x893 &  x899 &  x908 &  x911 &  x920 &  x947 &  x953 &  x986 &  x989 &  x992 &  x995 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1028 &  x1034 &  x1043 &  x1046 &  x1061 &  x1064 &  x1073 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1121 & ~x432 & ~x472 & ~x511 & ~x693 & ~x756 & ~x795 & ~x834 & ~x873;
assign c5164 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x26 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x68 &  x71 &  x74 &  x80 &  x83 &  x86 &  x89 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x125 &  x128 &  x134 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x161 &  x164 &  x167 &  x170 &  x173 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x209 &  x212 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x323 &  x326 &  x329 &  x332 &  x335 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x380 &  x383 &  x386 &  x389 &  x392 &  x404 &  x407 &  x410 &  x413 &  x422 &  x428 &  x434 &  x437 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x542 &  x545 &  x548 &  x550 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x589 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x626 &  x629 &  x632 &  x635 &  x641 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x668 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x700 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x752 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x845 &  x848 &  x851 &  x857 &  x860 &  x863 &  x866 &  x872 &  x875 &  x878 &  x881 &  x884 &  x893 &  x895 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x928 &  x929 &  x932 &  x934 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x955 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1072 &  x1073 &  x1076 &  x1078 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x141 & ~x180 & ~x219 & ~x600 & ~x639 & ~x678 & ~x819 & ~x1041 & ~x1080;
assign c5166 =  x2 &  x8 &  x11 &  x14 &  x32 &  x38 &  x44 &  x50 &  x53 &  x56 &  x59 &  x62 &  x74 &  x77 &  x83 &  x92 &  x98 &  x101 &  x104 &  x107 &  x119 &  x122 &  x134 &  x137 &  x146 &  x152 &  x155 &  x158 &  x176 &  x182 &  x190 &  x203 &  x212 &  x218 &  x221 &  x227 &  x248 &  x254 &  x257 &  x269 &  x278 &  x287 &  x293 &  x311 &  x314 &  x329 &  x335 &  x338 &  x341 &  x350 &  x356 &  x359 &  x362 &  x365 &  x379 &  x380 &  x392 &  x404 &  x413 &  x418 &  x422 &  x425 &  x428 &  x440 &  x443 &  x446 &  x455 &  x464 &  x467 &  x473 &  x479 &  x485 &  x490 &  x500 &  x506 &  x512 &  x515 &  x518 &  x524 &  x527 &  x530 &  x542 &  x548 &  x554 &  x557 &  x563 &  x566 &  x568 &  x572 &  x599 &  x602 &  x605 &  x608 &  x611 &  x617 &  x632 &  x635 &  x641 &  x647 &  x650 &  x671 &  x680 &  x683 &  x707 &  x710 &  x716 &  x719 &  x731 &  x737 &  x740 &  x752 &  x755 &  x758 &  x767 &  x770 &  x785 &  x788 &  x791 &  x797 &  x806 &  x815 &  x820 &  x821 &  x827 &  x836 &  x842 &  x845 &  x848 &  x854 &  x857 &  x860 &  x869 &  x875 &  x881 &  x896 &  x917 &  x926 &  x935 &  x940 &  x944 &  x950 &  x953 &  x965 &  x968 &  x971 &  x974 &  x980 &  x986 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1106 &  x1109 &  x1118 &  x1121 &  x1130 & ~x363 & ~x480 & ~x519 & ~x525 & ~x597 & ~x603 & ~x714 & ~x720 & ~x792 & ~x831 & ~x837;
assign c5168 =  x2 &  x5 &  x11 &  x14 &  x20 &  x44 &  x47 &  x56 &  x61 &  x62 &  x68 &  x74 &  x89 &  x92 &  x95 &  x98 &  x100 &  x107 &  x119 &  x134 &  x149 &  x152 &  x179 &  x182 &  x188 &  x191 &  x197 &  x203 &  x206 &  x218 &  x224 &  x227 &  x230 &  x236 &  x242 &  x245 &  x248 &  x254 &  x263 &  x269 &  x272 &  x284 &  x299 &  x302 &  x305 &  x319 &  x326 &  x335 &  x344 &  x347 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x389 &  x392 &  x407 &  x413 &  x428 &  x437 &  x440 &  x449 &  x452 &  x461 &  x464 &  x476 &  x485 &  x488 &  x491 &  x500 &  x503 &  x508 &  x509 &  x515 &  x518 &  x533 &  x536 &  x539 &  x551 &  x560 &  x569 &  x572 &  x599 &  x605 &  x611 &  x617 &  x620 &  x623 &  x626 &  x635 &  x638 &  x653 &  x677 &  x683 &  x686 &  x698 &  x707 &  x713 &  x716 &  x722 &  x725 &  x731 &  x737 &  x745 &  x746 &  x749 &  x758 &  x773 &  x784 &  x791 &  x797 &  x800 &  x803 &  x818 &  x821 &  x827 &  x833 &  x842 &  x854 &  x863 &  x869 &  x881 &  x884 &  x899 &  x902 &  x926 &  x929 &  x932 &  x935 &  x941 &  x944 &  x947 &  x965 &  x977 &  x986 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1022 &  x1028 &  x1034 &  x1055 &  x1064 &  x1070 &  x1073 &  x1088 &  x1094 &  x1103 &  x1115 &  x1121 &  x1127 &  x1130 & ~x402 & ~x519 & ~x597 & ~x598 & ~x636;
assign c5170 =  x5 &  x11 &  x20 &  x26 &  x35 &  x41 &  x65 &  x68 &  x83 &  x89 &  x119 &  x122 &  x161 &  x179 &  x212 &  x230 &  x245 &  x260 &  x281 &  x302 &  x320 &  x326 &  x344 &  x347 &  x371 &  x377 &  x398 &  x419 &  x422 &  x428 &  x431 &  x449 &  x458 &  x485 &  x503 &  x506 &  x542 &  x560 &  x566 &  x584 &  x599 &  x608 &  x611 &  x614 &  x620 &  x635 &  x650 &  x698 &  x703 &  x707 &  x743 &  x749 &  x773 &  x782 &  x791 &  x794 &  x812 &  x823 &  x827 &  x845 &  x848 &  x854 &  x857 &  x862 &  x875 &  x878 &  x889 &  x896 &  x902 &  x914 &  x929 &  x940 &  x953 &  x962 &  x965 &  x968 &  x971 &  x989 &  x1001 &  x1055 &  x1064 &  x1073 &  x1115 & ~x324 & ~x363 & ~x480 & ~x756 & ~x796;
assign c5172 =  x29 &  x38 &  x59 &  x65 &  x92 &  x128 &  x140 &  x154 &  x158 &  x167 &  x170 &  x188 &  x191 &  x206 &  x215 &  x239 &  x242 &  x245 &  x254 &  x266 &  x269 &  x302 &  x323 &  x326 &  x350 &  x359 &  x395 &  x401 &  x416 &  x419 &  x440 &  x445 &  x455 &  x458 &  x467 &  x512 &  x515 &  x539 &  x548 &  x554 &  x572 &  x581 &  x593 &  x608 &  x611 &  x617 &  x665 &  x674 &  x683 &  x692 &  x722 &  x725 &  x740 &  x746 &  x749 &  x770 &  x773 &  x776 &  x794 &  x797 &  x809 &  x845 &  x857 &  x860 &  x863 &  x875 &  x899 &  x920 &  x941 &  x956 &  x971 &  x977 &  x980 &  x1007 &  x1025 &  x1046 &  x1073 &  x1079 &  x1097 &  x1100 &  x1115 &  x1124 &  x1130 & ~x237 & ~x432 & ~x433 & ~x519 & ~x558 & ~x597 & ~x598 & ~x675 & ~x909;
assign c5174 =  x2 &  x8 &  x11 &  x17 &  x20 &  x22 &  x23 &  x29 &  x31 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x61 &  x62 &  x65 &  x70 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x458 &  x461 &  x464 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x491 &  x494 &  x497 &  x500 &  x506 &  x509 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x548 &  x551 &  x557 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x605 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x632 &  x635 &  x641 &  x644 &  x647 &  x649 &  x650 &  x653 &  x656 &  x662 &  x671 &  x674 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x701 &  x707 &  x713 &  x722 &  x725 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x758 &  x761 &  x764 &  x767 &  x770 &  x785 &  x788 &  x791 &  x794 &  x800 &  x803 &  x806 &  x812 &  x815 &  x818 &  x824 &  x827 &  x830 &  x833 &  x836 &  x842 &  x845 &  x851 &  x854 &  x857 &  x860 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x923 &  x926 &  x932 &  x935 &  x938 &  x944 &  x947 &  x950 &  x953 &  x959 &  x962 &  x971 &  x977 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x75 & ~x714 & ~x792 & ~x831 & ~x870 & ~x909 & ~x990 & ~x1029;
assign c5176 =  x1 &  x14 &  x26 &  x29 &  x32 &  x39 &  x40 &  x47 &  x56 &  x62 &  x65 &  x71 &  x74 &  x77 &  x78 &  x79 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x107 &  x110 &  x113 &  x117 &  x118 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x149 &  x155 &  x157 &  x161 &  x164 &  x167 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x195 &  x196 &  x197 &  x203 &  x206 &  x221 &  x227 &  x233 &  x236 &  x245 &  x248 &  x260 &  x263 &  x272 &  x274 &  x278 &  x287 &  x290 &  x293 &  x299 &  x311 &  x314 &  x316 &  x320 &  x329 &  x332 &  x335 &  x347 &  x353 &  x355 &  x356 &  x362 &  x365 &  x383 &  x386 &  x392 &  x413 &  x416 &  x422 &  x425 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x458 &  x461 &  x464 &  x467 &  x476 &  x482 &  x485 &  x488 &  x491 &  x497 &  x503 &  x512 &  x536 &  x539 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x572 &  x578 &  x581 &  x584 &  x587 &  x599 &  x605 &  x608 &  x614 &  x620 &  x632 &  x635 &  x647 &  x650 &  x653 &  x659 &  x665 &  x674 &  x680 &  x689 &  x698 &  x701 &  x707 &  x710 &  x716 &  x722 &  x725 &  x737 &  x740 &  x743 &  x746 &  x752 &  x755 &  x758 &  x764 &  x776 &  x782 &  x785 &  x791 &  x800 &  x803 &  x809 &  x815 &  x824 &  x833 &  x839 &  x842 &  x848 &  x851 &  x854 &  x866 &  x872 &  x878 &  x890 &  x893 &  x896 &  x899 &  x905 &  x908 &  x914 &  x917 &  x923 &  x929 &  x938 &  x941 &  x947 &  x950 &  x956 &  x959 &  x968 &  x971 &  x974 &  x977 &  x983 &  x986 &  x989 &  x998 &  x1001 &  x1004 &  x1013 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1046 &  x1049 &  x1055 &  x1058 &  x1061 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1118 &  x1124 &  x1127 & ~x3 & ~x42 & ~x43 & ~x81 & ~x90 & ~x91 & ~x168 & ~x246 & ~x252 & ~x585 & ~x624;
assign c5178 =  x8 &  x20 &  x26 &  x29 &  x38 &  x83 &  x92 &  x95 &  x122 &  x137 &  x146 &  x173 &  x206 &  x233 &  x242 &  x290 &  x308 &  x317 &  x335 &  x341 &  x344 &  x425 &  x428 &  x437 &  x449 &  x461 &  x464 &  x475 &  x506 &  x551 &  x553 &  x554 &  x560 &  x563 &  x575 &  x581 &  x586 &  x611 &  x625 &  x638 &  x665 &  x677 &  x702 &  x703 &  x707 &  x710 &  x731 &  x752 &  x767 &  x770 &  x781 &  x785 &  x854 &  x862 &  x875 &  x899 &  x901 &  x902 &  x914 &  x980 &  x986 &  x998 &  x1007 &  x1019 &  x1040 &  x1043 &  x1046 &  x1067 &  x1070 &  x1082 &  x1088 &  x1100 &  x1103 &  x1109 &  x1115 &  x1118 &  x1124 & ~x472 & ~x693 & ~x756 & ~x834 & ~x873;
assign c5180 =  x5 &  x17 &  x20 &  x29 &  x44 &  x53 &  x83 &  x86 &  x98 &  x104 &  x167 &  x173 &  x179 &  x248 &  x269 &  x278 &  x314 &  x320 &  x347 &  x359 &  x389 &  x392 &  x407 &  x419 &  x422 &  x443 &  x461 &  x476 &  x482 &  x491 &  x503 &  x527 &  x533 &  x545 &  x581 &  x635 &  x638 &  x644 &  x668 &  x683 &  x698 &  x707 &  x710 &  x737 &  x752 &  x767 &  x779 &  x803 &  x809 &  x824 &  x842 &  x851 &  x860 &  x878 &  x881 &  x893 &  x953 &  x956 &  x983 &  x989 &  x1004 &  x1007 &  x1052 &  x1056 &  x1064 &  x1085 &  x1088 &  x1091 &  x1094 &  x1096 &  x1103 & ~x312 & ~x429 & ~x628 & ~x667 & ~x816 & ~x870 & ~x987 & ~x1066;
assign c5182 =  x5 &  x17 &  x35 &  x41 &  x47 &  x62 &  x74 &  x77 &  x80 &  x83 &  x89 &  x107 &  x113 &  x131 &  x134 &  x167 &  x170 &  x176 &  x194 &  x197 &  x200 &  x218 &  x242 &  x251 &  x254 &  x281 &  x284 &  x305 &  x308 &  x338 &  x341 &  x353 &  x356 &  x359 &  x362 &  x374 &  x377 &  x380 &  x383 &  x386 &  x395 &  x398 &  x401 &  x422 &  x449 &  x458 &  x464 &  x469 &  x491 &  x497 &  x506 &  x512 &  x515 &  x521 &  x530 &  x584 &  x590 &  x593 &  x599 &  x605 &  x608 &  x620 &  x623 &  x635 &  x644 &  x665 &  x667 &  x698 &  x701 &  x706 &  x710 &  x728 &  x737 &  x746 &  x749 &  x758 &  x761 &  x767 &  x779 &  x785 &  x794 &  x806 &  x809 &  x824 &  x827 &  x839 &  x851 &  x854 &  x863 &  x887 &  x905 &  x923 &  x935 &  x980 &  x1007 &  x1025 &  x1028 &  x1040 &  x1055 &  x1058 &  x1064 &  x1067 &  x1073 &  x1091 &  x1094 &  x1109 &  x1112 &  x1115 & ~x237 & ~x276 & ~x277 & ~x285 & ~x316 & ~x324 & ~x519 & ~x678;
assign c5184 =  x11 &  x14 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x65 &  x68 &  x89 &  x95 &  x98 &  x104 &  x113 &  x116 &  x119 &  x122 &  x128 &  x140 &  x182 &  x185 &  x197 &  x203 &  x206 &  x209 &  x218 &  x221 &  x230 &  x242 &  x245 &  x254 &  x257 &  x260 &  x263 &  x266 &  x272 &  x275 &  x281 &  x290 &  x299 &  x311 &  x326 &  x344 &  x347 &  x350 &  x353 &  x362 &  x365 &  x374 &  x383 &  x386 &  x422 &  x425 &  x467 &  x475 &  x488 &  x497 &  x512 &  x514 &  x524 &  x527 &  x533 &  x536 &  x551 &  x557 &  x566 &  x578 &  x593 &  x596 &  x599 &  x611 &  x626 &  x638 &  x641 &  x647 &  x677 &  x689 &  x701 &  x704 &  x713 &  x716 &  x722 &  x725 &  x749 &  x767 &  x773 &  x776 &  x788 &  x794 &  x803 &  x818 &  x836 &  x848 &  x854 &  x860 &  x872 &  x884 &  x887 &  x890 &  x893 &  x898 &  x899 &  x914 &  x926 &  x941 &  x950 &  x956 &  x959 &  x962 &  x968 &  x983 &  x995 &  x998 &  x1004 &  x1031 &  x1037 &  x1046 &  x1055 &  x1058 &  x1073 &  x1076 &  x1088 &  x1109 &  x1121 &  x1124 & ~x72 & ~x195 & ~x273 & ~x628 & ~x987;
assign c5186 =  x8 &  x17 &  x38 &  x47 &  x71 &  x92 &  x104 &  x107 &  x113 &  x116 &  x119 &  x125 &  x149 &  x152 &  x167 &  x179 &  x191 &  x203 &  x209 &  x212 &  x215 &  x218 &  x221 &  x227 &  x245 &  x248 &  x251 &  x266 &  x269 &  x275 &  x284 &  x293 &  x299 &  x305 &  x317 &  x346 &  x362 &  x365 &  x380 &  x407 &  x413 &  x416 &  x425 &  x452 &  x455 &  x464 &  x479 &  x497 &  x503 &  x506 &  x508 &  x509 &  x521 &  x524 &  x533 &  x539 &  x542 &  x548 &  x551 &  x560 &  x569 &  x581 &  x586 &  x599 &  x608 &  x611 &  x623 &  x632 &  x641 &  x644 &  x662 &  x667 &  x668 &  x671 &  x683 &  x704 &  x705 &  x713 &  x716 &  x737 &  x745 &  x755 &  x758 &  x764 &  x770 &  x776 &  x779 &  x785 &  x791 &  x794 &  x806 &  x812 &  x815 &  x821 &  x823 &  x833 &  x863 &  x899 &  x914 &  x917 &  x920 &  x923 &  x938 &  x941 &  x947 &  x959 &  x974 &  x986 &  x989 &  x992 &  x1010 &  x1019 &  x1025 &  x1040 &  x1046 &  x1049 &  x1055 &  x1058 &  x1082 &  x1097 &  x1100 &  x1106 &  x1112 &  x1118 &  x1124 &  x1130 & ~x354 & ~x355;
assign c5188 =  x32 &  x56 &  x65 &  x71 &  x77 &  x80 &  x86 &  x95 &  x104 &  x191 &  x206 &  x221 &  x224 &  x296 &  x299 &  x302 &  x323 &  x332 &  x335 &  x356 &  x362 &  x374 &  x385 &  x395 &  x397 &  x401 &  x458 &  x463 &  x475 &  x515 &  x523 &  x533 &  x545 &  x557 &  x572 &  x602 &  x629 &  x644 &  x650 &  x662 &  x677 &  x728 &  x731 &  x740 &  x749 &  x761 &  x773 &  x782 &  x830 &  x839 &  x848 &  x860 &  x872 &  x920 &  x965 &  x1010 &  x1016 &  x1034 &  x1040 &  x1064 &  x1076 &  x1082 & ~x603 & ~x642 & ~x720 & ~x753 & ~x759 & ~x792 & ~x798 & ~x873 & ~x909;
assign c5190 =  x5 &  x14 &  x20 &  x26 &  x35 &  x38 &  x41 &  x50 &  x53 &  x56 &  x62 &  x79 &  x80 &  x95 &  x98 &  x101 &  x113 &  x118 &  x119 &  x125 &  x128 &  x131 &  x134 &  x143 &  x146 &  x152 &  x155 &  x161 &  x164 &  x173 &  x179 &  x188 &  x191 &  x197 &  x200 &  x209 &  x212 &  x218 &  x221 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x263 &  x266 &  x269 &  x274 &  x275 &  x284 &  x290 &  x302 &  x308 &  x314 &  x317 &  x326 &  x335 &  x338 &  x344 &  x355 &  x356 &  x365 &  x371 &  x377 &  x386 &  x395 &  x410 &  x422 &  x434 &  x437 &  x440 &  x446 &  x449 &  x464 &  x467 &  x470 &  x500 &  x503 &  x506 &  x509 &  x512 &  x518 &  x521 &  x532 &  x551 &  x554 &  x557 &  x560 &  x572 &  x575 &  x587 &  x590 &  x593 &  x596 &  x602 &  x605 &  x617 &  x620 &  x626 &  x629 &  x647 &  x653 &  x665 &  x671 &  x686 &  x695 &  x713 &  x716 &  x722 &  x737 &  x746 &  x749 &  x764 &  x773 &  x776 &  x782 &  x791 &  x797 &  x800 &  x803 &  x806 &  x815 &  x821 &  x824 &  x833 &  x838 &  x848 &  x851 &  x863 &  x866 &  x872 &  x875 &  x877 &  x878 &  x881 &  x884 &  x890 &  x902 &  x908 &  x914 &  x916 &  x920 &  x926 &  x932 &  x941 &  x950 &  x959 &  x962 &  x965 &  x971 &  x995 &  x1001 &  x1004 &  x1010 &  x1022 &  x1031 &  x1034 &  x1037 &  x1055 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1085 &  x1106 &  x1118 &  x1127 &  x1130 & ~x81 & ~x246 & ~x327 & ~x366 & ~x405 & ~x507 & ~x546 & ~x633 & ~x672 & ~x711 & ~x828;
assign c5192 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x41 &  x44 &  x47 &  x50 &  x56 &  x59 &  x65 &  x71 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x197 &  x203 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x383 &  x389 &  x392 &  x395 &  x398 &  x404 &  x407 &  x410 &  x413 &  x419 &  x422 &  x425 &  x428 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x476 &  x479 &  x482 &  x485 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x524 &  x527 &  x530 &  x533 &  x536 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x575 &  x578 &  x581 &  x587 &  x590 &  x596 &  x599 &  x602 &  x605 &  x608 &  x614 &  x617 &  x620 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x647 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x731 &  x734 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x770 &  x776 &  x779 &  x782 &  x788 &  x791 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x830 &  x833 &  x836 &  x838 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x881 &  x884 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x916 &  x923 &  x926 &  x929 &  x932 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1067 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130 & ~x42 & ~x81 & ~x168 & ~x169 & ~x207 & ~x246 & ~x247 & ~x285 & ~x324 & ~x363 & ~x402 & ~x441 & ~x480 & ~x519 & ~x558 & ~x597 & ~x828 & ~x867;
assign c5194 =  x11 &  x23 &  x47 &  x53 &  x59 &  x80 &  x83 &  x92 &  x98 &  x101 &  x113 &  x125 &  x128 &  x131 &  x137 &  x149 &  x152 &  x197 &  x206 &  x212 &  x215 &  x224 &  x236 &  x245 &  x272 &  x305 &  x308 &  x350 &  x383 &  x392 &  x404 &  x419 &  x440 &  x458 &  x482 &  x500 &  x515 &  x518 &  x524 &  x533 &  x542 &  x551 &  x557 &  x563 &  x580 &  x584 &  x590 &  x605 &  x629 &  x635 &  x644 &  x650 &  x671 &  x674 &  x677 &  x680 &  x689 &  x698 &  x701 &  x707 &  x710 &  x716 &  x749 &  x770 &  x779 &  x781 &  x782 &  x818 &  x820 &  x857 &  x866 &  x872 &  x878 &  x899 &  x902 &  x914 &  x917 &  x923 &  x929 &  x932 &  x935 &  x941 &  x944 &  x974 &  x980 &  x986 &  x992 &  x1022 &  x1025 &  x1054 &  x1091 &  x1096 &  x1106 &  x1121 & ~x273 & ~x312 & ~x429 & ~x666 & ~x667 & ~x948 & ~x1026;
assign c5196 =  x56 &  x71 &  x74 &  x89 &  x110 &  x113 &  x116 &  x124 &  x128 &  x131 &  x146 &  x191 &  x200 &  x206 &  x218 &  x221 &  x230 &  x242 &  x248 &  x272 &  x275 &  x344 &  x362 &  x377 &  x398 &  x407 &  x428 &  x440 &  x446 &  x449 &  x467 &  x476 &  x482 &  x500 &  x503 &  x506 &  x524 &  x533 &  x572 &  x653 &  x692 &  x719 &  x725 &  x743 &  x782 &  x803 &  x809 &  x833 &  x845 &  x866 &  x872 &  x884 &  x914 &  x923 &  x929 &  x944 &  x983 &  x1010 &  x1043 &  x1052 &  x1067 &  x1097 &  x1106 &  x1121 &  x1127 & ~x408 & ~x433;
assign c5198 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x44 &  x53 &  x59 &  x62 &  x68 &  x77 &  x83 &  x89 &  x92 &  x107 &  x119 &  x122 &  x125 &  x128 &  x140 &  x143 &  x146 &  x164 &  x167 &  x191 &  x194 &  x200 &  x206 &  x212 &  x218 &  x227 &  x230 &  x233 &  x236 &  x263 &  x266 &  x281 &  x302 &  x308 &  x311 &  x323 &  x335 &  x347 &  x350 &  x353 &  x356 &  x362 &  x368 &  x371 &  x374 &  x377 &  x380 &  x389 &  x401 &  x407 &  x416 &  x419 &  x422 &  x431 &  x437 &  x443 &  x452 &  x455 &  x458 &  x461 &  x467 &  x470 &  x473 &  x476 &  x485 &  x488 &  x494 &  x500 &  x506 &  x515 &  x521 &  x539 &  x542 &  x551 &  x563 &  x581 &  x584 &  x590 &  x593 &  x599 &  x602 &  x605 &  x608 &  x611 &  x617 &  x620 &  x623 &  x626 &  x632 &  x644 &  x647 &  x650 &  x659 &  x662 &  x677 &  x692 &  x695 &  x701 &  x704 &  x707 &  x713 &  x719 &  x731 &  x737 &  x740 &  x745 &  x752 &  x755 &  x770 &  x773 &  x776 &  x784 &  x791 &  x794 &  x800 &  x812 &  x815 &  x821 &  x823 &  x824 &  x842 &  x851 &  x854 &  x857 &  x860 &  x862 &  x866 &  x875 &  x878 &  x881 &  x890 &  x895 &  x899 &  x901 &  x902 &  x905 &  x920 &  x926 &  x929 &  x932 &  x941 &  x944 &  x947 &  x950 &  x959 &  x965 &  x968 &  x977 &  x983 &  x1001 &  x1004 &  x1010 &  x1016 &  x1022 &  x1034 &  x1037 &  x1040 &  x1055 &  x1058 &  x1070 &  x1076 &  x1091 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130 & ~x315 & ~x354 & ~x537 & ~x756 & ~x1074 & ~x1086;
assign c5200 =  x5 &  x8 &  x11 &  x14 &  x17 &  x26 &  x29 &  x32 &  x35 &  x44 &  x47 &  x50 &  x56 &  x65 &  x68 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x110 &  x116 &  x122 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x155 &  x158 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x188 &  x191 &  x194 &  x200 &  x203 &  x212 &  x215 &  x218 &  x224 &  x233 &  x236 &  x239 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x278 &  x281 &  x284 &  x290 &  x293 &  x305 &  x308 &  x317 &  x323 &  x326 &  x332 &  x335 &  x344 &  x347 &  x350 &  x356 &  x359 &  x362 &  x368 &  x371 &  x374 &  x380 &  x383 &  x389 &  x392 &  x395 &  x398 &  x404 &  x407 &  x410 &  x413 &  x419 &  x422 &  x428 &  x434 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x464 &  x476 &  x482 &  x488 &  x494 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x527 &  x536 &  x539 &  x542 &  x545 &  x551 &  x557 &  x569 &  x572 &  x575 &  x590 &  x593 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x656 &  x662 &  x668 &  x674 &  x677 &  x683 &  x689 &  x692 &  x695 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x731 &  x737 &  x746 &  x758 &  x761 &  x767 &  x773 &  x776 &  x779 &  x788 &  x791 &  x797 &  x800 &  x809 &  x812 &  x821 &  x824 &  x827 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x857 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x884 &  x887 &  x893 &  x896 &  x899 &  x911 &  x914 &  x920 &  x926 &  x932 &  x935 &  x944 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1064 &  x1067 &  x1076 &  x1079 &  x1082 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x120 & ~x159 & ~x237 & ~x238 & ~x276 & ~x315 & ~x324 & ~x354 & ~x363 & ~x369 & ~x447 & ~x526 & ~x564;
assign c5202 =  x2 &  x5 &  x11 &  x17 &  x20 &  x26 &  x32 &  x35 &  x41 &  x47 &  x50 &  x56 &  x59 &  x62 &  x65 &  x68 &  x77 &  x80 &  x92 &  x95 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x128 &  x134 &  x146 &  x152 &  x155 &  x161 &  x167 &  x170 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x218 &  x221 &  x227 &  x230 &  x235 &  x242 &  x245 &  x260 &  x263 &  x266 &  x272 &  x274 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x313 &  x314 &  x317 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x344 &  x353 &  x356 &  x359 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x410 &  x413 &  x425 &  x430 &  x431 &  x434 &  x440 &  x443 &  x446 &  x449 &  x461 &  x467 &  x469 &  x470 &  x476 &  x482 &  x494 &  x500 &  x506 &  x508 &  x509 &  x518 &  x521 &  x527 &  x545 &  x547 &  x548 &  x551 &  x554 &  x557 &  x569 &  x575 &  x581 &  x587 &  x596 &  x602 &  x605 &  x608 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x638 &  x650 &  x656 &  x662 &  x665 &  x668 &  x677 &  x680 &  x686 &  x692 &  x695 &  x698 &  x704 &  x707 &  x713 &  x716 &  x722 &  x728 &  x731 &  x737 &  x740 &  x746 &  x755 &  x758 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x784 &  x788 &  x791 &  x800 &  x803 &  x809 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x851 &  x854 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x884 &  x887 &  x902 &  x905 &  x908 &  x914 &  x917 &  x920 &  x923 &  x929 &  x935 &  x938 &  x944 &  x950 &  x953 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x989 &  x992 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1037 &  x1046 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1084 &  x1088 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 & ~x198 & ~x237 & ~x276 & ~x277 & ~x558;
assign c5204 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x35 &  x38 &  x41 &  x50 &  x53 &  x56 &  x59 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x128 &  x137 &  x140 &  x143 &  x146 &  x149 &  x155 &  x158 &  x167 &  x170 &  x176 &  x197 &  x200 &  x203 &  x206 &  x212 &  x215 &  x218 &  x221 &  x227 &  x230 &  x233 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x263 &  x269 &  x272 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x302 &  x305 &  x311 &  x314 &  x320 &  x323 &  x326 &  x329 &  x335 &  x338 &  x341 &  x350 &  x353 &  x356 &  x362 &  x365 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x443 &  x446 &  x458 &  x461 &  x467 &  x470 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x509 &  x512 &  x518 &  x521 &  x524 &  x533 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x560 &  x566 &  x572 &  x578 &  x581 &  x584 &  x587 &  x590 &  x596 &  x599 &  x605 &  x608 &  x611 &  x614 &  x623 &  x629 &  x632 &  x635 &  x641 &  x650 &  x653 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x686 &  x695 &  x698 &  x704 &  x707 &  x710 &  x713 &  x716 &  x722 &  x725 &  x731 &  x734 &  x737 &  x740 &  x743 &  x749 &  x758 &  x761 &  x764 &  x776 &  x788 &  x791 &  x794 &  x797 &  x800 &  x806 &  x809 &  x815 &  x818 &  x821 &  x824 &  x827 &  x833 &  x836 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x872 &  x878 &  x881 &  x884 &  x887 &  x896 &  x899 &  x902 &  x911 &  x914 &  x920 &  x923 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x950 &  x956 &  x959 &  x962 &  x968 &  x971 &  x974 &  x977 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1028 &  x1034 &  x1037 &  x1043 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1073 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 & ~x3 & ~x4 & ~x12 & ~x42 & ~x43 & ~x51 & ~x63 & ~x90 & ~x108 & ~x129 & ~x168 & ~x207 & ~x246 & ~x285 & ~x324 & ~x639 & ~x678 & ~x717 & ~x819 & ~x846 & ~x858 & ~x885 & ~x897 & ~x924 & ~x936 & ~x1047 & ~x1086;
assign c5206 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x44 &  x47 &  x50 &  x53 &  x56 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x89 &  x92 &  x95 &  x98 &  x101 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x164 &  x167 &  x170 &  x176 &  x197 &  x206 &  x215 &  x218 &  x221 &  x224 &  x230 &  x233 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x278 &  x284 &  x296 &  x302 &  x308 &  x311 &  x314 &  x320 &  x329 &  x332 &  x335 &  x341 &  x347 &  x356 &  x359 &  x362 &  x365 &  x371 &  x377 &  x380 &  x401 &  x404 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x479 &  x482 &  x485 &  x488 &  x497 &  x509 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x584 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x623 &  x626 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x659 &  x668 &  x671 &  x674 &  x680 &  x683 &  x686 &  x688 &  x692 &  x695 &  x698 &  x707 &  x710 &  x716 &  x719 &  x722 &  x725 &  x728 &  x734 &  x740 &  x743 &  x758 &  x764 &  x770 &  x773 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x803 &  x806 &  x809 &  x812 &  x818 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x845 &  x848 &  x854 &  x857 &  x863 &  x866 &  x869 &  x872 &  x875 &  x884 &  x890 &  x896 &  x905 &  x911 &  x920 &  x926 &  x947 &  x950 &  x953 &  x956 &  x959 &  x961 &  x962 &  x971 &  x977 &  x980 &  x986 &  x989 &  x992 &  x998 &  x1004 &  x1007 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1049 &  x1064 &  x1067 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1121 &  x1127 & ~x42 & ~x81 & ~x120 & ~x121 & ~x207 & ~x246 & ~x285 & ~x324 & ~x402 & ~x423 & ~x483;
assign c5208 =  x5 &  x20 &  x41 &  x59 &  x74 &  x77 &  x80 &  x98 &  x107 &  x113 &  x116 &  x122 &  x128 &  x131 &  x140 &  x143 &  x152 &  x155 &  x161 &  x167 &  x176 &  x179 &  x182 &  x200 &  x209 &  x212 &  x215 &  x218 &  x221 &  x233 &  x242 &  x272 &  x284 &  x287 &  x293 &  x305 &  x323 &  x331 &  x335 &  x347 &  x362 &  x371 &  x383 &  x395 &  x401 &  x409 &  x416 &  x431 &  x458 &  x464 &  x479 &  x485 &  x488 &  x503 &  x509 &  x512 &  x524 &  x527 &  x536 &  x545 &  x548 &  x557 &  x566 &  x574 &  x578 &  x587 &  x590 &  x599 &  x629 &  x635 &  x638 &  x641 &  x646 &  x647 &  x656 &  x665 &  x701 &  x707 &  x713 &  x722 &  x767 &  x776 &  x782 &  x785 &  x818 &  x827 &  x830 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x893 &  x908 &  x920 &  x926 &  x944 &  x950 &  x962 &  x965 &  x968 &  x979 &  x980 &  x1013 &  x1016 &  x1025 &  x1028 &  x1031 &  x1034 &  x1058 &  x1096 &  x1100 &  x1124 & ~x354 & ~x393 & ~x570 & ~x648;
assign c5210 =  x2 &  x5 &  x14 &  x23 &  x35 &  x44 &  x59 &  x65 &  x68 &  x73 &  x74 &  x77 &  x79 &  x92 &  x98 &  x101 &  x104 &  x113 &  x118 &  x119 &  x125 &  x143 &  x146 &  x151 &  x155 &  x158 &  x167 &  x172 &  x173 &  x184 &  x191 &  x200 &  x206 &  x209 &  x212 &  x215 &  x227 &  x230 &  x233 &  x239 &  x242 &  x245 &  x248 &  x260 &  x263 &  x266 &  x272 &  x275 &  x281 &  x287 &  x290 &  x299 &  x308 &  x323 &  x326 &  x332 &  x335 &  x344 &  x347 &  x359 &  x362 &  x365 &  x371 &  x377 &  x389 &  x392 &  x395 &  x398 &  x404 &  x422 &  x431 &  x434 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x464 &  x467 &  x473 &  x479 &  x494 &  x497 &  x500 &  x503 &  x506 &  x518 &  x521 &  x530 &  x539 &  x563 &  x566 &  x572 &  x575 &  x577 &  x578 &  x581 &  x584 &  x590 &  x596 &  x599 &  x605 &  x608 &  x614 &  x617 &  x638 &  x647 &  x656 &  x662 &  x665 &  x668 &  x680 &  x686 &  x689 &  x701 &  x704 &  x707 &  x722 &  x734 &  x740 &  x752 &  x755 &  x758 &  x763 &  x767 &  x782 &  x791 &  x803 &  x806 &  x808 &  x809 &  x815 &  x818 &  x821 &  x830 &  x833 &  x836 &  x857 &  x860 &  x863 &  x869 &  x878 &  x881 &  x899 &  x905 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x944 &  x947 &  x950 &  x962 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x992 &  x998 &  x1007 &  x1016 &  x1022 &  x1025 &  x1034 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1061 &  x1070 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1100 &  x1106 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x441 & ~x480 & ~x558 & ~x597 & ~x714;
assign c5212 =  x2 &  x14 &  x53 &  x62 &  x65 &  x71 &  x77 &  x92 &  x134 &  x137 &  x143 &  x149 &  x158 &  x170 &  x185 &  x188 &  x215 &  x218 &  x221 &  x227 &  x236 &  x239 &  x242 &  x245 &  x251 &  x275 &  x284 &  x287 &  x296 &  x302 &  x323 &  x359 &  x368 &  x374 &  x395 &  x422 &  x436 &  x443 &  x449 &  x476 &  x479 &  x491 &  x503 &  x518 &  x536 &  x575 &  x584 &  x599 &  x614 &  x629 &  x647 &  x653 &  x662 &  x668 &  x677 &  x680 &  x683 &  x740 &  x749 &  x761 &  x767 &  x773 &  x776 &  x791 &  x794 &  x803 &  x821 &  x830 &  x836 &  x842 &  x845 &  x860 &  x866 &  x872 &  x892 &  x901 &  x926 &  x932 &  x940 &  x950 &  x956 &  x959 &  x968 &  x974 &  x995 &  x1016 &  x1031 &  x1043 &  x1064 &  x1067 &  x1103 &  x1112 &  x1118 &  x1121 &  x1124 & ~x315 & ~x354 & ~x393 & ~x432 & ~x471 & ~x597 & ~x615 & ~x873 & ~x909;
assign c5214 =  x8 &  x11 &  x14 &  x20 &  x23 &  x29 &  x35 &  x41 &  x44 &  x53 &  x59 &  x65 &  x74 &  x83 &  x86 &  x89 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x122 &  x128 &  x131 &  x137 &  x149 &  x152 &  x155 &  x161 &  x164 &  x170 &  x173 &  x176 &  x179 &  x191 &  x194 &  x197 &  x206 &  x215 &  x218 &  x221 &  x227 &  x242 &  x251 &  x254 &  x260 &  x263 &  x278 &  x281 &  x290 &  x293 &  x296 &  x299 &  x302 &  x308 &  x311 &  x317 &  x322 &  x332 &  x335 &  x338 &  x341 &  x344 &  x353 &  x356 &  x359 &  x361 &  x362 &  x371 &  x374 &  x380 &  x383 &  x392 &  x395 &  x398 &  x401 &  x407 &  x413 &  x416 &  x419 &  x425 &  x431 &  x437 &  x446 &  x452 &  x458 &  x461 &  x464 &  x473 &  x476 &  x479 &  x482 &  x491 &  x494 &  x497 &  x500 &  x503 &  x512 &  x518 &  x521 &  x524 &  x527 &  x533 &  x539 &  x542 &  x545 &  x551 &  x554 &  x557 &  x566 &  x569 &  x575 &  x578 &  x584 &  x587 &  x590 &  x608 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x638 &  x647 &  x650 &  x653 &  x656 &  x659 &  x668 &  x671 &  x677 &  x683 &  x686 &  x692 &  x695 &  x698 &  x704 &  x710 &  x716 &  x722 &  x725 &  x731 &  x743 &  x749 &  x752 &  x755 &  x761 &  x764 &  x767 &  x773 &  x782 &  x785 &  x788 &  x791 &  x797 &  x800 &  x806 &  x809 &  x812 &  x815 &  x821 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x845 &  x848 &  x854 &  x857 &  x872 &  x875 &  x878 &  x881 &  x884 &  x890 &  x893 &  x896 &  x902 &  x905 &  x908 &  x911 &  x920 &  x926 &  x929 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x956 &  x962 &  x968 &  x971 &  x974 &  x977 &  x980 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1064 &  x1079 &  x1082 &  x1088 &  x1091 &  x1097 &  x1106 &  x1109 &  x1112 &  x1124 &  x1127 &  x1130 & ~x207 & ~x288 & ~x585 & ~x639 & ~x657 & ~x678 & ~x852 & ~x891 & ~x918 & ~x930 & ~x969 & ~x996 & ~x1008 & ~x1029 & ~x1047 & ~x1068;
assign c5216 =  x2 &  x5 &  x8 &  x11 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x44 &  x50 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x80 &  x83 &  x86 &  x98 &  x107 &  x110 &  x116 &  x118 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x203 &  x206 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x236 &  x239 &  x242 &  x248 &  x257 &  x260 &  x263 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x341 &  x344 &  x347 &  x350 &  x356 &  x359 &  x362 &  x368 &  x371 &  x374 &  x380 &  x383 &  x386 &  x392 &  x395 &  x398 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x434 &  x437 &  x440 &  x443 &  x446 &  x455 &  x458 &  x467 &  x473 &  x476 &  x479 &  x482 &  x488 &  x491 &  x494 &  x500 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x554 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x590 &  x596 &  x599 &  x602 &  x605 &  x608 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x635 &  x638 &  x641 &  x644 &  x647 &  x653 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x683 &  x688 &  x689 &  x692 &  x695 &  x698 &  x704 &  x706 &  x713 &  x716 &  x719 &  x722 &  x731 &  x734 &  x737 &  x740 &  x743 &  x749 &  x752 &  x755 &  x758 &  x761 &  x766 &  x767 &  x770 &  x773 &  x779 &  x782 &  x784 &  x785 &  x788 &  x794 &  x797 &  x800 &  x803 &  x805 &  x812 &  x815 &  x818 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x844 &  x845 &  x851 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x917 &  x920 &  x922 &  x923 &  x926 &  x932 &  x935 &  x941 &  x944 &  x947 &  x950 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1000 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1027 &  x1031 &  x1033 &  x1034 &  x1037 &  x1040 &  x1045 &  x1046 &  x1049 &  x1051 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1072 &  x1073 &  x1076 &  x1085 &  x1094 &  x1099 &  x1100 &  x1103 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x42;
assign c5218 =  x2 &  x5 &  x14 &  x23 &  x38 &  x41 &  x44 &  x50 &  x53 &  x56 &  x58 &  x68 &  x71 &  x77 &  x80 &  x86 &  x97 &  x104 &  x110 &  x113 &  x116 &  x122 &  x128 &  x134 &  x140 &  x143 &  x146 &  x179 &  x182 &  x209 &  x215 &  x227 &  x230 &  x242 &  x245 &  x254 &  x278 &  x287 &  x290 &  x293 &  x296 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x326 &  x335 &  x341 &  x344 &  x356 &  x359 &  x365 &  x371 &  x386 &  x389 &  x392 &  x395 &  x401 &  x407 &  x422 &  x425 &  x437 &  x446 &  x452 &  x458 &  x461 &  x464 &  x467 &  x476 &  x488 &  x491 &  x494 &  x518 &  x521 &  x524 &  x527 &  x536 &  x539 &  x554 &  x560 &  x566 &  x569 &  x575 &  x590 &  x599 &  x614 &  x617 &  x623 &  x626 &  x629 &  x638 &  x641 &  x644 &  x662 &  x665 &  x683 &  x706 &  x707 &  x710 &  x716 &  x719 &  x731 &  x749 &  x755 &  x758 &  x761 &  x764 &  x776 &  x785 &  x791 &  x823 &  x824 &  x839 &  x857 &  x863 &  x866 &  x875 &  x881 &  x887 &  x905 &  x911 &  x917 &  x926 &  x935 &  x950 &  x953 &  x965 &  x974 &  x977 &  x998 &  x1013 &  x1016 &  x1022 &  x1025 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1064 &  x1070 &  x1076 &  x1094 &  x1097 &  x1100 &  x1106 &  x1112 &  x1118 &  x1124 &  x1127 &  x1130 & ~x198 & ~x276 & ~x316 & ~x375 & ~x531;
assign c5220 =  x2 &  x5 &  x14 &  x23 &  x56 &  x83 &  x89 &  x95 &  x113 &  x131 &  x140 &  x158 &  x164 &  x176 &  x179 &  x194 &  x230 &  x236 &  x254 &  x266 &  x269 &  x272 &  x308 &  x320 &  x371 &  x398 &  x407 &  x410 &  x485 &  x497 &  x506 &  x521 &  x536 &  x581 &  x608 &  x614 &  x626 &  x635 &  x653 &  x671 &  x677 &  x689 &  x698 &  x746 &  x761 &  x770 &  x773 &  x782 &  x785 &  x797 &  x806 &  x818 &  x824 &  x845 &  x860 &  x869 &  x875 &  x896 &  x923 &  x935 &  x941 &  x947 &  x953 &  x959 &  x977 &  x1013 &  x1028 &  x1043 &  x1046 &  x1049 &  x1052 &  x1061 &  x1082 &  x1085 &  x1088 &  x1097 &  x1124 &  x1130 & ~x39 & ~x315 & ~x433 & ~x492 & ~x531 & ~x1062 & ~x1101;
assign c5222 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x56 &  x59 &  x68 &  x71 &  x74 &  x77 &  x79 &  x80 &  x83 &  x89 &  x92 &  x98 &  x104 &  x107 &  x110 &  x116 &  x118 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x157 &  x158 &  x161 &  x164 &  x173 &  x176 &  x179 &  x182 &  x185 &  x191 &  x194 &  x195 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x224 &  x230 &  x233 &  x235 &  x236 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x274 &  x275 &  x278 &  x290 &  x293 &  x296 &  x308 &  x311 &  x313 &  x314 &  x317 &  x320 &  x326 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x356 &  x359 &  x365 &  x368 &  x371 &  x377 &  x383 &  x386 &  x389 &  x398 &  x401 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x437 &  x440 &  x443 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x473 &  x476 &  x485 &  x497 &  x500 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x530 &  x533 &  x536 &  x539 &  x545 &  x548 &  x554 &  x566 &  x572 &  x578 &  x581 &  x587 &  x590 &  x596 &  x599 &  x602 &  x608 &  x614 &  x617 &  x620 &  x623 &  x626 &  x632 &  x638 &  x641 &  x644 &  x653 &  x656 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x683 &  x689 &  x692 &  x695 &  x698 &  x701 &  x710 &  x713 &  x716 &  x722 &  x728 &  x734 &  x737 &  x743 &  x749 &  x755 &  x758 &  x764 &  x767 &  x770 &  x773 &  x779 &  x782 &  x785 &  x788 &  x794 &  x800 &  x803 &  x806 &  x812 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x884 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x911 &  x914 &  x920 &  x926 &  x929 &  x935 &  x938 &  x947 &  x950 &  x959 &  x962 &  x965 &  x968 &  x971 &  x977 &  x983 &  x986 &  x989 &  x995 &  x1004 &  x1007 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1073 &  x1076 &  x1094 &  x1097 &  x1106 &  x1112 &  x1121 &  x1124 &  x1127 & ~x81 & ~x82 & ~x168 & ~x330 & ~x363 & ~x627 & ~x780 & ~x819;
assign c5224 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x50 &  x53 &  x56 &  x59 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x431 &  x434 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x590 &  x593 &  x596 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x628 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x698 &  x701 &  x704 &  x707 &  x713 &  x716 &  x722 &  x725 &  x728 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x761 &  x764 &  x767 &  x773 &  x776 &  x779 &  x782 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x854 &  x857 &  x860 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x929 &  x938 &  x941 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1039 &  x1040 &  x1046 &  x1049 &  x1055 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1078 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 &  x1130 & ~x159 & ~x198 & ~x199 & ~x237 & ~x246 & ~x324 & ~x402 & ~x780 & ~x819 & ~x858 & ~x897 & ~x936 & ~x1014 & ~x1047 & ~x1053 & ~x1086 & ~x1092 & ~x1125;
assign c5226 =  x5 &  x14 &  x23 &  x32 &  x38 &  x41 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x101 &  x107 &  x113 &  x116 &  x119 &  x128 &  x131 &  x134 &  x146 &  x149 &  x152 &  x155 &  x158 &  x167 &  x173 &  x179 &  x185 &  x191 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x233 &  x236 &  x245 &  x248 &  x251 &  x254 &  x257 &  x263 &  x269 &  x272 &  x274 &  x275 &  x278 &  x284 &  x287 &  x296 &  x305 &  x311 &  x317 &  x320 &  x323 &  x326 &  x335 &  x341 &  x344 &  x350 &  x362 &  x365 &  x368 &  x371 &  x374 &  x380 &  x386 &  x389 &  x392 &  x398 &  x407 &  x410 &  x413 &  x419 &  x425 &  x428 &  x434 &  x437 &  x440 &  x443 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x470 &  x476 &  x479 &  x482 &  x485 &  x488 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x545 &  x557 &  x575 &  x581 &  x584 &  x587 &  x589 &  x593 &  x596 &  x605 &  x608 &  x610 &  x611 &  x614 &  x616 &  x617 &  x620 &  x632 &  x638 &  x641 &  x644 &  x650 &  x655 &  x656 &  x665 &  x668 &  x671 &  x677 &  x680 &  x683 &  x689 &  x692 &  x694 &  x695 &  x698 &  x701 &  x704 &  x710 &  x719 &  x722 &  x725 &  x728 &  x731 &  x737 &  x740 &  x746 &  x752 &  x755 &  x758 &  x764 &  x766 &  x767 &  x770 &  x772 &  x785 &  x794 &  x800 &  x803 &  x806 &  x809 &  x815 &  x818 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x845 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x869 &  x875 &  x878 &  x887 &  x890 &  x893 &  x896 &  x908 &  x911 &  x914 &  x923 &  x926 &  x929 &  x944 &  x947 &  x950 &  x956 &  x959 &  x965 &  x974 &  x980 &  x983 &  x989 &  x992 &  x1001 &  x1004 &  x1010 &  x1013 &  x1021 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1091 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1118 &  x1121 &  x1127 & ~x519 & ~x558 & ~x561 & ~x600 & ~x639 & ~x741;
assign c5228 =  x8 &  x11 &  x14 &  x20 &  x35 &  x47 &  x50 &  x62 &  x74 &  x80 &  x83 &  x89 &  x98 &  x107 &  x110 &  x119 &  x128 &  x137 &  x140 &  x143 &  x161 &  x170 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x206 &  x215 &  x218 &  x224 &  x230 &  x233 &  x236 &  x248 &  x254 &  x257 &  x263 &  x272 &  x275 &  x278 &  x284 &  x287 &  x296 &  x302 &  x311 &  x313 &  x323 &  x332 &  x335 &  x344 &  x356 &  x359 &  x371 &  x374 &  x391 &  x401 &  x407 &  x410 &  x422 &  x434 &  x437 &  x440 &  x443 &  x464 &  x470 &  x488 &  x494 &  x497 &  x500 &  x512 &  x518 &  x521 &  x524 &  x527 &  x542 &  x545 &  x551 &  x554 &  x569 &  x572 &  x584 &  x590 &  x593 &  x596 &  x599 &  x605 &  x608 &  x614 &  x620 &  x626 &  x632 &  x635 &  x638 &  x650 &  x671 &  x677 &  x683 &  x704 &  x707 &  x710 &  x716 &  x725 &  x728 &  x731 &  x734 &  x737 &  x752 &  x755 &  x764 &  x767 &  x776 &  x779 &  x785 &  x797 &  x803 &  x830 &  x839 &  x842 &  x848 &  x851 &  x878 &  x881 &  x893 &  x896 &  x899 &  x902 &  x914 &  x920 &  x932 &  x941 &  x944 &  x950 &  x959 &  x965 &  x983 &  x986 &  x989 &  x992 &  x1001 &  x1004 &  x1010 &  x1013 &  x1018 &  x1022 &  x1025 &  x1034 &  x1043 &  x1046 &  x1073 &  x1079 &  x1091 &  x1094 &  x1106 &  x1112 &  x1115 &  x1118 &  x1130 & ~x18 & ~x57 & ~x114 & ~x135 & ~x231 & ~x270 & ~x336 & ~x363 & ~x480 & ~x558 & ~x564 & ~x753 & ~x792;
assign c5230 =  x2 &  x8 &  x14 &  x20 &  x29 &  x44 &  x77 &  x89 &  x98 &  x101 &  x116 &  x125 &  x143 &  x164 &  x170 &  x176 &  x203 &  x215 &  x218 &  x230 &  x236 &  x248 &  x260 &  x278 &  x293 &  x311 &  x314 &  x323 &  x326 &  x332 &  x347 &  x353 &  x362 &  x371 &  x374 &  x380 &  x392 &  x410 &  x431 &  x443 &  x449 &  x476 &  x479 &  x497 &  x512 &  x530 &  x542 &  x563 &  x566 &  x596 &  x602 &  x605 &  x608 &  x614 &  x629 &  x644 &  x656 &  x662 &  x665 &  x674 &  x683 &  x689 &  x692 &  x695 &  x701 &  x719 &  x740 &  x758 &  x764 &  x800 &  x803 &  x818 &  x833 &  x839 &  x842 &  x869 &  x890 &  x908 &  x917 &  x923 &  x926 &  x935 &  x940 &  x941 &  x986 &  x989 &  x1001 &  x1007 &  x1013 &  x1016 &  x1031 &  x1040 &  x1046 &  x1052 &  x1061 &  x1064 &  x1067 &  x1073 &  x1091 &  x1100 &  x1103 &  x1118 &  x1124 &  x1127 & ~x246 & ~x363 & ~x375 & ~x381 & ~x643;
assign c5232 =  x8 &  x11 &  x20 &  x26 &  x29 &  x32 &  x35 &  x41 &  x50 &  x53 &  x56 &  x65 &  x71 &  x74 &  x77 &  x80 &  x89 &  x95 &  x98 &  x104 &  x107 &  x113 &  x116 &  x125 &  x128 &  x131 &  x143 &  x149 &  x157 &  x161 &  x170 &  x176 &  x188 &  x191 &  x194 &  x196 &  x197 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x274 &  x275 &  x278 &  x284 &  x287 &  x290 &  x296 &  x299 &  x308 &  x311 &  x313 &  x314 &  x317 &  x323 &  x326 &  x329 &  x332 &  x338 &  x344 &  x347 &  x352 &  x368 &  x377 &  x380 &  x383 &  x386 &  x395 &  x404 &  x407 &  x410 &  x416 &  x425 &  x428 &  x431 &  x440 &  x461 &  x464 &  x470 &  x482 &  x485 &  x491 &  x494 &  x497 &  x500 &  x509 &  x512 &  x518 &  x524 &  x527 &  x530 &  x536 &  x542 &  x551 &  x554 &  x566 &  x572 &  x578 &  x581 &  x584 &  x590 &  x593 &  x599 &  x602 &  x605 &  x610 &  x611 &  x614 &  x623 &  x626 &  x629 &  x644 &  x647 &  x656 &  x668 &  x677 &  x683 &  x686 &  x695 &  x707 &  x710 &  x719 &  x727 &  x728 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x761 &  x776 &  x788 &  x791 &  x794 &  x797 &  x800 &  x809 &  x821 &  x824 &  x839 &  x842 &  x845 &  x848 &  x860 &  x869 &  x881 &  x890 &  x893 &  x902 &  x908 &  x920 &  x923 &  x929 &  x938 &  x947 &  x953 &  x968 &  x974 &  x980 &  x989 &  x992 &  x1007 &  x1016 &  x1028 &  x1031 &  x1043 &  x1046 &  x1049 &  x1055 &  x1061 &  x1067 &  x1070 &  x1073 &  x1079 &  x1100 &  x1103 & ~x42 & ~x81 & ~x82 & ~x141 & ~x180 & ~x225 & ~x264 & ~x265 & ~x303 & ~x369 & ~x444 & ~x861;
assign c5234 =  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x40 &  x41 &  x44 &  x47 &  x50 &  x53 &  x59 &  x65 &  x68 &  x71 &  x74 &  x77 &  x79 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x101 &  x104 &  x107 &  x113 &  x116 &  x118 &  x119 &  x122 &  x125 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x157 &  x161 &  x164 &  x170 &  x173 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x195 &  x196 &  x197 &  x203 &  x206 &  x209 &  x212 &  x218 &  x221 &  x227 &  x230 &  x233 &  x234 &  x235 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x272 &  x273 &  x274 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x311 &  x313 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x431 &  x433 &  x434 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x464 &  x467 &  x470 &  x472 &  x473 &  x479 &  x482 &  x485 &  x491 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x527 &  x530 &  x536 &  x539 &  x545 &  x551 &  x554 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x659 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x728 &  x731 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x770 &  x776 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x833 &  x836 &  x839 &  x842 &  x845 &  x851 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x959 &  x968 &  x971 &  x977 &  x980 &  x983 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x24 & ~x42 & ~x63 & ~x141 & ~x147 & ~x148 & ~x180 & ~x186 & ~x207 & ~x225 & ~x246 & ~x264 & ~x444;
assign c5236 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x23 &  x29 &  x41 &  x44 &  x47 &  x50 &  x53 &  x59 &  x62 &  x65 &  x71 &  x74 &  x77 &  x86 &  x89 &  x95 &  x98 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x146 &  x152 &  x155 &  x158 &  x161 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x275 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x335 &  x341 &  x350 &  x352 &  x353 &  x356 &  x362 &  x365 &  x368 &  x371 &  x374 &  x383 &  x386 &  x389 &  x391 &  x392 &  x395 &  x398 &  x401 &  x404 &  x410 &  x413 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x440 &  x452 &  x455 &  x458 &  x464 &  x467 &  x469 &  x473 &  x476 &  x479 &  x482 &  x485 &  x491 &  x494 &  x500 &  x503 &  x508 &  x509 &  x512 &  x515 &  x521 &  x527 &  x530 &  x533 &  x536 &  x539 &  x545 &  x547 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x584 &  x587 &  x590 &  x593 &  x599 &  x602 &  x608 &  x611 &  x617 &  x620 &  x623 &  x626 &  x628 &  x629 &  x632 &  x635 &  x638 &  x644 &  x647 &  x650 &  x653 &  x656 &  x662 &  x665 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x722 &  x725 &  x728 &  x737 &  x740 &  x743 &  x749 &  x758 &  x761 &  x767 &  x770 &  x776 &  x779 &  x782 &  x785 &  x794 &  x797 &  x800 &  x806 &  x809 &  x824 &  x827 &  x830 &  x839 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x881 &  x884 &  x887 &  x890 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x956 &  x959 &  x965 &  x968 &  x971 &  x977 &  x980 &  x983 &  x989 &  x992 &  x998 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1067 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 & ~x198 & ~x237 & ~x238 & ~x276 & ~x277 & ~x316 & ~x354 & ~x600 & ~x603;
assign c5238 =  x50 &  x89 &  x92 &  x110 &  x152 &  x179 &  x212 &  x242 &  x260 &  x335 &  x344 &  x398 &  x444 &  x457 &  x461 &  x509 &  x539 &  x557 &  x581 &  x584 &  x614 &  x623 &  x626 &  x629 &  x635 &  x659 &  x665 &  x710 &  x716 &  x743 &  x749 &  x752 &  x794 &  x848 &  x872 &  x896 &  x899 &  x911 &  x920 &  x986 &  x1004 &  x1018 &  x1076 &  x1106 & ~x471 & ~x477 & ~x570 & ~x831 & ~x870;
assign c5240 =  x32 &  x38 &  x44 &  x47 &  x65 &  x77 &  x95 &  x98 &  x128 &  x137 &  x149 &  x158 &  x188 &  x197 &  x218 &  x224 &  x290 &  x320 &  x335 &  x338 &  x404 &  x416 &  x497 &  x536 &  x542 &  x551 &  x608 &  x644 &  x668 &  x689 &  x701 &  x722 &  x734 &  x737 &  x740 &  x788 &  x823 &  x830 &  x845 &  x889 &  x905 &  x929 &  x968 &  x980 &  x1010 &  x1031 &  x1100 & ~x237 & ~x324 & ~x453 & ~x480 & ~x519 & ~x678 & ~x795 & ~x796;
assign c5242 =  x2 &  x14 &  x17 &  x44 &  x59 &  x137 &  x149 &  x203 &  x206 &  x215 &  x227 &  x257 &  x269 &  x293 &  x305 &  x332 &  x341 &  x347 &  x350 &  x359 &  x398 &  x419 &  x422 &  x449 &  x482 &  x503 &  x566 &  x596 &  x602 &  x611 &  x614 &  x638 &  x644 &  x653 &  x656 &  x659 &  x674 &  x701 &  x713 &  x728 &  x737 &  x740 &  x761 &  x764 &  x776 &  x803 &  x821 &  x857 &  x860 &  x863 &  x866 &  x950 &  x977 &  x989 &  x995 &  x1004 &  x1007 &  x1013 &  x1015 &  x1022 &  x1056 &  x1058 &  x1064 &  x1076 & ~x195 & ~x546 & ~x549 & ~x628 & ~x714 & ~x987;
assign c5244 =  x2 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x74 &  x77 &  x80 &  x89 &  x92 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x125 &  x128 &  x131 &  x137 &  x140 &  x143 &  x152 &  x155 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x194 &  x197 &  x200 &  x203 &  x209 &  x212 &  x215 &  x218 &  x221 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x260 &  x263 &  x266 &  x272 &  x275 &  x278 &  x290 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x314 &  x317 &  x320 &  x323 &  x326 &  x332 &  x335 &  x338 &  x344 &  x350 &  x353 &  x359 &  x362 &  x365 &  x368 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x404 &  x407 &  x410 &  x413 &  x419 &  x425 &  x428 &  x431 &  x437 &  x443 &  x446 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x479 &  x482 &  x488 &  x494 &  x497 &  x503 &  x506 &  x509 &  x524 &  x527 &  x533 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x587 &  x590 &  x593 &  x602 &  x605 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x731 &  x734 &  x737 &  x740 &  x743 &  x755 &  x758 &  x761 &  x770 &  x773 &  x779 &  x785 &  x788 &  x791 &  x794 &  x797 &  x803 &  x806 &  x809 &  x812 &  x815 &  x821 &  x824 &  x827 &  x830 &  x833 &  x842 &  x845 &  x851 &  x857 &  x860 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x902 &  x905 &  x908 &  x920 &  x923 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x950 &  x953 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x3 & ~x4 & ~x42 & ~x43 & ~x90 & ~x129 & ~x168 & ~x169 & ~x208 & ~x246 & ~x324 & ~x325 & ~x402 & ~x639 & ~x741 & ~x819 & ~x858 & ~x897 & ~x936 & ~x1053;
assign c5246 =  x2 &  x5 &  x14 &  x17 &  x23 &  x29 &  x32 &  x41 &  x44 &  x56 &  x59 &  x62 &  x65 &  x68 &  x79 &  x83 &  x89 &  x92 &  x95 &  x101 &  x107 &  x125 &  x131 &  x146 &  x149 &  x152 &  x155 &  x157 &  x158 &  x161 &  x164 &  x167 &  x173 &  x182 &  x188 &  x194 &  x196 &  x197 &  x203 &  x206 &  x212 &  x221 &  x227 &  x230 &  x236 &  x248 &  x251 &  x254 &  x257 &  x263 &  x266 &  x272 &  x274 &  x275 &  x296 &  x308 &  x311 &  x313 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x356 &  x362 &  x365 &  x371 &  x383 &  x386 &  x389 &  x398 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x428 &  x431 &  x440 &  x446 &  x452 &  x461 &  x464 &  x473 &  x479 &  x482 &  x485 &  x488 &  x491 &  x497 &  x506 &  x509 &  x521 &  x524 &  x527 &  x545 &  x548 &  x551 &  x557 &  x566 &  x571 &  x572 &  x578 &  x581 &  x587 &  x590 &  x596 &  x602 &  x610 &  x614 &  x620 &  x623 &  x629 &  x635 &  x638 &  x649 &  x650 &  x653 &  x656 &  x659 &  x662 &  x671 &  x686 &  x689 &  x692 &  x698 &  x701 &  x704 &  x707 &  x713 &  x716 &  x719 &  x727 &  x731 &  x737 &  x743 &  x749 &  x755 &  x758 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x812 &  x815 &  x821 &  x830 &  x836 &  x845 &  x850 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x884 &  x887 &  x893 &  x911 &  x914 &  x923 &  x929 &  x932 &  x938 &  x947 &  x950 &  x953 &  x965 &  x968 &  x977 &  x980 &  x986 &  x992 &  x998 &  x1001 &  x1007 &  x1010 &  x1016 &  x1019 &  x1022 &  x1031 &  x1037 &  x1046 &  x1049 &  x1052 &  x1058 &  x1067 &  x1073 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1112 &  x1121 &  x1124 &  x1130 & ~x36 & ~x42 & ~x594 & ~x633 & ~x672 & ~x711 & ~x741 & ~x780 & ~x858;
assign c5248 =  x8 &  x17 &  x29 &  x35 &  x38 &  x41 &  x44 &  x50 &  x53 &  x56 &  x59 &  x65 &  x68 &  x71 &  x79 &  x80 &  x86 &  x92 &  x98 &  x101 &  x107 &  x110 &  x118 &  x119 &  x122 &  x125 &  x131 &  x137 &  x140 &  x146 &  x149 &  x155 &  x158 &  x161 &  x167 &  x170 &  x173 &  x176 &  x182 &  x185 &  x191 &  x194 &  x195 &  x196 &  x200 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x233 &  x235 &  x236 &  x245 &  x248 &  x257 &  x260 &  x263 &  x266 &  x274 &  x278 &  x281 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x314 &  x317 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x368 &  x371 &  x392 &  x395 &  x398 &  x401 &  x404 &  x410 &  x416 &  x431 &  x440 &  x446 &  x452 &  x455 &  x464 &  x470 &  x473 &  x479 &  x485 &  x488 &  x497 &  x500 &  x506 &  x512 &  x518 &  x521 &  x524 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x590 &  x596 &  x599 &  x602 &  x605 &  x608 &  x614 &  x617 &  x626 &  x629 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x665 &  x680 &  x683 &  x695 &  x698 &  x713 &  x725 &  x728 &  x731 &  x740 &  x743 &  x746 &  x752 &  x755 &  x764 &  x773 &  x785 &  x788 &  x797 &  x800 &  x803 &  x806 &  x812 &  x821 &  x830 &  x833 &  x838 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x866 &  x872 &  x878 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x917 &  x926 &  x929 &  x932 &  x944 &  x947 &  x950 &  x956 &  x959 &  x968 &  x977 &  x980 &  x986 &  x989 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1034 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1105 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 & ~x12 & ~x13 & ~x52 & ~x90 & ~x192 & ~x207 & ~x246 & ~x247 & ~x285 & ~x324 & ~x325;
assign c5250 =  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x56 &  x65 &  x74 &  x83 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x116 &  x128 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x158 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x203 &  x206 &  x212 &  x221 &  x224 &  x230 &  x233 &  x236 &  x242 &  x245 &  x248 &  x254 &  x266 &  x269 &  x272 &  x275 &  x278 &  x284 &  x287 &  x290 &  x293 &  x296 &  x302 &  x305 &  x308 &  x311 &  x314 &  x320 &  x323 &  x335 &  x338 &  x341 &  x347 &  x359 &  x362 &  x368 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x395 &  x404 &  x407 &  x419 &  x422 &  x425 &  x434 &  x443 &  x446 &  x449 &  x452 &  x458 &  x467 &  x470 &  x476 &  x479 &  x485 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x524 &  x530 &  x536 &  x539 &  x542 &  x551 &  x560 &  x563 &  x566 &  x569 &  x572 &  x574 &  x578 &  x590 &  x593 &  x596 &  x599 &  x605 &  x608 &  x611 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x638 &  x641 &  x644 &  x653 &  x659 &  x662 &  x665 &  x668 &  x677 &  x680 &  x683 &  x692 &  x698 &  x701 &  x704 &  x713 &  x719 &  x722 &  x725 &  x728 &  x740 &  x743 &  x755 &  x758 &  x761 &  x767 &  x773 &  x776 &  x779 &  x782 &  x784 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x812 &  x815 &  x821 &  x827 &  x830 &  x833 &  x839 &  x842 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x875 &  x878 &  x881 &  x887 &  x890 &  x896 &  x899 &  x908 &  x917 &  x920 &  x929 &  x932 &  x941 &  x944 &  x953 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1094 &  x1100 &  x1106 &  x1112 &  x1130 & ~x198 & ~x441 & ~x442 & ~x480 & ~x481 & ~x519 & ~x520 & ~x756 & ~x795;
assign c5252 =  x8 &  x23 &  x29 &  x44 &  x80 &  x125 &  x140 &  x143 &  x146 &  x221 &  x242 &  x290 &  x296 &  x302 &  x308 &  x320 &  x326 &  x347 &  x350 &  x398 &  x425 &  x431 &  x452 &  x485 &  x488 &  x515 &  x533 &  x542 &  x560 &  x575 &  x578 &  x581 &  x599 &  x638 &  x647 &  x650 &  x668 &  x683 &  x701 &  x704 &  x707 &  x713 &  x764 &  x775 &  x776 &  x781 &  x785 &  x815 &  x830 &  x842 &  x893 &  x902 &  x938 &  x959 &  x968 &  x974 &  x983 &  x1040 &  x1055 &  x1067 &  x1073 &  x1085 & ~x315 & ~x589 & ~x714 & ~x831 & ~x849 & ~x870 & ~x909 & ~x910 & ~x987;
assign c5254 =  x2 &  x8 &  x11 &  x14 &  x20 &  x29 &  x38 &  x44 &  x47 &  x68 &  x74 &  x80 &  x83 &  x86 &  x92 &  x95 &  x103 &  x107 &  x119 &  x122 &  x128 &  x131 &  x137 &  x143 &  x155 &  x167 &  x173 &  x179 &  x182 &  x185 &  x191 &  x209 &  x212 &  x233 &  x242 &  x260 &  x275 &  x281 &  x284 &  x287 &  x290 &  x299 &  x302 &  x311 &  x323 &  x329 &  x332 &  x335 &  x338 &  x356 &  x362 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x389 &  x392 &  x395 &  x401 &  x416 &  x434 &  x437 &  x464 &  x473 &  x479 &  x485 &  x494 &  x497 &  x503 &  x509 &  x512 &  x518 &  x527 &  x530 &  x533 &  x539 &  x542 &  x548 &  x566 &  x569 &  x572 &  x587 &  x596 &  x602 &  x608 &  x617 &  x623 &  x632 &  x644 &  x647 &  x653 &  x662 &  x665 &  x695 &  x704 &  x710 &  x719 &  x722 &  x734 &  x737 &  x755 &  x758 &  x764 &  x773 &  x776 &  x785 &  x806 &  x809 &  x815 &  x818 &  x833 &  x836 &  x839 &  x842 &  x845 &  x854 &  x857 &  x863 &  x878 &  x881 &  x884 &  x890 &  x896 &  x899 &  x902 &  x908 &  x911 &  x920 &  x929 &  x932 &  x944 &  x968 &  x971 &  x974 &  x977 &  x986 &  x1001 &  x1004 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1028 &  x1037 &  x1046 &  x1049 &  x1055 &  x1058 &  x1067 &  x1076 &  x1088 &  x1091 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 & ~x27 & ~x78 & ~x156 & ~x276 & ~x324 & ~x354 & ~x355 & ~x393 & ~x486 & ~x525 & ~x564;
assign c5256 =  x23 &  x32 &  x47 &  x65 &  x68 &  x71 &  x80 &  x83 &  x89 &  x92 &  x101 &  x104 &  x152 &  x155 &  x173 &  x233 &  x260 &  x287 &  x296 &  x302 &  x326 &  x335 &  x389 &  x395 &  x398 &  x401 &  x410 &  x431 &  x446 &  x464 &  x476 &  x482 &  x485 &  x494 &  x503 &  x509 &  x533 &  x536 &  x578 &  x608 &  x638 &  x641 &  x668 &  x680 &  x698 &  x706 &  x707 &  x710 &  x719 &  x734 &  x737 &  x746 &  x749 &  x761 &  x764 &  x782 &  x824 &  x842 &  x851 &  x866 &  x869 &  x878 &  x895 &  x905 &  x914 &  x920 &  x932 &  x938 &  x944 &  x947 &  x956 &  x977 &  x986 &  x992 &  x998 &  x1007 &  x1025 &  x1040 &  x1046 &  x1061 &  x1067 &  x1091 &  x1094 &  x1118 & ~x394 & ~x408 & ~x486 & ~x603 & ~x717;
assign c5258 =  x23 &  x26 &  x29 &  x41 &  x59 &  x68 &  x74 &  x80 &  x95 &  x140 &  x143 &  x182 &  x206 &  x230 &  x233 &  x242 &  x251 &  x305 &  x341 &  x365 &  x395 &  x401 &  x405 &  x407 &  x416 &  x431 &  x437 &  x440 &  x452 &  x470 &  x482 &  x488 &  x491 &  x497 &  x500 &  x506 &  x512 &  x518 &  x524 &  x527 &  x539 &  x557 &  x563 &  x566 &  x572 &  x578 &  x599 &  x626 &  x629 &  x635 &  x656 &  x662 &  x674 &  x677 &  x686 &  x689 &  x701 &  x707 &  x710 &  x722 &  x725 &  x728 &  x740 &  x746 &  x752 &  x764 &  x767 &  x779 &  x812 &  x839 &  x869 &  x878 &  x917 &  x926 &  x929 &  x992 &  x998 &  x1001 &  x1013 &  x1022 &  x1031 &  x1043 &  x1064 &  x1073 &  x1082 &  x1091 &  x1094 &  x1103 &  x1106 &  x1109 &  x1121 &  x1130 & ~x273 & ~x354 & ~x390 & ~x1068;
assign c5260 =  x11 &  x14 &  x26 &  x29 &  x32 &  x41 &  x56 &  x59 &  x83 &  x95 &  x104 &  x110 &  x116 &  x128 &  x140 &  x173 &  x176 &  x191 &  x212 &  x230 &  x233 &  x236 &  x248 &  x257 &  x284 &  x299 &  x302 &  x311 &  x314 &  x317 &  x320 &  x329 &  x335 &  x344 &  x347 &  x356 &  x362 &  x380 &  x404 &  x407 &  x410 &  x413 &  x416 &  x425 &  x428 &  x437 &  x440 &  x452 &  x458 &  x469 &  x479 &  x494 &  x506 &  x548 &  x554 &  x557 &  x566 &  x569 &  x578 &  x589 &  x599 &  x605 &  x614 &  x620 &  x632 &  x665 &  x677 &  x695 &  x704 &  x706 &  x707 &  x713 &  x719 &  x728 &  x743 &  x758 &  x761 &  x764 &  x766 &  x782 &  x812 &  x824 &  x827 &  x851 &  x854 &  x890 &  x908 &  x926 &  x947 &  x959 &  x980 &  x983 &  x1004 &  x1007 &  x1010 &  x1019 &  x1052 &  x1070 &  x1073 &  x1097 &  x1112 & ~x160 & ~x198 & ~x231 & ~x246 & ~x297 & ~x519;
assign c5262 =  x5 &  x8 &  x20 &  x23 &  x26 &  x29 &  x35 &  x38 &  x40 &  x41 &  x50 &  x59 &  x62 &  x67 &  x68 &  x71 &  x72 &  x73 &  x74 &  x79 &  x80 &  x86 &  x89 &  x92 &  x101 &  x107 &  x119 &  x122 &  x128 &  x134 &  x140 &  x143 &  x157 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x182 &  x194 &  x196 &  x197 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x227 &  x235 &  x239 &  x245 &  x251 &  x257 &  x260 &  x272 &  x274 &  x281 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x313 &  x320 &  x323 &  x326 &  x329 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x368 &  x377 &  x389 &  x392 &  x395 &  x401 &  x413 &  x431 &  x434 &  x440 &  x443 &  x449 &  x455 &  x461 &  x470 &  x482 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x521 &  x524 &  x527 &  x530 &  x539 &  x557 &  x560 &  x563 &  x566 &  x572 &  x575 &  x590 &  x593 &  x599 &  x602 &  x608 &  x611 &  x617 &  x620 &  x622 &  x632 &  x635 &  x638 &  x650 &  x653 &  x659 &  x662 &  x671 &  x680 &  x689 &  x692 &  x698 &  x707 &  x713 &  x731 &  x740 &  x749 &  x758 &  x764 &  x767 &  x770 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x797 &  x800 &  x806 &  x821 &  x827 &  x830 &  x833 &  x839 &  x841 &  x842 &  x848 &  x851 &  x854 &  x857 &  x866 &  x869 &  x872 &  x878 &  x881 &  x884 &  x887 &  x896 &  x899 &  x902 &  x905 &  x911 &  x917 &  x920 &  x926 &  x928 &  x929 &  x944 &  x950 &  x956 &  x959 &  x962 &  x965 &  x967 &  x968 &  x974 &  x977 &  x983 &  x986 &  x989 &  x998 &  x1004 &  x1007 &  x1010 &  x1013 &  x1019 &  x1025 &  x1028 &  x1030 &  x1034 &  x1037 &  x1040 &  x1043 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1069 &  x1070 &  x1073 &  x1076 &  x1082 &  x1094 &  x1097 &  x1100 &  x1103 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x477 & ~x516 & ~x555;
assign c5264 =  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x44 &  x47 &  x50 &  x53 &  x62 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x118 &  x119 &  x125 &  x128 &  x134 &  x140 &  x146 &  x149 &  x152 &  x155 &  x157 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x179 &  x182 &  x185 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x224 &  x230 &  x233 &  x235 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x269 &  x272 &  x275 &  x278 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x311 &  x312 &  x313 &  x314 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x341 &  x347 &  x350 &  x352 &  x353 &  x362 &  x368 &  x371 &  x377 &  x383 &  x386 &  x389 &  x391 &  x392 &  x395 &  x398 &  x404 &  x410 &  x413 &  x419 &  x422 &  x428 &  x433 &  x434 &  x437 &  x440 &  x443 &  x446 &  x452 &  x455 &  x458 &  x464 &  x467 &  x470 &  x472 &  x473 &  x479 &  x482 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x509 &  x511 &  x512 &  x515 &  x518 &  x521 &  x530 &  x536 &  x539 &  x542 &  x550 &  x551 &  x563 &  x566 &  x569 &  x572 &  x575 &  x581 &  x584 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x635 &  x638 &  x644 &  x647 &  x650 &  x653 &  x656 &  x668 &  x674 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x701 &  x704 &  x707 &  x710 &  x716 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x776 &  x779 &  x782 &  x788 &  x791 &  x794 &  x797 &  x803 &  x806 &  x809 &  x812 &  x818 &  x821 &  x824 &  x827 &  x833 &  x839 &  x845 &  x848 &  x854 &  x857 &  x863 &  x875 &  x878 &  x881 &  x884 &  x887 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x917 &  x920 &  x923 &  x926 &  x932 &  x938 &  x941 &  x947 &  x950 &  x953 &  x956 &  x959 &  x965 &  x968 &  x974 &  x977 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1124 &  x1130 & ~x159 & ~x160 & ~x483 & ~x523 & ~x561 & ~x600;
assign c5266 =  x5 &  x11 &  x17 &  x20 &  x26 &  x29 &  x40 &  x50 &  x59 &  x62 &  x68 &  x74 &  x77 &  x79 &  x83 &  x89 &  x95 &  x98 &  x104 &  x110 &  x116 &  x118 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x155 &  x157 &  x164 &  x167 &  x170 &  x182 &  x185 &  x191 &  x194 &  x196 &  x200 &  x203 &  x206 &  x209 &  x218 &  x221 &  x224 &  x227 &  x233 &  x242 &  x257 &  x260 &  x266 &  x272 &  x275 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x314 &  x317 &  x320 &  x323 &  x326 &  x332 &  x341 &  x344 &  x350 &  x353 &  x356 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x389 &  x401 &  x404 &  x407 &  x413 &  x422 &  x428 &  x431 &  x434 &  x446 &  x449 &  x455 &  x461 &  x464 &  x467 &  x470 &  x473 &  x482 &  x485 &  x488 &  x494 &  x497 &  x500 &  x506 &  x512 &  x515 &  x521 &  x524 &  x527 &  x530 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x563 &  x566 &  x584 &  x587 &  x593 &  x596 &  x608 &  x614 &  x617 &  x623 &  x629 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x662 &  x665 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x704 &  x710 &  x716 &  x737 &  x743 &  x749 &  x752 &  x755 &  x767 &  x773 &  x779 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x806 &  x809 &  x818 &  x827 &  x830 &  x833 &  x836 &  x842 &  x845 &  x848 &  x851 &  x854 &  x860 &  x866 &  x872 &  x881 &  x884 &  x887 &  x899 &  x902 &  x905 &  x908 &  x911 &  x917 &  x920 &  x923 &  x926 &  x941 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1016 &  x1019 &  x1022 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1052 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1091 &  x1094 &  x1097 &  x1100 &  x1112 &  x1118 &  x1127 & ~x42 & ~x148 & ~x186 & ~x187 & ~x225 & ~x246 & ~x264 & ~x288 & ~x327 & ~x366 & ~x367 & ~x405 & ~x406 & ~x444 & ~x483 & ~x633 & ~x741 & ~x780 & ~x819;
assign c5268 =  x2 &  x11 &  x50 &  x62 &  x68 &  x80 &  x104 &  x110 &  x122 &  x161 &  x176 &  x182 &  x185 &  x233 &  x239 &  x248 &  x254 &  x257 &  x263 &  x272 &  x275 &  x284 &  x296 &  x302 &  x308 &  x317 &  x341 &  x353 &  x368 &  x383 &  x401 &  x407 &  x434 &  x440 &  x467 &  x479 &  x488 &  x503 &  x515 &  x533 &  x551 &  x560 &  x563 &  x572 &  x578 &  x599 &  x623 &  x638 &  x647 &  x662 &  x670 &  x734 &  x749 &  x773 &  x782 &  x797 &  x809 &  x820 &  x821 &  x830 &  x839 &  x857 &  x858 &  x890 &  x898 &  x902 &  x908 &  x914 &  x917 &  x938 &  x941 &  x947 &  x956 &  x971 &  x974 &  x989 &  x1001 &  x1007 &  x1010 &  x1016 &  x1017 &  x1018 &  x1022 &  x1052 &  x1070 &  x1082 &  x1085 &  x1088 &  x1100 &  x1103 &  x1121 &  x1127 & ~x399 & ~x429 & ~x667 & ~x948;
assign c5270 =  x38 &  x41 &  x71 &  x158 &  x167 &  x188 &  x242 &  x269 &  x296 &  x332 &  x344 &  x407 &  x437 &  x440 &  x452 &  x473 &  x522 &  x527 &  x599 &  x701 &  x716 &  x752 &  x755 &  x836 &  x896 &  x911 &  x923 &  x983 &  x998 &  x1061 &  x1096 &  x1106 & ~x165 & ~x351 & ~x510 & ~x550 & ~x792;
assign c5272 =  x8 &  x14 &  x68 &  x83 &  x95 &  x116 &  x125 &  x170 &  x197 &  x200 &  x202 &  x215 &  x233 &  x245 &  x251 &  x269 &  x281 &  x299 &  x314 &  x317 &  x352 &  x362 &  x368 &  x377 &  x404 &  x407 &  x416 &  x422 &  x430 &  x440 &  x443 &  x452 &  x470 &  x473 &  x485 &  x548 &  x557 &  x587 &  x605 &  x628 &  x638 &  x671 &  x674 &  x716 &  x722 &  x734 &  x746 &  x749 &  x761 &  x773 &  x809 &  x824 &  x836 &  x845 &  x848 &  x851 &  x878 &  x890 &  x902 &  x920 &  x926 &  x935 &  x953 &  x986 &  x995 &  x1004 &  x1034 &  x1058 &  x1094 &  x1103 &  x1109 &  x1115 &  x1124 & ~x355;
assign c5274 =  x2 &  x14 &  x29 &  x44 &  x50 &  x56 &  x59 &  x74 &  x80 &  x89 &  x101 &  x110 &  x113 &  x149 &  x179 &  x191 &  x200 &  x209 &  x212 &  x239 &  x245 &  x251 &  x260 &  x266 &  x272 &  x293 &  x338 &  x350 &  x371 &  x380 &  x386 &  x392 &  x407 &  x422 &  x440 &  x475 &  x482 &  x500 &  x503 &  x509 &  x518 &  x521 &  x530 &  x536 &  x542 &  x551 &  x553 &  x563 &  x572 &  x581 &  x592 &  x593 &  x602 &  x605 &  x608 &  x617 &  x650 &  x653 &  x683 &  x689 &  x692 &  x701 &  x722 &  x728 &  x742 &  x743 &  x764 &  x791 &  x797 &  x800 &  x803 &  x806 &  x815 &  x818 &  x860 &  x866 &  x869 &  x875 &  x881 &  x887 &  x899 &  x902 &  x926 &  x932 &  x940 &  x941 &  x968 &  x979 &  x1007 &  x1016 &  x1025 &  x1034 &  x1037 &  x1046 &  x1049 &  x1061 &  x1064 &  x1076 &  x1079 &  x1085 &  x1097 &  x1100 &  x1106 &  x1115 &  x1121 &  x1127 & ~x273 & ~x351 & ~x471 & ~x550 & ~x621;
assign c5276 =  x1 &  x5 &  x8 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x40 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x79 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x101 &  x104 &  x110 &  x116 &  x118 &  x122 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x161 &  x164 &  x167 &  x170 &  x176 &  x179 &  x188 &  x191 &  x194 &  x196 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x235 &  x236 &  x239 &  x245 &  x248 &  x251 &  x257 &  x260 &  x263 &  x269 &  x272 &  x274 &  x275 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x308 &  x311 &  x313 &  x314 &  x317 &  x320 &  x323 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x355 &  x356 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x433 &  x434 &  x440 &  x443 &  x446 &  x452 &  x458 &  x461 &  x467 &  x473 &  x476 &  x479 &  x482 &  x488 &  x491 &  x494 &  x503 &  x506 &  x509 &  x512 &  x515 &  x527 &  x530 &  x536 &  x542 &  x548 &  x551 &  x554 &  x560 &  x563 &  x566 &  x569 &  x575 &  x581 &  x584 &  x587 &  x590 &  x602 &  x605 &  x608 &  x611 &  x617 &  x620 &  x623 &  x626 &  x629 &  x635 &  x638 &  x641 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x698 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x815 &  x818 &  x821 &  x824 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x854 &  x857 &  x860 &  x866 &  x869 &  x872 &  x878 &  x881 &  x884 &  x887 &  x890 &  x899 &  x902 &  x905 &  x908 &  x911 &  x917 &  x920 &  x923 &  x926 &  x929 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1097 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130 & ~x42 & ~x207 & ~x246 & ~x285 & ~x300 & ~x324 & ~x339 & ~x363 & ~x445 & ~x484;
assign c5278 =  x14 &  x41 &  x62 &  x65 &  x86 &  x92 &  x104 &  x107 &  x110 &  x113 &  x134 &  x164 &  x173 &  x185 &  x200 &  x215 &  x218 &  x227 &  x245 &  x269 &  x293 &  x320 &  x329 &  x353 &  x374 &  x377 &  x380 &  x401 &  x404 &  x410 &  x419 &  x422 &  x425 &  x436 &  x469 &  x473 &  x485 &  x497 &  x509 &  x542 &  x569 &  x575 &  x578 &  x596 &  x620 &  x623 &  x641 &  x680 &  x692 &  x707 &  x734 &  x745 &  x746 &  x773 &  x776 &  x806 &  x809 &  x821 &  x941 &  x973 &  x974 &  x980 &  x998 &  x1010 &  x1013 &  x1040 &  x1052 &  x1091 &  x1106 &  x1115 &  x1121 &  x1124 & ~x237 & ~x480 & ~x675;
assign c5280 =  x2 &  x11 &  x14 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x62 &  x65 &  x71 &  x74 &  x77 &  x79 &  x80 &  x83 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x118 &  x119 &  x122 &  x125 &  x131 &  x137 &  x140 &  x146 &  x149 &  x152 &  x155 &  x157 &  x158 &  x161 &  x164 &  x170 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x196 &  x197 &  x203 &  x206 &  x209 &  x215 &  x221 &  x224 &  x227 &  x230 &  x235 &  x242 &  x248 &  x257 &  x263 &  x266 &  x269 &  x274 &  x275 &  x278 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x314 &  x317 &  x320 &  x326 &  x329 &  x332 &  x335 &  x338 &  x344 &  x347 &  x350 &  x353 &  x355 &  x356 &  x359 &  x365 &  x371 &  x374 &  x377 &  x383 &  x386 &  x392 &  x394 &  x395 &  x398 &  x401 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x433 &  x437 &  x440 &  x443 &  x446 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x524 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x566 &  x569 &  x575 &  x578 &  x581 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x644 &  x647 &  x650 &  x653 &  x656 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x686 &  x689 &  x692 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x725 &  x728 &  x731 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x824 &  x827 &  x830 &  x836 &  x842 &  x845 &  x848 &  x854 &  x857 &  x860 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x893 &  x896 &  x899 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x953 &  x959 &  x962 &  x965 &  x968 &  x971 &  x977 &  x980 &  x983 &  x992 &  x995 &  x998 &  x1007 &  x1010 &  x1013 &  x1022 &  x1025 &  x1028 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1070 &  x1072 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x3 & ~x42 & ~x81 & ~x82 & ~x252 & ~x330 & ~x369 & ~x405 & ~x585 & ~x624 & ~x663 & ~x666 & ~x702 & ~x705;
assign c5282 =  x5 &  x65 &  x86 &  x110 &  x143 &  x173 &  x203 &  x278 &  x293 &  x296 &  x308 &  x326 &  x350 &  x374 &  x392 &  x395 &  x413 &  x449 &  x452 &  x482 &  x515 &  x527 &  x575 &  x581 &  x614 &  x647 &  x686 &  x719 &  x731 &  x737 &  x767 &  x797 &  x803 &  x827 &  x833 &  x842 &  x887 &  x893 &  x899 &  x944 &  x992 &  x1010 &  x1013 &  x1025 &  x1067 &  x1085 &  x1106 &  x1127 & ~x126 & ~x273 & ~x453 & ~x718 & ~x835 & ~x1041;
assign c5284 =  x5 &  x17 &  x20 &  x35 &  x41 &  x44 &  x46 &  x71 &  x74 &  x79 &  x85 &  x95 &  x119 &  x123 &  x140 &  x155 &  x158 &  x163 &  x164 &  x167 &  x170 &  x173 &  x176 &  x185 &  x203 &  x206 &  x233 &  x245 &  x269 &  x275 &  x278 &  x281 &  x284 &  x296 &  x299 &  x308 &  x317 &  x323 &  x329 &  x347 &  x350 &  x353 &  x362 &  x386 &  x389 &  x401 &  x407 &  x410 &  x416 &  x419 &  x437 &  x440 &  x455 &  x458 &  x467 &  x476 &  x500 &  x515 &  x530 &  x551 &  x554 &  x566 &  x569 &  x572 &  x587 &  x593 &  x599 &  x614 &  x620 &  x635 &  x638 &  x647 &  x650 &  x653 &  x656 &  x677 &  x680 &  x686 &  x710 &  x713 &  x722 &  x728 &  x734 &  x749 &  x755 &  x758 &  x767 &  x773 &  x782 &  x800 &  x809 &  x815 &  x818 &  x821 &  x824 &  x830 &  x850 &  x863 &  x866 &  x869 &  x872 &  x881 &  x884 &  x887 &  x893 &  x899 &  x905 &  x911 &  x923 &  x926 &  x932 &  x935 &  x953 &  x971 &  x974 &  x992 &  x998 &  x1004 &  x1007 &  x1019 &  x1034 &  x1037 &  x1049 &  x1058 &  x1073 &  x1076 &  x1079 &  x1088 &  x1118 &  x1121 & ~x159 & ~x264 & ~x819;
assign c5286 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x56 &  x59 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x122 &  x125 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x338 &  x341 &  x347 &  x350 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x542 &  x545 &  x548 &  x551 &  x557 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x656 &  x659 &  x662 &  x665 &  x668 &  x674 &  x677 &  x680 &  x686 &  x688 &  x689 &  x692 &  x695 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x727 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x773 &  x779 &  x782 &  x785 &  x788 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x838 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x893 &  x896 &  x899 &  x902 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x953 &  x956 &  x959 &  x962 &  x965 &  x971 &  x974 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x3 & ~x42 & ~x129 & ~x169 & ~x246 & ~x285 & ~x324 & ~x363 & ~x402 & ~x444 & ~x522 & ~x600 & ~x639 & ~x750;
assign c5288 =  x5 &  x11 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x59 &  x62 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x89 &  x92 &  x94 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x118 &  x119 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x145 &  x146 &  x149 &  x152 &  x155 &  x157 &  x161 &  x164 &  x170 &  x172 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x206 &  x209 &  x211 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x235 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x257 &  x263 &  x269 &  x274 &  x281 &  x284 &  x287 &  x289 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x344 &  x347 &  x350 &  x352 &  x353 &  x356 &  x365 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x391 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x443 &  x446 &  x452 &  x455 &  x458 &  x461 &  x464 &  x470 &  x473 &  x476 &  x479 &  x491 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x542 &  x545 &  x548 &  x551 &  x557 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x602 &  x605 &  x608 &  x614 &  x620 &  x623 &  x626 &  x629 &  x632 &  x638 &  x641 &  x644 &  x646 &  x647 &  x650 &  x653 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x737 &  x740 &  x743 &  x746 &  x755 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x812 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x854 &  x857 &  x860 &  x863 &  x866 &  x872 &  x878 &  x884 &  x887 &  x890 &  x896 &  x899 &  x902 &  x905 &  x908 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x120 & ~x159 & ~x198 & ~x363 & ~x402 & ~x403 & ~x441 & ~x480 & ~x519 & ~x597;
assign c5290 =  x2 &  x8 &  x14 &  x20 &  x26 &  x32 &  x33 &  x34 &  x40 &  x47 &  x59 &  x68 &  x71 &  x73 &  x74 &  x79 &  x83 &  x89 &  x112 &  x122 &  x125 &  x131 &  x137 &  x140 &  x143 &  x146 &  x151 &  x152 &  x157 &  x158 &  x161 &  x182 &  x188 &  x197 &  x206 &  x212 &  x215 &  x230 &  x235 &  x239 &  x251 &  x263 &  x266 &  x274 &  x284 &  x287 &  x296 &  x299 &  x326 &  x335 &  x338 &  x347 &  x353 &  x389 &  x395 &  x410 &  x413 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x452 &  x464 &  x467 &  x470 &  x473 &  x479 &  x488 &  x493 &  x494 &  x497 &  x503 &  x506 &  x515 &  x518 &  x524 &  x536 &  x542 &  x548 &  x551 &  x557 &  x560 &  x563 &  x566 &  x578 &  x581 &  x584 &  x587 &  x596 &  x602 &  x605 &  x608 &  x614 &  x622 &  x626 &  x629 &  x635 &  x638 &  x641 &  x649 &  x650 &  x665 &  x674 &  x677 &  x680 &  x685 &  x692 &  x695 &  x707 &  x710 &  x719 &  x722 &  x725 &  x734 &  x740 &  x743 &  x749 &  x755 &  x758 &  x770 &  x778 &  x785 &  x800 &  x809 &  x815 &  x817 &  x818 &  x821 &  x830 &  x833 &  x842 &  x845 &  x847 &  x851 &  x872 &  x875 &  x878 &  x884 &  x890 &  x893 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x938 &  x944 &  x947 &  x950 &  x971 &  x980 &  x989 &  x995 &  x998 &  x1004 &  x1007 &  x1013 &  x1028 &  x1034 &  x1037 &  x1040 &  x1055 &  x1064 &  x1070 &  x1076 &  x1079 &  x1085 &  x1088 &  x1096 &  x1100 &  x1103 &  x1112 &  x1118 &  x1127 & ~x285 & ~x324 & ~x666;
assign c5292 =  x0 &  x5 &  x14 &  x17 &  x34 &  x39 &  x41 &  x47 &  x67 &  x77 &  x83 &  x86 &  x98 &  x116 &  x119 &  x134 &  x137 &  x143 &  x149 &  x161 &  x176 &  x185 &  x191 &  x196 &  x206 &  x221 &  x230 &  x233 &  x242 &  x245 &  x248 &  x260 &  x269 &  x275 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x323 &  x341 &  x344 &  x353 &  x395 &  x401 &  x407 &  x425 &  x437 &  x446 &  x449 &  x461 &  x482 &  x530 &  x569 &  x578 &  x581 &  x590 &  x593 &  x617 &  x620 &  x623 &  x626 &  x710 &  x725 &  x740 &  x749 &  x758 &  x764 &  x769 &  x779 &  x782 &  x833 &  x839 &  x842 &  x869 &  x878 &  x890 &  x905 &  x917 &  x944 &  x950 &  x968 &  x986 &  x989 &  x992 &  x995 &  x997 &  x1006 &  x1016 &  x1018 &  x1052 &  x1061 &  x1076 &  x1096 &  x1106 &  x1112 & ~x438 & ~x672;
assign c5294 =  x5 &  x17 &  x38 &  x41 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x83 &  x86 &  x89 &  x101 &  x107 &  x119 &  x122 &  x125 &  x137 &  x149 &  x152 &  x164 &  x170 &  x176 &  x188 &  x194 &  x209 &  x212 &  x227 &  x233 &  x236 &  x251 &  x254 &  x257 &  x260 &  x272 &  x278 &  x287 &  x293 &  x302 &  x308 &  x311 &  x314 &  x317 &  x320 &  x326 &  x329 &  x338 &  x344 &  x356 &  x377 &  x380 &  x383 &  x401 &  x410 &  x413 &  x422 &  x425 &  x430 &  x443 &  x446 &  x452 &  x461 &  x469 &  x473 &  x482 &  x485 &  x491 &  x506 &  x518 &  x521 &  x524 &  x530 &  x533 &  x539 &  x545 &  x551 &  x557 &  x563 &  x566 &  x569 &  x575 &  x578 &  x587 &  x590 &  x593 &  x605 &  x611 &  x617 &  x623 &  x626 &  x628 &  x635 &  x656 &  x665 &  x667 &  x680 &  x686 &  x695 &  x710 &  x722 &  x728 &  x734 &  x737 &  x740 &  x746 &  x752 &  x755 &  x758 &  x767 &  x784 &  x821 &  x824 &  x827 &  x830 &  x839 &  x845 &  x851 &  x857 &  x862 &  x878 &  x881 &  x884 &  x887 &  x893 &  x901 &  x902 &  x911 &  x923 &  x935 &  x938 &  x959 &  x968 &  x971 &  x977 &  x980 &  x986 &  x989 &  x995 &  x1007 &  x1010 &  x1025 &  x1034 &  x1040 &  x1046 &  x1058 &  x1070 &  x1073 &  x1079 &  x1085 &  x1091 &  x1109 & ~x237 & ~x603 & ~x642 & ~x678 & ~x681;
assign c5296 =  x2 &  x5 &  x17 &  x20 &  x35 &  x38 &  x53 &  x65 &  x80 &  x86 &  x113 &  x116 &  x143 &  x155 &  x167 &  x170 &  x202 &  x212 &  x215 &  x218 &  x224 &  x245 &  x248 &  x257 &  x260 &  x269 &  x284 &  x319 &  x326 &  x329 &  x332 &  x344 &  x347 &  x353 &  x356 &  x362 &  x368 &  x371 &  x380 &  x392 &  x401 &  x410 &  x419 &  x431 &  x437 &  x440 &  x449 &  x455 &  x467 &  x485 &  x497 &  x506 &  x515 &  x524 &  x539 &  x545 &  x554 &  x572 &  x575 &  x581 &  x587 &  x590 &  x593 &  x599 &  x605 &  x623 &  x641 &  x653 &  x674 &  x689 &  x692 &  x701 &  x710 &  x728 &  x734 &  x740 &  x749 &  x773 &  x776 &  x779 &  x800 &  x812 &  x815 &  x818 &  x824 &  x830 &  x833 &  x845 &  x857 &  x860 &  x863 &  x866 &  x869 &  x881 &  x884 &  x887 &  x899 &  x929 &  x932 &  x935 &  x941 &  x947 &  x950 &  x956 &  x962 &  x974 &  x995 &  x998 &  x1001 &  x1004 &  x1018 &  x1025 &  x1031 &  x1040 &  x1046 &  x1049 &  x1082 &  x1106 &  x1118 &  x1121 & ~x237 & ~x291 & ~x316 & ~x636 & ~x675 & ~x714;
assign c5298 =  x5 &  x8 &  x14 &  x35 &  x47 &  x53 &  x59 &  x62 &  x80 &  x89 &  x110 &  x116 &  x122 &  x134 &  x137 &  x155 &  x170 &  x188 &  x194 &  x200 &  x203 &  x215 &  x224 &  x242 &  x245 &  x272 &  x275 &  x296 &  x305 &  x311 &  x335 &  x341 &  x347 &  x371 &  x380 &  x389 &  x395 &  x404 &  x413 &  x416 &  x431 &  x446 &  x482 &  x488 &  x500 &  x515 &  x533 &  x551 &  x557 &  x560 &  x572 &  x578 &  x581 &  x584 &  x590 &  x596 &  x605 &  x635 &  x656 &  x659 &  x686 &  x695 &  x698 &  x722 &  x728 &  x731 &  x742 &  x749 &  x776 &  x779 &  x794 &  x797 &  x806 &  x818 &  x827 &  x854 &  x860 &  x866 &  x875 &  x878 &  x881 &  x896 &  x908 &  x911 &  x938 &  x939 &  x941 &  x947 &  x953 &  x979 &  x1004 &  x1013 &  x1028 &  x1043 &  x1046 &  x1058 &  x1076 &  x1079 &  x1088 &  x1091 &  x1094 &  x1112 &  x1130 & ~x234 & ~x312 & ~x351 & ~x471 & ~x511 & ~x621 & ~x792 & ~x831 & ~x837;
assign c51 =  x50 &  x56 &  x170 &  x308 &  x632 &  x683 &  x746 &  x770 &  x845 &  x1052 & ~x505 & ~x1050;
assign c53 =  x20 &  x29 &  x35 &  x38 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x74 &  x77 &  x80 &  x89 &  x104 &  x110 &  x122 &  x128 &  x134 &  x161 &  x170 &  x175 &  x179 &  x181 &  x182 &  x188 &  x191 &  x203 &  x212 &  x215 &  x224 &  x227 &  x239 &  x272 &  x281 &  x287 &  x290 &  x299 &  x302 &  x314 &  x317 &  x323 &  x332 &  x335 &  x341 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x386 &  x392 &  x394 &  x401 &  x404 &  x413 &  x419 &  x422 &  x430 &  x433 &  x437 &  x443 &  x449 &  x452 &  x469 &  x470 &  x472 &  x479 &  x485 &  x500 &  x503 &  x508 &  x518 &  x521 &  x524 &  x533 &  x536 &  x542 &  x545 &  x554 &  x557 &  x566 &  x572 &  x575 &  x578 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x614 &  x623 &  x626 &  x629 &  x632 &  x641 &  x653 &  x671 &  x674 &  x680 &  x683 &  x686 &  x695 &  x707 &  x716 &  x719 &  x722 &  x734 &  x737 &  x749 &  x755 &  x764 &  x770 &  x773 &  x776 &  x797 &  x803 &  x806 &  x851 &  x860 &  x863 &  x872 &  x878 &  x881 &  x899 &  x908 &  x914 &  x923 &  x929 &  x932 &  x938 &  x947 &  x974 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1016 &  x1025 &  x1040 &  x1046 &  x1052 &  x1058 &  x1061 &  x1064 &  x1070 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x195 & ~x513;
assign c55 =  x4 &  x23 &  x50 &  x59 &  x95 &  x128 &  x152 &  x199 &  x272 &  x308 &  x341 &  x344 &  x347 &  x353 &  x404 &  x443 &  x452 &  x485 &  x494 &  x563 &  x566 &  x587 &  x641 &  x647 &  x671 &  x677 &  x701 &  x740 &  x757 &  x761 &  x782 &  x881 &  x932 &  x938 &  x968 &  x1013 &  x1055 &  x1064 &  x1091 &  x1121 & ~x642 & ~x900;
assign c57 =  x20 &  x47 &  x158 &  x188 &  x206 &  x218 &  x236 &  x308 &  x326 &  x353 &  x398 &  x410 &  x449 &  x461 &  x515 &  x566 &  x569 &  x578 &  x599 &  x629 &  x658 &  x668 &  x686 &  x719 &  x782 &  x791 &  x962 &  x974 &  x992 &  x1007 &  x1115 &  x1130 & ~x264 & ~x822 & ~x862 & ~x1095;
assign c59 =  x5 &  x14 &  x20 &  x29 &  x41 &  x44 &  x56 &  x65 &  x68 &  x77 &  x80 &  x83 &  x98 &  x101 &  x104 &  x113 &  x121 &  x122 &  x125 &  x128 &  x131 &  x137 &  x140 &  x143 &  x152 &  x158 &  x170 &  x173 &  x194 &  x196 &  x199 &  x203 &  x209 &  x215 &  x218 &  x224 &  x227 &  x235 &  x236 &  x248 &  x251 &  x254 &  x257 &  x260 &  x266 &  x269 &  x274 &  x284 &  x287 &  x290 &  x299 &  x320 &  x323 &  x329 &  x332 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x374 &  x383 &  x395 &  x398 &  x404 &  x413 &  x422 &  x425 &  x428 &  x431 &  x440 &  x443 &  x446 &  x449 &  x455 &  x458 &  x461 &  x464 &  x470 &  x473 &  x476 &  x482 &  x491 &  x497 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x527 &  x533 &  x536 &  x545 &  x548 &  x560 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x587 &  x593 &  x599 &  x602 &  x605 &  x608 &  x617 &  x626 &  x635 &  x638 &  x644 &  x647 &  x653 &  x665 &  x668 &  x671 &  x674 &  x680 &  x686 &  x701 &  x704 &  x707 &  x710 &  x713 &  x719 &  x722 &  x731 &  x740 &  x746 &  x749 &  x752 &  x760 &  x764 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x818 &  x827 &  x830 &  x839 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x875 &  x878 &  x887 &  x893 &  x899 &  x902 &  x908 &  x914 &  x917 &  x926 &  x944 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1022 &  x1025 &  x1028 &  x1037 &  x1052 &  x1055 &  x1064 &  x1076 &  x1079 &  x1085 &  x1088 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x330 & ~x663 & ~x912 & ~x951;
assign c511 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x29 &  x32 &  x35 &  x41 &  x44 &  x50 &  x53 &  x59 &  x65 &  x74 &  x77 &  x86 &  x89 &  x98 &  x101 &  x110 &  x116 &  x125 &  x131 &  x140 &  x143 &  x146 &  x155 &  x158 &  x170 &  x176 &  x179 &  x182 &  x185 &  x191 &  x197 &  x200 &  x206 &  x208 &  x212 &  x215 &  x218 &  x227 &  x233 &  x236 &  x239 &  x247 &  x248 &  x254 &  x260 &  x266 &  x269 &  x272 &  x281 &  x296 &  x299 &  x308 &  x317 &  x332 &  x344 &  x350 &  x359 &  x371 &  x380 &  x383 &  x386 &  x395 &  x401 &  x413 &  x419 &  x422 &  x431 &  x434 &  x437 &  x446 &  x449 &  x452 &  x455 &  x461 &  x464 &  x467 &  x476 &  x482 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x509 &  x512 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x560 &  x563 &  x566 &  x575 &  x581 &  x587 &  x593 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x656 &  x659 &  x662 &  x671 &  x674 &  x677 &  x683 &  x686 &  x692 &  x695 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x740 &  x743 &  x752 &  x761 &  x764 &  x767 &  x770 &  x773 &  x779 &  x782 &  x790 &  x794 &  x797 &  x800 &  x803 &  x809 &  x824 &  x827 &  x830 &  x833 &  x835 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x869 &  x872 &  x875 &  x881 &  x887 &  x896 &  x899 &  x908 &  x911 &  x932 &  x935 &  x944 &  x950 &  x953 &  x956 &  x974 &  x989 &  x992 &  x995 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1040 &  x1043 &  x1049 &  x1055 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1082 &  x1085 &  x1088 &  x1091 &  x1106 &  x1109 &  x1115 &  x1118 &  x1127 & ~x201 & ~x240;
assign c513 =  x170 &  x205 &  x293 &  x335 &  x424 &  x434 &  x560 &  x593 &  x608 &  x721 &  x740 &  x746 &  x872 &  x1001 &  x1004 & ~x381 & ~x459 & ~x471 & ~x666 & ~x705;
assign c515 =  x11 &  x43 &  x47 &  x71 &  x82 &  x101 &  x122 &  x125 &  x131 &  x143 &  x155 &  x164 &  x170 &  x176 &  x185 &  x188 &  x191 &  x194 &  x199 &  x200 &  x203 &  x206 &  x209 &  x221 &  x227 &  x233 &  x245 &  x263 &  x269 &  x272 &  x275 &  x281 &  x287 &  x290 &  x308 &  x314 &  x329 &  x335 &  x338 &  x344 &  x350 &  x353 &  x356 &  x368 &  x374 &  x389 &  x392 &  x395 &  x410 &  x413 &  x419 &  x440 &  x461 &  x515 &  x527 &  x530 &  x536 &  x539 &  x560 &  x563 &  x569 &  x572 &  x575 &  x587 &  x608 &  x611 &  x617 &  x632 &  x644 &  x653 &  x662 &  x665 &  x668 &  x674 &  x686 &  x695 &  x707 &  x710 &  x719 &  x728 &  x734 &  x737 &  x740 &  x755 &  x788 &  x791 &  x799 &  x806 &  x812 &  x821 &  x827 &  x830 &  x848 &  x857 &  x869 &  x872 &  x875 &  x887 &  x899 &  x916 &  x917 &  x926 &  x935 &  x941 &  x944 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x980 &  x995 &  x998 &  x1001 &  x1004 &  x1006 &  x1019 &  x1028 &  x1037 &  x1043 &  x1045 &  x1049 &  x1052 &  x1055 &  x1058 &  x1073 &  x1094 &  x1121 &  x1124 &  x1130 & ~x705 & ~x822;
assign c517 =  x11 &  x13 &  x32 &  x71 &  x164 &  x199 &  x203 &  x254 &  x404 &  x407 &  x452 &  x461 &  x491 &  x575 &  x581 &  x605 &  x632 &  x748 &  x755 &  x845 &  x872 &  x929 & ~x72 & ~x858 & ~x1092;
assign c519 =  x19 &  x31 &  x125 &  x470 &  x500 &  x572 &  x720 &  x914 &  x1010 & ~x333;
assign c521 =  x32 &  x170 &  x272 &  x403 &  x409 &  x581 &  x628 &  x713 &  x946 &  x1001 & ~x165 & ~x282;
assign c523 =  x26 &  x88 &  x161 &  x173 &  x283 &  x409 &  x415 &  x448 &  x467 &  x473 &  x557 &  x559 &  x598 &  x623 &  x668 &  x671 &  x706 &  x764 &  x806 &  x839 &  x842 &  x929 &  x1025 & ~x468;
assign c525 =  x5 &  x53 &  x59 &  x68 &  x74 &  x77 &  x83 &  x86 &  x101 &  x155 &  x164 &  x185 &  x188 &  x206 &  x221 &  x233 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x263 &  x265 &  x269 &  x272 &  x314 &  x323 &  x338 &  x344 &  x350 &  x353 &  x359 &  x365 &  x380 &  x395 &  x401 &  x404 &  x410 &  x413 &  x419 &  x428 &  x437 &  x440 &  x446 &  x452 &  x470 &  x473 &  x476 &  x482 &  x512 &  x521 &  x530 &  x545 &  x557 &  x569 &  x584 &  x608 &  x620 &  x629 &  x632 &  x635 &  x653 &  x662 &  x686 &  x701 &  x707 &  x752 &  x764 &  x773 &  x776 &  x785 &  x800 &  x812 &  x821 &  x827 &  x845 &  x848 &  x854 &  x857 &  x860 &  x863 &  x866 &  x878 &  x890 &  x896 &  x905 &  x913 &  x917 &  x920 &  x923 &  x941 &  x944 &  x989 &  x998 &  x1001 &  x1019 &  x1037 &  x1043 &  x1049 &  x1064 &  x1103 &  x1112 &  x1115 & ~x372 & ~x606 & ~x1095;
assign c527 =  x5 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x44 &  x50 &  x53 &  x56 &  x62 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x101 &  x104 &  x110 &  x113 &  x119 &  x122 &  x125 &  x131 &  x134 &  x137 &  x140 &  x143 &  x154 &  x155 &  x164 &  x167 &  x170 &  x176 &  x179 &  x184 &  x187 &  x188 &  x191 &  x194 &  x197 &  x200 &  x206 &  x209 &  x220 &  x221 &  x223 &  x227 &  x233 &  x236 &  x242 &  x245 &  x248 &  x251 &  x259 &  x260 &  x263 &  x266 &  x269 &  x272 &  x290 &  x293 &  x296 &  x298 &  x302 &  x314 &  x317 &  x320 &  x323 &  x329 &  x335 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x374 &  x383 &  x386 &  x389 &  x392 &  x395 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x437 &  x440 &  x452 &  x455 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x506 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x542 &  x545 &  x551 &  x557 &  x560 &  x563 &  x566 &  x569 &  x581 &  x584 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x644 &  x647 &  x650 &  x653 &  x659 &  x662 &  x665 &  x668 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x701 &  x707 &  x713 &  x728 &  x734 &  x737 &  x740 &  x749 &  x752 &  x758 &  x770 &  x773 &  x788 &  x797 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x842 &  x851 &  x854 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x884 &  x887 &  x890 &  x896 &  x902 &  x905 &  x908 &  x911 &  x917 &  x920 &  x923 &  x926 &  x935 &  x941 &  x944 &  x950 &  x953 &  x956 &  x965 &  x968 &  x971 &  x974 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1022 &  x1025 &  x1028 &  x1034 &  x1037 &  x1040 &  x1046 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1109 &  x1115 &  x1121 &  x1130 & ~x120 & ~x195 & ~x198 & ~x273 & ~x522;
assign c529 =  x5 &  x23 &  x25 &  x44 &  x64 &  x71 &  x101 &  x107 &  x146 &  x155 &  x173 &  x179 &  x254 &  x311 &  x316 &  x326 &  x332 &  x355 &  x392 &  x404 &  x433 &  x524 &  x554 &  x569 &  x605 &  x650 &  x656 &  x659 &  x665 &  x713 &  x734 &  x806 &  x839 &  x872 &  x929 &  x932 &  x959 &  x965 &  x995 &  x1004 &  x1007 &  x1088 & ~x54 & ~x897;
assign c531 =  x64 &  x113 &  x355 &  x419 &  x446 &  x683 &  x800 &  x821 &  x953 &  x1007 &  x1031 &  x1094 & ~x0 & ~x40 & ~x93;
assign c533 =  x5 &  x23 &  x32 &  x35 &  x50 &  x53 &  x71 &  x92 &  x101 &  x125 &  x128 &  x131 &  x170 &  x173 &  x212 &  x245 &  x269 &  x272 &  x277 &  x290 &  x296 &  x314 &  x332 &  x335 &  x356 &  x374 &  x391 &  x413 &  x416 &  x443 &  x473 &  x476 &  x488 &  x491 &  x509 &  x527 &  x536 &  x560 &  x586 &  x590 &  x596 &  x599 &  x614 &  x620 &  x656 &  x713 &  x722 &  x737 &  x755 &  x845 &  x857 &  x860 &  x869 &  x872 &  x938 &  x968 &  x980 &  x1007 &  x1031 &  x1076 &  x1082 &  x1088 &  x1097 &  x1103 &  x1124 &  x1130 & ~x111 & ~x474;
assign c535 =  x2 &  x8 &  x14 &  x35 &  x44 &  x47 &  x50 &  x53 &  x68 &  x71 &  x74 &  x83 &  x86 &  x89 &  x95 &  x101 &  x122 &  x140 &  x143 &  x179 &  x191 &  x197 &  x203 &  x206 &  x209 &  x224 &  x230 &  x233 &  x254 &  x260 &  x266 &  x296 &  x320 &  x323 &  x326 &  x329 &  x332 &  x356 &  x365 &  x370 &  x374 &  x377 &  x389 &  x392 &  x403 &  x407 &  x409 &  x413 &  x415 &  x425 &  x428 &  x431 &  x446 &  x448 &  x449 &  x458 &  x473 &  x479 &  x482 &  x487 &  x512 &  x521 &  x533 &  x542 &  x545 &  x551 &  x560 &  x575 &  x581 &  x614 &  x626 &  x644 &  x659 &  x665 &  x674 &  x689 &  x706 &  x710 &  x725 &  x737 &  x743 &  x746 &  x752 &  x755 &  x758 &  x776 &  x788 &  x797 &  x800 &  x806 &  x809 &  x833 &  x848 &  x854 &  x869 &  x881 &  x887 &  x890 &  x893 &  x899 &  x905 &  x908 &  x911 &  x920 &  x932 &  x950 &  x971 &  x983 &  x986 &  x1001 &  x1010 &  x1016 &  x1022 &  x1034 &  x1037 &  x1061 &  x1085 &  x1100 &  x1109 &  x1118 &  x1127 &  x1130 & ~x843 & ~x960 & ~x1071;
assign c537 =  x8 &  x50 &  x82 &  x89 &  x95 &  x110 &  x131 &  x149 &  x170 &  x197 &  x203 &  x299 &  x302 &  x338 &  x395 &  x446 &  x479 &  x506 &  x509 &  x563 &  x641 &  x722 &  x737 &  x743 &  x752 &  x776 &  x791 &  x797 &  x811 &  x830 &  x845 &  x878 &  x941 &  x989 &  x995 &  x1004 &  x1007 &  x1040 &  x1051 &  x1084 &  x1106 &  x1121 &  x1123 & ~x306 & ~x858;
assign c539 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x278 &  x281 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x317 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x392 &  x395 &  x398 &  x400 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x442 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x509 &  x512 &  x515 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x626 &  x628 &  x629 &  x632 &  x635 &  x638 &  x644 &  x647 &  x650 &  x653 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x703 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x725 &  x728 &  x731 &  x734 &  x737 &  x742 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x806 &  x809 &  x812 &  x815 &  x818 &  x820 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x859 &  x863 &  x866 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x898 &  x899 &  x902 &  x908 &  x911 &  x917 &  x920 &  x926 &  x932 &  x935 &  x937 &  x938 &  x941 &  x944 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x976 &  x977 &  x980 &  x983 &  x986 &  x989 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1088 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1124 & ~x273 & ~x312 & ~x351;
assign c541 =  x89 &  x101 &  x212 &  x227 &  x236 &  x337 &  x359 &  x380 &  x389 &  x425 &  x452 &  x524 &  x542 &  x638 &  x827 &  x848 &  x875 &  x944 &  x1034 &  x1097 &  x1109 &  x1121 & ~x513 & ~x670 & ~x855 & ~x894;
assign c543 =  x5 &  x8 &  x11 &  x16 &  x59 &  x62 &  x74 &  x106 &  x119 &  x128 &  x131 &  x144 &  x152 &  x167 &  x176 &  x179 &  x188 &  x190 &  x194 &  x269 &  x299 &  x305 &  x326 &  x335 &  x347 &  x383 &  x403 &  x431 &  x437 &  x449 &  x464 &  x494 &  x500 &  x521 &  x533 &  x554 &  x557 &  x598 &  x605 &  x623 &  x626 &  x674 &  x695 &  x725 &  x737 &  x743 &  x752 &  x779 &  x788 &  x800 &  x821 &  x839 &  x869 &  x875 &  x878 &  x887 &  x896 &  x898 &  x908 &  x911 &  x923 &  x941 &  x971 &  x1001 &  x1046 &  x1055 &  x1058 &  x1076 &  x1079 &  x1112 &  x1127 & ~x51 & ~x90;
assign c545 =  x92 &  x367 & ~x687 & ~x901;
assign c547 =  x1 &  x2 &  x4 &  x8 &  x23 &  x40 &  x41 &  x53 &  x56 &  x68 &  x77 &  x79 &  x92 &  x113 &  x137 &  x152 &  x179 &  x196 &  x218 &  x221 &  x233 &  x242 &  x245 &  x266 &  x275 &  x284 &  x290 &  x299 &  x305 &  x320 &  x329 &  x332 &  x347 &  x356 &  x365 &  x389 &  x395 &  x404 &  x407 &  x410 &  x416 &  x419 &  x425 &  x449 &  x458 &  x467 &  x470 &  x488 &  x497 &  x503 &  x509 &  x512 &  x560 &  x566 &  x572 &  x587 &  x599 &  x605 &  x608 &  x620 &  x632 &  x638 &  x641 &  x647 &  x653 &  x659 &  x665 &  x668 &  x674 &  x677 &  x680 &  x689 &  x704 &  x710 &  x713 &  x716 &  x721 &  x722 &  x728 &  x743 &  x758 &  x761 &  x764 &  x767 &  x782 &  x785 &  x791 &  x800 &  x803 &  x806 &  x824 &  x833 &  x845 &  x857 &  x860 &  x863 &  x872 &  x875 &  x878 &  x887 &  x896 &  x911 &  x914 &  x917 &  x923 &  x929 &  x932 &  x944 &  x950 &  x953 &  x956 &  x974 &  x998 &  x1010 &  x1013 &  x1025 &  x1031 &  x1046 &  x1067 &  x1070 &  x1079 &  x1091 &  x1094 &  x1106 &  x1109 &  x1112 &  x1127 &  x1130 & ~x45 & ~x123 & ~x822 & ~x1059 & ~x1098;
assign c549 =  x17 &  x20 &  x29 &  x32 &  x35 &  x53 &  x56 &  x65 &  x82 &  x83 &  x92 &  x113 &  x119 &  x121 &  x122 &  x125 &  x134 &  x140 &  x149 &  x176 &  x179 &  x197 &  x199 &  x200 &  x218 &  x221 &  x227 &  x230 &  x235 &  x245 &  x251 &  x263 &  x266 &  x278 &  x287 &  x290 &  x314 &  x329 &  x338 &  x344 &  x347 &  x350 &  x359 &  x368 &  x374 &  x377 &  x380 &  x383 &  x386 &  x398 &  x407 &  x410 &  x428 &  x452 &  x461 &  x464 &  x479 &  x491 &  x497 &  x515 &  x521 &  x527 &  x530 &  x545 &  x560 &  x584 &  x593 &  x608 &  x614 &  x617 &  x629 &  x632 &  x635 &  x647 &  x650 &  x653 &  x668 &  x677 &  x692 &  x698 &  x701 &  x704 &  x716 &  x719 &  x722 &  x728 &  x731 &  x767 &  x773 &  x800 &  x803 &  x812 &  x818 &  x821 &  x854 &  x875 &  x878 &  x887 &  x899 &  x905 &  x908 &  x911 &  x914 &  x926 &  x929 &  x959 &  x968 &  x986 &  x992 &  x1013 &  x1019 &  x1025 &  x1034 &  x1037 &  x1043 &  x1052 &  x1055 &  x1058 &  x1082 &  x1088 &  x1118 &  x1121 &  x1124 &  x1130 & ~x264 & ~x303 & ~x783 & ~x1017;
assign c551 =  x35 &  x68 &  x95 &  x98 &  x118 &  x134 &  x137 &  x146 &  x194 &  x230 &  x274 &  x293 &  x299 &  x302 &  x305 &  x346 &  x395 &  x398 &  x431 &  x461 &  x479 &  x491 &  x503 &  x524 &  x542 &  x575 &  x584 &  x641 &  x671 &  x695 &  x704 &  x731 &  x743 &  x797 &  x803 &  x854 &  x869 &  x878 &  x919 &  x929 &  x941 &  x947 &  x958 &  x965 &  x968 &  x989 &  x997 &  x1061 &  x1088 &  x1103 & ~x627 & ~x666 & ~x669 & ~x708 & ~x744 & ~x1083;
assign c553 =  x2 &  x5 &  x8 &  x20 &  x23 &  x32 &  x35 &  x41 &  x44 &  x47 &  x50 &  x56 &  x62 &  x71 &  x77 &  x80 &  x83 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x131 &  x134 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x161 &  x164 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x212 &  x215 &  x221 &  x227 &  x230 &  x233 &  x236 &  x242 &  x245 &  x248 &  x254 &  x257 &  x260 &  x263 &  x266 &  x272 &  x278 &  x281 &  x290 &  x293 &  x305 &  x308 &  x311 &  x320 &  x326 &  x332 &  x335 &  x341 &  x344 &  x359 &  x362 &  x365 &  x371 &  x374 &  x383 &  x386 &  x392 &  x395 &  x398 &  x401 &  x404 &  x410 &  x413 &  x425 &  x428 &  x434 &  x440 &  x443 &  x455 &  x458 &  x461 &  x467 &  x470 &  x476 &  x479 &  x482 &  x488 &  x491 &  x494 &  x503 &  x518 &  x524 &  x527 &  x530 &  x533 &  x545 &  x548 &  x554 &  x563 &  x572 &  x575 &  x584 &  x587 &  x590 &  x599 &  x605 &  x608 &  x611 &  x620 &  x626 &  x629 &  x632 &  x638 &  x644 &  x647 &  x650 &  x656 &  x662 &  x664 &  x665 &  x668 &  x671 &  x674 &  x683 &  x689 &  x695 &  x698 &  x703 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x728 &  x734 &  x737 &  x740 &  x746 &  x749 &  x758 &  x761 &  x764 &  x767 &  x770 &  x781 &  x785 &  x797 &  x803 &  x806 &  x820 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x842 &  x845 &  x848 &  x859 &  x860 &  x863 &  x866 &  x869 &  x881 &  x893 &  x896 &  x898 &  x911 &  x914 &  x932 &  x935 &  x937 &  x941 &  x947 &  x950 &  x953 &  x962 &  x965 &  x968 &  x971 &  x974 &  x976 &  x977 &  x983 &  x989 &  x992 &  x995 &  x1007 &  x1010 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1052 &  x1055 &  x1058 &  x1061 &  x1076 &  x1079 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1124 &  x1127 & ~x426 & ~x513 & ~x801 & ~x879;
assign c555 =  x17 &  x77 &  x80 &  x83 &  x134 &  x140 &  x233 &  x236 &  x242 &  x248 &  x272 &  x284 &  x296 &  x298 &  x329 &  x374 &  x389 &  x416 &  x434 &  x442 &  x506 &  x515 &  x536 &  x563 &  x628 &  x641 &  x703 &  x737 &  x755 &  x776 &  x781 &  x791 &  x820 &  x823 &  x830 &  x866 &  x898 &  x905 &  x911 &  x946 &  x962 &  x985 &  x986 &  x1019 &  x1028 &  x1031 &  x1058 &  x1076 &  x1094 &  x1130;
assign c557 =  x2 &  x5 &  x44 &  x71 &  x92 &  x95 &  x110 &  x125 &  x131 &  x143 &  x161 &  x170 &  x188 &  x194 &  x212 &  x218 &  x245 &  x269 &  x275 &  x284 &  x299 &  x314 &  x323 &  x337 &  x356 &  x362 &  x386 &  x398 &  x407 &  x415 &  x422 &  x425 &  x455 &  x470 &  x503 &  x560 &  x569 &  x584 &  x587 &  x623 &  x635 &  x677 &  x698 &  x701 &  x706 &  x719 &  x725 &  x743 &  x749 &  x752 &  x770 &  x773 &  x785 &  x791 &  x809 &  x821 &  x842 &  x845 &  x857 &  x869 &  x887 &  x890 &  x917 &  x920 &  x935 &  x950 &  x965 &  x968 &  x971 &  x992 &  x1010 &  x1019 &  x1022 &  x1049 &  x1061 &  x1064 &  x1067 &  x1100 &  x1103 &  x1109 &  x1118 &  x1124 &  x1127 & ~x312 & ~x961 & ~x999 & ~x1077;
assign c559 =  x137 &  x275 &  x299 &  x332 &  x389 &  x605 &  x698 &  x706 &  x932 &  x941 &  x995 &  x1004 &  x1082 &  x1088 &  x1130 & ~x468 & ~x922 & ~x1038;
assign c561 =  x5 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x32 &  x41 &  x53 &  x56 &  x68 &  x71 &  x82 &  x86 &  x89 &  x92 &  x98 &  x107 &  x122 &  x125 &  x128 &  x137 &  x143 &  x146 &  x149 &  x167 &  x170 &  x173 &  x176 &  x179 &  x191 &  x197 &  x206 &  x209 &  x215 &  x221 &  x227 &  x236 &  x242 &  x245 &  x263 &  x275 &  x278 &  x281 &  x311 &  x320 &  x338 &  x347 &  x356 &  x359 &  x374 &  x377 &  x380 &  x383 &  x386 &  x398 &  x401 &  x404 &  x413 &  x416 &  x419 &  x422 &  x431 &  x434 &  x437 &  x449 &  x452 &  x467 &  x476 &  x491 &  x503 &  x512 &  x515 &  x527 &  x545 &  x548 &  x554 &  x557 &  x563 &  x595 &  x614 &  x617 &  x623 &  x629 &  x632 &  x635 &  x641 &  x650 &  x653 &  x662 &  x668 &  x671 &  x679 &  x683 &  x686 &  x689 &  x695 &  x704 &  x707 &  x722 &  x725 &  x737 &  x746 &  x767 &  x770 &  x782 &  x788 &  x791 &  x794 &  x800 &  x803 &  x809 &  x815 &  x830 &  x833 &  x836 &  x860 &  x863 &  x881 &  x884 &  x893 &  x896 &  x899 &  x917 &  x920 &  x926 &  x941 &  x950 &  x956 &  x983 &  x986 &  x989 &  x998 &  x1001 &  x1010 &  x1013 &  x1019 &  x1022 &  x1034 &  x1037 &  x1043 &  x1052 &  x1055 &  x1058 &  x1073 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1118 &  x1121 &  x1127 &  x1130 & ~x303 & ~x666 & ~x822;
assign c563 =  x5 &  x8 &  x11 &  x14 &  x17 &  x32 &  x41 &  x44 &  x47 &  x53 &  x62 &  x68 &  x74 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x107 &  x110 &  x113 &  x116 &  x137 &  x143 &  x149 &  x167 &  x173 &  x176 &  x182 &  x188 &  x191 &  x194 &  x209 &  x212 &  x221 &  x233 &  x236 &  x242 &  x248 &  x251 &  x260 &  x266 &  x275 &  x278 &  x281 &  x284 &  x287 &  x296 &  x299 &  x308 &  x314 &  x325 &  x326 &  x335 &  x338 &  x341 &  x344 &  x353 &  x359 &  x362 &  x368 &  x371 &  x374 &  x383 &  x386 &  x389 &  x392 &  x395 &  x401 &  x413 &  x416 &  x425 &  x428 &  x434 &  x437 &  x449 &  x455 &  x458 &  x467 &  x470 &  x476 &  x479 &  x482 &  x485 &  x491 &  x506 &  x509 &  x512 &  x530 &  x545 &  x551 &  x554 &  x569 &  x572 &  x575 &  x581 &  x584 &  x587 &  x589 &  x596 &  x599 &  x608 &  x611 &  x617 &  x620 &  x623 &  x641 &  x647 &  x656 &  x659 &  x668 &  x677 &  x680 &  x683 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x713 &  x725 &  x728 &  x731 &  x737 &  x749 &  x752 &  x761 &  x767 &  x785 &  x800 &  x803 &  x806 &  x809 &  x812 &  x827 &  x830 &  x842 &  x845 &  x851 &  x854 &  x860 &  x866 &  x869 &  x872 &  x878 &  x881 &  x887 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x917 &  x941 &  x944 &  x950 &  x962 &  x968 &  x971 &  x974 &  x980 &  x983 &  x986 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1037 &  x1040 &  x1046 &  x1055 &  x1058 &  x1064 &  x1067 &  x1073 &  x1097 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1124 &  x1130 & ~x39 & ~x42 & ~x81 & ~x159 & ~x195 & ~x276 & ~x306;
assign c565 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x44 &  x50 &  x56 &  x59 &  x62 &  x68 &  x74 &  x77 &  x86 &  x89 &  x92 &  x98 &  x101 &  x107 &  x113 &  x116 &  x119 &  x122 &  x125 &  x131 &  x134 &  x137 &  x140 &  x143 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x176 &  x179 &  x182 &  x185 &  x191 &  x197 &  x200 &  x203 &  x206 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x347 &  x350 &  x353 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x419 &  x422 &  x425 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x458 &  x464 &  x467 &  x470 &  x478 &  x479 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x545 &  x551 &  x554 &  x557 &  x560 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x589 &  x590 &  x596 &  x599 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x625 &  x626 &  x628 &  x629 &  x632 &  x635 &  x638 &  x644 &  x647 &  x656 &  x659 &  x664 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x703 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x734 &  x737 &  x740 &  x742 &  x746 &  x749 &  x752 &  x758 &  x761 &  x764 &  x770 &  x776 &  x779 &  x781 &  x782 &  x788 &  x791 &  x794 &  x797 &  x806 &  x818 &  x820 &  x824 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x854 &  x859 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x898 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x923 &  x926 &  x929 &  x932 &  x935 &  x937 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x962 &  x965 &  x971 &  x974 &  x976 &  x977 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1007 &  x1010 &  x1013 &  x1015 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1054 &  x1061 &  x1064 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x687 & ~x726 & ~x765;
assign c567 =  x2 &  x5 &  x8 &  x14 &  x17 &  x23 &  x26 &  x32 &  x35 &  x41 &  x47 &  x50 &  x59 &  x62 &  x68 &  x83 &  x86 &  x95 &  x101 &  x107 &  x119 &  x121 &  x122 &  x125 &  x131 &  x134 &  x140 &  x149 &  x152 &  x158 &  x160 &  x170 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x203 &  x206 &  x212 &  x215 &  x218 &  x224 &  x227 &  x236 &  x238 &  x245 &  x254 &  x260 &  x275 &  x281 &  x287 &  x293 &  x296 &  x302 &  x305 &  x308 &  x311 &  x326 &  x329 &  x338 &  x344 &  x347 &  x350 &  x356 &  x359 &  x365 &  x368 &  x377 &  x380 &  x386 &  x398 &  x404 &  x407 &  x413 &  x416 &  x425 &  x434 &  x437 &  x449 &  x455 &  x458 &  x461 &  x467 &  x470 &  x473 &  x476 &  x482 &  x485 &  x488 &  x497 &  x500 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x548 &  x554 &  x557 &  x563 &  x566 &  x569 &  x575 &  x581 &  x584 &  x590 &  x593 &  x614 &  x617 &  x623 &  x626 &  x629 &  x632 &  x635 &  x641 &  x644 &  x653 &  x656 &  x659 &  x665 &  x668 &  x674 &  x680 &  x683 &  x686 &  x689 &  x695 &  x698 &  x707 &  x710 &  x716 &  x719 &  x722 &  x728 &  x737 &  x743 &  x746 &  x749 &  x755 &  x757 &  x764 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x806 &  x809 &  x812 &  x818 &  x821 &  x824 &  x839 &  x845 &  x851 &  x854 &  x860 &  x863 &  x866 &  x869 &  x872 &  x878 &  x881 &  x884 &  x887 &  x902 &  x905 &  x908 &  x911 &  x914 &  x920 &  x923 &  x926 &  x929 &  x938 &  x941 &  x944 &  x959 &  x965 &  x974 &  x980 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1013 &  x1019 &  x1025 &  x1028 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1055 &  x1058 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1127 &  x1130 & ~x258 & ~x375 & ~x822 & ~x861 & ~x900 & ~x939;
assign c569 =  x13 &  x383 &  x597 &  x799 & ~x984;
assign c571 =  x43 &  x56 &  x82 &  x137 &  x143 &  x199 &  x311 &  x320 &  x365 &  x401 &  x410 &  x455 &  x467 &  x631 &  x835 & ~x414;
assign c573 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x38 &  x41 &  x44 &  x47 &  x53 &  x56 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x101 &  x107 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x206 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x275 &  x278 &  x281 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x337 &  x338 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x376 &  x377 &  x380 &  x383 &  x389 &  x392 &  x395 &  x401 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x425 &  x431 &  x434 &  x437 &  x440 &  x443 &  x449 &  x452 &  x455 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x511 &  x515 &  x518 &  x521 &  x533 &  x536 &  x542 &  x545 &  x548 &  x550 &  x554 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x589 &  x590 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x632 &  x635 &  x638 &  x641 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x667 &  x668 &  x671 &  x683 &  x686 &  x689 &  x698 &  x701 &  x703 &  x704 &  x710 &  x716 &  x719 &  x722 &  x725 &  x728 &  x734 &  x737 &  x742 &  x743 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x776 &  x779 &  x781 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x809 &  x812 &  x815 &  x818 &  x820 &  x821 &  x824 &  x827 &  x836 &  x839 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x878 &  x881 &  x884 &  x887 &  x893 &  x896 &  x902 &  x905 &  x908 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x983 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x195 & ~x234 & ~x273;
assign c575 =  x2 &  x8 &  x89 &  x143 &  x191 &  x275 &  x343 &  x356 &  x404 &  x424 &  x440 &  x515 &  x566 &  x581 &  x653 &  x794 &  x857 &  x877 &  x878 &  x908 &  x929 &  x1028 &  x1043 &  x1061 & ~x84 & ~x123 & ~x141 & ~x1104 & ~x1116;
assign c577 =  x2 &  x5 &  x11 &  x17 &  x20 &  x23 &  x26 &  x29 &  x35 &  x41 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x71 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x182 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x230 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x266 &  x275 &  x278 &  x281 &  x287 &  x290 &  x296 &  x299 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x332 &  x335 &  x337 &  x338 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x368 &  x370 &  x374 &  x376 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x419 &  x422 &  x428 &  x434 &  x440 &  x443 &  x446 &  x452 &  x461 &  x464 &  x467 &  x470 &  x476 &  x482 &  x488 &  x491 &  x494 &  x497 &  x500 &  x512 &  x515 &  x518 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x563 &  x566 &  x569 &  x575 &  x578 &  x581 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x611 &  x614 &  x617 &  x623 &  x626 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x656 &  x659 &  x662 &  x664 &  x665 &  x674 &  x677 &  x683 &  x689 &  x692 &  x698 &  x701 &  x703 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x764 &  x767 &  x770 &  x773 &  x776 &  x781 &  x785 &  x788 &  x794 &  x797 &  x800 &  x806 &  x809 &  x815 &  x818 &  x820 &  x821 &  x824 &  x830 &  x833 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x859 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x899 &  x902 &  x905 &  x908 &  x911 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x968 &  x974 &  x977 &  x980 &  x992 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1064 &  x1067 &  x1070 &  x1076 &  x1085 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x120 & ~x159 & ~x198 & ~x237 & ~x276 & ~x393 & ~x591 & ~x630 & ~x669 & ~x1011 & ~x1050;
assign c579 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x169 &  x170 &  x173 &  x176 &  x179 &  x181 &  x182 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x248 &  x251 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x383 &  x386 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x641 &  x644 &  x650 &  x653 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x959 &  x962 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x81 & ~x384 & ~x435 & ~x474 & ~x513 & ~x552;
assign c581 =  x80 &  x107 &  x212 &  x257 &  x383 &  x389 &  x401 &  x524 &  x569 &  x683 &  x770 &  x827 &  x878 &  x953 &  x1076 &  x1079 &  x1115 &  x1118 & ~x123 & ~x138 & ~x540 & ~x669 & ~x747 & ~x786 & ~x1032;
assign c583 =  x86 &  x140 &  x185 &  x212 &  x326 &  x440 &  x488 &  x527 &  x641 &  x664 &  x728 &  x758 &  x781 &  x796 &  x797 &  x835 &  x929 &  x937 &  x953 &  x989 &  x1029 &  x1034 &  x1055 &  x1068 & ~x84;
assign c585 =  x11 &  x29 &  x35 &  x47 &  x53 &  x71 &  x74 &  x89 &  x98 &  x104 &  x128 &  x137 &  x155 &  x164 &  x166 &  x173 &  x176 &  x179 &  x200 &  x212 &  x215 &  x218 &  x233 &  x236 &  x245 &  x257 &  x260 &  x262 &  x263 &  x284 &  x287 &  x293 &  x296 &  x302 &  x305 &  x320 &  x326 &  x335 &  x341 &  x350 &  x362 &  x365 &  x377 &  x383 &  x386 &  x395 &  x404 &  x413 &  x416 &  x452 &  x458 &  x461 &  x464 &  x470 &  x488 &  x509 &  x515 &  x518 &  x524 &  x545 &  x572 &  x578 &  x587 &  x596 &  x605 &  x614 &  x620 &  x629 &  x641 &  x653 &  x665 &  x668 &  x671 &  x677 &  x679 &  x680 &  x686 &  x689 &  x695 &  x710 &  x713 &  x716 &  x722 &  x731 &  x740 &  x749 &  x755 &  x797 &  x806 &  x812 &  x824 &  x827 &  x830 &  x833 &  x842 &  x848 &  x857 &  x860 &  x869 &  x872 &  x875 &  x881 &  x887 &  x899 &  x911 &  x923 &  x932 &  x935 &  x941 &  x956 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x992 &  x1004 &  x1013 &  x1019 &  x1025 &  x1031 &  x1034 &  x1058 &  x1061 &  x1064 &  x1070 &  x1076 &  x1082 &  x1091 &  x1118 &  x1130 & ~x276 & ~x705 & ~x744 & ~x783 & ~x822 & ~x939 & ~x978 & ~x1056;
assign c587 =  x8 &  x20 &  x50 &  x71 &  x89 &  x95 &  x98 &  x116 &  x137 &  x176 &  x179 &  x197 &  x215 &  x233 &  x338 &  x346 &  x347 &  x404 &  x416 &  x455 &  x488 &  x494 &  x503 &  x539 &  x545 &  x608 &  x611 &  x620 &  x626 &  x671 &  x713 &  x716 &  x734 &  x764 &  x776 &  x785 &  x803 &  x842 &  x868 &  x875 &  x887 &  x920 &  x929 &  x944 &  x946 &  x952 &  x971 &  x976 &  x1034 &  x1061 &  x1073 &  x1076 &  x1088 &  x1115 & ~x123 & ~x474 & ~x1059 & ~x1098;
assign c589 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x181 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x220 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x247 &  x248 &  x251 &  x254 &  x257 &  x259 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x299 &  x302 &  x308 &  x311 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x371 &  x377 &  x380 &  x383 &  x389 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x433 &  x434 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x511 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x550 &  x551 &  x557 &  x560 &  x563 &  x566 &  x572 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x589 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x617 &  x620 &  x623 &  x626 &  x629 &  x635 &  x641 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x195 & ~x234;
assign c591 =  x29 &  x82 &  x110 &  x121 &  x160 &  x199 &  x254 &  x269 &  x273 &  x281 &  x302 &  x605 &  x686 &  x794 &  x812 &  x827 &  x848 &  x866 &  x869 &  x881 &  x1010 & ~x111;
assign c593 =  x20 &  x35 &  x41 &  x68 &  x83 &  x92 &  x104 &  x128 &  x143 &  x146 &  x158 &  x167 &  x176 &  x179 &  x221 &  x230 &  x245 &  x248 &  x272 &  x290 &  x296 &  x311 &  x314 &  x320 &  x323 &  x356 &  x389 &  x395 &  x407 &  x419 &  x425 &  x440 &  x442 &  x449 &  x455 &  x478 &  x479 &  x500 &  x515 &  x527 &  x554 &  x563 &  x566 &  x569 &  x575 &  x587 &  x605 &  x611 &  x656 &  x664 &  x665 &  x674 &  x683 &  x686 &  x703 &  x704 &  x707 &  x710 &  x719 &  x722 &  x745 &  x767 &  x776 &  x779 &  x785 &  x820 &  x830 &  x836 &  x872 &  x893 &  x898 &  x920 &  x941 &  x947 &  x956 &  x971 &  x976 &  x980 &  x983 &  x995 &  x1010 &  x1015 &  x1040 &  x1049 &  x1073 &  x1097 &  x1103 &  x1127 & ~x708 & ~x1044 & ~x1083;
assign c595 =  x2 &  x14 &  x17 &  x20 &  x29 &  x44 &  x53 &  x56 &  x65 &  x68 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x110 &  x119 &  x122 &  x125 &  x137 &  x140 &  x155 &  x158 &  x161 &  x164 &  x185 &  x188 &  x197 &  x203 &  x209 &  x218 &  x221 &  x227 &  x230 &  x236 &  x239 &  x245 &  x248 &  x251 &  x263 &  x266 &  x269 &  x272 &  x275 &  x284 &  x296 &  x299 &  x308 &  x317 &  x323 &  x326 &  x332 &  x338 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x364 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x392 &  x395 &  x398 &  x407 &  x410 &  x416 &  x425 &  x428 &  x434 &  x437 &  x443 &  x449 &  x458 &  x461 &  x464 &  x470 &  x473 &  x476 &  x482 &  x485 &  x488 &  x494 &  x497 &  x503 &  x512 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x557 &  x560 &  x572 &  x575 &  x578 &  x584 &  x587 &  x593 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x623 &  x626 &  x628 &  x629 &  x632 &  x638 &  x641 &  x647 &  x656 &  x659 &  x662 &  x665 &  x671 &  x677 &  x689 &  x695 &  x698 &  x701 &  x706 &  x710 &  x713 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x743 &  x745 &  x749 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x784 &  x785 &  x791 &  x794 &  x797 &  x803 &  x812 &  x815 &  x818 &  x821 &  x824 &  x836 &  x839 &  x842 &  x845 &  x857 &  x860 &  x866 &  x878 &  x884 &  x887 &  x890 &  x893 &  x902 &  x908 &  x911 &  x914 &  x917 &  x923 &  x938 &  x950 &  x956 &  x965 &  x974 &  x983 &  x986 &  x992 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1025 &  x1031 &  x1034 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1073 &  x1076 &  x1079 &  x1082 &  x1088 &  x1100 &  x1103 &  x1109 &  x1112 &  x1118 &  x1124 &  x1127 & ~x195 & ~x237 & ~x384 & ~x456;
assign c597 =  x4 &  x5 &  x11 &  x80 &  x107 &  x121 &  x167 &  x212 &  x237 &  x239 &  x263 &  x308 &  x317 &  x323 &  x329 &  x503 &  x602 &  x632 &  x806 &  x851 &  x1025 &  x1124 & ~x1092;
assign c599 =  x35 &  x71 &  x77 &  x164 &  x200 &  x224 &  x245 &  x278 &  x287 &  x293 &  x311 &  x335 &  x401 &  x455 &  x467 &  x488 &  x491 &  x509 &  x548 &  x554 &  x569 &  x593 &  x644 &  x658 &  x677 &  x679 &  x689 &  x773 &  x788 &  x836 &  x857 &  x866 &  x887 &  x977 &  x1055 &  x1091 & ~x69 & ~x588 & ~x609 & ~x939;
assign c5101 =  x14 &  x32 &  x71 &  x80 &  x101 &  x107 &  x122 &  x161 &  x209 &  x248 &  x250 &  x323 &  x350 &  x359 &  x377 &  x452 &  x470 &  x485 &  x497 &  x512 &  x554 &  x560 &  x578 &  x584 &  x596 &  x599 &  x602 &  x641 &  x671 &  x698 &  x725 &  x728 &  x743 &  x779 &  x842 &  x875 &  x887 &  x896 &  x905 &  x908 &  x914 &  x959 &  x989 &  x995 &  x1025 &  x1031 &  x1034 &  x1091 &  x1106 &  x1130 & ~x147 & ~x246 & ~x315 & ~x471 & ~x549 & ~x1056 & ~x1095;
assign c5103 =  x17 &  x248 &  x275 &  x314 &  x343 &  x569 & ~x321 & ~x352 & ~x462 & ~x639 & ~x1077;
assign c5105 =  x23 &  x29 &  x44 &  x56 &  x146 &  x173 &  x179 &  x194 &  x236 &  x248 &  x344 &  x356 &  x382 &  x415 &  x442 &  x470 &  x485 &  x493 &  x512 &  x554 &  x584 &  x590 &  x623 &  x635 &  x674 &  x677 &  x680 &  x695 &  x704 &  x719 &  x734 &  x740 &  x743 &  x770 &  x784 &  x836 &  x839 &  x848 &  x866 &  x875 &  x878 &  x917 &  x920 &  x1004 &  x1019 &  x1040 &  x1058 &  x1103 &  x1112 & ~x81 & ~x657;
assign c5107 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x128 &  x131 &  x134 &  x137 &  x140 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x167 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x220 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x383 &  x389 &  x392 &  x395 &  x401 &  x404 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x458 &  x461 &  x464 &  x467 &  x470 &  x472 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x506 &  x509 &  x511 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x550 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x581 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x703 &  x704 &  x707 &  x710 &  x713 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x749 &  x752 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x829 &  x830 &  x833 &  x839 &  x842 &  x845 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x992 &  x995 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x195 & ~x234;
assign c5109 =  x31 &  x35 &  x41 &  x56 &  x70 &  x77 &  x104 &  x122 &  x164 &  x169 &  x218 &  x236 &  x257 &  x290 &  x302 &  x311 &  x316 &  x355 &  x394 &  x395 &  x446 &  x497 &  x509 &  x512 &  x533 &  x542 &  x626 &  x650 &  x659 &  x794 &  x806 &  x872 &  x911 &  x950 &  x1079 &  x1112 &  x1118 & ~x39;
assign c5111 =  x41 &  x89 &  x140 &  x197 &  x284 &  x296 &  x308 &  x401 &  x422 &  x443 &  x464 &  x518 &  x526 &  x569 &  x572 &  x584 &  x656 &  x671 &  x686 &  x714 &  x770 &  x776 &  x830 &  x833 &  x899 &  x932 &  x953 &  x1010 &  x1043 &  x1049 &  x1073 &  x1082 &  x1100 & ~x1077 & ~x1116;
assign c5113 =  x5 &  x17 &  x20 &  x26 &  x43 &  x44 &  x71 &  x74 &  x82 &  x92 &  x104 &  x122 &  x131 &  x156 &  x167 &  x194 &  x212 &  x233 &  x245 &  x248 &  x260 &  x269 &  x272 &  x290 &  x302 &  x410 &  x413 &  x419 &  x425 &  x428 &  x449 &  x461 &  x467 &  x470 &  x482 &  x497 &  x536 &  x557 &  x578 &  x587 &  x590 &  x599 &  x632 &  x644 &  x665 &  x668 &  x689 &  x740 &  x818 &  x827 &  x851 &  x947 &  x971 &  x974 &  x1013 &  x1016 &  x1022 &  x1043 &  x1049 &  x1058 &  x1076 & ~x72;
assign c5115 =  x11 &  x50 &  x104 &  x110 &  x116 &  x170 &  x197 &  x269 &  x293 &  x308 &  x326 &  x392 &  x425 &  x428 &  x443 &  x446 &  x448 &  x449 &  x461 &  x473 &  x493 &  x494 &  x530 &  x542 &  x563 &  x596 &  x605 &  x611 &  x614 &  x689 &  x704 &  x710 &  x740 &  x745 &  x755 &  x758 &  x784 &  x791 &  x824 &  x833 &  x860 &  x866 &  x890 &  x965 &  x989 &  x1043 &  x1055 &  x1058 &  x1061 &  x1067 &  x1103 &  x1124 & ~x276 & ~x390 & ~x393 & ~x430 & ~x468 & ~x469 & ~x540 & ~x657;
assign c5117 =  x23 &  x32 &  x41 &  x47 &  x56 &  x86 &  x107 &  x143 &  x152 &  x197 &  x203 &  x236 &  x242 &  x263 &  x341 &  x368 &  x380 &  x382 &  x383 &  x386 &  x443 &  x460 &  x487 &  x488 &  x500 &  x515 &  x532 &  x605 &  x617 &  x623 &  x641 &  x644 &  x692 &  x716 &  x746 &  x749 &  x755 &  x776 &  x784 &  x785 &  x788 &  x800 &  x809 &  x842 &  x878 &  x893 &  x899 &  x902 &  x920 &  x974 &  x980 &  x1001 &  x1013 &  x1025 &  x1049 &  x1054 &  x1076 &  x1094 &  x1118 & ~x312 & ~x555;
assign c5119 =  x298 &  x403 &  x1040 & ~x514;
assign c5121 =  x26 &  x32 &  x47 &  x98 &  x116 &  x128 &  x176 &  x188 &  x194 &  x239 &  x254 &  x259 &  x278 &  x281 &  x290 &  x296 &  x302 &  x329 &  x350 &  x356 &  x374 &  x389 &  x410 &  x425 &  x433 &  x437 &  x449 &  x472 &  x482 &  x508 &  x524 &  x563 &  x587 &  x653 &  x662 &  x665 &  x668 &  x680 &  x698 &  x728 &  x758 &  x791 &  x800 &  x851 &  x854 &  x857 &  x869 &  x872 &  x887 &  x899 &  x947 &  x971 &  x998 &  x1013 &  x1025 &  x1073 &  x1091 &  x1127 & ~x165 & ~x195 & ~x234 & ~x513;
assign c5123 =  x29 &  x32 &  x44 &  x50 &  x68 &  x86 &  x110 &  x131 &  x137 &  x254 &  x266 &  x275 &  x317 &  x320 &  x323 &  x341 &  x350 &  x353 &  x376 &  x389 &  x443 &  x448 &  x461 &  x464 &  x473 &  x482 &  x493 &  x559 &  x569 &  x593 &  x620 &  x668 &  x686 &  x689 &  x706 &  x719 &  x785 &  x836 &  x839 &  x851 &  x863 &  x923 &  x950 &  x965 &  x977 &  x1013 &  x1016 &  x1031 & ~x120 & ~x198 & ~x312 & ~x1083;
assign c5125 =  x52 &  x152 &  x161 &  x176 &  x181 &  x239 &  x281 &  x296 &  x551 &  x584 &  x689 &  x794 &  x877 &  x887 &  x974 &  x1022 &  x1115 & ~x171 & ~x405;
assign c5127 =  x17 &  x23 &  x32 &  x41 &  x44 &  x80 &  x101 &  x119 &  x137 &  x140 &  x158 &  x169 &  x173 &  x179 &  x194 &  x207 &  x209 &  x212 &  x227 &  x246 &  x247 &  x266 &  x275 &  x286 &  x325 &  x332 &  x374 &  x386 &  x392 &  x398 &  x410 &  x437 &  x455 &  x470 &  x473 &  x497 &  x506 &  x509 &  x515 &  x536 &  x542 &  x548 &  x551 &  x554 &  x557 &  x560 &  x584 &  x599 &  x605 &  x611 &  x635 &  x647 &  x671 &  x680 &  x686 &  x689 &  x692 &  x701 &  x707 &  x719 &  x728 &  x770 &  x785 &  x797 &  x803 &  x818 &  x821 &  x830 &  x845 &  x869 &  x884 &  x893 &  x911 &  x932 &  x935 &  x959 &  x977 &  x998 &  x1010 &  x1028 &  x1046 &  x1049 &  x1058 &  x1064 &  x1067 &  x1073 &  x1076 &  x1088 &  x1103 &  x1109 &  x1121 &  x1130 & ~x858;
assign c5129 =  x8 &  x17 &  x26 &  x32 &  x35 &  x38 &  x41 &  x44 &  x53 &  x56 &  x59 &  x68 &  x71 &  x82 &  x83 &  x92 &  x101 &  x110 &  x113 &  x116 &  x119 &  x122 &  x128 &  x131 &  x137 &  x140 &  x146 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x179 &  x182 &  x197 &  x200 &  x203 &  x209 &  x212 &  x215 &  x218 &  x224 &  x233 &  x239 &  x245 &  x248 &  x251 &  x254 &  x257 &  x269 &  x272 &  x278 &  x283 &  x284 &  x296 &  x299 &  x302 &  x305 &  x317 &  x320 &  x329 &  x332 &  x344 &  x347 &  x353 &  x359 &  x365 &  x368 &  x383 &  x386 &  x392 &  x395 &  x398 &  x407 &  x413 &  x416 &  x419 &  x422 &  x431 &  x434 &  x437 &  x443 &  x449 &  x455 &  x458 &  x467 &  x470 &  x476 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x506 &  x509 &  x512 &  x515 &  x524 &  x527 &  x536 &  x539 &  x545 &  x557 &  x572 &  x575 &  x584 &  x590 &  x593 &  x596 &  x599 &  x602 &  x608 &  x611 &  x620 &  x626 &  x632 &  x635 &  x644 &  x647 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x683 &  x686 &  x689 &  x701 &  x704 &  x707 &  x710 &  x713 &  x719 &  x725 &  x728 &  x731 &  x740 &  x746 &  x752 &  x755 &  x757 &  x758 &  x773 &  x776 &  x779 &  x791 &  x794 &  x796 &  x797 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x835 &  x839 &  x842 &  x845 &  x857 &  x860 &  x863 &  x875 &  x878 &  x884 &  x887 &  x890 &  x893 &  x902 &  x908 &  x911 &  x914 &  x923 &  x932 &  x941 &  x950 &  x953 &  x956 &  x962 &  x965 &  x968 &  x971 &  x974 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1028 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1076 &  x1082 &  x1085 &  x1088 &  x1094 &  x1100 &  x1102 &  x1103 &  x1106 &  x1121 &  x1124 &  x1127 &  x1130 & ~x264 & ~x588;
assign c5131 =  x2 &  x5 &  x11 &  x14 &  x17 &  x43 &  x47 &  x53 &  x77 &  x80 &  x83 &  x86 &  x101 &  x110 &  x113 &  x119 &  x121 &  x131 &  x140 &  x143 &  x149 &  x152 &  x155 &  x164 &  x170 &  x176 &  x179 &  x191 &  x206 &  x212 &  x221 &  x224 &  x227 &  x230 &  x248 &  x254 &  x260 &  x263 &  x281 &  x284 &  x287 &  x296 &  x299 &  x305 &  x317 &  x320 &  x323 &  x329 &  x332 &  x338 &  x344 &  x350 &  x353 &  x359 &  x362 &  x368 &  x374 &  x386 &  x389 &  x392 &  x422 &  x425 &  x428 &  x434 &  x440 &  x458 &  x485 &  x494 &  x500 &  x506 &  x509 &  x530 &  x536 &  x542 &  x548 &  x557 &  x563 &  x569 &  x572 &  x578 &  x587 &  x590 &  x593 &  x608 &  x611 &  x629 &  x647 &  x656 &  x665 &  x668 &  x674 &  x677 &  x689 &  x692 &  x701 &  x710 &  x722 &  x734 &  x740 &  x752 &  x755 &  x757 &  x761 &  x770 &  x782 &  x788 &  x796 &  x812 &  x827 &  x833 &  x835 &  x842 &  x854 &  x878 &  x893 &  x902 &  x926 &  x932 &  x935 &  x941 &  x947 &  x956 &  x959 &  x965 &  x980 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1016 &  x1025 &  x1028 &  x1030 &  x1034 &  x1043 &  x1046 &  x1064 &  x1069 &  x1076 &  x1085 &  x1088 &  x1094 &  x1108 &  x1118 &  x1124 &  x1130 & ~x414;
assign c5133 =  x20 &  x26 &  x32 &  x56 &  x59 &  x128 &  x170 &  x203 &  x209 &  x230 &  x272 &  x284 &  x296 &  x305 &  x331 &  x344 &  x353 &  x356 &  x382 &  x388 &  x404 &  x409 &  x416 &  x425 &  x428 &  x455 &  x482 &  x485 &  x493 &  x494 &  x530 &  x536 &  x544 &  x551 &  x569 &  x596 &  x608 &  x626 &  x743 &  x779 &  x806 &  x809 &  x812 &  x823 &  x824 &  x839 &  x842 &  x851 &  x869 &  x875 &  x926 &  x944 &  x947 &  x959 &  x962 &  x1013 &  x1028 &  x1049 &  x1061 &  x1067 &  x1088 &  x1094 &  x1097 &  x1130 & ~x390 & ~x469 & ~x618;
assign c5135 =  x32 &  x35 &  x53 &  x59 &  x65 &  x98 &  x137 &  x176 &  x239 &  x257 &  x278 &  x305 &  x314 &  x350 &  x365 &  x409 &  x415 &  x425 &  x434 &  x527 &  x557 &  x590 &  x667 &  x706 &  x791 &  x815 &  x827 &  x833 &  x836 &  x842 &  x860 &  x866 &  x869 &  x881 &  x1010 &  x1013 &  x1016 &  x1103 & ~x765 & ~x766;
assign c5137 =  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x35 &  x37 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x136 &  x137 &  x140 &  x143 &  x146 &  x148 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x185 &  x187 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x214 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x232 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x337 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x403 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x820 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x976 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x3 & ~x39 & ~x42 & ~x78 & ~x81 & ~x117 & ~x156 & ~x195 & ~x198 & ~x234 & ~x237 & ~x276 & ~x315;
assign c5139 =  x68 &  x80 &  x83 &  x91 &  x230 &  x233 &  x395 &  x488 &  x548 &  x563 &  x578 &  x593 &  x602 &  x707 &  x767 &  x779 &  x830 &  x833 &  x835 &  x1019 & ~x648 & ~x900 & ~x1056;
assign c5141 =  x2 &  x5 &  x8 &  x11 &  x14 &  x23 &  x26 &  x29 &  x32 &  x41 &  x47 &  x50 &  x53 &  x56 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x92 &  x98 &  x101 &  x107 &  x113 &  x116 &  x119 &  x125 &  x128 &  x131 &  x137 &  x140 &  x143 &  x149 &  x152 &  x155 &  x161 &  x164 &  x167 &  x170 &  x173 &  x182 &  x188 &  x191 &  x194 &  x200 &  x203 &  x206 &  x215 &  x218 &  x221 &  x224 &  x227 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x269 &  x275 &  x278 &  x281 &  x290 &  x293 &  x302 &  x305 &  x308 &  x311 &  x314 &  x320 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x383 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x428 &  x431 &  x434 &  x437 &  x443 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x473 &  x476 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x506 &  x509 &  x511 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x548 &  x551 &  x554 &  x560 &  x566 &  x569 &  x575 &  x587 &  x593 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x635 &  x641 &  x644 &  x650 &  x653 &  x656 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x716 &  x719 &  x722 &  x728 &  x731 &  x734 &  x737 &  x740 &  x746 &  x749 &  x751 &  x752 &  x761 &  x764 &  x767 &  x773 &  x776 &  x779 &  x782 &  x790 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x818 &  x824 &  x827 &  x828 &  x829 &  x830 &  x833 &  x839 &  x842 &  x848 &  x851 &  x854 &  x860 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x896 &  x902 &  x905 &  x908 &  x911 &  x923 &  x926 &  x929 &  x932 &  x935 &  x941 &  x944 &  x950 &  x953 &  x956 &  x959 &  x962 &  x968 &  x974 &  x986 &  x992 &  x1001 &  x1007 &  x1010 &  x1013 &  x1022 &  x1025 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1097 &  x1103 &  x1106 &  x1109 &  x1118 &  x1124 &  x1127 &  x1130 & ~x156;
assign c5143 =  x47 &  x56 &  x80 &  x179 &  x191 &  x194 &  x287 &  x292 &  x299 &  x308 &  x332 &  x392 &  x419 &  x431 &  x453 &  x458 &  x464 &  x481 &  x494 &  x515 &  x530 &  x536 &  x542 &  x581 &  x584 &  x596 &  x617 &  x644 &  x686 &  x742 &  x770 &  x824 &  x866 &  x881 &  x893 &  x905 &  x941 &  x1016 &  x1025 &  x1049 &  x1115 &  x1130 & ~x630;
assign c5145 =  x2 &  x5 &  x8 &  x11 &  x23 &  x26 &  x43 &  x50 &  x77 &  x82 &  x83 &  x86 &  x95 &  x98 &  x101 &  x110 &  x118 &  x121 &  x122 &  x128 &  x137 &  x149 &  x157 &  x160 &  x164 &  x167 &  x179 &  x182 &  x206 &  x218 &  x221 &  x227 &  x233 &  x248 &  x251 &  x266 &  x272 &  x275 &  x287 &  x293 &  x323 &  x347 &  x362 &  x368 &  x371 &  x392 &  x407 &  x416 &  x431 &  x434 &  x437 &  x443 &  x452 &  x464 &  x485 &  x494 &  x497 &  x506 &  x515 &  x518 &  x524 &  x533 &  x536 &  x554 &  x572 &  x575 &  x578 &  x581 &  x590 &  x596 &  x608 &  x626 &  x635 &  x647 &  x653 &  x656 &  x659 &  x686 &  x689 &  x710 &  x719 &  x728 &  x743 &  x749 &  x755 &  x809 &  x821 &  x827 &  x836 &  x848 &  x854 &  x857 &  x878 &  x893 &  x905 &  x911 &  x914 &  x920 &  x959 &  x968 &  x971 &  x1016 &  x1019 &  x1025 &  x1031 &  x1034 &  x1037 &  x1046 &  x1049 &  x1052 &  x1070 &  x1073 &  x1076 &  x1088 &  x1112 &  x1121 &  x1124 &  x1127 & ~x585 & ~x624 & ~x663 & ~x702 & ~x858 & ~x873 & ~x912;
assign c5147 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x74 &  x83 &  x86 &  x89 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x119 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x173 &  x179 &  x182 &  x185 &  x191 &  x194 &  x200 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x245 &  x248 &  x251 &  x257 &  x260 &  x263 &  x266 &  x269 &  x275 &  x278 &  x281 &  x284 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x320 &  x326 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x401 &  x404 &  x407 &  x410 &  x422 &  x424 &  x425 &  x428 &  x431 &  x434 &  x440 &  x443 &  x446 &  x449 &  x455 &  x461 &  x464 &  x467 &  x470 &  x476 &  x485 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x521 &  x524 &  x530 &  x533 &  x539 &  x545 &  x551 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x626 &  x632 &  x635 &  x638 &  x641 &  x650 &  x653 &  x662 &  x665 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x698 &  x704 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x776 &  x782 &  x800 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x830 &  x836 &  x839 &  x845 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x938 &  x941 &  x950 &  x953 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x980 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1061 &  x1064 &  x1073 &  x1076 &  x1079 &  x1085 &  x1094 &  x1100 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x471 & ~x666 & ~x705 & ~x744 & ~x900 & ~x939 & ~x978 & ~x1017 & ~x1032 & ~x1056 & ~x1065 & ~x1071 & ~x1095;
assign c5149 =  x1 &  x2 &  x4 &  x26 &  x62 &  x65 &  x71 &  x77 &  x80 &  x86 &  x89 &  x92 &  x119 &  x125 &  x131 &  x140 &  x146 &  x149 &  x152 &  x156 &  x157 &  x160 &  x161 &  x164 &  x176 &  x179 &  x185 &  x194 &  x221 &  x235 &  x245 &  x266 &  x269 &  x281 &  x293 &  x296 &  x302 &  x305 &  x323 &  x326 &  x329 &  x335 &  x341 &  x356 &  x374 &  x392 &  x401 &  x407 &  x410 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x458 &  x467 &  x470 &  x473 &  x479 &  x491 &  x503 &  x515 &  x530 &  x551 &  x581 &  x608 &  x626 &  x629 &  x632 &  x635 &  x641 &  x659 &  x662 &  x674 &  x686 &  x698 &  x716 &  x725 &  x728 &  x731 &  x743 &  x755 &  x758 &  x764 &  x773 &  x779 &  x809 &  x815 &  x818 &  x851 &  x860 &  x878 &  x884 &  x890 &  x902 &  x908 &  x926 &  x932 &  x935 &  x947 &  x950 &  x959 &  x968 &  x980 &  x998 &  x1010 &  x1055 &  x1064 &  x1088 &  x1100 &  x1103 &  x1112 &  x1115 &  x1118 &  x1121 & ~x141 & ~x180 & ~x624;
assign c5151 =  x8 &  x11 &  x14 &  x17 &  x23 &  x26 &  x32 &  x38 &  x50 &  x53 &  x65 &  x71 &  x77 &  x83 &  x86 &  x104 &  x110 &  x113 &  x116 &  x122 &  x131 &  x137 &  x140 &  x143 &  x149 &  x161 &  x173 &  x176 &  x179 &  x182 &  x185 &  x194 &  x200 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x251 &  x253 &  x257 &  x260 &  x265 &  x269 &  x304 &  x305 &  x311 &  x317 &  x320 &  x323 &  x325 &  x332 &  x335 &  x337 &  x338 &  x350 &  x356 &  x368 &  x374 &  x380 &  x383 &  x392 &  x398 &  x407 &  x413 &  x419 &  x446 &  x449 &  x455 &  x458 &  x467 &  x470 &  x482 &  x485 &  x488 &  x491 &  x497 &  x503 &  x506 &  x509 &  x518 &  x533 &  x539 &  x542 &  x548 &  x554 &  x557 &  x563 &  x584 &  x587 &  x590 &  x596 &  x605 &  x614 &  x620 &  x650 &  x653 &  x656 &  x662 &  x668 &  x680 &  x686 &  x695 &  x704 &  x710 &  x716 &  x719 &  x731 &  x734 &  x746 &  x752 &  x758 &  x767 &  x770 &  x773 &  x779 &  x791 &  x806 &  x809 &  x812 &  x815 &  x836 &  x839 &  x842 &  x848 &  x854 &  x857 &  x860 &  x869 &  x878 &  x881 &  x887 &  x914 &  x962 &  x965 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1004 &  x1007 &  x1010 &  x1016 &  x1022 &  x1031 &  x1034 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1070 &  x1079 &  x1085 &  x1097 &  x1112 &  x1127 &  x1130 & ~x3 & ~x42 & ~x234 & ~x237 & ~x312 & ~x501 & ~x540;
assign c5153 =  x2 &  x5 &  x32 &  x41 &  x47 &  x53 &  x62 &  x65 &  x74 &  x77 &  x92 &  x104 &  x116 &  x119 &  x125 &  x137 &  x146 &  x149 &  x161 &  x194 &  x212 &  x215 &  x221 &  x224 &  x227 &  x236 &  x248 &  x251 &  x257 &  x281 &  x284 &  x296 &  x302 &  x314 &  x335 &  x344 &  x347 &  x356 &  x362 &  x374 &  x401 &  x407 &  x409 &  x416 &  x419 &  x428 &  x440 &  x449 &  x458 &  x464 &  x470 &  x482 &  x486 &  x487 &  x494 &  x500 &  x521 &  x533 &  x557 &  x560 &  x584 &  x596 &  x599 &  x629 &  x632 &  x638 &  x641 &  x644 &  x647 &  x650 &  x662 &  x667 &  x677 &  x689 &  x695 &  x707 &  x722 &  x728 &  x731 &  x734 &  x745 &  x749 &  x758 &  x761 &  x776 &  x784 &  x797 &  x803 &  x821 &  x823 &  x845 &  x872 &  x893 &  x914 &  x932 &  x959 &  x962 &  x971 &  x974 &  x995 &  x998 &  x1007 &  x1019 &  x1022 &  x1037 &  x1046 &  x1067 &  x1076 &  x1085 &  x1100 &  x1103 &  x1115 &  x1121 & ~x399 & ~x438 & ~x477;
assign c5155 =  x664 &  x742 &  x781 &  x820 &  x859 &  x898 &  x929 & ~x513 & ~x514 & ~x553 & ~x606;
assign c5157 =  x5 &  x8 &  x14 &  x26 &  x44 &  x47 &  x50 &  x53 &  x56 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x89 &  x92 &  x95 &  x101 &  x104 &  x110 &  x119 &  x131 &  x140 &  x149 &  x152 &  x158 &  x173 &  x179 &  x182 &  x188 &  x206 &  x209 &  x212 &  x215 &  x227 &  x236 &  x248 &  x263 &  x266 &  x281 &  x289 &  x296 &  x299 &  x308 &  x311 &  x317 &  x323 &  x332 &  x341 &  x347 &  x353 &  x356 &  x359 &  x362 &  x367 &  x374 &  x385 &  x386 &  x395 &  x401 &  x404 &  x413 &  x425 &  x431 &  x434 &  x452 &  x455 &  x458 &  x470 &  x476 &  x479 &  x484 &  x488 &  x497 &  x500 &  x506 &  x512 &  x521 &  x524 &  x527 &  x530 &  x545 &  x548 &  x551 &  x560 &  x563 &  x569 &  x572 &  x587 &  x596 &  x599 &  x605 &  x608 &  x611 &  x614 &  x617 &  x629 &  x635 &  x644 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x674 &  x677 &  x680 &  x686 &  x692 &  x701 &  x704 &  x707 &  x716 &  x718 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x752 &  x757 &  x761 &  x764 &  x767 &  x770 &  x785 &  x788 &  x796 &  x797 &  x806 &  x827 &  x830 &  x833 &  x835 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x868 &  x869 &  x875 &  x881 &  x893 &  x896 &  x905 &  x907 &  x911 &  x914 &  x920 &  x923 &  x932 &  x935 &  x938 &  x941 &  x962 &  x971 &  x974 &  x977 &  x980 &  x983 &  x991 &  x998 &  x1013 &  x1016 &  x1019 &  x1025 &  x1052 &  x1067 &  x1070 &  x1073 &  x1079 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1102 &  x1112 &  x1124 &  x1130;
assign c5159 =  x4 &  x43 &  x59 &  x62 &  x92 &  x101 &  x121 &  x155 &  x170 &  x182 &  x197 &  x199 &  x200 &  x215 &  x238 &  x254 &  x277 &  x287 &  x293 &  x353 &  x395 &  x458 &  x464 &  x485 &  x488 &  x524 &  x527 &  x536 &  x569 &  x572 &  x632 &  x653 &  x665 &  x686 &  x704 &  x719 &  x728 &  x737 &  x743 &  x746 &  x767 &  x773 &  x782 &  x791 &  x818 &  x824 &  x827 &  x866 &  x884 &  x965 &  x971 &  x1040 &  x1064 &  x1067 &  x1076 &  x1115 & ~x303 & ~x304;
assign c5161 =  x4 &  x11 &  x20 &  x107 &  x143 &  x167 &  x170 &  x257 &  x260 &  x293 &  x302 &  x308 &  x338 &  x341 &  x356 &  x392 &  x410 &  x427 &  x452 &  x473 &  x482 &  x494 &  x512 &  x527 &  x545 &  x572 &  x575 &  x578 &  x581 &  x617 &  x662 &  x677 &  x704 &  x716 &  x767 &  x809 &  x839 &  x893 &  x899 &  x1064 &  x1088 &  x1100 &  x1109 & ~x153 & ~x921 & ~x939;
assign c5163 =  x29 &  x38 &  x86 &  x89 &  x104 &  x121 &  x131 &  x149 &  x160 &  x199 &  x200 &  x212 &  x230 &  x257 &  x269 &  x278 &  x290 &  x326 &  x338 &  x347 &  x353 &  x356 &  x359 &  x362 &  x398 &  x401 &  x407 &  x464 &  x467 &  x470 &  x479 &  x485 &  x503 &  x506 &  x515 &  x566 &  x575 &  x578 &  x581 &  x584 &  x602 &  x623 &  x629 &  x641 &  x659 &  x671 &  x674 &  x680 &  x686 &  x695 &  x731 &  x737 &  x746 &  x758 &  x767 &  x815 &  x851 &  x884 &  x905 &  x908 &  x929 &  x944 &  x956 &  x992 &  x1031 &  x1049 &  x1064 &  x1070 &  x1085 &  x1109 &  x1112 & ~x333 & ~x1017;
assign c5165 =  x20 &  x26 &  x29 &  x47 &  x74 &  x89 &  x104 &  x116 &  x137 &  x140 &  x149 &  x161 &  x167 &  x179 &  x191 &  x238 &  x251 &  x278 &  x308 &  x365 &  x386 &  x407 &  x431 &  x434 &  x440 &  x443 &  x467 &  x473 &  x491 &  x494 &  x515 &  x587 &  x596 &  x614 &  x619 &  x623 &  x641 &  x647 &  x674 &  x707 &  x710 &  x746 &  x752 &  x809 &  x833 &  x845 &  x854 &  x875 &  x983 &  x989 &  x1103 &  x1109 &  x1121 & ~x111 & ~x1053;
assign c5167 =  x4 &  x41 &  x59 &  x89 &  x161 &  x200 &  x221 &  x238 &  x347 &  x452 &  x494 &  x497 &  x506 &  x626 &  x680 &  x728 &  x758 &  x776 &  x851 &  x869 &  x947 &  x1016 &  x1052 &  x1076 &  x1079 & ~x111 & ~x1056;
assign c5169 =  x8 &  x20 &  x35 &  x38 &  x41 &  x53 &  x83 &  x125 &  x134 &  x137 &  x146 &  x158 &  x161 &  x167 &  x176 &  x179 &  x185 &  x194 &  x212 &  x218 &  x236 &  x256 &  x266 &  x346 &  x350 &  x370 &  x374 &  x404 &  x427 &  x440 &  x452 &  x467 &  x479 &  x512 &  x602 &  x611 &  x625 &  x626 &  x632 &  x638 &  x743 &  x749 &  x752 &  x761 &  x788 &  x881 &  x911 &  x917 &  x920 &  x923 &  x929 &  x938 &  x1007 &  x1025 &  x1034 &  x1043 &  x1088 &  x1106 &  x1109 &  x1124 &  x1127 & ~x129 & ~x474;
assign c5171 =  x2 &  x5 &  x8 &  x17 &  x23 &  x26 &  x47 &  x56 &  x74 &  x110 &  x125 &  x140 &  x158 &  x176 &  x182 &  x188 &  x191 &  x200 &  x203 &  x209 &  x215 &  x224 &  x236 &  x242 &  x245 &  x329 &  x353 &  x356 &  x362 &  x392 &  x404 &  x434 &  x458 &  x509 &  x512 &  x554 &  x563 &  x569 &  x581 &  x590 &  x599 &  x602 &  x620 &  x677 &  x683 &  x701 &  x704 &  x752 &  x755 &  x758 &  x773 &  x800 &  x842 &  x866 &  x887 &  x896 &  x899 &  x908 &  x911 &  x926 &  x938 &  x980 &  x989 &  x992 &  x1004 &  x1007 &  x1010 &  x1022 &  x1037 &  x1046 &  x1049 &  x1067 &  x1079 &  x1088 &  x1094 &  x1106 & ~x213 & ~x240 & ~x318 & ~x319 & ~x358 & ~x432;
assign c5173 =  x2 &  x5 &  x20 &  x23 &  x29 &  x32 &  x35 &  x50 &  x53 &  x59 &  x62 &  x65 &  x74 &  x77 &  x86 &  x89 &  x95 &  x98 &  x101 &  x110 &  x113 &  x116 &  x119 &  x134 &  x137 &  x140 &  x149 &  x155 &  x158 &  x161 &  x167 &  x176 &  x182 &  x185 &  x191 &  x197 &  x203 &  x206 &  x209 &  x212 &  x215 &  x224 &  x230 &  x233 &  x239 &  x248 &  x251 &  x254 &  x263 &  x266 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x299 &  x302 &  x305 &  x308 &  x311 &  x335 &  x338 &  x341 &  x347 &  x350 &  x356 &  x365 &  x371 &  x374 &  x383 &  x389 &  x392 &  x415 &  x416 &  x419 &  x422 &  x425 &  x431 &  x442 &  x449 &  x452 &  x470 &  x473 &  x482 &  x488 &  x494 &  x500 &  x506 &  x512 &  x518 &  x536 &  x542 &  x545 &  x554 &  x556 &  x557 &  x560 &  x566 &  x569 &  x572 &  x578 &  x581 &  x587 &  x590 &  x593 &  x599 &  x611 &  x614 &  x620 &  x623 &  x626 &  x629 &  x635 &  x641 &  x644 &  x647 &  x650 &  x659 &  x664 &  x680 &  x683 &  x689 &  x695 &  x701 &  x704 &  x707 &  x710 &  x713 &  x722 &  x734 &  x737 &  x742 &  x746 &  x749 &  x752 &  x761 &  x764 &  x767 &  x770 &  x776 &  x779 &  x781 &  x784 &  x785 &  x788 &  x794 &  x803 &  x806 &  x809 &  x812 &  x815 &  x824 &  x833 &  x836 &  x842 &  x848 &  x851 &  x854 &  x857 &  x859 &  x863 &  x866 &  x869 &  x872 &  x875 &  x881 &  x884 &  x893 &  x896 &  x898 &  x908 &  x911 &  x920 &  x932 &  x937 &  x938 &  x941 &  x944 &  x947 &  x959 &  x968 &  x971 &  x974 &  x977 &  x983 &  x986 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1031 &  x1034 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1094 &  x1100 &  x1118 &  x1124 &  x1130 & ~x273 & ~x276 & ~x351 & ~x354 & ~x393 & ~x432;
assign c5175 =  x56 &  x82 &  x89 &  x92 &  x98 &  x230 &  x238 &  x248 &  x254 &  x257 &  x277 &  x290 &  x326 &  x362 &  x395 &  x404 &  x431 &  x449 &  x455 &  x479 &  x491 &  x509 &  x536 &  x539 &  x545 &  x554 &  x599 &  x602 &  x644 &  x662 &  x674 &  x698 &  x710 &  x743 &  x749 &  x757 &  x767 &  x773 &  x788 &  x791 &  x796 &  x797 &  x962 &  x986 &  x989 &  x1004 &  x1010 &  x1073 &  x1085 & ~x453 & ~x492;
assign c5177 =  x13 &  x20 &  x25 &  x26 &  x29 &  x52 &  x146 &  x182 &  x238 &  x245 &  x277 &  x302 &  x316 &  x338 &  x341 &  x377 &  x500 &  x545 &  x575 &  x581 &  x611 &  x614 &  x650 &  x665 &  x692 &  x737 &  x749 &  x761 &  x887 &  x932 &  x980 &  x989 &  x992 &  x1028 &  x1085 &  x1088 & ~x858 & ~x1014 & ~x1092;
assign c5179 =  x5 &  x26 &  x59 &  x65 &  x68 &  x80 &  x98 &  x101 &  x116 &  x134 &  x143 &  x155 &  x203 &  x215 &  x218 &  x224 &  x239 &  x245 &  x251 &  x254 &  x260 &  x272 &  x287 &  x290 &  x302 &  x314 &  x350 &  x353 &  x365 &  x370 &  x386 &  x410 &  x413 &  x433 &  x443 &  x452 &  x482 &  x488 &  x503 &  x509 &  x515 &  x518 &  x524 &  x542 &  x554 &  x563 &  x569 &  x578 &  x581 &  x623 &  x628 &  x638 &  x644 &  x653 &  x659 &  x662 &  x695 &  x713 &  x722 &  x734 &  x740 &  x743 &  x764 &  x767 &  x776 &  x812 &  x824 &  x833 &  x842 &  x857 &  x866 &  x881 &  x890 &  x923 &  x932 &  x944 &  x953 &  x962 &  x965 &  x995 &  x998 &  x1025 &  x1031 &  x1058 &  x1070 &  x1100 &  x1130 & ~x390 & ~x771 & ~x810;
assign c5181 =  x4 & ~x162 & ~x711 & ~x858;
assign c5183 =  x2 &  x5 &  x8 &  x11 &  x17 &  x20 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x50 &  x56 &  x62 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x170 &  x173 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x203 &  x206 &  x212 &  x218 &  x221 &  x230 &  x236 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x272 &  x275 &  x278 &  x281 &  x284 &  x290 &  x293 &  x299 &  x302 &  x305 &  x308 &  x314 &  x317 &  x320 &  x323 &  x326 &  x332 &  x335 &  x338 &  x350 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x377 &  x380 &  x383 &  x392 &  x398 &  x404 &  x407 &  x410 &  x419 &  x422 &  x425 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x458 &  x467 &  x469 &  x470 &  x476 &  x488 &  x494 &  x503 &  x506 &  x507 &  x508 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x545 &  x547 &  x548 &  x551 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x581 &  x584 &  x586 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x617 &  x620 &  x623 &  x625 &  x626 &  x629 &  x632 &  x635 &  x638 &  x644 &  x647 &  x650 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x716 &  x719 &  x722 &  x725 &  x728 &  x734 &  x737 &  x740 &  x743 &  x746 &  x755 &  x758 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x845 &  x848 &  x851 &  x857 &  x860 &  x863 &  x866 &  x875 &  x881 &  x884 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x941 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x195 & ~x435 & ~x492 & ~x570 & ~x726;
assign c5185 =  x2 &  x5 &  x8 &  x17 &  x26 &  x32 &  x35 &  x38 &  x41 &  x47 &  x50 &  x59 &  x62 &  x65 &  x77 &  x83 &  x92 &  x95 &  x98 &  x110 &  x119 &  x122 &  x125 &  x128 &  x131 &  x140 &  x143 &  x146 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x227 &  x239 &  x245 &  x257 &  x266 &  x272 &  x278 &  x284 &  x302 &  x308 &  x311 &  x316 &  x317 &  x323 &  x326 &  x329 &  x341 &  x344 &  x347 &  x356 &  x359 &  x362 &  x371 &  x374 &  x377 &  x383 &  x389 &  x395 &  x398 &  x401 &  x416 &  x422 &  x425 &  x431 &  x433 &  x443 &  x449 &  x455 &  x464 &  x470 &  x479 &  x494 &  x497 &  x503 &  x509 &  x521 &  x536 &  x542 &  x548 &  x551 &  x557 &  x560 &  x566 &  x569 &  x572 &  x575 &  x581 &  x593 &  x599 &  x602 &  x605 &  x611 &  x620 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x674 &  x680 &  x686 &  x692 &  x698 &  x701 &  x704 &  x707 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x743 &  x746 &  x752 &  x764 &  x767 &  x773 &  x782 &  x788 &  x791 &  x797 &  x800 &  x806 &  x809 &  x812 &  x818 &  x821 &  x833 &  x839 &  x845 &  x848 &  x851 &  x860 &  x875 &  x878 &  x881 &  x884 &  x890 &  x893 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x926 &  x932 &  x938 &  x941 &  x947 &  x956 &  x959 &  x962 &  x965 &  x971 &  x974 &  x977 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1034 &  x1037 &  x1043 &  x1049 &  x1052 &  x1064 &  x1076 &  x1079 &  x1082 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 &  x1115 &  x1118 &  x1124 &  x1127 &  x1130 & ~x39 & ~x54 & ~x78 & ~x228 & ~x741 & ~x780 & ~x819 & ~x858;
assign c5187 =  x77 &  x83 &  x95 &  x107 &  x122 &  x130 &  x208 &  x247 &  x263 &  x275 &  x341 &  x383 &  x392 &  x431 &  x488 &  x587 &  x608 &  x671 &  x683 &  x770 &  x797 &  x809 &  x836 &  x881 &  x932 &  x947 &  x956 &  x983 &  x998 &  x1064 & ~x222 & ~x255 & ~x741;
assign c5189 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x158 &  x161 &  x164 &  x170 &  x173 &  x175 &  x176 &  x179 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x305 &  x308 &  x311 &  x314 &  x316 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x428 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x464 &  x467 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x569 &  x575 &  x578 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x857 &  x860 &  x863 &  x866 &  x869 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 &  x1130 & ~x3 & ~x42 & ~x78 & ~x81 & ~x117;
assign c5191 =  x169 &  x566 & ~x111 & ~x183 & ~x216 & ~x702 & ~x858 & ~x897 & ~x936 & ~x1092;
assign c5193 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x83 &  x86 &  x92 &  x98 &  x104 &  x107 &  x110 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x140 &  x146 &  x155 &  x161 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x197 &  x200 &  x203 &  x206 &  x209 &  x215 &  x230 &  x233 &  x236 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x275 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x308 &  x311 &  x314 &  x317 &  x320 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x353 &  x359 &  x362 &  x365 &  x368 &  x371 &  x376 &  x380 &  x383 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x413 &  x415 &  x416 &  x419 &  x422 &  x428 &  x437 &  x449 &  x452 &  x458 &  x464 &  x467 &  x470 &  x476 &  x479 &  x482 &  x488 &  x497 &  x503 &  x506 &  x509 &  x512 &  x515 &  x521 &  x524 &  x527 &  x533 &  x539 &  x542 &  x545 &  x551 &  x554 &  x557 &  x560 &  x569 &  x578 &  x584 &  x587 &  x589 &  x590 &  x593 &  x599 &  x602 &  x608 &  x614 &  x620 &  x623 &  x626 &  x628 &  x629 &  x632 &  x635 &  x638 &  x641 &  x650 &  x653 &  x656 &  x659 &  x668 &  x671 &  x680 &  x683 &  x689 &  x692 &  x695 &  x698 &  x701 &  x703 &  x707 &  x710 &  x713 &  x716 &  x719 &  x728 &  x734 &  x737 &  x742 &  x743 &  x746 &  x749 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x779 &  x781 &  x782 &  x785 &  x788 &  x791 &  x797 &  x803 &  x806 &  x809 &  x815 &  x818 &  x820 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x857 &  x859 &  x866 &  x872 &  x875 &  x884 &  x887 &  x890 &  x896 &  x905 &  x914 &  x920 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x977 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1015 &  x1016 &  x1019 &  x1022 &  x1024 &  x1034 &  x1037 &  x1040 &  x1049 &  x1052 &  x1054 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1093 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x273 & ~x312 & ~x351;
assign c5195 =  x41 &  x47 &  x65 &  x68 &  x86 &  x98 &  x101 &  x110 &  x116 &  x134 &  x137 &  x140 &  x143 &  x158 &  x176 &  x185 &  x191 &  x212 &  x215 &  x218 &  x221 &  x236 &  x263 &  x269 &  x281 &  x284 &  x287 &  x296 &  x302 &  x308 &  x326 &  x329 &  x338 &  x347 &  x353 &  x356 &  x365 &  x370 &  x377 &  x380 &  x398 &  x425 &  x440 &  x445 &  x485 &  x491 &  x500 &  x503 &  x506 &  x512 &  x515 &  x533 &  x551 &  x557 &  x572 &  x587 &  x593 &  x596 &  x626 &  x629 &  x635 &  x641 &  x671 &  x677 &  x698 &  x719 &  x722 &  x740 &  x746 &  x785 &  x794 &  x797 &  x800 &  x845 &  x866 &  x878 &  x881 &  x893 &  x908 &  x923 &  x941 &  x953 &  x956 &  x983 &  x1013 &  x1067 &  x1082 &  x1094 &  x1106 &  x1108 &  x1115 &  x1127 &  x1130 & ~x84 & ~x162 & ~x474 & ~x513 & ~x816;
assign c5197 =  x4 &  x14 &  x35 &  x38 &  x43 &  x47 &  x82 &  x104 &  x110 &  x125 &  x128 &  x146 &  x155 &  x170 &  x197 &  x206 &  x248 &  x263 &  x277 &  x284 &  x296 &  x308 &  x323 &  x332 &  x362 &  x365 &  x383 &  x389 &  x395 &  x407 &  x419 &  x443 &  x461 &  x467 &  x500 &  x506 &  x515 &  x524 &  x542 &  x551 &  x566 &  x629 &  x632 &  x638 &  x644 &  x653 &  x656 &  x680 &  x683 &  x692 &  x695 &  x698 &  x707 &  x719 &  x743 &  x755 &  x767 &  x773 &  x779 &  x812 &  x818 &  x824 &  x830 &  x835 &  x839 &  x842 &  x845 &  x851 &  x857 &  x860 &  x920 &  x926 &  x941 &  x944 &  x950 &  x956 &  x968 &  x998 &  x1013 &  x1019 &  x1046 &  x1061 &  x1070 &  x1073 &  x1082 &  x1097 & ~x936 & ~x1014;
assign c5199 =  x14 &  x26 &  x50 &  x59 &  x86 &  x89 &  x95 &  x98 &  x101 &  x107 &  x113 &  x119 &  x121 &  x125 &  x134 &  x137 &  x140 &  x158 &  x173 &  x176 &  x185 &  x194 &  x199 &  x236 &  x239 &  x245 &  x263 &  x266 &  x284 &  x293 &  x305 &  x308 &  x311 &  x314 &  x323 &  x329 &  x344 &  x350 &  x371 &  x374 &  x389 &  x395 &  x398 &  x401 &  x404 &  x413 &  x437 &  x440 &  x452 &  x455 &  x461 &  x467 &  x469 &  x470 &  x473 &  x479 &  x491 &  x509 &  x521 &  x527 &  x530 &  x551 &  x554 &  x557 &  x563 &  x581 &  x593 &  x596 &  x599 &  x608 &  x629 &  x644 &  x653 &  x659 &  x662 &  x671 &  x674 &  x677 &  x680 &  x683 &  x719 &  x725 &  x728 &  x764 &  x773 &  x776 &  x779 &  x782 &  x791 &  x800 &  x818 &  x824 &  x845 &  x848 &  x854 &  x863 &  x872 &  x878 &  x884 &  x887 &  x911 &  x920 &  x923 &  x935 &  x938 &  x941 &  x962 &  x977 &  x980 &  x992 &  x1013 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1043 &  x1061 &  x1073 &  x1091 &  x1097 &  x1103 &  x1106 &  x1115 &  x1118 & ~x666 & ~x681 & ~x705 & ~x744 & ~x783 & ~x822 & ~x939;
assign c5201 =  x2 &  x8 &  x14 &  x17 &  x23 &  x32 &  x38 &  x41 &  x47 &  x59 &  x65 &  x71 &  x77 &  x83 &  x86 &  x95 &  x116 &  x125 &  x128 &  x134 &  x146 &  x155 &  x161 &  x167 &  x170 &  x173 &  x176 &  x182 &  x191 &  x194 &  x203 &  x227 &  x230 &  x236 &  x239 &  x245 &  x247 &  x260 &  x263 &  x269 &  x275 &  x287 &  x290 &  x292 &  x293 &  x329 &  x332 &  x335 &  x344 &  x359 &  x365 &  x380 &  x386 &  x389 &  x392 &  x410 &  x413 &  x416 &  x419 &  x431 &  x434 &  x440 &  x443 &  x446 &  x452 &  x455 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x497 &  x509 &  x518 &  x521 &  x533 &  x539 &  x548 &  x557 &  x563 &  x569 &  x572 &  x581 &  x596 &  x599 &  x608 &  x614 &  x617 &  x641 &  x653 &  x656 &  x659 &  x674 &  x680 &  x701 &  x710 &  x716 &  x719 &  x722 &  x728 &  x734 &  x746 &  x749 &  x752 &  x758 &  x764 &  x776 &  x779 &  x800 &  x821 &  x824 &  x827 &  x830 &  x833 &  x835 &  x836 &  x860 &  x863 &  x866 &  x874 &  x878 &  x884 &  x890 &  x893 &  x896 &  x899 &  x905 &  x908 &  x911 &  x914 &  x929 &  x932 &  x935 &  x953 &  x956 &  x974 &  x992 &  x995 &  x1001 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1034 &  x1037 &  x1040 &  x1046 &  x1055 &  x1058 &  x1070 &  x1082 &  x1085 &  x1094 &  x1100 &  x1106 &  x1121 &  x1124 & ~x81 & ~x1056;
assign c5203 =  x26 &  x29 &  x38 &  x41 &  x53 &  x56 &  x68 &  x74 &  x77 &  x80 &  x86 &  x95 &  x98 &  x104 &  x113 &  x125 &  x128 &  x131 &  x140 &  x149 &  x158 &  x197 &  x203 &  x209 &  x212 &  x226 &  x242 &  x248 &  x251 &  x257 &  x265 &  x266 &  x290 &  x293 &  x298 &  x299 &  x314 &  x317 &  x335 &  x337 &  x344 &  x376 &  x383 &  x395 &  x398 &  x404 &  x419 &  x437 &  x440 &  x452 &  x464 &  x509 &  x512 &  x515 &  x521 &  x524 &  x536 &  x557 &  x566 &  x578 &  x611 &  x617 &  x623 &  x626 &  x629 &  x635 &  x656 &  x659 &  x671 &  x692 &  x706 &  x737 &  x740 &  x761 &  x767 &  x776 &  x785 &  x794 &  x818 &  x863 &  x884 &  x899 &  x902 &  x905 &  x914 &  x932 &  x968 &  x974 &  x989 &  x992 &  x1013 &  x1028 &  x1034 &  x1085 &  x1100 &  x1121 &  x1124 & ~x120 & ~x273 & ~x405;
assign c5205 =  x11 &  x14 &  x17 &  x20 &  x26 &  x50 &  x65 &  x71 &  x86 &  x91 &  x95 &  x101 &  x116 &  x128 &  x131 &  x134 &  x140 &  x143 &  x161 &  x170 &  x173 &  x185 &  x188 &  x191 &  x197 &  x200 &  x209 &  x224 &  x242 &  x245 &  x248 &  x254 &  x257 &  x269 &  x296 &  x302 &  x316 &  x317 &  x338 &  x347 &  x353 &  x365 &  x368 &  x374 &  x392 &  x395 &  x398 &  x413 &  x419 &  x425 &  x428 &  x446 &  x452 &  x458 &  x461 &  x464 &  x467 &  x470 &  x503 &  x509 &  x512 &  x524 &  x542 &  x545 &  x548 &  x557 &  x560 &  x578 &  x596 &  x599 &  x602 &  x611 &  x614 &  x623 &  x653 &  x671 &  x698 &  x716 &  x722 &  x725 &  x737 &  x752 &  x755 &  x791 &  x818 &  x821 &  x830 &  x848 &  x854 &  x860 &  x863 &  x866 &  x875 &  x881 &  x893 &  x899 &  x932 &  x944 &  x947 &  x950 &  x959 &  x965 &  x968 &  x977 &  x980 &  x992 &  x1001 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1055 &  x1067 &  x1076 &  x1124 & ~x39 & ~x117 & ~x228 & ~x1092;
assign c5207 =  x164 &  x167 &  x184 &  x227 &  x305 &  x323 &  x418 &  x419 &  x481 &  x518 &  x595 &  x597 &  x598 &  x602 &  x614 &  x620 &  x656 &  x665 &  x839 &  x863 &  x902 &  x917 &  x998 & ~x276;
assign c5209 =  x62 &  x65 &  x113 &  x134 &  x143 &  x245 &  x305 &  x401 &  x476 &  x518 &  x536 &  x587 &  x589 &  x647 &  x683 &  x1007 &  x1046 &  x1100 & ~x313 & ~x384 & ~x444;
assign c5211 =  x8 &  x170 &  x242 &  x287 &  x304 &  x317 &  x335 &  x347 &  x380 &  x385 &  x416 &  x422 &  x481 &  x521 &  x545 &  x764 &  x833 &  x908 &  x965 &  x1082 &  x1127 & ~x474 & ~x513 & ~x708 & ~x894 & ~x1077;
assign c5213 =  x2 &  x32 &  x35 &  x41 &  x59 &  x77 &  x161 &  x200 &  x278 &  x314 &  x335 &  x349 &  x401 &  x407 &  x410 &  x413 &  x452 &  x461 &  x554 &  x593 &  x623 &  x806 &  x842 &  x914 &  x920 &  x923 &  x980 &  x1030 &  x1040 &  x1061 &  x1069 &  x1070 &  x1108 &  x1109 & ~x273 & ~x1038;
assign c5215 =  x358 &  x376 &  x409 &  x524 &  x667 &  x706 &  x1022 & ~x117 & ~x391 & ~x501;
assign c5217 =  x2 &  x5 &  x8 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x50 &  x59 &  x68 &  x83 &  x89 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x122 &  x125 &  x128 &  x146 &  x149 &  x155 &  x164 &  x200 &  x206 &  x245 &  x248 &  x254 &  x263 &  x266 &  x269 &  x272 &  x278 &  x284 &  x287 &  x293 &  x311 &  x317 &  x332 &  x338 &  x344 &  x359 &  x365 &  x374 &  x377 &  x380 &  x395 &  x398 &  x407 &  x425 &  x434 &  x437 &  x440 &  x452 &  x458 &  x473 &  x476 &  x482 &  x485 &  x488 &  x491 &  x503 &  x524 &  x533 &  x542 &  x545 &  x546 &  x557 &  x569 &  x575 &  x581 &  x584 &  x586 &  x587 &  x602 &  x614 &  x626 &  x635 &  x638 &  x650 &  x656 &  x662 &  x665 &  x671 &  x674 &  x698 &  x710 &  x728 &  x734 &  x764 &  x767 &  x770 &  x776 &  x781 &  x782 &  x788 &  x815 &  x818 &  x827 &  x833 &  x839 &  x848 &  x851 &  x854 &  x860 &  x863 &  x869 &  x872 &  x905 &  x911 &  x917 &  x920 &  x926 &  x938 &  x944 &  x950 &  x980 &  x986 &  x992 &  x1001 &  x1007 &  x1010 &  x1028 &  x1037 &  x1043 &  x1046 &  x1049 &  x1055 &  x1058 &  x1067 &  x1082 &  x1091 &  x1100 &  x1115 &  x1118 &  x1124 &  x1130 & ~x195 & ~x474 & ~x513 & ~x927;
assign c5219 =  x5 &  x8 &  x11 &  x17 &  x47 &  x65 &  x77 &  x80 &  x107 &  x119 &  x149 &  x152 &  x170 &  x179 &  x194 &  x203 &  x221 &  x233 &  x248 &  x269 &  x299 &  x305 &  x308 &  x311 &  x320 &  x323 &  x329 &  x338 &  x347 &  x353 &  x380 &  x410 &  x449 &  x494 &  x527 &  x530 &  x545 &  x551 &  x557 &  x560 &  x575 &  x599 &  x602 &  x644 &  x653 &  x659 &  x677 &  x680 &  x683 &  x692 &  x719 &  x728 &  x740 &  x749 &  x755 &  x758 &  x794 &  x803 &  x824 &  x842 &  x860 &  x908 &  x920 &  x935 &  x941 &  x956 &  x959 &  x962 &  x983 &  x1004 &  x1025 &  x1028 &  x1043 &  x1046 &  x1064 &  x1088 &  x1100 &  x1118 & ~x687 & ~x688 & ~x900 & ~x939 & ~x1017 & ~x1095;
assign c5221 =  x2 &  x20 &  x116 &  x134 &  x200 &  x205 &  x212 &  x230 &  x248 &  x260 &  x269 &  x275 &  x296 &  x386 &  x392 &  x398 &  x407 &  x424 &  x425 &  x461 &  x506 &  x539 &  x551 &  x575 &  x596 &  x611 &  x650 &  x653 &  x680 &  x758 &  x761 &  x779 &  x782 &  x788 &  x794 &  x812 &  x821 &  x827 &  x860 &  x878 &  x908 &  x931 &  x941 &  x968 &  x1076 &  x1100 & ~x381 & ~x459 & ~x471 & ~x627 & ~x666 & ~x822;
assign c5223 =  x20 &  x32 &  x53 &  x62 &  x68 &  x83 &  x86 &  x107 &  x122 &  x134 &  x152 &  x160 &  x164 &  x182 &  x185 &  x197 &  x206 &  x257 &  x269 &  x277 &  x278 &  x290 &  x293 &  x305 &  x329 &  x332 &  x341 &  x344 &  x368 &  x371 &  x383 &  x392 &  x401 &  x416 &  x431 &  x437 &  x455 &  x461 &  x500 &  x536 &  x554 &  x566 &  x611 &  x614 &  x644 &  x668 &  x683 &  x710 &  x734 &  x737 &  x749 &  x752 &  x761 &  x776 &  x785 &  x794 &  x812 &  x815 &  x839 &  x848 &  x851 &  x854 &  x881 &  x920 &  x932 &  x935 &  x959 &  x962 &  x989 &  x1010 &  x1040 &  x1043 &  x1079 & ~x336 & ~x460;
assign c5225 =  x5 &  x14 &  x22 &  x29 &  x35 &  x38 &  x44 &  x47 &  x53 &  x55 &  x62 &  x65 &  x71 &  x80 &  x95 &  x100 &  x104 &  x110 &  x116 &  x118 &  x119 &  x122 &  x131 &  x143 &  x144 &  x146 &  x149 &  x152 &  x158 &  x161 &  x164 &  x167 &  x176 &  x184 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x212 &  x218 &  x221 &  x224 &  x227 &  x230 &  x236 &  x239 &  x245 &  x263 &  x278 &  x284 &  x296 &  x311 &  x347 &  x350 &  x353 &  x356 &  x359 &  x368 &  x371 &  x380 &  x392 &  x395 &  x398 &  x401 &  x410 &  x413 &  x419 &  x428 &  x437 &  x449 &  x452 &  x461 &  x470 &  x476 &  x479 &  x482 &  x488 &  x497 &  x500 &  x509 &  x521 &  x524 &  x527 &  x536 &  x548 &  x557 &  x572 &  x575 &  x596 &  x598 &  x599 &  x602 &  x605 &  x617 &  x623 &  x641 &  x644 &  x647 &  x653 &  x659 &  x665 &  x668 &  x677 &  x680 &  x683 &  x692 &  x695 &  x701 &  x707 &  x710 &  x713 &  x716 &  x719 &  x728 &  x731 &  x734 &  x740 &  x743 &  x746 &  x755 &  x764 &  x770 &  x776 &  x785 &  x788 &  x791 &  x797 &  x800 &  x803 &  x809 &  x818 &  x833 &  x845 &  x848 &  x851 &  x854 &  x857 &  x863 &  x869 &  x878 &  x884 &  x890 &  x893 &  x896 &  x902 &  x908 &  x914 &  x920 &  x923 &  x935 &  x938 &  x941 &  x956 &  x959 &  x962 &  x968 &  x977 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1013 &  x1016 &  x1019 &  x1025 &  x1034 &  x1037 &  x1043 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1085 &  x1094 &  x1109 &  x1115 &  x1118 &  x1130 & ~x1011 & ~x1050;
assign c5227 =  x230 & ~x123 & ~x162 & ~x201 & ~x321;
assign c5229 =  x17 &  x41 &  x44 &  x56 &  x62 &  x65 &  x74 &  x83 &  x122 &  x131 &  x134 &  x143 &  x161 &  x164 &  x170 &  x176 &  x185 &  x191 &  x203 &  x209 &  x221 &  x230 &  x233 &  x236 &  x239 &  x245 &  x254 &  x263 &  x269 &  x272 &  x287 &  x293 &  x308 &  x311 &  x320 &  x323 &  x329 &  x338 &  x344 &  x347 &  x371 &  x377 &  x380 &  x395 &  x401 &  x407 &  x410 &  x437 &  x449 &  x455 &  x506 &  x536 &  x545 &  x551 &  x554 &  x557 &  x575 &  x578 &  x590 &  x596 &  x617 &  x632 &  x659 &  x671 &  x674 &  x707 &  x713 &  x722 &  x728 &  x746 &  x749 &  x752 &  x757 &  x764 &  x773 &  x779 &  x782 &  x788 &  x796 &  x797 &  x800 &  x803 &  x809 &  x821 &  x839 &  x851 &  x854 &  x857 &  x887 &  x908 &  x911 &  x983 &  x997 &  x1001 &  x1016 &  x1019 &  x1028 &  x1031 &  x1034 &  x1040 &  x1061 &  x1076 &  x1082 &  x1088 &  x1091 &  x1100 &  x1112 &  x1130 & ~x471 & ~x570 & ~x588 & ~x627 & ~x648 & ~x744 & ~x861;
assign c5231 =  x52 &  x92 &  x110 &  x128 &  x161 &  x182 &  x197 &  x212 &  x221 &  x236 &  x254 &  x257 &  x263 &  x272 &  x305 &  x368 &  x380 &  x401 &  x433 &  x461 &  x497 &  x521 &  x563 &  x593 &  x644 &  x689 &  x728 &  x791 &  x809 &  x851 &  x860 &  x863 &  x866 &  x881 &  x932 &  x983 &  x1022 &  x1034 &  x1058 &  x1061 &  x1064 &  x1097 &  x1121 & ~x72 & ~x261 & ~x267 & ~x897 & ~x975;
assign c5233 =  x17 &  x449 &  x698 &  x706 &  x740 &  x781 &  x857 &  x859 &  x1049 &  x1124 & ~x393 & ~x432 & ~x450 & ~x462 & ~x540;
assign c5235 =  x62 &  x71 &  x113 &  x253 &  x578 &  x586 &  x995 & ~x345 & ~x553;
assign c5237 =  x5 &  x8 &  x41 &  x47 &  x65 &  x68 &  x92 &  x101 &  x107 &  x110 &  x113 &  x119 &  x122 &  x134 &  x137 &  x176 &  x269 &  x290 &  x296 &  x302 &  x308 &  x326 &  x338 &  x371 &  x389 &  x392 &  x394 &  x395 &  x401 &  x428 &  x431 &  x434 &  x440 &  x443 &  x464 &  x479 &  x485 &  x497 &  x524 &  x530 &  x548 &  x557 &  x575 &  x578 &  x608 &  x614 &  x620 &  x623 &  x626 &  x644 &  x647 &  x683 &  x695 &  x707 &  x722 &  x725 &  x734 &  x737 &  x746 &  x794 &  x809 &  x830 &  x836 &  x842 &  x845 &  x848 &  x857 &  x872 &  x884 &  x890 &  x917 &  x971 &  x974 &  x1016 &  x1040 &  x1043 &  x1055 &  x1073 &  x1082 &  x1094 &  x1103 &  x1112 &  x1121 & ~x583 & ~x1050;
assign c5239 =  x20 &  x41 &  x65 &  x80 &  x83 &  x101 &  x107 &  x125 &  x143 &  x146 &  x152 &  x161 &  x188 &  x197 &  x200 &  x215 &  x218 &  x236 &  x239 &  x242 &  x251 &  x254 &  x257 &  x260 &  x263 &  x275 &  x296 &  x305 &  x332 &  x338 &  x359 &  x371 &  x374 &  x389 &  x410 &  x428 &  x443 &  x446 &  x449 &  x470 &  x479 &  x482 &  x491 &  x521 &  x530 &  x551 &  x557 &  x563 &  x581 &  x584 &  x596 &  x608 &  x617 &  x620 &  x626 &  x632 &  x638 &  x641 &  x662 &  x677 &  x683 &  x704 &  x713 &  x716 &  x731 &  x755 &  x764 &  x776 &  x785 &  x794 &  x800 &  x809 &  x812 &  x818 &  x821 &  x836 &  x845 &  x848 &  x857 &  x863 &  x869 &  x875 &  x878 &  x893 &  x911 &  x917 &  x920 &  x923 &  x938 &  x941 &  x983 &  x998 &  x1004 &  x1016 &  x1019 &  x1022 &  x1034 &  x1040 &  x1061 &  x1070 &  x1079 &  x1082 &  x1085 &  x1091 &  x1097 &  x1112 &  x1121 &  x1130 & ~x249 & ~x354 & ~x570 & ~x687 & ~x783 & ~x822 & ~x900 & ~x978;
assign c5241 =  x59 &  x71 &  x131 &  x152 &  x218 &  x335 &  x341 &  x347 &  x350 &  x359 &  x368 &  x377 &  x440 &  x442 &  x443 &  x452 &  x485 &  x515 &  x524 &  x527 &  x542 &  x575 &  x623 &  x635 &  x665 &  x701 &  x706 &  x761 &  x770 &  x779 &  x784 &  x785 &  x821 &  x845 &  x881 &  x890 &  x893 &  x923 &  x962 &  x971 &  x1025 &  x1073 &  x1109 &  x1118 & ~x120 & ~x198 & ~x246 & ~x285 & ~x312 & ~x921;
assign c5243 =  x14 &  x25 &  x52 &  x64 &  x91 &  x182 &  x209 &  x323 &  x401 &  x425 &  x608 &  x722 &  x838 &  x926 &  x971 &  x1027 &  x1070 & ~x357;
assign c5245 =  x20 &  x32 &  x74 &  x77 &  x100 &  x113 &  x152 &  x206 &  x223 &  x242 &  x254 &  x278 &  x317 &  x323 &  x338 &  x356 &  x359 &  x364 &  x400 &  x406 &  x458 &  x554 &  x584 &  x614 &  x698 &  x755 &  x770 &  x779 &  x784 &  x818 &  x890 &  x905 &  x917 &  x971 &  x976 &  x1076 &  x1088 &  x1106 & ~x351;
assign c5247 =  x8 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x47 &  x53 &  x59 &  x65 &  x68 &  x74 &  x80 &  x104 &  x110 &  x116 &  x125 &  x128 &  x158 &  x167 &  x170 &  x173 &  x176 &  x182 &  x194 &  x197 &  x200 &  x203 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x248 &  x257 &  x275 &  x287 &  x290 &  x302 &  x305 &  x311 &  x314 &  x317 &  x323 &  x329 &  x341 &  x353 &  x359 &  x368 &  x380 &  x395 &  x398 &  x401 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x433 &  x437 &  x440 &  x446 &  x455 &  x464 &  x467 &  x472 &  x473 &  x491 &  x494 &  x497 &  x500 &  x503 &  x511 &  x515 &  x518 &  x524 &  x530 &  x533 &  x536 &  x548 &  x557 &  x560 &  x569 &  x578 &  x584 &  x587 &  x589 &  x593 &  x596 &  x599 &  x605 &  x623 &  x626 &  x632 &  x638 &  x647 &  x650 &  x656 &  x665 &  x668 &  x671 &  x689 &  x695 &  x698 &  x701 &  x707 &  x716 &  x719 &  x722 &  x740 &  x749 &  x752 &  x761 &  x767 &  x773 &  x779 &  x788 &  x794 &  x797 &  x803 &  x806 &  x809 &  x812 &  x818 &  x827 &  x836 &  x839 &  x842 &  x860 &  x866 &  x872 &  x875 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x902 &  x905 &  x908 &  x911 &  x917 &  x920 &  x926 &  x929 &  x935 &  x938 &  x953 &  x956 &  x965 &  x977 &  x980 &  x983 &  x989 &  x995 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1043 &  x1046 &  x1055 &  x1064 &  x1070 &  x1073 &  x1094 &  x1100 &  x1103 &  x1112 &  x1124 &  x1127 & ~x273 & ~x312 & ~x537 & ~x576 & ~x615;
assign c5249 =  x44 &  x121 &  x160 & ~x66 & ~x333 & ~x522;
assign c5251 =  x128 &  x187 &  x292 &  x422 &  x488 &  x692 &  x760 &  x794 &  x799 & ~x204 & ~x366 & ~x522;
assign c5253 =  x59 &  x107 &  x200 &  x215 &  x239 &  x419 &  x512 &  x605 &  x608 &  x614 &  x632 &  x665 &  x677 &  x686 &  x878 &  x890 &  x1064 &  x1070 &  x1073 & ~x844 & ~x960 & ~x1011 & ~x1050 & ~x1095;
assign c5255 =  x4 &  x14 &  x134 &  x146 &  x188 &  x199 &  x238 &  x281 &  x371 &  x392 &  x422 &  x464 &  x503 &  x506 &  x641 &  x644 &  x662 &  x689 &  x707 &  x721 &  x734 &  x743 &  x746 &  x760 &  x773 &  x863 &  x875 &  x908 &  x965 &  x989 &  x1034 &  x1067 &  x1088 &  x1097 & ~x414 & ~x663 & ~x741;
assign c5257 =  x5 &  x74 &  x86 &  x104 &  x167 &  x179 &  x191 &  x200 &  x206 &  x239 &  x245 &  x365 &  x374 &  x433 &  x472 &  x485 &  x530 &  x569 &  x589 &  x625 &  x628 &  x647 &  x653 &  x665 &  x707 &  x710 &  x731 &  x743 &  x788 &  x806 &  x822 &  x869 &  x932 &  x953 &  x1034 &  x1046 &  x1115;
assign c5259 =  x5 &  x20 &  x32 &  x38 &  x50 &  x62 &  x68 &  x74 &  x92 &  x98 &  x119 &  x125 &  x131 &  x134 &  x146 &  x149 &  x173 &  x176 &  x185 &  x188 &  x224 &  x233 &  x236 &  x272 &  x281 &  x284 &  x304 &  x311 &  x314 &  x317 &  x329 &  x332 &  x374 &  x383 &  x392 &  x407 &  x415 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x448 &  x452 &  x454 &  x461 &  x473 &  x476 &  x479 &  x488 &  x493 &  x494 &  x497 &  x521 &  x527 &  x539 &  x545 &  x548 &  x551 &  x557 &  x563 &  x566 &  x584 &  x587 &  x590 &  x593 &  x599 &  x602 &  x611 &  x620 &  x623 &  x632 &  x644 &  x647 &  x656 &  x674 &  x680 &  x686 &  x689 &  x701 &  x704 &  x713 &  x745 &  x749 &  x752 &  x758 &  x764 &  x788 &  x794 &  x800 &  x806 &  x821 &  x827 &  x833 &  x836 &  x839 &  x854 &  x875 &  x878 &  x884 &  x887 &  x893 &  x905 &  x914 &  x917 &  x935 &  x941 &  x950 &  x977 &  x980 &  x983 &  x989 &  x995 &  x1004 &  x1013 &  x1016 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1061 &  x1070 &  x1073 &  x1085 &  x1106 &  x1112 &  x1127 & ~x156 & ~x391 & ~x429 & ~x430 & ~x468 & ~x469 & ~x507 & ~x540 & ~x546;
assign c5261 =  x43 &  x121 &  x260 &  x326 &  x383 &  x419 &  x749 &  x883 &  x917 &  x922 &  x1040 &  x1091 & ~x294 & ~x702 & ~x858 & ~x975;
assign c5263 =  x131 &  x181 &  x221 &  x287 &  x316 &  x355 &  x394 &  x472 &  x536 &  x589 &  x627 &  x671 &  x686 &  x908 &  x917 &  x1013;
assign c5265 =  x2 &  x20 &  x32 &  x35 &  x77 &  x86 &  x137 &  x155 &  x176 &  x194 &  x209 &  x221 &  x224 &  x242 &  x251 &  x266 &  x287 &  x296 &  x323 &  x338 &  x353 &  x371 &  x386 &  x389 &  x416 &  x440 &  x458 &  x464 &  x467 &  x482 &  x497 &  x503 &  x506 &  x530 &  x533 &  x551 &  x560 &  x563 &  x587 &  x596 &  x608 &  x611 &  x617 &  x620 &  x638 &  x668 &  x671 &  x713 &  x725 &  x746 &  x764 &  x773 &  x788 &  x818 &  x821 &  x824 &  x836 &  x839 &  x848 &  x863 &  x866 &  x884 &  x887 &  x890 &  x896 &  x902 &  x923 &  x935 &  x941 &  x944 &  x952 &  x959 &  x962 &  x989 &  x1025 &  x1040 &  x1043 &  x1067 &  x1073 &  x1094 &  x1109 &  x1124 & ~x84 & ~x123 & ~x177 & ~x255 & ~x588;
assign c5267 =  x53 &  x86 &  x122 &  x137 &  x161 &  x236 &  x263 &  x278 &  x290 &  x293 &  x302 &  x362 &  x464 &  x467 &  x602 &  x623 &  x653 &  x674 &  x679 &  x686 &  x701 &  x713 &  x743 &  x758 &  x764 &  x803 &  x824 &  x854 &  x857 &  x875 &  x887 &  x890 &  x893 &  x941 &  x944 &  x953 &  x959 &  x977 &  x980 &  x1019 &  x1049 & ~x378 & ~x379 & ~x418;
assign c5269 =  x11 &  x71 &  x116 &  x209 &  x296 &  x356 &  x464 &  x635 &  x785 &  x848 &  x956 &  x1055 & ~x378 & ~x573 & ~x652 & ~x730 & ~x808 & ~x885;
assign c5271 =  x14 &  x43 &  x44 &  x82 &  x86 &  x104 &  x107 &  x110 &  x134 &  x137 &  x140 &  x149 &  x155 &  x156 &  x161 &  x191 &  x248 &  x287 &  x299 &  x365 &  x425 &  x452 &  x461 &  x476 &  x503 &  x518 &  x524 &  x530 &  x545 &  x554 &  x557 &  x563 &  x575 &  x608 &  x617 &  x632 &  x638 &  x659 &  x662 &  x680 &  x692 &  x695 &  x701 &  x704 &  x716 &  x725 &  x749 &  x755 &  x764 &  x776 &  x794 &  x803 &  x884 &  x893 &  x899 &  x932 &  x950 &  x959 &  x968 &  x983 &  x1013 &  x1040 &  x1055 &  x1070 &  x1118 & ~x84 & ~x123 & ~x258 & ~x783;
assign c5273 =  x35 &  x191 &  x224 &  x269 &  x299 &  x314 &  x374 &  x407 &  x425 &  x443 &  x485 &  x488 &  x500 &  x506 &  x526 &  x548 &  x745 &  x770 &  x773 &  x784 &  x902 &  x962 &  x1061 & ~x469 & ~x507 & ~x547 & ~x843;
assign c5275 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x29 &  x41 &  x53 &  x56 &  x65 &  x68 &  x71 &  x80 &  x83 &  x86 &  x95 &  x98 &  x104 &  x116 &  x125 &  x128 &  x134 &  x140 &  x146 &  x161 &  x164 &  x176 &  x185 &  x188 &  x203 &  x206 &  x209 &  x212 &  x218 &  x221 &  x233 &  x248 &  x251 &  x272 &  x275 &  x284 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x314 &  x320 &  x326 &  x335 &  x338 &  x347 &  x350 &  x353 &  x362 &  x368 &  x374 &  x377 &  x380 &  x386 &  x389 &  x404 &  x410 &  x413 &  x416 &  x419 &  x422 &  x431 &  x434 &  x440 &  x443 &  x449 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x485 &  x488 &  x497 &  x521 &  x527 &  x548 &  x551 &  x554 &  x560 &  x572 &  x581 &  x587 &  x590 &  x602 &  x620 &  x623 &  x626 &  x632 &  x635 &  x638 &  x641 &  x647 &  x653 &  x656 &  x674 &  x680 &  x683 &  x686 &  x689 &  x695 &  x698 &  x710 &  x719 &  x722 &  x725 &  x728 &  x734 &  x740 &  x743 &  x755 &  x758 &  x761 &  x764 &  x767 &  x779 &  x782 &  x788 &  x797 &  x806 &  x809 &  x812 &  x824 &  x827 &  x830 &  x836 &  x842 &  x845 &  x854 &  x860 &  x863 &  x866 &  x869 &  x874 &  x875 &  x884 &  x890 &  x899 &  x902 &  x905 &  x911 &  x917 &  x920 &  x923 &  x926 &  x941 &  x952 &  x962 &  x989 &  x992 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1034 &  x1037 &  x1046 &  x1049 &  x1058 &  x1064 &  x1070 &  x1088 &  x1097 &  x1103 &  x1106 &  x1109 &  x1115 & ~x354 & ~x393 & ~x432 & ~x570 & ~x726 & ~x765 & ~x1056;
assign c5277 =  x11 &  x104 &  x187 &  x245 &  x275 &  x332 &  x476 &  x479 &  x545 &  x565 &  x635 &  x779 &  x791 &  x812 &  x887 & ~x396 & ~x435 & ~x513 & ~x594 & ~x1008;
assign c5279 =  x17 &  x116 &  x173 &  x239 &  x242 &  x251 &  x287 &  x376 &  x415 &  x431 &  x448 &  x454 &  x481 &  x623 &  x659 &  x677 &  x704 &  x745 &  x823 &  x869 &  x929 &  x950 &  x959 &  x1076 &  x1115 &  x1118 & ~x273 & ~x429 & ~x618 & ~x1077;
assign c5281 =  x32 &  x89 &  x116 &  x128 &  x145 &  x158 &  x215 &  x224 &  x227 &  x242 &  x281 &  x293 &  x295 &  x341 &  x376 &  x403 &  x422 &  x443 &  x458 &  x497 &  x536 &  x554 &  x644 &  x689 &  x710 &  x713 &  x749 &  x767 &  x866 &  x893 &  x902 &  x926 &  x935 &  x983 &  x1079 & ~x81 & ~x120 & ~x276 & ~x312 & ~x354 & ~x1050;
assign c5283 =  x101 &  x325 &  x406 &  x480 &  x871 &  x949;
assign c5285 =  x2 &  x359 &  x497 &  x589 &  x664 & ~x429 & ~x1077;
assign c5287 =  x26 &  x89 &  x95 &  x113 &  x128 &  x143 &  x152 &  x158 &  x221 &  x224 &  x230 &  x233 &  x239 &  x251 &  x281 &  x314 &  x320 &  x323 &  x344 &  x362 &  x380 &  x404 &  x410 &  x419 &  x427 &  x470 &  x491 &  x494 &  x503 &  x515 &  x524 &  x527 &  x548 &  x590 &  x620 &  x632 &  x644 &  x647 &  x664 &  x683 &  x701 &  x728 &  x731 &  x742 &  x743 &  x746 &  x773 &  x776 &  x779 &  x785 &  x797 &  x803 &  x821 &  x851 &  x863 &  x914 &  x917 &  x926 &  x938 &  x953 &  x968 &  x971 &  x1001 &  x1055 &  x1067 &  x1079 & ~x648 & ~x894 & ~x993 & ~x1050;
assign c5289 =  x2 &  x8 &  x11 &  x26 &  x32 &  x38 &  x41 &  x47 &  x50 &  x53 &  x62 &  x65 &  x68 &  x74 &  x82 &  x86 &  x89 &  x95 &  x98 &  x101 &  x110 &  x113 &  x116 &  x131 &  x146 &  x149 &  x179 &  x188 &  x194 &  x197 &  x199 &  x200 &  x206 &  x209 &  x218 &  x227 &  x242 &  x251 &  x254 &  x257 &  x260 &  x266 &  x269 &  x272 &  x281 &  x284 &  x290 &  x317 &  x323 &  x332 &  x335 &  x344 &  x356 &  x368 &  x374 &  x377 &  x392 &  x407 &  x416 &  x431 &  x437 &  x449 &  x458 &  x464 &  x470 &  x479 &  x491 &  x500 &  x503 &  x509 &  x515 &  x521 &  x524 &  x530 &  x533 &  x536 &  x545 &  x554 &  x560 &  x566 &  x590 &  x593 &  x599 &  x611 &  x620 &  x632 &  x635 &  x638 &  x644 &  x647 &  x656 &  x661 &  x662 &  x674 &  x689 &  x698 &  x725 &  x731 &  x740 &  x746 &  x749 &  x752 &  x761 &  x764 &  x785 &  x794 &  x815 &  x818 &  x821 &  x824 &  x827 &  x836 &  x839 &  x842 &  x850 &  x857 &  x860 &  x884 &  x890 &  x929 &  x938 &  x962 &  x980 &  x986 &  x992 &  x998 &  x1007 &  x1016 &  x1022 &  x1031 &  x1034 &  x1058 &  x1070 &  x1079 &  x1085 &  x1088 &  x1103 &  x1109 &  x1112 &  x1121 & ~x975 & ~x1014;
assign c5291 =  x8 &  x416 &  x781 &  x800 & ~x570 & ~x1057;
assign c5293 =  x50 &  x70 &  x77 &  x119 &  x176 &  x251 &  x277 &  x290 &  x620 &  x662 &  x686 &  x719 &  x728 &  x974 &  x1037 &  x1103 &  x1127 & ~x387 & ~x408 & ~x531;
assign c5295 =  x17 &  x23 &  x62 &  x80 &  x134 &  x154 &  x215 &  x226 &  x248 &  x272 &  x311 &  x323 &  x329 &  x362 &  x433 &  x443 &  x476 &  x569 &  x589 &  x617 &  x629 &  x664 &  x704 &  x725 &  x781 &  x820 &  x845 &  x884 &  x902 &  x905 &  x917 &  x932 &  x959 &  x986 &  x989 &  x1058;
assign c5297 =  x11 &  x41 &  x50 &  x64 &  x65 &  x71 &  x86 &  x91 &  x119 &  x128 &  x182 &  x188 &  x191 &  x209 &  x239 &  x254 &  x263 &  x266 &  x269 &  x277 &  x278 &  x281 &  x316 &  x368 &  x389 &  x413 &  x419 &  x425 &  x433 &  x446 &  x449 &  x473 &  x497 &  x509 &  x518 &  x533 &  x536 &  x554 &  x560 &  x566 &  x611 &  x614 &  x644 &  x719 &  x752 &  x758 &  x788 &  x794 &  x818 &  x833 &  x851 &  x875 &  x905 &  x932 &  x938 &  x949 &  x953 &  x971 &  x989 &  x1004 &  x1076 &  x1094 &  x1109 &  x1118;
assign c5299 =  x62 &  x77 &  x95 &  x107 &  x110 &  x125 &  x143 &  x164 &  x173 &  x209 &  x212 &  x218 &  x239 &  x251 &  x257 &  x290 &  x302 &  x316 &  x317 &  x326 &  x344 &  x350 &  x368 &  x371 &  x398 &  x407 &  x413 &  x419 &  x425 &  x443 &  x446 &  x464 &  x482 &  x500 &  x515 &  x524 &  x545 &  x554 &  x560 &  x575 &  x590 &  x593 &  x626 &  x629 &  x638 &  x647 &  x659 &  x674 &  x701 &  x707 &  x719 &  x722 &  x725 &  x728 &  x734 &  x737 &  x746 &  x764 &  x773 &  x788 &  x821 &  x830 &  x836 &  x863 &  x875 &  x878 &  x890 &  x896 &  x923 &  x947 &  x977 &  x1007 &  x1043 &  x1046 &  x1049 &  x1055 &  x1076 &  x1109 &  x1115 &  x1121 & ~x39 & ~x117 & ~x435 & ~x1092;
assign c60 =  x2 &  x5 &  x8 &  x11 &  x20 &  x26 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x125 &  x131 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x206 &  x212 &  x218 &  x221 &  x227 &  x230 &  x233 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x377 &  x380 &  x386 &  x388 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x427 &  x428 &  x431 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x466 &  x470 &  x473 &  x476 &  x479 &  x485 &  x488 &  x491 &  x497 &  x503 &  x506 &  x509 &  x512 &  x518 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x740 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x977 &  x980 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1013 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 &  x1130 & ~x438 & ~x477 & ~x516 & ~x519 & ~x552 & ~x555 & ~x591 & ~x630 & ~x633 & ~x669 & ~x792 & ~x981 & ~x1020 & ~x1059;
assign c62 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x532 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x571 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x610 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x649 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x688 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x716 &  x719 &  x722 &  x727 &  x728 &  x731 &  x734 &  x737 &  x740 &  x742 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x785 &  x788 &  x790 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x901 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x940 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1018 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x507 & ~x771 & ~x849 & ~x1005;
assign c64 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x119 &  x122 &  x125 &  x131 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x349 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x388 &  x392 &  x395 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x479 &  x482 &  x485 &  x491 &  x494 &  x497 &  x500 &  x503 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x632 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x722 &  x725 &  x728 &  x731 &  x734 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x767 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x863 &  x866 &  x872 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 &  x1130 & ~x195 & ~x273 & ~x312 & ~x351 & ~x444 & ~x483 & ~x484 & ~x522 & ~x523 & ~x561 & ~x562 & ~x601 & ~x603 & ~x639 & ~x678;
assign c66 =  x5 &  x7 &  x8 &  x11 &  x14 &  x17 &  x20 &  x32 &  x35 &  x38 &  x41 &  x44 &  x46 &  x47 &  x50 &  x53 &  x56 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x85 &  x86 &  x89 &  x92 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x124 &  x128 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x161 &  x163 &  x164 &  x167 &  x170 &  x176 &  x181 &  x182 &  x185 &  x188 &  x191 &  x197 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x220 &  x221 &  x230 &  x239 &  x241 &  x242 &  x245 &  x251 &  x254 &  x257 &  x259 &  x260 &  x265 &  x266 &  x272 &  x275 &  x278 &  x280 &  x284 &  x287 &  x290 &  x293 &  x296 &  x298 &  x302 &  x305 &  x308 &  x311 &  x317 &  x319 &  x320 &  x323 &  x329 &  x335 &  x337 &  x344 &  x347 &  x349 &  x350 &  x353 &  x356 &  x362 &  x368 &  x371 &  x374 &  x376 &  x377 &  x380 &  x383 &  x386 &  x388 &  x392 &  x395 &  x404 &  x415 &  x416 &  x419 &  x422 &  x425 &  x427 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x449 &  x454 &  x458 &  x461 &  x466 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x493 &  x494 &  x500 &  x503 &  x506 &  x518 &  x521 &  x530 &  x536 &  x545 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x572 &  x578 &  x584 &  x587 &  x593 &  x596 &  x602 &  x608 &  x614 &  x623 &  x626 &  x629 &  x632 &  x638 &  x641 &  x644 &  x647 &  x649 &  x653 &  x656 &  x659 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x722 &  x725 &  x727 &  x728 &  x734 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x761 &  x764 &  x766 &  x767 &  x773 &  x779 &  x782 &  x791 &  x794 &  x797 &  x803 &  x809 &  x812 &  x815 &  x821 &  x824 &  x827 &  x830 &  x836 &  x842 &  x845 &  x854 &  x857 &  x863 &  x866 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x914 &  x923 &  x926 &  x929 &  x932 &  x938 &  x941 &  x947 &  x950 &  x959 &  x968 &  x971 &  x974 &  x977 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1016 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1049 &  x1052 &  x1058 &  x1061 &  x1067 &  x1073 &  x1076 &  x1082 &  x1085 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x312 & ~x717;
assign c68 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x34 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x73 &  x74 &  x77 &  x80 &  x82 &  x83 &  x89 &  x92 &  x95 &  x101 &  x104 &  x107 &  x110 &  x112 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x155 &  x158 &  x161 &  x167 &  x170 &  x173 &  x179 &  x182 &  x185 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x260 &  x263 &  x266 &  x268 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x299 &  x302 &  x305 &  x307 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x332 &  x335 &  x341 &  x344 &  x346 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x413 &  x415 &  x416 &  x419 &  x422 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x454 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x479 &  x482 &  x485 &  x488 &  x491 &  x493 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x521 &  x524 &  x527 &  x530 &  x532 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x571 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x610 &  x611 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x649 &  x653 &  x656 &  x659 &  x662 &  x668 &  x674 &  x680 &  x682 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x713 &  x716 &  x719 &  x721 &  x722 &  x725 &  x727 &  x728 &  x731 &  x733 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x760 &  x761 &  x764 &  x766 &  x767 &  x770 &  x772 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x827 &  x830 &  x836 &  x842 &  x845 &  x848 &  x851 &  x853 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x890 &  x896 &  x899 &  x902 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x977 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1007 &  x1013 &  x1016 &  x1019 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x858 & ~x897;
assign c610 =  x2 &  x5 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x176 &  x179 &  x182 &  x185 &  x188 &  x194 &  x197 &  x203 &  x209 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x329 &  x332 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x376 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x397 &  x398 &  x401 &  x404 &  x413 &  x415 &  x416 &  x419 &  x422 &  x428 &  x431 &  x434 &  x436 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x460 &  x461 &  x464 &  x467 &  x473 &  x476 &  x482 &  x485 &  x487 &  x488 &  x491 &  x493 &  x494 &  x497 &  x499 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x526 &  x527 &  x530 &  x533 &  x538 &  x539 &  x542 &  x544 &  x545 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x572 &  x575 &  x581 &  x583 &  x584 &  x587 &  x593 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x622 &  x629 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x725 &  x731 &  x734 &  x737 &  x740 &  x749 &  x752 &  x755 &  x758 &  x767 &  x773 &  x779 &  x782 &  x785 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x824 &  x830 &  x833 &  x836 &  x839 &  x845 &  x848 &  x854 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x944 &  x947 &  x953 &  x956 &  x959 &  x962 &  x965 &  x971 &  x974 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1058 &  x1061 &  x1064 &  x1076 &  x1079 &  x1082 &  x1085 &  x1094 &  x1096 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x312 & ~x351 & ~x390 & ~x429 & ~x432 & ~x468 & ~x471 & ~x510 & ~x549 & ~x753 & ~x792 & ~x834 & ~x948 & ~x987 & ~x1026 & ~x1104;
assign c612 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x292 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x934 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1111 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x273 & ~x282 & ~x312 & ~x321 & ~x483 & ~x936 & ~x975;
assign c614 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x22 &  x23 &  x26 &  x32 &  x35 &  x38 &  x40 &  x41 &  x44 &  x50 &  x56 &  x59 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x100 &  x104 &  x110 &  x113 &  x116 &  x118 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x139 &  x140 &  x143 &  x146 &  x152 &  x155 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x212 &  x217 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x242 &  x245 &  x248 &  x251 &  x257 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x293 &  x299 &  x302 &  x305 &  x314 &  x317 &  x320 &  x323 &  x326 &  x335 &  x341 &  x344 &  x356 &  x359 &  x362 &  x374 &  x377 &  x380 &  x383 &  x385 &  x386 &  x392 &  x404 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x437 &  x440 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x467 &  x473 &  x476 &  x479 &  x482 &  x485 &  x491 &  x497 &  x500 &  x502 &  x506 &  x515 &  x518 &  x521 &  x524 &  x530 &  x533 &  x536 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x587 &  x590 &  x596 &  x602 &  x605 &  x611 &  x620 &  x623 &  x632 &  x635 &  x644 &  x653 &  x658 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x680 &  x686 &  x688 &  x689 &  x692 &  x698 &  x701 &  x704 &  x707 &  x710 &  x719 &  x725 &  x728 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x775 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x809 &  x812 &  x814 &  x815 &  x818 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x841 &  x842 &  x845 &  x848 &  x851 &  x854 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x896 &  x899 &  x905 &  x908 &  x911 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x971 &  x974 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1037 &  x1043 &  x1046 &  x1049 &  x1055 &  x1061 &  x1064 &  x1070 &  x1076 &  x1082 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x252 & ~x282 & ~x285 & ~x336 & ~x375 & ~x441;
assign c616 =  x5 &  x8 &  x11 &  x17 &  x23 &  x41 &  x53 &  x56 &  x68 &  x76 &  x80 &  x83 &  x86 &  x98 &  x104 &  x110 &  x119 &  x125 &  x131 &  x137 &  x143 &  x146 &  x158 &  x161 &  x179 &  x182 &  x185 &  x194 &  x197 &  x200 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x239 &  x251 &  x254 &  x260 &  x263 &  x269 &  x293 &  x296 &  x311 &  x317 &  x320 &  x332 &  x338 &  x341 &  x344 &  x350 &  x359 &  x362 &  x365 &  x368 &  x374 &  x380 &  x386 &  x395 &  x404 &  x407 &  x410 &  x413 &  x428 &  x440 &  x443 &  x464 &  x467 &  x470 &  x473 &  x482 &  x485 &  x494 &  x500 &  x512 &  x518 &  x521 &  x524 &  x539 &  x542 &  x545 &  x548 &  x557 &  x569 &  x581 &  x590 &  x596 &  x599 &  x602 &  x608 &  x611 &  x617 &  x623 &  x629 &  x638 &  x644 &  x647 &  x650 &  x653 &  x668 &  x674 &  x677 &  x680 &  x683 &  x689 &  x695 &  x698 &  x701 &  x719 &  x722 &  x725 &  x728 &  x734 &  x755 &  x761 &  x764 &  x773 &  x776 &  x779 &  x782 &  x788 &  x791 &  x800 &  x803 &  x805 &  x809 &  x815 &  x821 &  x826 &  x842 &  x845 &  x848 &  x851 &  x857 &  x863 &  x865 &  x866 &  x869 &  x872 &  x875 &  x878 &  x883 &  x884 &  x893 &  x902 &  x920 &  x926 &  x932 &  x935 &  x938 &  x941 &  x947 &  x955 &  x961 &  x965 &  x980 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1016 &  x1019 &  x1022 &  x1025 &  x1027 &  x1031 &  x1037 &  x1043 &  x1051 &  x1058 &  x1064 &  x1067 &  x1082 &  x1085 &  x1088 &  x1090 &  x1091 &  x1094 &  x1097 &  x1100 &  x1109 &  x1115 &  x1121 &  x1127 &  x1130 & ~x327 & ~x444 & ~x483 & ~x549;
assign c618 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x56 &  x62 &  x65 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x263 &  x266 &  x269 &  x272 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x379 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x674 &  x677 &  x680 &  x683 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x827 &  x830 &  x833 &  x841 &  x842 &  x845 &  x848 &  x851 &  x854 &  x856 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x880 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x934 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x6 & ~x480 & ~x483 & ~x486 & ~x522 & ~x525;
assign c620 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x25 &  x26 &  x29 &  x32 &  x38 &  x50 &  x53 &  x56 &  x62 &  x64 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x95 &  x98 &  x101 &  x103 &  x104 &  x110 &  x113 &  x119 &  x122 &  x125 &  x128 &  x134 &  x140 &  x143 &  x149 &  x152 &  x155 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x230 &  x233 &  x239 &  x242 &  x245 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x350 &  x353 &  x359 &  x368 &  x371 &  x380 &  x386 &  x389 &  x392 &  x395 &  x401 &  x404 &  x407 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x446 &  x449 &  x455 &  x461 &  x470 &  x476 &  x485 &  x488 &  x491 &  x497 &  x503 &  x506 &  x509 &  x512 &  x515 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x545 &  x548 &  x551 &  x554 &  x560 &  x563 &  x566 &  x569 &  x575 &  x578 &  x581 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x794 &  x797 &  x800 &  x803 &  x809 &  x812 &  x815 &  x821 &  x824 &  x827 &  x830 &  x836 &  x838 &  x839 &  x842 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x875 &  x887 &  x890 &  x896 &  x902 &  x905 &  x908 &  x914 &  x916 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x980 &  x983 &  x986 &  x989 &  x994 &  x995 &  x998 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1033 &  x1034 &  x1037 &  x1039 &  x1040 &  x1043 &  x1046 &  x1049 &  x1051 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1078 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1109 &  x1117 &  x1118 &  x1130 & ~x246 & ~x285 & ~x477 & ~x780 & ~x897;
assign c622 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x80 &  x83 &  x86 &  x89 &  x95 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x209 &  x212 &  x218 &  x221 &  x224 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x464 &  x467 &  x470 &  x473 &  x476 &  x482 &  x485 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x515 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x599 &  x605 &  x614 &  x617 &  x620 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x857 &  x860 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x273 & ~x312 & ~x315 & ~x351 & ~x354 & ~x393 & ~x399 & ~x432 & ~x438 & ~x477 & ~x516 & ~x636 & ~x637 & ~x675 & ~x676 & ~x678 & ~x714 & ~x717 & ~x753 & ~x756 & ~x792 & ~x831;
assign c624 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x83 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x262 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x454 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x532 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x683 &  x686 &  x689 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x776 &  x779 &  x782 &  x785 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x812 &  x815 &  x818 &  x821 &  x823 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x941 &  x944 &  x947 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x977 &  x979 &  x980 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1018 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1096 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x360 & ~x399 & ~x438 & ~x477 & ~x546 & ~x756 & ~x759 & ~x795 & ~x798 & ~x837 & ~x876 & ~x915;
assign c626 =  x2 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x68 &  x71 &  x77 &  x80 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x185 &  x188 &  x194 &  x197 &  x200 &  x206 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x239 &  x242 &  x245 &  x248 &  x251 &  x257 &  x263 &  x266 &  x269 &  x275 &  x278 &  x287 &  x290 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x320 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x355 &  x356 &  x359 &  x368 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x446 &  x452 &  x455 &  x458 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x566 &  x569 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x632 &  x635 &  x638 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x674 &  x680 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x761 &  x764 &  x767 &  x773 &  x776 &  x782 &  x785 &  x788 &  x791 &  x794 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x832 &  x836 &  x839 &  x842 &  x845 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x929 &  x938 &  x941 &  x944 &  x950 &  x953 &  x959 &  x962 &  x965 &  x968 &  x977 &  x980 &  x983 &  x986 &  x988 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1037 &  x1040 &  x1043 &  x1045 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1097 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x249 & ~x288 & ~x363 & ~x402 & ~x441 & ~x483 & ~x522 & ~x624 & ~x666 & ~x702 & ~x705 & ~x741 & ~x744 & ~x780 & ~x783 & ~x822 & ~x858 & ~x897 & ~x1014 & ~x1053;
assign c628 =  x2 &  x8 &  x14 &  x26 &  x35 &  x38 &  x41 &  x47 &  x50 &  x62 &  x68 &  x71 &  x77 &  x79 &  x80 &  x112 &  x113 &  x119 &  x128 &  x131 &  x137 &  x139 &  x152 &  x155 &  x157 &  x164 &  x179 &  x197 &  x200 &  x203 &  x218 &  x224 &  x230 &  x236 &  x242 &  x251 &  x254 &  x260 &  x263 &  x269 &  x272 &  x281 &  x293 &  x299 &  x305 &  x311 &  x314 &  x317 &  x323 &  x326 &  x341 &  x344 &  x350 &  x368 &  x371 &  x374 &  x386 &  x395 &  x404 &  x410 &  x413 &  x416 &  x424 &  x428 &  x431 &  x449 &  x476 &  x485 &  x488 &  x491 &  x518 &  x548 &  x554 &  x557 &  x560 &  x571 &  x587 &  x608 &  x614 &  x626 &  x635 &  x647 &  x650 &  x656 &  x674 &  x689 &  x692 &  x698 &  x704 &  x710 &  x716 &  x728 &  x731 &  x734 &  x755 &  x767 &  x769 &  x773 &  x785 &  x794 &  x809 &  x836 &  x842 &  x854 &  x860 &  x863 &  x866 &  x875 &  x878 &  x908 &  x941 &  x944 &  x965 &  x974 &  x980 &  x1010 &  x1025 &  x1043 &  x1049 &  x1052 &  x1055 &  x1067 &  x1082 &  x1097 &  x1100 &  x1103 &  x1106 &  x1118 & ~x12 & ~x285 & ~x363 & ~x402 & ~x864 & ~x1020 & ~x1059 & ~x1071 & ~x1098 & ~x1104;
assign c630 =  x4 &  x8 &  x11 &  x26 &  x32 &  x35 &  x38 &  x41 &  x47 &  x50 &  x53 &  x59 &  x77 &  x80 &  x83 &  x89 &  x92 &  x95 &  x98 &  x100 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x137 &  x139 &  x140 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x176 &  x178 &  x179 &  x182 &  x185 &  x191 &  x200 &  x203 &  x212 &  x215 &  x217 &  x218 &  x227 &  x236 &  x239 &  x242 &  x245 &  x251 &  x257 &  x260 &  x263 &  x266 &  x278 &  x284 &  x287 &  x295 &  x299 &  x302 &  x314 &  x317 &  x323 &  x334 &  x335 &  x341 &  x344 &  x350 &  x359 &  x362 &  x371 &  x372 &  x373 &  x380 &  x386 &  x389 &  x392 &  x398 &  x404 &  x407 &  x412 &  x416 &  x419 &  x422 &  x425 &  x431 &  x437 &  x440 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x463 &  x476 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x512 &  x515 &  x518 &  x527 &  x530 &  x536 &  x542 &  x548 &  x551 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x605 &  x611 &  x617 &  x623 &  x626 &  x632 &  x641 &  x644 &  x647 &  x650 &  x653 &  x662 &  x665 &  x668 &  x671 &  x674 &  x680 &  x683 &  x692 &  x695 &  x698 &  x701 &  x710 &  x719 &  x724 &  x725 &  x737 &  x740 &  x743 &  x749 &  x752 &  x763 &  x767 &  x776 &  x779 &  x802 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x827 &  x830 &  x833 &  x842 &  x845 &  x854 &  x857 &  x869 &  x872 &  x883 &  x884 &  x886 &  x899 &  x905 &  x914 &  x923 &  x926 &  x929 &  x932 &  x944 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x980 &  x986 &  x995 &  x998 &  x1001 &  x1007 &  x1019 &  x1022 &  x1037 &  x1043 &  x1049 &  x1055 &  x1058 &  x1064 &  x1067 &  x1073 &  x1078 &  x1079 &  x1085 &  x1091 &  x1094 &  x1100 &  x1112 &  x1121 &  x1127;
assign c632 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x35 &  x38 &  x41 &  x44 &  x47 &  x59 &  x62 &  x65 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x104 &  x110 &  x113 &  x119 &  x122 &  x125 &  x128 &  x131 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x164 &  x173 &  x176 &  x182 &  x185 &  x191 &  x197 &  x200 &  x203 &  x209 &  x212 &  x215 &  x224 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x263 &  x266 &  x269 &  x278 &  x281 &  x284 &  x287 &  x290 &  x296 &  x314 &  x317 &  x320 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x365 &  x368 &  x374 &  x377 &  x383 &  x386 &  x389 &  x392 &  x401 &  x404 &  x407 &  x413 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x446 &  x449 &  x452 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x485 &  x488 &  x491 &  x494 &  x497 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x806 &  x809 &  x815 &  x818 &  x821 &  x824 &  x830 &  x833 &  x836 &  x848 &  x851 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x902 &  x905 &  x908 &  x914 &  x923 &  x929 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x968 &  x971 &  x979 &  x983 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1052 &  x1055 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1088 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x555 & ~x594 & ~x633 & ~x765 & ~x792 & ~x960 & ~x999 & ~x1000 & ~x1020 & ~x1038 & ~x1059;
assign c634 =  x2 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x206 &  x209 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x254 &  x257 &  x260 &  x263 &  x269 &  x272 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x317 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x377 &  x383 &  x386 &  x389 &  x392 &  x401 &  x407 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x434 &  x437 &  x440 &  x443 &  x449 &  x452 &  x455 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x487 &  x491 &  x493 &  x494 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x553 &  x554 &  x557 &  x566 &  x571 &  x572 &  x575 &  x578 &  x581 &  x583 &  x587 &  x592 &  x596 &  x599 &  x602 &  x608 &  x610 &  x611 &  x614 &  x620 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x647 &  x649 &  x650 &  x653 &  x656 &  x661 &  x662 &  x665 &  x668 &  x671 &  x677 &  x680 &  x682 &  x683 &  x686 &  x688 &  x692 &  x698 &  x704 &  x707 &  x710 &  x713 &  x719 &  x725 &  x727 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x788 &  x791 &  x797 &  x800 &  x803 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x839 &  x845 &  x851 &  x854 &  x860 &  x866 &  x869 &  x875 &  x878 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1114 &  x1115 &  x1118 &  x1121 &  x1124 & ~x471 & ~x477 & ~x510 & ~x516 & ~x549 & ~x555 & ~x588 & ~x594 & ~x627 & ~x633 & ~x672;
assign c636 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x43 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x121 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x158 &  x160 &  x161 &  x164 &  x167 &  x170 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x236 &  x238 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x277 &  x278 &  x281 &  x287 &  x290 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x316 &  x317 &  x320 &  x329 &  x347 &  x350 &  x353 &  x355 &  x356 &  x359 &  x371 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x428 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x494 &  x497 &  x503 &  x509 &  x512 &  x518 &  x521 &  x527 &  x530 &  x536 &  x538 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x563 &  x565 &  x566 &  x569 &  x572 &  x575 &  x577 &  x578 &  x581 &  x583 &  x584 &  x587 &  x590 &  x593 &  x599 &  x602 &  x604 &  x605 &  x611 &  x617 &  x620 &  x622 &  x623 &  x626 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x671 &  x674 &  x677 &  x682 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x734 &  x737 &  x740 &  x746 &  x752 &  x758 &  x760 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x785 &  x788 &  x791 &  x794 &  x800 &  x803 &  x809 &  x812 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x838 &  x839 &  x842 &  x845 &  x851 &  x854 &  x857 &  x860 &  x872 &  x875 &  x877 &  x881 &  x884 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x935 &  x941 &  x944 &  x947 &  x953 &  x959 &  x962 &  x968 &  x971 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1012 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1130 & ~x438 & ~x477 & ~x516 & ~x555 & ~x594 & ~x633 & ~x672;
assign c638 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x29 &  x35 &  x41 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x95 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x128 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x164 &  x167 &  x173 &  x176 &  x179 &  x191 &  x194 &  x197 &  x203 &  x209 &  x212 &  x215 &  x218 &  x224 &  x227 &  x232 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x263 &  x272 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x308 &  x317 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x350 &  x353 &  x356 &  x359 &  x362 &  x371 &  x374 &  x380 &  x389 &  x392 &  x394 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x431 &  x433 &  x434 &  x443 &  x446 &  x455 &  x461 &  x467 &  x470 &  x473 &  x476 &  x485 &  x488 &  x491 &  x494 &  x500 &  x506 &  x515 &  x518 &  x521 &  x524 &  x530 &  x533 &  x536 &  x539 &  x545 &  x548 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x632 &  x635 &  x638 &  x641 &  x644 &  x653 &  x656 &  x659 &  x662 &  x680 &  x686 &  x689 &  x692 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x749 &  x752 &  x761 &  x764 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x794 &  x797 &  x799 &  x800 &  x806 &  x812 &  x815 &  x818 &  x821 &  x830 &  x833 &  x836 &  x838 &  x839 &  x842 &  x845 &  x848 &  x851 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x914 &  x917 &  x920 &  x929 &  x932 &  x935 &  x938 &  x941 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x977 &  x980 &  x986 &  x992 &  x995 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130 & ~x210 & ~x363 & ~x441 & ~x519 & ~x633 & ~x672 & ~x741 & ~x780 & ~x858 & ~x897 & ~x1014 & ~x1053;
assign c640 =  x2 &  x5 &  x8 &  x11 &  x13 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x44 &  x50 &  x52 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x91 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x130 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x164 &  x167 &  x169 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x203 &  x206 &  x208 &  x209 &  x212 &  x218 &  x221 &  x227 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x251 &  x254 &  x257 &  x259 &  x260 &  x263 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x298 &  x299 &  x302 &  x305 &  x308 &  x310 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x337 &  x341 &  x344 &  x347 &  x349 &  x350 &  x353 &  x356 &  x359 &  x362 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x388 &  x389 &  x395 &  x401 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x674 &  x677 &  x683 &  x686 &  x689 &  x692 &  x698 &  x701 &  x704 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x752 &  x755 &  x758 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x845 &  x848 &  x857 &  x860 &  x862 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x901 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x932 &  x935 &  x938 &  x940 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x156 & ~x195 & ~x234 & ~x273 & ~x312 & ~x636 & ~x678 & ~x717;
assign c642 =  x2 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x32 &  x35 &  x41 &  x44 &  x47 &  x50 &  x62 &  x65 &  x74 &  x77 &  x86 &  x89 &  x104 &  x107 &  x113 &  x119 &  x122 &  x125 &  x128 &  x134 &  x137 &  x146 &  x149 &  x157 &  x167 &  x173 &  x209 &  x212 &  x215 &  x218 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x257 &  x260 &  x263 &  x269 &  x278 &  x284 &  x290 &  x296 &  x308 &  x314 &  x317 &  x320 &  x329 &  x335 &  x338 &  x341 &  x371 &  x377 &  x380 &  x383 &  x386 &  x392 &  x395 &  x398 &  x410 &  x416 &  x431 &  x434 &  x437 &  x440 &  x446 &  x458 &  x467 &  x470 &  x473 &  x476 &  x479 &  x488 &  x491 &  x497 &  x512 &  x527 &  x536 &  x545 &  x548 &  x554 &  x560 &  x563 &  x569 &  x581 &  x587 &  x593 &  x596 &  x599 &  x602 &  x611 &  x620 &  x626 &  x629 &  x635 &  x638 &  x640 &  x641 &  x643 &  x644 &  x646 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x677 &  x680 &  x682 &  x683 &  x686 &  x689 &  x692 &  x695 &  x701 &  x704 &  x713 &  x716 &  x721 &  x722 &  x725 &  x731 &  x737 &  x746 &  x749 &  x755 &  x757 &  x758 &  x760 &  x767 &  x770 &  x776 &  x782 &  x785 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x832 &  x833 &  x835 &  x842 &  x848 &  x853 &  x854 &  x857 &  x874 &  x877 &  x878 &  x881 &  x884 &  x890 &  x893 &  x899 &  x902 &  x905 &  x911 &  x916 &  x920 &  x928 &  x929 &  x932 &  x938 &  x947 &  x950 &  x956 &  x959 &  x962 &  x965 &  x971 &  x977 &  x983 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1027 &  x1031 &  x1034 &  x1037 &  x1043 &  x1052 &  x1064 &  x1082 &  x1085 &  x1094 &  x1105 &  x1106 &  x1109 &  x1112 &  x1130 & ~x207 & ~x822;
assign c644 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x646 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x273 & ~x312 & ~x351 & ~x405 & ~x444 & ~x483 & ~x522 & ~x561 & ~x600 & ~x639 & ~x640 & ~x678 & ~x717;
assign c646 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x137 &  x140 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x494 &  x497 &  x500 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x695 &  x698 &  x701 &  x704 &  x707 &  x713 &  x716 &  x719 &  x725 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x821 &  x824 &  x827 &  x830 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x210 & ~x288 & ~x402 & ~x435 & ~x441 & ~x474 & ~x480 & ~x519 & ~x558 & ~x597 & ~x636 & ~x675 & ~x678 & ~x714 & ~x717 & ~x792 & ~x795 & ~x831 & ~x834 & ~x903 & ~x942;
assign c648 =  x2 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x35 &  x41 &  x44 &  x47 &  x50 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x131 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x155 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x251 &  x257 &  x263 &  x266 &  x272 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x310 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x353 &  x356 &  x362 &  x365 &  x368 &  x374 &  x377 &  x380 &  x389 &  x392 &  x395 &  x398 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x427 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x466 &  x467 &  x470 &  x476 &  x482 &  x488 &  x494 &  x497 &  x500 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x548 &  x551 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x578 &  x587 &  x593 &  x605 &  x608 &  x611 &  x617 &  x620 &  x623 &  x626 &  x632 &  x635 &  x638 &  x641 &  x647 &  x650 &  x653 &  x656 &  x662 &  x665 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x713 &  x716 &  x719 &  x722 &  x725 &  x734 &  x737 &  x746 &  x752 &  x755 &  x758 &  x761 &  x767 &  x770 &  x773 &  x779 &  x782 &  x785 &  x788 &  x794 &  x797 &  x800 &  x803 &  x809 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x869 &  x875 &  x878 &  x881 &  x884 &  x887 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x926 &  x932 &  x938 &  x944 &  x947 &  x950 &  x953 &  x956 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x995 &  x998 &  x1004 &  x1010 &  x1013 &  x1016 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1094 &  x1097 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130 & ~x54 & ~x93 & ~x132 & ~x171 & ~x306 & ~x327 & ~x366 & ~x444 & ~x483 & ~x561 & ~x756 & ~x795 & ~x969 & ~x1125;
assign c650 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x191 &  x194 &  x197 &  x200 &  x203 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x269 &  x272 &  x275 &  x277 &  x278 &  x283 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x305 &  x308 &  x311 &  x314 &  x316 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x353 &  x355 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x610 &  x611 &  x614 &  x617 &  x620 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x890 &  x893 &  x896 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x132 & ~x507 & ~x546 & ~x549 & ~x585 & ~x588 & ~x618 & ~x627 & ~x657 & ~x666 & ~x696 & ~x702 & ~x705 & ~x735 & ~x744 & ~x783 & ~x822 & ~x861;
assign c652 =  x2 &  x8 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x131 &  x134 &  x137 &  x140 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x233 &  x236 &  x245 &  x248 &  x254 &  x263 &  x266 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x314 &  x317 &  x323 &  x329 &  x335 &  x338 &  x341 &  x347 &  x350 &  x353 &  x356 &  x365 &  x368 &  x371 &  x377 &  x383 &  x386 &  x389 &  x392 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x515 &  x518 &  x521 &  x524 &  x533 &  x536 &  x539 &  x542 &  x545 &  x551 &  x554 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x587 &  x590 &  x593 &  x599 &  x605 &  x611 &  x614 &  x620 &  x623 &  x626 &  x629 &  x632 &  x638 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x668 &  x671 &  x677 &  x680 &  x683 &  x689 &  x695 &  x698 &  x704 &  x707 &  x713 &  x716 &  x719 &  x722 &  x728 &  x731 &  x734 &  x740 &  x743 &  x746 &  x749 &  x758 &  x770 &  x773 &  x776 &  x782 &  x788 &  x791 &  x797 &  x800 &  x803 &  x812 &  x815 &  x821 &  x827 &  x830 &  x833 &  x836 &  x839 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x953 &  x956 &  x959 &  x962 &  x965 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x998 &  x1004 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1100 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x108 & ~x147 & ~x186 & ~x237 & ~x315 & ~x480 & ~x513 & ~x519 & ~x552 & ~x597 & ~x870 & ~x1065 & ~x1080;
assign c654 =  x2 &  x11 &  x14 &  x17 &  x20 &  x26 &  x29 &  x35 &  x38 &  x41 &  x44 &  x47 &  x53 &  x59 &  x62 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x98 &  x101 &  x104 &  x107 &  x110 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x188 &  x191 &  x194 &  x197 &  x200 &  x206 &  x209 &  x212 &  x215 &  x217 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x256 &  x257 &  x260 &  x263 &  x266 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x293 &  x295 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x322 &  x323 &  x328 &  x329 &  x335 &  x338 &  x344 &  x350 &  x353 &  x356 &  x365 &  x368 &  x371 &  x376 &  x377 &  x380 &  x386 &  x389 &  x392 &  x395 &  x398 &  x400 &  x401 &  x404 &  x407 &  x410 &  x413 &  x415 &  x416 &  x419 &  x421 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x439 &  x443 &  x446 &  x449 &  x452 &  x454 &  x455 &  x458 &  x460 &  x461 &  x467 &  x470 &  x473 &  x478 &  x479 &  x485 &  x488 &  x491 &  x494 &  x497 &  x499 &  x500 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x530 &  x536 &  x539 &  x542 &  x545 &  x548 &  x554 &  x560 &  x563 &  x566 &  x572 &  x575 &  x578 &  x584 &  x587 &  x590 &  x596 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x677 &  x680 &  x683 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x734 &  x737 &  x740 &  x743 &  x749 &  x752 &  x758 &  x761 &  x770 &  x773 &  x779 &  x782 &  x785 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x818 &  x821 &  x827 &  x830 &  x839 &  x842 &  x845 &  x848 &  x857 &  x860 &  x863 &  x866 &  x875 &  x878 &  x881 &  x884 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x935 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x962 &  x965 &  x968 &  x971 &  x974 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x714 & ~x753 & ~x792 & ~x831 & ~x888;
assign c656 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x56 &  x59 &  x65 &  x70 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x95 &  x101 &  x104 &  x107 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x188 &  x194 &  x200 &  x203 &  x206 &  x212 &  x215 &  x218 &  x224 &  x227 &  x230 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x263 &  x266 &  x281 &  x284 &  x290 &  x296 &  x298 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x329 &  x338 &  x341 &  x347 &  x353 &  x365 &  x368 &  x371 &  x374 &  x376 &  x377 &  x380 &  x386 &  x389 &  x392 &  x401 &  x407 &  x410 &  x413 &  x416 &  x425 &  x433 &  x434 &  x440 &  x443 &  x446 &  x452 &  x461 &  x467 &  x470 &  x473 &  x482 &  x485 &  x488 &  x494 &  x497 &  x503 &  x509 &  x515 &  x521 &  x524 &  x527 &  x533 &  x536 &  x542 &  x545 &  x548 &  x551 &  x554 &  x560 &  x563 &  x569 &  x572 &  x575 &  x581 &  x584 &  x590 &  x593 &  x599 &  x602 &  x608 &  x614 &  x617 &  x623 &  x632 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x665 &  x668 &  x671 &  x674 &  x686 &  x689 &  x692 &  x698 &  x701 &  x704 &  x710 &  x713 &  x716 &  x719 &  x728 &  x740 &  x749 &  x755 &  x764 &  x767 &  x770 &  x776 &  x779 &  x782 &  x791 &  x794 &  x809 &  x815 &  x824 &  x827 &  x836 &  x839 &  x851 &  x857 &  x860 &  x869 &  x878 &  x881 &  x887 &  x890 &  x899 &  x902 &  x908 &  x911 &  x914 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x965 &  x967 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x998 &  x1004 &  x1006 &  x1007 &  x1010 &  x1016 &  x1019 &  x1025 &  x1028 &  x1037 &  x1040 &  x1043 &  x1045 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1100 &  x1109 &  x1112 &  x1118 &  x1124 &  x1127 &  x1130 & ~x405 & ~x480 & ~x702 & ~x780 & ~x819 & ~x897;
assign c658 =  x5 &  x8 &  x11 &  x14 &  x17 &  x26 &  x29 &  x32 &  x35 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x65 &  x68 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x128 &  x131 &  x134 &  x137 &  x146 &  x149 &  x152 &  x155 &  x158 &  x164 &  x167 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x206 &  x212 &  x215 &  x218 &  x221 &  x227 &  x230 &  x233 &  x236 &  x239 &  x251 &  x254 &  x257 &  x260 &  x263 &  x272 &  x275 &  x278 &  x281 &  x287 &  x290 &  x296 &  x305 &  x308 &  x311 &  x314 &  x320 &  x323 &  x326 &  x329 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x356 &  x362 &  x365 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x416 &  x422 &  x428 &  x431 &  x434 &  x443 &  x446 &  x457 &  x458 &  x461 &  x464 &  x466 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x506 &  x509 &  x521 &  x524 &  x530 &  x536 &  x539 &  x542 &  x545 &  x551 &  x554 &  x566 &  x569 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x602 &  x608 &  x611 &  x614 &  x617 &  x623 &  x626 &  x632 &  x635 &  x641 &  x644 &  x650 &  x656 &  x659 &  x662 &  x665 &  x671 &  x674 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x701 &  x704 &  x707 &  x713 &  x716 &  x719 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x749 &  x752 &  x755 &  x758 &  x761 &  x767 &  x773 &  x776 &  x779 &  x782 &  x784 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x824 &  x827 &  x830 &  x845 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x911 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x940 &  x941 &  x944 &  x947 &  x956 &  x959 &  x962 &  x977 &  x979 &  x983 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1018 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1058 &  x1061 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1096 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 & ~x306 & ~x354 & ~x390 & ~x429 & ~x468 & ~x756 & ~x757 & ~x796 & ~x870;
assign c660 =  x5 &  x8 &  x11 &  x17 &  x20 &  x23 &  x26 &  x29 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x107 &  x116 &  x119 &  x122 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x155 &  x158 &  x161 &  x163 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x188 &  x194 &  x197 &  x200 &  x202 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x241 &  x242 &  x245 &  x248 &  x254 &  x257 &  x260 &  x263 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x353 &  x356 &  x358 &  x359 &  x362 &  x368 &  x371 &  x376 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x415 &  x416 &  x422 &  x425 &  x427 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x449 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x488 &  x491 &  x493 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x532 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x590 &  x593 &  x596 &  x602 &  x605 &  x608 &  x614 &  x617 &  x620 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x653 &  x656 &  x659 &  x665 &  x668 &  x671 &  x674 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x782 &  x785 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x890 &  x893 &  x899 &  x902 &  x905 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x931 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x959 &  x965 &  x968 &  x971 &  x977 &  x980 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x675 & ~x714 & ~x831 & ~x870;
assign c662 =  x5 &  x8 &  x14 &  x20 &  x26 &  x29 &  x38 &  x41 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x107 &  x110 &  x113 &  x115 &  x116 &  x119 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x149 &  x152 &  x155 &  x161 &  x170 &  x173 &  x179 &  x182 &  x185 &  x191 &  x203 &  x209 &  x218 &  x221 &  x224 &  x233 &  x239 &  x248 &  x251 &  x254 &  x263 &  x266 &  x272 &  x275 &  x278 &  x281 &  x287 &  x293 &  x296 &  x302 &  x308 &  x311 &  x314 &  x320 &  x326 &  x329 &  x335 &  x338 &  x344 &  x350 &  x353 &  x355 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x395 &  x401 &  x404 &  x410 &  x416 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x449 &  x452 &  x458 &  x461 &  x464 &  x467 &  x470 &  x472 &  x476 &  x479 &  x482 &  x485 &  x494 &  x497 &  x500 &  x506 &  x509 &  x512 &  x518 &  x521 &  x524 &  x530 &  x533 &  x542 &  x548 &  x557 &  x563 &  x572 &  x575 &  x578 &  x581 &  x584 &  x596 &  x602 &  x605 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x680 &  x683 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x716 &  x727 &  x734 &  x743 &  x746 &  x752 &  x760 &  x761 &  x764 &  x779 &  x791 &  x793 &  x799 &  x800 &  x806 &  x815 &  x818 &  x821 &  x824 &  x830 &  x836 &  x839 &  x845 &  x848 &  x851 &  x857 &  x860 &  x866 &  x869 &  x875 &  x878 &  x881 &  x884 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x950 &  x961 &  x962 &  x965 &  x967 &  x971 &  x974 &  x977 &  x980 &  x989 &  x992 &  x998 &  x1000 &  x1001 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1028 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1106 &  x1112 &  x1118 &  x1124 &  x1130 & ~x366 & ~x402 & ~x405 & ~x441 & ~x480 & ~x663 & ~x741 & ~x780 & ~x819 & ~x858 & ~x897;
assign c664 =  x5 &  x8 &  x20 &  x29 &  x35 &  x38 &  x50 &  x56 &  x59 &  x62 &  x68 &  x74 &  x77 &  x86 &  x89 &  x95 &  x98 &  x119 &  x128 &  x131 &  x140 &  x149 &  x161 &  x164 &  x167 &  x182 &  x188 &  x200 &  x209 &  x215 &  x218 &  x224 &  x230 &  x239 &  x242 &  x251 &  x260 &  x281 &  x308 &  x311 &  x314 &  x320 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x359 &  x383 &  x389 &  x392 &  x395 &  x401 &  x407 &  x410 &  x416 &  x422 &  x428 &  x434 &  x443 &  x446 &  x449 &  x452 &  x458 &  x461 &  x464 &  x470 &  x473 &  x488 &  x491 &  x493 &  x494 &  x497 &  x500 &  x503 &  x506 &  x524 &  x533 &  x536 &  x539 &  x542 &  x551 &  x557 &  x566 &  x571 &  x584 &  x596 &  x608 &  x611 &  x614 &  x623 &  x638 &  x649 &  x662 &  x665 &  x674 &  x695 &  x710 &  x713 &  x716 &  x728 &  x740 &  x746 &  x749 &  x752 &  x755 &  x773 &  x782 &  x785 &  x800 &  x803 &  x812 &  x818 &  x821 &  x833 &  x836 &  x839 &  x848 &  x851 &  x863 &  x866 &  x869 &  x872 &  x878 &  x890 &  x893 &  x899 &  x920 &  x923 &  x926 &  x929 &  x935 &  x944 &  x947 &  x956 &  x971 &  x974 &  x986 &  x992 &  x1001 &  x1004 &  x1010 &  x1016 &  x1025 &  x1028 &  x1031 &  x1034 &  x1043 &  x1058 &  x1061 &  x1064 &  x1067 &  x1091 &  x1094 &  x1103 &  x1112 &  x1121 &  x1127 & ~x210 & ~x225 & ~x477 & ~x633 & ~x672 & ~x711 & ~x789 & ~x828 & ~x906 & ~x945 & ~x946 & ~x984;
assign c666 =  x2 &  x5 &  x8 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x47 &  x50 &  x53 &  x62 &  x71 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x140 &  x149 &  x152 &  x158 &  x164 &  x167 &  x170 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x206 &  x209 &  x212 &  x218 &  x221 &  x224 &  x230 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x263 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x293 &  x296 &  x299 &  x308 &  x311 &  x317 &  x320 &  x323 &  x326 &  x329 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x374 &  x380 &  x386 &  x392 &  x395 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x437 &  x440 &  x443 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x518 &  x521 &  x524 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x554 &  x557 &  x560 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x587 &  x590 &  x593 &  x599 &  x602 &  x614 &  x617 &  x623 &  x626 &  x629 &  x632 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x794 &  x797 &  x803 &  x806 &  x809 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x845 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x934 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x156 & ~x195 & ~x196 & ~x288 & ~x561 & ~x741 & ~x780 & ~x783;
assign c668 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x38 &  x41 &  x44 &  x53 &  x56 &  x59 &  x62 &  x65 &  x74 &  x80 &  x83 &  x86 &  x95 &  x98 &  x101 &  x104 &  x107 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x155 &  x158 &  x161 &  x170 &  x176 &  x179 &  x185 &  x188 &  x194 &  x197 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x230 &  x236 &  x239 &  x242 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x314 &  x320 &  x323 &  x326 &  x329 &  x335 &  x338 &  x344 &  x347 &  x350 &  x353 &  x359 &  x362 &  x365 &  x368 &  x371 &  x377 &  x379 &  x380 &  x386 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x417 &  x418 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x446 &  x452 &  x455 &  x457 &  x458 &  x461 &  x464 &  x470 &  x473 &  x476 &  x482 &  x485 &  x488 &  x491 &  x494 &  x496 &  x497 &  x503 &  x506 &  x509 &  x512 &  x515 &  x521 &  x524 &  x527 &  x533 &  x535 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x590 &  x596 &  x599 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x665 &  x668 &  x671 &  x674 &  x677 &  x689 &  x698 &  x701 &  x710 &  x716 &  x722 &  x725 &  x728 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x961 &  x962 &  x968 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1000 &  x1004 &  x1007 &  x1010 &  x1013 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 & ~x480 & ~x513 & ~x519 & ~x558 & ~x597;
assign c670 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x35 &  x38 &  x44 &  x53 &  x56 &  x59 &  x62 &  x65 &  x71 &  x77 &  x80 &  x83 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x125 &  x127 &  x128 &  x131 &  x137 &  x140 &  x143 &  x152 &  x155 &  x161 &  x164 &  x166 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x194 &  x197 &  x200 &  x206 &  x209 &  x215 &  x218 &  x221 &  x224 &  x230 &  x233 &  x236 &  x242 &  x245 &  x247 &  x248 &  x254 &  x263 &  x266 &  x269 &  x272 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x323 &  x326 &  x329 &  x332 &  x335 &  x341 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x383 &  x386 &  x388 &  x389 &  x392 &  x395 &  x398 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x427 &  x428 &  x434 &  x437 &  x443 &  x446 &  x449 &  x455 &  x458 &  x461 &  x466 &  x467 &  x470 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x505 &  x506 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x572 &  x578 &  x581 &  x587 &  x590 &  x593 &  x605 &  x608 &  x611 &  x614 &  x617 &  x623 &  x629 &  x644 &  x647 &  x650 &  x656 &  x659 &  x665 &  x668 &  x674 &  x677 &  x680 &  x683 &  x689 &  x695 &  x698 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x746 &  x749 &  x752 &  x755 &  x758 &  x764 &  x767 &  x770 &  x773 &  x776 &  x782 &  x788 &  x791 &  x794 &  x797 &  x803 &  x806 &  x809 &  x812 &  x818 &  x821 &  x824 &  x830 &  x833 &  x836 &  x839 &  x842 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x908 &  x911 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x156 & ~x195 & ~x234 & ~x273 & ~x312 & ~x600 & ~x639 & ~x678 & ~x1068;
assign c672 =  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x44 &  x50 &  x53 &  x56 &  x65 &  x68 &  x74 &  x77 &  x83 &  x89 &  x92 &  x95 &  x98 &  x101 &  x107 &  x110 &  x113 &  x122 &  x128 &  x134 &  x137 &  x146 &  x152 &  x155 &  x158 &  x161 &  x167 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x200 &  x203 &  x209 &  x212 &  x218 &  x221 &  x224 &  x227 &  x236 &  x239 &  x245 &  x248 &  x251 &  x254 &  x260 &  x263 &  x269 &  x284 &  x287 &  x293 &  x296 &  x305 &  x311 &  x314 &  x317 &  x320 &  x326 &  x329 &  x332 &  x338 &  x341 &  x362 &  x365 &  x368 &  x371 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x404 &  x407 &  x410 &  x413 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x443 &  x446 &  x449 &  x455 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x494 &  x497 &  x506 &  x509 &  x512 &  x521 &  x529 &  x530 &  x533 &  x536 &  x538 &  x542 &  x554 &  x557 &  x560 &  x563 &  x566 &  x568 &  x569 &  x575 &  x578 &  x584 &  x587 &  x590 &  x593 &  x596 &  x605 &  x611 &  x614 &  x617 &  x623 &  x629 &  x632 &  x638 &  x644 &  x647 &  x650 &  x659 &  x662 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x737 &  x740 &  x743 &  x752 &  x755 &  x761 &  x764 &  x767 &  x770 &  x773 &  x784 &  x785 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x821 &  x823 &  x827 &  x836 &  x839 &  x845 &  x848 &  x851 &  x866 &  x875 &  x878 &  x881 &  x899 &  x902 &  x905 &  x908 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x938 &  x941 &  x944 &  x947 &  x950 &  x956 &  x959 &  x962 &  x965 &  x968 &  x977 &  x979 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1013 &  x1016 &  x1018 &  x1019 &  x1025 &  x1028 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1057 &  x1058 &  x1061 &  x1067 &  x1070 &  x1076 &  x1082 &  x1091 &  x1094 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1130 & ~x351 & ~x390 & ~x391 & ~x714 & ~x756 & ~x792 & ~x873;
assign c674 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x661 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x700 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x93 & ~x132 & ~x171 & ~x210 & ~x249 & ~x288 & ~x327 & ~x366 & ~x402 & ~x441 & ~x480 & ~x624 & ~x663 & ~x702 & ~x741 & ~x780 & ~x783 & ~x819 & ~x858 & ~x897 & ~x936 & ~x939 & ~x975 & ~x978 & ~x1014 & ~x1053 & ~x1092;
assign c676 =  x2 &  x8 &  x11 &  x14 &  x17 &  x23 &  x26 &  x35 &  x38 &  x41 &  x44 &  x50 &  x53 &  x56 &  x59 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x106 &  x107 &  x110 &  x113 &  x116 &  x119 &  x125 &  x131 &  x134 &  x137 &  x139 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x167 &  x170 &  x173 &  x176 &  x178 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x217 &  x218 &  x221 &  x223 &  x227 &  x230 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x256 &  x260 &  x263 &  x266 &  x272 &  x275 &  x281 &  x284 &  x290 &  x293 &  x295 &  x296 &  x299 &  x302 &  x305 &  x308 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x340 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x361 &  x362 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x416 &  x419 &  x421 &  x425 &  x428 &  x431 &  x434 &  x437 &  x443 &  x446 &  x451 &  x452 &  x455 &  x457 &  x458 &  x461 &  x464 &  x476 &  x479 &  x482 &  x485 &  x488 &  x493 &  x494 &  x496 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x524 &  x527 &  x529 &  x530 &  x532 &  x533 &  x535 &  x539 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x568 &  x569 &  x575 &  x578 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x607 &  x608 &  x611 &  x613 &  x614 &  x620 &  x623 &  x626 &  x629 &  x635 &  x638 &  x641 &  x644 &  x646 &  x647 &  x653 &  x656 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x691 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x730 &  x734 &  x737 &  x740 &  x746 &  x749 &  x752 &  x758 &  x761 &  x763 &  x764 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x802 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x827 &  x830 &  x833 &  x836 &  x839 &  x845 &  x848 &  x851 &  x854 &  x857 &  x863 &  x866 &  x872 &  x875 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x958 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x980 &  x983 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1025 &  x1028 &  x1034 &  x1036 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1061 &  x1064 &  x1073 &  x1075 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1114 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130;
assign c678 =  x2 &  x5 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x74 &  x77 &  x79 &  x80 &  x83 &  x86 &  x89 &  x95 &  x101 &  x107 &  x110 &  x113 &  x119 &  x122 &  x125 &  x134 &  x143 &  x146 &  x152 &  x155 &  x158 &  x161 &  x163 &  x167 &  x170 &  x173 &  x179 &  x182 &  x191 &  x200 &  x203 &  x206 &  x209 &  x212 &  x218 &  x221 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x257 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x293 &  x296 &  x299 &  x302 &  x307 &  x311 &  x317 &  x323 &  x329 &  x341 &  x344 &  x347 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x389 &  x392 &  x395 &  x397 &  x398 &  x401 &  x404 &  x410 &  x413 &  x415 &  x416 &  x422 &  x425 &  x428 &  x436 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x464 &  x467 &  x470 &  x476 &  x479 &  x491 &  x493 &  x497 &  x505 &  x509 &  x512 &  x515 &  x521 &  x524 &  x527 &  x530 &  x532 &  x533 &  x536 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x584 &  x587 &  x590 &  x602 &  x605 &  x608 &  x610 &  x611 &  x614 &  x617 &  x620 &  x623 &  x629 &  x632 &  x635 &  x641 &  x644 &  x649 &  x650 &  x653 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x680 &  x686 &  x688 &  x689 &  x695 &  x698 &  x704 &  x707 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x734 &  x737 &  x740 &  x746 &  x752 &  x755 &  x758 &  x773 &  x775 &  x776 &  x782 &  x788 &  x791 &  x794 &  x800 &  x802 &  x803 &  x806 &  x809 &  x812 &  x815 &  x821 &  x824 &  x827 &  x833 &  x836 &  x841 &  x842 &  x845 &  x848 &  x851 &  x857 &  x860 &  x863 &  x866 &  x869 &  x880 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x935 &  x944 &  x947 &  x953 &  x962 &  x965 &  x968 &  x971 &  x974 &  x976 &  x983 &  x989 &  x995 &  x997 &  x1001 &  x1007 &  x1010 &  x1015 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1043 &  x1049 &  x1052 &  x1054 &  x1058 &  x1061 &  x1064 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1103 &  x1106 &  x1109 &  x1112 &  x1114 &  x1115 &  x1118 &  x1124 &  x1127;
assign c680 =  x5 &  x8 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x59 &  x62 &  x68 &  x71 &  x74 &  x77 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x107 &  x110 &  x113 &  x116 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x218 &  x224 &  x227 &  x233 &  x236 &  x239 &  x248 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x317 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x353 &  x356 &  x362 &  x365 &  x368 &  x374 &  x377 &  x380 &  x383 &  x386 &  x392 &  x395 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x458 &  x467 &  x470 &  x473 &  x476 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x656 &  x659 &  x661 &  x662 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x707 &  x710 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x761 &  x770 &  x773 &  x778 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x815 &  x817 &  x818 &  x821 &  x824 &  x827 &  x833 &  x836 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x866 &  x869 &  x875 &  x878 &  x884 &  x887 &  x893 &  x896 &  x899 &  x905 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x935 &  x938 &  x941 &  x944 &  x947 &  x953 &  x956 &  x959 &  x962 &  x965 &  x971 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 &  x1130 & ~x78 & ~x171 & ~x288 & ~x327 & ~x366 & ~x405 & ~x468 & ~x549 & ~x1101;
assign c682 =  x1 &  x5 &  x11 &  x16 &  x17 &  x20 &  x29 &  x35 &  x44 &  x47 &  x67 &  x71 &  x74 &  x92 &  x95 &  x104 &  x110 &  x113 &  x119 &  x122 &  x131 &  x137 &  x140 &  x143 &  x152 &  x158 &  x161 &  x179 &  x185 &  x191 &  x197 &  x206 &  x209 &  x217 &  x223 &  x224 &  x236 &  x251 &  x256 &  x262 &  x275 &  x287 &  x301 &  x302 &  x314 &  x317 &  x326 &  x339 &  x340 &  x344 &  x347 &  x350 &  x356 &  x362 &  x365 &  x378 &  x392 &  x401 &  x412 &  x431 &  x443 &  x451 &  x461 &  x464 &  x470 &  x473 &  x476 &  x485 &  x490 &  x494 &  x512 &  x518 &  x528 &  x536 &  x545 &  x548 &  x566 &  x568 &  x575 &  x578 &  x593 &  x617 &  x638 &  x656 &  x659 &  x665 &  x674 &  x695 &  x698 &  x719 &  x734 &  x737 &  x755 &  x764 &  x779 &  x791 &  x797 &  x800 &  x802 &  x814 &  x821 &  x836 &  x841 &  x860 &  x866 &  x869 &  x878 &  x880 &  x881 &  x893 &  x899 &  x902 &  x932 &  x947 &  x958 &  x959 &  x992 &  x997 &  x1013 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1049 &  x1055 &  x1058 &  x1061 &  x1076 &  x1079 &  x1082 &  x1088 &  x1112 &  x1115 &  x1118;
assign c684 =  x8 &  x17 &  x23 &  x29 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x71 &  x77 &  x82 &  x83 &  x92 &  x101 &  x107 &  x110 &  x113 &  x116 &  x121 &  x125 &  x128 &  x131 &  x137 &  x140 &  x146 &  x155 &  x158 &  x160 &  x161 &  x164 &  x167 &  x179 &  x182 &  x197 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x236 &  x239 &  x245 &  x248 &  x254 &  x257 &  x260 &  x266 &  x277 &  x281 &  x284 &  x293 &  x299 &  x305 &  x314 &  x320 &  x323 &  x335 &  x338 &  x341 &  x344 &  x356 &  x362 &  x365 &  x368 &  x371 &  x374 &  x380 &  x383 &  x392 &  x395 &  x398 &  x401 &  x416 &  x419 &  x422 &  x425 &  x437 &  x440 &  x446 &  x455 &  x463 &  x464 &  x473 &  x479 &  x488 &  x491 &  x509 &  x512 &  x515 &  x518 &  x524 &  x527 &  x536 &  x551 &  x557 &  x560 &  x563 &  x569 &  x575 &  x581 &  x584 &  x587 &  x593 &  x602 &  x605 &  x614 &  x620 &  x622 &  x632 &  x635 &  x641 &  x644 &  x650 &  x653 &  x656 &  x659 &  x661 &  x665 &  x674 &  x677 &  x704 &  x707 &  x710 &  x716 &  x719 &  x728 &  x731 &  x740 &  x749 &  x752 &  x764 &  x767 &  x773 &  x785 &  x788 &  x791 &  x800 &  x806 &  x809 &  x817 &  x821 &  x824 &  x833 &  x842 &  x851 &  x856 &  x857 &  x866 &  x875 &  x877 &  x878 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x911 &  x914 &  x929 &  x935 &  x938 &  x947 &  x956 &  x965 &  x968 &  x974 &  x980 &  x986 &  x1001 &  x1013 &  x1016 &  x1025 &  x1028 &  x1034 &  x1037 &  x1052 &  x1058 &  x1064 &  x1079 &  x1088 &  x1094 &  x1097 &  x1100 &  x1106 &  x1121 & ~x54 & ~x93 & ~x249 & ~x393;
assign c686 =  x5 &  x17 &  x23 &  x62 &  x68 &  x74 &  x77 &  x92 &  x95 &  x101 &  x122 &  x125 &  x134 &  x140 &  x149 &  x161 &  x164 &  x170 &  x179 &  x194 &  x218 &  x221 &  x236 &  x242 &  x245 &  x254 &  x260 &  x263 &  x269 &  x271 &  x272 &  x275 &  x287 &  x299 &  x329 &  x335 &  x338 &  x341 &  x350 &  x355 &  x356 &  x362 &  x368 &  x377 &  x383 &  x389 &  x392 &  x394 &  x401 &  x404 &  x407 &  x422 &  x428 &  x437 &  x440 &  x443 &  x452 &  x464 &  x467 &  x482 &  x509 &  x533 &  x536 &  x539 &  x545 &  x548 &  x569 &  x572 &  x578 &  x584 &  x596 &  x602 &  x611 &  x617 &  x620 &  x623 &  x635 &  x641 &  x650 &  x653 &  x665 &  x701 &  x704 &  x716 &  x719 &  x725 &  x728 &  x731 &  x734 &  x737 &  x752 &  x770 &  x782 &  x794 &  x797 &  x800 &  x803 &  x806 &  x818 &  x836 &  x854 &  x860 &  x866 &  x869 &  x872 &  x905 &  x908 &  x928 &  x938 &  x941 &  x944 &  x947 &  x950 &  x955 &  x956 &  x959 &  x961 &  x965 &  x973 &  x974 &  x995 &  x1000 &  x1013 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1052 &  x1055 &  x1067 &  x1070 &  x1072 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1097 &  x1100 &  x1103 &  x1115 &  x1127 &  x1130 & ~x54 & ~x444 & ~x741 & ~x744 & ~x780 & ~x822 & ~x897 & ~x936 & ~x975;
assign c688 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x38 &  x41 &  x44 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x74 &  x77 &  x80 &  x89 &  x92 &  x95 &  x104 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x191 &  x194 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x242 &  x245 &  x251 &  x254 &  x260 &  x263 &  x266 &  x272 &  x275 &  x278 &  x284 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x338 &  x341 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x377 &  x380 &  x383 &  x389 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x446 &  x455 &  x458 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x485 &  x488 &  x491 &  x494 &  x497 &  x512 &  x515 &  x527 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x599 &  x602 &  x605 &  x608 &  x614 &  x620 &  x623 &  x629 &  x641 &  x650 &  x653 &  x659 &  x662 &  x665 &  x674 &  x680 &  x683 &  x686 &  x689 &  x695 &  x698 &  x704 &  x710 &  x713 &  x719 &  x722 &  x731 &  x740 &  x743 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x821 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x896 &  x899 &  x902 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1013 &  x1016 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1085 &  x1088 &  x1091 &  x1094 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1130 & ~x195 & ~x198 & ~x234 & ~x237 & ~x273 & ~x312 & ~x444 & ~x483 & ~x522 & ~x561 & ~x897 & ~x948 & ~x981 & ~x987 & ~x1020 & ~x1059;
assign c690 =  x5 &  x8 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x59 &  x62 &  x65 &  x71 &  x77 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x104 &  x110 &  x113 &  x119 &  x122 &  x125 &  x128 &  x131 &  x137 &  x140 &  x146 &  x152 &  x155 &  x158 &  x170 &  x173 &  x176 &  x179 &  x188 &  x191 &  x194 &  x200 &  x206 &  x212 &  x224 &  x227 &  x230 &  x233 &  x242 &  x248 &  x251 &  x254 &  x260 &  x263 &  x266 &  x269 &  x271 &  x272 &  x275 &  x278 &  x281 &  x284 &  x290 &  x293 &  x299 &  x302 &  x305 &  x308 &  x314 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x347 &  x350 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x380 &  x398 &  x401 &  x404 &  x407 &  x413 &  x416 &  x419 &  x422 &  x425 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x467 &  x470 &  x476 &  x482 &  x488 &  x494 &  x497 &  x503 &  x506 &  x509 &  x512 &  x518 &  x521 &  x524 &  x530 &  x533 &  x536 &  x539 &  x544 &  x545 &  x548 &  x551 &  x554 &  x557 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x583 &  x584 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x614 &  x620 &  x622 &  x623 &  x626 &  x629 &  x638 &  x641 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x671 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x728 &  x731 &  x734 &  x740 &  x743 &  x746 &  x749 &  x752 &  x761 &  x773 &  x776 &  x779 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x809 &  x812 &  x815 &  x818 &  x827 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x854 &  x856 &  x857 &  x860 &  x863 &  x866 &  x872 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x947 &  x950 &  x953 &  x962 &  x965 &  x968 &  x974 &  x980 &  x989 &  x992 &  x995 &  x1001 &  x1007 &  x1013 &  x1016 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1112 &  x1118 &  x1124 &  x1130 & ~x210 & ~x234 & ~x1017;
assign c692 =  x2 &  x5 &  x8 &  x14 &  x17 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x53 &  x56 &  x62 &  x65 &  x71 &  x74 &  x80 &  x83 &  x92 &  x98 &  x104 &  x107 &  x113 &  x122 &  x125 &  x128 &  x134 &  x137 &  x143 &  x149 &  x155 &  x158 &  x161 &  x173 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x239 &  x242 &  x245 &  x251 &  x257 &  x260 &  x266 &  x277 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x302 &  x305 &  x308 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x341 &  x344 &  x347 &  x350 &  x353 &  x365 &  x368 &  x377 &  x383 &  x386 &  x389 &  x392 &  x401 &  x404 &  x410 &  x413 &  x422 &  x434 &  x437 &  x440 &  x449 &  x452 &  x455 &  x458 &  x461 &  x467 &  x470 &  x473 &  x482 &  x488 &  x494 &  x497 &  x500 &  x503 &  x506 &  x512 &  x515 &  x518 &  x521 &  x524 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x575 &  x578 &  x581 &  x584 &  x590 &  x593 &  x596 &  x602 &  x605 &  x611 &  x614 &  x617 &  x620 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x653 &  x656 &  x665 &  x671 &  x677 &  x683 &  x686 &  x695 &  x701 &  x710 &  x719 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x767 &  x770 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x812 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x869 &  x872 &  x875 &  x877 &  x896 &  x916 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x944 &  x950 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x983 &  x986 &  x992 &  x1001 &  x1004 &  x1010 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1040 &  x1046 &  x1049 &  x1052 &  x1058 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1123 & ~x93 & ~x132 & ~x171 & ~x210 & ~x249 & ~x288 & ~x468 & ~x507 & ~x546 & ~x549 & ~x588 & ~x834 & ~x873;
assign c694 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x86 &  x89 &  x92 &  x98 &  x101 &  x104 &  x107 &  x113 &  x116 &  x119 &  x125 &  x128 &  x131 &  x134 &  x137 &  x143 &  x146 &  x149 &  x152 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x368 &  x374 &  x377 &  x380 &  x383 &  x389 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x491 &  x494 &  x497 &  x500 &  x509 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x671 &  x674 &  x680 &  x686 &  x689 &  x692 &  x698 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x761 &  x764 &  x767 &  x770 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x833 &  x836 &  x839 &  x842 &  x845 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x875 &  x878 &  x881 &  x890 &  x893 &  x896 &  x899 &  x908 &  x911 &  x913 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x940 &  x941 &  x944 &  x947 &  x950 &  x953 &  x959 &  x962 &  x965 &  x968 &  x974 &  x977 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1010 &  x1013 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x48 & ~x282 & ~x402 & ~x441 & ~x474 & ~x480 & ~x513 & ~x519;
assign c696 =  x1 &  x11 &  x20 &  x23 &  x35 &  x40 &  x47 &  x50 &  x53 &  x59 &  x62 &  x65 &  x68 &  x80 &  x86 &  x92 &  x95 &  x98 &  x100 &  x104 &  x110 &  x112 &  x113 &  x116 &  x119 &  x131 &  x139 &  x140 &  x143 &  x149 &  x152 &  x161 &  x164 &  x167 &  x170 &  x176 &  x178 &  x179 &  x190 &  x197 &  x203 &  x218 &  x236 &  x245 &  x251 &  x254 &  x260 &  x266 &  x269 &  x272 &  x278 &  x281 &  x284 &  x287 &  x290 &  x295 &  x296 &  x299 &  x305 &  x308 &  x320 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x365 &  x374 &  x392 &  x395 &  x401 &  x410 &  x413 &  x425 &  x428 &  x434 &  x440 &  x443 &  x446 &  x455 &  x458 &  x467 &  x473 &  x476 &  x479 &  x482 &  x491 &  x494 &  x500 &  x503 &  x506 &  x512 &  x539 &  x542 &  x545 &  x548 &  x551 &  x560 &  x566 &  x572 &  x578 &  x587 &  x590 &  x605 &  x608 &  x611 &  x623 &  x626 &  x647 &  x650 &  x653 &  x658 &  x662 &  x665 &  x668 &  x671 &  x683 &  x689 &  x710 &  x713 &  x719 &  x722 &  x731 &  x737 &  x743 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x782 &  x785 &  x791 &  x800 &  x803 &  x806 &  x818 &  x821 &  x824 &  x830 &  x833 &  x836 &  x839 &  x841 &  x860 &  x863 &  x866 &  x869 &  x878 &  x880 &  x890 &  x893 &  x899 &  x908 &  x911 &  x920 &  x926 &  x932 &  x938 &  x950 &  x956 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1010 &  x1025 &  x1028 &  x1034 &  x1037 &  x1040 &  x1049 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1130 & ~x321 & ~x441 & ~x519 & ~x597 & ~x642;
assign c698 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x29 &  x32 &  x38 &  x44 &  x47 &  x50 &  x53 &  x56 &  x62 &  x68 &  x71 &  x74 &  x77 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x110 &  x113 &  x116 &  x119 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x158 &  x161 &  x167 &  x170 &  x173 &  x176 &  x179 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x233 &  x245 &  x248 &  x251 &  x257 &  x260 &  x266 &  x269 &  x272 &  x278 &  x281 &  x284 &  x290 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x323 &  x329 &  x332 &  x338 &  x341 &  x343 &  x344 &  x350 &  x353 &  x359 &  x362 &  x365 &  x368 &  x371 &  x380 &  x386 &  x389 &  x392 &  x395 &  x398 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x428 &  x431 &  x437 &  x440 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x476 &  x479 &  x482 &  x488 &  x491 &  x494 &  x497 &  x499 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x527 &  x530 &  x533 &  x537 &  x538 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x560 &  x563 &  x566 &  x569 &  x581 &  x583 &  x584 &  x587 &  x596 &  x599 &  x602 &  x608 &  x611 &  x617 &  x622 &  x623 &  x629 &  x635 &  x638 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x661 &  x662 &  x665 &  x668 &  x671 &  x680 &  x683 &  x686 &  x692 &  x695 &  x707 &  x716 &  x719 &  x722 &  x725 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x761 &  x764 &  x767 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x803 &  x806 &  x812 &  x821 &  x823 &  x824 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x953 &  x956 &  x959 &  x962 &  x968 &  x971 &  x974 &  x977 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1018 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1055 &  x1057 &  x1058 &  x1061 &  x1067 &  x1069 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1096 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x471;
assign c6100 =  x2 &  x5 &  x8 &  x14 &  x17 &  x23 &  x29 &  x32 &  x35 &  x38 &  x41 &  x47 &  x50 &  x53 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x92 &  x110 &  x113 &  x116 &  x131 &  x143 &  x152 &  x155 &  x158 &  x167 &  x170 &  x173 &  x179 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x212 &  x230 &  x236 &  x239 &  x245 &  x248 &  x254 &  x263 &  x266 &  x269 &  x275 &  x278 &  x281 &  x290 &  x293 &  x296 &  x302 &  x305 &  x308 &  x311 &  x317 &  x323 &  x326 &  x329 &  x332 &  x335 &  x341 &  x344 &  x347 &  x353 &  x365 &  x368 &  x371 &  x374 &  x377 &  x383 &  x388 &  x389 &  x395 &  x398 &  x401 &  x404 &  x416 &  x421 &  x422 &  x425 &  x427 &  x431 &  x434 &  x440 &  x443 &  x455 &  x460 &  x461 &  x464 &  x466 &  x470 &  x473 &  x476 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x509 &  x512 &  x515 &  x530 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x557 &  x560 &  x563 &  x571 &  x572 &  x578 &  x584 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x623 &  x626 &  x635 &  x641 &  x647 &  x650 &  x653 &  x656 &  x659 &  x665 &  x671 &  x677 &  x680 &  x683 &  x689 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x722 &  x725 &  x731 &  x740 &  x743 &  x749 &  x764 &  x767 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x800 &  x806 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x845 &  x848 &  x851 &  x854 &  x860 &  x866 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x908 &  x914 &  x920 &  x926 &  x932 &  x938 &  x944 &  x953 &  x956 &  x965 &  x968 &  x971 &  x979 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1019 &  x1022 &  x1025 &  x1028 &  x1043 &  x1049 &  x1055 &  x1058 &  x1061 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 & ~x273 & ~x312 & ~x351 & ~x390 & ~x391 & ~x430 & ~x438 & ~x507 & ~x717 & ~x753 & ~x756 & ~x795 & ~x834 & ~x873;
assign c6102 =  x2 &  x5 &  x8 &  x11 &  x20 &  x23 &  x29 &  x32 &  x35 &  x38 &  x44 &  x47 &  x50 &  x53 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x317 &  x320 &  x326 &  x329 &  x332 &  x335 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x386 &  x389 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x566 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x614 &  x617 &  x620 &  x623 &  x626 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x728 &  x731 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x989 &  x992 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x9 & ~x48 & ~x171 & ~x210 & ~x249 & ~x288 & ~x438 & ~x444 & ~x483 & ~x516 & ~x756 & ~x858 & ~x897 & ~x906 & ~x945 & ~x951 & ~x984 & ~x990 & ~x1023 & ~x1068 & ~x1107;
assign c6104 =  x2 &  x8 &  x11 &  x20 &  x29 &  x32 &  x38 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x77 &  x86 &  x92 &  x98 &  x101 &  x104 &  x107 &  x113 &  x116 &  x122 &  x131 &  x134 &  x143 &  x164 &  x170 &  x173 &  x182 &  x185 &  x188 &  x194 &  x215 &  x224 &  x233 &  x236 &  x239 &  x248 &  x251 &  x254 &  x260 &  x263 &  x272 &  x275 &  x284 &  x290 &  x296 &  x299 &  x308 &  x320 &  x323 &  x329 &  x347 &  x353 &  x359 &  x371 &  x377 &  x380 &  x386 &  x392 &  x398 &  x401 &  x404 &  x407 &  x418 &  x422 &  x428 &  x431 &  x443 &  x446 &  x455 &  x458 &  x476 &  x482 &  x485 &  x491 &  x494 &  x503 &  x506 &  x509 &  x521 &  x524 &  x527 &  x542 &  x545 &  x550 &  x557 &  x560 &  x563 &  x566 &  x575 &  x581 &  x587 &  x602 &  x605 &  x611 &  x626 &  x632 &  x641 &  x647 &  x653 &  x659 &  x665 &  x677 &  x680 &  x686 &  x692 &  x698 &  x704 &  x710 &  x716 &  x725 &  x728 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x764 &  x767 &  x779 &  x788 &  x797 &  x809 &  x815 &  x824 &  x827 &  x833 &  x839 &  x845 &  x875 &  x878 &  x887 &  x914 &  x917 &  x920 &  x926 &  x935 &  x938 &  x944 &  x956 &  x968 &  x977 &  x989 &  x998 &  x1001 &  x1007 &  x1010 &  x1019 &  x1028 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1064 &  x1073 &  x1079 &  x1088 &  x1091 &  x1097 &  x1106 &  x1118 &  x1121 &  x1124 & ~x234 & ~x273 & ~x561 & ~x603 & ~x735 & ~x780 & ~x867 & ~x906;
assign c6106 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x44 &  x50 &  x56 &  x59 &  x62 &  x65 &  x68 &  x77 &  x80 &  x83 &  x86 &  x89 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x119 &  x122 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x275 &  x278 &  x281 &  x284 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x347 &  x353 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x395 &  x401 &  x407 &  x410 &  x413 &  x419 &  x422 &  x425 &  x428 &  x431 &  x440 &  x443 &  x446 &  x452 &  x455 &  x461 &  x467 &  x470 &  x479 &  x485 &  x491 &  x494 &  x497 &  x500 &  x509 &  x512 &  x515 &  x518 &  x527 &  x530 &  x533 &  x536 &  x539 &  x545 &  x551 &  x554 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x584 &  x587 &  x590 &  x593 &  x596 &  x602 &  x605 &  x611 &  x614 &  x617 &  x620 &  x623 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x677 &  x680 &  x686 &  x689 &  x692 &  x698 &  x704 &  x707 &  x710 &  x713 &  x716 &  x722 &  x725 &  x728 &  x731 &  x737 &  x743 &  x746 &  x749 &  x752 &  x758 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x803 &  x806 &  x809 &  x818 &  x821 &  x824 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x854 &  x857 &  x860 &  x866 &  x869 &  x872 &  x875 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x908 &  x914 &  x917 &  x926 &  x929 &  x932 &  x935 &  x944 &  x950 &  x956 &  x962 &  x965 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1073 &  x1079 &  x1082 &  x1085 &  x1091 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 &  x1130 & ~x132 & ~x210 & ~x249 & ~x288 & ~x327 & ~x363 & ~x364 & ~x366 & ~x402 & ~x441 & ~x444 & ~x480 & ~x483 & ~x663 & ~x795 & ~x867 & ~x873 & ~x906 & ~x912;
assign c6108 =  x8 &  x14 &  x23 &  x26 &  x35 &  x44 &  x47 &  x56 &  x65 &  x68 &  x77 &  x83 &  x89 &  x98 &  x101 &  x107 &  x119 &  x125 &  x128 &  x131 &  x137 &  x140 &  x143 &  x146 &  x161 &  x164 &  x170 &  x179 &  x182 &  x185 &  x191 &  x194 &  x200 &  x209 &  x218 &  x221 &  x239 &  x242 &  x245 &  x248 &  x257 &  x263 &  x269 &  x275 &  x284 &  x287 &  x290 &  x296 &  x311 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x341 &  x344 &  x347 &  x350 &  x353 &  x365 &  x368 &  x371 &  x374 &  x380 &  x383 &  x395 &  x410 &  x413 &  x416 &  x425 &  x428 &  x431 &  x437 &  x440 &  x443 &  x449 &  x458 &  x461 &  x467 &  x470 &  x473 &  x476 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x515 &  x524 &  x527 &  x530 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x560 &  x566 &  x572 &  x575 &  x578 &  x590 &  x593 &  x599 &  x605 &  x611 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x641 &  x647 &  x653 &  x665 &  x668 &  x680 &  x683 &  x692 &  x695 &  x698 &  x701 &  x704 &  x710 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x773 &  x779 &  x788 &  x797 &  x800 &  x809 &  x824 &  x827 &  x830 &  x836 &  x839 &  x845 &  x848 &  x851 &  x857 &  x860 &  x872 &  x875 &  x878 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x911 &  x914 &  x917 &  x920 &  x929 &  x935 &  x938 &  x941 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x971 &  x980 &  x983 &  x986 &  x992 &  x1001 &  x1004 &  x1013 &  x1019 &  x1022 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1127 & ~x9 & ~x48 & ~x87 & ~x126 & ~x165 & ~x363 & ~x405 & ~x441 & ~x489 & ~x528 & ~x567 & ~x597 & ~x603 & ~x606;
assign c6110 =  x8 &  x11 &  x20 &  x25 &  x44 &  x50 &  x59 &  x62 &  x64 &  x71 &  x86 &  x92 &  x95 &  x103 &  x104 &  x113 &  x119 &  x149 &  x154 &  x158 &  x179 &  x185 &  x188 &  x191 &  x194 &  x212 &  x218 &  x224 &  x230 &  x236 &  x245 &  x248 &  x263 &  x269 &  x278 &  x281 &  x287 &  x290 &  x305 &  x308 &  x311 &  x314 &  x317 &  x334 &  x335 &  x338 &  x341 &  x350 &  x356 &  x359 &  x368 &  x373 &  x395 &  x401 &  x410 &  x416 &  x419 &  x425 &  x437 &  x443 &  x455 &  x458 &  x461 &  x470 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x503 &  x515 &  x536 &  x539 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x581 &  x596 &  x599 &  x605 &  x608 &  x614 &  x617 &  x620 &  x626 &  x632 &  x635 &  x644 &  x647 &  x659 &  x662 &  x665 &  x668 &  x689 &  x710 &  x716 &  x719 &  x722 &  x724 &  x734 &  x740 &  x743 &  x761 &  x791 &  x800 &  x806 &  x812 &  x818 &  x824 &  x833 &  x836 &  x839 &  x841 &  x851 &  x860 &  x866 &  x872 &  x878 &  x879 &  x880 &  x883 &  x893 &  x896 &  x899 &  x902 &  x905 &  x911 &  x917 &  x920 &  x922 &  x932 &  x935 &  x938 &  x944 &  x950 &  x953 &  x961 &  x962 &  x965 &  x968 &  x977 &  x980 &  x986 &  x989 &  x1000 &  x1007 &  x1025 &  x1043 &  x1046 &  x1052 &  x1067 &  x1070 &  x1073 &  x1091 &  x1100 &  x1109 &  x1121 &  x1124 &  x1127;
assign c6112 =  x2 &  x14 &  x20 &  x23 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x62 &  x65 &  x68 &  x80 &  x83 &  x86 &  x89 &  x92 &  x98 &  x104 &  x110 &  x115 &  x116 &  x128 &  x131 &  x134 &  x140 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x179 &  x182 &  x185 &  x197 &  x200 &  x203 &  x212 &  x218 &  x221 &  x227 &  x230 &  x233 &  x239 &  x242 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x302 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x335 &  x338 &  x341 &  x344 &  x350 &  x353 &  x359 &  x362 &  x368 &  x380 &  x386 &  x389 &  x392 &  x401 &  x404 &  x407 &  x410 &  x413 &  x419 &  x422 &  x425 &  x428 &  x434 &  x440 &  x443 &  x446 &  x452 &  x455 &  x458 &  x464 &  x467 &  x470 &  x473 &  x476 &  x485 &  x488 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x524 &  x527 &  x530 &  x533 &  x542 &  x548 &  x551 &  x557 &  x560 &  x563 &  x566 &  x569 &  x575 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x602 &  x605 &  x608 &  x611 &  x617 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x656 &  x662 &  x665 &  x668 &  x671 &  x680 &  x689 &  x692 &  x695 &  x698 &  x704 &  x707 &  x713 &  x716 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x809 &  x812 &  x815 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x851 &  x854 &  x860 &  x863 &  x866 &  x872 &  x875 &  x881 &  x884 &  x890 &  x896 &  x899 &  x902 &  x908 &  x911 &  x914 &  x917 &  x920 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x956 &  x959 &  x962 &  x965 &  x971 &  x977 &  x983 &  x986 &  x989 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1031 &  x1040 &  x1046 &  x1049 &  x1055 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1130 & ~x3 & ~x39 & ~x78 & ~x249 & ~x285 & ~x288 & ~x289 & ~x327 & ~x328 & ~x366 & ~x444 & ~x483 & ~x858 & ~x897 & ~x936 & ~x975 & ~x1014 & ~x1053;
assign c6114 =  x2 &  x5 &  x20 &  x26 &  x29 &  x32 &  x35 &  x44 &  x47 &  x53 &  x56 &  x62 &  x68 &  x71 &  x74 &  x77 &  x83 &  x86 &  x89 &  x92 &  x95 &  x101 &  x107 &  x113 &  x116 &  x119 &  x125 &  x128 &  x131 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x178 &  x179 &  x182 &  x185 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x239 &  x242 &  x245 &  x251 &  x254 &  x256 &  x260 &  x263 &  x266 &  x269 &  x272 &  x278 &  x281 &  x284 &  x290 &  x293 &  x295 &  x296 &  x299 &  x302 &  x305 &  x308 &  x314 &  x320 &  x323 &  x326 &  x332 &  x334 &  x335 &  x338 &  x341 &  x344 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x373 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x412 &  x413 &  x416 &  x422 &  x425 &  x431 &  x434 &  x437 &  x440 &  x443 &  x449 &  x451 &  x452 &  x455 &  x458 &  x464 &  x467 &  x470 &  x476 &  x479 &  x482 &  x485 &  x490 &  x494 &  x497 &  x506 &  x509 &  x515 &  x521 &  x524 &  x527 &  x529 &  x530 &  x533 &  x542 &  x545 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x568 &  x572 &  x575 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x656 &  x659 &  x668 &  x671 &  x674 &  x677 &  x683 &  x689 &  x692 &  x695 &  x698 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x725 &  x731 &  x734 &  x737 &  x740 &  x743 &  x752 &  x758 &  x763 &  x764 &  x773 &  x776 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x802 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x872 &  x878 &  x881 &  x884 &  x887 &  x893 &  x896 &  x899 &  x902 &  x908 &  x923 &  x926 &  x929 &  x935 &  x938 &  x941 &  x947 &  x950 &  x953 &  x958 &  x959 &  x962 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x997 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1025 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1114 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x276 & ~x357 & ~x396 & ~x825 & ~x864;
assign c6116 =  x5 &  x8 &  x11 &  x14 &  x17 &  x23 &  x35 &  x38 &  x40 &  x41 &  x44 &  x47 &  x62 &  x65 &  x68 &  x71 &  x77 &  x79 &  x80 &  x83 &  x86 &  x98 &  x104 &  x107 &  x113 &  x116 &  x118 &  x119 &  x122 &  x125 &  x134 &  x146 &  x152 &  x155 &  x158 &  x164 &  x173 &  x185 &  x191 &  x200 &  x206 &  x212 &  x217 &  x218 &  x224 &  x227 &  x229 &  x233 &  x251 &  x257 &  x260 &  x262 &  x275 &  x284 &  x293 &  x295 &  x296 &  x302 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x362 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x386 &  x392 &  x395 &  x398 &  x401 &  x407 &  x419 &  x427 &  x428 &  x431 &  x434 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x482 &  x485 &  x488 &  x494 &  x497 &  x500 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x527 &  x530 &  x536 &  x539 &  x542 &  x548 &  x551 &  x554 &  x557 &  x563 &  x569 &  x572 &  x574 &  x575 &  x581 &  x587 &  x590 &  x596 &  x605 &  x613 &  x614 &  x620 &  x623 &  x632 &  x635 &  x644 &  x650 &  x652 &  x653 &  x662 &  x668 &  x683 &  x689 &  x692 &  x701 &  x713 &  x716 &  x722 &  x731 &  x734 &  x746 &  x749 &  x752 &  x763 &  x764 &  x769 &  x770 &  x779 &  x785 &  x802 &  x806 &  x808 &  x812 &  x818 &  x821 &  x833 &  x839 &  x842 &  x848 &  x851 &  x853 &  x857 &  x863 &  x872 &  x878 &  x884 &  x887 &  x896 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x929 &  x938 &  x946 &  x950 &  x956 &  x958 &  x962 &  x965 &  x971 &  x974 &  x977 &  x986 &  x989 &  x992 &  x1004 &  x1013 &  x1019 &  x1028 &  x1031 &  x1036 &  x1037 &  x1055 &  x1067 &  x1070 &  x1073 &  x1075 &  x1076 &  x1085 &  x1088 &  x1091 &  x1100 &  x1109 &  x1112 &  x1115 &  x1121 &  x1127 & ~x354 & ~x432;
assign c6118 =  x20 &  x26 &  x29 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x83 &  x86 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x125 &  x128 &  x131 &  x134 &  x140 &  x143 &  x149 &  x158 &  x161 &  x173 &  x179 &  x182 &  x188 &  x191 &  x194 &  x203 &  x206 &  x209 &  x212 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x257 &  x260 &  x266 &  x269 &  x272 &  x278 &  x284 &  x290 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x326 &  x332 &  x337 &  x341 &  x344 &  x347 &  x350 &  x353 &  x359 &  x368 &  x371 &  x377 &  x380 &  x383 &  x386 &  x392 &  x395 &  x398 &  x401 &  x407 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x434 &  x437 &  x443 &  x446 &  x452 &  x455 &  x458 &  x464 &  x470 &  x476 &  x479 &  x482 &  x485 &  x493 &  x494 &  x503 &  x506 &  x515 &  x518 &  x524 &  x530 &  x532 &  x533 &  x536 &  x539 &  x545 &  x548 &  x551 &  x554 &  x563 &  x566 &  x569 &  x572 &  x575 &  x581 &  x584 &  x596 &  x599 &  x605 &  x608 &  x611 &  x614 &  x623 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x677 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x704 &  x719 &  x722 &  x725 &  x728 &  x734 &  x740 &  x746 &  x749 &  x752 &  x761 &  x764 &  x767 &  x770 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x803 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x832 &  x833 &  x836 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x896 &  x899 &  x902 &  x905 &  x908 &  x914 &  x917 &  x920 &  x923 &  x929 &  x935 &  x941 &  x944 &  x947 &  x953 &  x959 &  x965 &  x968 &  x974 &  x980 &  x983 &  x986 &  x989 &  x992 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1019 &  x1022 &  x1028 &  x1037 &  x1040 &  x1046 &  x1052 &  x1058 &  x1064 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1127 & ~x54 & ~x93 & ~x249 & ~x444 & ~x780 & ~x813 & ~x819 & ~x820 & ~x858 & ~x897 & ~x906;
assign c6120 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x383 &  x386 &  x389 &  x395 &  x398 &  x401 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x282 & ~x321 & ~x441 & ~x474 & ~x483 & ~x618 & ~x942 & ~x981 & ~x1080 & ~x1110 & ~x1119;
assign c6122 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x89 &  x92 &  x98 &  x101 &  x104 &  x107 &  x110 &  x119 &  x122 &  x125 &  x128 &  x131 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x260 &  x269 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x368 &  x371 &  x374 &  x380 &  x383 &  x388 &  x392 &  x395 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x500 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x542 &  x545 &  x548 &  x554 &  x557 &  x560 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x599 &  x605 &  x608 &  x611 &  x620 &  x623 &  x628 &  x629 &  x632 &  x638 &  x641 &  x644 &  x647 &  x650 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x761 &  x764 &  x767 &  x770 &  x776 &  x782 &  x785 &  x788 &  x791 &  x803 &  x809 &  x815 &  x818 &  x821 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x860 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x935 &  x938 &  x941 &  x944 &  x947 &  x953 &  x956 &  x959 &  x962 &  x968 &  x971 &  x974 &  x977 &  x980 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1025 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1079 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x72 & ~x111 & ~x195 & ~x234 & ~x273 & ~x282 & ~x441 & ~x480 & ~x483 & ~x519 & ~x522 & ~x561 & ~x597 & ~x675;
assign c6124 =  x17 &  x20 &  x26 &  x32 &  x38 &  x41 &  x47 &  x56 &  x59 &  x77 &  x80 &  x89 &  x95 &  x110 &  x113 &  x119 &  x131 &  x140 &  x143 &  x146 &  x149 &  x158 &  x161 &  x164 &  x167 &  x170 &  x179 &  x185 &  x191 &  x197 &  x203 &  x206 &  x209 &  x212 &  x218 &  x221 &  x227 &  x230 &  x233 &  x236 &  x239 &  x248 &  x257 &  x260 &  x263 &  x272 &  x275 &  x278 &  x281 &  x287 &  x293 &  x299 &  x308 &  x311 &  x316 &  x317 &  x323 &  x326 &  x332 &  x341 &  x344 &  x347 &  x353 &  x355 &  x356 &  x362 &  x368 &  x386 &  x392 &  x401 &  x407 &  x410 &  x422 &  x428 &  x431 &  x449 &  x452 &  x461 &  x467 &  x470 &  x476 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x503 &  x509 &  x515 &  x524 &  x533 &  x539 &  x557 &  x566 &  x569 &  x575 &  x578 &  x584 &  x593 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x632 &  x635 &  x638 &  x641 &  x656 &  x659 &  x668 &  x674 &  x677 &  x683 &  x689 &  x692 &  x707 &  x710 &  x716 &  x722 &  x731 &  x746 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x779 &  x782 &  x788 &  x794 &  x800 &  x806 &  x809 &  x818 &  x821 &  x824 &  x827 &  x832 &  x833 &  x836 &  x863 &  x869 &  x872 &  x875 &  x883 &  x893 &  x896 &  x908 &  x910 &  x917 &  x922 &  x923 &  x926 &  x944 &  x947 &  x950 &  x956 &  x962 &  x968 &  x983 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1019 &  x1022 &  x1034 &  x1039 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1064 &  x1067 &  x1070 &  x1073 &  x1082 &  x1085 &  x1091 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 & ~x54 & ~x132 & ~x171 & ~x213 & ~x246 & ~x249 & ~x285 & ~x324 & ~x363 & ~x627 & ~x858 & ~x936;
assign c6126 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x26 &  x35 &  x38 &  x41 &  x47 &  x50 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x104 &  x110 &  x119 &  x125 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x155 &  x158 &  x164 &  x170 &  x173 &  x176 &  x188 &  x191 &  x197 &  x200 &  x209 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x242 &  x245 &  x248 &  x251 &  x257 &  x263 &  x266 &  x269 &  x275 &  x281 &  x284 &  x287 &  x293 &  x296 &  x311 &  x320 &  x323 &  x332 &  x335 &  x338 &  x341 &  x344 &  x350 &  x353 &  x359 &  x362 &  x368 &  x371 &  x374 &  x376 &  x377 &  x383 &  x389 &  x392 &  x395 &  x401 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x428 &  x434 &  x440 &  x443 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x479 &  x488 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x524 &  x536 &  x539 &  x542 &  x545 &  x554 &  x557 &  x560 &  x563 &  x566 &  x572 &  x575 &  x587 &  x590 &  x593 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x626 &  x629 &  x635 &  x638 &  x641 &  x644 &  x653 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x713 &  x716 &  x719 &  x722 &  x725 &  x731 &  x737 &  x743 &  x746 &  x752 &  x755 &  x758 &  x764 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x797 &  x809 &  x815 &  x818 &  x821 &  x824 &  x827 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x863 &  x872 &  x875 &  x881 &  x884 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x917 &  x923 &  x929 &  x932 &  x941 &  x947 &  x950 &  x953 &  x959 &  x965 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1043 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1079 &  x1088 &  x1091 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 & ~x78 & ~x234 & ~x273 & ~x282 & ~x480 & ~x513 & ~x519 & ~x636 & ~x1014 & ~x1053;
assign c6128 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x583 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x901 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x940 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1018 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1057 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1096 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x165 & ~x399 & ~x405 & ~x438 & ~x477 & ~x516 & ~x555 & ~x594 & ~x633 & ~x714 & ~x753 & ~x792 & ~x831;
assign c6130 =  x8 &  x11 &  x20 &  x23 &  x26 &  x32 &  x35 &  x38 &  x47 &  x50 &  x68 &  x74 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x125 &  x146 &  x149 &  x158 &  x161 &  x164 &  x167 &  x170 &  x176 &  x179 &  x182 &  x191 &  x203 &  x209 &  x212 &  x218 &  x233 &  x239 &  x242 &  x257 &  x260 &  x269 &  x275 &  x278 &  x287 &  x290 &  x299 &  x308 &  x320 &  x332 &  x335 &  x338 &  x356 &  x359 &  x365 &  x368 &  x374 &  x377 &  x389 &  x410 &  x413 &  x425 &  x428 &  x431 &  x437 &  x443 &  x452 &  x455 &  x458 &  x461 &  x467 &  x476 &  x479 &  x491 &  x497 &  x503 &  x509 &  x515 &  x518 &  x521 &  x524 &  x530 &  x536 &  x542 &  x548 &  x557 &  x575 &  x581 &  x587 &  x596 &  x599 &  x602 &  x605 &  x608 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x635 &  x644 &  x647 &  x653 &  x662 &  x668 &  x671 &  x680 &  x683 &  x686 &  x689 &  x695 &  x698 &  x710 &  x722 &  x725 &  x731 &  x734 &  x737 &  x740 &  x752 &  x758 &  x761 &  x764 &  x767 &  x770 &  x776 &  x782 &  x785 &  x803 &  x806 &  x812 &  x821 &  x824 &  x830 &  x833 &  x839 &  x848 &  x854 &  x857 &  x866 &  x869 &  x872 &  x878 &  x896 &  x905 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x938 &  x944 &  x950 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x977 &  x983 &  x986 &  x992 &  x995 &  x1001 &  x1013 &  x1022 &  x1025 &  x1037 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1112 &  x1121 &  x1127 & ~x27 & ~x54 & ~x132 & ~x171 & ~x210 & ~x501 & ~x540 & ~x546 & ~x579 & ~x580 & ~x585 & ~x618 & ~x625 & ~x672;
assign c6132 =  x5 &  x14 &  x17 &  x20 &  x32 &  x35 &  x38 &  x47 &  x53 &  x62 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x170 &  x173 &  x176 &  x179 &  x182 &  x188 &  x191 &  x197 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x284 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x326 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x389 &  x392 &  x395 &  x398 &  x401 &  x410 &  x416 &  x419 &  x422 &  x428 &  x434 &  x443 &  x446 &  x461 &  x464 &  x470 &  x473 &  x476 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x512 &  x515 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x548 &  x554 &  x557 &  x560 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x629 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x665 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x695 &  x707 &  x710 &  x713 &  x719 &  x722 &  x725 &  x728 &  x731 &  x740 &  x749 &  x752 &  x755 &  x758 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x797 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x902 &  x905 &  x908 &  x917 &  x923 &  x926 &  x935 &  x938 &  x944 &  x953 &  x956 &  x962 &  x968 &  x971 &  x977 &  x980 &  x989 &  x992 &  x998 &  x1004 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1082 &  x1088 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 & ~x132 & ~x171 & ~x306 & ~x429 & ~x438 & ~x468 & ~x510 & ~x756 & ~x795 & ~x846 & ~x873 & ~x885 & ~x912 & ~x924 & ~x951 & ~x963 & ~x1002 & ~x1041 & ~x1062 & ~x1119;
assign c6134 =  x5 &  x14 &  x23 &  x29 &  x32 &  x41 &  x44 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x77 &  x80 &  x86 &  x104 &  x107 &  x110 &  x113 &  x116 &  x125 &  x128 &  x131 &  x134 &  x140 &  x143 &  x146 &  x149 &  x161 &  x167 &  x173 &  x176 &  x179 &  x181 &  x191 &  x193 &  x194 &  x197 &  x200 &  x203 &  x206 &  x215 &  x218 &  x221 &  x227 &  x232 &  x233 &  x239 &  x242 &  x248 &  x251 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x293 &  x296 &  x298 &  x299 &  x302 &  x308 &  x314 &  x326 &  x332 &  x337 &  x338 &  x341 &  x344 &  x347 &  x350 &  x359 &  x365 &  x368 &  x374 &  x377 &  x380 &  x383 &  x389 &  x392 &  x395 &  x398 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x458 &  x461 &  x479 &  x482 &  x488 &  x497 &  x500 &  x503 &  x506 &  x515 &  x518 &  x521 &  x527 &  x533 &  x536 &  x557 &  x563 &  x566 &  x569 &  x575 &  x581 &  x587 &  x589 &  x596 &  x602 &  x605 &  x608 &  x614 &  x620 &  x623 &  x626 &  x629 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x680 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x788 &  x794 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x824 &  x830 &  x833 &  x839 &  x842 &  x845 &  x848 &  x857 &  x860 &  x866 &  x875 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x902 &  x908 &  x914 &  x917 &  x920 &  x926 &  x932 &  x935 &  x941 &  x944 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1064 &  x1076 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1115 &  x1117 &  x1118 & ~x195 & ~x523 & ~x561 & ~x562 & ~x600 & ~x819 & ~x975;
assign c6136 =  x5 &  x11 &  x20 &  x23 &  x56 &  x77 &  x80 &  x83 &  x98 &  x101 &  x125 &  x127 &  x158 &  x161 &  x167 &  x176 &  x182 &  x185 &  x188 &  x203 &  x209 &  x221 &  x223 &  x278 &  x283 &  x287 &  x293 &  x298 &  x301 &  x302 &  x305 &  x323 &  x325 &  x326 &  x328 &  x334 &  x335 &  x343 &  x344 &  x361 &  x374 &  x380 &  x383 &  x398 &  x410 &  x422 &  x437 &  x443 &  x452 &  x454 &  x461 &  x494 &  x533 &  x536 &  x542 &  x551 &  x590 &  x593 &  x596 &  x611 &  x620 &  x634 &  x647 &  x650 &  x653 &  x662 &  x686 &  x701 &  x710 &  x712 &  x728 &  x749 &  x751 &  x776 &  x785 &  x790 &  x797 &  x800 &  x809 &  x812 &  x827 &  x857 &  x868 &  x878 &  x886 &  x890 &  x907 &  x950 &  x968 &  x998 &  x1004 &  x1016 &  x1034 &  x1043 &  x1064 &  x1070 &  x1073 &  x1082 &  x1085 &  x1094 &  x1103 &  x1114 &  x1124;
assign c6138 =  x5 &  x11 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x59 &  x62 &  x68 &  x74 &  x79 &  x83 &  x86 &  x89 &  x92 &  x95 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x134 &  x140 &  x143 &  x152 &  x155 &  x158 &  x161 &  x167 &  x173 &  x182 &  x191 &  x194 &  x200 &  x203 &  x206 &  x215 &  x227 &  x233 &  x245 &  x248 &  x251 &  x254 &  x257 &  x269 &  x281 &  x287 &  x299 &  x302 &  x305 &  x317 &  x320 &  x322 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x350 &  x356 &  x359 &  x371 &  x374 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x404 &  x407 &  x410 &  x419 &  x421 &  x422 &  x431 &  x443 &  x446 &  x449 &  x455 &  x461 &  x473 &  x479 &  x482 &  x488 &  x491 &  x494 &  x500 &  x503 &  x512 &  x521 &  x527 &  x530 &  x533 &  x542 &  x545 &  x548 &  x554 &  x557 &  x560 &  x569 &  x571 &  x572 &  x587 &  x602 &  x608 &  x617 &  x623 &  x635 &  x641 &  x650 &  x659 &  x665 &  x683 &  x698 &  x701 &  x707 &  x710 &  x713 &  x731 &  x734 &  x746 &  x755 &  x758 &  x767 &  x773 &  x776 &  x782 &  x794 &  x797 &  x800 &  x802 &  x803 &  x812 &  x815 &  x827 &  x830 &  x842 &  x851 &  x854 &  x860 &  x866 &  x869 &  x872 &  x880 &  x893 &  x896 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x938 &  x941 &  x947 &  x950 &  x956 &  x962 &  x965 &  x968 &  x980 &  x983 &  x986 &  x992 &  x1001 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1040 &  x1043 &  x1049 &  x1052 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1097 &  x1100 &  x1103 &  x1112 &  x1115 &  x1121 &  x1124 & ~x90 & ~x96 & ~x225 & ~x627;
assign c6140 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x26 &  x29 &  x38 &  x41 &  x44 &  x50 &  x59 &  x65 &  x71 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x119 &  x122 &  x125 &  x137 &  x140 &  x143 &  x149 &  x155 &  x158 &  x161 &  x164 &  x170 &  x179 &  x182 &  x185 &  x188 &  x194 &  x200 &  x203 &  x215 &  x218 &  x220 &  x221 &  x224 &  x227 &  x230 &  x236 &  x242 &  x245 &  x248 &  x251 &  x254 &  x259 &  x260 &  x263 &  x272 &  x275 &  x278 &  x287 &  x290 &  x293 &  x302 &  x305 &  x311 &  x314 &  x317 &  x319 &  x329 &  x332 &  x335 &  x337 &  x347 &  x350 &  x356 &  x359 &  x365 &  x368 &  x371 &  x377 &  x380 &  x386 &  x389 &  x395 &  x401 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x425 &  x437 &  x440 &  x443 &  x449 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x476 &  x479 &  x482 &  x488 &  x491 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x545 &  x554 &  x557 &  x563 &  x566 &  x569 &  x578 &  x587 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x626 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x683 &  x686 &  x689 &  x692 &  x707 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x743 &  x746 &  x752 &  x755 &  x758 &  x761 &  x770 &  x773 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x845 &  x851 &  x854 &  x860 &  x875 &  x878 &  x880 &  x881 &  x887 &  x890 &  x896 &  x902 &  x905 &  x908 &  x911 &  x914 &  x920 &  x938 &  x950 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x989 &  x995 &  x1001 &  x1004 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1040 &  x1043 &  x1052 &  x1055 &  x1061 &  x1067 &  x1073 &  x1076 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1106 &  x1115 &  x1127 &  x1130 & ~x78 & ~x234 & ~x273 & ~x399 & ~x483 & ~x561 & ~x678;
assign c6142 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x155 &  x158 &  x161 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x280 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x310 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x419 &  x422 &  x425 &  x428 &  x431 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x497 &  x500 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x593 &  x596 &  x599 &  x605 &  x608 &  x611 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x911 &  x914 &  x917 &  x920 &  x926 &  x929 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x968 &  x971 &  x977 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 &  x1130 & ~x126 & ~x195 & ~x204 & ~x234 & ~x243 & ~x273 & ~x282 & ~x321 & ~x405 & ~x444 & ~x483 & ~x522 & ~x561 & ~x600 & ~x678 & ~x702 & ~x741;
assign c6144 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1045 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x156 & ~x195 & ~x198 & ~x402 & ~x441 & ~x666 & ~x705 & ~x744 & ~x783 & ~x822 & ~x897 & ~x936 & ~x975 & ~x1014 & ~x1053 & ~x1092;
assign c6146 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x263 &  x272 &  x275 &  x278 &  x281 &  x284 &  x290 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x317 &  x320 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x368 &  x371 &  x374 &  x377 &  x383 &  x386 &  x389 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x434 &  x440 &  x443 &  x449 &  x455 &  x458 &  x461 &  x464 &  x466 &  x467 &  x473 &  x476 &  x479 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x521 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x650 &  x653 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x695 &  x698 &  x701 &  x704 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x740 &  x743 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x857 &  x860 &  x863 &  x869 &  x881 &  x884 &  x887 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x351 & ~x390 & ~x405 & ~x429 & ~x430 & ~x438 & ~x444 & ~x468 & ~x477 & ~x507 & ~x516 & ~x594 & ~x756 & ~x951 & ~x981 & ~x984;
assign c6148 =  x2 &  x5 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x71 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x176 &  x179 &  x182 &  x185 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x281 &  x284 &  x287 &  x291 &  x292 &  x293 &  x296 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x323 &  x326 &  x329 &  x332 &  x335 &  x341 &  x344 &  x350 &  x353 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x380 &  x383 &  x386 &  x388 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x466 &  x467 &  x470 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x611 &  x614 &  x617 &  x623 &  x626 &  x629 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x662 &  x668 &  x671 &  x674 &  x677 &  x680 &  x686 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x737 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x884 &  x887 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x977 &  x980 &  x983 &  x986 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1055 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1111 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x273 & ~x276 & ~x312 & ~x639 & ~x678 & ~x717;
assign c6150 =  x2 &  x5 &  x11 &  x14 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x50 &  x56 &  x58 &  x59 &  x62 &  x65 &  x68 &  x74 &  x77 &  x83 &  x89 &  x92 &  x95 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x131 &  x134 &  x137 &  x140 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x173 &  x175 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x206 &  x212 &  x215 &  x218 &  x221 &  x224 &  x233 &  x239 &  x242 &  x245 &  x248 &  x251 &  x257 &  x260 &  x263 &  x266 &  x272 &  x281 &  x284 &  x290 &  x293 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x329 &  x332 &  x347 &  x350 &  x356 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x380 &  x383 &  x386 &  x392 &  x398 &  x401 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x485 &  x491 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x572 &  x575 &  x578 &  x584 &  x587 &  x590 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x656 &  x659 &  x662 &  x668 &  x671 &  x677 &  x680 &  x683 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x713 &  x716 &  x719 &  x725 &  x728 &  x731 &  x734 &  x737 &  x743 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x866 &  x872 &  x878 &  x881 &  x884 &  x890 &  x893 &  x896 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x940 &  x941 &  x950 &  x959 &  x962 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1016 &  x1018 &  x1019 &  x1025 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1070 &  x1073 &  x1076 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x78 & ~x156 & ~x195 & ~x321 & ~x327 & ~x366 & ~x405 & ~x444 & ~x483 & ~x600 & ~x678 & ~x1092;
assign c6152 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x386 &  x388 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x485 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x548 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x596 &  x599 &  x605 &  x608 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x273 & ~x321 & ~x360 & ~x399 & ~x438 & ~x477 & ~x639 & ~x642 & ~x678 & ~x717 & ~x756 & ~x759 & ~x795 & ~x798 & ~x924;
assign c6154 =  x1 &  x5 &  x8 &  x11 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x40 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x110 &  x116 &  x119 &  x128 &  x137 &  x140 &  x143 &  x146 &  x151 &  x152 &  x155 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x188 &  x191 &  x200 &  x212 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x260 &  x263 &  x266 &  x275 &  x284 &  x290 &  x293 &  x296 &  x302 &  x305 &  x307 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x335 &  x338 &  x341 &  x344 &  x350 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x395 &  x407 &  x413 &  x416 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x464 &  x470 &  x476 &  x482 &  x485 &  x488 &  x490 &  x494 &  x497 &  x500 &  x503 &  x509 &  x512 &  x518 &  x521 &  x524 &  x527 &  x529 &  x533 &  x539 &  x542 &  x545 &  x551 &  x554 &  x563 &  x566 &  x568 &  x569 &  x572 &  x575 &  x580 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x607 &  x608 &  x611 &  x614 &  x617 &  x619 &  x620 &  x623 &  x626 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x671 &  x677 &  x683 &  x685 &  x686 &  x689 &  x692 &  x697 &  x698 &  x701 &  x704 &  x710 &  x713 &  x719 &  x724 &  x725 &  x731 &  x734 &  x736 &  x737 &  x740 &  x743 &  x746 &  x758 &  x760 &  x763 &  x764 &  x773 &  x775 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x806 &  x809 &  x812 &  x814 &  x815 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x851 &  x857 &  x863 &  x866 &  x878 &  x881 &  x890 &  x899 &  x905 &  x908 &  x911 &  x914 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x953 &  x956 &  x959 &  x962 &  x965 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1019 &  x1022 &  x1025 &  x1034 &  x1037 &  x1043 &  x1049 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1075 &  x1076 &  x1079 &  x1082 &  x1085 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x51 & ~x90 & ~x321 & ~x360 & ~x399;
assign c6156 =  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x59 &  x62 &  x68 &  x71 &  x74 &  x77 &  x80 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x140 &  x143 &  x146 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x251 &  x260 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x349 &  x353 &  x356 &  x359 &  x362 &  x368 &  x371 &  x374 &  x380 &  x386 &  x395 &  x401 &  x404 &  x407 &  x409 &  x410 &  x416 &  x419 &  x422 &  x425 &  x431 &  x434 &  x440 &  x446 &  x448 &  x449 &  x452 &  x458 &  x464 &  x466 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x509 &  x512 &  x515 &  x518 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x551 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x587 &  x593 &  x596 &  x605 &  x608 &  x614 &  x617 &  x620 &  x623 &  x626 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x779 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x809 &  x812 &  x815 &  x818 &  x827 &  x833 &  x836 &  x839 &  x842 &  x845 &  x851 &  x854 &  x860 &  x863 &  x866 &  x875 &  x878 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x914 &  x917 &  x920 &  x923 &  x932 &  x935 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x962 &  x965 &  x968 &  x971 &  x977 &  x980 &  x983 &  x986 &  x995 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x156 & ~x195 & ~x234 & ~x273 & ~x312 & ~x351 & ~x354 & ~x390 & ~x391 & ~x393 & ~x429 & ~x522 & ~x561 & ~x600 & ~x639 & ~x678 & ~x717 & ~x756 & ~x795 & ~x831;
assign c6158 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x26 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x155 &  x158 &  x164 &  x167 &  x170 &  x173 &  x176 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x353 &  x355 &  x356 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x422 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x458 &  x461 &  x464 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x584 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x698 &  x701 &  x704 &  x710 &  x713 &  x719 &  x721 &  x725 &  x728 &  x731 &  x733 &  x734 &  x737 &  x740 &  x749 &  x752 &  x755 &  x758 &  x761 &  x770 &  x776 &  x782 &  x785 &  x788 &  x794 &  x797 &  x799 &  x800 &  x803 &  x806 &  x809 &  x811 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x850 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x916 &  x917 &  x920 &  x923 &  x926 &  x928 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x955 &  x956 &  x959 &  x961 &  x962 &  x965 &  x967 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x988 &  x989 &  x992 &  x994 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1090 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x93 & ~x213 & ~x291 & ~x663 & ~x666 & ~x705 & ~x741 & ~x780 & ~x783 & ~x789 & ~x819 & ~x822 & ~x858 & ~x897 & ~x936 & ~x975 & ~x1014 & ~x1053;
assign c6160 =  x1 &  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x40 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x67 &  x68 &  x71 &  x74 &  x77 &  x79 &  x83 &  x86 &  x92 &  x95 &  x101 &  x104 &  x106 &  x107 &  x110 &  x113 &  x116 &  x118 &  x119 &  x122 &  x125 &  x128 &  x134 &  x137 &  x140 &  x145 &  x146 &  x149 &  x152 &  x161 &  x164 &  x167 &  x170 &  x176 &  x179 &  x182 &  x188 &  x191 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x254 &  x257 &  x260 &  x266 &  x272 &  x274 &  x275 &  x281 &  x284 &  x290 &  x296 &  x299 &  x305 &  x308 &  x311 &  x313 &  x314 &  x320 &  x323 &  x335 &  x338 &  x341 &  x350 &  x352 &  x365 &  x368 &  x374 &  x377 &  x380 &  x383 &  x389 &  x391 &  x395 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x419 &  x422 &  x428 &  x430 &  x431 &  x434 &  x437 &  x443 &  x446 &  x449 &  x452 &  x455 &  x464 &  x467 &  x469 &  x473 &  x476 &  x482 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x548 &  x551 &  x554 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x623 &  x626 &  x632 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x716 &  x722 &  x725 &  x728 &  x731 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x760 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x785 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x848 &  x854 &  x857 &  x860 &  x866 &  x869 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x971 &  x974 &  x977 &  x983 &  x986 &  x998 &  x1001 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1058 &  x1064 &  x1067 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x285 & ~x303 & ~x342 & ~x363 & ~x402 & ~x1011 & ~x1032 & ~x1044 & ~x1071 & ~x1110 & ~x1122 & ~x1128;
assign c6162 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x271 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x292 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x331 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x349 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x529 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x931 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x399 & ~x438 & ~x477 & ~x516 & ~x597 & ~x636 & ~x675;
assign c6164 =  x2 &  x5 &  x8 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x50 &  x53 &  x56 &  x59 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x128 &  x134 &  x137 &  x140 &  x143 &  x146 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x191 &  x194 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x251 &  x254 &  x257 &  x263 &  x266 &  x269 &  x272 &  x275 &  x281 &  x284 &  x290 &  x293 &  x299 &  x302 &  x308 &  x311 &  x314 &  x317 &  x320 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x356 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x398 &  x401 &  x404 &  x407 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x446 &  x449 &  x452 &  x458 &  x461 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x494 &  x497 &  x500 &  x506 &  x509 &  x515 &  x518 &  x530 &  x536 &  x539 &  x551 &  x554 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x578 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x614 &  x617 &  x620 &  x623 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x661 &  x665 &  x677 &  x683 &  x686 &  x695 &  x698 &  x700 &  x701 &  x713 &  x716 &  x719 &  x722 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x767 &  x773 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x827 &  x833 &  x836 &  x839 &  x842 &  x848 &  x851 &  x854 &  x857 &  x863 &  x866 &  x872 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x902 &  x905 &  x908 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x327 & ~x438 & ~x468 & ~x477 & ~x507 & ~x516 & ~x546 & ~x549 & ~x555 & ~x585 & ~x594 & ~x624 & ~x951 & ~x990 & ~x1029 & ~x1068 & ~x1104 & ~x1107;
assign c6166 =  x2 &  x5 &  x8 &  x11 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x368 &  x371 &  x374 &  x377 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x491 &  x494 &  x497 &  x500 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x688 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x731 &  x734 &  x740 &  x743 &  x746 &  x749 &  x755 &  x758 &  x760 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x893 &  x896 &  x902 &  x908 &  x911 &  x917 &  x920 &  x922 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x965 &  x971 &  x974 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1123 &  x1124 &  x1127 &  x1130 & ~x285 & ~x288 & ~x324 & ~x396 & ~x441 & ~x783 & ~x858 & ~x861 & ~x897 & ~x900 & ~x936 & ~x939 & ~x1053 & ~x1092;
assign c6168 =  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x83 &  x86 &  x89 &  x92 &  x98 &  x101 &  x104 &  x107 &  x113 &  x122 &  x125 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x161 &  x167 &  x170 &  x176 &  x182 &  x185 &  x188 &  x197 &  x200 &  x206 &  x209 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x257 &  x260 &  x263 &  x266 &  x268 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x293 &  x299 &  x305 &  x307 &  x308 &  x311 &  x320 &  x326 &  x329 &  x335 &  x338 &  x343 &  x344 &  x346 &  x347 &  x350 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x376 &  x377 &  x380 &  x382 &  x386 &  x389 &  x395 &  x398 &  x401 &  x404 &  x410 &  x413 &  x415 &  x416 &  x419 &  x422 &  x425 &  x428 &  x434 &  x440 &  x443 &  x446 &  x449 &  x452 &  x454 &  x455 &  x464 &  x466 &  x467 &  x482 &  x488 &  x491 &  x493 &  x494 &  x497 &  x500 &  x502 &  x503 &  x505 &  x506 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x581 &  x584 &  x587 &  x590 &  x593 &  x599 &  x605 &  x608 &  x611 &  x614 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x646 &  x647 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x680 &  x683 &  x692 &  x695 &  x698 &  x701 &  x710 &  x716 &  x719 &  x722 &  x725 &  x728 &  x734 &  x737 &  x740 &  x743 &  x749 &  x752 &  x755 &  x758 &  x761 &  x770 &  x776 &  x779 &  x782 &  x788 &  x791 &  x794 &  x800 &  x818 &  x821 &  x824 &  x827 &  x830 &  x836 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x875 &  x878 &  x887 &  x890 &  x893 &  x896 &  x902 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x938 &  x941 &  x944 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1022 &  x1025 &  x1031 &  x1034 &  x1043 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1109 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x591 & ~x717;
assign c6170 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x466 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x497 &  x500 &  x503 &  x505 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x312 & ~x351 & ~x354 & ~x393 & ~x561 & ~x600 & ~x601 & ~x639 & ~x675 & ~x678 & ~x714 & ~x717;
assign c6172 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x50 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x202 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x488 &  x491 &  x494 &  x500 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x689 &  x692 &  x698 &  x701 &  x704 &  x707 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x766 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x799 &  x803 &  x805 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x838 &  x839 &  x842 &  x844 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x871 &  x872 &  x875 &  x877 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x922 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x961 &  x962 &  x965 &  x968 &  x971 &  x974 &  x980 &  x983 &  x986 &  x988 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x249 & ~x402 & ~x480 & ~x519 & ~x663 & ~x702 & ~x741 & ~x780 & ~x858 & ~x897 & ~x936 & ~x975 & ~x1014 & ~x1053;
assign c6174 =  x2 &  x5 &  x8 &  x14 &  x20 &  x26 &  x29 &  x32 &  x38 &  x44 &  x50 &  x56 &  x59 &  x65 &  x68 &  x77 &  x83 &  x86 &  x95 &  x98 &  x107 &  x113 &  x116 &  x119 &  x122 &  x125 &  x131 &  x134 &  x140 &  x146 &  x152 &  x155 &  x158 &  x161 &  x167 &  x173 &  x179 &  x182 &  x188 &  x191 &  x197 &  x203 &  x206 &  x209 &  x218 &  x221 &  x224 &  x227 &  x230 &  x239 &  x242 &  x254 &  x257 &  x263 &  x272 &  x281 &  x284 &  x299 &  x302 &  x305 &  x311 &  x314 &  x323 &  x326 &  x329 &  x332 &  x338 &  x344 &  x350 &  x362 &  x365 &  x368 &  x371 &  x377 &  x386 &  x392 &  x395 &  x401 &  x404 &  x416 &  x419 &  x434 &  x440 &  x443 &  x458 &  x470 &  x482 &  x485 &  x494 &  x503 &  x509 &  x518 &  x521 &  x527 &  x533 &  x542 &  x548 &  x551 &  x554 &  x569 &  x578 &  x581 &  x584 &  x587 &  x596 &  x602 &  x605 &  x608 &  x611 &  x623 &  x626 &  x629 &  x632 &  x650 &  x653 &  x656 &  x662 &  x668 &  x671 &  x674 &  x677 &  x680 &  x688 &  x689 &  x695 &  x713 &  x725 &  x728 &  x734 &  x737 &  x740 &  x743 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x773 &  x776 &  x779 &  x782 &  x788 &  x791 &  x797 &  x806 &  x809 &  x824 &  x827 &  x833 &  x836 &  x842 &  x848 &  x860 &  x863 &  x866 &  x869 &  x881 &  x884 &  x890 &  x893 &  x896 &  x899 &  x908 &  x911 &  x914 &  x920 &  x926 &  x935 &  x938 &  x947 &  x959 &  x962 &  x965 &  x968 &  x974 &  x980 &  x992 &  x995 &  x1001 &  x1007 &  x1016 &  x1022 &  x1025 &  x1031 &  x1034 &  x1040 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1082 &  x1085 &  x1097 &  x1109 &  x1112 &  x1115 &  x1124 &  x1127 &  x1130 & ~x195 & ~x210 & ~x249 & ~x288 & ~x327 & ~x405 & ~x522 & ~x624 & ~x885 & ~x918 & ~x1014 & ~x1047;
assign c6176 =  x2 &  x11 &  x26 &  x29 &  x32 &  x35 &  x41 &  x47 &  x53 &  x56 &  x59 &  x65 &  x68 &  x71 &  x77 &  x83 &  x86 &  x92 &  x98 &  x101 &  x104 &  x110 &  x116 &  x119 &  x122 &  x128 &  x131 &  x134 &  x140 &  x143 &  x155 &  x158 &  x161 &  x167 &  x176 &  x188 &  x191 &  x194 &  x197 &  x218 &  x221 &  x227 &  x230 &  x239 &  x242 &  x245 &  x248 &  x254 &  x257 &  x263 &  x266 &  x275 &  x281 &  x283 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x301 &  x305 &  x314 &  x317 &  x320 &  x323 &  x332 &  x335 &  x341 &  x356 &  x359 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x386 &  x389 &  x395 &  x398 &  x410 &  x413 &  x421 &  x425 &  x428 &  x431 &  x443 &  x449 &  x452 &  x458 &  x460 &  x463 &  x464 &  x466 &  x467 &  x479 &  x482 &  x491 &  x494 &  x505 &  x506 &  x509 &  x512 &  x515 &  x518 &  x524 &  x527 &  x533 &  x539 &  x542 &  x545 &  x548 &  x554 &  x560 &  x563 &  x572 &  x575 &  x581 &  x587 &  x590 &  x593 &  x596 &  x599 &  x605 &  x608 &  x611 &  x614 &  x617 &  x623 &  x632 &  x635 &  x644 &  x646 &  x653 &  x665 &  x671 &  x674 &  x677 &  x680 &  x683 &  x685 &  x686 &  x689 &  x695 &  x704 &  x707 &  x710 &  x719 &  x724 &  x725 &  x728 &  x734 &  x752 &  x755 &  x758 &  x763 &  x764 &  x769 &  x779 &  x788 &  x797 &  x800 &  x803 &  x809 &  x815 &  x818 &  x821 &  x827 &  x833 &  x836 &  x848 &  x851 &  x857 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x890 &  x896 &  x899 &  x902 &  x911 &  x914 &  x920 &  x923 &  x932 &  x950 &  x953 &  x958 &  x959 &  x962 &  x965 &  x968 &  x977 &  x983 &  x989 &  x995 &  x997 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1024 &  x1034 &  x1036 &  x1037 &  x1042 &  x1048 &  x1049 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1075 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1097 &  x1106 &  x1109 &  x1112 &  x1114 &  x1115 &  x1121 &  x1124 &  x1127;
assign c6178 =  x5 &  x8 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x191 &  x194 &  x197 &  x203 &  x209 &  x212 &  x215 &  x218 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x260 &  x263 &  x269 &  x275 &  x287 &  x290 &  x293 &  x299 &  x302 &  x305 &  x308 &  x317 &  x320 &  x329 &  x337 &  x338 &  x341 &  x347 &  x350 &  x353 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x380 &  x383 &  x386 &  x389 &  x395 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x431 &  x437 &  x440 &  x446 &  x452 &  x455 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x554 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x581 &  x584 &  x587 &  x593 &  x596 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x667 &  x671 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x716 &  x719 &  x722 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x788 &  x791 &  x794 &  x797 &  x806 &  x812 &  x818 &  x821 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x899 &  x902 &  x905 &  x908 &  x911 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x938 &  x944 &  x947 &  x950 &  x953 &  x956 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x979 &  x983 &  x986 &  x989 &  x995 &  x1001 &  x1007 &  x1016 &  x1018 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1070 &  x1073 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1100 &  x1106 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 & ~x273 & ~x405 & ~x600 & ~x636 & ~x675 & ~x678 & ~x714 & ~x717 & ~x753 & ~x756 & ~x792 & ~x795 & ~x810 & ~x831 & ~x834;
assign c6180 =  x2 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x83 &  x86 &  x92 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x146 &  x149 &  x152 &  x158 &  x161 &  x164 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x209 &  x212 &  x215 &  x218 &  x220 &  x221 &  x224 &  x227 &  x230 &  x233 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x293 &  x296 &  x302 &  x305 &  x311 &  x314 &  x317 &  x320 &  x329 &  x335 &  x338 &  x341 &  x344 &  x347 &  x349 &  x350 &  x353 &  x356 &  x359 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x386 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x488 &  x491 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x649 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x686 &  x688 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x746 &  x749 &  x752 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x805 &  x806 &  x812 &  x818 &  x821 &  x824 &  x827 &  x833 &  x836 &  x842 &  x844 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x875 &  x878 &  x881 &  x884 &  x887 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x923 &  x926 &  x929 &  x935 &  x938 &  x941 &  x944 &  x950 &  x953 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x980 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1051 &  x1052 &  x1058 &  x1061 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130 & ~x147 & ~x720;
assign c6182 =  x11 &  x14 &  x17 &  x29 &  x35 &  x47 &  x50 &  x59 &  x62 &  x74 &  x83 &  x86 &  x89 &  x92 &  x110 &  x113 &  x116 &  x119 &  x143 &  x146 &  x164 &  x167 &  x170 &  x182 &  x188 &  x203 &  x206 &  x209 &  x233 &  x236 &  x248 &  x254 &  x257 &  x263 &  x269 &  x278 &  x281 &  x284 &  x290 &  x308 &  x311 &  x332 &  x347 &  x350 &  x368 &  x374 &  x377 &  x389 &  x392 &  x395 &  x398 &  x401 &  x407 &  x410 &  x416 &  x425 &  x434 &  x446 &  x455 &  x458 &  x461 &  x467 &  x473 &  x476 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x506 &  x518 &  x530 &  x536 &  x539 &  x545 &  x551 &  x560 &  x566 &  x578 &  x587 &  x593 &  x599 &  x602 &  x605 &  x608 &  x617 &  x626 &  x632 &  x656 &  x665 &  x677 &  x686 &  x695 &  x698 &  x704 &  x728 &  x737 &  x743 &  x746 &  x752 &  x755 &  x758 &  x764 &  x767 &  x770 &  x785 &  x794 &  x800 &  x803 &  x806 &  x809 &  x818 &  x830 &  x833 &  x836 &  x842 &  x848 &  x857 &  x860 &  x869 &  x872 &  x884 &  x887 &  x890 &  x893 &  x902 &  x917 &  x920 &  x923 &  x935 &  x944 &  x953 &  x959 &  x962 &  x965 &  x971 &  x974 &  x977 &  x983 &  x986 &  x992 &  x995 &  x1004 &  x1010 &  x1019 &  x1031 &  x1043 &  x1046 &  x1055 &  x1058 &  x1064 &  x1070 &  x1073 &  x1079 &  x1085 &  x1091 &  x1094 &  x1109 &  x1115 &  x1124 & ~x12 & ~x51 & ~x246 & ~x282 & ~x285 & ~x360 & ~x402 & ~x480 & ~x597 & ~x636 & ~x783 & ~x825 & ~x861 & ~x867 & ~x903 & ~x942 & ~x1104;
assign c6184 =  x23 &  x35 &  x41 &  x47 &  x50 &  x53 &  x68 &  x71 &  x83 &  x86 &  x89 &  x104 &  x110 &  x116 &  x119 &  x122 &  x128 &  x131 &  x146 &  x152 &  x170 &  x176 &  x182 &  x197 &  x200 &  x218 &  x221 &  x230 &  x233 &  x236 &  x251 &  x260 &  x269 &  x272 &  x275 &  x278 &  x284 &  x293 &  x302 &  x314 &  x323 &  x329 &  x335 &  x338 &  x341 &  x344 &  x350 &  x359 &  x371 &  x377 &  x386 &  x389 &  x398 &  x428 &  x434 &  x443 &  x449 &  x452 &  x461 &  x482 &  x485 &  x494 &  x497 &  x515 &  x518 &  x524 &  x527 &  x542 &  x551 &  x563 &  x587 &  x590 &  x593 &  x596 &  x602 &  x614 &  x620 &  x623 &  x626 &  x632 &  x638 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x698 &  x701 &  x707 &  x713 &  x725 &  x728 &  x734 &  x746 &  x755 &  x758 &  x761 &  x773 &  x776 &  x779 &  x782 &  x791 &  x794 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x845 &  x857 &  x860 &  x866 &  x881 &  x893 &  x896 &  x917 &  x923 &  x929 &  x938 &  x941 &  x968 &  x974 &  x977 &  x992 &  x1010 &  x1034 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1079 &  x1085 &  x1094 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 & ~x3 & ~x9 & ~x84 & ~x129 & ~x246 & ~x249 & ~x252 & ~x285 & ~x366 & ~x939;
assign c6186 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x343 &  x344 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x382 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x421 &  x422 &  x425 &  x428 &  x431 &  x437 &  x440 &  x443 &  x446 &  x452 &  x455 &  x458 &  x460 &  x461 &  x464 &  x470 &  x473 &  x479 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x616 &  x620 &  x623 &  x626 &  x629 &  x635 &  x638 &  x641 &  x644 &  x646 &  x647 &  x650 &  x653 &  x655 &  x656 &  x662 &  x671 &  x674 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x890 &  x893 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x552 & ~x555 & ~x591 & ~x627 & ~x666 & ~x753 & ~x792;
assign c6188 =  x2 &  x5 &  x8 &  x14 &  x20 &  x23 &  x29 &  x32 &  x38 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x64 &  x65 &  x71 &  x74 &  x83 &  x86 &  x89 &  x92 &  x101 &  x103 &  x104 &  x107 &  x119 &  x122 &  x128 &  x131 &  x134 &  x142 &  x143 &  x152 &  x155 &  x167 &  x173 &  x179 &  x182 &  x185 &  x188 &  x194 &  x203 &  x209 &  x215 &  x224 &  x227 &  x236 &  x239 &  x245 &  x248 &  x254 &  x257 &  x259 &  x260 &  x269 &  x272 &  x275 &  x278 &  x281 &  x287 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x326 &  x329 &  x332 &  x335 &  x337 &  x344 &  x350 &  x353 &  x356 &  x362 &  x365 &  x368 &  x371 &  x380 &  x389 &  x392 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x415 &  x419 &  x425 &  x428 &  x431 &  x434 &  x440 &  x443 &  x449 &  x454 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x485 &  x494 &  x497 &  x503 &  x506 &  x509 &  x512 &  x515 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x554 &  x557 &  x563 &  x572 &  x587 &  x590 &  x596 &  x602 &  x605 &  x610 &  x617 &  x623 &  x629 &  x632 &  x638 &  x641 &  x647 &  x650 &  x662 &  x665 &  x668 &  x677 &  x683 &  x686 &  x689 &  x698 &  x701 &  x707 &  x710 &  x716 &  x719 &  x746 &  x755 &  x761 &  x764 &  x767 &  x776 &  x782 &  x788 &  x791 &  x794 &  x803 &  x809 &  x812 &  x815 &  x818 &  x830 &  x833 &  x836 &  x842 &  x851 &  x854 &  x860 &  x863 &  x872 &  x884 &  x890 &  x893 &  x899 &  x905 &  x911 &  x914 &  x917 &  x922 &  x926 &  x929 &  x941 &  x947 &  x953 &  x956 &  x959 &  x961 &  x962 &  x965 &  x971 &  x977 &  x980 &  x983 &  x989 &  x992 &  x998 &  x1000 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1038 &  x1039 &  x1043 &  x1049 &  x1055 &  x1073 &  x1076 &  x1078 &  x1079 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1117 &  x1118 &  x1121 &  x1127 &  x1130 & ~x117 & ~x897;
assign c6190 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x181 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x220 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x259 &  x260 &  x263 &  x265 &  x266 &  x269 &  x271 &  x272 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x298 &  x299 &  x302 &  x310 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x337 &  x338 &  x341 &  x344 &  x347 &  x349 &  x350 &  x353 &  x359 &  x362 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x386 &  x388 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x427 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x466 &  x467 &  x470 &  x473 &  x479 &  x482 &  x485 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x958 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1090 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x561 & ~x600 & ~x639 & ~x678 & ~x717;
assign c6192 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x44 &  x53 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x83 &  x89 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x128 &  x131 &  x134 &  x137 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x179 &  x182 &  x185 &  x191 &  x197 &  x200 &  x203 &  x209 &  x212 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x281 &  x284 &  x290 &  x299 &  x302 &  x314 &  x317 &  x323 &  x326 &  x329 &  x332 &  x338 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x407 &  x413 &  x416 &  x425 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x455 &  x458 &  x461 &  x470 &  x473 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x548 &  x551 &  x554 &  x560 &  x563 &  x569 &  x572 &  x578 &  x581 &  x584 &  x590 &  x596 &  x599 &  x602 &  x605 &  x611 &  x620 &  x623 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x659 &  x662 &  x668 &  x671 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x707 &  x710 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x776 &  x784 &  x788 &  x791 &  x797 &  x800 &  x803 &  x809 &  x812 &  x815 &  x818 &  x821 &  x823 &  x824 &  x827 &  x836 &  x839 &  x845 &  x848 &  x851 &  x857 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x920 &  x926 &  x929 &  x935 &  x940 &  x941 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x979 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1010 &  x1013 &  x1018 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1049 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x237 & ~x276 & ~x282 & ~x321 & ~x360 & ~x399 & ~x444 & ~x522 & ~x675 & ~x714 & ~x753 & ~x948 & ~x1026;
assign c6194 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x115 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x154 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x181 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x553 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x799 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x838 &  x839 &  x842 &  x845 &  x848 &  x850 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x877 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x916 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x994 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1033 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x210 & ~x288 & ~x780 & ~x819 & ~x858 & ~x897 & ~x936 & ~x975 & ~x1014 & ~x1053;
assign c6196 =  x2 &  x5 &  x8 &  x14 &  x17 &  x26 &  x29 &  x35 &  x38 &  x41 &  x44 &  x47 &  x56 &  x68 &  x74 &  x77 &  x80 &  x89 &  x101 &  x112 &  x119 &  x143 &  x152 &  x167 &  x170 &  x176 &  x179 &  x191 &  x200 &  x203 &  x209 &  x212 &  x224 &  x229 &  x239 &  x245 &  x254 &  x268 &  x269 &  x281 &  x284 &  x290 &  x296 &  x302 &  x305 &  x308 &  x320 &  x329 &  x335 &  x340 &  x344 &  x350 &  x353 &  x362 &  x368 &  x373 &  x377 &  x383 &  x386 &  x392 &  x395 &  x398 &  x407 &  x410 &  x412 &  x413 &  x425 &  x434 &  x446 &  x449 &  x458 &  x464 &  x470 &  x476 &  x479 &  x482 &  x488 &  x491 &  x500 &  x503 &  x506 &  x521 &  x524 &  x533 &  x535 &  x563 &  x572 &  x584 &  x590 &  x596 &  x599 &  x605 &  x608 &  x620 &  x631 &  x638 &  x641 &  x644 &  x670 &  x671 &  x680 &  x683 &  x692 &  x698 &  x701 &  x704 &  x707 &  x713 &  x716 &  x734 &  x740 &  x746 &  x752 &  x755 &  x761 &  x770 &  x773 &  x776 &  x782 &  x785 &  x790 &  x791 &  x794 &  x797 &  x800 &  x802 &  x824 &  x836 &  x839 &  x842 &  x854 &  x857 &  x866 &  x872 &  x875 &  x878 &  x881 &  x884 &  x886 &  x893 &  x896 &  x899 &  x902 &  x911 &  x920 &  x929 &  x935 &  x938 &  x941 &  x944 &  x950 &  x958 &  x959 &  x971 &  x974 &  x977 &  x980 &  x989 &  x995 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1040 &  x1061 &  x1067 &  x1070 &  x1085 &  x1094 &  x1115 &  x1124 &  x1127 &  x1130 & ~x354 & ~x393 & ~x549;
assign c6198 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x54 & ~x93 & ~x132 & ~x144 & ~x168 & ~x171 & ~x183 & ~x207 & ~x210 & ~x222 & ~x246 & ~x249 & ~x285 & ~x286 & ~x288 & ~x324 & ~x363 & ~x546 & ~x585 & ~x594 & ~x618;
assign c6200 =  x17 &  x26 &  x35 &  x38 &  x40 &  x47 &  x53 &  x56 &  x59 &  x65 &  x74 &  x80 &  x98 &  x101 &  x104 &  x110 &  x119 &  x125 &  x134 &  x140 &  x146 &  x155 &  x167 &  x170 &  x173 &  x178 &  x179 &  x182 &  x194 &  x197 &  x200 &  x205 &  x209 &  x212 &  x217 &  x218 &  x223 &  x230 &  x233 &  x239 &  x248 &  x284 &  x287 &  x305 &  x308 &  x311 &  x341 &  x344 &  x350 &  x359 &  x362 &  x368 &  x395 &  x410 &  x416 &  x419 &  x434 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x457 &  x458 &  x464 &  x476 &  x479 &  x506 &  x509 &  x515 &  x518 &  x530 &  x551 &  x557 &  x566 &  x575 &  x593 &  x602 &  x608 &  x611 &  x623 &  x626 &  x629 &  x644 &  x671 &  x674 &  x677 &  x680 &  x683 &  x689 &  x695 &  x704 &  x724 &  x737 &  x749 &  x764 &  x767 &  x770 &  x773 &  x785 &  x788 &  x791 &  x800 &  x803 &  x812 &  x818 &  x827 &  x830 &  x839 &  x842 &  x845 &  x848 &  x851 &  x860 &  x863 &  x881 &  x890 &  x911 &  x932 &  x935 &  x941 &  x950 &  x962 &  x974 &  x983 &  x986 &  x995 &  x1001 &  x1004 &  x1007 &  x1034 &  x1052 &  x1076 &  x1079 &  x1082 &  x1091 &  x1106 &  x1121 &  x1127 & ~x75 & ~x588 & ~x627 & ~x666 & ~x705 & ~x1032;
assign c6202 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x41 &  x44 &  x47 &  x59 &  x62 &  x65 &  x68 &  x77 &  x80 &  x83 &  x92 &  x95 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x152 &  x155 &  x158 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x236 &  x242 &  x244 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x283 &  x284 &  x287 &  x290 &  x296 &  x299 &  x305 &  x308 &  x311 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x341 &  x344 &  x347 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x386 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x415 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x439 &  x440 &  x446 &  x451 &  x455 &  x458 &  x460 &  x461 &  x473 &  x478 &  x479 &  x482 &  x485 &  x488 &  x489 &  x491 &  x494 &  x497 &  x500 &  x509 &  x512 &  x515 &  x524 &  x529 &  x530 &  x533 &  x539 &  x542 &  x545 &  x554 &  x557 &  x563 &  x566 &  x568 &  x569 &  x572 &  x575 &  x578 &  x581 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x614 &  x617 &  x620 &  x635 &  x638 &  x641 &  x644 &  x647 &  x653 &  x659 &  x662 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x688 &  x689 &  x692 &  x695 &  x698 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x727 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x752 &  x755 &  x758 &  x764 &  x766 &  x767 &  x770 &  x773 &  x776 &  x779 &  x785 &  x788 &  x791 &  x794 &  x803 &  x805 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x881 &  x884 &  x887 &  x890 &  x896 &  x902 &  x908 &  x911 &  x917 &  x920 &  x926 &  x929 &  x932 &  x938 &  x941 &  x944 &  x950 &  x953 &  x959 &  x968 &  x971 &  x974 &  x977 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x705 & ~x744;
assign c6204 =  x8 &  x14 &  x17 &  x20 &  x23 &  x32 &  x38 &  x41 &  x49 &  x56 &  x59 &  x68 &  x74 &  x80 &  x86 &  x92 &  x95 &  x98 &  x101 &  x107 &  x110 &  x119 &  x125 &  x131 &  x137 &  x139 &  x155 &  x161 &  x164 &  x167 &  x170 &  x173 &  x179 &  x184 &  x188 &  x190 &  x206 &  x209 &  x212 &  x215 &  x217 &  x224 &  x227 &  x229 &  x230 &  x233 &  x239 &  x245 &  x248 &  x257 &  x260 &  x262 &  x263 &  x269 &  x272 &  x278 &  x284 &  x293 &  x295 &  x299 &  x308 &  x320 &  x329 &  x334 &  x338 &  x341 &  x347 &  x350 &  x359 &  x367 &  x368 &  x371 &  x380 &  x383 &  x386 &  x397 &  x401 &  x404 &  x413 &  x427 &  x431 &  x436 &  x440 &  x443 &  x446 &  x455 &  x458 &  x466 &  x476 &  x482 &  x490 &  x494 &  x503 &  x505 &  x524 &  x527 &  x530 &  x545 &  x551 &  x560 &  x566 &  x569 &  x572 &  x575 &  x584 &  x587 &  x593 &  x596 &  x602 &  x608 &  x611 &  x614 &  x617 &  x629 &  x632 &  x644 &  x653 &  x656 &  x659 &  x662 &  x674 &  x677 &  x680 &  x686 &  x689 &  x692 &  x707 &  x710 &  x713 &  x725 &  x728 &  x734 &  x743 &  x749 &  x752 &  x758 &  x764 &  x767 &  x770 &  x773 &  x782 &  x785 &  x788 &  x794 &  x797 &  x800 &  x802 &  x803 &  x818 &  x833 &  x839 &  x841 &  x842 &  x848 &  x854 &  x860 &  x869 &  x875 &  x880 &  x881 &  x884 &  x899 &  x905 &  x908 &  x911 &  x917 &  x919 &  x926 &  x932 &  x935 &  x941 &  x944 &  x947 &  x953 &  x956 &  x958 &  x962 &  x980 &  x995 &  x1001 &  x1007 &  x1013 &  x1028 &  x1031 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1064 &  x1070 &  x1079 &  x1082 &  x1085 &  x1097 &  x1100 &  x1103 &  x1109 &  x1118 &  x1121 &  x1127 & ~x354 & ~x393;
assign c6206 =  x5 &  x11 &  x14 &  x23 &  x26 &  x32 &  x35 &  x38 &  x44 &  x47 &  x50 &  x53 &  x59 &  x68 &  x77 &  x80 &  x83 &  x86 &  x89 &  x95 &  x98 &  x101 &  x116 &  x122 &  x128 &  x134 &  x137 &  x149 &  x152 &  x158 &  x161 &  x170 &  x176 &  x179 &  x194 &  x206 &  x209 &  x215 &  x218 &  x221 &  x227 &  x230 &  x233 &  x242 &  x245 &  x248 &  x251 &  x254 &  x260 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x314 &  x317 &  x326 &  x329 &  x332 &  x335 &  x338 &  x344 &  x350 &  x359 &  x365 &  x368 &  x374 &  x377 &  x383 &  x389 &  x392 &  x395 &  x398 &  x416 &  x425 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x455 &  x461 &  x464 &  x470 &  x476 &  x485 &  x488 &  x494 &  x500 &  x503 &  x509 &  x515 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x542 &  x545 &  x548 &  x551 &  x557 &  x560 &  x563 &  x566 &  x569 &  x578 &  x584 &  x587 &  x590 &  x596 &  x599 &  x602 &  x605 &  x617 &  x620 &  x629 &  x635 &  x641 &  x644 &  x650 &  x653 &  x656 &  x665 &  x671 &  x674 &  x680 &  x695 &  x698 &  x701 &  x704 &  x728 &  x737 &  x740 &  x752 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x800 &  x806 &  x812 &  x815 &  x818 &  x824 &  x827 &  x830 &  x833 &  x842 &  x848 &  x854 &  x863 &  x866 &  x869 &  x875 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x908 &  x911 &  x914 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x941 &  x944 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x995 &  x1004 &  x1010 &  x1019 &  x1022 &  x1028 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1061 &  x1067 &  x1070 &  x1076 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x273 & ~x312 & ~x321 & ~x351 & ~x444 & ~x474 & ~x483 & ~x484 & ~x513 & ~x523 & ~x561 & ~x600 & ~x603 & ~x639;
assign c6208 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x29 &  x32 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x71 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x137 &  x140 &  x152 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x182 &  x188 &  x191 &  x197 &  x200 &  x203 &  x206 &  x212 &  x215 &  x218 &  x221 &  x230 &  x233 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x260 &  x263 &  x272 &  x278 &  x281 &  x284 &  x287 &  x290 &  x296 &  x302 &  x308 &  x317 &  x320 &  x326 &  x335 &  x338 &  x344 &  x347 &  x350 &  x353 &  x362 &  x365 &  x371 &  x374 &  x380 &  x383 &  x386 &  x389 &  x392 &  x398 &  x404 &  x407 &  x410 &  x419 &  x422 &  x431 &  x437 &  x440 &  x443 &  x446 &  x449 &  x454 &  x455 &  x461 &  x464 &  x467 &  x470 &  x476 &  x479 &  x482 &  x488 &  x491 &  x494 &  x506 &  x509 &  x512 &  x515 &  x518 &  x524 &  x533 &  x536 &  x539 &  x542 &  x545 &  x554 &  x557 &  x560 &  x563 &  x566 &  x578 &  x581 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x617 &  x620 &  x623 &  x626 &  x629 &  x641 &  x647 &  x650 &  x653 &  x656 &  x659 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x695 &  x698 &  x701 &  x713 &  x716 &  x722 &  x725 &  x728 &  x734 &  x737 &  x743 &  x746 &  x752 &  x755 &  x758 &  x764 &  x767 &  x770 &  x773 &  x779 &  x782 &  x785 &  x788 &  x791 &  x800 &  x806 &  x812 &  x814 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x842 &  x848 &  x853 &  x854 &  x860 &  x863 &  x869 &  x878 &  x881 &  x884 &  x887 &  x890 &  x896 &  x902 &  x905 &  x908 &  x923 &  x929 &  x935 &  x938 &  x940 &  x944 &  x947 &  x953 &  x956 &  x959 &  x962 &  x965 &  x971 &  x977 &  x980 &  x989 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1022 &  x1034 &  x1037 &  x1043 &  x1046 &  x1052 &  x1055 &  x1070 &  x1073 &  x1076 &  x1082 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 & ~x390 & ~x399 & ~x438 & ~x516 & ~x555 & ~x678 & ~x717 & ~x1020;
assign c6210 =  x5 &  x11 &  x14 &  x26 &  x29 &  x32 &  x35 &  x44 &  x50 &  x56 &  x62 &  x65 &  x68 &  x80 &  x83 &  x89 &  x95 &  x101 &  x104 &  x110 &  x113 &  x119 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x146 &  x155 &  x158 &  x164 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x200 &  x206 &  x224 &  x230 &  x236 &  x245 &  x248 &  x254 &  x257 &  x263 &  x266 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x299 &  x305 &  x308 &  x311 &  x314 &  x317 &  x323 &  x335 &  x338 &  x341 &  x344 &  x350 &  x353 &  x359 &  x362 &  x365 &  x368 &  x371 &  x377 &  x380 &  x386 &  x389 &  x392 &  x395 &  x398 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x440 &  x443 &  x455 &  x461 &  x473 &  x479 &  x482 &  x485 &  x488 &  x497 &  x503 &  x506 &  x512 &  x518 &  x521 &  x524 &  x533 &  x542 &  x545 &  x551 &  x557 &  x560 &  x566 &  x572 &  x575 &  x578 &  x581 &  x587 &  x593 &  x599 &  x608 &  x614 &  x620 &  x638 &  x641 &  x650 &  x653 &  x656 &  x662 &  x674 &  x680 &  x689 &  x692 &  x695 &  x698 &  x701 &  x707 &  x710 &  x713 &  x716 &  x719 &  x725 &  x728 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x761 &  x764 &  x767 &  x773 &  x776 &  x782 &  x788 &  x791 &  x794 &  x800 &  x806 &  x812 &  x830 &  x836 &  x842 &  x845 &  x854 &  x857 &  x866 &  x875 &  x881 &  x884 &  x893 &  x896 &  x899 &  x902 &  x923 &  x929 &  x938 &  x944 &  x947 &  x950 &  x956 &  x959 &  x962 &  x974 &  x977 &  x980 &  x986 &  x989 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1037 &  x1043 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1082 &  x1091 &  x1097 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1130 & ~x93 & ~x132 & ~x210 & ~x249 & ~x327 & ~x366 & ~x516 & ~x594 & ~x624 & ~x627 & ~x633 & ~x651 & ~x663 & ~x664 & ~x666 & ~x690 & ~x702 & ~x729 & ~x780 & ~x781;
assign c6212 =  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x95 &  x98 &  x101 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x131 &  x134 &  x137 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x203 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x263 &  x275 &  x281 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x353 &  x356 &  x359 &  x365 &  x368 &  x371 &  x374 &  x377 &  x383 &  x392 &  x395 &  x398 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x434 &  x437 &  x443 &  x446 &  x449 &  x455 &  x458 &  x461 &  x470 &  x473 &  x476 &  x479 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x509 &  x515 &  x521 &  x524 &  x527 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x569 &  x572 &  x575 &  x578 &  x587 &  x590 &  x593 &  x596 &  x605 &  x608 &  x611 &  x614 &  x620 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x674 &  x677 &  x683 &  x688 &  x689 &  x692 &  x695 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x725 &  x728 &  x734 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x767 &  x776 &  x782 &  x785 &  x788 &  x791 &  x794 &  x800 &  x803 &  x806 &  x809 &  x812 &  x821 &  x824 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x980 &  x983 &  x986 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1022 &  x1025 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1067 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x6 & ~x90 & ~x123 & ~x168 & ~x207 & ~x513 & ~x663 & ~x702 & ~x741 & ~x825 & ~x864 & ~x870 & ~x981 & ~x1020;
assign c6214 =  x2 &  x5 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x142 &  x143 &  x146 &  x149 &  x152 &  x154 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x181 &  x182 &  x185 &  x188 &  x191 &  x193 &  x194 &  x197 &  x200 &  x203 &  x206 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x232 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x263 &  x269 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x298 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x337 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x542 &  x545 &  x548 &  x551 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x856 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x895 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x934 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x962 &  x965 &  x968 &  x971 &  x973 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1012 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1051 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x441 & ~x444 & ~x483 & ~x522 & ~x561;
assign c6216 =  x2 &  x5 &  x11 &  x14 &  x17 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x53 &  x59 &  x65 &  x68 &  x71 &  x74 &  x77 &  x83 &  x86 &  x95 &  x104 &  x110 &  x113 &  x122 &  x128 &  x140 &  x149 &  x152 &  x155 &  x158 &  x176 &  x179 &  x182 &  x185 &  x191 &  x197 &  x206 &  x209 &  x215 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x248 &  x251 &  x260 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x302 &  x304 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x337 &  x338 &  x356 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x383 &  x386 &  x388 &  x392 &  x395 &  x398 &  x401 &  x407 &  x415 &  x419 &  x422 &  x427 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x452 &  x454 &  x455 &  x458 &  x464 &  x467 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x527 &  x530 &  x533 &  x535 &  x542 &  x545 &  x554 &  x557 &  x560 &  x569 &  x572 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x635 &  x638 &  x641 &  x650 &  x656 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x770 &  x776 &  x779 &  x782 &  x785 &  x791 &  x797 &  x800 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x827 &  x833 &  x836 &  x842 &  x845 &  x848 &  x851 &  x854 &  x860 &  x863 &  x866 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x953 &  x959 &  x965 &  x968 &  x974 &  x980 &  x983 &  x989 &  x992 &  x995 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1028 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1055 &  x1058 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x0 & ~x39 & ~x156 & ~x195 & ~x234 & ~x312 & ~x351 & ~x678 & ~x717 & ~x753 & ~x756 & ~x795 & ~x831;
assign c6218 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x26 &  x35 &  x41 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x197 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x236 &  x245 &  x248 &  x251 &  x254 &  x257 &  x263 &  x266 &  x269 &  x272 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x394 &  x398 &  x401 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x476 &  x479 &  x482 &  x485 &  x488 &  x494 &  x497 &  x500 &  x503 &  x506 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x551 &  x553 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x584 &  x587 &  x590 &  x596 &  x599 &  x602 &  x605 &  x608 &  x614 &  x617 &  x620 &  x623 &  x629 &  x632 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x842 &  x845 &  x848 &  x851 &  x854 &  x856 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x878 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x910 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x928 &  x929 &  x932 &  x938 &  x941 &  x947 &  x950 &  x956 &  x959 &  x962 &  x968 &  x971 &  x973 &  x974 &  x977 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1012 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1051 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1090 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x441 & ~x588 & ~x627 & ~x666 & ~x705 & ~x744 & ~x783 & ~x789 & ~x822 & ~x861 & ~x900 & ~x939 & ~x978;
assign c6220 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x76 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x895 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x934 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x973 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1049 &  x1051 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x285 & ~x288 & ~x327 & ~x366 & ~x405 & ~x438 & ~x477 & ~x516 & ~x555 & ~x594 & ~x633 & ~x672 & ~x984;
assign c6222 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x22 &  x23 &  x26 &  x29 &  x32 &  x34 &  x35 &  x38 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x61 &  x62 &  x65 &  x71 &  x73 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x112 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x139 &  x140 &  x143 &  x151 &  x152 &  x155 &  x158 &  x164 &  x167 &  x170 &  x176 &  x178 &  x179 &  x182 &  x185 &  x188 &  x190 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x229 &  x230 &  x236 &  x239 &  x242 &  x245 &  x248 &  x254 &  x257 &  x260 &  x266 &  x268 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x307 &  x308 &  x311 &  x314 &  x317 &  x320 &  x326 &  x329 &  x335 &  x338 &  x341 &  x344 &  x346 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x532 &  x533 &  x539 &  x542 &  x545 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x571 &  x572 &  x575 &  x578 &  x580 &  x581 &  x584 &  x587 &  x590 &  x593 &  x599 &  x602 &  x605 &  x608 &  x610 &  x611 &  x614 &  x617 &  x619 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x656 &  x658 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x697 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x721 &  x722 &  x725 &  x728 &  x733 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x760 &  x761 &  x764 &  x766 &  x767 &  x769 &  x770 &  x772 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x805 &  x806 &  x809 &  x811 &  x812 &  x815 &  x817 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x856 &  x857 &  x863 &  x866 &  x869 &  x872 &  x875 &  x881 &  x884 &  x887 &  x890 &  x893 &  x895 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x934 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130;
assign c6224 =  x8 &  x11 &  x17 &  x23 &  x32 &  x35 &  x38 &  x44 &  x47 &  x62 &  x65 &  x68 &  x71 &  x77 &  x83 &  x86 &  x89 &  x92 &  x95 &  x104 &  x107 &  x110 &  x116 &  x122 &  x125 &  x131 &  x140 &  x142 &  x143 &  x149 &  x152 &  x158 &  x167 &  x173 &  x181 &  x191 &  x194 &  x203 &  x206 &  x209 &  x212 &  x218 &  x224 &  x227 &  x230 &  x233 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x263 &  x269 &  x272 &  x278 &  x281 &  x284 &  x299 &  x302 &  x305 &  x311 &  x314 &  x320 &  x326 &  x329 &  x332 &  x335 &  x344 &  x353 &  x356 &  x365 &  x368 &  x374 &  x377 &  x386 &  x389 &  x395 &  x398 &  x401 &  x407 &  x410 &  x416 &  x431 &  x434 &  x440 &  x443 &  x446 &  x461 &  x464 &  x467 &  x473 &  x476 &  x485 &  x491 &  x494 &  x497 &  x500 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x532 &  x533 &  x536 &  x539 &  x542 &  x551 &  x554 &  x560 &  x566 &  x571 &  x572 &  x575 &  x581 &  x584 &  x587 &  x590 &  x596 &  x599 &  x602 &  x605 &  x608 &  x610 &  x611 &  x614 &  x617 &  x623 &  x626 &  x629 &  x632 &  x635 &  x647 &  x650 &  x656 &  x659 &  x665 &  x671 &  x674 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x701 &  x704 &  x707 &  x713 &  x716 &  x722 &  x728 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x773 &  x776 &  x779 &  x782 &  x788 &  x791 &  x803 &  x806 &  x809 &  x824 &  x826 &  x827 &  x833 &  x842 &  x845 &  x851 &  x865 &  x866 &  x869 &  x872 &  x875 &  x881 &  x884 &  x896 &  x902 &  x904 &  x905 &  x914 &  x917 &  x923 &  x926 &  x932 &  x938 &  x944 &  x947 &  x950 &  x953 &  x955 &  x956 &  x959 &  x962 &  x965 &  x971 &  x974 &  x977 &  x980 &  x983 &  x989 &  x994 &  x995 &  x998 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1085 &  x1094 &  x1097 &  x1100 &  x1103 &  x1115 &  x1117 &  x1118 &  x1121 &  x1127 &  x1130 & ~x210 & ~x249 & ~x327 & ~x405 & ~x444 & ~x858 & ~x1053;
assign c6226 =  x2 &  x5 &  x11 &  x14 &  x17 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x272 &  x275 &  x278 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x304 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x479 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x544 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x583 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x695 &  x701 &  x704 &  x707 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x740 &  x743 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x778 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x195 & ~x234 & ~x243 & ~x636 & ~x675 & ~x936 & ~x969 & ~x975;
assign c6228 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x250 &  x251 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x377 &  x380 &  x382 &  x383 &  x386 &  x388 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x653 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x790 &  x791 &  x794 &  x797 &  x803 &  x806 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x893 &  x896 &  x899 &  x905 &  x908 &  x911 &  x914 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x953 &  x956 &  x962 &  x965 &  x968 &  x974 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1007 &  x1010 &  x1018 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1124 &  x1127 &  x1130 & ~x198 & ~x237 & ~x600 & ~x636 & ~x675;
assign c6230 =  x1 &  x2 &  x8 &  x11 &  x14 &  x20 &  x22 &  x23 &  x26 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x61 &  x62 &  x65 &  x67 &  x68 &  x71 &  x74 &  x77 &  x79 &  x80 &  x83 &  x89 &  x95 &  x98 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x139 &  x145 &  x146 &  x149 &  x151 &  x152 &  x155 &  x158 &  x161 &  x164 &  x170 &  x173 &  x176 &  x178 &  x179 &  x182 &  x184 &  x185 &  x188 &  x190 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x223 &  x224 &  x227 &  x230 &  x233 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x262 &  x263 &  x266 &  x268 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x305 &  x308 &  x314 &  x320 &  x323 &  x329 &  x332 &  x335 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x365 &  x371 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x458 &  x461 &  x464 &  x467 &  x473 &  x476 &  x479 &  x485 &  x488 &  x494 &  x497 &  x500 &  x503 &  x515 &  x518 &  x521 &  x524 &  x530 &  x533 &  x536 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x584 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x680 &  x683 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x731 &  x734 &  x737 &  x740 &  x743 &  x749 &  x755 &  x758 &  x761 &  x763 &  x764 &  x767 &  x769 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x797 &  x805 &  x806 &  x809 &  x812 &  x814 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x853 &  x854 &  x860 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x886 &  x887 &  x890 &  x892 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x920 &  x923 &  x925 &  x926 &  x929 &  x932 &  x941 &  x944 &  x947 &  x950 &  x953 &  x959 &  x962 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1034 &  x1037 &  x1043 &  x1049 &  x1052 &  x1055 &  x1058 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x246 & ~x285 & ~x324 & ~x363 & ~x441 & ~x1032;
assign c6232 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x137 &  x143 &  x146 &  x149 &  x152 &  x154 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x235 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x275 &  x277 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x316 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x355 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x605 &  x608 &  x611 &  x617 &  x620 &  x623 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x916 &  x917 &  x920 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x994 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1033 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x207 & ~x246 & ~x285 & ~x288 & ~x324 & ~x325 & ~x327 & ~x363 & ~x366 & ~x405 & ~x444 & ~x585 & ~x588 & ~x858 & ~x897 & ~x936;
assign c6234 =  x2 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x116 &  x122 &  x128 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x179 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x275 &  x278 &  x281 &  x284 &  x290 &  x293 &  x299 &  x305 &  x308 &  x311 &  x314 &  x323 &  x326 &  x332 &  x335 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x368 &  x374 &  x377 &  x383 &  x386 &  x392 &  x395 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x427 &  x434 &  x437 &  x440 &  x443 &  x446 &  x452 &  x455 &  x461 &  x464 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x494 &  x497 &  x500 &  x503 &  x506 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x584 &  x586 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x641 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x671 &  x674 &  x677 &  x680 &  x689 &  x695 &  x701 &  x704 &  x707 &  x710 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x872 &  x875 &  x878 &  x884 &  x890 &  x893 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x926 &  x929 &  x932 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x959 &  x965 &  x968 &  x971 &  x974 &  x977 &  x979 &  x980 &  x983 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x195 & ~x273 & ~x282 & ~x321 & ~x351 & ~x354 & ~x360 & ~x390 & ~x522;
assign c6236 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x337 &  x338 &  x341 &  x347 &  x349 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x376 &  x377 &  x380 &  x383 &  x386 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x415 &  x416 &  x419 &  x422 &  x425 &  x427 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x454 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x527 &  x530 &  x536 &  x539 &  x542 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x665 &  x671 &  x674 &  x680 &  x683 &  x689 &  x692 &  x698 &  x701 &  x704 &  x706 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x806 &  x809 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x117 & ~x675 & ~x891 & ~x930 & ~x969 & ~x984;
assign c6238 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x379 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x418 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x457 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x806 &  x809 &  x815 &  x818 &  x824 &  x827 &  x833 &  x836 &  x839 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x926 &  x929 &  x932 &  x935 &  x937 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x976 &  x977 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1018 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x273 & ~x312 & ~x351 & ~x600 & ~x678 & ~x717 & ~x756 & ~x948 & ~x987 & ~x999 & ~x1026;
assign c6240 =  x2 &  x5 &  x8 &  x14 &  x17 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x163 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x202 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x265 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x299 &  x302 &  x304 &  x305 &  x308 &  x311 &  x314 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x337 &  x338 &  x341 &  x343 &  x344 &  x347 &  x349 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x382 &  x383 &  x386 &  x388 &  x389 &  x392 &  x395 &  x398 &  x401 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x427 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x466 &  x467 &  x470 &  x473 &  x479 &  x482 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x542 &  x545 &  x548 &  x554 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x941 &  x944 &  x950 &  x953 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x195 & ~x234 & ~x276 & ~x312 & ~x639 & ~x678 & ~x717 & ~x756 & ~x795 & ~x831 & ~x834 & ~x990;
assign c6242 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x47 &  x50 &  x56 &  x62 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x113 &  x116 &  x119 &  x122 &  x128 &  x131 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x197 &  x200 &  x203 &  x206 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x257 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x290 &  x296 &  x302 &  x305 &  x308 &  x311 &  x314 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x359 &  x362 &  x365 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x431 &  x434 &  x440 &  x446 &  x449 &  x452 &  x455 &  x461 &  x467 &  x473 &  x476 &  x479 &  x482 &  x488 &  x491 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x647 &  x650 &  x653 &  x659 &  x661 &  x662 &  x665 &  x668 &  x674 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x700 &  x701 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x770 &  x773 &  x776 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x809 &  x812 &  x815 &  x818 &  x821 &  x827 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x863 &  x866 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x950 &  x953 &  x956 &  x959 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x315 & ~x354 & ~x360 & ~x399 & ~x432 & ~x714 & ~x753 & ~x786 & ~x792 & ~x870 & ~x903 & ~x909 & ~x948 & ~x981 & ~x987 & ~x1026 & ~x1044;
assign c6244 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x649 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x384 & ~x663 & ~x669 & ~x708 & ~x747 & ~x786 & ~x825 & ~x927 & ~x942 & ~x1026;
assign c6246 =  x2 &  x11 &  x17 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x61 &  x62 &  x68 &  x77 &  x83 &  x92 &  x98 &  x101 &  x112 &  x116 &  x119 &  x125 &  x134 &  x139 &  x140 &  x143 &  x146 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x178 &  x185 &  x194 &  x197 &  x200 &  x209 &  x217 &  x224 &  x230 &  x233 &  x236 &  x239 &  x242 &  x248 &  x251 &  x256 &  x260 &  x268 &  x269 &  x272 &  x281 &  x295 &  x307 &  x308 &  x311 &  x323 &  x326 &  x329 &  x335 &  x344 &  x365 &  x368 &  x374 &  x377 &  x380 &  x383 &  x395 &  x401 &  x410 &  x413 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x440 &  x449 &  x452 &  x455 &  x461 &  x464 &  x470 &  x476 &  x479 &  x482 &  x485 &  x488 &  x500 &  x503 &  x512 &  x515 &  x521 &  x527 &  x530 &  x532 &  x535 &  x539 &  x542 &  x545 &  x548 &  x563 &  x569 &  x574 &  x587 &  x596 &  x599 &  x605 &  x610 &  x611 &  x614 &  x620 &  x629 &  x632 &  x638 &  x644 &  x649 &  x653 &  x668 &  x674 &  x677 &  x680 &  x683 &  x688 &  x689 &  x695 &  x698 &  x707 &  x719 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x755 &  x758 &  x761 &  x767 &  x776 &  x779 &  x782 &  x785 &  x788 &  x794 &  x797 &  x800 &  x818 &  x824 &  x827 &  x833 &  x836 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x863 &  x869 &  x887 &  x892 &  x896 &  x899 &  x902 &  x905 &  x911 &  x917 &  x923 &  x926 &  x932 &  x938 &  x941 &  x944 &  x950 &  x953 &  x956 &  x958 &  x959 &  x962 &  x968 &  x971 &  x977 &  x980 &  x983 &  x992 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1028 &  x1031 &  x1037 &  x1040 &  x1061 &  x1064 &  x1076 &  x1085 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 & ~x432 & ~x471 & ~x510 & ~x549 & ~x870 & ~x1059 & ~x1098;
assign c6248 =  x2 &  x5 &  x20 &  x23 &  x26 &  x32 &  x35 &  x41 &  x44 &  x59 &  x62 &  x68 &  x80 &  x86 &  x98 &  x101 &  x107 &  x116 &  x119 &  x122 &  x125 &  x134 &  x140 &  x142 &  x143 &  x149 &  x152 &  x155 &  x158 &  x164 &  x170 &  x173 &  x182 &  x191 &  x194 &  x200 &  x209 &  x212 &  x215 &  x218 &  x224 &  x233 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x263 &  x269 &  x272 &  x275 &  x281 &  x284 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x317 &  x323 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x383 &  x386 &  x389 &  x395 &  x401 &  x416 &  x422 &  x428 &  x431 &  x434 &  x440 &  x443 &  x449 &  x455 &  x458 &  x461 &  x466 &  x467 &  x470 &  x473 &  x476 &  x482 &  x485 &  x491 &  x494 &  x500 &  x503 &  x505 &  x506 &  x509 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x538 &  x539 &  x542 &  x545 &  x551 &  x557 &  x563 &  x569 &  x572 &  x575 &  x578 &  x584 &  x590 &  x593 &  x596 &  x599 &  x608 &  x622 &  x623 &  x626 &  x635 &  x638 &  x641 &  x647 &  x656 &  x671 &  x674 &  x677 &  x689 &  x692 &  x695 &  x701 &  x704 &  x707 &  x710 &  x716 &  x725 &  x731 &  x734 &  x737 &  x758 &  x761 &  x764 &  x767 &  x770 &  x776 &  x791 &  x794 &  x800 &  x803 &  x806 &  x809 &  x815 &  x821 &  x824 &  x830 &  x833 &  x848 &  x857 &  x862 &  x863 &  x878 &  x890 &  x893 &  x896 &  x901 &  x902 &  x905 &  x911 &  x917 &  x920 &  x923 &  x926 &  x940 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x968 &  x971 &  x980 &  x986 &  x989 &  x998 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1043 &  x1049 &  x1052 &  x1058 &  x1064 &  x1067 &  x1070 &  x1076 &  x1082 &  x1088 &  x1093 &  x1097 &  x1100 &  x1103 &  x1106 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130 & ~x117 & ~x312 & ~x393 & ~x429 & ~x792 & ~x831 & ~x834 & ~x873 & ~x876;
assign c6250 =  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x25 &  x29 &  x32 &  x41 &  x47 &  x65 &  x74 &  x77 &  x83 &  x86 &  x89 &  x95 &  x98 &  x101 &  x119 &  x122 &  x128 &  x131 &  x134 &  x140 &  x142 &  x143 &  x146 &  x149 &  x152 &  x158 &  x173 &  x181 &  x182 &  x185 &  x194 &  x203 &  x209 &  x212 &  x218 &  x224 &  x226 &  x230 &  x233 &  x236 &  x239 &  x245 &  x254 &  x257 &  x259 &  x263 &  x265 &  x266 &  x275 &  x278 &  x281 &  x287 &  x302 &  x308 &  x332 &  x335 &  x337 &  x347 &  x350 &  x353 &  x356 &  x359 &  x365 &  x368 &  x371 &  x376 &  x380 &  x395 &  x398 &  x404 &  x407 &  x413 &  x422 &  x431 &  x434 &  x443 &  x452 &  x455 &  x461 &  x467 &  x479 &  x491 &  x494 &  x500 &  x506 &  x509 &  x512 &  x515 &  x518 &  x524 &  x527 &  x545 &  x551 &  x557 &  x560 &  x566 &  x569 &  x572 &  x575 &  x581 &  x593 &  x596 &  x602 &  x608 &  x614 &  x617 &  x623 &  x635 &  x647 &  x662 &  x667 &  x668 &  x674 &  x677 &  x689 &  x695 &  x704 &  x710 &  x712 &  x713 &  x719 &  x734 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x763 &  x770 &  x776 &  x779 &  x782 &  x791 &  x797 &  x806 &  x815 &  x830 &  x836 &  x842 &  x851 &  x860 &  x866 &  x875 &  x878 &  x884 &  x887 &  x896 &  x899 &  x902 &  x908 &  x911 &  x914 &  x920 &  x923 &  x926 &  x935 &  x941 &  x959 &  x962 &  x965 &  x974 &  x980 &  x989 &  x998 &  x1000 &  x1001 &  x1004 &  x1007 &  x1028 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1070 &  x1073 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1112 &  x1115 &  x1118 &  x1121 & ~x897;
assign c6252 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x35 &  x38 &  x50 &  x53 &  x56 &  x62 &  x65 &  x71 &  x77 &  x89 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x119 &  x122 &  x125 &  x128 &  x140 &  x146 &  x155 &  x164 &  x173 &  x179 &  x188 &  x191 &  x194 &  x197 &  x206 &  x209 &  x212 &  x224 &  x227 &  x230 &  x239 &  x245 &  x248 &  x254 &  x257 &  x260 &  x269 &  x272 &  x275 &  x281 &  x287 &  x296 &  x302 &  x308 &  x314 &  x317 &  x320 &  x323 &  x326 &  x332 &  x335 &  x344 &  x347 &  x350 &  x353 &  x356 &  x362 &  x368 &  x377 &  x383 &  x392 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x437 &  x440 &  x443 &  x446 &  x452 &  x455 &  x461 &  x464 &  x470 &  x479 &  x482 &  x485 &  x491 &  x494 &  x497 &  x503 &  x506 &  x509 &  x512 &  x533 &  x542 &  x545 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x587 &  x590 &  x602 &  x605 &  x608 &  x611 &  x620 &  x623 &  x629 &  x632 &  x635 &  x644 &  x656 &  x668 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x698 &  x701 &  x704 &  x707 &  x710 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x737 &  x743 &  x746 &  x749 &  x761 &  x764 &  x776 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x836 &  x842 &  x854 &  x860 &  x863 &  x872 &  x878 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x911 &  x914 &  x920 &  x922 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x953 &  x956 &  x961 &  x965 &  x967 &  x968 &  x971 &  x974 &  x977 &  x980 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1010 &  x1022 &  x1034 &  x1039 &  x1043 &  x1046 &  x1049 &  x1055 &  x1058 &  x1061 &  x1064 &  x1073 &  x1079 &  x1082 &  x1085 &  x1094 &  x1100 &  x1103 &  x1106 &  x1121 &  x1127 &  x1130 & ~x93 & ~x94 & ~x172 & ~x210 & ~x213 & ~x249 & ~x366 & ~x702 & ~x741 & ~x780 & ~x783 & ~x819 & ~x897 & ~x936 & ~x975 & ~x1014 & ~x1053;
assign c6254 =  x5 &  x8 &  x14 &  x17 &  x26 &  x32 &  x35 &  x38 &  x44 &  x47 &  x50 &  x53 &  x56 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x116 &  x122 &  x131 &  x134 &  x140 &  x143 &  x146 &  x149 &  x155 &  x158 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x362 &  x371 &  x374 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x428 &  x431 &  x434 &  x437 &  x440 &  x446 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x560 &  x563 &  x566 &  x569 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x605 &  x608 &  x611 &  x617 &  x620 &  x623 &  x629 &  x632 &  x635 &  x641 &  x644 &  x647 &  x653 &  x656 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x704 &  x710 &  x713 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x863 &  x866 &  x869 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x905 &  x908 &  x914 &  x920 &  x923 &  x926 &  x929 &  x932 &  x938 &  x941 &  x947 &  x953 &  x956 &  x959 &  x965 &  x968 &  x974 &  x980 &  x983 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1130 & ~x48 & ~x159 & ~x198 & ~x204 & ~x321 & ~x360 & ~x480 & ~x558 & ~x597 & ~x642 & ~x675 & ~x693 & ~x714 & ~x720 & ~x732 & ~x759 & ~x831 & ~x870 & ~x1005;
assign c6256 =  x2 &  x5 &  x8 &  x11 &  x17 &  x20 &  x23 &  x29 &  x32 &  x35 &  x38 &  x41 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x71 &  x76 &  x83 &  x86 &  x89 &  x92 &  x101 &  x110 &  x113 &  x119 &  x122 &  x125 &  x134 &  x143 &  x146 &  x155 &  x158 &  x161 &  x167 &  x173 &  x176 &  x179 &  x182 &  x188 &  x191 &  x197 &  x200 &  x203 &  x209 &  x212 &  x218 &  x224 &  x227 &  x230 &  x239 &  x242 &  x248 &  x257 &  x260 &  x263 &  x275 &  x284 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x317 &  x320 &  x323 &  x326 &  x332 &  x341 &  x344 &  x347 &  x350 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x413 &  x416 &  x422 &  x428 &  x431 &  x437 &  x443 &  x446 &  x449 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x485 &  x488 &  x491 &  x493 &  x494 &  x500 &  x503 &  x506 &  x509 &  x515 &  x521 &  x524 &  x527 &  x530 &  x532 &  x533 &  x548 &  x551 &  x557 &  x566 &  x572 &  x575 &  x578 &  x581 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x611 &  x614 &  x629 &  x632 &  x635 &  x638 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x665 &  x668 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x704 &  x707 &  x710 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x805 &  x806 &  x812 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x844 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x869 &  x872 &  x875 &  x878 &  x883 &  x887 &  x890 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x921 &  x922 &  x923 &  x926 &  x929 &  x932 &  x941 &  x947 &  x950 &  x953 &  x956 &  x961 &  x962 &  x965 &  x968 &  x974 &  x977 &  x980 &  x989 &  x992 &  x998 &  x1000 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x171 & ~x210 & ~x249 & ~x288 & ~x327 & ~x462;
assign c6258 =  x2 &  x5 &  x8 &  x11 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x41 &  x44 &  x47 &  x50 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x940 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1018 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x237 & ~x276 & ~x405 & ~x522 & ~x558 & ~x597 & ~x675 & ~x714 & ~x753 & ~x831 & ~x870 & ~x942 & ~x1005 & ~x1026;
assign c6260 =  x2 &  x5 &  x8 &  x11 &  x20 &  x23 &  x29 &  x35 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x71 &  x74 &  x80 &  x86 &  x89 &  x98 &  x101 &  x110 &  x113 &  x115 &  x116 &  x119 &  x131 &  x134 &  x140 &  x143 &  x146 &  x149 &  x152 &  x154 &  x155 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x194 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x233 &  x236 &  x239 &  x248 &  x251 &  x260 &  x269 &  x272 &  x278 &  x281 &  x287 &  x296 &  x314 &  x317 &  x320 &  x341 &  x344 &  x347 &  x355 &  x356 &  x365 &  x371 &  x374 &  x377 &  x395 &  x398 &  x407 &  x413 &  x416 &  x422 &  x431 &  x434 &  x440 &  x446 &  x455 &  x464 &  x467 &  x473 &  x476 &  x485 &  x491 &  x497 &  x506 &  x515 &  x524 &  x527 &  x530 &  x533 &  x536 &  x542 &  x548 &  x551 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x587 &  x593 &  x599 &  x602 &  x605 &  x611 &  x614 &  x617 &  x623 &  x629 &  x635 &  x638 &  x644 &  x650 &  x662 &  x665 &  x674 &  x677 &  x680 &  x683 &  x695 &  x704 &  x707 &  x710 &  x713 &  x716 &  x725 &  x728 &  x734 &  x740 &  x746 &  x749 &  x752 &  x761 &  x767 &  x770 &  x773 &  x779 &  x782 &  x785 &  x788 &  x794 &  x797 &  x806 &  x809 &  x811 &  x827 &  x833 &  x850 &  x851 &  x857 &  x863 &  x866 &  x872 &  x877 &  x878 &  x889 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x914 &  x923 &  x926 &  x932 &  x938 &  x944 &  x953 &  x956 &  x959 &  x962 &  x965 &  x967 &  x971 &  x974 &  x980 &  x983 &  x986 &  x992 &  x994 &  x995 &  x998 &  x1001 &  x1006 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1031 &  x1033 &  x1034 &  x1037 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1066 &  x1070 &  x1073 &  x1079 &  x1084 &  x1085 &  x1088 &  x1091 &  x1106 &  x1112 &  x1115 &  x1121 &  x1127 & ~x249 & ~x288 & ~x327 & ~x405 & ~x444 & ~x483 & ~x897 & ~x936 & ~x975 & ~x1014;
assign c6262 =  x2 &  x8 &  x11 &  x14 &  x17 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x113 &  x116 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x185 &  x188 &  x200 &  x203 &  x206 &  x212 &  x215 &  x218 &  x221 &  x224 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x302 &  x305 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x335 &  x341 &  x344 &  x347 &  x353 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x458 &  x461 &  x467 &  x470 &  x473 &  x476 &  x482 &  x488 &  x491 &  x497 &  x503 &  x506 &  x509 &  x515 &  x521 &  x527 &  x530 &  x536 &  x539 &  x542 &  x545 &  x548 &  x550 &  x551 &  x554 &  x557 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x686 &  x689 &  x692 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x761 &  x764 &  x770 &  x776 &  x779 &  x782 &  x788 &  x791 &  x794 &  x797 &  x800 &  x806 &  x809 &  x818 &  x821 &  x827 &  x830 &  x836 &  x839 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x878 &  x884 &  x887 &  x890 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1016 &  x1019 &  x1022 &  x1025 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 & ~x99 & ~x105 & ~x138 & ~x435 & ~x519 & ~x558 & ~x597 & ~x636 & ~x729 & ~x822;
assign c6264 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x542 &  x548 &  x551 &  x554 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x809 &  x812 &  x815 &  x818 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x159 & ~x165 & ~x195 & ~x249 & ~x288 & ~x327 & ~x405 & ~x444 & ~x484 & ~x522 & ~x523 & ~x780 & ~x819 & ~x1023;
assign c6266 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x22 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x61 &  x65 &  x68 &  x74 &  x77 &  x79 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x128 &  x131 &  x134 &  x137 &  x139 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x178 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x217 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x256 &  x257 &  x263 &  x266 &  x269 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x295 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x334 &  x335 &  x338 &  x341 &  x347 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x398 &  x401 &  x407 &  x410 &  x412 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x449 &  x451 &  x452 &  x455 &  x458 &  x461 &  x464 &  x470 &  x473 &  x476 &  x479 &  x482 &  x488 &  x490 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x524 &  x529 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x560 &  x563 &  x566 &  x568 &  x569 &  x572 &  x575 &  x578 &  x580 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x607 &  x608 &  x611 &  x614 &  x617 &  x619 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x644 &  x646 &  x650 &  x653 &  x656 &  x658 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x685 &  x686 &  x688 &  x689 &  x692 &  x695 &  x697 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x724 &  x725 &  x728 &  x731 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x758 &  x760 &  x763 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x788 &  x791 &  x794 &  x797 &  x802 &  x803 &  x806 &  x809 &  x812 &  x814 &  x815 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x841 &  x842 &  x845 &  x848 &  x851 &  x853 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x892 &  x896 &  x899 &  x902 &  x905 &  x911 &  x914 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x441 & ~x480 & ~x519;
assign c6268 =  x2 &  x5 &  x11 &  x14 &  x17 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x320 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x355 &  x356 &  x359 &  x362 &  x368 &  x371 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x394 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x452 &  x455 &  x461 &  x464 &  x467 &  x473 &  x476 &  x479 &  x482 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x662 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x698 &  x701 &  x707 &  x710 &  x713 &  x716 &  x719 &  x721 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x752 &  x755 &  x760 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x797 &  x799 &  x806 &  x809 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x838 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1127 &  x1130 & ~x9 & ~x171 & ~x342 & ~x363 & ~x405 & ~x408 & ~x663 & ~x672 & ~x702 & ~x741;
assign c6270 =  x2 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x281 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x419 &  x422 &  x425 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x653 &  x656 &  x659 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x719 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x838 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x955 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x994 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x0 & ~x9 & ~x39 & ~x78 & ~x132 & ~x171 & ~x366 & ~x405 & ~x406 & ~x444 & ~x445 & ~x483 & ~x522 & ~x663 & ~x702 & ~x819 & ~x858 & ~x936 & ~x975 & ~x1053;
assign c6272 =  x2 &  x5 &  x17 &  x20 &  x23 &  x32 &  x35 &  x38 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x80 &  x83 &  x86 &  x95 &  x98 &  x101 &  x107 &  x110 &  x113 &  x116 &  x122 &  x125 &  x128 &  x131 &  x134 &  x140 &  x142 &  x143 &  x146 &  x152 &  x158 &  x164 &  x170 &  x173 &  x176 &  x182 &  x185 &  x194 &  x197 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x230 &  x233 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x278 &  x284 &  x287 &  x290 &  x298 &  x299 &  x305 &  x308 &  x310 &  x311 &  x320 &  x326 &  x329 &  x337 &  x338 &  x344 &  x350 &  x353 &  x356 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x379 &  x389 &  x392 &  x395 &  x398 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x434 &  x440 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x473 &  x476 &  x482 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x548 &  x551 &  x554 &  x557 &  x560 &  x566 &  x572 &  x578 &  x581 &  x584 &  x587 &  x593 &  x596 &  x599 &  x602 &  x611 &  x614 &  x623 &  x629 &  x632 &  x635 &  x638 &  x647 &  x650 &  x656 &  x665 &  x668 &  x674 &  x677 &  x680 &  x686 &  x701 &  x710 &  x713 &  x716 &  x719 &  x725 &  x728 &  x731 &  x740 &  x743 &  x746 &  x749 &  x751 &  x752 &  x755 &  x758 &  x767 &  x770 &  x776 &  x779 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x851 &  x857 &  x866 &  x869 &  x872 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x926 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x971 &  x974 &  x977 &  x980 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1028 &  x1034 &  x1040 &  x1043 &  x1049 &  x1055 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 & ~x195 & ~x600 & ~x714 & ~x831 & ~x870;
assign c6274 =  x2 &  x11 &  x14 &  x38 &  x50 &  x59 &  x71 &  x80 &  x89 &  x116 &  x131 &  x134 &  x140 &  x143 &  x152 &  x164 &  x185 &  x191 &  x200 &  x206 &  x239 &  x254 &  x260 &  x275 &  x281 &  x287 &  x293 &  x299 &  x302 &  x314 &  x326 &  x338 &  x341 &  x377 &  x386 &  x407 &  x416 &  x431 &  x440 &  x446 &  x452 &  x464 &  x476 &  x482 &  x485 &  x491 &  x500 &  x512 &  x545 &  x548 &  x554 &  x557 &  x608 &  x620 &  x632 &  x635 &  x644 &  x668 &  x671 &  x683 &  x695 &  x701 &  x704 &  x728 &  x734 &  x773 &  x788 &  x800 &  x809 &  x827 &  x830 &  x857 &  x859 &  x860 &  x863 &  x875 &  x893 &  x899 &  x905 &  x920 &  x923 &  x940 &  x956 &  x968 &  x971 &  x976 &  x979 &  x1001 &  x1013 &  x1016 &  x1018 &  x1019 &  x1034 &  x1057 &  x1067 &  x1082 &  x1091 &  x1094 &  x1096 &  x1103 &  x1118 &  x1121 &  x1130 & ~x135 & ~x438 & ~x471 & ~x510 & ~x630 & ~x864 & ~x870 & ~x888 & ~x909;
assign c6276 =  x2 &  x5 &  x20 &  x23 &  x25 &  x26 &  x29 &  x32 &  x35 &  x50 &  x59 &  x62 &  x68 &  x83 &  x86 &  x95 &  x98 &  x101 &  x103 &  x110 &  x128 &  x134 &  x140 &  x155 &  x158 &  x161 &  x164 &  x170 &  x176 &  x181 &  x187 &  x188 &  x191 &  x194 &  x206 &  x209 &  x215 &  x226 &  x227 &  x248 &  x265 &  x275 &  x281 &  x287 &  x293 &  x296 &  x302 &  x320 &  x326 &  x332 &  x347 &  x350 &  x356 &  x359 &  x362 &  x374 &  x377 &  x383 &  x389 &  x395 &  x401 &  x407 &  x415 &  x419 &  x421 &  x425 &  x427 &  x437 &  x440 &  x443 &  x446 &  x454 &  x455 &  x464 &  x466 &  x467 &  x476 &  x482 &  x488 &  x500 &  x527 &  x530 &  x533 &  x544 &  x545 &  x560 &  x563 &  x566 &  x575 &  x581 &  x582 &  x584 &  x590 &  x593 &  x599 &  x605 &  x608 &  x611 &  x617 &  x622 &  x623 &  x626 &  x629 &  x638 &  x650 &  x653 &  x662 &  x674 &  x680 &  x683 &  x698 &  x704 &  x710 &  x719 &  x734 &  x737 &  x740 &  x749 &  x755 &  x761 &  x764 &  x773 &  x776 &  x785 &  x788 &  x791 &  x818 &  x827 &  x836 &  x842 &  x845 &  x848 &  x857 &  x860 &  x863 &  x866 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x893 &  x899 &  x905 &  x908 &  x911 &  x914 &  x929 &  x935 &  x938 &  x941 &  x950 &  x953 &  x956 &  x967 &  x983 &  x986 &  x992 &  x1001 &  x1019 &  x1022 &  x1025 &  x1031 &  x1040 &  x1046 &  x1055 &  x1061 &  x1079 &  x1082 &  x1088 &  x1094 &  x1100 &  x1103 &  x1118 &  x1124 &  x1130;
assign c6278 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x56 &  x59 &  x62 &  x65 &  x71 &  x77 &  x80 &  x83 &  x89 &  x95 &  x98 &  x101 &  x104 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x163 &  x167 &  x173 &  x176 &  x179 &  x182 &  x185 &  x191 &  x194 &  x197 &  x200 &  x206 &  x209 &  x212 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x241 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x266 &  x269 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x299 &  x302 &  x304 &  x305 &  x308 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x337 &  x338 &  x341 &  x343 &  x344 &  x347 &  x349 &  x350 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x382 &  x383 &  x386 &  x388 &  x389 &  x392 &  x395 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x421 &  x422 &  x425 &  x427 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x455 &  x458 &  x460 &  x461 &  x464 &  x467 &  x473 &  x476 &  x479 &  x482 &  x485 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x554 &  x557 &  x560 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x734 &  x737 &  x740 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x851 &  x857 &  x863 &  x866 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x911 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x974 &  x977 &  x979 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1057 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1127 &  x1130 & ~x195 & ~x273 & ~x312 & ~x351 & ~x522 & ~x678 & ~x714 & ~x717 & ~x756;
assign c6280 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x119 &  x122 &  x125 &  x131 &  x134 &  x143 &  x146 &  x149 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x206 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x689 &  x692 &  x695 &  x698 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x6 & ~x12 & ~x51 & ~x84 & ~x90 & ~x123 & ~x129 & ~x168 & ~x201 & ~x207 & ~x240 & ~x279 & ~x285 & ~x324 & ~x363 & ~x396 & ~x402 & ~x435 & ~x441 & ~x480 & ~x519 & ~x558 & ~x597 & ~x630 & ~x636 & ~x669 & ~x675 & ~x714 & ~x753 & ~x792 & ~x825 & ~x831 & ~x864 & ~x870 & ~x903 & ~x942 & ~x948 & ~x981 & ~x1011 & ~x1098;
assign c6282 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x275 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x234 & ~x321 & ~x441 & ~x444 & ~x483 & ~x522 & ~x600 & ~x639 & ~x678 & ~x741 & ~x780 & ~x819 & ~x858 & ~x897 & ~x906 & ~x936 & ~x945 & ~x975 & ~x1053;
assign c6284 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x82 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x121 &  x122 &  x125 &  x128 &  x131 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x160 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x260 &  x263 &  x272 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x344 &  x347 &  x350 &  x353 &  x356 &  x362 &  x365 &  x368 &  x371 &  x374 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x440 &  x443 &  x449 &  x452 &  x454 &  x455 &  x458 &  x461 &  x464 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x491 &  x494 &  x500 &  x503 &  x506 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x557 &  x560 &  x563 &  x566 &  x568 &  x569 &  x572 &  x575 &  x581 &  x584 &  x590 &  x593 &  x595 &  x596 &  x599 &  x602 &  x605 &  x608 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x634 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x655 &  x656 &  x659 &  x662 &  x665 &  x668 &  x673 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x707 &  x713 &  x716 &  x719 &  x722 &  x728 &  x731 &  x737 &  x740 &  x746 &  x752 &  x755 &  x758 &  x761 &  x764 &  x770 &  x773 &  x776 &  x779 &  x782 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x881 &  x884 &  x887 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x956 &  x962 &  x965 &  x968 &  x971 &  x974 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x345 & ~x366;
assign c6286 =  x5 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x68 &  x71 &  x74 &  x77 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x122 &  x125 &  x128 &  x131 &  x134 &  x140 &  x143 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x188 &  x194 &  x197 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x233 &  x239 &  x245 &  x248 &  x251 &  x254 &  x260 &  x263 &  x269 &  x278 &  x281 &  x283 &  x284 &  x287 &  x290 &  x299 &  x305 &  x308 &  x311 &  x317 &  x322 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x449 &  x452 &  x454 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x509 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x532 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x571 &  x575 &  x578 &  x581 &  x584 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x610 &  x613 &  x614 &  x617 &  x620 &  x626 &  x629 &  x632 &  x635 &  x641 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x671 &  x674 &  x680 &  x683 &  x685 &  x686 &  x692 &  x695 &  x698 &  x704 &  x707 &  x710 &  x719 &  x722 &  x723 &  x725 &  x727 &  x731 &  x743 &  x746 &  x749 &  x752 &  x758 &  x761 &  x763 &  x764 &  x767 &  x773 &  x776 &  x779 &  x782 &  x791 &  x794 &  x797 &  x800 &  x802 &  x803 &  x805 &  x806 &  x809 &  x812 &  x818 &  x824 &  x829 &  x833 &  x836 &  x841 &  x842 &  x848 &  x851 &  x854 &  x857 &  x863 &  x866 &  x869 &  x872 &  x881 &  x883 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x908 &  x917 &  x920 &  x923 &  x929 &  x932 &  x938 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x977 &  x980 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130;
assign c6288 =  x8 &  x20 &  x26 &  x29 &  x32 &  x38 &  x44 &  x47 &  x50 &  x53 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x98 &  x104 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x137 &  x140 &  x149 &  x152 &  x155 &  x158 &  x173 &  x176 &  x179 &  x182 &  x197 &  x203 &  x206 &  x209 &  x215 &  x224 &  x227 &  x230 &  x238 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x263 &  x266 &  x269 &  x272 &  x277 &  x278 &  x284 &  x287 &  x290 &  x293 &  x299 &  x308 &  x311 &  x314 &  x320 &  x329 &  x338 &  x344 &  x350 &  x356 &  x362 &  x374 &  x383 &  x392 &  x395 &  x404 &  x407 &  x410 &  x416 &  x419 &  x428 &  x440 &  x443 &  x446 &  x455 &  x458 &  x461 &  x467 &  x479 &  x485 &  x488 &  x494 &  x500 &  x509 &  x512 &  x515 &  x524 &  x530 &  x539 &  x545 &  x548 &  x554 &  x560 &  x563 &  x566 &  x569 &  x571 &  x578 &  x581 &  x590 &  x593 &  x596 &  x599 &  x602 &  x610 &  x614 &  x617 &  x620 &  x623 &  x629 &  x647 &  x649 &  x653 &  x662 &  x665 &  x671 &  x674 &  x676 &  x683 &  x689 &  x692 &  x698 &  x701 &  x704 &  x709 &  x713 &  x727 &  x728 &  x731 &  x737 &  x740 &  x746 &  x755 &  x757 &  x761 &  x764 &  x767 &  x770 &  x776 &  x779 &  x782 &  x793 &  x794 &  x803 &  x806 &  x815 &  x818 &  x821 &  x824 &  x830 &  x832 &  x839 &  x842 &  x848 &  x851 &  x857 &  x860 &  x863 &  x866 &  x869 &  x875 &  x878 &  x883 &  x884 &  x890 &  x893 &  x896 &  x905 &  x911 &  x920 &  x923 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x949 &  x950 &  x953 &  x956 &  x959 &  x968 &  x971 &  x974 &  x977 &  x983 &  x988 &  x989 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1046 &  x1052 &  x1061 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1103 &  x1109 &  x1112 &  x1115 &  x1127 & ~x132 & ~x510 & ~x549 & ~x585 & ~x588 & ~x663 & ~x705 & ~x741 & ~x744 & ~x858 & ~x861 & ~x897 & ~x936 & ~x975;
assign c6290 =  x11 &  x32 &  x59 &  x71 &  x83 &  x86 &  x92 &  x113 &  x122 &  x131 &  x134 &  x179 &  x209 &  x215 &  x227 &  x230 &  x233 &  x239 &  x248 &  x275 &  x287 &  x293 &  x308 &  x314 &  x332 &  x335 &  x355 &  x356 &  x386 &  x389 &  x407 &  x410 &  x428 &  x434 &  x458 &  x467 &  x485 &  x491 &  x503 &  x509 &  x542 &  x545 &  x560 &  x572 &  x578 &  x581 &  x593 &  x599 &  x620 &  x632 &  x644 &  x647 &  x656 &  x659 &  x671 &  x680 &  x698 &  x746 &  x749 &  x752 &  x755 &  x761 &  x764 &  x799 &  x800 &  x803 &  x806 &  x815 &  x827 &  x838 &  x854 &  x863 &  x866 &  x875 &  x896 &  x899 &  x902 &  x916 &  x922 &  x923 &  x961 &  x974 &  x1000 &  x1016 &  x1022 &  x1039 &  x1052 &  x1079 &  x1091 &  x1118 & ~x3 & ~x93 & ~x132 & ~x249 & ~x289 & ~x327 & ~x549 & ~x588 & ~x897 & ~x1053;
assign c6292 =  x8 &  x11 &  x32 &  x59 &  x62 &  x68 &  x77 &  x80 &  x100 &  x101 &  x104 &  x113 &  x118 &  x122 &  x143 &  x146 &  x167 &  x173 &  x182 &  x184 &  x188 &  x191 &  x194 &  x197 &  x200 &  x209 &  x215 &  x223 &  x224 &  x230 &  x239 &  x245 &  x254 &  x257 &  x266 &  x269 &  x272 &  x281 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x311 &  x317 &  x320 &  x326 &  x332 &  x341 &  x350 &  x356 &  x365 &  x368 &  x371 &  x374 &  x383 &  x386 &  x389 &  x404 &  x410 &  x416 &  x428 &  x437 &  x440 &  x443 &  x455 &  x467 &  x473 &  x478 &  x491 &  x494 &  x500 &  x506 &  x509 &  x515 &  x533 &  x551 &  x554 &  x557 &  x575 &  x578 &  x587 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x632 &  x641 &  x644 &  x647 &  x656 &  x659 &  x662 &  x665 &  x686 &  x689 &  x698 &  x701 &  x707 &  x710 &  x713 &  x716 &  x725 &  x734 &  x749 &  x752 &  x758 &  x761 &  x764 &  x773 &  x779 &  x791 &  x806 &  x809 &  x812 &  x815 &  x821 &  x830 &  x833 &  x836 &  x848 &  x851 &  x857 &  x863 &  x866 &  x884 &  x893 &  x896 &  x899 &  x914 &  x923 &  x926 &  x932 &  x941 &  x944 &  x950 &  x953 &  x956 &  x959 &  x968 &  x977 &  x983 &  x986 &  x989 &  x1001 &  x1007 &  x1010 &  x1022 &  x1025 &  x1037 &  x1040 &  x1043 &  x1055 &  x1058 &  x1064 &  x1067 &  x1073 &  x1076 &  x1097 &  x1100 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 &  x1130 & ~x84 & ~x123 & ~x129 & ~x246 & ~x369 & ~x441 & ~x636 & ~x1083 & ~x1104;
assign c6294 =  x1 &  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x29 &  x35 &  x38 &  x41 &  x47 &  x53 &  x59 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x98 &  x100 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x128 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x167 &  x170 &  x173 &  x185 &  x188 &  x200 &  x206 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x260 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x338 &  x341 &  x350 &  x356 &  x365 &  x368 &  x374 &  x377 &  x383 &  x386 &  x392 &  x395 &  x398 &  x401 &  x413 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x443 &  x449 &  x452 &  x458 &  x461 &  x464 &  x470 &  x473 &  x482 &  x491 &  x493 &  x506 &  x512 &  x518 &  x521 &  x524 &  x530 &  x533 &  x539 &  x542 &  x551 &  x554 &  x560 &  x563 &  x568 &  x578 &  x581 &  x584 &  x587 &  x593 &  x599 &  x617 &  x619 &  x620 &  x626 &  x641 &  x643 &  x644 &  x650 &  x653 &  x655 &  x658 &  x659 &  x665 &  x671 &  x674 &  x677 &  x680 &  x686 &  x694 &  x695 &  x701 &  x704 &  x707 &  x710 &  x716 &  x719 &  x722 &  x728 &  x740 &  x743 &  x749 &  x752 &  x758 &  x761 &  x770 &  x773 &  x779 &  x782 &  x788 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x821 &  x824 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x854 &  x863 &  x866 &  x872 &  x875 &  x878 &  x884 &  x896 &  x899 &  x902 &  x911 &  x920 &  x926 &  x932 &  x935 &  x938 &  x941 &  x947 &  x953 &  x962 &  x965 &  x968 &  x974 &  x977 &  x989 &  x992 &  x995 &  x1001 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1067 &  x1070 &  x1076 &  x1088 &  x1094 &  x1097 &  x1115 &  x1124 &  x1127 &  x1130 & ~x84 & ~x90 & ~x207 & ~x426;
assign c6296 =  x2 &  x11 &  x14 &  x26 &  x35 &  x50 &  x53 &  x56 &  x59 &  x62 &  x77 &  x80 &  x86 &  x107 &  x122 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x164 &  x167 &  x182 &  x185 &  x188 &  x191 &  x197 &  x203 &  x212 &  x218 &  x221 &  x230 &  x232 &  x233 &  x236 &  x260 &  x263 &  x272 &  x281 &  x290 &  x329 &  x344 &  x347 &  x353 &  x359 &  x362 &  x371 &  x377 &  x389 &  x394 &  x407 &  x410 &  x413 &  x419 &  x434 &  x437 &  x440 &  x443 &  x446 &  x455 &  x461 &  x470 &  x472 &  x473 &  x476 &  x482 &  x485 &  x491 &  x497 &  x500 &  x506 &  x511 &  x518 &  x521 &  x524 &  x527 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x560 &  x572 &  x578 &  x581 &  x596 &  x602 &  x608 &  x614 &  x626 &  x629 &  x632 &  x635 &  x644 &  x653 &  x656 &  x665 &  x668 &  x671 &  x680 &  x698 &  x704 &  x707 &  x746 &  x749 &  x761 &  x773 &  x782 &  x788 &  x791 &  x799 &  x806 &  x827 &  x830 &  x836 &  x845 &  x850 &  x866 &  x875 &  x878 &  x884 &  x889 &  x893 &  x899 &  x905 &  x917 &  x920 &  x929 &  x932 &  x944 &  x950 &  x959 &  x962 &  x968 &  x977 &  x986 &  x995 &  x1000 &  x1004 &  x1007 &  x1013 &  x1019 &  x1022 &  x1028 &  x1037 &  x1040 &  x1067 &  x1076 &  x1079 &  x1091 &  x1097 &  x1115 &  x1127 &  x1130 & ~x9 & ~x366 & ~x702 & ~x741 & ~x750 & ~x897;
assign c6298 =  x5 &  x14 &  x17 &  x20 &  x29 &  x35 &  x38 &  x41 &  x44 &  x50 &  x56 &  x68 &  x74 &  x77 &  x80 &  x86 &  x89 &  x92 &  x107 &  x113 &  x118 &  x119 &  x122 &  x125 &  x137 &  x143 &  x145 &  x146 &  x151 &  x155 &  x157 &  x164 &  x170 &  x179 &  x185 &  x196 &  x200 &  x209 &  x212 &  x215 &  x221 &  x229 &  x230 &  x233 &  x236 &  x239 &  x242 &  x251 &  x266 &  x275 &  x293 &  x296 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x326 &  x335 &  x341 &  x344 &  x350 &  x356 &  x365 &  x368 &  x380 &  x383 &  x389 &  x398 &  x416 &  x422 &  x425 &  x428 &  x434 &  x437 &  x440 &  x446 &  x449 &  x458 &  x461 &  x470 &  x473 &  x482 &  x485 &  x497 &  x503 &  x506 &  x518 &  x527 &  x536 &  x539 &  x542 &  x547 &  x548 &  x551 &  x557 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x586 &  x587 &  x590 &  x593 &  x599 &  x602 &  x605 &  x617 &  x619 &  x620 &  x623 &  x625 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x659 &  x668 &  x674 &  x680 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x785 &  x794 &  x800 &  x803 &  x806 &  x812 &  x815 &  x818 &  x820 &  x824 &  x827 &  x830 &  x836 &  x839 &  x845 &  x848 &  x854 &  x860 &  x866 &  x869 &  x878 &  x884 &  x887 &  x890 &  x896 &  x898 &  x905 &  x911 &  x917 &  x926 &  x929 &  x937 &  x941 &  x950 &  x965 &  x974 &  x989 &  x991 &  x998 &  x1004 &  x1007 &  x1019 &  x1022 &  x1025 &  x1030 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1061 &  x1067 &  x1073 &  x1076 &  x1082 &  x1088 &  x1094 &  x1097 &  x1100 &  x1106 &  x1118 &  x1121 &  x1127 &  x1130 & ~x30 & ~x246 & ~x285 & ~x363 & ~x402 & ~x441 & ~x597 & ~x636 & ~x675 & ~x714 & ~x753;
assign c61 =  x549 &  x705 &  x744 & ~x1041;
assign c63 =  x1059 & ~x1000;
assign c65 =  x265 &  x601 &  x796 & ~x817;
assign c67 =  x14 &  x95 &  x188 &  x194 &  x265 &  x266 &  x601 &  x611 &  x715 &  x833 &  x863 &  x869 &  x896 &  x898 &  x1103 & ~x849 & ~x888 & ~x996;
assign c69 =  x211 &  x250 &  x282 &  x289 &  x352 &  x508;
assign c611 =  x820 & ~x610;
assign c613 =  x627 &  x666 &  x744 & ~x498 & ~x1041;
assign c615 =  x1000 & ~x142 & ~x177 & ~x202;
assign c617 =  x781 & ~x195 & ~x762;
assign c619 =  x391 &  x468 &  x586 & ~x514;
assign c621 =  x17 &  x142 &  x241 &  x272 &  x368 &  x466 &  x476 &  x505 &  x520 &  x563 &  x605 &  x650 &  x656 &  x728 &  x812 &  x836 &  x935 &  x953 & ~x624 & ~x702 & ~x780 & ~x1074;
assign c623 =  x447 &  x508 &  x520;
assign c625 =  x44 &  x148 &  x220 &  x253 &  x394 &  x472 &  x806 &  x809 & ~x51;
assign c627 = ~x869;
assign c629 =  x669 & ~x127 & ~x879;
assign c631 =  x313 &  x391 &  x469 &  x509 &  x566 &  x751 & ~x298 & ~x936;
assign c633 =  x265 &  x496 &  x640 &  x819 &  x1093 & ~x648;
assign c635 =  x157 &  x196 &  x274 &  x352 &  x391 &  x556 &  x655 &  x732 & ~x429;
assign c637 =  x481 & ~x493;
assign c639 =  x288 &  x430 &  x1048 &  x1123;
assign c641 =  x175 &  x286 &  x404 &  x559 &  x637 &  x757 & ~x1080;
assign c643 =  x63 &  x108 &  x469 &  x625;
assign c645 =  x17 &  x88 &  x313 & ~x220 & ~x279 & ~x819 & ~x1053;
assign c647 =  x196 &  x313 &  x377 &  x383 &  x857 & ~x192 & ~x298 & ~x858;
assign c649 =  x304 &  x342 &  x562 &  x601 &  x757;
assign c651 = ~x348 & ~x412;
assign c653 =  x586 &  x664 & ~x423 & ~x673;
assign c655 = ~x271 & ~x412;
assign c657 =  x37 &  x469 & ~x514;
assign c659 =  x484 &  x666 &  x744 & ~x621 & ~x924;
assign c661 =  x523 &  x742 & ~x655 & ~x837;
assign c663 =  x175 &  x742 & ~x622;
assign c665 =  x468 & ~x382;
assign c667 =  x169 &  x208 &  x233 &  x253 &  x526 &  x542 &  x603 &  x613 &  x793 &  x872;
assign c669 =  x200 &  x278 &  x313 &  x352 &  x391 &  x469 &  x1078 & ~x231 & ~x378 & ~x978;
assign c671 =  x47 &  x161 &  x435 &  x475 &  x513 &  x695 &  x908 &  x938 &  x1115 & ~x468 & ~x639 & ~x780 & ~x1029 & ~x1041;
assign c673 =  x37 &  x547 &  x625 &  x1091 & ~x117 & ~x156 & ~x426 & ~x594;
assign c675 =  x481 &  x678 & ~x726;
assign c677 =  x664 &  x666 & ~x45 & ~x673;
assign c679 =  x211 &  x352 &  x391 &  x747 &  x786 & ~x339;
assign c681 =  x117 &  x195 &  x352 &  x452 &  x650 &  x778 & ~x624 & ~x858;
assign c683 =  x351 & ~x271;
assign c685 =  x546 & ~x466;
assign c687 =  x280 &  x409 &  x445 &  x781 & ~x12 & ~x1111;
assign c689 =  x147 & ~x84 & ~x735;
assign c691 =  x742 & ~x610;
assign c693 =  x11 &  x14 &  x80 &  x98 &  x161 &  x203 &  x221 &  x239 &  x293 &  x350 &  x374 &  x398 &  x403 &  x410 &  x425 &  x494 &  x500 &  x524 &  x563 &  x569 &  x578 &  x593 &  x602 &  x653 &  x677 &  x749 &  x797 &  x830 &  x907 &  x917 &  x920 &  x932 &  x1085 &  x1100 & ~x243 & ~x840 & ~x996 & ~x1002;
assign c695 =  x208 &  x470 &  x674 & ~x529 & ~x567 & ~x609;
assign c697 =  x53 &  x71 &  x176 &  x191 &  x196 &  x233 &  x352 &  x353 &  x380 &  x391 &  x497 &  x539 &  x560 &  x599 &  x623 &  x695 &  x716 &  x770 &  x788 &  x833 &  x883 &  x929 &  x965 &  x974 &  x992 &  x1025 &  x1043 &  x1046 &  x1055 & ~x259 & ~x298 & ~x624 & ~x897;
assign c699 =  x471 &  x552;
assign c6101 =  x62 &  x80 &  x140 &  x143 &  x164 &  x176 &  x353 &  x377 &  x404 &  x446 &  x586 &  x617 &  x625 &  x629 &  x695 &  x701 &  x742 &  x761 &  x824 &  x926 &  x938 &  x1088 & ~x117 & ~x156 & ~x459 & ~x495 & ~x498;
assign c6103 =  x549 & ~x781 & ~x820;
assign c6105 =  x559 & ~x570 & ~x649;
assign c6107 =  x79 &  x94 &  x195 &  x234 &  x557 &  x803 &  x811 &  x917 &  x1013 &  x1058 &  x1088 &  x1112 & ~x180 & ~x192 & ~x258 & ~x900;
assign c6109 =  x94 &  x157 &  x203 &  x218 &  x234 &  x260 &  x287 &  x488 &  x548 &  x587 &  x680 &  x758 &  x778 &  x812 &  x821 &  x914 &  x1001 &  x1052 & ~x624 & ~x819 & ~x858;
assign c6111 =  x480 &  x549;
assign c6113 =  x230 &  x481 &  x509 &  x620 &  x641 &  x698 &  x898 &  x976 &  x1023 & ~x687;
assign c6115 =  x132 &  x967 & ~x343;
assign c6117 =  x253 &  x438 & ~x429;
assign c6119 =  x461 &  x664 &  x742 &  x820 &  x898 &  x1054 &  x1093 & ~x414 & ~x649;
assign c6121 =  x110 &  x191 &  x236 &  x304 &  x640 &  x791 &  x893 &  x897 & ~x168 & ~x237 & ~x243 & ~x276;
assign c6123 =  x358 &  x981 & ~x1030;
assign c6125 =  x859 &  x897 & ~x129 & ~x234;
assign c6127 =  x234 &  x1117 & ~x114 & ~x142 & ~x180 & ~x279;
assign c6129 =  x194 &  x251 &  x352 &  x359 &  x380 &  x527 &  x536 &  x692 &  x728 &  x827 &  x866 &  x872 &  x971 &  x989 & ~x231 & ~x262 & ~x819;
assign c6131 =  x438 &  x481 & ~x390;
assign c6133 =  x109 &  x403 & ~x727;
assign c6135 =  x187 &  x625 &  x703 &  x742 &  x820 & ~x787;
assign c6137 =  x549 &  x666 & ~x387 & ~x426 & ~x723;
assign c6139 =  x390 & ~x270 & ~x336 & ~x436;
assign c6141 =  x520 & ~x610 & ~x688;
assign c6143 =  x559 &  x637 & ~x684 & ~x687 & ~x912;
assign c6145 =  x204 & ~x337;
assign c6147 =  x897 &  x1053 & ~x883;
assign c6149 =  x897 & ~x156 & ~x777;
assign c6151 =  x227 &  x304 &  x488 &  x703 &  x781 &  x820 &  x859 &  x890 &  x1019 & ~x765 & ~x895;
assign c6153 =  x328 &  x942 & ~x243 & ~x780 & ~x1041;
assign c6155 =  x522 & ~x733;
assign c6157 =  x25 &  x313 &  x352 &  x469 &  x503 &  x547 &  x581 & ~x537 & ~x990;
assign c6159 =  x367 &  x484 &  x1024 &  x1061 &  x1101 & ~x648;
assign c6161 =  x526 &  x611 &  x637 &  x672 &  x1073 & ~x195 & ~x234;
assign c6163 =  x9 &  x195 &  x700 & ~x525;
assign c6165 =  x9 &  x195 &  x313 &  x734 & ~x180 & ~x741 & ~x819 & ~x820 & ~x1014;
assign c6167 =  x238 & ~x531 & ~x862;
assign c6169 =  x41 &  x209 &  x470 &  x479 &  x559 &  x560 &  x594 &  x598 &  x758 & ~x609;
assign c6171 = ~x426 & ~x492 & ~x529 & ~x777;
assign c6173 =  x16 &  x62 &  x78 &  x117 &  x234 &  x308 &  x623 &  x818 &  x833 &  x967 & ~x858;
assign c6175 =  x5 &  x35 &  x38 &  x86 &  x92 &  x215 &  x263 &  x275 &  x308 &  x314 &  x329 &  x332 &  x335 &  x350 &  x353 &  x362 &  x458 &  x473 &  x476 &  x481 &  x509 &  x516 &  x533 &  x563 &  x566 &  x611 &  x644 &  x674 &  x779 &  x833 &  x866 &  x878 &  x902 &  x908 &  x935 &  x1016 &  x1043 &  x1127 & ~x528;
assign c6177 =  x274 &  x549;
assign c6179 =  x209 &  x227 &  x352 &  x549 &  x569 &  x584 &  x653 &  x743 & ~x0;
assign c6181 =  x14 &  x20 &  x26 &  x29 &  x32 &  x78 &  x110 &  x140 &  x195 &  x215 &  x218 &  x245 &  x274 &  x278 &  x305 &  x308 &  x313 &  x314 &  x329 &  x365 &  x377 &  x386 &  x401 &  x416 &  x431 &  x449 &  x452 &  x467 &  x509 &  x518 &  x539 &  x578 &  x592 &  x629 &  x641 &  x674 &  x728 &  x731 &  x740 &  x839 &  x845 &  x890 &  x896 &  x905 &  x929 &  x989 &  x994 &  x1001 &  x1004 &  x1028 &  x1034 &  x1046 &  x1055 &  x1070 &  x1094 &  x1100 & ~x102 & ~x114 & ~x141 & ~x180;
assign c6183 =  x945 & ~x307;
assign c6185 =  x718 &  x781 & ~x276 & ~x777 & ~x817;
assign c6187 =  x628 &  x906 &  x943 & ~x918;
assign c6189 =  x1 &  x32 &  x40 &  x74 &  x79 &  x117 &  x134 &  x156 &  x157 &  x195 &  x196 &  x206 &  x224 &  x234 &  x274 &  x314 &  x332 &  x359 &  x443 &  x455 &  x503 &  x506 &  x542 &  x572 &  x596 &  x611 &  x641 &  x644 &  x680 &  x778 &  x845 &  x881 &  x908 &  x914 &  x929 &  x962 &  x995 &  x1013 &  x1094 & ~x141 & ~x666 & ~x897;
assign c6191 =  x104 &  x549 &  x627 &  x666 &  x725 &  x744 &  x1040 &  x1091;
assign c6193 =  x444 &  x483 &  x586;
assign c6195 =  x3 &  x209 &  x904 & ~x163 & ~x705;
assign c6197 =  x718 &  x859 & ~x778 & ~x903;
assign c6199 =  x23 &  x26 &  x53 &  x56 &  x62 &  x71 &  x74 &  x77 &  x80 &  x89 &  x92 &  x95 &  x125 &  x140 &  x158 &  x161 &  x182 &  x191 &  x224 &  x263 &  x269 &  x281 &  x290 &  x296 &  x302 &  x317 &  x353 &  x356 &  x362 &  x392 &  x394 &  x398 &  x401 &  x410 &  x416 &  x431 &  x440 &  x443 &  x446 &  x455 &  x458 &  x461 &  x464 &  x467 &  x472 &  x473 &  x476 &  x494 &  x515 &  x550 &  x551 &  x554 &  x559 &  x563 &  x589 &  x590 &  x608 &  x611 &  x620 &  x623 &  x626 &  x629 &  x632 &  x665 &  x668 &  x675 &  x683 &  x695 &  x701 &  x712 &  x715 &  x716 &  x725 &  x728 &  x743 &  x754 &  x767 &  x770 &  x788 &  x812 &  x839 &  x848 &  x851 &  x869 &  x878 &  x881 &  x884 &  x896 &  x899 &  x905 &  x926 &  x932 &  x950 &  x956 &  x971 &  x983 &  x1007 &  x1022 &  x1031 &  x1034 &  x1037 &  x1043 &  x1055 &  x1058 &  x1061 &  x1067 &  x1070 &  x1079 &  x1088 &  x1097 &  x1109 &  x1118;
assign c6201 =  x391 & ~x193 & ~x684;
assign c6203 =  x14 &  x143 &  x214 &  x253 &  x290 &  x403 &  x695 &  x710 &  x734 &  x910 & ~x624 & ~x762 & ~x1029 & ~x1068;
assign c6205 =  x32 &  x44 &  x56 &  x65 &  x89 &  x137 &  x140 &  x170 &  x188 &  x194 &  x212 &  x288 &  x289 &  x296 &  x302 &  x308 &  x311 &  x352 &  x367 &  x380 &  x386 &  x395 &  x413 &  x455 &  x485 &  x494 &  x503 &  x506 &  x509 &  x533 &  x545 &  x560 &  x566 &  x608 &  x626 &  x641 &  x656 &  x689 &  x692 &  x713 &  x737 &  x743 &  x773 &  x776 &  x794 &  x824 &  x836 &  x839 &  x893 &  x908 &  x914 &  x929 &  x950 &  x986 &  x995 &  x1016 &  x1019 &  x1064 &  x1123 & ~x576;
assign c6207 =  x110 &  x122 &  x236 &  x275 &  x305 &  x448 &  x464 &  x484 &  x596 &  x626 &  x782 &  x953 &  x1010 &  x1067 &  x1084 &  x1100 & ~x576;
assign c6209 =  x94 &  x234 &  x273 &  x430 & ~x154 & ~x1056;
assign c6211 =  x136 &  x1003 & ~x760;
assign c6213 =  x130 &  x952 & ~x862;
assign c6215 =  x304 &  x900 & ~x739;
assign c6217 =  x522 &  x625 & ~x912;
assign c6219 = ~x95;
assign c6221 =  x157 &  x471 &  x700 &  x817;
assign c6223 =  x78 & ~x63 & ~x409;
assign c6225 =  x187 &  x625 &  x780 &  x858 & ~x234;
assign c6227 =  x9 &  x156 & ~x142 & ~x858;
assign c6229 =  x265 &  x304 &  x637 &  x781 &  x820 &  x898 &  x1031 &  x1085 & ~x273 & ~x699 & ~x804;
assign c6231 =  x481 &  x594 & ~x612;
assign c6233 =  x70 &  x523 &  x586 & ~x537 & ~x873;
assign c6235 =  x167 &  x187 &  x193 &  x239 &  x319 &  x395 &  x562 &  x589 &  x716 &  x743 &  x781 &  x839 &  x899 &  x998 &  x1094 & ~x315;
assign c6237 =  x5 &  x11 &  x155 &  x167 &  x179 &  x187 &  x308 &  x374 &  x745 &  x749 &  x890 &  x1067 & ~x699 & ~x1111;
assign c6239 =  x61 &  x94 &  x409 &  x556 &  x679 &  x791 &  x897;
assign c6241 =  x939 & ~x195 & ~x958;
assign c6243 =  x158 &  x282 &  x586 &  x1007 & ~x414;
assign c6245 =  x196 &  x471 &  x771 &  x841;
assign c6247 =  x148 &  x430 &  x744;
assign c6249 =  x165 &  x313 &  x391 &  x908 & ~x192;
assign c6251 =  x196 &  x390 &  x401 &  x602 &  x746 &  x752 &  x794 &  x1082 & ~x232 & ~x357;
assign c6253 =  x52 &  x483 & ~x291;
assign c6255 = ~x379 & ~x382 & ~x681;
assign c6257 = ~x617;
assign c6259 =  x277 & ~x804 & ~x862;
assign c6261 =  x430 &  x585 &  x663 &  x963;
assign c6263 =  x664 &  x906 & ~x535;
assign c6265 =  x62 &  x98 &  x104 &  x115 &  x173 &  x209 &  x218 &  x224 &  x241 &  x242 &  x311 &  x377 &  x398 &  x467 &  x472 &  x581 &  x589 &  x590 &  x659 &  x677 &  x680 &  x701 &  x713 &  x749 &  x764 &  x770 &  x839 &  x902 &  x932 &  x947 &  x1034 & ~x51 & ~x120 & ~x717;
assign c6267 =  x364 & ~x427;
assign c6269 =  x271 &  x406 &  x664 &  x859 &  x900 & ~x354;
assign c6271 =  x25 &  x227 &  x413 &  x523 &  x547 & ~x681;
assign c6273 =  x936 & ~x661 & ~x787;
assign c6275 =  x19 &  x37 &  x484 & ~x543 & ~x567;
assign c6277 = ~x415 & ~x901;
assign c6279 =  x282 & ~x420;
assign c6281 =  x97 &  x484 &  x508 &  x617 &  x869 & ~x459 & ~x495;
assign c6283 =  x273 &  x430 & ~x154 & ~x231 & ~x1059;
assign c6285 =  x664 &  x744 & ~x661 & ~x723;
assign c6287 =  x588 & ~x490 & ~x573;
assign c6289 =  x324;
assign c6291 =  x364 &  x586 &  x625 & ~x427;
assign c6293 = ~x76 & ~x241 & ~x492;
assign c6295 =  x741 & ~x649 & ~x709;
assign c6297 =  x897 & ~x699 & ~x805;
assign c6299 =  x31 &  x70 &  x187 &  x703 & ~x51 & ~x955;
assign c70 =  x2 &  x5 &  x11 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x80 &  x83 &  x89 &  x92 &  x95 &  x98 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x170 &  x176 &  x179 &  x182 &  x185 &  x188 &  x194 &  x197 &  x203 &  x212 &  x221 &  x224 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x251 &  x254 &  x257 &  x260 &  x263 &  x272 &  x275 &  x278 &  x281 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x317 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x371 &  x374 &  x377 &  x383 &  x386 &  x391 &  x395 &  x398 &  x401 &  x407 &  x413 &  x419 &  x425 &  x431 &  x440 &  x446 &  x449 &  x455 &  x458 &  x461 &  x464 &  x470 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x506 &  x512 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x545 &  x548 &  x551 &  x560 &  x566 &  x569 &  x572 &  x578 &  x581 &  x584 &  x590 &  x593 &  x596 &  x602 &  x605 &  x608 &  x614 &  x617 &  x620 &  x623 &  x626 &  x632 &  x635 &  x638 &  x647 &  x653 &  x656 &  x659 &  x665 &  x668 &  x670 &  x671 &  x674 &  x680 &  x683 &  x692 &  x695 &  x698 &  x701 &  x709 &  x713 &  x716 &  x719 &  x725 &  x728 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x758 &  x761 &  x767 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x932 &  x935 &  x938 &  x941 &  x944 &  x950 &  x953 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x980 &  x983 &  x986 &  x989 &  x992 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1031 &  x1037 &  x1040 &  x1043 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1118 &  x1127 & ~x369 & ~x408 & ~x447 & ~x486 & ~x531 & ~x564 & ~x570 & ~x627 & ~x666 & ~x702 & ~x706 & ~x741 & ~x744 & ~x745 & ~x780 & ~x783 & ~x861 & ~x900 & ~x936 & ~x939 & ~x975 & ~x1053;
assign c72 =  x2 &  x5 &  x11 &  x14 &  x26 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x104 &  x110 &  x113 &  x116 &  x122 &  x125 &  x131 &  x140 &  x143 &  x149 &  x155 &  x158 &  x161 &  x164 &  x165 &  x167 &  x170 &  x173 &  x182 &  x185 &  x188 &  x191 &  x194 &  x196 &  x197 &  x205 &  x209 &  x212 &  x215 &  x227 &  x230 &  x233 &  x234 &  x238 &  x239 &  x248 &  x254 &  x266 &  x272 &  x273 &  x275 &  x278 &  x281 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x320 &  x323 &  x332 &  x335 &  x347 &  x350 &  x352 &  x356 &  x362 &  x365 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x391 &  x392 &  x395 &  x398 &  x404 &  x410 &  x416 &  x422 &  x425 &  x428 &  x430 &  x434 &  x455 &  x461 &  x464 &  x473 &  x485 &  x488 &  x494 &  x506 &  x509 &  x530 &  x536 &  x539 &  x545 &  x557 &  x560 &  x569 &  x572 &  x578 &  x581 &  x587 &  x590 &  x593 &  x599 &  x602 &  x605 &  x608 &  x614 &  x617 &  x620 &  x623 &  x629 &  x635 &  x641 &  x650 &  x653 &  x656 &  x659 &  x674 &  x677 &  x680 &  x689 &  x695 &  x701 &  x710 &  x713 &  x716 &  x719 &  x728 &  x734 &  x740 &  x743 &  x746 &  x752 &  x755 &  x767 &  x770 &  x776 &  x779 &  x782 &  x788 &  x791 &  x812 &  x818 &  x821 &  x827 &  x830 &  x833 &  x839 &  x848 &  x854 &  x860 &  x866 &  x875 &  x878 &  x884 &  x887 &  x890 &  x896 &  x899 &  x902 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x947 &  x956 &  x962 &  x965 &  x968 &  x974 &  x977 &  x980 &  x992 &  x1004 &  x1016 &  x1022 &  x1025 &  x1034 &  x1037 &  x1040 &  x1043 &  x1073 &  x1076 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1118 &  x1124 &  x1127 & ~x162 & ~x240 & ~x241 & ~x336 & ~x375 & ~x519 & ~x666;
assign c74 =  x2 &  x8 &  x11 &  x17 &  x20 &  x23 &  x26 &  x44 &  x47 &  x50 &  x59 &  x62 &  x68 &  x71 &  x77 &  x86 &  x89 &  x91 &  x92 &  x95 &  x101 &  x104 &  x107 &  x110 &  x116 &  x122 &  x128 &  x130 &  x131 &  x134 &  x137 &  x140 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x170 &  x173 &  x179 &  x185 &  x188 &  x194 &  x197 &  x203 &  x206 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x239 &  x242 &  x245 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x278 &  x281 &  x284 &  x287 &  x290 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x338 &  x341 &  x344 &  x350 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x380 &  x383 &  x389 &  x392 &  x395 &  x401 &  x404 &  x407 &  x413 &  x416 &  x419 &  x422 &  x428 &  x431 &  x434 &  x437 &  x443 &  x446 &  x455 &  x458 &  x464 &  x467 &  x470 &  x473 &  x476 &  x485 &  x494 &  x506 &  x509 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x547 &  x548 &  x554 &  x557 &  x560 &  x563 &  x572 &  x575 &  x578 &  x581 &  x584 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x617 &  x620 &  x623 &  x629 &  x632 &  x635 &  x644 &  x647 &  x650 &  x656 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x689 &  x692 &  x695 &  x698 &  x704 &  x707 &  x710 &  x713 &  x716 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x752 &  x755 &  x758 &  x761 &  x773 &  x776 &  x779 &  x782 &  x794 &  x797 &  x800 &  x802 &  x806 &  x809 &  x815 &  x818 &  x821 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x851 &  x854 &  x857 &  x863 &  x869 &  x872 &  x875 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x919 &  x923 &  x926 &  x929 &  x935 &  x938 &  x941 &  x944 &  x947 &  x953 &  x956 &  x959 &  x965 &  x968 &  x977 &  x980 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130 & ~x279 & ~x666 & ~x667 & ~x705 & ~x706 & ~x744 & ~x745 & ~x783 & ~x784 & ~x823 & ~x900 & ~x939;
assign c76 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x399 &  x400 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x430 &  x431 &  x437 &  x438 &  x439 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x469 &  x470 &  x473 &  x476 &  x478 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x507 &  x508 &  x509 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x547 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x625 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x662 &  x664 &  x665 &  x668 &  x671 &  x674 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x703 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x742 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x926 &  x929 &  x932 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x396 & ~x435 & ~x474 & ~x531 & ~x570 & ~x609 & ~x648 & ~x687 & ~x744 & ~x783 & ~x784 & ~x822 & ~x823 & ~x861;
assign c78 =  x17 &  x23 &  x26 &  x38 &  x44 &  x47 &  x50 &  x56 &  x65 &  x68 &  x71 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x110 &  x119 &  x128 &  x131 &  x143 &  x152 &  x155 &  x158 &  x161 &  x170 &  x176 &  x185 &  x188 &  x200 &  x203 &  x212 &  x215 &  x224 &  x227 &  x239 &  x248 &  x251 &  x260 &  x266 &  x275 &  x281 &  x305 &  x314 &  x320 &  x323 &  x326 &  x328 &  x329 &  x335 &  x338 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x377 &  x383 &  x386 &  x389 &  x398 &  x404 &  x410 &  x419 &  x425 &  x431 &  x434 &  x437 &  x443 &  x446 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x488 &  x491 &  x497 &  x509 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x542 &  x545 &  x548 &  x554 &  x557 &  x560 &  x572 &  x575 &  x578 &  x581 &  x590 &  x601 &  x602 &  x611 &  x617 &  x620 &  x635 &  x638 &  x641 &  x650 &  x656 &  x659 &  x668 &  x671 &  x677 &  x679 &  x689 &  x692 &  x695 &  x701 &  x707 &  x713 &  x716 &  x718 &  x719 &  x722 &  x724 &  x728 &  x740 &  x746 &  x752 &  x761 &  x773 &  x785 &  x788 &  x794 &  x800 &  x803 &  x806 &  x815 &  x827 &  x830 &  x833 &  x836 &  x842 &  x845 &  x848 &  x857 &  x863 &  x866 &  x872 &  x884 &  x890 &  x899 &  x911 &  x914 &  x917 &  x923 &  x926 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x956 &  x959 &  x965 &  x968 &  x971 &  x977 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1013 &  x1028 &  x1031 &  x1040 &  x1058 &  x1064 &  x1067 &  x1079 &  x1082 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1112 &  x1118 &  x1121 &  x1124 &  x1130 & ~x498 & ~x537 & ~x570 & ~x576 & ~x627 & ~x636 & ~x666 & ~x667 & ~x675 & ~x705 & ~x706 & ~x714 & ~x745 & ~x783 & ~x822;
assign c710 =  x11 &  x20 &  x26 &  x29 &  x35 &  x38 &  x41 &  x47 &  x50 &  x56 &  x65 &  x71 &  x77 &  x80 &  x83 &  x86 &  x89 &  x95 &  x101 &  x107 &  x110 &  x113 &  x119 &  x122 &  x125 &  x131 &  x134 &  x143 &  x149 &  x152 &  x155 &  x158 &  x164 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x197 &  x200 &  x203 &  x206 &  x209 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x251 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x281 &  x284 &  x286 &  x292 &  x296 &  x299 &  x302 &  x304 &  x305 &  x308 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x331 &  x332 &  x338 &  x347 &  x353 &  x356 &  x362 &  x365 &  x368 &  x370 &  x371 &  x374 &  x377 &  x380 &  x389 &  x392 &  x395 &  x398 &  x401 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x434 &  x437 &  x440 &  x442 &  x446 &  x452 &  x461 &  x464 &  x467 &  x473 &  x476 &  x479 &  x481 &  x482 &  x485 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x515 &  x520 &  x521 &  x524 &  x530 &  x533 &  x536 &  x539 &  x545 &  x548 &  x551 &  x559 &  x560 &  x563 &  x566 &  x569 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x637 &  x638 &  x644 &  x647 &  x650 &  x653 &  x662 &  x665 &  x668 &  x671 &  x677 &  x680 &  x683 &  x689 &  x695 &  x698 &  x701 &  x703 &  x704 &  x707 &  x710 &  x719 &  x722 &  x728 &  x731 &  x734 &  x742 &  x746 &  x752 &  x755 &  x758 &  x761 &  x764 &  x770 &  x773 &  x776 &  x779 &  x782 &  x791 &  x797 &  x800 &  x803 &  x812 &  x815 &  x818 &  x827 &  x833 &  x836 &  x839 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x874 &  x875 &  x881 &  x884 &  x887 &  x890 &  x896 &  x898 &  x899 &  x902 &  x908 &  x911 &  x913 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x937 &  x938 &  x941 &  x947 &  x950 &  x952 &  x953 &  x956 &  x959 &  x962 &  x965 &  x971 &  x974 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1016 &  x1019 &  x1022 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1097 &  x1106 &  x1112 &  x1115 &  x1121 & ~x978 & ~x1017;
assign c712 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x320 &  x323 &  x326 &  x329 &  x335 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x362 &  x371 &  x374 &  x380 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x473 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x503 &  x506 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x557 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x596 &  x599 &  x601 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x625 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x668 &  x674 &  x677 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x703 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x734 &  x737 &  x740 &  x742 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x781 &  x782 &  x785 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x814 &  x815 &  x818 &  x820 &  x824 &  x830 &  x833 &  x836 &  x839 &  x845 &  x848 &  x851 &  x854 &  x857 &  x859 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x892 &  x893 &  x896 &  x898 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x952 &  x953 &  x956 &  x959 &  x962 &  x968 &  x971 &  x974 &  x977 &  x983 &  x986 &  x989 &  x992 &  x995 &  x997 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x570 & ~x609 & ~x648 & ~x649 & ~x687 & ~x726 & ~x765 & ~x804 & ~x978;
assign c714 =  x2 &  x5 &  x11 &  x14 &  x20 &  x26 &  x29 &  x35 &  x38 &  x41 &  x44 &  x50 &  x59 &  x65 &  x74 &  x77 &  x80 &  x86 &  x92 &  x95 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x122 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x247 &  x248 &  x251 &  x257 &  x260 &  x263 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x286 &  x287 &  x290 &  x293 &  x296 &  x305 &  x308 &  x311 &  x314 &  x323 &  x325 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x364 &  x365 &  x374 &  x377 &  x383 &  x389 &  x392 &  x395 &  x398 &  x401 &  x403 &  x404 &  x407 &  x410 &  x413 &  x419 &  x422 &  x434 &  x437 &  x440 &  x441 &  x442 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x467 &  x473 &  x476 &  x479 &  x481 &  x482 &  x485 &  x491 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x520 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x559 &  x560 &  x566 &  x569 &  x572 &  x575 &  x578 &  x584 &  x587 &  x590 &  x596 &  x598 &  x599 &  x605 &  x608 &  x611 &  x614 &  x617 &  x626 &  x629 &  x632 &  x635 &  x644 &  x647 &  x650 &  x659 &  x662 &  x665 &  x668 &  x680 &  x686 &  x689 &  x692 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x728 &  x734 &  x737 &  x740 &  x743 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x796 &  x797 &  x803 &  x806 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x835 &  x836 &  x839 &  x842 &  x848 &  x851 &  x854 &  x857 &  x863 &  x869 &  x872 &  x875 &  x878 &  x884 &  x887 &  x890 &  x893 &  x896 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x968 &  x974 &  x980 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1124 &  x1127 & ~x195 & ~x204 & ~x273 & ~x312 & ~x351 & ~x861 & ~x900 & ~x939 & ~x978;
assign c716 =  x8 &  x11 &  x13 &  x17 &  x20 &  x26 &  x29 &  x41 &  x44 &  x50 &  x59 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x98 &  x101 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x143 &  x155 &  x158 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x188 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x218 &  x224 &  x230 &  x236 &  x239 &  x245 &  x248 &  x254 &  x257 &  x260 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x290 &  x296 &  x299 &  x305 &  x308 &  x314 &  x323 &  x332 &  x335 &  x341 &  x347 &  x350 &  x356 &  x362 &  x365 &  x368 &  x371 &  x374 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x434 &  x437 &  x440 &  x443 &  x446 &  x455 &  x461 &  x464 &  x470 &  x473 &  x482 &  x485 &  x488 &  x494 &  x497 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x530 &  x536 &  x545 &  x548 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x584 &  x590 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x644 &  x647 &  x665 &  x668 &  x671 &  x674 &  x677 &  x683 &  x686 &  x689 &  x692 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x755 &  x767 &  x773 &  x779 &  x782 &  x785 &  x788 &  x791 &  x800 &  x803 &  x806 &  x809 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x854 &  x857 &  x863 &  x866 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x905 &  x908 &  x911 &  x914 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1010 &  x1013 &  x1019 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1088 &  x1091 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1127 &  x1130 & ~x180 & ~x393 & ~x394 & ~x432 & ~x433 & ~x471 & ~x510 & ~x585 & ~x663 & ~x702 & ~x741 & ~x774 & ~x813 & ~x891;
assign c718 =  x2 &  x5 &  x17 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x47 &  x53 &  x62 &  x74 &  x77 &  x80 &  x86 &  x89 &  x98 &  x104 &  x107 &  x113 &  x116 &  x119 &  x125 &  x131 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x173 &  x179 &  x182 &  x185 &  x188 &  x194 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x226 &  x230 &  x233 &  x242 &  x245 &  x254 &  x257 &  x260 &  x263 &  x266 &  x272 &  x275 &  x278 &  x281 &  x290 &  x293 &  x296 &  x302 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x338 &  x350 &  x353 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x382 &  x383 &  x386 &  x395 &  x398 &  x401 &  x407 &  x413 &  x419 &  x421 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x446 &  x449 &  x458 &  x461 &  x467 &  x470 &  x473 &  x479 &  x485 &  x488 &  x497 &  x500 &  x506 &  x512 &  x518 &  x521 &  x524 &  x529 &  x530 &  x536 &  x539 &  x542 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x584 &  x590 &  x593 &  x598 &  x599 &  x602 &  x605 &  x608 &  x611 &  x617 &  x626 &  x638 &  x644 &  x650 &  x653 &  x656 &  x659 &  x665 &  x668 &  x671 &  x674 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x707 &  x716 &  x719 &  x734 &  x743 &  x746 &  x755 &  x758 &  x761 &  x767 &  x770 &  x779 &  x794 &  x797 &  x806 &  x809 &  x815 &  x821 &  x824 &  x827 &  x833 &  x839 &  x842 &  x848 &  x851 &  x857 &  x863 &  x866 &  x872 &  x875 &  x884 &  x887 &  x890 &  x902 &  x905 &  x914 &  x917 &  x923 &  x926 &  x938 &  x944 &  x953 &  x956 &  x959 &  x962 &  x971 &  x974 &  x977 &  x986 &  x989 &  x995 &  x1004 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1055 &  x1058 &  x1061 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1097 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x351 & ~x354 & ~x390 & ~x393 & ~x432 & ~x1018 & ~x1095;
assign c720 =  x2 &  x5 &  x11 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x44 &  x47 &  x50 &  x56 &  x59 &  x62 &  x68 &  x74 &  x83 &  x86 &  x89 &  x92 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x119 &  x122 &  x125 &  x128 &  x131 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x200 &  x206 &  x212 &  x215 &  x218 &  x221 &  x224 &  x230 &  x233 &  x239 &  x245 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x275 &  x278 &  x281 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x317 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x353 &  x356 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x395 &  x398 &  x401 &  x404 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x434 &  x437 &  x440 &  x443 &  x452 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x491 &  x494 &  x497 &  x500 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x545 &  x548 &  x551 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x584 &  x587 &  x590 &  x602 &  x605 &  x611 &  x620 &  x623 &  x626 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x656 &  x662 &  x668 &  x674 &  x680 &  x683 &  x689 &  x692 &  x698 &  x701 &  x704 &  x716 &  x719 &  x722 &  x728 &  x731 &  x737 &  x740 &  x746 &  x749 &  x752 &  x761 &  x764 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x797 &  x800 &  x803 &  x806 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x836 &  x842 &  x845 &  x848 &  x851 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x890 &  x893 &  x896 &  x899 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x950 &  x959 &  x962 &  x965 &  x968 &  x974 &  x977 &  x980 &  x983 &  x989 &  x992 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1025 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1070 &  x1073 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x33 & ~x72 & ~x111 & ~x112 & ~x150 & ~x177 & ~x189 & ~x192 & ~x216 & ~x240 & ~x279 & ~x294 & ~x297 & ~x333 & ~x336 & ~x375 & ~x414 & ~x492 & ~x531;
assign c722 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x49 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x397 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x436 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x475 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x578 &  x584 &  x587 &  x590 &  x593 &  x596 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x626 &  x632 &  x635 &  x638 &  x640 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x754 &  x755 &  x758 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x793 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x827 &  x830 &  x832 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x956 &  x959 &  x962 &  x965 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x393 & ~x432 & ~x433 & ~x472 & ~x510 & ~x549 & ~x550 & ~x588 & ~x589 & ~x627 & ~x666 & ~x918 & ~x957 & ~x996;
assign c724 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x95 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x170 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x206 &  x209 &  x212 &  x218 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x275 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x317 &  x320 &  x322 &  x323 &  x325 &  x326 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x377 &  x383 &  x386 &  x389 &  x391 &  x392 &  x395 &  x398 &  x401 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x430 &  x431 &  x437 &  x440 &  x443 &  x446 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x508 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x530 &  x533 &  x536 &  x539 &  x542 &  x548 &  x551 &  x554 &  x557 &  x560 &  x569 &  x572 &  x575 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x605 &  x611 &  x614 &  x617 &  x620 &  x623 &  x629 &  x632 &  x635 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x689 &  x692 &  x695 &  x698 &  x701 &  x710 &  x713 &  x716 &  x719 &  x722 &  x728 &  x737 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x830 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x860 &  x863 &  x866 &  x869 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x968 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x117 & ~x156 & ~x195 & ~x357 & ~x358 & ~x396 & ~x397 & ~x435 & ~x450 & ~x666 & ~x705 & ~x744 & ~x745 & ~x784 & ~x822;
assign c726 =  x2 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x283 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x322 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x631 &  x632 &  x635 &  x638 &  x644 &  x647 &  x650 &  x653 &  x656 &  x658 &  x659 &  x662 &  x665 &  x668 &  x669 &  x670 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x691 &  x692 &  x695 &  x697 &  x698 &  x701 &  x704 &  x707 &  x708 &  x709 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x730 &  x731 &  x734 &  x736 &  x737 &  x743 &  x746 &  x748 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x769 &  x770 &  x773 &  x775 &  x776 &  x779 &  x782 &  x785 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x633 & ~x672;
assign c728 =  x2 &  x5 &  x8 &  x11 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x59 &  x62 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x119 &  x122 &  x125 &  x127 &  x128 &  x131 &  x134 &  x137 &  x140 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x314 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x352 &  x353 &  x356 &  x362 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x389 &  x391 &  x392 &  x395 &  x401 &  x404 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x452 &  x455 &  x461 &  x464 &  x467 &  x469 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x494 &  x497 &  x500 &  x503 &  x506 &  x508 &  x509 &  x512 &  x515 &  x518 &  x521 &  x523 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x547 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x596 &  x599 &  x600 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x640 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x679 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x710 &  x718 &  x719 &  x722 &  x725 &  x731 &  x734 &  x737 &  x740 &  x743 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x857 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 &  x1130 & ~x201 & ~x240 & ~x342 & ~x381 & ~x675 & ~x714 & ~x744 & ~x753 & ~x783 & ~x822 & ~x861 & ~x939;
assign c730 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x107 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x155 &  x158 &  x161 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x281 &  x284 &  x290 &  x292 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x338 &  x344 &  x347 &  x350 &  x356 &  x359 &  x362 &  x365 &  x368 &  x370 &  x371 &  x374 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x439 &  x440 &  x442 &  x443 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x473 &  x476 &  x479 &  x481 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x509 &  x512 &  x518 &  x520 &  x521 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x559 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x598 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x623 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x671 &  x674 &  x677 &  x683 &  x686 &  x689 &  x692 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x722 &  x725 &  x728 &  x731 &  x737 &  x746 &  x752 &  x755 &  x758 &  x761 &  x764 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x803 &  x806 &  x812 &  x815 &  x818 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x941 &  x944 &  x947 &  x950 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130 & ~x195 & ~x234 & ~x273 & ~x312 & ~x351 & ~x900 & ~x939 & ~x940 & ~x978 & ~x979 & ~x1017;
assign c732 =  x29 &  x38 &  x44 &  x53 &  x65 &  x74 &  x77 &  x83 &  x86 &  x92 &  x104 &  x107 &  x128 &  x134 &  x143 &  x152 &  x155 &  x173 &  x179 &  x185 &  x197 &  x212 &  x218 &  x221 &  x233 &  x248 &  x251 &  x257 &  x260 &  x263 &  x275 &  x293 &  x302 &  x317 &  x335 &  x350 &  x353 &  x359 &  x362 &  x377 &  x383 &  x386 &  x404 &  x425 &  x428 &  x431 &  x434 &  x446 &  x452 &  x479 &  x497 &  x500 &  x506 &  x512 &  x518 &  x530 &  x545 &  x554 &  x581 &  x599 &  x602 &  x608 &  x614 &  x626 &  x634 &  x638 &  x650 &  x656 &  x659 &  x662 &  x674 &  x683 &  x695 &  x698 &  x701 &  x713 &  x715 &  x718 &  x743 &  x758 &  x764 &  x779 &  x785 &  x788 &  x791 &  x794 &  x800 &  x806 &  x812 &  x821 &  x824 &  x842 &  x845 &  x848 &  x890 &  x896 &  x897 &  x902 &  x905 &  x914 &  x917 &  x920 &  x937 &  x941 &  x947 &  x950 &  x953 &  x956 &  x962 &  x975 &  x977 &  x992 &  x1004 &  x1015 &  x1019 &  x1022 &  x1034 &  x1043 &  x1046 &  x1049 &  x1053 &  x1054 &  x1058 &  x1097 &  x1100 &  x1106 &  x1108 &  x1124 & ~x312 & ~x315 & ~x393 & ~x429 & ~x432 & ~x510 & ~x588 & ~x627 & ~x960;
assign c734 =  x1 &  x10 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x40 &  x41 &  x44 &  x47 &  x49 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x78 &  x79 &  x80 &  x83 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x117 &  x118 &  x122 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x156 &  x157 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x188 &  x194 &  x195 &  x196 &  x197 &  x200 &  x203 &  x209 &  x212 &  x215 &  x218 &  x224 &  x227 &  x230 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x269 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x317 &  x320 &  x329 &  x332 &  x335 &  x338 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x428 &  x431 &  x434 &  x437 &  x446 &  x449 &  x455 &  x461 &  x464 &  x467 &  x470 &  x473 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x560 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x599 &  x602 &  x608 &  x611 &  x617 &  x620 &  x626 &  x629 &  x632 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x665 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x758 &  x761 &  x767 &  x770 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x842 &  x848 &  x851 &  x854 &  x857 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x935 &  x941 &  x944 &  x947 &  x950 &  x956 &  x959 &  x962 &  x965 &  x971 &  x974 &  x977 &  x983 &  x986 &  x989 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1052 &  x1055 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 &  x1130 & ~x63 & ~x75 & ~x84 & ~x102 & ~x123 & ~x162 & ~x180 & ~x219 & ~x297 & ~x298 & ~x336 & ~x393 & ~x414 & ~x432 & ~x471 & ~x588;
assign c736 =  x2 &  x11 &  x14 &  x17 &  x23 &  x26 &  x29 &  x35 &  x38 &  x41 &  x47 &  x50 &  x65 &  x68 &  x74 &  x77 &  x86 &  x98 &  x101 &  x107 &  x110 &  x116 &  x119 &  x122 &  x125 &  x131 &  x137 &  x140 &  x143 &  x149 &  x152 &  x158 &  x161 &  x164 &  x166 &  x167 &  x170 &  x185 &  x188 &  x191 &  x194 &  x196 &  x197 &  x200 &  x203 &  x215 &  x227 &  x235 &  x239 &  x242 &  x251 &  x254 &  x263 &  x266 &  x273 &  x274 &  x278 &  x284 &  x287 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x344 &  x350 &  x352 &  x356 &  x374 &  x377 &  x380 &  x386 &  x389 &  x391 &  x392 &  x395 &  x398 &  x410 &  x413 &  x416 &  x419 &  x422 &  x430 &  x431 &  x434 &  x440 &  x443 &  x446 &  x452 &  x455 &  x458 &  x461 &  x469 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x503 &  x506 &  x512 &  x524 &  x530 &  x533 &  x539 &  x542 &  x545 &  x551 &  x554 &  x557 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x587 &  x593 &  x599 &  x602 &  x608 &  x614 &  x617 &  x623 &  x626 &  x638 &  x647 &  x653 &  x665 &  x668 &  x677 &  x680 &  x683 &  x686 &  x695 &  x698 &  x701 &  x707 &  x719 &  x737 &  x740 &  x743 &  x749 &  x755 &  x758 &  x764 &  x770 &  x776 &  x779 &  x782 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x827 &  x830 &  x833 &  x836 &  x839 &  x848 &  x860 &  x866 &  x869 &  x881 &  x884 &  x890 &  x899 &  x905 &  x908 &  x911 &  x914 &  x929 &  x932 &  x938 &  x941 &  x947 &  x950 &  x962 &  x965 &  x977 &  x980 &  x992 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1046 &  x1055 &  x1061 &  x1067 &  x1076 &  x1079 &  x1082 &  x1091 &  x1097 &  x1100 &  x1103 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 & ~x162 & ~x297 & ~x336 & ~x402 & ~x441 & ~x480 & ~x519 & ~x520 & ~x558 & ~x783;
assign c738 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x26 &  x29 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x146 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x197 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x224 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x317 &  x320 &  x323 &  x329 &  x332 &  x335 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x413 &  x416 &  x422 &  x425 &  x428 &  x430 &  x431 &  x434 &  x437 &  x440 &  x443 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x695 &  x697 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x743 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x788 &  x791 &  x794 &  x797 &  x800 &  x809 &  x812 &  x815 &  x818 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x309 & ~x348 & ~x492 & ~x594 & ~x633 & ~x648 & ~x666 & ~x672 & ~x687 & ~x705 & ~x711 & ~x726 & ~x750 & ~x789 & ~x790 & ~x828 & ~x867 & ~x906;
assign c740 =  x17 &  x29 &  x32 &  x35 &  x38 &  x41 &  x48 &  x53 &  x56 &  x71 &  x74 &  x83 &  x88 &  x89 &  x98 &  x113 &  x116 &  x128 &  x131 &  x134 &  x137 &  x143 &  x146 &  x161 &  x173 &  x179 &  x196 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x227 &  x230 &  x234 &  x239 &  x242 &  x245 &  x251 &  x257 &  x266 &  x274 &  x284 &  x287 &  x290 &  x302 &  x313 &  x320 &  x323 &  x335 &  x344 &  x350 &  x365 &  x371 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x413 &  x440 &  x445 &  x464 &  x467 &  x473 &  x479 &  x485 &  x491 &  x506 &  x512 &  x515 &  x524 &  x527 &  x533 &  x542 &  x545 &  x554 &  x557 &  x566 &  x572 &  x581 &  x587 &  x590 &  x596 &  x599 &  x602 &  x614 &  x623 &  x629 &  x635 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x674 &  x677 &  x680 &  x683 &  x686 &  x692 &  x698 &  x701 &  x704 &  x713 &  x716 &  x719 &  x725 &  x728 &  x737 &  x746 &  x749 &  x752 &  x758 &  x761 &  x764 &  x770 &  x791 &  x815 &  x821 &  x824 &  x833 &  x839 &  x842 &  x848 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x875 &  x881 &  x893 &  x896 &  x902 &  x905 &  x911 &  x917 &  x920 &  x923 &  x929 &  x932 &  x938 &  x941 &  x950 &  x959 &  x962 &  x974 &  x977 &  x983 &  x992 &  x1007 &  x1010 &  x1019 &  x1022 &  x1025 &  x1028 &  x1037 &  x1040 &  x1046 &  x1049 &  x1055 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 & ~x84 & ~x144 & ~x183 & ~x219 & ~x369 & ~x408 & ~x432 & ~x471 & ~x549 & ~x588;
assign c742 =  x8 &  x20 &  x23 &  x38 &  x44 &  x68 &  x80 &  x92 &  x95 &  x98 &  x110 &  x116 &  x119 &  x122 &  x134 &  x137 &  x140 &  x152 &  x167 &  x173 &  x176 &  x179 &  x182 &  x185 &  x194 &  x212 &  x215 &  x218 &  x224 &  x227 &  x239 &  x245 &  x254 &  x269 &  x275 &  x281 &  x293 &  x296 &  x308 &  x323 &  x326 &  x329 &  x335 &  x347 &  x350 &  x353 &  x368 &  x376 &  x395 &  x401 &  x413 &  x419 &  x434 &  x437 &  x440 &  x443 &  x446 &  x473 &  x479 &  x482 &  x494 &  x518 &  x521 &  x524 &  x527 &  x530 &  x539 &  x545 &  x548 &  x551 &  x554 &  x563 &  x584 &  x596 &  x602 &  x611 &  x617 &  x620 &  x623 &  x632 &  x644 &  x647 &  x653 &  x656 &  x665 &  x668 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x713 &  x722 &  x725 &  x731 &  x737 &  x742 &  x752 &  x755 &  x767 &  x773 &  x781 &  x788 &  x794 &  x797 &  x809 &  x812 &  x815 &  x818 &  x820 &  x848 &  x854 &  x860 &  x872 &  x878 &  x884 &  x887 &  x893 &  x905 &  x908 &  x911 &  x923 &  x932 &  x935 &  x944 &  x947 &  x950 &  x956 &  x962 &  x968 &  x974 &  x977 &  x980 &  x989 &  x998 &  x1022 &  x1025 &  x1043 &  x1049 &  x1064 &  x1070 &  x1076 &  x1082 &  x1085 &  x1094 &  x1100 &  x1127 & ~x393 & ~x432 & ~x882 & ~x922 & ~x994 & ~x1017 & ~x1032 & ~x1071 & ~x1072;
assign c744 =  x2 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x29 &  x32 &  x35 &  x41 &  x44 &  x47 &  x50 &  x53 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x83 &  x86 &  x89 &  x92 &  x107 &  x110 &  x119 &  x122 &  x128 &  x131 &  x134 &  x137 &  x140 &  x152 &  x164 &  x167 &  x170 &  x173 &  x176 &  x185 &  x191 &  x194 &  x197 &  x200 &  x206 &  x212 &  x218 &  x221 &  x227 &  x230 &  x239 &  x248 &  x251 &  x254 &  x257 &  x263 &  x266 &  x269 &  x278 &  x281 &  x283 &  x287 &  x299 &  x302 &  x305 &  x308 &  x317 &  x321 &  x322 &  x323 &  x326 &  x329 &  x332 &  x335 &  x341 &  x344 &  x347 &  x352 &  x356 &  x359 &  x361 &  x362 &  x365 &  x371 &  x383 &  x389 &  x391 &  x392 &  x401 &  x404 &  x407 &  x410 &  x413 &  x419 &  x422 &  x425 &  x428 &  x430 &  x431 &  x440 &  x443 &  x446 &  x449 &  x455 &  x464 &  x467 &  x469 &  x470 &  x473 &  x476 &  x479 &  x485 &  x488 &  x491 &  x494 &  x503 &  x508 &  x509 &  x512 &  x515 &  x521 &  x524 &  x530 &  x533 &  x536 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x581 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x638 &  x653 &  x656 &  x659 &  x668 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x695 &  x698 &  x701 &  x704 &  x707 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x743 &  x746 &  x749 &  x752 &  x755 &  x761 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x794 &  x800 &  x803 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x836 &  x839 &  x842 &  x848 &  x851 &  x857 &  x866 &  x875 &  x878 &  x881 &  x887 &  x893 &  x896 &  x899 &  x902 &  x908 &  x911 &  x914 &  x917 &  x919 &  x920 &  x923 &  x926 &  x929 &  x935 &  x950 &  x953 &  x956 &  x959 &  x962 &  x968 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x998 &  x1007 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1037 &  x1043 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1115 &  x1118 &  x1124 &  x1130 & ~x357 & ~x396 & ~x435 & ~x489 & ~x492 & ~x531 & ~x705 & ~x706 & ~x744 & ~x745 & ~x783 & ~x822 & ~x861;
assign c746 =  x5 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x83 &  x86 &  x89 &  x92 &  x98 &  x101 &  x104 &  x110 &  x113 &  x119 &  x122 &  x125 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x167 &  x170 &  x173 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x230 &  x239 &  x242 &  x245 &  x248 &  x257 &  x260 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x380 &  x383 &  x389 &  x395 &  x398 &  x401 &  x403 &  x404 &  x407 &  x410 &  x413 &  x416 &  x425 &  x428 &  x434 &  x437 &  x440 &  x442 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x481 &  x485 &  x488 &  x491 &  x497 &  x500 &  x503 &  x509 &  x512 &  x518 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x554 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x578 &  x584 &  x587 &  x593 &  x596 &  x599 &  x602 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x644 &  x647 &  x650 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x689 &  x701 &  x704 &  x707 &  x710 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x743 &  x746 &  x749 &  x758 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x818 &  x821 &  x824 &  x830 &  x833 &  x836 &  x842 &  x848 &  x851 &  x854 &  x860 &  x866 &  x869 &  x878 &  x887 &  x890 &  x893 &  x896 &  x899 &  x905 &  x908 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x965 &  x968 &  x974 &  x977 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x156 & ~x234 & ~x687 & ~x726 & ~x861 & ~x901 & ~x939 & ~x940 & ~x978 & ~x987 & ~x1026 & ~x1056 & ~x1065 & ~x1104;
assign c748 =  x2 &  x5 &  x8 &  x14 &  x17 &  x23 &  x29 &  x32 &  x35 &  x38 &  x41 &  x47 &  x50 &  x53 &  x59 &  x62 &  x65 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x314 &  x317 &  x320 &  x323 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x391 &  x392 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x446 &  x452 &  x458 &  x461 &  x467 &  x469 &  x470 &  x473 &  x476 &  x479 &  x485 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x554 &  x557 &  x560 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x623 &  x626 &  x629 &  x632 &  x635 &  x640 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x680 &  x683 &  x686 &  x689 &  x692 &  x697 &  x701 &  x704 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x730 &  x734 &  x737 &  x740 &  x746 &  x749 &  x755 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x794 &  x800 &  x803 &  x812 &  x814 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x842 &  x845 &  x848 &  x851 &  x857 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x917 &  x920 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x950 &  x956 &  x959 &  x965 &  x968 &  x971 &  x977 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1058 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x201 & ~x279 & ~x318 & ~x357 & ~x411 & ~x627 & ~x666 & ~x667 & ~x705 & ~x706 & ~x744 & ~x745 & ~x783 & ~x822 & ~x849;
assign c750 =  x2 &  x5 &  x8 &  x11 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x53 &  x59 &  x65 &  x71 &  x74 &  x77 &  x86 &  x92 &  x95 &  x98 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x149 &  x152 &  x155 &  x158 &  x164 &  x173 &  x179 &  x182 &  x185 &  x191 &  x194 &  x197 &  x206 &  x215 &  x221 &  x236 &  x239 &  x242 &  x248 &  x251 &  x257 &  x260 &  x269 &  x272 &  x275 &  x293 &  x296 &  x299 &  x302 &  x305 &  x320 &  x332 &  x335 &  x338 &  x344 &  x347 &  x353 &  x365 &  x368 &  x374 &  x377 &  x386 &  x389 &  x395 &  x401 &  x407 &  x428 &  x431 &  x437 &  x440 &  x455 &  x458 &  x461 &  x470 &  x473 &  x479 &  x482 &  x485 &  x491 &  x500 &  x506 &  x515 &  x520 &  x521 &  x527 &  x536 &  x545 &  x554 &  x560 &  x572 &  x575 &  x578 &  x581 &  x587 &  x590 &  x593 &  x596 &  x602 &  x605 &  x608 &  x614 &  x617 &  x620 &  x623 &  x626 &  x635 &  x638 &  x644 &  x659 &  x662 &  x671 &  x674 &  x677 &  x683 &  x686 &  x695 &  x701 &  x710 &  x716 &  x719 &  x722 &  x725 &  x737 &  x740 &  x742 &  x743 &  x755 &  x758 &  x764 &  x767 &  x770 &  x773 &  x779 &  x785 &  x788 &  x797 &  x803 &  x809 &  x812 &  x815 &  x820 &  x830 &  x836 &  x845 &  x854 &  x857 &  x866 &  x869 &  x875 &  x881 &  x887 &  x890 &  x896 &  x899 &  x902 &  x905 &  x911 &  x913 &  x914 &  x920 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x953 &  x959 &  x962 &  x977 &  x992 &  x998 &  x1010 &  x1013 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1052 &  x1055 &  x1058 &  x1060 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1099 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 & ~x234 & ~x312 & ~x540 & ~x939 & ~x978 & ~x993;
assign c752 =  x2 &  x5 &  x8 &  x14 &  x20 &  x23 &  x26 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x62 &  x65 &  x71 &  x95 &  x98 &  x104 &  x116 &  x119 &  x128 &  x131 &  x137 &  x143 &  x146 &  x152 &  x155 &  x161 &  x170 &  x173 &  x176 &  x179 &  x188 &  x200 &  x206 &  x209 &  x221 &  x230 &  x236 &  x242 &  x245 &  x254 &  x257 &  x275 &  x278 &  x293 &  x299 &  x302 &  x338 &  x344 &  x350 &  x359 &  x362 &  x365 &  x368 &  x383 &  x386 &  x392 &  x401 &  x407 &  x419 &  x422 &  x431 &  x437 &  x440 &  x446 &  x449 &  x470 &  x482 &  x485 &  x488 &  x500 &  x503 &  x506 &  x509 &  x512 &  x518 &  x527 &  x539 &  x545 &  x548 &  x554 &  x560 &  x563 &  x581 &  x587 &  x593 &  x596 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x635 &  x637 &  x641 &  x647 &  x653 &  x665 &  x674 &  x683 &  x692 &  x698 &  x713 &  x719 &  x722 &  x725 &  x728 &  x752 &  x761 &  x767 &  x773 &  x806 &  x809 &  x812 &  x818 &  x820 &  x824 &  x830 &  x833 &  x836 &  x842 &  x860 &  x866 &  x869 &  x896 &  x898 &  x905 &  x914 &  x917 &  x920 &  x923 &  x932 &  x937 &  x956 &  x965 &  x976 &  x977 &  x980 &  x983 &  x986 &  x995 &  x1010 &  x1013 &  x1015 &  x1016 &  x1019 &  x1025 &  x1031 &  x1034 &  x1040 &  x1046 &  x1061 &  x1067 &  x1070 &  x1076 &  x1082 &  x1087 &  x1088 &  x1091 &  x1093 &  x1094 &  x1106 &  x1121 &  x1124 &  x1127 &  x1130 & ~x273 & ~x276 & ~x390 & ~x432 & ~x471 & ~x915 & ~x922 & ~x954 & ~x961 & ~x993 & ~x999 & ~x1000 & ~x1039 & ~x1110 & ~x1116;
assign c754 =  x2 &  x11 &  x17 &  x20 &  x26 &  x35 &  x47 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x95 &  x101 &  x107 &  x110 &  x116 &  x119 &  x128 &  x131 &  x137 &  x143 &  x149 &  x155 &  x164 &  x170 &  x173 &  x179 &  x182 &  x185 &  x188 &  x194 &  x200 &  x203 &  x206 &  x218 &  x226 &  x230 &  x239 &  x248 &  x251 &  x257 &  x260 &  x293 &  x304 &  x311 &  x317 &  x329 &  x338 &  x344 &  x347 &  x356 &  x365 &  x368 &  x377 &  x380 &  x383 &  x401 &  x415 &  x419 &  x422 &  x427 &  x428 &  x431 &  x443 &  x446 &  x449 &  x458 &  x461 &  x464 &  x494 &  x503 &  x506 &  x509 &  x524 &  x536 &  x539 &  x542 &  x563 &  x566 &  x575 &  x578 &  x581 &  x587 &  x590 &  x601 &  x605 &  x611 &  x614 &  x617 &  x626 &  x637 &  x638 &  x644 &  x650 &  x653 &  x665 &  x673 &  x704 &  x707 &  x711 &  x713 &  x716 &  x719 &  x725 &  x728 &  x731 &  x734 &  x746 &  x755 &  x761 &  x764 &  x767 &  x773 &  x791 &  x794 &  x800 &  x803 &  x809 &  x812 &  x815 &  x821 &  x824 &  x827 &  x839 &  x845 &  x857 &  x859 &  x860 &  x866 &  x872 &  x875 &  x884 &  x887 &  x898 &  x899 &  x908 &  x911 &  x914 &  x935 &  x941 &  x950 &  x956 &  x965 &  x968 &  x976 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1019 &  x1028 &  x1031 &  x1040 &  x1054 &  x1091 &  x1097 &  x1130 & ~x234 & ~x273 & ~x390 & ~x468 & ~x507 & ~x960;
assign c756 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x391 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x430 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x469 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x631 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x669 &  x670 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x708 &  x709 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x747 &  x748 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x787 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x826 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x851 &  x854 &  x857 &  x860 &  x863 &  x865 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x453 & ~x531 & ~x564 & ~x570 & ~x666 & ~x667 & ~x705 & ~x706 & ~x744 & ~x783 & ~x822;
assign c758 =  x5 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x47 &  x50 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x80 &  x89 &  x92 &  x95 &  x98 &  x104 &  x113 &  x116 &  x119 &  x125 &  x128 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x185 &  x188 &  x194 &  x197 &  x200 &  x203 &  x212 &  x218 &  x221 &  x227 &  x230 &  x233 &  x239 &  x251 &  x257 &  x260 &  x266 &  x269 &  x278 &  x281 &  x287 &  x290 &  x299 &  x302 &  x304 &  x305 &  x308 &  x311 &  x326 &  x332 &  x335 &  x337 &  x341 &  x343 &  x356 &  x359 &  x362 &  x365 &  x368 &  x377 &  x380 &  x383 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x409 &  x410 &  x413 &  x422 &  x428 &  x443 &  x446 &  x448 &  x458 &  x461 &  x473 &  x476 &  x479 &  x481 &  x485 &  x488 &  x491 &  x497 &  x503 &  x506 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x560 &  x566 &  x569 &  x575 &  x578 &  x581 &  x584 &  x587 &  x593 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x629 &  x638 &  x653 &  x659 &  x665 &  x668 &  x671 &  x672 &  x673 &  x674 &  x677 &  x680 &  x683 &  x689 &  x692 &  x698 &  x701 &  x712 &  x713 &  x716 &  x719 &  x725 &  x734 &  x737 &  x749 &  x761 &  x764 &  x770 &  x773 &  x776 &  x791 &  x794 &  x809 &  x812 &  x815 &  x827 &  x833 &  x836 &  x848 &  x854 &  x857 &  x866 &  x884 &  x893 &  x896 &  x899 &  x905 &  x908 &  x917 &  x923 &  x929 &  x935 &  x941 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x989 &  x1001 &  x1010 &  x1022 &  x1030 &  x1031 &  x1040 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1069 &  x1079 &  x1082 &  x1085 &  x1091 &  x1100 &  x1103 &  x1108 &  x1124 &  x1127 &  x1130 & ~x1056;
assign c760 =  x2 &  x5 &  x8 &  x11 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x152 &  x155 &  x158 &  x161 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x631 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x670 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x708 &  x709 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x747 &  x748 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x787 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x865 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x192 & ~x372 & ~x411 & ~x666 & ~x705 & ~x706 & ~x744 & ~x745 & ~x783 & ~x822 & ~x861;
assign c762 =  x5 &  x11 &  x23 &  x26 &  x32 &  x47 &  x53 &  x68 &  x74 &  x77 &  x80 &  x101 &  x113 &  x116 &  x119 &  x128 &  x134 &  x137 &  x140 &  x146 &  x149 &  x158 &  x164 &  x170 &  x179 &  x191 &  x194 &  x197 &  x200 &  x206 &  x218 &  x227 &  x239 &  x242 &  x245 &  x254 &  x257 &  x259 &  x272 &  x284 &  x287 &  x290 &  x308 &  x314 &  x323 &  x326 &  x329 &  x335 &  x341 &  x353 &  x356 &  x359 &  x362 &  x365 &  x374 &  x380 &  x386 &  x395 &  x398 &  x412 &  x416 &  x419 &  x425 &  x434 &  x437 &  x442 &  x446 &  x458 &  x464 &  x476 &  x488 &  x494 &  x499 &  x503 &  x509 &  x515 &  x518 &  x521 &  x533 &  x548 &  x554 &  x560 &  x575 &  x581 &  x602 &  x608 &  x611 &  x614 &  x629 &  x632 &  x637 &  x638 &  x650 &  x653 &  x656 &  x659 &  x665 &  x671 &  x676 &  x692 &  x707 &  x713 &  x716 &  x718 &  x725 &  x737 &  x740 &  x746 &  x749 &  x752 &  x754 &  x755 &  x758 &  x785 &  x788 &  x791 &  x797 &  x815 &  x818 &  x824 &  x845 &  x851 &  x854 &  x860 &  x866 &  x872 &  x878 &  x881 &  x884 &  x896 &  x897 &  x898 &  x911 &  x914 &  x917 &  x935 &  x938 &  x941 &  x956 &  x965 &  x968 &  x974 &  x975 &  x976 &  x983 &  x991 &  x992 &  x995 &  x998 &  x1013 &  x1022 &  x1028 &  x1034 &  x1040 &  x1046 &  x1049 &  x1052 &  x1061 &  x1069 &  x1076 &  x1088 &  x1107 &  x1112 &  x1124 &  x1127 & ~x354 & ~x471;
assign c764 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x176 &  x179 &  x182 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x266 &  x269 &  x272 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x389 &  x395 &  x398 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x569 &  x572 &  x578 &  x581 &  x584 &  x590 &  x593 &  x599 &  x602 &  x608 &  x611 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x701 &  x704 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x866 &  x869 &  x872 &  x874 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x896 &  x899 &  x902 &  x905 &  x908 &  x913 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x609 & ~x648 & ~x687 & ~x726 & ~x750 & ~x765 & ~x789 & ~x828 & ~x829 & ~x843 & ~x861 & ~x867 & ~x868 & ~x882 & ~x906 & ~x907 & ~x921 & ~x945 & ~x960 & ~x984 & ~x999 & ~x1011;
assign c766 =  x2 &  x5 &  x17 &  x23 &  x26 &  x29 &  x32 &  x35 &  x47 &  x56 &  x59 &  x65 &  x74 &  x80 &  x92 &  x98 &  x107 &  x110 &  x113 &  x137 &  x143 &  x161 &  x167 &  x170 &  x173 &  x182 &  x185 &  x200 &  x239 &  x245 &  x248 &  x251 &  x259 &  x260 &  x278 &  x281 &  x293 &  x298 &  x311 &  x314 &  x329 &  x332 &  x335 &  x343 &  x350 &  x353 &  x359 &  x368 &  x376 &  x380 &  x383 &  x395 &  x401 &  x413 &  x416 &  x431 &  x452 &  x455 &  x458 &  x467 &  x473 &  x476 &  x482 &  x488 &  x497 &  x506 &  x509 &  x515 &  x524 &  x527 &  x557 &  x563 &  x566 &  x584 &  x587 &  x590 &  x593 &  x596 &  x605 &  x608 &  x620 &  x635 &  x638 &  x641 &  x647 &  x659 &  x662 &  x671 &  x686 &  x692 &  x695 &  x698 &  x704 &  x707 &  x710 &  x716 &  x719 &  x728 &  x731 &  x749 &  x755 &  x761 &  x767 &  x770 &  x788 &  x803 &  x809 &  x830 &  x836 &  x848 &  x854 &  x866 &  x884 &  x887 &  x890 &  x896 &  x902 &  x908 &  x929 &  x938 &  x944 &  x950 &  x953 &  x956 &  x962 &  x965 &  x974 &  x980 &  x982 &  x986 &  x992 &  x995 &  x1001 &  x1007 &  x1021 &  x1022 &  x1034 &  x1037 &  x1040 &  x1043 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1094 &  x1099 &  x1100 &  x1109 &  x1112 &  x1115 &  x1127 & ~x312 & ~x351 & ~x837 & ~x843 & ~x882 & ~x978 & ~x1116;
assign c768 =  x2 &  x5 &  x8 &  x13 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x50 &  x52 &  x53 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x89 &  x91 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x146 &  x149 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x208 &  x209 &  x212 &  x215 &  x218 &  x224 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x254 &  x257 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x437 &  x440 &  x443 &  x449 &  x455 &  x458 &  x464 &  x467 &  x470 &  x473 &  x475 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x514 &  x515 &  x518 &  x521 &  x523 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x560 &  x562 &  x563 &  x566 &  x569 &  x572 &  x575 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x640 &  x641 &  x644 &  x647 &  x649 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x688 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x728 &  x731 &  x737 &  x740 &  x743 &  x746 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x812 &  x818 &  x821 &  x824 &  x827 &  x830 &  x836 &  x839 &  x845 &  x848 &  x851 &  x854 &  x857 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1127 &  x1130 & ~x471 & ~x510 & ~x744 & ~x780 & ~x783 & ~x1002 & ~x1041;
assign c770 =  x2 &  x5 &  x8 &  x14 &  x17 &  x26 &  x41 &  x44 &  x47 &  x52 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x86 &  x92 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x119 &  x122 &  x134 &  x149 &  x152 &  x155 &  x161 &  x173 &  x182 &  x185 &  x188 &  x191 &  x194 &  x200 &  x203 &  x206 &  x212 &  x215 &  x218 &  x227 &  x233 &  x239 &  x245 &  x248 &  x254 &  x272 &  x274 &  x275 &  x284 &  x287 &  x293 &  x305 &  x311 &  x313 &  x314 &  x320 &  x323 &  x326 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x356 &  x362 &  x365 &  x371 &  x374 &  x377 &  x383 &  x386 &  x395 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x452 &  x455 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x485 &  x488 &  x491 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x524 &  x527 &  x533 &  x536 &  x539 &  x545 &  x548 &  x551 &  x554 &  x557 &  x563 &  x569 &  x572 &  x575 &  x581 &  x584 &  x587 &  x590 &  x593 &  x599 &  x605 &  x608 &  x614 &  x623 &  x626 &  x629 &  x632 &  x641 &  x644 &  x650 &  x652 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x674 &  x677 &  x686 &  x689 &  x695 &  x698 &  x701 &  x704 &  x707 &  x716 &  x719 &  x722 &  x728 &  x731 &  x734 &  x740 &  x743 &  x749 &  x752 &  x755 &  x758 &  x761 &  x767 &  x770 &  x773 &  x779 &  x785 &  x788 &  x800 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x833 &  x839 &  x845 &  x848 &  x851 &  x857 &  x860 &  x863 &  x866 &  x872 &  x875 &  x878 &  x881 &  x893 &  x899 &  x902 &  x908 &  x911 &  x914 &  x920 &  x926 &  x932 &  x941 &  x947 &  x950 &  x953 &  x956 &  x965 &  x968 &  x971 &  x974 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1034 &  x1037 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1070 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1115 &  x1121 &  x1124 &  x1127 & ~x297 & ~x336 & ~x453 & ~x492 & ~x531 & ~x588 & ~x628 & ~x666 & ~x741 & ~x819 & ~x858 & ~x897 & ~x912 & ~x936 & ~x951 & ~x1107;
assign c772 =  x2 &  x8 &  x11 &  x14 &  x20 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x56 &  x65 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x107 &  x110 &  x122 &  x128 &  x134 &  x140 &  x143 &  x146 &  x149 &  x155 &  x161 &  x164 &  x167 &  x173 &  x179 &  x188 &  x191 &  x197 &  x212 &  x215 &  x221 &  x227 &  x233 &  x236 &  x239 &  x245 &  x254 &  x257 &  x260 &  x269 &  x272 &  x275 &  x278 &  x281 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x329 &  x332 &  x341 &  x350 &  x356 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x380 &  x383 &  x389 &  x395 &  x398 &  x401 &  x404 &  x407 &  x413 &  x416 &  x425 &  x428 &  x431 &  x434 &  x437 &  x446 &  x449 &  x458 &  x461 &  x464 &  x467 &  x479 &  x482 &  x485 &  x491 &  x497 &  x500 &  x503 &  x506 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x542 &  x545 &  x548 &  x557 &  x560 &  x566 &  x572 &  x581 &  x584 &  x590 &  x596 &  x599 &  x605 &  x608 &  x611 &  x614 &  x635 &  x638 &  x644 &  x647 &  x650 &  x656 &  x662 &  x664 &  x665 &  x668 &  x671 &  x677 &  x683 &  x692 &  x698 &  x701 &  x703 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x734 &  x743 &  x752 &  x755 &  x770 &  x779 &  x782 &  x788 &  x791 &  x794 &  x803 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x839 &  x842 &  x848 &  x854 &  x860 &  x863 &  x869 &  x884 &  x887 &  x905 &  x911 &  x914 &  x917 &  x923 &  x932 &  x938 &  x944 &  x947 &  x959 &  x965 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x992 &  x998 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1025 &  x1031 &  x1034 &  x1046 &  x1049 &  x1070 &  x1073 &  x1076 &  x1079 &  x1088 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1118 &  x1124 &  x1130 & ~x3 & ~x42 & ~x81 & ~x120 & ~x159 & ~x198 & ~x276 & ~x315 & ~x393 & ~x471 & ~x645 & ~x684 & ~x726 & ~x804 & ~x843 & ~x882 & ~x939 & ~x940 & ~x1095;
assign c774 =  x2 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x87 &  x88 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x127 &  x128 &  x131 &  x134 &  x137 &  x143 &  x146 &  x149 &  x152 &  x155 &  x157 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x185 &  x188 &  x191 &  x194 &  x196 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x235 &  x236 &  x239 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x272 &  x274 &  x275 &  x278 &  x281 &  x284 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x317 &  x320 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x392 &  x395 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x566 &  x569 &  x572 &  x575 &  x587 &  x593 &  x596 &  x599 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x632 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x740 &  x743 &  x746 &  x749 &  x755 &  x758 &  x767 &  x773 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x857 &  x863 &  x866 &  x869 &  x872 &  x875 &  x881 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x911 &  x914 &  x920 &  x923 &  x926 &  x929 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x983 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1064 &  x1067 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x177 & ~x180 & ~x219 & ~x255 & ~x294 & ~x297 & ~x330 & ~x369 & ~x375 & ~x408 & ~x471 & ~x510 & ~x549 & ~x550 & ~x588 & ~x627 & ~x663 & ~x783 & ~x822;
assign c776 =  x2 &  x8 &  x11 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x62 &  x74 &  x77 &  x80 &  x83 &  x88 &  x92 &  x95 &  x104 &  x107 &  x110 &  x113 &  x125 &  x140 &  x143 &  x146 &  x155 &  x158 &  x164 &  x170 &  x179 &  x182 &  x194 &  x196 &  x197 &  x200 &  x206 &  x221 &  x227 &  x235 &  x242 &  x245 &  x251 &  x260 &  x272 &  x278 &  x281 &  x287 &  x293 &  x299 &  x302 &  x311 &  x313 &  x314 &  x323 &  x335 &  x338 &  x344 &  x353 &  x365 &  x368 &  x377 &  x380 &  x383 &  x386 &  x395 &  x401 &  x407 &  x419 &  x428 &  x431 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x467 &  x470 &  x473 &  x479 &  x482 &  x488 &  x491 &  x494 &  x503 &  x506 &  x512 &  x521 &  x524 &  x529 &  x530 &  x533 &  x536 &  x551 &  x554 &  x557 &  x560 &  x562 &  x563 &  x568 &  x569 &  x572 &  x578 &  x584 &  x587 &  x590 &  x596 &  x599 &  x617 &  x629 &  x632 &  x638 &  x644 &  x646 &  x650 &  x656 &  x662 &  x665 &  x668 &  x680 &  x683 &  x689 &  x692 &  x698 &  x701 &  x704 &  x710 &  x713 &  x716 &  x719 &  x731 &  x758 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x794 &  x806 &  x815 &  x818 &  x824 &  x830 &  x833 &  x839 &  x842 &  x848 &  x854 &  x857 &  x863 &  x869 &  x872 &  x875 &  x881 &  x893 &  x896 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x926 &  x935 &  x938 &  x947 &  x953 &  x956 &  x959 &  x962 &  x965 &  x974 &  x977 &  x980 &  x986 &  x992 &  x995 &  x1010 &  x1013 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1061 &  x1073 &  x1076 &  x1079 &  x1085 &  x1091 &  x1094 &  x1097 &  x1103 &  x1115 &  x1118 & ~x201 & ~x219 & ~x258 & ~x297 & ~x336 & ~x337 & ~x510 & ~x549 & ~x550 & ~x588 & ~x705 & ~x936;
assign c778 =  x5 &  x8 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x50 &  x56 &  x59 &  x62 &  x65 &  x71 &  x77 &  x83 &  x89 &  x92 &  x95 &  x101 &  x104 &  x107 &  x122 &  x125 &  x131 &  x137 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x212 &  x215 &  x221 &  x236 &  x245 &  x254 &  x257 &  x260 &  x263 &  x272 &  x278 &  x281 &  x284 &  x285 &  x286 &  x287 &  x290 &  x293 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x325 &  x329 &  x332 &  x338 &  x350 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x394 &  x395 &  x401 &  x404 &  x410 &  x413 &  x419 &  x422 &  x429 &  x430 &  x431 &  x440 &  x443 &  x449 &  x452 &  x455 &  x458 &  x464 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x503 &  x508 &  x509 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x539 &  x545 &  x547 &  x548 &  x551 &  x563 &  x572 &  x575 &  x581 &  x584 &  x590 &  x593 &  x596 &  x599 &  x617 &  x623 &  x626 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x701 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x743 &  x749 &  x752 &  x758 &  x764 &  x767 &  x770 &  x776 &  x782 &  x785 &  x791 &  x794 &  x797 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x830 &  x836 &  x839 &  x842 &  x845 &  x854 &  x860 &  x863 &  x866 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x941 &  x944 &  x950 &  x953 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x989 &  x992 &  x998 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 & ~x318 & ~x357 & ~x666 & ~x705 & ~x706 & ~x744 & ~x745 & ~x783 & ~x784;
assign c780 =  x5 &  x8 &  x11 &  x17 &  x20 &  x26 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x49 &  x53 &  x59 &  x65 &  x68 &  x77 &  x86 &  x98 &  x107 &  x113 &  x116 &  x117 &  x118 &  x119 &  x122 &  x128 &  x134 &  x143 &  x146 &  x155 &  x156 &  x157 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x182 &  x188 &  x194 &  x196 &  x203 &  x206 &  x209 &  x230 &  x233 &  x239 &  x242 &  x254 &  x257 &  x260 &  x263 &  x266 &  x272 &  x278 &  x281 &  x284 &  x287 &  x293 &  x299 &  x302 &  x305 &  x311 &  x317 &  x323 &  x326 &  x335 &  x344 &  x350 &  x359 &  x362 &  x368 &  x374 &  x395 &  x410 &  x416 &  x419 &  x422 &  x428 &  x431 &  x437 &  x446 &  x452 &  x455 &  x457 &  x458 &  x461 &  x464 &  x473 &  x476 &  x479 &  x485 &  x491 &  x497 &  x500 &  x503 &  x512 &  x515 &  x536 &  x539 &  x545 &  x548 &  x551 &  x554 &  x557 &  x563 &  x566 &  x578 &  x584 &  x587 &  x593 &  x596 &  x602 &  x605 &  x614 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x656 &  x659 &  x662 &  x665 &  x671 &  x674 &  x677 &  x689 &  x692 &  x695 &  x701 &  x707 &  x713 &  x721 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x746 &  x755 &  x760 &  x767 &  x770 &  x773 &  x776 &  x782 &  x788 &  x791 &  x794 &  x797 &  x806 &  x809 &  x812 &  x815 &  x821 &  x824 &  x827 &  x833 &  x836 &  x845 &  x848 &  x851 &  x854 &  x863 &  x866 &  x875 &  x878 &  x881 &  x890 &  x896 &  x902 &  x905 &  x908 &  x914 &  x917 &  x920 &  x926 &  x932 &  x938 &  x941 &  x950 &  x953 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x992 &  x1004 &  x1010 &  x1019 &  x1022 &  x1031 &  x1034 &  x1037 &  x1046 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1076 &  x1079 &  x1082 &  x1094 &  x1097 &  x1103 &  x1109 &  x1112 &  x1121 &  x1130 & ~x141 & ~x174 & ~x180 & ~x297 & ~x369 & ~x408 & ~x432 & ~x433 & ~x472 & ~x510 & ~x511 & ~x549 & ~x588 & ~x663 & ~x666 & ~x705 & ~x858;
assign c782 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x360 &  x361 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x400 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x430 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x469 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x508 &  x509 &  x512 &  x518 &  x521 &  x524 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x547 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x623 &  x626 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x863 &  x866 &  x869 &  x875 &  x878 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x950 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x78 & ~x117 & ~x156 & ~x195 & ~x396 & ~x411 & ~x435 & ~x450 & ~x489 & ~x705 & ~x744 & ~x783 & ~x784 & ~x822 & ~x861;
assign c784 =  x2 &  x8 &  x11 &  x14 &  x20 &  x26 &  x50 &  x53 &  x59 &  x62 &  x71 &  x83 &  x95 &  x113 &  x122 &  x125 &  x134 &  x137 &  x140 &  x143 &  x152 &  x173 &  x176 &  x182 &  x191 &  x200 &  x203 &  x218 &  x221 &  x224 &  x236 &  x242 &  x260 &  x266 &  x278 &  x287 &  x299 &  x320 &  x324 &  x326 &  x329 &  x335 &  x338 &  x341 &  x347 &  x356 &  x360 &  x362 &  x371 &  x380 &  x383 &  x392 &  x401 &  x404 &  x413 &  x416 &  x419 &  x422 &  x430 &  x434 &  x442 &  x443 &  x452 &  x467 &  x476 &  x482 &  x500 &  x506 &  x508 &  x512 &  x515 &  x533 &  x547 &  x554 &  x557 &  x560 &  x572 &  x584 &  x599 &  x602 &  x608 &  x614 &  x620 &  x625 &  x632 &  x635 &  x641 &  x659 &  x662 &  x677 &  x680 &  x689 &  x701 &  x703 &  x704 &  x707 &  x713 &  x716 &  x719 &  x725 &  x731 &  x737 &  x743 &  x749 &  x752 &  x764 &  x767 &  x791 &  x794 &  x800 &  x815 &  x818 &  x821 &  x827 &  x830 &  x836 &  x863 &  x884 &  x887 &  x890 &  x905 &  x917 &  x920 &  x923 &  x935 &  x941 &  x944 &  x947 &  x959 &  x962 &  x968 &  x980 &  x983 &  x986 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1019 &  x1022 &  x1025 &  x1028 &  x1034 &  x1043 &  x1055 &  x1058 &  x1064 &  x1067 &  x1082 &  x1085 &  x1091 &  x1097 &  x1100 &  x1106 &  x1118 &  x1127 & ~x426 & ~x744 & ~x784 & ~x822 & ~x861;
assign c786 =  x5 &  x17 &  x23 &  x26 &  x29 &  x32 &  x35 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x65 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x97 &  x98 &  x101 &  x107 &  x110 &  x113 &  x116 &  x119 &  x125 &  x130 &  x131 &  x137 &  x140 &  x143 &  x146 &  x149 &  x155 &  x158 &  x161 &  x164 &  x167 &  x169 &  x173 &  x176 &  x188 &  x194 &  x203 &  x204 &  x206 &  x209 &  x212 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x243 &  x244 &  x245 &  x247 &  x248 &  x251 &  x254 &  x260 &  x266 &  x275 &  x283 &  x284 &  x287 &  x293 &  x299 &  x302 &  x308 &  x311 &  x326 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x419 &  x425 &  x428 &  x431 &  x434 &  x440 &  x443 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x473 &  x476 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x518 &  x521 &  x530 &  x536 &  x539 &  x542 &  x551 &  x554 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x587 &  x593 &  x596 &  x602 &  x605 &  x614 &  x620 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x680 &  x686 &  x695 &  x698 &  x704 &  x707 &  x716 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x770 &  x779 &  x788 &  x791 &  x794 &  x803 &  x806 &  x809 &  x812 &  x815 &  x824 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x854 &  x863 &  x884 &  x890 &  x893 &  x896 &  x899 &  x911 &  x914 &  x929 &  x932 &  x935 &  x938 &  x947 &  x950 &  x962 &  x968 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1031 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1064 &  x1067 &  x1073 &  x1082 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 &  x1130 & ~x264 & ~x306 & ~x627 & ~x705 & ~x706 & ~x783 & ~x822;
assign c788 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x59 &  x62 &  x65 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x439 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x478 &  x479 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x625 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x703 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x742 &  x743 &  x746 &  x749 &  x752 &  x755 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x781 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x820 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x859 &  x860 &  x863 &  x866 &  x869 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x315 & ~x354 & ~x393 & ~x432 & ~x471 & ~x513 & ~x552 & ~x591 & ~x606 & ~x726 & ~x765 & ~x900 & ~x939 & ~x940 & ~x978 & ~x979 & ~x1056;
assign c790 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x166 &  x167 &  x170 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x205 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x235 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x274 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x391 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x430 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x548 &  x551 &  x552 &  x553 &  x554 &  x557 &  x560 &  x562 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x592 &  x593 &  x596 &  x599 &  x601 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x631 &  x632 &  x635 &  x638 &  x640 &  x641 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x670 &  x671 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x330 & ~x369 & ~x408 & ~x510 & ~x549 & ~x588 & ~x627 & ~x666;
assign c792 =  x26 &  x32 &  x41 &  x50 &  x59 &  x65 &  x68 &  x71 &  x74 &  x83 &  x107 &  x110 &  x113 &  x119 &  x125 &  x128 &  x131 &  x143 &  x146 &  x149 &  x155 &  x161 &  x173 &  x176 &  x182 &  x185 &  x194 &  x197 &  x203 &  x230 &  x236 &  x242 &  x257 &  x266 &  x275 &  x278 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x323 &  x332 &  x338 &  x341 &  x347 &  x350 &  x359 &  x362 &  x365 &  x371 &  x374 &  x380 &  x389 &  x398 &  x401 &  x410 &  x413 &  x419 &  x422 &  x425 &  x431 &  x437 &  x440 &  x446 &  x449 &  x452 &  x455 &  x461 &  x464 &  x467 &  x473 &  x482 &  x485 &  x488 &  x494 &  x503 &  x509 &  x512 &  x515 &  x518 &  x542 &  x551 &  x554 &  x569 &  x572 &  x581 &  x584 &  x587 &  x602 &  x608 &  x611 &  x614 &  x617 &  x623 &  x626 &  x629 &  x632 &  x637 &  x638 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x668 &  x671 &  x674 &  x689 &  x692 &  x695 &  x698 &  x704 &  x716 &  x722 &  x737 &  x743 &  x746 &  x749 &  x752 &  x755 &  x764 &  x767 &  x776 &  x779 &  x785 &  x791 &  x800 &  x806 &  x812 &  x815 &  x820 &  x821 &  x827 &  x830 &  x833 &  x842 &  x854 &  x859 &  x860 &  x863 &  x869 &  x878 &  x881 &  x884 &  x890 &  x893 &  x896 &  x905 &  x908 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x937 &  x944 &  x959 &  x962 &  x968 &  x977 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1015 &  x1016 &  x1022 &  x1025 &  x1043 &  x1046 &  x1053 &  x1054 &  x1058 &  x1061 &  x1070 &  x1073 &  x1082 &  x1092 &  x1093 &  x1097 &  x1100 &  x1103 &  x1109 &  x1118 &  x1121 &  x1124 &  x1126 &  x1127 & ~x579 & ~x882 & ~x960 & ~x1038 & ~x1077 & ~x1083 & ~x1116 & ~x1117 & ~x1122;
assign c794 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x23 &  x25 &  x26 &  x29 &  x32 &  x41 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x64 &  x65 &  x68 &  x71 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x130 &  x131 &  x134 &  x137 &  x140 &  x143 &  x145 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x167 &  x169 &  x170 &  x173 &  x176 &  x182 &  x184 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x208 &  x209 &  x212 &  x215 &  x221 &  x223 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x247 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x272 &  x275 &  x278 &  x281 &  x284 &  x286 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x317 &  x323 &  x325 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x364 &  x365 &  x370 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x403 &  x404 &  x407 &  x409 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x481 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x520 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x554 &  x557 &  x560 &  x566 &  x569 &  x572 &  x575 &  x578 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x617 &  x620 &  x623 &  x626 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x653 &  x656 &  x662 &  x665 &  x668 &  x671 &  x673 &  x674 &  x677 &  x680 &  x683 &  x689 &  x692 &  x695 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x751 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x833 &  x836 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x881 &  x884 &  x890 &  x893 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x959 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x117 & ~x1116;
assign c796 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x148 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x176 &  x182 &  x185 &  x187 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x226 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x359 &  x362 &  x364 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x386 &  x392 &  x398 &  x401 &  x403 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x315 & ~x354 & ~x426 & ~x465 & ~x504 & ~x744 & ~x783 & ~x822 & ~x823 & ~x861 & ~x862 & ~x900 & ~x901;
assign c798 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x130 &  x131 &  x134 &  x137 &  x140 &  x146 &  x149 &  x152 &  x155 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x199 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x238 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x269 &  x272 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x391 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x464 &  x467 &  x469 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x562 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x590 &  x593 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x640 &  x641 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x757 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x844 &  x845 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x883 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x961 &  x962 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x597 & ~x627 & ~x636 & ~x744 & ~x783 & ~x822;
assign c7100 =  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x92 &  x95 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x167 &  x173 &  x176 &  x179 &  x182 &  x185 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x227 &  x230 &  x233 &  x236 &  x239 &  x245 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x290 &  x293 &  x296 &  x299 &  x302 &  x308 &  x314 &  x317 &  x320 &  x326 &  x329 &  x332 &  x335 &  x338 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x401 &  x403 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x461 &  x470 &  x479 &  x482 &  x485 &  x488 &  x494 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x524 &  x527 &  x530 &  x533 &  x539 &  x541 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x575 &  x578 &  x580 &  x584 &  x587 &  x590 &  x593 &  x596 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x644 &  x647 &  x656 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x697 &  x701 &  x707 &  x710 &  x713 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x736 &  x737 &  x743 &  x746 &  x764 &  x767 &  x770 &  x773 &  x776 &  x782 &  x785 &  x791 &  x794 &  x797 &  x800 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x833 &  x836 &  x839 &  x842 &  x845 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x884 &  x887 &  x893 &  x896 &  x902 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x941 &  x944 &  x947 &  x950 &  x952 &  x953 &  x956 &  x962 &  x968 &  x971 &  x974 &  x977 &  x986 &  x995 &  x1001 &  x1004 &  x1019 &  x1022 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1121 &  x1124 &  x1127 &  x1130 & ~x531 & ~x570 & ~x603 & ~x642 & ~x681 & ~x720 & ~x765 & ~x1017;
assign c7102 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x26 &  x29 &  x38 &  x41 &  x44 &  x50 &  x53 &  x56 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x127 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x157 &  x158 &  x173 &  x176 &  x185 &  x188 &  x191 &  x197 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x233 &  x236 &  x242 &  x245 &  x248 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x274 &  x278 &  x281 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x314 &  x317 &  x320 &  x323 &  x326 &  x332 &  x335 &  x347 &  x352 &  x353 &  x362 &  x365 &  x371 &  x380 &  x386 &  x389 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x452 &  x455 &  x458 &  x464 &  x467 &  x470 &  x475 &  x479 &  x482 &  x491 &  x497 &  x503 &  x506 &  x509 &  x521 &  x524 &  x527 &  x533 &  x539 &  x542 &  x548 &  x551 &  x553 &  x562 &  x572 &  x578 &  x581 &  x593 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x641 &  x647 &  x650 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x683 &  x701 &  x704 &  x707 &  x713 &  x716 &  x722 &  x725 &  x728 &  x737 &  x743 &  x749 &  x752 &  x755 &  x761 &  x770 &  x773 &  x776 &  x779 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x806 &  x809 &  x812 &  x818 &  x821 &  x830 &  x836 &  x842 &  x845 &  x851 &  x857 &  x863 &  x866 &  x869 &  x872 &  x878 &  x884 &  x887 &  x893 &  x899 &  x902 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x992 &  x998 &  x1010 &  x1013 &  x1022 &  x1028 &  x1034 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1061 &  x1064 &  x1070 &  x1079 &  x1088 &  x1091 &  x1094 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x219 & ~x258 & ~x259 & ~x297 & ~x298 & ~x330 & ~x510 & ~x511 & ~x549 & ~x588 & ~x627 & ~x744;
assign c7104 =  x8 &  x11 &  x26 &  x38 &  x56 &  x74 &  x80 &  x104 &  x122 &  x131 &  x137 &  x146 &  x155 &  x164 &  x170 &  x176 &  x188 &  x203 &  x242 &  x269 &  x278 &  x287 &  x296 &  x317 &  x323 &  x353 &  x365 &  x371 &  x377 &  x389 &  x401 &  x404 &  x407 &  x419 &  x422 &  x425 &  x428 &  x478 &  x497 &  x512 &  x536 &  x539 &  x542 &  x557 &  x602 &  x641 &  x653 &  x656 &  x674 &  x686 &  x713 &  x716 &  x743 &  x767 &  x794 &  x797 &  x821 &  x833 &  x848 &  x857 &  x892 &  x896 &  x899 &  x938 &  x953 &  x974 &  x980 &  x1004 &  x1016 &  x1019 &  x1028 &  x1061 &  x1076 &  x1087 &  x1097 &  x1121 & ~x195 & ~x234 & ~x315 & ~x354 & ~x861 & ~x901 & ~x939;
assign c7106 =  x2 &  x5 &  x8 &  x11 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x53 &  x56 &  x59 &  x65 &  x68 &  x77 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x116 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x143 &  x149 &  x167 &  x170 &  x176 &  x179 &  x182 &  x185 &  x188 &  x194 &  x197 &  x200 &  x206 &  x209 &  x215 &  x218 &  x221 &  x224 &  x233 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x266 &  x269 &  x272 &  x278 &  x284 &  x287 &  x290 &  x293 &  x296 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x338 &  x344 &  x347 &  x350 &  x353 &  x359 &  x362 &  x365 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x395 &  x398 &  x407 &  x410 &  x413 &  x416 &  x422 &  x428 &  x431 &  x434 &  x437 &  x443 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x488 &  x491 &  x494 &  x497 &  x500 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x554 &  x557 &  x560 &  x563 &  x569 &  x572 &  x578 &  x581 &  x587 &  x593 &  x596 &  x599 &  x605 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x635 &  x638 &  x641 &  x644 &  x647 &  x653 &  x659 &  x662 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x719 &  x722 &  x725 &  x728 &  x731 &  x740 &  x743 &  x746 &  x749 &  x752 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x779 &  x782 &  x785 &  x788 &  x794 &  x797 &  x800 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x863 &  x866 &  x869 &  x872 &  x878 &  x881 &  x890 &  x893 &  x896 &  x899 &  x905 &  x908 &  x914 &  x920 &  x923 &  x929 &  x932 &  x935 &  x937 &  x938 &  x941 &  x944 &  x947 &  x956 &  x958 &  x959 &  x962 &  x965 &  x968 &  x970 &  x971 &  x974 &  x977 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1010 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1034 &  x1040 &  x1043 &  x1046 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1130 & ~x687 & ~x726 & ~x727 & ~x766 & ~x804 & ~x805 & ~x843 & ~x882 & ~x900 & ~x921 & ~x939 & ~x978 & ~x1017;
assign c7108 =  x5 &  x14 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x65 &  x68 &  x71 &  x74 &  x83 &  x86 &  x95 &  x104 &  x107 &  x110 &  x119 &  x125 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x155 &  x161 &  x167 &  x170 &  x173 &  x179 &  x182 &  x191 &  x197 &  x203 &  x206 &  x215 &  x218 &  x221 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x286 &  x287 &  x290 &  x293 &  x299 &  x305 &  x308 &  x311 &  x323 &  x325 &  x326 &  x332 &  x335 &  x347 &  x350 &  x356 &  x359 &  x365 &  x371 &  x374 &  x377 &  x392 &  x395 &  x398 &  x407 &  x416 &  x431 &  x437 &  x440 &  x446 &  x452 &  x455 &  x458 &  x464 &  x467 &  x473 &  x479 &  x485 &  x488 &  x491 &  x497 &  x500 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x530 &  x533 &  x539 &  x542 &  x545 &  x548 &  x551 &  x557 &  x560 &  x566 &  x569 &  x572 &  x578 &  x584 &  x594 &  x595 &  x599 &  x602 &  x605 &  x608 &  x614 &  x617 &  x623 &  x625 &  x635 &  x647 &  x650 &  x653 &  x656 &  x664 &  x665 &  x674 &  x680 &  x689 &  x692 &  x698 &  x704 &  x707 &  x710 &  x719 &  x722 &  x725 &  x728 &  x737 &  x740 &  x743 &  x746 &  x752 &  x755 &  x767 &  x770 &  x779 &  x782 &  x785 &  x788 &  x791 &  x797 &  x800 &  x809 &  x815 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x854 &  x857 &  x860 &  x863 &  x875 &  x878 &  x884 &  x896 &  x899 &  x902 &  x905 &  x911 &  x926 &  x929 &  x932 &  x935 &  x938 &  x944 &  x953 &  x959 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x1001 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1034 &  x1040 &  x1043 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1091 &  x1097 &  x1100 &  x1103 &  x1115 &  x1118 &  x1121 &  x1127 & ~x315 & ~x354 & ~x432 & ~x471 & ~x552 & ~x669 & ~x939;
assign c7110 =  x11 &  x14 &  x17 &  x26 &  x29 &  x35 &  x38 &  x41 &  x47 &  x49 &  x50 &  x53 &  x56 &  x59 &  x62 &  x77 &  x79 &  x80 &  x88 &  x95 &  x98 &  x107 &  x110 &  x113 &  x118 &  x119 &  x122 &  x128 &  x137 &  x143 &  x149 &  x155 &  x157 &  x160 &  x167 &  x170 &  x182 &  x188 &  x196 &  x197 &  x200 &  x212 &  x221 &  x227 &  x230 &  x235 &  x236 &  x239 &  x242 &  x251 &  x254 &  x260 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x293 &  x296 &  x299 &  x308 &  x313 &  x314 &  x326 &  x338 &  x341 &  x344 &  x356 &  x362 &  x365 &  x368 &  x374 &  x383 &  x386 &  x392 &  x398 &  x407 &  x413 &  x428 &  x437 &  x443 &  x455 &  x463 &  x464 &  x470 &  x473 &  x479 &  x482 &  x500 &  x503 &  x512 &  x515 &  x521 &  x527 &  x530 &  x536 &  x548 &  x551 &  x554 &  x557 &  x563 &  x572 &  x593 &  x596 &  x602 &  x605 &  x608 &  x614 &  x617 &  x620 &  x632 &  x638 &  x641 &  x644 &  x650 &  x653 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x683 &  x689 &  x698 &  x701 &  x707 &  x710 &  x713 &  x716 &  x719 &  x725 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x748 &  x755 &  x758 &  x761 &  x773 &  x776 &  x785 &  x788 &  x794 &  x797 &  x806 &  x809 &  x815 &  x824 &  x826 &  x833 &  x836 &  x842 &  x844 &  x848 &  x854 &  x860 &  x866 &  x869 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x896 &  x905 &  x908 &  x916 &  x920 &  x923 &  x929 &  x932 &  x941 &  x944 &  x950 &  x956 &  x965 &  x968 &  x980 &  x986 &  x989 &  x995 &  x1001 &  x1004 &  x1007 &  x1016 &  x1025 &  x1028 &  x1037 &  x1043 &  x1049 &  x1052 &  x1064 &  x1076 &  x1085 &  x1088 &  x1091 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 & ~x84 & ~x123 & ~x162 & ~x375 & ~x393 & ~x432 & ~x433 & ~x472 & ~x511 & ~x549 & ~x627;
assign c7112 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x130 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x169 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x196 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x235 &  x236 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x274 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x391 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x469 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x541 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x580 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x971 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x258 & ~x297 & ~x336 & ~x510 & ~x549 & ~x550 & ~x588 & ~x589 & ~x627 & ~x628 & ~x666 & ~x667 & ~x705 & ~x780 & ~x858 & ~x897 & ~x936 & ~x975 & ~x1092;
assign c7114 =  x2 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x98 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x131 &  x134 &  x137 &  x140 &  x145 &  x152 &  x155 &  x158 &  x161 &  x167 &  x179 &  x182 &  x188 &  x191 &  x194 &  x197 &  x200 &  x209 &  x212 &  x215 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x272 &  x275 &  x281 &  x284 &  x293 &  x296 &  x299 &  x302 &  x308 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x380 &  x386 &  x389 &  x392 &  x395 &  x398 &  x400 &  x410 &  x413 &  x422 &  x425 &  x428 &  x431 &  x434 &  x439 &  x440 &  x443 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x473 &  x476 &  x482 &  x485 &  x494 &  x500 &  x503 &  x506 &  x512 &  x518 &  x521 &  x524 &  x530 &  x536 &  x539 &  x542 &  x545 &  x548 &  x554 &  x557 &  x560 &  x566 &  x575 &  x578 &  x581 &  x584 &  x590 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x625 &  x626 &  x629 &  x635 &  x638 &  x647 &  x650 &  x653 &  x656 &  x659 &  x668 &  x671 &  x674 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x701 &  x703 &  x704 &  x710 &  x713 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x740 &  x742 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x785 &  x788 &  x791 &  x800 &  x803 &  x806 &  x812 &  x815 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x875 &  x887 &  x890 &  x893 &  x899 &  x905 &  x911 &  x914 &  x917 &  x920 &  x923 &  x929 &  x935 &  x938 &  x941 &  x944 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x977 &  x980 &  x983 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1025 &  x1028 &  x1031 &  x1034 &  x1046 &  x1049 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x474 & ~x792 & ~x822 & ~x831 & ~x861 & ~x862 & ~x870 & ~x901 & ~x939 & ~x948 & ~x978 & ~x1065;
assign c7116 =  x13 &  x23 &  x32 &  x35 &  x48 &  x49 &  x50 &  x53 &  x56 &  x65 &  x68 &  x71 &  x74 &  x79 &  x83 &  x88 &  x95 &  x101 &  x113 &  x118 &  x125 &  x131 &  x152 &  x155 &  x164 &  x179 &  x188 &  x191 &  x194 &  x195 &  x200 &  x203 &  x209 &  x215 &  x224 &  x227 &  x230 &  x245 &  x248 &  x254 &  x263 &  x269 &  x293 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x317 &  x320 &  x323 &  x335 &  x338 &  x341 &  x350 &  x371 &  x389 &  x398 &  x407 &  x419 &  x428 &  x443 &  x449 &  x458 &  x461 &  x467 &  x479 &  x488 &  x500 &  x518 &  x521 &  x530 &  x536 &  x545 &  x548 &  x551 &  x560 &  x569 &  x575 &  x578 &  x587 &  x590 &  x593 &  x614 &  x623 &  x626 &  x638 &  x653 &  x659 &  x665 &  x668 &  x683 &  x686 &  x689 &  x692 &  x704 &  x719 &  x722 &  x734 &  x737 &  x743 &  x746 &  x755 &  x770 &  x773 &  x776 &  x779 &  x797 &  x800 &  x803 &  x806 &  x815 &  x824 &  x827 &  x833 &  x845 &  x851 &  x854 &  x857 &  x860 &  x881 &  x896 &  x914 &  x920 &  x932 &  x944 &  x950 &  x956 &  x959 &  x962 &  x980 &  x983 &  x986 &  x1004 &  x1010 &  x1013 &  x1019 &  x1034 &  x1043 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1082 &  x1088 &  x1091 &  x1097 &  x1109 & ~x123 & ~x162 & ~x471 & ~x472 & ~x511 & ~x819;
assign c7118 =  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x47 &  x50 &  x59 &  x62 &  x65 &  x68 &  x71 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x125 &  x130 &  x131 &  x134 &  x137 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x167 &  x169 &  x176 &  x182 &  x185 &  x188 &  x194 &  x197 &  x200 &  x203 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x266 &  x269 &  x274 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x305 &  x308 &  x311 &  x313 &  x317 &  x320 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x352 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x380 &  x383 &  x386 &  x389 &  x391 &  x392 &  x395 &  x398 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x430 &  x431 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x464 &  x467 &  x469 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x494 &  x500 &  x503 &  x506 &  x509 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x547 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x611 &  x617 &  x623 &  x626 &  x629 &  x635 &  x644 &  x653 &  x656 &  x658 &  x659 &  x662 &  x665 &  x668 &  x671 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x749 &  x752 &  x755 &  x758 &  x761 &  x767 &  x770 &  x776 &  x782 &  x785 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x821 &  x824 &  x827 &  x836 &  x842 &  x848 &  x854 &  x857 &  x860 &  x866 &  x869 &  x875 &  x878 &  x887 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x986 &  x989 &  x992 &  x995 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x279 & ~x336 & ~x375 & ~x588 & ~x666 & ~x705 & ~x706 & ~x741 & ~x819;
assign c7120 =  x5 &  x8 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x52 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x83 &  x89 &  x91 &  x92 &  x101 &  x104 &  x107 &  x110 &  x116 &  x119 &  x122 &  x125 &  x131 &  x140 &  x143 &  x149 &  x152 &  x155 &  x158 &  x164 &  x167 &  x170 &  x173 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x196 &  x197 &  x203 &  x206 &  x209 &  x212 &  x218 &  x230 &  x236 &  x239 &  x242 &  x248 &  x251 &  x260 &  x263 &  x266 &  x269 &  x278 &  x284 &  x287 &  x290 &  x293 &  x299 &  x302 &  x305 &  x308 &  x313 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x344 &  x347 &  x350 &  x352 &  x353 &  x356 &  x359 &  x362 &  x368 &  x371 &  x374 &  x377 &  x383 &  x386 &  x389 &  x391 &  x395 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x430 &  x431 &  x434 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x500 &  x503 &  x506 &  x509 &  x514 &  x515 &  x521 &  x524 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x553 &  x554 &  x557 &  x560 &  x563 &  x566 &  x572 &  x575 &  x578 &  x581 &  x584 &  x590 &  x593 &  x596 &  x599 &  x605 &  x611 &  x614 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x695 &  x698 &  x704 &  x707 &  x710 &  x719 &  x722 &  x725 &  x731 &  x734 &  x737 &  x740 &  x746 &  x749 &  x752 &  x755 &  x761 &  x764 &  x767 &  x773 &  x776 &  x779 &  x785 &  x788 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x875 &  x881 &  x884 &  x887 &  x893 &  x902 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x258 & ~x408 & ~x510 & ~x549 & ~x550 & ~x588 & ~x589 & ~x627 & ~x663 & ~x702 & ~x705 & ~x741 & ~x819 & ~x858;
assign c7122 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x26 &  x29 &  x32 &  x35 &  x41 &  x44 &  x47 &  x50 &  x53 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x83 &  x95 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x149 &  x152 &  x161 &  x164 &  x170 &  x173 &  x179 &  x182 &  x188 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x275 &  x278 &  x281 &  x284 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x314 &  x317 &  x320 &  x323 &  x326 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x362 &  x365 &  x371 &  x374 &  x377 &  x383 &  x386 &  x389 &  x395 &  x398 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x431 &  x434 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x520 &  x524 &  x527 &  x530 &  x533 &  x536 &  x545 &  x548 &  x551 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x719 &  x731 &  x734 &  x737 &  x743 &  x746 &  x749 &  x752 &  x755 &  x757 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x788 &  x791 &  x796 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x893 &  x896 &  x899 &  x902 &  x905 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x938 &  x941 &  x947 &  x950 &  x953 &  x956 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1013 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1127 &  x1130 & ~x120 & ~x198 & ~x237 & ~x276 & ~x315 & ~x435 & ~x765 & ~x861 & ~x900 & ~x901 & ~x940 & ~x978 & ~x1017 & ~x1056;
assign c7124 =  x8 &  x14 &  x20 &  x26 &  x29 &  x38 &  x44 &  x47 &  x56 &  x77 &  x80 &  x92 &  x95 &  x98 &  x134 &  x137 &  x152 &  x197 &  x200 &  x206 &  x227 &  x230 &  x239 &  x251 &  x254 &  x259 &  x260 &  x263 &  x269 &  x290 &  x293 &  x296 &  x305 &  x311 &  x323 &  x332 &  x343 &  x359 &  x362 &  x370 &  x374 &  x377 &  x380 &  x382 &  x392 &  x395 &  x406 &  x410 &  x413 &  x428 &  x434 &  x448 &  x464 &  x467 &  x479 &  x485 &  x487 &  x491 &  x497 &  x500 &  x506 &  x512 &  x515 &  x521 &  x533 &  x536 &  x548 &  x557 &  x569 &  x572 &  x581 &  x584 &  x587 &  x593 &  x596 &  x605 &  x611 &  x614 &  x634 &  x644 &  x650 &  x656 &  x659 &  x668 &  x680 &  x686 &  x689 &  x698 &  x712 &  x716 &  x728 &  x734 &  x740 &  x743 &  x746 &  x750 &  x758 &  x779 &  x782 &  x785 &  x791 &  x794 &  x800 &  x806 &  x809 &  x818 &  x819 &  x827 &  x836 &  x839 &  x859 &  x863 &  x866 &  x869 &  x872 &  x884 &  x898 &  x899 &  x902 &  x905 &  x917 &  x929 &  x935 &  x937 &  x953 &  x962 &  x968 &  x974 &  x976 &  x977 &  x980 &  x1001 &  x1025 &  x1031 &  x1034 &  x1037 &  x1061 &  x1064 &  x1067 &  x1079 &  x1088 &  x1118 &  x1124 &  x1130;
assign c7126 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x904 &  x905 &  x908 &  x911 &  x914 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x982 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1020 &  x1021 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1060 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1099 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x99 & ~x138 & ~x189 & ~x228 & ~x267 & ~x345 & ~x900 & ~x939 & ~x978 & ~x1017;
assign c7128 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x59 &  x62 &  x68 &  x71 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x302 &  x305 &  x308 &  x311 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x403 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x481 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x608 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x637 &  x638 &  x641 &  x644 &  x650 &  x653 &  x659 &  x662 &  x664 &  x665 &  x668 &  x671 &  x674 &  x676 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x703 &  x707 &  x710 &  x713 &  x715 &  x716 &  x719 &  x722 &  x725 &  x728 &  x734 &  x737 &  x740 &  x742 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x827 &  x830 &  x833 &  x835 &  x842 &  x845 &  x848 &  x851 &  x854 &  x860 &  x863 &  x865 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x902 &  x904 &  x905 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x938 &  x941 &  x943 &  x944 &  x947 &  x950 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1121 &  x1124 &  x1130 & ~x609 & ~x648 & ~x687 & ~x726 & ~x861 & ~x939 & ~x978;
assign c7130 =  x2 &  x8 &  x11 &  x17 &  x20 &  x23 &  x35 &  x41 &  x53 &  x59 &  x62 &  x65 &  x74 &  x77 &  x83 &  x92 &  x104 &  x107 &  x116 &  x119 &  x131 &  x140 &  x149 &  x155 &  x158 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x191 &  x194 &  x197 &  x200 &  x203 &  x212 &  x224 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x265 &  x266 &  x269 &  x281 &  x284 &  x290 &  x293 &  x296 &  x299 &  x302 &  x304 &  x308 &  x311 &  x314 &  x326 &  x329 &  x332 &  x335 &  x338 &  x344 &  x347 &  x353 &  x356 &  x368 &  x371 &  x374 &  x377 &  x383 &  x392 &  x401 &  x410 &  x413 &  x419 &  x422 &  x428 &  x443 &  x449 &  x452 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x500 &  x503 &  x518 &  x527 &  x530 &  x533 &  x548 &  x554 &  x557 &  x559 &  x560 &  x563 &  x578 &  x581 &  x584 &  x587 &  x593 &  x596 &  x602 &  x605 &  x608 &  x617 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x650 &  x656 &  x664 &  x677 &  x695 &  x698 &  x701 &  x703 &  x704 &  x707 &  x710 &  x713 &  x719 &  x725 &  x728 &  x734 &  x737 &  x742 &  x746 &  x752 &  x758 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x791 &  x794 &  x797 &  x803 &  x818 &  x820 &  x821 &  x830 &  x836 &  x842 &  x854 &  x860 &  x869 &  x872 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x923 &  x932 &  x935 &  x947 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x983 &  x989 &  x998 &  x1004 &  x1019 &  x1022 &  x1025 &  x1031 &  x1037 &  x1049 &  x1058 &  x1061 &  x1064 &  x1067 &  x1079 &  x1082 &  x1091 &  x1094 &  x1106 &  x1112 &  x1121 &  x1124 &  x1127 &  x1130 & ~x315 & ~x354 & ~x393 & ~x432 & ~x471 & ~x606 & ~x630 & ~x645 & ~x939 & ~x960 & ~x978 & ~x1017 & ~x1056 & ~x1095;
assign c7132 =  x2 &  x11 &  x17 &  x23 &  x26 &  x41 &  x44 &  x47 &  x53 &  x59 &  x62 &  x65 &  x68 &  x74 &  x77 &  x89 &  x92 &  x98 &  x101 &  x107 &  x113 &  x119 &  x122 &  x125 &  x128 &  x134 &  x140 &  x152 &  x158 &  x161 &  x167 &  x170 &  x188 &  x194 &  x203 &  x212 &  x215 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x251 &  x254 &  x260 &  x263 &  x272 &  x278 &  x284 &  x287 &  x296 &  x314 &  x317 &  x323 &  x326 &  x332 &  x335 &  x338 &  x344 &  x347 &  x359 &  x371 &  x377 &  x380 &  x386 &  x392 &  x395 &  x398 &  x401 &  x404 &  x410 &  x416 &  x422 &  x425 &  x431 &  x434 &  x437 &  x440 &  x443 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x473 &  x479 &  x485 &  x488 &  x491 &  x506 &  x509 &  x515 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x548 &  x557 &  x560 &  x566 &  x578 &  x584 &  x599 &  x605 &  x629 &  x632 &  x635 &  x644 &  x647 &  x653 &  x659 &  x668 &  x671 &  x680 &  x683 &  x686 &  x692 &  x710 &  x713 &  x716 &  x719 &  x722 &  x731 &  x737 &  x743 &  x746 &  x752 &  x770 &  x776 &  x779 &  x785 &  x788 &  x797 &  x800 &  x803 &  x820 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x842 &  x848 &  x851 &  x854 &  x857 &  x859 &  x860 &  x863 &  x872 &  x875 &  x878 &  x884 &  x893 &  x896 &  x898 &  x902 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x931 &  x938 &  x941 &  x952 &  x953 &  x956 &  x962 &  x965 &  x968 &  x970 &  x976 &  x977 &  x989 &  x997 &  x1015 &  x1016 &  x1019 &  x1030 &  x1031 &  x1036 &  x1037 &  x1040 &  x1043 &  x1046 &  x1054 &  x1055 &  x1064 &  x1069 &  x1073 &  x1076 &  x1082 &  x1091 &  x1093 &  x1094 &  x1100 &  x1106 &  x1112 &  x1115 &  x1118 &  x1124 &  x1130 & ~x837 & ~x876 & ~x915 & ~x916 & ~x921 & ~x960 & ~x978 & ~x1032 & ~x1071;
assign c7134 =  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x179 &  x182 &  x191 &  x194 &  x197 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x320 &  x323 &  x326 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x592 &  x593 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x631 &  x632 &  x635 &  x640 &  x641 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x670 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x691 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x746 &  x748 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x803 &  x806 &  x809 &  x812 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x953 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x369 & ~x414 & ~x453 & ~x492 & ~x531 & ~x555 & ~x594 & ~x624 & ~x633 & ~x663 & ~x672 & ~x702 & ~x711 & ~x741 & ~x750 & ~x780 & ~x819 & ~x858 & ~x897;
assign c7136 =  x11 &  x14 &  x20 &  x22 &  x32 &  x34 &  x50 &  x53 &  x61 &  x62 &  x65 &  x74 &  x77 &  x92 &  x107 &  x119 &  x137 &  x146 &  x149 &  x152 &  x161 &  x173 &  x211 &  x218 &  x221 &  x224 &  x227 &  x236 &  x250 &  x251 &  x254 &  x260 &  x263 &  x266 &  x268 &  x287 &  x290 &  x293 &  x299 &  x307 &  x317 &  x329 &  x353 &  x359 &  x362 &  x365 &  x371 &  x383 &  x410 &  x412 &  x413 &  x431 &  x440 &  x443 &  x445 &  x446 &  x455 &  x458 &  x461 &  x464 &  x485 &  x488 &  x491 &  x500 &  x509 &  x518 &  x527 &  x536 &  x539 &  x554 &  x557 &  x575 &  x581 &  x584 &  x587 &  x593 &  x595 &  x634 &  x638 &  x647 &  x659 &  x662 &  x671 &  x674 &  x677 &  x698 &  x710 &  x713 &  x715 &  x716 &  x719 &  x725 &  x740 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x781 &  x794 &  x812 &  x818 &  x824 &  x839 &  x848 &  x851 &  x860 &  x866 &  x872 &  x881 &  x892 &  x920 &  x926 &  x931 &  x935 &  x970 &  x971 &  x975 &  x983 &  x992 &  x998 &  x1007 &  x1014 &  x1019 &  x1028 &  x1031 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1073 &  x1076 &  x1085 &  x1091 &  x1106 & ~x354 & ~x393 & ~x1128;
assign c7138 =  x5 &  x11 &  x23 &  x41 &  x43 &  x47 &  x62 &  x65 &  x68 &  x71 &  x77 &  x79 &  x86 &  x89 &  x92 &  x104 &  x110 &  x113 &  x116 &  x118 &  x119 &  x122 &  x137 &  x158 &  x164 &  x170 &  x182 &  x194 &  x197 &  x203 &  x218 &  x239 &  x242 &  x245 &  x248 &  x250 &  x254 &  x257 &  x260 &  x269 &  x281 &  x284 &  x287 &  x289 &  x302 &  x305 &  x326 &  x329 &  x340 &  x350 &  x356 &  x359 &  x367 &  x371 &  x374 &  x380 &  x383 &  x386 &  x389 &  x395 &  x407 &  x416 &  x428 &  x437 &  x446 &  x449 &  x452 &  x455 &  x458 &  x470 &  x479 &  x482 &  x485 &  x491 &  x506 &  x509 &  x518 &  x524 &  x533 &  x536 &  x539 &  x548 &  x551 &  x562 &  x563 &  x575 &  x593 &  x608 &  x614 &  x623 &  x629 &  x635 &  x659 &  x665 &  x668 &  x671 &  x677 &  x683 &  x698 &  x701 &  x713 &  x722 &  x728 &  x737 &  x746 &  x752 &  x755 &  x758 &  x761 &  x767 &  x770 &  x773 &  x776 &  x782 &  x785 &  x788 &  x791 &  x794 &  x803 &  x806 &  x809 &  x815 &  x818 &  x824 &  x827 &  x830 &  x833 &  x839 &  x851 &  x866 &  x869 &  x872 &  x881 &  x887 &  x893 &  x902 &  x908 &  x911 &  x920 &  x926 &  x935 &  x941 &  x947 &  x953 &  x959 &  x962 &  x970 &  x971 &  x977 &  x983 &  x986 &  x997 &  x1004 &  x1013 &  x1025 &  x1028 &  x1034 &  x1037 &  x1040 &  x1049 &  x1064 &  x1073 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 & ~x1017 & ~x1018 & ~x1056;
assign c7140 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x929 &  x932 &  x938 &  x941 &  x947 &  x950 &  x953 &  x956 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x998 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130 & ~x15 & ~x27 & ~x54 & ~x66 & ~x93 & ~x99 & ~x105 & ~x144 & ~x183 & ~x189 & ~x411 & ~x531 & ~x570 & ~x783 & ~x822 & ~x861 & ~x867 & ~x900 & ~x906 & ~x945 & ~x978 & ~x984 & ~x1023 & ~x1062 & ~x1101;
assign c7142 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x65 &  x71 &  x74 &  x80 &  x83 &  x86 &  x89 &  x95 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x380 &  x382 &  x386 &  x389 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x421 &  x422 &  x425 &  x428 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x551 &  x554 &  x557 &  x559 &  x560 &  x563 &  x566 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x598 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x637 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x716 &  x719 &  x722 &  x725 &  x728 &  x734 &  x737 &  x740 &  x742 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x781 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x820 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x859 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x884 &  x890 &  x893 &  x896 &  x898 &  x899 &  x902 &  x905 &  x908 &  x914 &  x920 &  x923 &  x929 &  x932 &  x935 &  x937 &  x938 &  x941 &  x944 &  x947 &  x950 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1015 &  x1016 &  x1019 &  x1022 &  x1025 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1054 &  x1055 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1093 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1130 & ~x315 & ~x354 & ~x390 & ~x393 & ~x432 & ~x471 & ~x939 & ~x978 & ~x1017 & ~x1056 & ~x1104;
assign c7144 =  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x44 &  x47 &  x50 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x80 &  x82 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x113 &  x119 &  x121 &  x122 &  x125 &  x134 &  x137 &  x140 &  x146 &  x155 &  x157 &  x158 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x196 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x218 &  x224 &  x230 &  x233 &  x234 &  x235 &  x239 &  x248 &  x251 &  x257 &  x260 &  x263 &  x266 &  x269 &  x275 &  x278 &  x281 &  x284 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x317 &  x323 &  x326 &  x332 &  x338 &  x341 &  x347 &  x350 &  x352 &  x353 &  x356 &  x359 &  x362 &  x368 &  x371 &  x374 &  x377 &  x380 &  x389 &  x392 &  x395 &  x398 &  x401 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x430 &  x431 &  x434 &  x437 &  x440 &  x449 &  x455 &  x458 &  x461 &  x464 &  x469 &  x470 &  x473 &  x475 &  x476 &  x484 &  x485 &  x488 &  x491 &  x494 &  x500 &  x506 &  x509 &  x514 &  x515 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x542 &  x545 &  x548 &  x553 &  x557 &  x562 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x605 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x653 &  x656 &  x659 &  x665 &  x671 &  x674 &  x677 &  x680 &  x686 &  x692 &  x695 &  x701 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x758 &  x761 &  x764 &  x767 &  x773 &  x776 &  x779 &  x782 &  x788 &  x791 &  x794 &  x800 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x902 &  x911 &  x914 &  x917 &  x920 &  x926 &  x929 &  x932 &  x935 &  x944 &  x947 &  x950 &  x953 &  x962 &  x965 &  x968 &  x974 &  x977 &  x980 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1058 &  x1061 &  x1064 &  x1070 &  x1079 &  x1082 &  x1088 &  x1091 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x114 & ~x162 & ~x219 & ~x297 & ~x432 & ~x471 & ~x510 & ~x519;
assign c7146 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x62 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x89 &  x91 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x130 &  x131 &  x137 &  x140 &  x143 &  x146 &  x149 &  x155 &  x158 &  x161 &  x164 &  x167 &  x169 &  x170 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x208 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x244 &  x245 &  x247 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x380 &  x383 &  x386 &  x389 &  x391 &  x392 &  x395 &  x401 &  x404 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x430 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x458 &  x464 &  x469 &  x470 &  x473 &  x476 &  x479 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x508 &  x512 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x587 &  x593 &  x596 &  x599 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x710 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x740 &  x743 &  x746 &  x749 &  x752 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x785 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x941 &  x944 &  x947 &  x950 &  x953 &  x959 &  x962 &  x965 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x315 & ~x706 & ~x783 & ~x822 & ~x861 & ~x939;
assign c7148 =  x5 &  x8 &  x11 &  x14 &  x17 &  x23 &  x26 &  x29 &  x32 &  x35 &  x41 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x91 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x113 &  x116 &  x119 &  x122 &  x128 &  x131 &  x134 &  x137 &  x140 &  x146 &  x152 &  x155 &  x158 &  x161 &  x164 &  x170 &  x173 &  x176 &  x179 &  x182 &  x188 &  x191 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x248 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x281 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x383 &  x386 &  x389 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x503 &  x506 &  x509 &  x512 &  x514 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x562 &  x563 &  x566 &  x569 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x629 &  x632 &  x635 &  x638 &  x640 &  x641 &  x644 &  x650 &  x653 &  x656 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x752 &  x755 &  x758 &  x761 &  x764 &  x770 &  x773 &  x776 &  x779 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x928 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x956 &  x959 &  x962 &  x965 &  x967 &  x968 &  x974 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1006 &  x1007 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x330 & ~x369 & ~x408 & ~x471 & ~x511 & ~x549 & ~x550 & ~x588 & ~x589 & ~x627 & ~x628 & ~x666 & ~x705 & ~x744 & ~x783;
assign c7150 =  x2 &  x5 &  x26 &  x29 &  x32 &  x41 &  x44 &  x47 &  x53 &  x62 &  x65 &  x68 &  x71 &  x77 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x122 &  x125 &  x134 &  x137 &  x140 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x176 &  x179 &  x185 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x224 &  x230 &  x236 &  x242 &  x245 &  x248 &  x257 &  x269 &  x272 &  x275 &  x278 &  x293 &  x296 &  x302 &  x305 &  x308 &  x320 &  x323 &  x335 &  x338 &  x341 &  x347 &  x353 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x383 &  x392 &  x398 &  x401 &  x404 &  x407 &  x416 &  x419 &  x434 &  x437 &  x440 &  x443 &  x455 &  x464 &  x467 &  x470 &  x473 &  x476 &  x485 &  x488 &  x491 &  x494 &  x497 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x533 &  x542 &  x545 &  x551 &  x557 &  x559 &  x560 &  x566 &  x569 &  x575 &  x581 &  x590 &  x596 &  x598 &  x599 &  x602 &  x611 &  x614 &  x617 &  x620 &  x629 &  x632 &  x635 &  x638 &  x641 &  x647 &  x653 &  x662 &  x665 &  x668 &  x671 &  x677 &  x683 &  x707 &  x728 &  x734 &  x737 &  x742 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x770 &  x776 &  x781 &  x794 &  x797 &  x803 &  x806 &  x820 &  x824 &  x827 &  x836 &  x839 &  x845 &  x848 &  x851 &  x857 &  x860 &  x869 &  x872 &  x875 &  x878 &  x890 &  x898 &  x899 &  x905 &  x908 &  x911 &  x929 &  x932 &  x935 &  x941 &  x947 &  x950 &  x953 &  x956 &  x965 &  x968 &  x971 &  x998 &  x1007 &  x1009 &  x1013 &  x1016 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1049 &  x1055 &  x1067 &  x1073 &  x1079 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1121 & ~x471 & ~x837 & ~x876 & ~x915 & ~x916 & ~x921 & ~x978 & ~x993 & ~x1017 & ~x1032 & ~x1056 & ~x1110 & ~x1111;
assign c7152 =  x5 &  x8 &  x14 &  x17 &  x29 &  x44 &  x50 &  x56 &  x59 &  x62 &  x65 &  x68 &  x74 &  x80 &  x89 &  x98 &  x101 &  x103 &  x104 &  x107 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x130 &  x134 &  x137 &  x143 &  x146 &  x152 &  x155 &  x158 &  x161 &  x164 &  x169 &  x170 &  x173 &  x176 &  x182 &  x191 &  x197 &  x206 &  x209 &  x212 &  x215 &  x224 &  x233 &  x236 &  x242 &  x245 &  x248 &  x254 &  x257 &  x260 &  x266 &  x269 &  x275 &  x278 &  x281 &  x284 &  x287 &  x293 &  x299 &  x305 &  x308 &  x311 &  x320 &  x323 &  x326 &  x332 &  x335 &  x338 &  x341 &  x347 &  x353 &  x362 &  x368 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x488 &  x497 &  x509 &  x512 &  x515 &  x518 &  x521 &  x527 &  x533 &  x536 &  x542 &  x545 &  x548 &  x551 &  x557 &  x560 &  x563 &  x569 &  x572 &  x578 &  x581 &  x584 &  x587 &  x593 &  x599 &  x608 &  x614 &  x617 &  x623 &  x626 &  x629 &  x635 &  x644 &  x646 &  x647 &  x650 &  x656 &  x659 &  x662 &  x665 &  x674 &  x677 &  x679 &  x683 &  x685 &  x689 &  x698 &  x701 &  x704 &  x707 &  x716 &  x718 &  x724 &  x725 &  x728 &  x734 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x757 &  x761 &  x763 &  x764 &  x767 &  x770 &  x773 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x802 &  x803 &  x809 &  x818 &  x821 &  x833 &  x835 &  x836 &  x841 &  x842 &  x845 &  x851 &  x854 &  x857 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x908 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x935 &  x938 &  x944 &  x950 &  x953 &  x956 &  x965 &  x968 &  x971 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1034 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1103 &  x1106 &  x1109 &  x1121 &  x1127 & ~x279 & ~x318 & ~x357 & ~x666 & ~x667 & ~x744 & ~x783 & ~x822;
assign c7154 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x703 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x742 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x796 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x904 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x943 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x237 & ~x276 & ~x354 & ~x393 & ~x471 & ~x510 & ~x549 & ~x726 & ~x900 & ~x939 & ~x940 & ~x978 & ~x979 & ~x1017 & ~x1018 & ~x1056 & ~x1095;
assign c7156 =  x14 &  x23 &  x26 &  x29 &  x41 &  x44 &  x62 &  x68 &  x71 &  x74 &  x83 &  x92 &  x95 &  x104 &  x113 &  x125 &  x131 &  x143 &  x146 &  x149 &  x164 &  x167 &  x170 &  x173 &  x185 &  x188 &  x200 &  x209 &  x212 &  x221 &  x224 &  x227 &  x245 &  x269 &  x275 &  x278 &  x284 &  x299 &  x302 &  x311 &  x323 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x359 &  x368 &  x377 &  x386 &  x398 &  x407 &  x413 &  x416 &  x419 &  x428 &  x434 &  x437 &  x440 &  x446 &  x464 &  x467 &  x473 &  x476 &  x488 &  x491 &  x497 &  x506 &  x515 &  x517 &  x518 &  x533 &  x536 &  x539 &  x545 &  x560 &  x569 &  x596 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x626 &  x638 &  x641 &  x662 &  x665 &  x674 &  x695 &  x698 &  x704 &  x707 &  x713 &  x719 &  x722 &  x725 &  x740 &  x746 &  x752 &  x755 &  x767 &  x770 &  x785 &  x797 &  x830 &  x845 &  x869 &  x884 &  x887 &  x896 &  x902 &  x923 &  x925 &  x935 &  x947 &  x950 &  x959 &  x962 &  x965 &  x968 &  x970 &  x980 &  x1003 &  x1004 &  x1010 &  x1013 &  x1022 &  x1028 &  x1040 &  x1048 &  x1055 &  x1064 &  x1067 &  x1070 &  x1079 &  x1103 &  x1109 &  x1112 &  x1118 &  x1124 &  x1127 &  x1130 & ~x189 & ~x567 & ~x606 & ~x726 & ~x798;
assign c7158 =  x5 &  x8 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x44 &  x50 &  x53 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x137 &  x140 &  x143 &  x146 &  x152 &  x164 &  x167 &  x170 &  x173 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x206 &  x209 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x239 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x284 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x317 &  x323 &  x326 &  x329 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x362 &  x365 &  x368 &  x377 &  x380 &  x389 &  x392 &  x398 &  x401 &  x406 &  x407 &  x410 &  x416 &  x419 &  x422 &  x431 &  x434 &  x437 &  x440 &  x443 &  x445 &  x446 &  x452 &  x455 &  x461 &  x464 &  x467 &  x476 &  x479 &  x484 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x524 &  x527 &  x530 &  x536 &  x542 &  x545 &  x548 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x587 &  x590 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x620 &  x623 &  x625 &  x626 &  x629 &  x632 &  x635 &  x638 &  x644 &  x656 &  x659 &  x662 &  x664 &  x665 &  x668 &  x674 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x703 &  x704 &  x707 &  x710 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x742 &  x743 &  x746 &  x749 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x781 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x815 &  x818 &  x820 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x845 &  x848 &  x851 &  x857 &  x859 &  x860 &  x863 &  x869 &  x872 &  x875 &  x878 &  x884 &  x887 &  x890 &  x896 &  x904 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x938 &  x941 &  x944 &  x947 &  x953 &  x956 &  x958 &  x959 &  x965 &  x968 &  x971 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x997 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130 & ~x276 & ~x354 & ~x861 & ~x940 & ~x978 & ~x1017;
assign c7160 =  x8 &  x20 &  x23 &  x35 &  x47 &  x50 &  x59 &  x62 &  x65 &  x80 &  x86 &  x107 &  x110 &  x113 &  x119 &  x131 &  x140 &  x149 &  x155 &  x167 &  x170 &  x179 &  x188 &  x206 &  x209 &  x224 &  x248 &  x260 &  x263 &  x266 &  x272 &  x275 &  x293 &  x305 &  x332 &  x344 &  x347 &  x359 &  x371 &  x380 &  x383 &  x392 &  x395 &  x404 &  x407 &  x413 &  x416 &  x419 &  x425 &  x443 &  x446 &  x452 &  x458 &  x467 &  x476 &  x485 &  x488 &  x491 &  x500 &  x503 &  x509 &  x515 &  x521 &  x524 &  x539 &  x554 &  x560 &  x575 &  x578 &  x581 &  x587 &  x593 &  x596 &  x602 &  x605 &  x608 &  x626 &  x629 &  x632 &  x635 &  x647 &  x650 &  x656 &  x674 &  x683 &  x692 &  x695 &  x701 &  x743 &  x749 &  x767 &  x791 &  x803 &  x809 &  x812 &  x815 &  x821 &  x827 &  x830 &  x833 &  x842 &  x845 &  x848 &  x851 &  x863 &  x869 &  x875 &  x878 &  x881 &  x884 &  x896 &  x899 &  x911 &  x917 &  x920 &  x923 &  x929 &  x935 &  x938 &  x947 &  x953 &  x968 &  x974 &  x977 &  x983 &  x989 &  x995 &  x998 &  x1004 &  x1007 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1034 &  x1046 &  x1076 &  x1079 &  x1085 &  x1091 &  x1097 &  x1103 &  x1115 &  x1130 & ~x150 & ~x414 & ~x415 & ~x453 & ~x531 & ~x532 & ~x570 & ~x571 & ~x609 & ~x648 & ~x732 & ~x783 & ~x1065;
assign c7162 =  x11 &  x20 &  x23 &  x26 &  x35 &  x38 &  x41 &  x44 &  x47 &  x53 &  x59 &  x62 &  x65 &  x68 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x101 &  x107 &  x110 &  x113 &  x122 &  x125 &  x146 &  x152 &  x155 &  x161 &  x164 &  x170 &  x179 &  x191 &  x209 &  x212 &  x221 &  x236 &  x254 &  x257 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x284 &  x290 &  x293 &  x308 &  x314 &  x320 &  x326 &  x329 &  x338 &  x341 &  x344 &  x350 &  x359 &  x362 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x395 &  x398 &  x404 &  x410 &  x413 &  x422 &  x425 &  x440 &  x443 &  x452 &  x455 &  x461 &  x464 &  x467 &  x470 &  x485 &  x494 &  x497 &  x500 &  x503 &  x509 &  x512 &  x518 &  x527 &  x533 &  x536 &  x548 &  x551 &  x554 &  x557 &  x566 &  x572 &  x578 &  x584 &  x587 &  x593 &  x599 &  x605 &  x608 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x659 &  x662 &  x665 &  x671 &  x683 &  x686 &  x689 &  x698 &  x704 &  x707 &  x710 &  x713 &  x719 &  x728 &  x734 &  x737 &  x740 &  x742 &  x746 &  x749 &  x755 &  x758 &  x761 &  x767 &  x770 &  x773 &  x776 &  x785 &  x788 &  x791 &  x797 &  x803 &  x809 &  x812 &  x815 &  x824 &  x830 &  x833 &  x839 &  x842 &  x845 &  x857 &  x866 &  x872 &  x881 &  x884 &  x893 &  x899 &  x902 &  x923 &  x926 &  x935 &  x944 &  x950 &  x953 &  x959 &  x962 &  x971 &  x986 &  x998 &  x1001 &  x1007 &  x1010 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1043 &  x1052 &  x1055 &  x1060 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1130 & ~x273 & ~x777 & ~x816 & ~x882 & ~x921 & ~x960 & ~x1011 & ~x1017 & ~x1018 & ~x1050 & ~x1089 & ~x1095 & ~x1128;
assign c7164 =  x10 &  x11 &  x14 &  x26 &  x29 &  x32 &  x40 &  x47 &  x49 &  x53 &  x62 &  x65 &  x68 &  x71 &  x74 &  x83 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x117 &  x118 &  x122 &  x131 &  x134 &  x140 &  x143 &  x149 &  x155 &  x156 &  x157 &  x158 &  x164 &  x170 &  x179 &  x185 &  x191 &  x194 &  x196 &  x203 &  x209 &  x212 &  x218 &  x221 &  x233 &  x245 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x274 &  x275 &  x278 &  x281 &  x287 &  x293 &  x296 &  x299 &  x314 &  x317 &  x329 &  x338 &  x341 &  x344 &  x347 &  x356 &  x359 &  x365 &  x368 &  x374 &  x377 &  x380 &  x383 &  x395 &  x401 &  x413 &  x422 &  x428 &  x431 &  x440 &  x443 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x473 &  x476 &  x482 &  x485 &  x488 &  x494 &  x497 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x548 &  x557 &  x560 &  x566 &  x569 &  x575 &  x587 &  x590 &  x593 &  x596 &  x608 &  x617 &  x626 &  x629 &  x632 &  x635 &  x638 &  x647 &  x650 &  x656 &  x671 &  x683 &  x692 &  x698 &  x701 &  x710 &  x713 &  x719 &  x722 &  x734 &  x740 &  x743 &  x749 &  x752 &  x755 &  x760 &  x761 &  x776 &  x785 &  x791 &  x794 &  x797 &  x799 &  x806 &  x815 &  x821 &  x827 &  x839 &  x842 &  x845 &  x863 &  x869 &  x872 &  x875 &  x887 &  x890 &  x893 &  x902 &  x911 &  x920 &  x923 &  x932 &  x944 &  x947 &  x953 &  x956 &  x959 &  x971 &  x980 &  x989 &  x992 &  x1001 &  x1004 &  x1022 &  x1028 &  x1040 &  x1046 &  x1061 &  x1064 &  x1067 &  x1079 &  x1085 &  x1088 &  x1103 &  x1106 &  x1109 &  x1118 &  x1124 &  x1127 & ~x85 & ~x180 & ~x219 & ~x258 & ~x394 & ~x432 & ~x741 & ~x780 & ~x819 & ~x858 & ~x897;
assign c7166 =  x2 &  x5 &  x8 &  x11 &  x17 &  x26 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x89 &  x95 &  x98 &  x104 &  x113 &  x119 &  x125 &  x128 &  x131 &  x134 &  x140 &  x143 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x197 &  x203 &  x206 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x251 &  x254 &  x260 &  x266 &  x272 &  x275 &  x278 &  x281 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x332 &  x335 &  x338 &  x341 &  x344 &  x350 &  x353 &  x356 &  x362 &  x371 &  x374 &  x380 &  x383 &  x386 &  x392 &  x395 &  x398 &  x401 &  x403 &  x404 &  x407 &  x413 &  x416 &  x419 &  x422 &  x431 &  x437 &  x440 &  x442 &  x446 &  x452 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x481 &  x482 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x523 &  x524 &  x527 &  x533 &  x536 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x572 &  x575 &  x581 &  x587 &  x590 &  x593 &  x599 &  x602 &  x605 &  x611 &  x617 &  x620 &  x623 &  x626 &  x632 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x662 &  x665 &  x674 &  x680 &  x683 &  x689 &  x692 &  x698 &  x701 &  x707 &  x713 &  x716 &  x719 &  x725 &  x728 &  x731 &  x734 &  x737 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x794 &  x796 &  x797 &  x806 &  x812 &  x818 &  x824 &  x827 &  x830 &  x833 &  x835 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x874 &  x875 &  x878 &  x881 &  x884 &  x890 &  x893 &  x896 &  x905 &  x908 &  x911 &  x917 &  x923 &  x926 &  x929 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x968 &  x971 &  x974 &  x980 &  x986 &  x992 &  x995 &  x1001 &  x1004 &  x1010 &  x1013 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1052 &  x1055 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x117 & ~x156 & ~x195 & ~x273 & ~x312 & ~x351 & ~x822 & ~x861 & ~x933 & ~x939 & ~x972 & ~x978;
assign c7168 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x23 &  x25 &  x26 &  x29 &  x35 &  x38 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x260 &  x266 &  x269 &  x275 &  x287 &  x290 &  x293 &  x296 &  x299 &  x305 &  x308 &  x314 &  x317 &  x320 &  x326 &  x332 &  x335 &  x338 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x398 &  x404 &  x407 &  x413 &  x416 &  x419 &  x422 &  x425 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x476 &  x479 &  x482 &  x488 &  x491 &  x494 &  x497 &  x500 &  x506 &  x509 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x599 &  x602 &  x608 &  x614 &  x617 &  x620 &  x623 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x674 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x713 &  x716 &  x719 &  x725 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x767 &  x770 &  x773 &  x775 &  x776 &  x779 &  x782 &  x788 &  x791 &  x794 &  x797 &  x800 &  x806 &  x812 &  x815 &  x821 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x863 &  x866 &  x869 &  x875 &  x878 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x914 &  x917 &  x920 &  x923 &  x929 &  x935 &  x950 &  x953 &  x956 &  x959 &  x962 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x1001 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 & ~x216 & ~x222 & ~x294 & ~x333 & ~x672 & ~x726 & ~x819 & ~x906;
assign c7170 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x29 &  x35 &  x38 &  x44 &  x50 &  x56 &  x59 &  x65 &  x71 &  x74 &  x80 &  x83 &  x89 &  x95 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x152 &  x155 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x233 &  x236 &  x239 &  x242 &  x248 &  x254 &  x257 &  x260 &  x265 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x290 &  x293 &  x296 &  x302 &  x304 &  x308 &  x311 &  x317 &  x320 &  x323 &  x329 &  x332 &  x341 &  x343 &  x344 &  x353 &  x356 &  x359 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x395 &  x398 &  x404 &  x410 &  x413 &  x416 &  x419 &  x431 &  x437 &  x440 &  x442 &  x443 &  x446 &  x449 &  x452 &  x455 &  x461 &  x464 &  x467 &  x479 &  x481 &  x482 &  x488 &  x491 &  x500 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x527 &  x533 &  x545 &  x548 &  x554 &  x562 &  x569 &  x575 &  x578 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x601 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x623 &  x626 &  x632 &  x635 &  x638 &  x640 &  x641 &  x644 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x674 &  x677 &  x679 &  x683 &  x686 &  x689 &  x692 &  x698 &  x701 &  x703 &  x707 &  x710 &  x713 &  x716 &  x718 &  x719 &  x722 &  x728 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x757 &  x761 &  x764 &  x767 &  x770 &  x773 &  x781 &  x788 &  x791 &  x796 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x820 &  x821 &  x824 &  x830 &  x833 &  x835 &  x836 &  x848 &  x854 &  x857 &  x859 &  x869 &  x872 &  x874 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x898 &  x899 &  x905 &  x908 &  x911 &  x913 &  x914 &  x920 &  x923 &  x929 &  x935 &  x937 &  x938 &  x941 &  x947 &  x953 &  x956 &  x965 &  x974 &  x989 &  x991 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1070 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x552 & ~x978;
assign c7172 =  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x74 &  x77 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x161 &  x164 &  x167 &  x173 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x218 &  x221 &  x224 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x251 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x292 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x329 &  x331 &  x332 &  x335 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x364 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x437 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x518 &  x524 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x635 &  x638 &  x641 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x703 &  x707 &  x710 &  x713 &  x716 &  x718 &  x719 &  x722 &  x725 &  x734 &  x737 &  x740 &  x743 &  x746 &  x748 &  x749 &  x752 &  x755 &  x757 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x787 &  x788 &  x791 &  x796 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x913 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x952 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x465 & ~x504 & ~x744 & ~x783 & ~x784 & ~x822 & ~x861;
assign c7174 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x52 &  x53 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x91 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x274 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x314 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x629 &  x632 &  x635 &  x638 &  x641 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x844 &  x845 &  x848 &  x851 &  x854 &  x860 &  x863 &  x866 &  x869 &  x872 &  x878 &  x881 &  x883 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x471 & ~x510 & ~x511 & ~x519 & ~x549 & ~x550 & ~x589 & ~x597 & ~x624 & ~x627 & ~x666 & ~x702 & ~x705 & ~x741 & ~x780 & ~x819;
assign c7176 =  x2 &  x5 &  x8 &  x11 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x242 &  x244 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x266 &  x269 &  x272 &  x274 &  x275 &  x278 &  x281 &  x282 &  x283 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x314 &  x317 &  x320 &  x322 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x356 &  x359 &  x361 &  x362 &  x365 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x391 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x430 &  x431 &  x434 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x469 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x508 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x547 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x656 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x333 & ~x372 & ~x411 & ~x519 & ~x627 & ~x666 & ~x667 & ~x705 & ~x706 & ~x744 & ~x783 & ~x822;
assign c7178 =  x5 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x34 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x74 &  x80 &  x83 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x167 &  x170 &  x179 &  x182 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x293 &  x299 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x365 &  x368 &  x371 &  x374 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x437 &  x440 &  x443 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x512 &  x515 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x551 &  x554 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x626 &  x629 &  x632 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x662 &  x664 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x695 &  x698 &  x701 &  x703 &  x704 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x770 &  x773 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x833 &  x836 &  x839 &  x842 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x878 &  x884 &  x887 &  x890 &  x893 &  x896 &  x902 &  x904 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x943 &  x944 &  x947 &  x956 &  x959 &  x962 &  x965 &  x971 &  x974 &  x980 &  x983 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1055 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1085 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1124 &  x1127 & ~x606 & ~x609 & ~x648 & ~x726 & ~x765 & ~x861 & ~x900 & ~x939 & ~x978;
assign c7180 =  x14 &  x23 &  x26 &  x32 &  x38 &  x41 &  x43 &  x50 &  x53 &  x56 &  x59 &  x62 &  x71 &  x74 &  x77 &  x80 &  x95 &  x113 &  x122 &  x128 &  x158 &  x170 &  x176 &  x185 &  x203 &  x206 &  x209 &  x233 &  x242 &  x254 &  x260 &  x266 &  x275 &  x281 &  x308 &  x317 &  x323 &  x326 &  x329 &  x332 &  x344 &  x347 &  x350 &  x367 &  x377 &  x392 &  x398 &  x404 &  x410 &  x416 &  x428 &  x434 &  x437 &  x440 &  x444 &  x446 &  x455 &  x470 &  x473 &  x476 &  x479 &  x483 &  x485 &  x497 &  x500 &  x506 &  x515 &  x518 &  x521 &  x522 &  x539 &  x545 &  x551 &  x554 &  x581 &  x584 &  x587 &  x590 &  x600 &  x608 &  x620 &  x623 &  x626 &  x629 &  x638 &  x680 &  x686 &  x707 &  x725 &  x728 &  x743 &  x746 &  x749 &  x752 &  x761 &  x770 &  x776 &  x788 &  x791 &  x797 &  x809 &  x818 &  x833 &  x836 &  x842 &  x845 &  x848 &  x851 &  x854 &  x863 &  x878 &  x887 &  x911 &  x914 &  x923 &  x926 &  x932 &  x944 &  x947 &  x953 &  x962 &  x971 &  x989 &  x1007 &  x1010 &  x1019 &  x1034 &  x1052 &  x1058 &  x1061 &  x1066 &  x1067 &  x1073 &  x1079 &  x1088 &  x1121 & ~x114 & ~x192 & ~x297;
assign c7182 =  x2 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x86 &  x89 &  x95 &  x98 &  x107 &  x110 &  x116 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x164 &  x167 &  x170 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x250 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x356 &  x359 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x391 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x443 &  x446 &  x449 &  x455 &  x458 &  x461 &  x464 &  x467 &  x469 &  x473 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x560 &  x563 &  x566 &  x569 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x671 &  x674 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x747 &  x748 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x773 &  x776 &  x779 &  x782 &  x785 &  x786 &  x787 &  x788 &  x791 &  x794 &  x797 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x826 &  x827 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x865 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x965 &  x971 &  x974 &  x977 &  x980 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x453 & ~x705 & ~x744 & ~x783 & ~x784 & ~x822 & ~x861;
assign c7184 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x148 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x170 &  x176 &  x179 &  x182 &  x185 &  x187 &  x188 &  x191 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x248 &  x251 &  x253 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x292 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x314 &  x317 &  x320 &  x323 &  x325 &  x326 &  x329 &  x332 &  x335 &  x338 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x403 &  x404 &  x407 &  x410 &  x413 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x442 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x509 &  x515 &  x518 &  x520 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x596 &  x599 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x653 &  x656 &  x659 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x695 &  x698 &  x704 &  x710 &  x713 &  x719 &  x722 &  x725 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x764 &  x767 &  x773 &  x775 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x806 &  x809 &  x812 &  x813 &  x814 &  x815 &  x818 &  x821 &  x824 &  x827 &  x833 &  x836 &  x845 &  x848 &  x851 &  x852 &  x853 &  x857 &  x860 &  x863 &  x869 &  x874 &  x875 &  x878 &  x884 &  x887 &  x890 &  x891 &  x892 &  x893 &  x899 &  x905 &  x908 &  x911 &  x913 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x931 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x952 &  x956 &  x962 &  x965 &  x968 &  x970 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1009 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1087 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130;
assign c7186 =  x8 &  x11 &  x26 &  x29 &  x35 &  x38 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x89 &  x92 &  x95 &  x98 &  x113 &  x116 &  x122 &  x125 &  x134 &  x146 &  x152 &  x158 &  x164 &  x173 &  x176 &  x179 &  x185 &  x188 &  x191 &  x194 &  x197 &  x215 &  x218 &  x221 &  x230 &  x236 &  x239 &  x242 &  x254 &  x257 &  x269 &  x281 &  x287 &  x299 &  x308 &  x311 &  x314 &  x317 &  x326 &  x329 &  x341 &  x344 &  x353 &  x356 &  x360 &  x362 &  x365 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x398 &  x400 &  x401 &  x404 &  x416 &  x422 &  x431 &  x437 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x464 &  x467 &  x473 &  x476 &  x479 &  x485 &  x488 &  x494 &  x503 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x548 &  x551 &  x554 &  x560 &  x563 &  x566 &  x569 &  x572 &  x581 &  x584 &  x587 &  x593 &  x596 &  x602 &  x608 &  x614 &  x617 &  x623 &  x626 &  x629 &  x635 &  x638 &  x641 &  x647 &  x650 &  x653 &  x659 &  x668 &  x677 &  x679 &  x680 &  x683 &  x686 &  x689 &  x695 &  x698 &  x701 &  x704 &  x707 &  x716 &  x718 &  x719 &  x722 &  x724 &  x731 &  x740 &  x743 &  x749 &  x752 &  x755 &  x758 &  x770 &  x773 &  x779 &  x785 &  x791 &  x809 &  x812 &  x815 &  x821 &  x824 &  x830 &  x845 &  x851 &  x854 &  x860 &  x866 &  x869 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x905 &  x917 &  x926 &  x932 &  x938 &  x941 &  x947 &  x950 &  x962 &  x971 &  x977 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1013 &  x1016 &  x1028 &  x1034 &  x1037 &  x1052 &  x1055 &  x1064 &  x1067 &  x1085 &  x1088 &  x1094 &  x1097 &  x1103 &  x1106 &  x1115 &  x1121 & ~x384 & ~x396 & ~x435 & ~x705 & ~x745 & ~x771 & ~x783;
assign c7188 =  x5 &  x8 &  x11 &  x14 &  x17 &  x26 &  x32 &  x35 &  x41 &  x44 &  x56 &  x59 &  x62 &  x65 &  x68 &  x77 &  x83 &  x86 &  x89 &  x95 &  x101 &  x104 &  x107 &  x110 &  x113 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x149 &  x155 &  x158 &  x164 &  x167 &  x176 &  x182 &  x185 &  x196 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x224 &  x227 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x275 &  x284 &  x287 &  x296 &  x302 &  x305 &  x311 &  x314 &  x317 &  x320 &  x323 &  x332 &  x335 &  x347 &  x356 &  x368 &  x371 &  x377 &  x380 &  x383 &  x392 &  x395 &  x401 &  x407 &  x410 &  x419 &  x425 &  x431 &  x434 &  x440 &  x443 &  x452 &  x467 &  x470 &  x476 &  x479 &  x488 &  x491 &  x494 &  x500 &  x512 &  x515 &  x530 &  x539 &  x545 &  x548 &  x551 &  x557 &  x563 &  x569 &  x575 &  x578 &  x584 &  x587 &  x590 &  x593 &  x596 &  x602 &  x605 &  x608 &  x614 &  x635 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x668 &  x674 &  x677 &  x683 &  x686 &  x689 &  x692 &  x698 &  x710 &  x713 &  x740 &  x743 &  x749 &  x752 &  x761 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x797 &  x806 &  x815 &  x821 &  x824 &  x827 &  x833 &  x836 &  x839 &  x851 &  x860 &  x866 &  x869 &  x884 &  x890 &  x893 &  x899 &  x902 &  x911 &  x917 &  x920 &  x926 &  x932 &  x935 &  x938 &  x947 &  x950 &  x956 &  x962 &  x971 &  x977 &  x980 &  x983 &  x986 &  x992 &  x1019 &  x1022 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1115 &  x1121 &  x1127 & ~x201 & ~x297 & ~x336 & ~x453 & ~x525 & ~x564 & ~x565 & ~x603 & ~x609 & ~x705 & ~x753;
assign c7190 =  x5 &  x11 &  x14 &  x20 &  x23 &  x26 &  x29 &  x38 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x71 &  x74 &  x77 &  x83 &  x86 &  x92 &  x98 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x131 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x266 &  x278 &  x281 &  x284 &  x293 &  x299 &  x302 &  x314 &  x317 &  x320 &  x323 &  x325 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x353 &  x359 &  x362 &  x364 &  x371 &  x374 &  x377 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x403 &  x404 &  x407 &  x413 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x446 &  x449 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x494 &  x497 &  x500 &  x503 &  x506 &  x508 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x542 &  x545 &  x547 &  x548 &  x551 &  x554 &  x557 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x586 &  x587 &  x590 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x757 &  x761 &  x767 &  x770 &  x773 &  x776 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x803 &  x806 &  x809 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x835 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x887 &  x890 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x929 &  x935 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x971 &  x974 &  x977 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1037 &  x1040 &  x1043 &  x1049 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x603 & ~x666 & ~x681 & ~x720 & ~x759 & ~x822 & ~x823 & ~x861 & ~x862 & ~x900 & ~x939;
assign c7192 =  x8 &  x14 &  x17 &  x29 &  x32 &  x38 &  x44 &  x65 &  x68 &  x74 &  x77 &  x86 &  x92 &  x101 &  x104 &  x107 &  x110 &  x119 &  x137 &  x146 &  x149 &  x155 &  x158 &  x161 &  x173 &  x191 &  x200 &  x209 &  x221 &  x230 &  x239 &  x242 &  x244 &  x266 &  x269 &  x281 &  x286 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x317 &  x320 &  x325 &  x326 &  x338 &  x341 &  x347 &  x350 &  x352 &  x356 &  x371 &  x380 &  x383 &  x386 &  x392 &  x394 &  x401 &  x404 &  x407 &  x416 &  x419 &  x428 &  x430 &  x431 &  x434 &  x440 &  x452 &  x455 &  x467 &  x479 &  x482 &  x485 &  x488 &  x491 &  x518 &  x521 &  x527 &  x530 &  x533 &  x536 &  x542 &  x545 &  x551 &  x557 &  x569 &  x572 &  x580 &  x581 &  x587 &  x593 &  x596 &  x602 &  x608 &  x614 &  x626 &  x632 &  x641 &  x656 &  x662 &  x665 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x704 &  x713 &  x719 &  x728 &  x731 &  x734 &  x737 &  x746 &  x752 &  x755 &  x764 &  x767 &  x770 &  x782 &  x800 &  x803 &  x806 &  x827 &  x830 &  x839 &  x848 &  x857 &  x866 &  x881 &  x896 &  x905 &  x920 &  x923 &  x938 &  x953 &  x956 &  x965 &  x971 &  x977 &  x983 &  x989 &  x995 &  x998 &  x1004 &  x1013 &  x1037 &  x1052 &  x1058 &  x1067 &  x1073 &  x1076 &  x1091 &  x1097 &  x1100 &  x1124 & ~x397 & ~x666 & ~x705 & ~x706 & ~x744 & ~x745 & ~x784 & ~x822;
assign c7194 =  x8 &  x11 &  x20 &  x32 &  x35 &  x41 &  x47 &  x53 &  x71 &  x77 &  x83 &  x89 &  x101 &  x104 &  x107 &  x125 &  x131 &  x137 &  x140 &  x146 &  x152 &  x176 &  x182 &  x185 &  x188 &  x200 &  x206 &  x212 &  x224 &  x227 &  x236 &  x245 &  x254 &  x257 &  x275 &  x284 &  x287 &  x290 &  x296 &  x299 &  x308 &  x311 &  x314 &  x317 &  x320 &  x329 &  x341 &  x344 &  x350 &  x356 &  x362 &  x365 &  x368 &  x371 &  x377 &  x383 &  x386 &  x389 &  x395 &  x410 &  x416 &  x419 &  x422 &  x428 &  x437 &  x440 &  x443 &  x455 &  x458 &  x470 &  x476 &  x479 &  x500 &  x503 &  x512 &  x527 &  x539 &  x542 &  x551 &  x554 &  x556 &  x563 &  x569 &  x578 &  x584 &  x587 &  x596 &  x599 &  x614 &  x623 &  x635 &  x641 &  x647 &  x656 &  x662 &  x665 &  x674 &  x677 &  x692 &  x704 &  x716 &  x731 &  x737 &  x740 &  x742 &  x752 &  x755 &  x758 &  x764 &  x767 &  x773 &  x776 &  x779 &  x782 &  x794 &  x800 &  x812 &  x818 &  x824 &  x833 &  x842 &  x848 &  x851 &  x857 &  x863 &  x875 &  x878 &  x884 &  x887 &  x890 &  x893 &  x899 &  x908 &  x914 &  x917 &  x920 &  x923 &  x935 &  x941 &  x953 &  x959 &  x965 &  x995 &  x1010 &  x1013 &  x1016 &  x1025 &  x1031 &  x1037 &  x1040 &  x1046 &  x1076 &  x1082 &  x1085 &  x1091 &  x1097 &  x1103 &  x1109 &  x1114 &  x1124 &  x1130 & ~x234 & ~x390 & ~x921 & ~x1017 & ~x1018 & ~x1057 & ~x1095 & ~x1096;
assign c7196 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x23 &  x26 &  x32 &  x35 &  x38 &  x41 &  x43 &  x44 &  x47 &  x50 &  x53 &  x59 &  x62 &  x65 &  x71 &  x74 &  x77 &  x80 &  x82 &  x83 &  x89 &  x95 &  x98 &  x101 &  x107 &  x113 &  x119 &  x121 &  x122 &  x125 &  x127 &  x128 &  x131 &  x143 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x179 &  x182 &  x185 &  x188 &  x191 &  x203 &  x206 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x274 &  x275 &  x278 &  x281 &  x284 &  x287 &  x289 &  x290 &  x293 &  x299 &  x302 &  x305 &  x311 &  x314 &  x317 &  x323 &  x326 &  x328 &  x332 &  x338 &  x341 &  x350 &  x356 &  x359 &  x362 &  x365 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x401 &  x404 &  x406 &  x410 &  x412 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x437 &  x444 &  x445 &  x446 &  x452 &  x458 &  x461 &  x467 &  x473 &  x476 &  x479 &  x484 &  x488 &  x491 &  x497 &  x500 &  x503 &  x506 &  x512 &  x515 &  x518 &  x521 &  x523 &  x524 &  x527 &  x530 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x584 &  x587 &  x590 &  x596 &  x599 &  x601 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x623 &  x629 &  x632 &  x638 &  x640 &  x641 &  x644 &  x647 &  x656 &  x662 &  x665 &  x668 &  x670 &  x671 &  x674 &  x679 &  x680 &  x685 &  x686 &  x689 &  x695 &  x698 &  x701 &  x704 &  x707 &  x709 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x740 &  x746 &  x749 &  x755 &  x758 &  x761 &  x779 &  x782 &  x785 &  x791 &  x794 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x824 &  x833 &  x836 &  x842 &  x845 &  x848 &  x854 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x962 &  x968 &  x974 &  x977 &  x980 &  x983 &  x989 &  x992 &  x995 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1058 &  x1073 &  x1076 &  x1079 &  x1082 &  x1088 &  x1097 &  x1100 &  x1103 &  x1109 &  x1115 &  x1121 &  x1127 &  x1130 & ~x219 & ~x258 & ~x666 & ~x705 & ~x744;
assign c7198 =  x2 &  x5 &  x8 &  x11 &  x14 &  x20 &  x26 &  x32 &  x35 &  x38 &  x44 &  x47 &  x50 &  x53 &  x56 &  x62 &  x65 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x131 &  x134 &  x140 &  x143 &  x146 &  x149 &  x155 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x244 &  x245 &  x248 &  x254 &  x260 &  x263 &  x272 &  x275 &  x278 &  x281 &  x283 &  x284 &  x286 &  x287 &  x290 &  x293 &  x296 &  x299 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x322 &  x323 &  x324 &  x326 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x352 &  x353 &  x356 &  x359 &  x361 &  x362 &  x364 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x389 &  x391 &  x395 &  x398 &  x400 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x422 &  x428 &  x430 &  x431 &  x437 &  x440 &  x446 &  x449 &  x455 &  x458 &  x461 &  x464 &  x467 &  x469 &  x470 &  x473 &  x476 &  x479 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x508 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x545 &  x547 &  x548 &  x551 &  x554 &  x557 &  x560 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x674 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x704 &  x707 &  x713 &  x716 &  x719 &  x722 &  x725 &  x734 &  x737 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x770 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x815 &  x818 &  x821 &  x824 &  x827 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x453 & ~x492 & ~x531 & ~x666 & ~x705 & ~x706 & ~x744 & ~x745 & ~x783 & ~x784 & ~x822;
assign c7200 =  x8 &  x17 &  x23 &  x38 &  x44 &  x53 &  x56 &  x62 &  x65 &  x70 &  x71 &  x80 &  x86 &  x89 &  x92 &  x95 &  x97 &  x98 &  x101 &  x110 &  x119 &  x122 &  x128 &  x130 &  x131 &  x143 &  x149 &  x152 &  x167 &  x173 &  x179 &  x185 &  x191 &  x197 &  x200 &  x208 &  x212 &  x215 &  x221 &  x224 &  x233 &  x239 &  x248 &  x254 &  x257 &  x269 &  x272 &  x281 &  x290 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x329 &  x338 &  x341 &  x350 &  x353 &  x356 &  x359 &  x365 &  x377 &  x398 &  x401 &  x407 &  x422 &  x425 &  x431 &  x434 &  x437 &  x446 &  x449 &  x461 &  x473 &  x479 &  x482 &  x503 &  x506 &  x509 &  x512 &  x554 &  x557 &  x560 &  x563 &  x572 &  x587 &  x593 &  x596 &  x599 &  x602 &  x611 &  x614 &  x617 &  x626 &  x635 &  x638 &  x644 &  x650 &  x656 &  x659 &  x662 &  x665 &  x668 &  x674 &  x677 &  x686 &  x692 &  x695 &  x707 &  x728 &  x737 &  x743 &  x755 &  x764 &  x773 &  x779 &  x791 &  x794 &  x797 &  x806 &  x809 &  x812 &  x821 &  x824 &  x827 &  x839 &  x842 &  x845 &  x860 &  x863 &  x869 &  x890 &  x896 &  x899 &  x902 &  x908 &  x917 &  x923 &  x929 &  x935 &  x938 &  x950 &  x953 &  x956 &  x962 &  x971 &  x980 &  x983 &  x986 &  x989 &  x998 &  x1004 &  x1013 &  x1019 &  x1022 &  x1046 &  x1058 &  x1061 &  x1067 &  x1070 &  x1076 &  x1085 &  x1088 &  x1091 &  x1097 &  x1103 &  x1106 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 & ~x306 & ~x319 & ~x372 & ~x417 & ~x456;
assign c7202 =  x2 &  x5 &  x14 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x44 &  x47 &  x56 &  x59 &  x62 &  x65 &  x68 &  x77 &  x86 &  x89 &  x92 &  x95 &  x98 &  x104 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x131 &  x134 &  x140 &  x149 &  x152 &  x155 &  x161 &  x167 &  x170 &  x176 &  x179 &  x182 &  x188 &  x194 &  x197 &  x200 &  x203 &  x205 &  x206 &  x208 &  x209 &  x212 &  x215 &  x218 &  x221 &  x227 &  x230 &  x233 &  x235 &  x236 &  x239 &  x245 &  x248 &  x254 &  x257 &  x263 &  x266 &  x278 &  x281 &  x284 &  x299 &  x305 &  x308 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x338 &  x344 &  x350 &  x352 &  x353 &  x356 &  x359 &  x368 &  x371 &  x374 &  x380 &  x386 &  x389 &  x392 &  x398 &  x401 &  x404 &  x407 &  x413 &  x416 &  x419 &  x425 &  x431 &  x434 &  x440 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x476 &  x479 &  x482 &  x485 &  x488 &  x494 &  x497 &  x506 &  x512 &  x518 &  x521 &  x524 &  x527 &  x530 &  x539 &  x541 &  x542 &  x545 &  x548 &  x551 &  x557 &  x560 &  x563 &  x566 &  x572 &  x578 &  x580 &  x581 &  x584 &  x590 &  x593 &  x596 &  x599 &  x602 &  x608 &  x614 &  x620 &  x623 &  x626 &  x629 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x656 &  x659 &  x662 &  x670 &  x671 &  x677 &  x680 &  x683 &  x689 &  x695 &  x704 &  x707 &  x710 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x743 &  x746 &  x752 &  x755 &  x758 &  x764 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x800 &  x806 &  x809 &  x812 &  x815 &  x821 &  x824 &  x827 &  x833 &  x836 &  x839 &  x845 &  x848 &  x851 &  x854 &  x866 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x896 &  x899 &  x902 &  x905 &  x911 &  x914 &  x917 &  x920 &  x926 &  x929 &  x935 &  x938 &  x944 &  x947 &  x953 &  x956 &  x959 &  x968 &  x974 &  x986 &  x992 &  x998 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1031 &  x1043 &  x1049 &  x1055 &  x1058 &  x1064 &  x1070 &  x1079 &  x1082 &  x1088 &  x1094 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1121 &  x1127 &  x1130 & ~x666 & ~x705 & ~x741 & ~x1101;
assign c7204 =  x29 &  x32 &  x83 &  x89 &  x92 &  x107 &  x110 &  x134 &  x143 &  x185 &  x188 &  x197 &  x212 &  x215 &  x221 &  x224 &  x233 &  x239 &  x248 &  x254 &  x257 &  x275 &  x278 &  x308 &  x317 &  x347 &  x350 &  x371 &  x383 &  x398 &  x404 &  x437 &  x442 &  x455 &  x473 &  x479 &  x481 &  x482 &  x494 &  x509 &  x515 &  x524 &  x545 &  x563 &  x569 &  x601 &  x659 &  x680 &  x701 &  x704 &  x713 &  x758 &  x782 &  x785 &  x797 &  x806 &  x818 &  x827 &  x830 &  x833 &  x836 &  x842 &  x851 &  x863 &  x932 &  x937 &  x941 &  x962 &  x965 &  x992 &  x1021 &  x1025 &  x1029 &  x1037 &  x1052 &  x1064 &  x1067 &  x1085 &  x1088 &  x1091 &  x1106 &  x1108 &  x1109 & ~x765;
assign c7206 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x41 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x80 &  x83 &  x86 &  x89 &  x95 &  x98 &  x101 &  x110 &  x113 &  x116 &  x122 &  x125 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x158 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x227 &  x230 &  x233 &  x236 &  x245 &  x248 &  x251 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x296 &  x302 &  x305 &  x311 &  x317 &  x320 &  x323 &  x332 &  x335 &  x338 &  x344 &  x350 &  x353 &  x359 &  x361 &  x362 &  x365 &  x368 &  x371 &  x377 &  x383 &  x386 &  x392 &  x398 &  x400 &  x401 &  x404 &  x407 &  x413 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x439 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x470 &  x476 &  x478 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x530 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x575 &  x590 &  x593 &  x596 &  x599 &  x605 &  x608 &  x614 &  x617 &  x620 &  x625 &  x626 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x701 &  x703 &  x704 &  x707 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x737 &  x740 &  x742 &  x743 &  x746 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x776 &  x779 &  x781 &  x788 &  x794 &  x800 &  x803 &  x812 &  x815 &  x820 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x851 &  x854 &  x860 &  x863 &  x869 &  x872 &  x875 &  x881 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x914 &  x917 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x950 &  x953 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1016 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x396 & ~x435 & ~x648 & ~x831 & ~x861 & ~x870 & ~x909 & ~x948 & ~x987 & ~x988 & ~x1026;
assign c7208 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x88 &  x89 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x127 &  x128 &  x131 &  x134 &  x140 &  x143 &  x146 &  x149 &  x152 &  x157 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x196 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x234 &  x235 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x269 &  x272 &  x274 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x302 &  x305 &  x308 &  x311 &  x313 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x617 &  x620 &  x623 &  x626 &  x629 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x758 &  x761 &  x767 &  x770 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x968 &  x971 &  x974 &  x977 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x114 & ~x153 & ~x180 & ~x219 & ~x297 & ~x432 & ~x471 & ~x472 & ~x510 & ~x511 & ~x549 & ~x588 & ~x624 & ~x663 & ~x702 & ~x741 & ~x780 & ~x819;
assign c7210 =  x1 &  x5 &  x8 &  x20 &  x23 &  x26 &  x32 &  x35 &  x38 &  x40 &  x44 &  x49 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x79 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x110 &  x113 &  x116 &  x118 &  x119 &  x122 &  x125 &  x128 &  x131 &  x137 &  x140 &  x143 &  x149 &  x155 &  x157 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x185 &  x188 &  x191 &  x196 &  x197 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x266 &  x272 &  x275 &  x278 &  x284 &  x290 &  x293 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x368 &  x371 &  x380 &  x389 &  x392 &  x395 &  x398 &  x401 &  x407 &  x410 &  x413 &  x416 &  x428 &  x431 &  x434 &  x437 &  x440 &  x446 &  x449 &  x452 &  x455 &  x458 &  x467 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x497 &  x503 &  x506 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x545 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x587 &  x590 &  x593 &  x596 &  x599 &  x601 &  x602 &  x605 &  x611 &  x620 &  x623 &  x629 &  x632 &  x635 &  x638 &  x640 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x680 &  x683 &  x689 &  x692 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x770 &  x776 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x809 &  x812 &  x815 &  x821 &  x824 &  x830 &  x833 &  x839 &  x842 &  x845 &  x851 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x926 &  x938 &  x944 &  x947 &  x950 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x977 &  x980 &  x983 &  x989 &  x992 &  x995 &  x1007 &  x1010 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1037 &  x1043 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1076 &  x1079 &  x1082 &  x1091 &  x1100 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 & ~x7 & ~x24 & ~x84 & ~x85 & ~x102 & ~x123 & ~x135 & ~x162 & ~x174 & ~x180 & ~x258 & ~x297 & ~x336 & ~x354 & ~x375 & ~x393 & ~x414 & ~x783 & ~x822 & ~x861;
assign c7212 =  x2 &  x5 &  x11 &  x17 &  x20 &  x26 &  x32 &  x35 &  x38 &  x41 &  x44 &  x50 &  x53 &  x56 &  x59 &  x65 &  x68 &  x74 &  x80 &  x86 &  x89 &  x95 &  x101 &  x104 &  x107 &  x113 &  x116 &  x122 &  x125 &  x128 &  x134 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x230 &  x233 &  x236 &  x242 &  x245 &  x248 &  x251 &  x257 &  x266 &  x272 &  x290 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x332 &  x341 &  x347 &  x353 &  x359 &  x362 &  x365 &  x368 &  x377 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x404 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x467 &  x470 &  x473 &  x476 &  x488 &  x491 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x593 &  x596 &  x599 &  x605 &  x608 &  x611 &  x614 &  x617 &  x623 &  x626 &  x629 &  x632 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x674 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x710 &  x713 &  x716 &  x719 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x758 &  x761 &  x767 &  x779 &  x782 &  x791 &  x794 &  x797 &  x800 &  x806 &  x809 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x839 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x869 &  x872 &  x878 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x905 &  x911 &  x914 &  x920 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x962 &  x965 &  x968 &  x974 &  x977 &  x980 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1019 &  x1022 &  x1025 &  x1028 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1127 & ~x504 & ~x594 & ~x633 & ~x634 & ~x666 & ~x672 & ~x673 & ~x705 & ~x706 & ~x711 & ~x712 & ~x744 & ~x745 & ~x750 & ~x780 & ~x783 & ~x789 & ~x819 & ~x822 & ~x858 & ~x861 & ~x897 & ~x936 & ~x975;
assign c7214 =  x2 &  x5 &  x35 &  x44 &  x53 &  x62 &  x65 &  x71 &  x77 &  x83 &  x119 &  x140 &  x152 &  x170 &  x182 &  x188 &  x200 &  x209 &  x227 &  x239 &  x269 &  x272 &  x275 &  x287 &  x302 &  x311 &  x323 &  x324 &  x329 &  x332 &  x335 &  x338 &  x341 &  x356 &  x359 &  x365 &  x371 &  x377 &  x380 &  x386 &  x389 &  x392 &  x398 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x429 &  x452 &  x458 &  x479 &  x485 &  x488 &  x491 &  x497 &  x500 &  x503 &  x506 &  x524 &  x557 &  x566 &  x569 &  x586 &  x587 &  x590 &  x599 &  x602 &  x611 &  x617 &  x623 &  x629 &  x659 &  x665 &  x671 &  x683 &  x689 &  x692 &  x695 &  x698 &  x710 &  x713 &  x719 &  x728 &  x734 &  x740 &  x752 &  x776 &  x788 &  x800 &  x830 &  x836 &  x839 &  x845 &  x860 &  x890 &  x893 &  x899 &  x911 &  x914 &  x917 &  x923 &  x938 &  x944 &  x956 &  x959 &  x962 &  x965 &  x977 &  x989 &  x1010 &  x1019 &  x1025 &  x1028 &  x1031 &  x1037 &  x1052 &  x1058 &  x1067 &  x1073 &  x1088 &  x1091 &  x1094 &  x1097 &  x1109 &  x1115 &  x1118 &  x1130 & ~x318 & ~x666 & ~x667 & ~x706 & ~x744 & ~x745 & ~x783 & ~x822 & ~x861;
assign c7216 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x64 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x103 &  x104 &  x107 &  x110 &  x116 &  x119 &  x122 &  x128 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x175 &  x176 &  x179 &  x182 &  x185 &  x187 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x305 &  x308 &  x311 &  x314 &  x317 &  x323 &  x325 &  x326 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x364 &  x365 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x392 &  x395 &  x398 &  x403 &  x404 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x434 &  x437 &  x443 &  x446 &  x449 &  x455 &  x458 &  x461 &  x464 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x640 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x704 &  x707 &  x709 &  x713 &  x716 &  x719 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x785 &  x788 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x827 &  x833 &  x836 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x959 &  x965 &  x968 &  x971 &  x974 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x396 & ~x435 & ~x666 & ~x705 & ~x706 & ~x783 & ~x822;
assign c7218 =  x2 &  x8 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x35 &  x44 &  x47 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x104 &  x107 &  x113 &  x122 &  x131 &  x143 &  x146 &  x149 &  x155 &  x158 &  x161 &  x170 &  x182 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x227 &  x230 &  x233 &  x236 &  x248 &  x254 &  x260 &  x266 &  x272 &  x275 &  x281 &  x287 &  x293 &  x299 &  x308 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x335 &  x338 &  x347 &  x353 &  x365 &  x377 &  x380 &  x386 &  x392 &  x398 &  x413 &  x419 &  x422 &  x437 &  x439 &  x440 &  x442 &  x443 &  x452 &  x467 &  x473 &  x476 &  x477 &  x478 &  x479 &  x481 &  x482 &  x488 &  x491 &  x500 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x545 &  x547 &  x551 &  x554 &  x557 &  x560 &  x569 &  x584 &  x586 &  x587 &  x589 &  x590 &  x596 &  x599 &  x602 &  x605 &  x608 &  x625 &  x626 &  x632 &  x638 &  x644 &  x647 &  x650 &  x653 &  x659 &  x662 &  x664 &  x665 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x725 &  x731 &  x737 &  x740 &  x749 &  x752 &  x755 &  x761 &  x764 &  x770 &  x773 &  x776 &  x779 &  x782 &  x788 &  x797 &  x803 &  x806 &  x809 &  x812 &  x815 &  x824 &  x830 &  x836 &  x842 &  x845 &  x848 &  x854 &  x857 &  x866 &  x869 &  x872 &  x875 &  x878 &  x890 &  x896 &  x899 &  x902 &  x905 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x935 &  x941 &  x947 &  x953 &  x956 &  x959 &  x965 &  x971 &  x974 &  x980 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1076 &  x1082 &  x1091 &  x1103 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x552 & ~x591 & ~x592 & ~x900 & ~x939;
assign c7220 =  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x116 &  x119 &  x122 &  x125 &  x131 &  x140 &  x143 &  x146 &  x152 &  x158 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x257 &  x260 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x296 &  x299 &  x302 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x335 &  x338 &  x341 &  x344 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x380 &  x389 &  x392 &  x395 &  x404 &  x413 &  x419 &  x422 &  x425 &  x431 &  x434 &  x437 &  x442 &  x443 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x479 &  x481 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x506 &  x509 &  x512 &  x515 &  x518 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x581 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x611 &  x614 &  x617 &  x623 &  x626 &  x632 &  x638 &  x641 &  x644 &  x647 &  x650 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x683 &  x689 &  x698 &  x701 &  x710 &  x713 &  x716 &  x722 &  x728 &  x731 &  x734 &  x737 &  x743 &  x746 &  x752 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x800 &  x806 &  x809 &  x812 &  x815 &  x821 &  x827 &  x839 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x878 &  x881 &  x884 &  x887 &  x893 &  x899 &  x905 &  x908 &  x914 &  x917 &  x920 &  x926 &  x938 &  x947 &  x956 &  x959 &  x962 &  x970 &  x971 &  x974 &  x986 &  x989 &  x992 &  x998 &  x1004 &  x1007 &  x1013 &  x1016 &  x1022 &  x1025 &  x1031 &  x1036 &  x1037 &  x1040 &  x1043 &  x1046 &  x1048 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1087 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 & ~x15 & ~x54 & ~x93 & ~x132 & ~x171 & ~x234 & ~x273 & ~x312 & ~x978;
assign c7222 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x308 &  x311 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x452 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x796 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x874 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1069 &  x1070 &  x1073 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 & ~x21 & ~x60 & ~x99 & ~x138 & ~x189 & ~x276 & ~x315 & ~x354 & ~x432 & ~x471 & ~x510 & ~x588 & ~x627 & ~x846;
assign c7224 =  x38 &  x41 &  x74 &  x77 &  x80 &  x83 &  x86 &  x95 &  x98 &  x116 &  x122 &  x140 &  x143 &  x158 &  x161 &  x164 &  x182 &  x188 &  x206 &  x221 &  x227 &  x239 &  x257 &  x260 &  x272 &  x281 &  x290 &  x317 &  x344 &  x359 &  x368 &  x389 &  x392 &  x416 &  x419 &  x422 &  x446 &  x482 &  x491 &  x503 &  x509 &  x520 &  x521 &  x527 &  x530 &  x542 &  x548 &  x551 &  x554 &  x563 &  x578 &  x593 &  x608 &  x634 &  x647 &  x659 &  x662 &  x665 &  x673 &  x695 &  x701 &  x710 &  x716 &  x734 &  x740 &  x751 &  x752 &  x761 &  x767 &  x780 &  x782 &  x785 &  x800 &  x803 &  x815 &  x819 &  x820 &  x827 &  x833 &  x839 &  x845 &  x858 &  x859 &  x875 &  x878 &  x899 &  x911 &  x926 &  x944 &  x956 &  x965 &  x974 &  x980 &  x986 &  x992 &  x1028 &  x1037 &  x1058 &  x1064 &  x1069 &  x1073 &  x1085 &  x1121 & ~x237 & ~x276 & ~x471 & ~x978;
assign c7226 =  x2 &  x5 &  x11 &  x13 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x52 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x80 &  x86 &  x89 &  x91 &  x95 &  x98 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x128 &  x130 &  x131 &  x134 &  x137 &  x140 &  x146 &  x149 &  x152 &  x158 &  x161 &  x164 &  x167 &  x168 &  x169 &  x170 &  x173 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x205 &  x206 &  x207 &  x208 &  x212 &  x218 &  x221 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x247 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x274 &  x275 &  x284 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x350 &  x352 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x374 &  x380 &  x386 &  x389 &  x392 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x428 &  x431 &  x434 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x482 &  x485 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x521 &  x524 &  x530 &  x533 &  x536 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x580 &  x581 &  x587 &  x590 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x659 &  x662 &  x665 &  x668 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x698 &  x704 &  x707 &  x710 &  x713 &  x716 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x749 &  x752 &  x755 &  x758 &  x761 &  x770 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x824 &  x827 &  x833 &  x836 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x866 &  x869 &  x878 &  x881 &  x884 &  x887 &  x893 &  x896 &  x902 &  x905 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x959 &  x962 &  x965 &  x971 &  x974 &  x980 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1007 &  x1013 &  x1016 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 &  x1130 & ~x549 & ~x588 & ~x589 & ~x627 & ~x666;
assign c7228 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x38 &  x53 &  x56 &  x62 &  x65 &  x68 &  x74 &  x80 &  x86 &  x92 &  x98 &  x101 &  x104 &  x128 &  x133 &  x137 &  x140 &  x143 &  x152 &  x164 &  x170 &  x176 &  x179 &  x188 &  x194 &  x197 &  x200 &  x203 &  x209 &  x211 &  x227 &  x236 &  x251 &  x263 &  x269 &  x278 &  x284 &  x287 &  x293 &  x299 &  x305 &  x308 &  x314 &  x320 &  x323 &  x326 &  x338 &  x341 &  x347 &  x353 &  x359 &  x362 &  x365 &  x368 &  x377 &  x389 &  x392 &  x395 &  x404 &  x406 &  x416 &  x419 &  x425 &  x430 &  x443 &  x446 &  x449 &  x455 &  x458 &  x461 &  x469 &  x470 &  x479 &  x485 &  x491 &  x494 &  x497 &  x503 &  x515 &  x518 &  x527 &  x530 &  x533 &  x539 &  x542 &  x545 &  x548 &  x557 &  x560 &  x562 &  x563 &  x572 &  x578 &  x584 &  x587 &  x590 &  x596 &  x599 &  x601 &  x605 &  x608 &  x620 &  x638 &  x640 &  x644 &  x647 &  x662 &  x665 &  x677 &  x679 &  x680 &  x685 &  x686 &  x692 &  x710 &  x713 &  x716 &  x724 &  x725 &  x728 &  x740 &  x746 &  x749 &  x755 &  x756 &  x757 &  x761 &  x763 &  x764 &  x770 &  x773 &  x779 &  x785 &  x788 &  x791 &  x795 &  x797 &  x800 &  x809 &  x812 &  x814 &  x815 &  x821 &  x824 &  x827 &  x830 &  x834 &  x842 &  x851 &  x854 &  x860 &  x866 &  x869 &  x872 &  x873 &  x874 &  x887 &  x890 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x935 &  x950 &  x952 &  x956 &  x959 &  x971 &  x977 &  x986 &  x991 &  x998 &  x1016 &  x1025 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1064 &  x1070 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1106 &  x1112 &  x1115 &  x1127 &  x1130 & ~x396 & ~x783 & ~x822 & ~x861;
assign c7230 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x110 &  x113 &  x116 &  x119 &  x125 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x209 &  x212 &  x215 &  x221 &  x224 &  x227 &  x230 &  x233 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x317 &  x320 &  x323 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x452 &  x455 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x481 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x520 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x710 &  x716 &  x719 &  x722 &  x725 &  x734 &  x737 &  x740 &  x742 &  x743 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x773 &  x781 &  x782 &  x785 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x820 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x859 &  x863 &  x866 &  x869 &  x872 &  x875 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x898 &  x899 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x926 &  x929 &  x932 &  x935 &  x937 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x976 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x998 &  x1001 &  x1004 &  x1010 &  x1015 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1054 &  x1055 &  x1058 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1091 &  x1093 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x606 & ~x645 & ~x765 & ~x804 & ~x849 & ~x888 & ~x900 & ~x939 & ~x966 & ~x978 & ~x1017 & ~x1044 & ~x1056 & ~x1083 & ~x1095 & ~x1122;
assign c7232 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x95 &  x98 &  x101 &  x110 &  x113 &  x116 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x164 &  x167 &  x170 &  x173 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x266 &  x269 &  x272 &  x274 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x314 &  x317 &  x320 &  x329 &  x332 &  x335 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x443 &  x449 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x542 &  x551 &  x554 &  x557 &  x560 &  x563 &  x572 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x602 &  x611 &  x614 &  x617 &  x619 &  x620 &  x623 &  x626 &  x632 &  x635 &  x641 &  x644 &  x647 &  x653 &  x657 &  x658 &  x659 &  x662 &  x665 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x696 &  x697 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x728 &  x736 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x761 &  x764 &  x767 &  x770 &  x773 &  x775 &  x776 &  x779 &  x782 &  x785 &  x791 &  x794 &  x797 &  x800 &  x803 &  x809 &  x812 &  x814 &  x815 &  x818 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x845 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x872 &  x878 &  x881 &  x884 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x920 &  x923 &  x929 &  x932 &  x935 &  x941 &  x947 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x980 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1043 &  x1046 &  x1049 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1088 &  x1094 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x231 & ~x333 & ~x447 & ~x525 & ~x588 & ~x627 & ~x666 & ~x705 & ~x744 & ~x783;
assign c7234 =  x2 &  x5 &  x8 &  x11 &  x17 &  x29 &  x32 &  x35 &  x43 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x74 &  x77 &  x83 &  x86 &  x89 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x121 &  x122 &  x125 &  x131 &  x137 &  x143 &  x152 &  x155 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x188 &  x191 &  x194 &  x200 &  x203 &  x209 &  x212 &  x215 &  x221 &  x227 &  x233 &  x239 &  x251 &  x254 &  x257 &  x269 &  x272 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x302 &  x305 &  x311 &  x314 &  x317 &  x320 &  x329 &  x335 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x359 &  x365 &  x368 &  x371 &  x374 &  x377 &  x383 &  x386 &  x389 &  x392 &  x401 &  x404 &  x407 &  x416 &  x422 &  x428 &  x431 &  x434 &  x437 &  x449 &  x455 &  x458 &  x461 &  x470 &  x473 &  x476 &  x491 &  x497 &  x500 &  x503 &  x509 &  x512 &  x518 &  x530 &  x533 &  x536 &  x539 &  x548 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x590 &  x593 &  x596 &  x599 &  x605 &  x614 &  x617 &  x620 &  x623 &  x626 &  x638 &  x641 &  x647 &  x650 &  x653 &  x656 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x691 &  x698 &  x701 &  x707 &  x713 &  x716 &  x719 &  x725 &  x728 &  x734 &  x737 &  x743 &  x746 &  x749 &  x758 &  x760 &  x761 &  x767 &  x768 &  x770 &  x773 &  x779 &  x782 &  x788 &  x791 &  x797 &  x800 &  x806 &  x815 &  x818 &  x821 &  x827 &  x833 &  x836 &  x839 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x869 &  x878 &  x881 &  x884 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x917 &  x920 &  x923 &  x929 &  x938 &  x947 &  x953 &  x956 &  x959 &  x965 &  x968 &  x974 &  x980 &  x983 &  x986 &  x989 &  x1010 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1034 &  x1037 &  x1049 &  x1055 &  x1058 &  x1064 &  x1070 &  x1076 &  x1082 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1127 &  x1130 & ~x633 & ~x744 & ~x783 & ~x816 & ~x855 & ~x894;
assign c7236 =  x14 &  x20 &  x23 &  x26 &  x29 &  x41 &  x43 &  x44 &  x50 &  x53 &  x56 &  x82 &  x89 &  x107 &  x116 &  x131 &  x137 &  x158 &  x173 &  x197 &  x200 &  x218 &  x224 &  x230 &  x254 &  x265 &  x266 &  x287 &  x308 &  x311 &  x317 &  x335 &  x340 &  x341 &  x344 &  x347 &  x350 &  x362 &  x373 &  x379 &  x380 &  x397 &  x404 &  x416 &  x425 &  x461 &  x488 &  x491 &  x497 &  x519 &  x542 &  x566 &  x572 &  x587 &  x599 &  x602 &  x620 &  x641 &  x644 &  x656 &  x662 &  x677 &  x698 &  x701 &  x704 &  x707 &  x713 &  x722 &  x743 &  x746 &  x758 &  x770 &  x773 &  x776 &  x785 &  x797 &  x800 &  x836 &  x842 &  x848 &  x859 &  x872 &  x878 &  x896 &  x913 &  x914 &  x956 &  x959 &  x974 &  x983 &  x989 &  x998 &  x1004 &  x1007 &  x1022 &  x1040 &  x1046 &  x1052 &  x1085 &  x1088 &  x1094 &  x1100 &  x1130;
assign c7238 =  x5 &  x14 &  x20 &  x23 &  x26 &  x29 &  x35 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x74 &  x77 &  x86 &  x92 &  x104 &  x113 &  x128 &  x134 &  x146 &  x149 &  x152 &  x155 &  x161 &  x164 &  x170 &  x179 &  x182 &  x185 &  x191 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x224 &  x227 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x266 &  x272 &  x275 &  x278 &  x281 &  x284 &  x290 &  x296 &  x308 &  x311 &  x314 &  x323 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x362 &  x365 &  x368 &  x389 &  x392 &  x404 &  x413 &  x416 &  x422 &  x425 &  x428 &  x431 &  x434 &  x443 &  x446 &  x452 &  x461 &  x464 &  x470 &  x482 &  x488 &  x494 &  x497 &  x506 &  x512 &  x515 &  x524 &  x527 &  x536 &  x539 &  x542 &  x545 &  x554 &  x556 &  x557 &  x560 &  x569 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x595 &  x596 &  x602 &  x605 &  x608 &  x614 &  x617 &  x623 &  x632 &  x638 &  x641 &  x644 &  x650 &  x653 &  x656 &  x664 &  x665 &  x668 &  x674 &  x677 &  x683 &  x686 &  x695 &  x698 &  x701 &  x703 &  x710 &  x713 &  x716 &  x719 &  x722 &  x728 &  x731 &  x734 &  x742 &  x752 &  x755 &  x758 &  x761 &  x767 &  x770 &  x773 &  x779 &  x781 &  x782 &  x788 &  x791 &  x794 &  x797 &  x800 &  x812 &  x815 &  x821 &  x824 &  x839 &  x842 &  x845 &  x848 &  x854 &  x859 &  x863 &  x866 &  x869 &  x875 &  x884 &  x887 &  x890 &  x896 &  x898 &  x899 &  x905 &  x908 &  x917 &  x920 &  x926 &  x932 &  x937 &  x938 &  x941 &  x947 &  x950 &  x953 &  x962 &  x965 &  x974 &  x976 &  x986 &  x989 &  x992 &  x998 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1055 &  x1061 &  x1064 &  x1070 &  x1076 &  x1079 &  x1088 &  x1091 &  x1100 &  x1103 &  x1115 &  x1118 &  x1127 & ~x312 & ~x354 & ~x390 & ~x393 & ~x471 & ~x630 & ~x669 & ~x765 & ~x804 & ~x921 & ~x960 & ~x1056;
assign c7240 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x41 &  x47 &  x56 &  x59 &  x62 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x98 &  x101 &  x104 &  x107 &  x110 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x143 &  x146 &  x149 &  x155 &  x164 &  x167 &  x170 &  x173 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x209 &  x212 &  x215 &  x218 &  x230 &  x233 &  x236 &  x239 &  x242 &  x248 &  x251 &  x254 &  x257 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x359 &  x365 &  x371 &  x374 &  x377 &  x383 &  x386 &  x389 &  x392 &  x395 &  x401 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x440 &  x443 &  x446 &  x449 &  x455 &  x458 &  x461 &  x464 &  x467 &  x473 &  x476 &  x478 &  x479 &  x482 &  x491 &  x494 &  x497 &  x500 &  x503 &  x512 &  x515 &  x518 &  x521 &  x524 &  x530 &  x533 &  x536 &  x542 &  x545 &  x551 &  x554 &  x556 &  x557 &  x559 &  x563 &  x569 &  x572 &  x575 &  x587 &  x590 &  x595 &  x598 &  x599 &  x602 &  x605 &  x608 &  x614 &  x617 &  x620 &  x626 &  x629 &  x635 &  x638 &  x641 &  x647 &  x650 &  x653 &  x656 &  x662 &  x665 &  x668 &  x677 &  x680 &  x683 &  x686 &  x689 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x719 &  x725 &  x728 &  x734 &  x737 &  x742 &  x743 &  x752 &  x755 &  x761 &  x764 &  x767 &  x770 &  x776 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x806 &  x812 &  x818 &  x820 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x848 &  x851 &  x859 &  x863 &  x869 &  x872 &  x875 &  x881 &  x884 &  x890 &  x893 &  x896 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x926 &  x929 &  x932 &  x935 &  x937 &  x941 &  x944 &  x947 &  x953 &  x956 &  x959 &  x962 &  x968 &  x974 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1064 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1127 &  x1130 & ~x273 & ~x312 & ~x351 & ~x354 & ~x390 & ~x432 & ~x1017 & ~x1018 & ~x1057;
assign c7242 =  x2 &  x11 &  x17 &  x26 &  x32 &  x35 &  x38 &  x44 &  x50 &  x65 &  x68 &  x71 &  x77 &  x86 &  x95 &  x98 &  x107 &  x110 &  x113 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x173 &  x176 &  x179 &  x182 &  x191 &  x194 &  x197 &  x206 &  x212 &  x215 &  x218 &  x221 &  x224 &  x230 &  x233 &  x236 &  x242 &  x245 &  x248 &  x251 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x293 &  x296 &  x299 &  x305 &  x308 &  x314 &  x317 &  x320 &  x323 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x350 &  x356 &  x368 &  x374 &  x377 &  x380 &  x392 &  x395 &  x398 &  x407 &  x410 &  x416 &  x428 &  x431 &  x434 &  x442 &  x443 &  x446 &  x449 &  x455 &  x461 &  x464 &  x467 &  x470 &  x473 &  x479 &  x482 &  x488 &  x494 &  x500 &  x503 &  x506 &  x508 &  x509 &  x515 &  x518 &  x530 &  x533 &  x539 &  x542 &  x545 &  x547 &  x551 &  x554 &  x569 &  x572 &  x578 &  x581 &  x584 &  x586 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x617 &  x620 &  x623 &  x625 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x671 &  x674 &  x677 &  x695 &  x698 &  x701 &  x703 &  x704 &  x710 &  x719 &  x722 &  x725 &  x728 &  x731 &  x740 &  x742 &  x743 &  x749 &  x752 &  x755 &  x758 &  x761 &  x767 &  x773 &  x776 &  x779 &  x785 &  x794 &  x796 &  x800 &  x803 &  x806 &  x809 &  x815 &  x821 &  x827 &  x830 &  x834 &  x835 &  x839 &  x845 &  x854 &  x857 &  x860 &  x866 &  x869 &  x874 &  x884 &  x890 &  x893 &  x905 &  x908 &  x913 &  x914 &  x920 &  x923 &  x926 &  x932 &  x938 &  x947 &  x952 &  x956 &  x968 &  x971 &  x974 &  x980 &  x983 &  x986 &  x991 &  x992 &  x1010 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1052 &  x1055 &  x1061 &  x1067 &  x1070 &  x1073 &  x1085 &  x1091 &  x1094 &  x1100 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x354 & ~x393 & ~x513 & ~x552 & ~x831 & ~x870 & ~x978;
assign c7244 =  x5 &  x11 &  x14 &  x17 &  x23 &  x26 &  x32 &  x35 &  x38 &  x44 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x77 &  x83 &  x86 &  x92 &  x101 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x134 &  x137 &  x140 &  x143 &  x155 &  x158 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x191 &  x194 &  x203 &  x206 &  x212 &  x224 &  x227 &  x233 &  x239 &  x242 &  x245 &  x251 &  x257 &  x259 &  x266 &  x275 &  x290 &  x298 &  x299 &  x302 &  x305 &  x314 &  x317 &  x323 &  x326 &  x332 &  x337 &  x338 &  x344 &  x347 &  x353 &  x362 &  x371 &  x376 &  x380 &  x386 &  x404 &  x406 &  x416 &  x425 &  x437 &  x440 &  x446 &  x452 &  x455 &  x467 &  x470 &  x476 &  x485 &  x491 &  x500 &  x503 &  x512 &  x536 &  x545 &  x551 &  x563 &  x566 &  x575 &  x578 &  x581 &  x584 &  x587 &  x593 &  x598 &  x602 &  x605 &  x608 &  x617 &  x632 &  x635 &  x638 &  x640 &  x641 &  x644 &  x650 &  x665 &  x668 &  x674 &  x683 &  x686 &  x695 &  x707 &  x713 &  x716 &  x719 &  x728 &  x734 &  x740 &  x749 &  x752 &  x758 &  x761 &  x764 &  x767 &  x776 &  x779 &  x781 &  x791 &  x794 &  x806 &  x815 &  x820 &  x821 &  x824 &  x830 &  x833 &  x836 &  x839 &  x851 &  x854 &  x857 &  x859 &  x869 &  x872 &  x878 &  x881 &  x890 &  x896 &  x905 &  x923 &  x926 &  x935 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x962 &  x965 &  x976 &  x977 &  x983 &  x991 &  x992 &  x998 &  x1007 &  x1010 &  x1016 &  x1022 &  x1028 &  x1029 &  x1034 &  x1040 &  x1054 &  x1055 &  x1061 &  x1070 &  x1075 &  x1076 &  x1079 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1124 &  x1127 &  x1130 & ~x354 & ~x393 & ~x1095;
assign c7246 =  x8 &  x11 &  x14 &  x17 &  x23 &  x29 &  x32 &  x35 &  x38 &  x41 &  x47 &  x50 &  x53 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x83 &  x92 &  x95 &  x98 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x131 &  x134 &  x137 &  x146 &  x149 &  x155 &  x164 &  x170 &  x173 &  x176 &  x182 &  x185 &  x188 &  x194 &  x197 &  x200 &  x203 &  x209 &  x218 &  x221 &  x224 &  x227 &  x236 &  x248 &  x251 &  x254 &  x260 &  x266 &  x269 &  x274 &  x278 &  x281 &  x290 &  x293 &  x302 &  x311 &  x313 &  x314 &  x317 &  x320 &  x323 &  x332 &  x335 &  x338 &  x344 &  x347 &  x353 &  x356 &  x362 &  x365 &  x368 &  x377 &  x383 &  x386 &  x391 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x443 &  x446 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x476 &  x482 &  x488 &  x491 &  x497 &  x500 &  x509 &  x515 &  x521 &  x524 &  x527 &  x530 &  x536 &  x539 &  x541 &  x545 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x580 &  x581 &  x590 &  x593 &  x596 &  x605 &  x614 &  x617 &  x620 &  x623 &  x626 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x656 &  x658 &  x659 &  x662 &  x668 &  x670 &  x671 &  x674 &  x677 &  x680 &  x683 &  x692 &  x697 &  x701 &  x707 &  x709 &  x710 &  x713 &  x719 &  x722 &  x724 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x815 &  x827 &  x830 &  x836 &  x842 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x875 &  x878 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x932 &  x938 &  x944 &  x947 &  x950 &  x956 &  x965 &  x968 &  x971 &  x977 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1010 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1052 &  x1061 &  x1064 &  x1070 &  x1073 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1121 &  x1124 &  x1127 &  x1130 & ~x318 & ~x336 & ~x348 & ~x369 & ~x447 & ~x588 & ~x627 & ~x666 & ~x744 & ~x783 & ~x822;
assign c7248 =  x2 &  x5 &  x11 &  x17 &  x20 &  x26 &  x29 &  x32 &  x35 &  x38 &  x44 &  x50 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x236 &  x239 &  x245 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x338 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x413 &  x416 &  x425 &  x428 &  x431 &  x437 &  x438 &  x439 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x478 &  x479 &  x482 &  x485 &  x488 &  x491 &  x497 &  x500 &  x503 &  x509 &  x512 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x547 &  x548 &  x551 &  x554 &  x560 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x584 &  x587 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x614 &  x617 &  x620 &  x623 &  x625 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x650 &  x653 &  x656 &  x659 &  x662 &  x664 &  x665 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x779 &  x782 &  x785 &  x788 &  x794 &  x797 &  x800 &  x803 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x845 &  x851 &  x854 &  x857 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x892 &  x893 &  x896 &  x899 &  x902 &  x911 &  x914 &  x919 &  x923 &  x925 &  x926 &  x929 &  x931 &  x935 &  x938 &  x944 &  x950 &  x953 &  x958 &  x959 &  x964 &  x968 &  x970 &  x971 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1130 & ~x513 & ~x609 & ~x822 & ~x900 & ~x939 & ~x960;
assign c7250 =  x5 &  x8 &  x11 &  x17 &  x20 &  x29 &  x32 &  x35 &  x47 &  x50 &  x53 &  x71 &  x74 &  x77 &  x80 &  x83 &  x89 &  x91 &  x92 &  x98 &  x101 &  x110 &  x116 &  x119 &  x122 &  x128 &  x131 &  x137 &  x146 &  x152 &  x155 &  x158 &  x161 &  x164 &  x170 &  x173 &  x179 &  x182 &  x185 &  x191 &  x197 &  x200 &  x212 &  x218 &  x221 &  x230 &  x233 &  x236 &  x242 &  x245 &  x248 &  x254 &  x257 &  x260 &  x263 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x290 &  x296 &  x299 &  x308 &  x311 &  x313 &  x317 &  x320 &  x323 &  x326 &  x335 &  x338 &  x341 &  x344 &  x347 &  x352 &  x356 &  x359 &  x365 &  x377 &  x380 &  x383 &  x389 &  x392 &  x401 &  x404 &  x410 &  x416 &  x422 &  x425 &  x428 &  x430 &  x434 &  x437 &  x440 &  x449 &  x455 &  x461 &  x469 &  x473 &  x476 &  x482 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x512 &  x515 &  x518 &  x521 &  x527 &  x530 &  x536 &  x542 &  x545 &  x548 &  x551 &  x562 &  x569 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x592 &  x593 &  x599 &  x601 &  x602 &  x605 &  x611 &  x614 &  x617 &  x620 &  x626 &  x629 &  x632 &  x640 &  x641 &  x644 &  x647 &  x650 &  x662 &  x665 &  x668 &  x674 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x710 &  x713 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x743 &  x746 &  x752 &  x758 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x812 &  x821 &  x824 &  x827 &  x830 &  x839 &  x842 &  x845 &  x851 &  x854 &  x860 &  x863 &  x875 &  x878 &  x896 &  x902 &  x905 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x995 &  x1001 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1037 &  x1043 &  x1046 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1079 &  x1088 &  x1091 &  x1094 &  x1100 &  x1109 &  x1118 &  x1127 & ~x369 & ~x408 & ~x588 & ~x589 & ~x627 & ~x628 & ~x666 & ~x667 & ~x705 & ~x744 & ~x783 & ~x1101;
assign c7252 =  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x32 &  x38 &  x41 &  x44 &  x47 &  x53 &  x59 &  x62 &  x65 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x107 &  x110 &  x113 &  x122 &  x131 &  x134 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x164 &  x167 &  x169 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x197 &  x200 &  x203 &  x208 &  x212 &  x215 &  x218 &  x221 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x254 &  x257 &  x260 &  x263 &  x272 &  x278 &  x284 &  x290 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x326 &  x332 &  x338 &  x341 &  x347 &  x350 &  x353 &  x359 &  x362 &  x365 &  x371 &  x374 &  x380 &  x383 &  x392 &  x395 &  x401 &  x403 &  x404 &  x407 &  x410 &  x416 &  x422 &  x428 &  x431 &  x434 &  x437 &  x440 &  x442 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x467 &  x470 &  x476 &  x479 &  x482 &  x485 &  x491 &  x494 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x560 &  x566 &  x569 &  x578 &  x581 &  x584 &  x590 &  x593 &  x596 &  x599 &  x602 &  x608 &  x611 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x638 &  x641 &  x647 &  x650 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x698 &  x707 &  x710 &  x713 &  x719 &  x722 &  x728 &  x737 &  x740 &  x743 &  x752 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x800 &  x803 &  x806 &  x815 &  x818 &  x830 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x896 &  x899 &  x902 &  x905 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x950 &  x953 &  x956 &  x959 &  x965 &  x968 &  x974 &  x977 &  x983 &  x986 &  x989 &  x998 &  x1001 &  x1004 &  x1007 &  x1019 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1079 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x0 & ~x27 & ~x33 & ~x39 & ~x72 & ~x105 & ~x111 & ~x117 & ~x144 & ~x156 & ~x189 & ~x228 & ~x267 & ~x411 & ~x450 & ~x489 & ~x744 & ~x783 & ~x822;
assign c7254 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x35 &  x38 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x107 &  x110 &  x113 &  x116 &  x122 &  x125 &  x131 &  x137 &  x140 &  x146 &  x149 &  x155 &  x158 &  x161 &  x167 &  x170 &  x176 &  x179 &  x182 &  x185 &  x188 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x218 &  x221 &  x224 &  x227 &  x230 &  x245 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x308 &  x311 &  x314 &  x323 &  x329 &  x332 &  x338 &  x341 &  x344 &  x347 &  x353 &  x356 &  x365 &  x368 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x404 &  x407 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x446 &  x449 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x476 &  x482 &  x485 &  x488 &  x491 &  x497 &  x500 &  x503 &  x509 &  x512 &  x515 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x566 &  x569 &  x575 &  x578 &  x581 &  x584 &  x587 &  x593 &  x596 &  x602 &  x611 &  x614 &  x617 &  x620 &  x623 &  x629 &  x638 &  x641 &  x647 &  x650 &  x659 &  x665 &  x668 &  x674 &  x677 &  x680 &  x683 &  x686 &  x695 &  x704 &  x707 &  x710 &  x713 &  x716 &  x725 &  x731 &  x734 &  x737 &  x740 &  x743 &  x749 &  x752 &  x755 &  x761 &  x767 &  x770 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x851 &  x854 &  x857 &  x860 &  x866 &  x869 &  x872 &  x875 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x902 &  x905 &  x908 &  x911 &  x920 &  x923 &  x929 &  x932 &  x935 &  x938 &  x941 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x968 &  x971 &  x974 &  x980 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1100 &  x1103 &  x1115 &  x1127 &  x1130 & ~x315 & ~x354 & ~x393 & ~x432 & ~x471 & ~x867 & ~x960 & ~x984 & ~x1011 & ~x1023 & ~x1024 & ~x1056 & ~x1062 & ~x1063 & ~x1095 & ~x1102;
assign c7256 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x140 &  x143 &  x146 &  x149 &  x152 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x274 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x305 &  x308 &  x313 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x470 &  x473 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x523 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x541 &  x542 &  x545 &  x551 &  x554 &  x557 &  x560 &  x562 &  x566 &  x568 &  x569 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x601 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x626 &  x629 &  x632 &  x635 &  x638 &  x640 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x718 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x896 &  x899 &  x902 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1049 &  x1052 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x123 & ~x162 & ~x201 & ~x202 & ~x447 & ~x525 & ~x549 & ~x564 & ~x588 & ~x589 & ~x627 & ~x628 & ~x666 & ~x705 & ~x744 & ~x783 & ~x822 & ~x861 & ~x1101;
assign c7258 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x253 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x292 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x317 &  x320 &  x323 &  x325 &  x326 &  x329 &  x331 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x370 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x401 &  x404 &  x407 &  x409 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x556 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x590 &  x593 &  x594 &  x595 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x634 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x673 &  x674 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x983 &  x986 &  x989 &  x992 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x39 & ~x822 & ~x861 & ~x900;
assign c7260 =  x2 &  x5 &  x11 &  x14 &  x20 &  x23 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x80 &  x83 &  x86 &  x89 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x116 &  x119 &  x122 &  x128 &  x134 &  x137 &  x140 &  x146 &  x149 &  x155 &  x158 &  x161 &  x164 &  x167 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x284 &  x287 &  x290 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x317 &  x320 &  x323 &  x325 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x347 &  x350 &  x353 &  x359 &  x362 &  x364 &  x368 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x403 &  x407 &  x410 &  x413 &  x419 &  x422 &  x425 &  x428 &  x431 &  x437 &  x440 &  x442 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x506 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x980 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x78 & ~x117 & ~x156 & ~x228 & ~x345 & ~x384 & ~x423 & ~x450 & ~x513 & ~x837 & ~x876;
assign c7262 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x176 &  x179 &  x182 &  x185 &  x188 &  x194 &  x197 &  x200 &  x203 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x233 &  x236 &  x239 &  x245 &  x248 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x395 &  x398 &  x404 &  x407 &  x413 &  x416 &  x422 &  x425 &  x428 &  x434 &  x440 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x470 &  x473 &  x482 &  x485 &  x491 &  x494 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x551 &  x554 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x659 &  x662 &  x665 &  x668 &  x674 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x701 &  x704 &  x707 &  x710 &  x716 &  x719 &  x722 &  x725 &  x728 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x758 &  x761 &  x764 &  x770 &  x773 &  x776 &  x779 &  x781 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x820 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x857 &  x858 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x896 &  x897 &  x898 &  x899 &  x902 &  x905 &  x908 &  x911 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x936 &  x937 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x975 &  x976 &  x977 &  x980 &  x986 &  x989 &  x991 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1015 &  x1016 &  x1019 &  x1022 &  x1025 &  x1030 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1053 &  x1054 &  x1055 &  x1058 &  x1061 &  x1064 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1092 &  x1093 &  x1100 &  x1103 &  x1106 &  x1108 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x195 & ~x234 & ~x921 & ~x960 & ~x1056 & ~x1095;
assign c7264 =  x2 &  x5 &  x8 &  x14 &  x17 &  x23 &  x26 &  x41 &  x44 &  x49 &  x53 &  x56 &  x59 &  x65 &  x68 &  x71 &  x77 &  x89 &  x92 &  x95 &  x110 &  x118 &  x122 &  x125 &  x127 &  x128 &  x131 &  x134 &  x143 &  x146 &  x149 &  x161 &  x176 &  x182 &  x185 &  x188 &  x191 &  x200 &  x203 &  x206 &  x212 &  x230 &  x233 &  x245 &  x251 &  x254 &  x257 &  x269 &  x278 &  x284 &  x287 &  x293 &  x296 &  x299 &  x302 &  x311 &  x317 &  x323 &  x329 &  x338 &  x341 &  x347 &  x356 &  x362 &  x367 &  x368 &  x377 &  x380 &  x386 &  x389 &  x392 &  x398 &  x401 &  x406 &  x407 &  x428 &  x431 &  x437 &  x443 &  x445 &  x446 &  x455 &  x461 &  x464 &  x467 &  x473 &  x476 &  x479 &  x482 &  x484 &  x491 &  x514 &  x518 &  x521 &  x524 &  x527 &  x530 &  x542 &  x553 &  x560 &  x566 &  x578 &  x584 &  x587 &  x593 &  x611 &  x617 &  x626 &  x629 &  x635 &  x638 &  x644 &  x650 &  x656 &  x659 &  x668 &  x671 &  x677 &  x680 &  x683 &  x685 &  x692 &  x695 &  x707 &  x713 &  x718 &  x719 &  x722 &  x728 &  x731 &  x734 &  x740 &  x743 &  x746 &  x749 &  x752 &  x764 &  x767 &  x782 &  x785 &  x791 &  x794 &  x796 &  x797 &  x800 &  x803 &  x806 &  x815 &  x824 &  x827 &  x830 &  x836 &  x839 &  x851 &  x854 &  x866 &  x869 &  x872 &  x881 &  x893 &  x896 &  x899 &  x902 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x941 &  x953 &  x956 &  x959 &  x962 &  x971 &  x977 &  x983 &  x986 &  x989 &  x992 &  x998 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1046 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1088 &  x1091 &  x1097 &  x1103 &  x1112 &  x1130 & ~x393 & ~x666 & ~x702 & ~x705 & ~x741 & ~x744 & ~x780 & ~x861;
assign c7266 =  x2 &  x5 &  x8 &  x20 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x53 &  x59 &  x62 &  x65 &  x68 &  x74 &  x77 &  x83 &  x87 &  x88 &  x89 &  x95 &  x98 &  x101 &  x104 &  x107 &  x113 &  x118 &  x119 &  x128 &  x134 &  x149 &  x152 &  x155 &  x158 &  x161 &  x167 &  x173 &  x176 &  x179 &  x185 &  x188 &  x195 &  x196 &  x203 &  x206 &  x209 &  x212 &  x218 &  x224 &  x227 &  x230 &  x234 &  x236 &  x239 &  x242 &  x245 &  x248 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x274 &  x275 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x302 &  x311 &  x313 &  x317 &  x320 &  x323 &  x329 &  x335 &  x338 &  x347 &  x350 &  x352 &  x353 &  x356 &  x365 &  x371 &  x374 &  x377 &  x380 &  x383 &  x389 &  x391 &  x398 &  x407 &  x410 &  x419 &  x422 &  x428 &  x431 &  x434 &  x440 &  x443 &  x449 &  x452 &  x455 &  x458 &  x464 &  x470 &  x473 &  x475 &  x479 &  x485 &  x491 &  x494 &  x496 &  x497 &  x500 &  x503 &  x515 &  x518 &  x521 &  x527 &  x533 &  x536 &  x539 &  x542 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x596 &  x599 &  x602 &  x605 &  x617 &  x620 &  x626 &  x629 &  x632 &  x641 &  x644 &  x647 &  x656 &  x659 &  x662 &  x665 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x692 &  x695 &  x698 &  x701 &  x707 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x737 &  x740 &  x746 &  x752 &  x758 &  x761 &  x764 &  x767 &  x776 &  x779 &  x788 &  x791 &  x794 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x857 &  x860 &  x863 &  x881 &  x887 &  x890 &  x893 &  x905 &  x908 &  x914 &  x917 &  x920 &  x926 &  x932 &  x935 &  x938 &  x941 &  x947 &  x950 &  x953 &  x956 &  x959 &  x965 &  x968 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1010 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1043 &  x1049 &  x1052 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1085 &  x1091 &  x1094 &  x1100 &  x1103 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 & ~x180 & ~x219 & ~x220 & ~x297 & ~x433 & ~x471 & ~x510 & ~x588 & ~x666;
assign c7268 =  x2 &  x5 &  x8 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x308 &  x314 &  x317 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x476 &  x479 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x590 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x703 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x742 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x859 &  x860 &  x863 &  x866 &  x869 &  x872 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x898 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x935 &  x937 &  x938 &  x941 &  x944 &  x947 &  x950 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x976 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1007 &  x1009 &  x1013 &  x1015 &  x1016 &  x1019 &  x1022 &  x1025 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1048 &  x1049 &  x1052 &  x1054 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1087 &  x1091 &  x1093 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x276 & ~x315 & ~x354 & ~x393 & ~x432 & ~x471 & ~x510 & ~x549 & ~x588 & ~x843 & ~x882 & ~x921 & ~x939 & ~x960 & ~x978 & ~x999 & ~x1017 & ~x1018 & ~x1038 & ~x1056 & ~x1057 & ~x1095 & ~x1122;
assign c7270 =  x5 &  x20 &  x26 &  x38 &  x41 &  x50 &  x62 &  x71 &  x74 &  x86 &  x98 &  x113 &  x134 &  x140 &  x146 &  x152 &  x164 &  x167 &  x170 &  x173 &  x182 &  x188 &  x191 &  x194 &  x200 &  x206 &  x212 &  x224 &  x242 &  x245 &  x254 &  x260 &  x263 &  x275 &  x278 &  x287 &  x290 &  x293 &  x302 &  x308 &  x317 &  x322 &  x332 &  x338 &  x341 &  x344 &  x350 &  x362 &  x374 &  x383 &  x389 &  x398 &  x401 &  x406 &  x413 &  x416 &  x440 &  x443 &  x446 &  x458 &  x464 &  x476 &  x482 &  x485 &  x494 &  x506 &  x508 &  x512 &  x524 &  x530 &  x551 &  x554 &  x563 &  x572 &  x578 &  x581 &  x593 &  x596 &  x602 &  x605 &  x608 &  x623 &  x635 &  x653 &  x671 &  x674 &  x695 &  x704 &  x710 &  x716 &  x737 &  x749 &  x755 &  x767 &  x779 &  x782 &  x794 &  x797 &  x803 &  x809 &  x815 &  x818 &  x839 &  x845 &  x848 &  x851 &  x857 &  x860 &  x863 &  x887 &  x890 &  x893 &  x902 &  x905 &  x911 &  x926 &  x932 &  x935 &  x941 &  x947 &  x965 &  x977 &  x980 &  x986 &  x989 &  x998 &  x1004 &  x1022 &  x1040 &  x1049 &  x1061 &  x1076 &  x1085 &  x1088 & ~x453 & ~x532 & ~x570 & ~x714 & ~x744 & ~x792 & ~x823 & ~x861 & ~x870 & ~x900 & ~x909;
assign c7272 =  x11 &  x14 &  x17 &  x23 &  x32 &  x44 &  x47 &  x50 &  x56 &  x59 &  x62 &  x65 &  x71 &  x74 &  x77 &  x86 &  x89 &  x95 &  x104 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x137 &  x140 &  x143 &  x146 &  x152 &  x170 &  x173 &  x179 &  x185 &  x191 &  x197 &  x200 &  x203 &  x215 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x257 &  x260 &  x263 &  x269 &  x272 &  x275 &  x281 &  x284 &  x296 &  x299 &  x305 &  x311 &  x314 &  x317 &  x320 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x362 &  x365 &  x371 &  x374 &  x382 &  x383 &  x386 &  x392 &  x395 &  x407 &  x410 &  x413 &  x421 &  x422 &  x425 &  x428 &  x431 &  x434 &  x437 &  x443 &  x446 &  x452 &  x458 &  x461 &  x464 &  x470 &  x476 &  x482 &  x485 &  x491 &  x494 &  x497 &  x499 &  x500 &  x503 &  x506 &  x512 &  x515 &  x518 &  x533 &  x539 &  x542 &  x548 &  x557 &  x559 &  x566 &  x569 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x620 &  x623 &  x632 &  x635 &  x637 &  x638 &  x640 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x668 &  x671 &  x679 &  x680 &  x686 &  x689 &  x698 &  x707 &  x710 &  x716 &  x725 &  x728 &  x734 &  x737 &  x740 &  x743 &  x746 &  x752 &  x755 &  x761 &  x767 &  x770 &  x779 &  x782 &  x790 &  x791 &  x797 &  x803 &  x809 &  x812 &  x818 &  x820 &  x821 &  x830 &  x836 &  x839 &  x842 &  x845 &  x851 &  x854 &  x860 &  x866 &  x872 &  x878 &  x881 &  x884 &  x887 &  x893 &  x896 &  x898 &  x902 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x937 &  x944 &  x947 &  x950 &  x953 &  x956 &  x962 &  x965 &  x968 &  x974 &  x976 &  x977 &  x980 &  x986 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1015 &  x1016 &  x1022 &  x1028 &  x1031 &  x1037 &  x1040 &  x1043 &  x1049 &  x1052 &  x1054 &  x1055 &  x1058 &  x1061 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1091 &  x1093 &  x1094 &  x1108 &  x1118 &  x1124 & ~x312 & ~x351 & ~x390 & ~x429 & ~x432 & ~x888;
assign c7274 =  x5 &  x8 &  x11 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x269 &  x275 &  x281 &  x284 &  x286 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x314 &  x317 &  x323 &  x325 &  x326 &  x329 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x353 &  x356 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x391 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x419 &  x422 &  x425 &  x428 &  x430 &  x431 &  x440 &  x443 &  x446 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x469 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x494 &  x497 &  x503 &  x506 &  x508 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x605 &  x608 &  x611 &  x614 &  x623 &  x626 &  x629 &  x632 &  x638 &  x641 &  x644 &  x646 &  x647 &  x650 &  x653 &  x656 &  x665 &  x668 &  x671 &  x674 &  x677 &  x679 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x718 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x785 &  x788 &  x791 &  x796 &  x800 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x932 &  x935 &  x938 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1046 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1076 &  x1079 &  x1082 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x588 & ~x627 & ~x628 & ~x666 & ~x667 & ~x705 & ~x783 & ~x822 & ~x936 & ~x975 & ~x1014 & ~x1053;
assign c7276 =  x5 &  x8 &  x11 &  x14 &  x32 &  x35 &  x44 &  x47 &  x50 &  x53 &  x56 &  x62 &  x65 &  x74 &  x77 &  x80 &  x95 &  x98 &  x110 &  x116 &  x125 &  x131 &  x134 &  x143 &  x146 &  x149 &  x158 &  x164 &  x173 &  x176 &  x182 &  x185 &  x188 &  x191 &  x194 &  x203 &  x209 &  x215 &  x218 &  x221 &  x224 &  x242 &  x248 &  x251 &  x259 &  x265 &  x272 &  x278 &  x281 &  x284 &  x287 &  x293 &  x304 &  x305 &  x308 &  x311 &  x317 &  x337 &  x350 &  x353 &  x356 &  x362 &  x365 &  x374 &  x377 &  x380 &  x383 &  x398 &  x401 &  x404 &  x413 &  x419 &  x422 &  x425 &  x428 &  x434 &  x446 &  x458 &  x470 &  x476 &  x479 &  x482 &  x491 &  x500 &  x506 &  x512 &  x521 &  x524 &  x527 &  x530 &  x539 &  x542 &  x545 &  x548 &  x551 &  x556 &  x559 &  x560 &  x563 &  x566 &  x572 &  x575 &  x584 &  x595 &  x596 &  x598 &  x599 &  x602 &  x605 &  x608 &  x626 &  x629 &  x632 &  x635 &  x641 &  x650 &  x653 &  x662 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x692 &  x698 &  x710 &  x713 &  x716 &  x722 &  x725 &  x728 &  x734 &  x737 &  x743 &  x752 &  x755 &  x758 &  x761 &  x776 &  x779 &  x781 &  x788 &  x794 &  x797 &  x800 &  x809 &  x812 &  x818 &  x820 &  x821 &  x836 &  x839 &  x845 &  x854 &  x857 &  x872 &  x884 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x914 &  x926 &  x944 &  x947 &  x956 &  x959 &  x962 &  x971 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1010 &  x1013 &  x1019 &  x1022 &  x1034 &  x1037 &  x1046 &  x1055 &  x1079 &  x1091 &  x1097 &  x1103 &  x1115 &  x1124 & ~x273 & ~x312 & ~x393 & ~x471 & ~x630 & ~x669 & ~x978 & ~x1017;
assign c7278 =  x2 &  x11 &  x14 &  x23 &  x29 &  x41 &  x50 &  x56 &  x68 &  x80 &  x83 &  x86 &  x95 &  x101 &  x107 &  x125 &  x134 &  x140 &  x158 &  x167 &  x176 &  x179 &  x182 &  x194 &  x206 &  x209 &  x215 &  x224 &  x227 &  x233 &  x245 &  x257 &  x269 &  x275 &  x284 &  x305 &  x311 &  x320 &  x329 &  x332 &  x335 &  x338 &  x344 &  x347 &  x359 &  x377 &  x383 &  x386 &  x392 &  x398 &  x403 &  x406 &  x410 &  x419 &  x422 &  x428 &  x446 &  x449 &  x461 &  x470 &  x481 &  x488 &  x494 &  x506 &  x512 &  x533 &  x536 &  x557 &  x559 &  x572 &  x575 &  x586 &  x605 &  x611 &  x625 &  x629 &  x638 &  x647 &  x659 &  x664 &  x668 &  x692 &  x704 &  x713 &  x716 &  x758 &  x764 &  x773 &  x779 &  x797 &  x806 &  x815 &  x824 &  x827 &  x830 &  x833 &  x836 &  x851 &  x853 &  x854 &  x860 &  x884 &  x890 &  x892 &  x905 &  x911 &  x913 &  x920 &  x929 &  x944 &  x953 &  x958 &  x977 &  x980 &  x992 &  x1001 &  x1004 &  x1025 &  x1034 &  x1040 &  x1061 &  x1070 &  x1073 &  x1079 &  x1088 &  x1091 &  x1094 &  x1100 &  x1112 &  x1121 & ~x861 & ~x900 & ~x939 & ~x940;
assign c7280 =  x32 &  x47 &  x50 &  x56 &  x62 &  x89 &  x107 &  x110 &  x170 &  x176 &  x179 &  x203 &  x221 &  x236 &  x239 &  x248 &  x275 &  x302 &  x314 &  x320 &  x323 &  x359 &  x382 &  x395 &  x413 &  x437 &  x446 &  x467 &  x473 &  x491 &  x506 &  x512 &  x515 &  x521 &  x539 &  x545 &  x572 &  x584 &  x611 &  x620 &  x665 &  x714 &  x767 &  x806 &  x827 &  x839 &  x842 &  x863 &  x866 &  x881 &  x908 &  x920 &  x923 &  x959 &  x968 &  x974 &  x980 &  x992 &  x1010 &  x1013 &  x1034 &  x1040 &  x1049 &  x1052 &  x1082 &  x1103 &  x1106 & ~x393 & ~x471 & ~x510 & ~x546 & ~x846 & ~x886;
assign c7282 =  x2 &  x5 &  x8 &  x11 &  x17 &  x20 &  x23 &  x26 &  x29 &  x38 &  x41 &  x44 &  x47 &  x50 &  x56 &  x59 &  x62 &  x65 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x95 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x125 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x155 &  x158 &  x164 &  x165 &  x166 &  x167 &  x170 &  x173 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x196 &  x197 &  x200 &  x203 &  x205 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x227 &  x233 &  x235 &  x236 &  x239 &  x242 &  x245 &  x251 &  x257 &  x260 &  x263 &  x266 &  x274 &  x275 &  x278 &  x281 &  x287 &  x290 &  x293 &  x296 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x332 &  x335 &  x338 &  x341 &  x344 &  x347 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x386 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x413 &  x416 &  x419 &  x425 &  x428 &  x431 &  x434 &  x437 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x470 &  x473 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x530 &  x533 &  x536 &  x539 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x569 &  x575 &  x578 &  x580 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x613 &  x614 &  x620 &  x623 &  x626 &  x629 &  x632 &  x638 &  x641 &  x644 &  x647 &  x650 &  x652 &  x656 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x734 &  x737 &  x743 &  x749 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x803 &  x806 &  x809 &  x812 &  x818 &  x827 &  x833 &  x836 &  x839 &  x845 &  x848 &  x854 &  x857 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x902 &  x908 &  x911 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x986 &  x989 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1016 &  x1019 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1079 &  x1082 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x180 & ~x510 & ~x549 & ~x588 & ~x609 & ~x627 & ~x648 & ~x666 & ~x960;
assign c7284 =  x2 &  x11 &  x14 &  x17 &  x20 &  x32 &  x35 &  x38 &  x41 &  x47 &  x53 &  x56 &  x59 &  x62 &  x65 &  x68 &  x86 &  x107 &  x110 &  x122 &  x125 &  x128 &  x134 &  x146 &  x149 &  x152 &  x158 &  x170 &  x176 &  x185 &  x191 &  x203 &  x215 &  x221 &  x224 &  x230 &  x233 &  x236 &  x239 &  x242 &  x248 &  x251 &  x266 &  x272 &  x278 &  x287 &  x296 &  x308 &  x311 &  x326 &  x332 &  x338 &  x347 &  x353 &  x359 &  x371 &  x377 &  x386 &  x389 &  x398 &  x404 &  x407 &  x416 &  x422 &  x434 &  x437 &  x443 &  x455 &  x464 &  x476 &  x479 &  x482 &  x485 &  x488 &  x500 &  x503 &  x509 &  x512 &  x524 &  x527 &  x536 &  x539 &  x551 &  x587 &  x590 &  x593 &  x596 &  x599 &  x620 &  x623 &  x629 &  x634 &  x644 &  x653 &  x656 &  x659 &  x662 &  x680 &  x683 &  x686 &  x695 &  x698 &  x704 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x743 &  x749 &  x770 &  x785 &  x791 &  x800 &  x803 &  x818 &  x821 &  x836 &  x842 &  x857 &  x866 &  x869 &  x884 &  x911 &  x917 &  x947 &  x956 &  x962 &  x995 &  x1016 &  x1022 &  x1031 &  x1043 &  x1046 &  x1052 &  x1064 &  x1073 &  x1085 &  x1091 &  x1103 &  x1124 &  x1126 & ~x799 & ~x825 & ~x837 & ~x882 & ~x960 & ~x999 & ~x1011;
assign c7286 =  x5 &  x11 &  x14 &  x17 &  x23 &  x26 &  x35 &  x38 &  x41 &  x50 &  x59 &  x62 &  x71 &  x74 &  x80 &  x86 &  x89 &  x92 &  x98 &  x104 &  x107 &  x110 &  x122 &  x125 &  x128 &  x131 &  x137 &  x140 &  x143 &  x146 &  x152 &  x155 &  x164 &  x165 &  x166 &  x170 &  x176 &  x179 &  x182 &  x185 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x245 &  x248 &  x251 &  x254 &  x263 &  x266 &  x269 &  x272 &  x274 &  x275 &  x286 &  x287 &  x290 &  x293 &  x299 &  x305 &  x308 &  x314 &  x317 &  x320 &  x323 &  x325 &  x326 &  x332 &  x335 &  x344 &  x350 &  x352 &  x353 &  x356 &  x359 &  x368 &  x371 &  x374 &  x380 &  x383 &  x389 &  x391 &  x392 &  x395 &  x398 &  x407 &  x410 &  x416 &  x419 &  x422 &  x425 &  x428 &  x431 &  x437 &  x440 &  x446 &  x449 &  x455 &  x458 &  x464 &  x476 &  x482 &  x494 &  x500 &  x502 &  x503 &  x506 &  x509 &  x512 &  x515 &  x524 &  x527 &  x530 &  x533 &  x536 &  x539 &  x541 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x566 &  x569 &  x572 &  x580 &  x581 &  x587 &  x590 &  x593 &  x596 &  x599 &  x605 &  x611 &  x620 &  x623 &  x626 &  x635 &  x638 &  x641 &  x644 &  x650 &  x659 &  x662 &  x665 &  x668 &  x674 &  x677 &  x689 &  x695 &  x698 &  x701 &  x704 &  x707 &  x713 &  x719 &  x722 &  x725 &  x728 &  x731 &  x737 &  x740 &  x752 &  x761 &  x770 &  x773 &  x776 &  x779 &  x785 &  x791 &  x794 &  x797 &  x803 &  x809 &  x812 &  x815 &  x818 &  x821 &  x827 &  x833 &  x842 &  x848 &  x860 &  x875 &  x878 &  x884 &  x890 &  x893 &  x896 &  x899 &  x902 &  x905 &  x908 &  x911 &  x917 &  x920 &  x923 &  x929 &  x935 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1037 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1067 &  x1070 &  x1076 &  x1079 &  x1082 &  x1088 &  x1091 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1115 &  x1118 &  x1121 &  x1124 & ~x271 & ~x297 & ~x588 & ~x627 & ~x666 & ~x744 & ~x822;
assign c7288 =  x2 &  x5 &  x8 &  x10 &  x11 &  x17 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x47 &  x49 &  x53 &  x59 &  x62 &  x65 &  x68 &  x74 &  x77 &  x80 &  x83 &  x86 &  x88 &  x89 &  x95 &  x101 &  x104 &  x107 &  x110 &  x116 &  x118 &  x119 &  x122 &  x125 &  x128 &  x134 &  x140 &  x143 &  x146 &  x149 &  x152 &  x156 &  x158 &  x161 &  x164 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x195 &  x196 &  x199 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x227 &  x230 &  x235 &  x242 &  x245 &  x248 &  x251 &  x254 &  x260 &  x263 &  x266 &  x269 &  x272 &  x274 &  x275 &  x278 &  x281 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x313 &  x314 &  x317 &  x320 &  x323 &  x326 &  x335 &  x338 &  x341 &  x344 &  x350 &  x353 &  x356 &  x362 &  x365 &  x371 &  x374 &  x377 &  x383 &  x385 &  x386 &  x389 &  x392 &  x395 &  x398 &  x404 &  x410 &  x413 &  x416 &  x419 &  x424 &  x425 &  x428 &  x431 &  x434 &  x440 &  x443 &  x449 &  x452 &  x455 &  x458 &  x463 &  x464 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x494 &  x500 &  x503 &  x506 &  x509 &  x512 &  x518 &  x524 &  x527 &  x529 &  x533 &  x536 &  x539 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x562 &  x563 &  x566 &  x569 &  x575 &  x584 &  x590 &  x596 &  x599 &  x601 &  x605 &  x608 &  x611 &  x614 &  x617 &  x623 &  x626 &  x632 &  x641 &  x644 &  x647 &  x650 &  x653 &  x659 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x713 &  x716 &  x719 &  x722 &  x731 &  x734 &  x737 &  x743 &  x752 &  x755 &  x761 &  x764 &  x770 &  x773 &  x776 &  x779 &  x782 &  x791 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x872 &  x875 &  x878 &  x881 &  x890 &  x893 &  x899 &  x902 &  x905 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x944 &  x950 &  x953 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1022 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1058 &  x1061 &  x1070 &  x1076 &  x1079 &  x1082 &  x1094 &  x1097 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1130 & ~x84 & ~x162 & ~x219 & ~x258 & ~x297 & ~x471 & ~x472 & ~x511 & ~x588 & ~x627 & ~x819;
assign c7290 =  x2 &  x5 &  x10 &  x11 &  x14 &  x17 &  x26 &  x32 &  x38 &  x41 &  x44 &  x47 &  x49 &  x56 &  x59 &  x71 &  x74 &  x77 &  x79 &  x80 &  x83 &  x86 &  x88 &  x89 &  x95 &  x98 &  x101 &  x107 &  x110 &  x116 &  x118 &  x121 &  x125 &  x128 &  x134 &  x137 &  x140 &  x143 &  x146 &  x149 &  x155 &  x157 &  x158 &  x164 &  x167 &  x170 &  x176 &  x179 &  x188 &  x191 &  x196 &  x197 &  x200 &  x203 &  x209 &  x218 &  x224 &  x230 &  x235 &  x239 &  x245 &  x248 &  x251 &  x254 &  x257 &  x263 &  x266 &  x269 &  x272 &  x274 &  x275 &  x278 &  x281 &  x290 &  x293 &  x299 &  x302 &  x305 &  x311 &  x314 &  x323 &  x329 &  x332 &  x338 &  x341 &  x347 &  x356 &  x359 &  x365 &  x368 &  x371 &  x374 &  x377 &  x383 &  x386 &  x395 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x425 &  x428 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x457 &  x458 &  x470 &  x473 &  x476 &  x479 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x506 &  x512 &  x515 &  x518 &  x527 &  x536 &  x542 &  x545 &  x548 &  x551 &  x554 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x590 &  x599 &  x602 &  x608 &  x611 &  x617 &  x623 &  x626 &  x629 &  x635 &  x641 &  x644 &  x647 &  x650 &  x653 &  x662 &  x665 &  x668 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x688 &  x691 &  x695 &  x704 &  x710 &  x716 &  x722 &  x725 &  x728 &  x731 &  x734 &  x740 &  x743 &  x746 &  x749 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x782 &  x785 &  x788 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x836 &  x839 &  x842 &  x851 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x884 &  x887 &  x893 &  x899 &  x911 &  x914 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x950 &  x956 &  x959 &  x962 &  x965 &  x968 &  x974 &  x977 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1007 &  x1010 &  x1013 &  x1016 &  x1028 &  x1031 &  x1034 &  x1037 &  x1043 &  x1046 &  x1049 &  x1055 &  x1061 &  x1064 &  x1070 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1121 &  x1124 &  x1127 & ~x84 & ~x174 & ~x433 & ~x471 & ~x472 & ~x510 & ~x666 & ~x705 & ~x744 & ~x783 & ~x822;
assign c7292 =  x2 &  x5 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x62 &  x65 &  x71 &  x74 &  x77 &  x83 &  x86 &  x89 &  x95 &  x98 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x230 &  x233 &  x239 &  x242 &  x245 &  x248 &  x257 &  x260 &  x263 &  x269 &  x272 &  x275 &  x281 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x308 &  x311 &  x314 &  x317 &  x320 &  x323 &  x326 &  x329 &  x332 &  x341 &  x344 &  x347 &  x353 &  x356 &  x365 &  x371 &  x374 &  x380 &  x383 &  x389 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x413 &  x416 &  x422 &  x428 &  x431 &  x437 &  x439 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x467 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x542 &  x545 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x632 &  x638 &  x641 &  x644 &  x647 &  x653 &  x659 &  x662 &  x665 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x809 &  x812 &  x815 &  x818 &  x821 &  x824 &  x827 &  x830 &  x833 &  x836 &  x839 &  x845 &  x851 &  x854 &  x857 &  x860 &  x863 &  x866 &  x869 &  x872 &  x875 &  x878 &  x884 &  x887 &  x890 &  x893 &  x899 &  x902 &  x905 &  x911 &  x917 &  x920 &  x923 &  x929 &  x932 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x995 &  x998 &  x1007 &  x1010 &  x1013 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1115 &  x1121 &  x1124 &  x1127 &  x1130 & ~x78 & ~x117 & ~x195 & ~x306 & ~x315 & ~x345 & ~x699 & ~x744 & ~x783 & ~x822 & ~x823 & ~x861 & ~x900 & ~x939;
assign c7294 =  x8 &  x14 &  x29 &  x35 &  x47 &  x56 &  x68 &  x80 &  x83 &  x98 &  x113 &  x122 &  x128 &  x140 &  x146 &  x158 &  x179 &  x203 &  x209 &  x218 &  x236 &  x239 &  x245 &  x260 &  x269 &  x275 &  x278 &  x287 &  x299 &  x302 &  x308 &  x323 &  x326 &  x335 &  x338 &  x344 &  x362 &  x365 &  x380 &  x383 &  x395 &  x401 &  x410 &  x416 &  x422 &  x461 &  x473 &  x476 &  x482 &  x485 &  x503 &  x512 &  x518 &  x530 &  x545 &  x547 &  x551 &  x578 &  x581 &  x584 &  x599 &  x605 &  x614 &  x617 &  x623 &  x641 &  x653 &  x668 &  x671 &  x677 &  x680 &  x686 &  x704 &  x710 &  x719 &  x722 &  x734 &  x767 &  x785 &  x794 &  x809 &  x815 &  x821 &  x833 &  x851 &  x863 &  x869 &  x881 &  x893 &  x896 &  x899 &  x905 &  x929 &  x935 &  x941 &  x956 &  x1013 &  x1016 &  x1019 &  x1022 &  x1058 &  x1064 &  x1076 &  x1079 &  x1085 &  x1091 &  x1103 &  x1112 &  x1115 & ~x78 & ~x156 & ~x823 & ~x861 & ~x862 & ~x901 & ~x939 & ~x979 & ~x1018;
assign c7296 =  x2 &  x5 &  x11 &  x14 &  x17 &  x20 &  x23 &  x26 &  x29 &  x32 &  x35 &  x38 &  x41 &  x44 &  x47 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x74 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x98 &  x101 &  x104 &  x107 &  x110 &  x113 &  x116 &  x119 &  x122 &  x125 &  x128 &  x131 &  x137 &  x140 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x161 &  x164 &  x167 &  x170 &  x173 &  x176 &  x179 &  x182 &  x185 &  x188 &  x191 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x215 &  x218 &  x221 &  x224 &  x227 &  x230 &  x233 &  x236 &  x239 &  x242 &  x244 &  x245 &  x248 &  x251 &  x254 &  x257 &  x260 &  x263 &  x266 &  x269 &  x272 &  x275 &  x278 &  x281 &  x283 &  x284 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x308 &  x311 &  x314 &  x317 &  x321 &  x322 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x344 &  x347 &  x350 &  x353 &  x356 &  x359 &  x361 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x380 &  x386 &  x389 &  x391 &  x392 &  x395 &  x398 &  x401 &  x404 &  x407 &  x413 &  x419 &  x422 &  x425 &  x428 &  x430 &  x431 &  x437 &  x440 &  x443 &  x446 &  x449 &  x452 &  x455 &  x458 &  x461 &  x464 &  x467 &  x469 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x512 &  x515 &  x518 &  x521 &  x524 &  x527 &  x530 &  x533 &  x536 &  x542 &  x545 &  x548 &  x554 &  x557 &  x560 &  x563 &  x566 &  x569 &  x572 &  x575 &  x578 &  x581 &  x584 &  x587 &  x590 &  x593 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x617 &  x620 &  x623 &  x626 &  x629 &  x632 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x653 &  x656 &  x659 &  x662 &  x665 &  x668 &  x670 &  x671 &  x674 &  x677 &  x680 &  x683 &  x686 &  x689 &  x692 &  x695 &  x698 &  x701 &  x704 &  x707 &  x709 &  x710 &  x713 &  x716 &  x719 &  x722 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x748 &  x749 &  x752 &  x755 &  x758 &  x761 &  x763 &  x764 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x787 &  x788 &  x791 &  x794 &  x797 &  x800 &  x802 &  x806 &  x809 &  x812 &  x815 &  x818 &  x824 &  x826 &  x827 &  x830 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x863 &  x865 &  x866 &  x869 &  x872 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x896 &  x899 &  x905 &  x908 &  x911 &  x914 &  x917 &  x920 &  x923 &  x926 &  x929 &  x932 &  x935 &  x938 &  x941 &  x947 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x968 &  x971 &  x974 &  x977 &  x980 &  x983 &  x986 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1010 &  x1013 &  x1016 &  x1019 &  x1025 &  x1028 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1058 &  x1061 &  x1064 &  x1067 &  x1070 &  x1073 &  x1079 &  x1082 &  x1088 &  x1091 &  x1097 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1121 &  x1124 &  x1127 & ~x336 & ~x357 & ~x414 & ~x453 & ~x666 & ~x705 & ~x744 & ~x745 & ~x783 & ~x822 & ~x861;
assign c7298 =  x5 &  x14 &  x17 &  x29 &  x44 &  x47 &  x62 &  x65 &  x74 &  x77 &  x89 &  x92 &  x119 &  x122 &  x128 &  x131 &  x134 &  x137 &  x140 &  x143 &  x146 &  x164 &  x191 &  x203 &  x206 &  x209 &  x218 &  x224 &  x233 &  x236 &  x257 &  x293 &  x296 &  x299 &  x323 &  x347 &  x350 &  x371 &  x377 &  x395 &  x401 &  x416 &  x425 &  x434 &  x437 &  x452 &  x455 &  x464 &  x482 &  x485 &  x494 &  x497 &  x512 &  x515 &  x524 &  x527 &  x557 &  x560 &  x563 &  x590 &  x593 &  x611 &  x617 &  x620 &  x629 &  x632 &  x650 &  x656 &  x674 &  x683 &  x710 &  x728 &  x755 &  x761 &  x764 &  x773 &  x779 &  x782 &  x785 &  x806 &  x809 &  x815 &  x827 &  x851 &  x854 &  x863 &  x884 &  x902 &  x914 &  x926 &  x929 &  x941 &  x950 &  x962 &  x974 &  x977 &  x983 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1019 &  x1021 &  x1055 &  x1060 &  x1061 &  x1067 &  x1076 &  x1085 &  x1088 &  x1103 &  x1124 & ~x39 & ~x78 & ~x237 & ~x354 & ~x393 & ~x765 & ~x1018;
assign c71 =  x472 &  x511 &  x790 & ~x601;
assign c73 =  x2 &  x23 &  x62 &  x95 &  x191 &  x302 &  x305 &  x341 &  x355 &  x380 &  x398 &  x413 &  x464 &  x503 &  x515 &  x518 &  x527 &  x560 &  x578 &  x593 &  x602 &  x620 &  x623 &  x634 &  x656 &  x662 &  x692 &  x695 &  x704 &  x715 &  x718 &  x722 &  x743 &  x758 &  x773 &  x794 &  x853 &  x875 &  x934 &  x956 &  x1001 &  x1007 &  x1027 &  x1106 &  x1121 & ~x744 & ~x861;
assign c75 =  x50 &  x341 &  x374 &  x554 &  x745 &  x823 &  x1049 & ~x51 & ~x636 & ~x1098;
assign c77 =  x939 & ~x1108;
assign c79 =  x8 &  x53 &  x65 &  x68 &  x80 &  x104 &  x116 &  x122 &  x131 &  x134 &  x143 &  x152 &  x155 &  x158 &  x182 &  x200 &  x227 &  x236 &  x239 &  x248 &  x269 &  x273 &  x274 &  x278 &  x281 &  x299 &  x305 &  x313 &  x329 &  x350 &  x404 &  x416 &  x422 &  x434 &  x455 &  x473 &  x479 &  x482 &  x488 &  x500 &  x527 &  x530 &  x536 &  x539 &  x572 &  x602 &  x605 &  x623 &  x626 &  x641 &  x650 &  x653 &  x655 &  x656 &  x662 &  x668 &  x673 &  x683 &  x698 &  x722 &  x740 &  x758 &  x779 &  x794 &  x800 &  x809 &  x830 &  x851 &  x866 &  x887 &  x890 &  x902 &  x926 &  x938 &  x947 &  x950 &  x968 &  x977 &  x992 &  x995 &  x1001 &  x1022 &  x1028 &  x1037 &  x1049 &  x1052 &  x1055 &  x1058 &  x1064 &  x1067 &  x1085 &  x1088 &  x1094 &  x1097 &  x1100 &  x1130 & ~x168 & ~x207 & ~x246;
assign c711 =  x14 &  x47 &  x272 &  x314 &  x332 &  x353 &  x380 &  x398 &  x407 &  x502 &  x506 &  x554 &  x656 &  x701 &  x740 &  x761 &  x833 &  x848 &  x920 &  x953 &  x1004 &  x1018 &  x1043 &  x1057 &  x1076 &  x1118 & ~x87 & ~x282 & ~x726;
assign c713 =  x68 &  x83 &  x98 &  x355 &  x368 &  x389 &  x394 &  x754 &  x791 &  x799 &  x844 & ~x696;
assign c715 =  x586 &  x784 &  x979 &  x1058 & ~x195 & ~x198;
assign c717 =  x217 &  x784 &  x901 &  x1101 & ~x120;
assign c719 =  x297 &  x475 & ~x477 & ~x633 & ~x711;
assign c721 =  x155 &  x167 &  x230 &  x251 &  x344 &  x380 &  x473 &  x539 &  x617 &  x632 &  x680 &  x742 &  x803 &  x859 &  x905 &  x1025 &  x1057 &  x1102 & ~x360 & ~x549 & ~x588 & ~x660 & ~x777 & ~x804;
assign c723 =  x328 &  x939 & ~x235 & ~x313;
assign c725 =  x499 & ~x312 & ~x637;
assign c727 =  x391 &  x550 & ~x403;
assign c729 =  x17 &  x29 &  x35 &  x38 &  x44 &  x53 &  x71 &  x83 &  x86 &  x89 &  x95 &  x98 &  x101 &  x119 &  x134 &  x152 &  x173 &  x179 &  x182 &  x194 &  x203 &  x206 &  x209 &  x236 &  x269 &  x272 &  x277 &  x278 &  x287 &  x302 &  x316 &  x323 &  x326 &  x347 &  x353 &  x359 &  x368 &  x389 &  x392 &  x407 &  x410 &  x413 &  x419 &  x428 &  x437 &  x452 &  x461 &  x470 &  x494 &  x500 &  x518 &  x524 &  x530 &  x533 &  x539 &  x545 &  x557 &  x566 &  x578 &  x590 &  x595 &  x608 &  x614 &  x617 &  x620 &  x626 &  x644 &  x656 &  x676 &  x692 &  x695 &  x698 &  x704 &  x728 &  x731 &  x740 &  x752 &  x779 &  x796 &  x803 &  x842 &  x848 &  x899 &  x917 &  x935 &  x959 &  x968 &  x980 &  x983 &  x992 &  x1007 &  x1010 &  x1028 &  x1052 &  x1076 &  x1085 &  x1100 & ~x663 & ~x703;
assign c731 =  x112 &  x784 & ~x120 & ~x597;
assign c733 =  x13 &  x511 &  x838 & ~x405 & ~x858;
assign c735 =  x68 &  x215 &  x272 &  x320 &  x397 &  x569 &  x590 &  x664 &  x671 &  x680 &  x692 &  x707 &  x728 &  x797 &  x1010 & ~x159 & ~x477 & ~x516 & ~x603 & ~x837;
assign c737 =  x26 &  x92 &  x116 &  x341 &  x355 &  x365 &  x368 &  x394 &  x476 &  x524 &  x530 &  x566 &  x581 &  x668 &  x698 &  x715 &  x793 &  x797 &  x799 &  x806 &  x821 &  x844 &  x869 &  x914 & ~x735;
assign c739 =  x325 &  x442 &  x940 &  x1057 & ~x391 & ~x810 & ~x849;
assign c741 =  x1021 & ~x48 & ~x552 & ~x664;
assign c743 =  x169 &  x550 & ~x441 & ~x519 & ~x840;
assign c745 =  x29 &  x44 &  x92 &  x107 &  x110 &  x122 &  x137 &  x164 &  x170 &  x173 &  x185 &  x188 &  x254 &  x296 &  x326 &  x332 &  x347 &  x353 &  x392 &  x407 &  x410 &  x452 &  x500 &  x503 &  x527 &  x560 &  x572 &  x578 &  x605 &  x623 &  x638 &  x671 &  x707 &  x779 &  x791 &  x794 &  x805 &  x815 &  x851 &  x863 &  x866 &  x875 &  x911 &  x913 &  x917 &  x1037 &  x1055 &  x1100 &  x1103 &  x1112 &  x1121 &  x1127 & ~x396 & ~x561 & ~x723 & ~x1098;
assign c747 =  x134 &  x209 &  x277 &  x299 &  x347 &  x355 &  x725 &  x754 &  x821 &  x1091 & ~x819 & ~x864 & ~x978 & ~x1017 & ~x1056;
assign c749 =  x137 &  x393 &  x832 & ~x1056;
assign c751 = ~x815;
assign c753 =  x196 &  x277 & ~x129 & ~x247 & ~x936;
assign c755 =  x95 &  x98 &  x124 &  x128 &  x143 &  x209 &  x217 &  x452 &  x461 &  x515 &  x551 &  x563 &  x566 &  x593 &  x685 &  x686 &  x692 &  x752 &  x788 &  x812 &  x815 &  x827 &  x893 &  x920 &  x950 &  x980 &  x1040 &  x1073 &  x1079 &  x1121 & ~x282 & ~x867 & ~x1098;
assign c757 =  x276 &  x394 & ~x247;
assign c759 =  x11 &  x29 &  x41 &  x50 &  x53 &  x62 &  x71 &  x98 &  x101 &  x116 &  x119 &  x137 &  x161 &  x167 &  x182 &  x218 &  x221 &  x233 &  x260 &  x272 &  x280 &  x299 &  x326 &  x335 &  x353 &  x362 &  x383 &  x392 &  x395 &  x407 &  x419 &  x431 &  x437 &  x440 &  x461 &  x470 &  x488 &  x509 &  x530 &  x533 &  x542 &  x551 &  x569 &  x584 &  x590 &  x593 &  x599 &  x602 &  x617 &  x625 &  x626 &  x650 &  x680 &  x686 &  x719 &  x749 &  x785 &  x797 &  x800 &  x833 &  x839 &  x848 &  x854 &  x866 &  x881 &  x890 &  x917 &  x920 &  x947 &  x965 &  x992 &  x1004 &  x1025 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1064 &  x1088 &  x1103 & ~x516 & ~x555 & ~x594 & ~x669 & ~x687 & ~x786;
assign c763 =  x978 &  x1056 & ~x973;
assign c765 =  x331 &  x617 &  x662 &  x956 &  x979 & ~x390 & ~x432 & ~x711;
assign c767 =  x167 &  x377 &  x497 &  x611 &  x656 &  x667 &  x692 &  x743 &  x1076 &  x1094 & ~x558 & ~x636 & ~x864 & ~x1056;
assign c769 =  x273 &  x394 & ~x207 & ~x507;
assign c771 =  x17 &  x134 &  x179 &  x200 &  x203 &  x290 &  x299 &  x335 &  x338 &  x446 &  x467 &  x472 &  x490 &  x593 &  x596 &  x620 &  x800 &  x821 &  x845 &  x851 &  x905 &  x929 &  x941 &  x974 &  x994 &  x1043 &  x1103 &  x1130 & ~x483;
assign c773 =  x308 &  x355 &  x401 &  x524 &  x548 &  x680 &  x692 &  x869 &  x956 &  x1025 &  x1073 & ~x600 & ~x729 & ~x897 & ~x936 & ~x1095;
assign c775 =  x322 &  x586 &  x589 &  x745 &  x916 & ~x654;
assign c777 =  x72 &  x262 &  x436 &  x585 &  x868 & ~x675;
assign c779 =  x115 &  x176 &  x179 &  x218 &  x263 &  x464 &  x470 &  x479 &  x524 &  x592 &  x599 &  x731 &  x743 &  x823 &  x899 &  x995 &  x1019 &  x1100 & ~x1125;
assign c781 =  x985 & ~x102 & ~x328 & ~x585;
assign c783 =  x2 &  x14 &  x47 &  x50 &  x56 &  x59 &  x83 &  x89 &  x101 &  x104 &  x110 &  x116 &  x119 &  x122 &  x125 &  x131 &  x146 &  x152 &  x158 &  x170 &  x173 &  x188 &  x215 &  x218 &  x221 &  x233 &  x253 &  x278 &  x287 &  x292 &  x305 &  x308 &  x320 &  x332 &  x335 &  x371 &  x377 &  x380 &  x398 &  x407 &  x410 &  x416 &  x431 &  x434 &  x443 &  x452 &  x461 &  x476 &  x479 &  x482 &  x491 &  x497 &  x506 &  x524 &  x533 &  x536 &  x539 &  x545 &  x548 &  x581 &  x587 &  x596 &  x608 &  x611 &  x617 &  x623 &  x638 &  x641 &  x656 &  x677 &  x692 &  x698 &  x737 &  x743 &  x749 &  x773 &  x779 &  x788 &  x791 &  x794 &  x797 &  x812 &  x818 &  x851 &  x854 &  x869 &  x884 &  x887 &  x890 &  x899 &  x917 &  x935 &  x938 &  x944 &  x956 &  x971 &  x976 &  x983 &  x1001 &  x1025 &  x1034 &  x1040 &  x1046 &  x1049 &  x1064 &  x1070 &  x1073 &  x1076 &  x1088 &  x1106 &  x1118 &  x1127 &  x1130 & ~x282 & ~x594 & ~x672 & ~x747 & ~x786;
assign c785 =  x17 &  x23 &  x44 &  x56 &  x65 &  x92 &  x101 &  x104 &  x164 &  x167 &  x170 &  x176 &  x179 &  x188 &  x194 &  x197 &  x208 &  x209 &  x212 &  x221 &  x230 &  x254 &  x260 &  x275 &  x286 &  x296 &  x308 &  x320 &  x356 &  x359 &  x365 &  x380 &  x395 &  x401 &  x410 &  x416 &  x443 &  x452 &  x470 &  x482 &  x488 &  x503 &  x530 &  x533 &  x551 &  x554 &  x557 &  x575 &  x584 &  x602 &  x611 &  x632 &  x650 &  x659 &  x662 &  x677 &  x686 &  x698 &  x701 &  x707 &  x731 &  x737 &  x752 &  x764 &  x770 &  x773 &  x776 &  x779 &  x781 &  x794 &  x803 &  x818 &  x820 &  x821 &  x827 &  x839 &  x901 &  x917 &  x932 &  x938 &  x941 &  x947 &  x950 &  x971 &  x977 &  x980 &  x983 &  x989 &  x995 &  x1001 &  x1007 &  x1034 &  x1040 &  x1057 &  x1070 &  x1096 &  x1121 &  x1127 & ~x198 & ~x276 & ~x354 & ~x471;
assign c787 =  x34 &  x119 &  x140 &  x262 &  x338 &  x389 &  x412 &  x452 &  x475 &  x551 &  x635 &  x644 &  x746 &  x781 &  x923 &  x1010 &  x1054 &  x1102 & ~x276 & ~x714 & ~x825 & ~x903;
assign c789 =  x354 &  x1027 & ~x1095;
assign c791 =  x433 &  x490 & ~x484;
assign c793 =  x241 &  x280 &  x319 &  x433 & ~x441 & ~x498 & ~x705;
assign c795 =  x610 &  x883 & ~x562;
assign c797 =  x445 &  x470 &  x710 &  x862 &  x938 &  x940 &  x1057 & ~x195 & ~x315 & ~x690;
assign c799 =  x217 &  x334 &  x380 &  x698 & ~x438 & ~x444 & ~x1059;
assign c7101 =  x53 &  x131 &  x161 &  x248 &  x251 &  x383 &  x430 &  x469 &  x470 &  x502 &  x581 &  x584 &  x626 &  x647 &  x683 &  x701 &  x743 &  x827 &  x907 &  x932 &  x971 &  x1001 &  x1052 &  x1127 &  x1130 & ~x3 & ~x129 & ~x324 & ~x708 & ~x825 & ~x1059 & ~x1098;
assign c7103 =  x14 &  x26 &  x50 &  x53 &  x62 &  x65 &  x74 &  x77 &  x86 &  x95 &  x98 &  x101 &  x104 &  x119 &  x128 &  x137 &  x143 &  x146 &  x170 &  x173 &  x176 &  x179 &  x182 &  x188 &  x197 &  x206 &  x218 &  x221 &  x227 &  x248 &  x254 &  x281 &  x287 &  x290 &  x308 &  x311 &  x319 &  x332 &  x335 &  x338 &  x353 &  x356 &  x365 &  x377 &  x380 &  x389 &  x392 &  x394 &  x398 &  x410 &  x416 &  x428 &  x458 &  x461 &  x473 &  x479 &  x509 &  x515 &  x533 &  x539 &  x542 &  x548 &  x551 &  x554 &  x557 &  x566 &  x587 &  x602 &  x605 &  x623 &  x629 &  x632 &  x641 &  x647 &  x653 &  x674 &  x680 &  x683 &  x686 &  x689 &  x692 &  x704 &  x710 &  x713 &  x719 &  x740 &  x752 &  x755 &  x758 &  x761 &  x773 &  x794 &  x803 &  x812 &  x818 &  x821 &  x827 &  x830 &  x838 &  x842 &  x845 &  x854 &  x857 &  x869 &  x875 &  x878 &  x881 &  x884 &  x893 &  x902 &  x905 &  x907 &  x911 &  x917 &  x923 &  x932 &  x935 &  x944 &  x950 &  x953 &  x956 &  x959 &  x962 &  x965 &  x971 &  x986 &  x995 &  x1007 &  x1019 &  x1031 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1058 &  x1064 &  x1073 &  x1076 &  x1079 &  x1091 &  x1094 &  x1100 &  x1103 &  x1121 &  x1124 & ~x261;
assign c7105 =  x488 &  x494 &  x581 &  x625 &  x706 &  x707 &  x851 &  x901 &  x946 &  x974 &  x977 &  x1010 & ~x120 & ~x237;
assign c7107 =  x276 &  x433 & ~x703 & ~x1092;
assign c7109 =  x628 &  x667 & ~x480 & ~x963 & ~x1059 & ~x1080;
assign c7111 =  x358 &  x401 &  x925 &  x1053 &  x1102 & ~x198 & ~x825;
assign c7113 =  x14 &  x32 &  x77 &  x233 &  x302 &  x491 &  x503 &  x572 &  x638 &  x668 &  x790 &  x832 &  x988 &  x1066 & ~x693;
assign c7115 =  x44 &  x110 &  x155 &  x176 &  x257 &  x298 &  x319 &  x569 &  x917 &  x956 &  x986 &  x1040 &  x1082 &  x1112 & ~x198 & ~x519 & ~x558 & ~x708 & ~x726 & ~x1059;
assign c7117 =  x193 &  x823 &  x861 &  x1057 & ~x603;
assign c7119 =  x588 &  x744;
assign c7121 =  x312 & ~x247 & ~x289;
assign c7123 =  x28 &  x77 &  x133 &  x347 &  x389 &  x614 &  x725 &  x737 &  x745 &  x776 &  x784 &  x791 &  x1018 &  x1057 & ~x492;
assign c7125 =  x202 &  x586 & ~x207 & ~x498 & ~x1098;
assign c7127 =  x784 &  x1018 & ~x273 & ~x792 & ~x810;
assign c7129 =  x355 &  x532 &  x973 & ~x186 & ~x483 & ~x900;
assign c7131 =  x396 &  x433 &  x547;
assign c7133 =  x2 &  x5 &  x7 &  x8 &  x17 &  x20 &  x23 &  x26 &  x32 &  x35 &  x44 &  x47 &  x50 &  x53 &  x56 &  x59 &  x65 &  x68 &  x77 &  x83 &  x86 &  x92 &  x98 &  x101 &  x107 &  x122 &  x125 &  x134 &  x137 &  x143 &  x146 &  x152 &  x155 &  x164 &  x167 &  x176 &  x179 &  x185 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x215 &  x218 &  x227 &  x230 &  x236 &  x239 &  x251 &  x257 &  x263 &  x269 &  x275 &  x278 &  x281 &  x287 &  x299 &  x302 &  x314 &  x317 &  x323 &  x326 &  x329 &  x335 &  x338 &  x341 &  x344 &  x347 &  x350 &  x356 &  x359 &  x362 &  x365 &  x368 &  x371 &  x374 &  x377 &  x383 &  x386 &  x392 &  x398 &  x401 &  x404 &  x407 &  x410 &  x413 &  x416 &  x425 &  x428 &  x431 &  x434 &  x437 &  x443 &  x449 &  x452 &  x455 &  x458 &  x464 &  x470 &  x473 &  x476 &  x479 &  x485 &  x488 &  x491 &  x494 &  x497 &  x500 &  x503 &  x506 &  x509 &  x515 &  x518 &  x521 &  x524 &  x527 &  x533 &  x536 &  x539 &  x542 &  x548 &  x551 &  x554 &  x557 &  x560 &  x563 &  x566 &  x572 &  x575 &  x578 &  x584 &  x587 &  x590 &  x593 &  x596 &  x599 &  x602 &  x605 &  x608 &  x611 &  x614 &  x620 &  x626 &  x629 &  x635 &  x644 &  x647 &  x650 &  x656 &  x659 &  x662 &  x665 &  x671 &  x674 &  x680 &  x683 &  x689 &  x692 &  x695 &  x701 &  x704 &  x707 &  x710 &  x713 &  x716 &  x719 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x746 &  x752 &  x770 &  x773 &  x776 &  x779 &  x782 &  x785 &  x788 &  x791 &  x794 &  x797 &  x800 &  x803 &  x806 &  x812 &  x815 &  x818 &  x821 &  x830 &  x833 &  x836 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x860 &  x866 &  x869 &  x872 &  x887 &  x893 &  x896 &  x902 &  x908 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x941 &  x944 &  x950 &  x959 &  x965 &  x968 &  x971 &  x974 &  x977 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1004 &  x1013 &  x1019 &  x1031 &  x1034 &  x1037 &  x1040 &  x1043 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1118 &  x1124 & ~x129 & ~x672 & ~x747 & ~x864;
assign c7135 =  x34 &  x319 &  x758 &  x821 &  x1024 & ~x633 & ~x669 & ~x876 & ~x1059;
assign c7137 =  x217 &  x784 &  x979 & ~x834;
assign c7139 =  x769 &  x985 & ~x159 & ~x402 & ~x708 & ~x1071;
assign c7141 =  x433 &  x955 &  x973 &  x983 & ~x363 & ~x630 & ~x900;
assign c7143 =  x32 &  x194 &  x233 &  x347 &  x419 &  x791 &  x890 &  x911 &  x1022 &  x1037 &  x1085 & ~x246 & ~x265 & ~x396 & ~x747;
assign c7145 =  x154 &  x232 &  x685 &  x779 &  x784 & ~x828;
assign c7147 =  x250 &  x745 &  x1024 & ~x492 & ~x531;
assign c7149 =  x8 &  x14 &  x20 &  x26 &  x29 &  x32 &  x38 &  x41 &  x44 &  x50 &  x53 &  x59 &  x116 &  x119 &  x122 &  x139 &  x146 &  x164 &  x178 &  x224 &  x239 &  x260 &  x262 &  x281 &  x295 &  x334 &  x347 &  x353 &  x359 &  x386 &  x389 &  x401 &  x443 &  x452 &  x464 &  x470 &  x476 &  x482 &  x491 &  x494 &  x500 &  x503 &  x506 &  x512 &  x557 &  x575 &  x578 &  x599 &  x626 &  x653 &  x671 &  x692 &  x701 &  x728 &  x794 &  x803 &  x821 &  x857 &  x862 &  x863 &  x911 &  x914 &  x965 &  x974 &  x986 &  x989 &  x1043 &  x1057 &  x1073 &  x1100 &  x1103 &  x1109 &  x1114 & ~x471;
assign c7151 =  x699 & ~x834 & ~x1086;
assign c7153 =  x823 & ~x121 & ~x1107;
assign c7155 =  x217 &  x745 & ~x81 & ~x453 & ~x1059;
assign c7157 =  x564 &  x732 &  x888;
assign c7159 = ~x278;
assign c7161 =  x550 &  x628 &  x844 & ~x654 & ~x717;
assign c7163 =  x23 &  x56 &  x71 &  x86 &  x98 &  x155 &  x157 &  x178 &  x188 &  x230 &  x235 &  x242 &  x347 &  x377 &  x380 &  x434 &  x455 &  x461 &  x476 &  x482 &  x494 &  x515 &  x521 &  x593 &  x596 &  x646 &  x683 &  x685 &  x730 &  x755 &  x761 &  x806 &  x829 &  x839 &  x848 &  x863 &  x908 &  x911 &  x935 &  x965 &  x986 &  x989 &  x1013 &  x1025 &  x1121 & ~x285 & ~x324 & ~x900 & ~x1017 & ~x1098;
assign c7165 =  x34 &  x397 &  x454 &  x475 &  x719 &  x938 & ~x168 & ~x636 & ~x876 & ~x1059;
assign c7167 =  x8 &  x11 &  x23 &  x29 &  x35 &  x38 &  x47 &  x59 &  x71 &  x74 &  x89 &  x92 &  x95 &  x107 &  x110 &  x116 &  x131 &  x158 &  x161 &  x176 &  x179 &  x194 &  x196 &  x209 &  x212 &  x215 &  x248 &  x254 &  x274 &  x281 &  x299 &  x311 &  x317 &  x347 &  x368 &  x371 &  x377 &  x395 &  x398 &  x413 &  x419 &  x428 &  x434 &  x446 &  x464 &  x491 &  x509 &  x512 &  x521 &  x524 &  x527 &  x530 &  x533 &  x539 &  x548 &  x569 &  x593 &  x599 &  x617 &  x623 &  x632 &  x656 &  x671 &  x701 &  x710 &  x722 &  x737 &  x749 &  x767 &  x773 &  x776 &  x806 &  x832 &  x842 &  x845 &  x866 &  x869 &  x871 &  x872 &  x875 &  x887 &  x902 &  x908 &  x935 &  x941 &  x947 &  x956 &  x974 &  x977 &  x983 &  x992 &  x995 &  x1016 &  x1022 &  x1034 &  x1040 &  x1046 &  x1061 &  x1067 &  x1073 &  x1079 &  x1085 &  x1091 &  x1103 &  x1112 &  x1121 &  x1127 & ~x129 & ~x435 & ~x666 & ~x975;
assign c7169 =  x115 &  x822 &  x940 &  x1057;
assign c7171 =  x29 &  x277 &  x556 &  x559 &  x637 &  x878 &  x1001 & ~x624 & ~x664 & ~x897;
assign c7173 =  x486 &  x838 &  x844 &  x850 &  x1042;
assign c7175 =  x40 &  x269 &  x460 &  x782 &  x845 &  x1034 &  x1081 &  x1092 &  x1102 &  x1112 & ~x903 & ~x1083 & ~x1116;
assign c7177 =  x85 &  x98 &  x104 &  x116 &  x122 &  x124 &  x131 &  x163 &  x185 &  x299 &  x319 &  x326 &  x341 &  x599 &  x686 &  x707 &  x836 &  x881 &  x899 &  x901 &  x905 &  x947 &  x953 &  x974 &  x1004 &  x1021 &  x1025 &  x1096 & ~x471;
assign c7179 =  x73 &  x106 &  x745 &  x784 & ~x24 & ~x1099;
assign c7181 =  x351 & ~x51 & ~x324 & ~x325 & ~x747;
assign c7183 =  x478 &  x940 & ~x234 & ~x1047;
assign c7185 =  x277 &  x532 &  x883 & ~x129 & ~x247;
assign c7187 =  x76 &  x939 &  x978 & ~x351 & ~x867;
assign c7189 =  x62 &  x143 &  x245 &  x266 &  x359 &  x395 &  x419 &  x446 &  x470 &  x494 &  x502 &  x503 &  x533 &  x635 &  x659 &  x704 &  x836 &  x938 &  x959 &  x965 &  x977 &  x1115 & ~x48 & ~x708 & ~x840 & ~x1035;
assign c7191 =  x415 &  x799 &  x883 & ~x742;
assign c7193 =  x5 &  x11 &  x14 &  x32 &  x41 &  x44 &  x47 &  x50 &  x56 &  x62 &  x71 &  x83 &  x92 &  x107 &  x113 &  x116 &  x119 &  x122 &  x125 &  x146 &  x152 &  x161 &  x164 &  x167 &  x182 &  x185 &  x200 &  x209 &  x251 &  x254 &  x260 &  x266 &  x272 &  x290 &  x293 &  x296 &  x299 &  x305 &  x311 &  x326 &  x332 &  x347 &  x371 &  x374 &  x401 &  x404 &  x407 &  x410 &  x419 &  x425 &  x431 &  x434 &  x437 &  x440 &  x443 &  x446 &  x472 &  x476 &  x479 &  x482 &  x485 &  x491 &  x494 &  x497 &  x500 &  x509 &  x511 &  x512 &  x515 &  x533 &  x536 &  x539 &  x548 &  x550 &  x551 &  x560 &  x569 &  x584 &  x587 &  x590 &  x599 &  x602 &  x608 &  x611 &  x617 &  x620 &  x632 &  x638 &  x641 &  x644 &  x656 &  x659 &  x668 &  x689 &  x695 &  x698 &  x701 &  x704 &  x713 &  x725 &  x731 &  x743 &  x746 &  x755 &  x764 &  x770 &  x824 &  x830 &  x833 &  x845 &  x848 &  x860 &  x863 &  x872 &  x884 &  x890 &  x908 &  x926 &  x932 &  x938 &  x944 &  x962 &  x968 &  x971 &  x980 &  x983 &  x989 &  x995 &  x998 &  x1004 &  x1013 &  x1016 &  x1019 &  x1025 &  x1031 &  x1037 &  x1049 &  x1052 &  x1055 &  x1061 &  x1073 &  x1082 &  x1088 &  x1097 &  x1106 &  x1115 &  x1130 & ~x3 & ~x360 & ~x900;
assign c7195 =  x315 &  x595 &  x793 &  x1066;
assign c7197 =  x44 &  x145 &  x170 &  x538 &  x617 &  x623 &  x685 &  x809 &  x824 &  x953 &  x1013 & ~x180 & ~x582 & ~x708 & ~x1098;
assign c7199 =  x445 &  x978 & ~x312 & ~x351 & ~x870;
assign c7201 =  x17 &  x146 &  x163 &  x202 &  x217 &  x224 &  x299 &  x344 &  x398 &  x401 &  x464 &  x841 &  x872 &  x1028 &  x1100 & ~x615 & ~x942 & ~x981;
assign c7203 =  x74 &  x634 &  x727 &  x799 &  x929 &  x1081 &  x1102;
assign c7205 = ~x803;
assign c7207 =  x198 & ~x286;
assign c7209 =  x783 &  x945;
assign c7211 =  x237 & ~x208;
assign c7213 =  x433 &  x544 &  x647 &  x692 &  x794 &  x854 &  x899 & ~x324 & ~x858 & ~x939;
assign c7215 =  x155 &  x511 &  x628 &  x667 &  x740 &  x784 & ~x855;
assign c7217 =  x177 &  x1024 & ~x246;
assign c7219 =  x11 &  x14 &  x17 &  x32 &  x38 &  x41 &  x53 &  x59 &  x62 &  x68 &  x71 &  x80 &  x83 &  x92 &  x95 &  x104 &  x110 &  x116 &  x119 &  x131 &  x140 &  x146 &  x155 &  x158 &  x164 &  x173 &  x176 &  x194 &  x200 &  x206 &  x209 &  x212 &  x215 &  x224 &  x227 &  x239 &  x245 &  x260 &  x266 &  x272 &  x275 &  x284 &  x296 &  x299 &  x302 &  x311 &  x320 &  x323 &  x338 &  x341 &  x344 &  x347 &  x353 &  x362 &  x365 &  x383 &  x389 &  x395 &  x404 &  x410 &  x413 &  x416 &  x419 &  x422 &  x428 &  x434 &  x458 &  x485 &  x491 &  x497 &  x506 &  x515 &  x518 &  x521 &  x524 &  x527 &  x533 &  x536 &  x542 &  x548 &  x554 &  x563 &  x572 &  x578 &  x584 &  x587 &  x593 &  x602 &  x608 &  x611 &  x620 &  x626 &  x632 &  x635 &  x638 &  x641 &  x656 &  x662 &  x665 &  x668 &  x677 &  x680 &  x689 &  x707 &  x710 &  x716 &  x719 &  x722 &  x725 &  x740 &  x743 &  x746 &  x752 &  x755 &  x770 &  x773 &  x779 &  x785 &  x791 &  x794 &  x800 &  x806 &  x812 &  x818 &  x821 &  x827 &  x833 &  x848 &  x854 &  x863 &  x866 &  x884 &  x887 &  x893 &  x908 &  x911 &  x920 &  x923 &  x932 &  x935 &  x938 &  x941 &  x947 &  x962 &  x965 &  x974 &  x977 &  x980 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1007 &  x1010 &  x1016 &  x1022 &  x1025 &  x1037 &  x1055 &  x1061 &  x1067 &  x1070 &  x1073 &  x1076 &  x1082 &  x1094 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1118 &  x1130 & ~x81 & ~x120 & ~x159 & ~x165 & ~x198 & ~x204 & ~x519 & ~x633 & ~x672 & ~x747;
assign c7221 =  x358 &  x445 &  x978 &  x1057;
assign c7223 =  x742 &  x784 &  x860 &  x884 &  x945 &  x988;
assign c7225 =  x23 &  x50 &  x80 &  x89 &  x98 &  x101 &  x107 &  x119 &  x122 &  x143 &  x146 &  x158 &  x197 &  x239 &  x242 &  x251 &  x263 &  x266 &  x275 &  x281 &  x314 &  x317 &  x323 &  x335 &  x359 &  x380 &  x407 &  x422 &  x428 &  x455 &  x467 &  x485 &  x491 &  x494 &  x512 &  x521 &  x527 &  x533 &  x539 &  x566 &  x569 &  x572 &  x590 &  x605 &  x611 &  x614 &  x617 &  x626 &  x629 &  x635 &  x641 &  x647 &  x665 &  x668 &  x683 &  x701 &  x722 &  x728 &  x734 &  x740 &  x779 &  x791 &  x794 &  x812 &  x820 &  x824 &  x833 &  x860 &  x896 &  x908 &  x914 &  x923 &  x926 &  x929 &  x940 &  x941 &  x971 &  x979 &  x986 &  x998 &  x1010 &  x1018 &  x1040 &  x1058 &  x1067 &  x1070 &  x1076 &  x1112 &  x1118 & ~x81 & ~x120 & ~x198 & ~x237 & ~x471 & ~x549 & ~x759;
assign c7227 =  x76 &  x391 &  x394 & ~x552;
assign c7229 =  x65 &  x128 &  x152 &  x155 &  x266 &  x287 &  x350 &  x394 &  x464 &  x488 &  x494 &  x503 &  x578 &  x617 &  x715 &  x755 &  x764 &  x800 &  x832 &  x838 &  x842 &  x895 &  x914 &  x944 &  x953 &  x1019 &  x1088 & ~x822 & ~x861 & ~x1056 & ~x1095;
assign c7231 =  x237 &  x478 &  x637 & ~x303;
assign c7233 =  x550 &  x949 & ~x963 & ~x1093;
assign c7235 =  x5 &  x26 &  x92 &  x170 &  x335 &  x374 &  x395 &  x422 &  x473 &  x584 &  x644 &  x797 &  x940 &  x968 &  x1018 & ~x120 & ~x198 & ~x354 & ~x390 & ~x792 & ~x870;
assign c7237 =  x85 &  x263 &  x379 &  x485 & ~x438 & ~x672 & ~x1044;
assign c7239 =  x901 &  x1057 &  x1101 & ~x120;
assign c7241 =  x667 & ~x78 & ~x516 & ~x780;
assign c7243 =  x469 &  x472 &  x701 &  x818 &  x884 & ~x441 & ~x531 & ~x669;
assign c7245 =  x40 &  x163 & ~x90 & ~x1098;
assign c7247 =  x592 &  x823 & ~x234 & ~x315 & ~x636;
assign c7249 =  x883 & ~x562;
assign c7251 =  x315 & ~x591 & ~x975 & ~x1095;
assign c7253 =  x1096 & ~x399 & ~x817 & ~x870 & ~x876;
assign c7255 =  x5 &  x17 &  x26 &  x38 &  x56 &  x68 &  x104 &  x116 &  x119 &  x122 &  x137 &  x167 &  x176 &  x182 &  x194 &  x200 &  x209 &  x230 &  x257 &  x272 &  x275 &  x284 &  x296 &  x308 &  x316 &  x355 &  x365 &  x374 &  x377 &  x386 &  x389 &  x395 &  x410 &  x416 &  x422 &  x425 &  x428 &  x449 &  x464 &  x470 &  x497 &  x527 &  x545 &  x557 &  x566 &  x569 &  x590 &  x617 &  x629 &  x638 &  x653 &  x656 &  x662 &  x665 &  x674 &  x677 &  x701 &  x715 &  x731 &  x740 &  x785 &  x818 &  x821 &  x827 &  x833 &  x839 &  x845 &  x848 &  x863 &  x869 &  x872 &  x881 &  x884 &  x893 &  x902 &  x914 &  x917 &  x920 &  x926 &  x938 &  x947 &  x962 &  x971 &  x974 &  x986 &  x1001 &  x1004 &  x1010 &  x1028 &  x1031 &  x1043 &  x1055 &  x1061 &  x1085 &  x1097 &  x1103 &  x1112 &  x1124 & ~x225 & ~x303 & ~x342 & ~x405 & ~x861 & ~x939 & ~x1014 & ~x1017 & ~x1053 & ~x1056;
assign c7257 =  x472 &  x560 &  x608 &  x1100 & ~x645 & ~x723 & ~x780 & ~x786 & ~x1095;
assign c7259 =  x664 & ~x162 & ~x195 & ~x312 & ~x441 & ~x675 & ~x864;
assign c7261 =  x472 & ~x325 & ~x858;
assign c7263 =  x178 &  x598 & ~x462 & ~x664;
assign c7265 =  x110 &  x200 &  x251 &  x469 &  x593 &  x596 &  x740 &  x868 &  x893 & ~x552 & ~x582 & ~x741 & ~x813;
assign c7267 =  x478 &  x901 &  x1024 & ~x87 & ~x726;
assign c7269 =  x164 &  x260 &  x296 &  x323 &  x472 &  x511 &  x751 &  x812 &  x986 &  x1004 &  x1066 &  x1106 & ~x303 & ~x741;
assign c7271 =  x22 &  x77 &  x104 &  x161 &  x190 &  x284 &  x320 &  x326 &  x356 &  x485 &  x503 &  x539 &  x737 &  x794 &  x905 &  x907 &  x989 &  x1091 & ~x597 & ~x708;
assign c7273 =  x978 & ~x273 & ~x390 & ~x870;
assign c7275 =  x664 &  x823 &  x980 &  x1091 & ~x354 & ~x636 & ~x693;
assign c7277 =  x2 &  x8 &  x62 &  x71 &  x113 &  x128 &  x143 &  x209 &  x218 &  x320 &  x323 &  x350 &  x355 &  x386 &  x413 &  x425 &  x433 &  x443 &  x476 &  x482 &  x512 &  x554 &  x557 &  x581 &  x584 &  x596 &  x608 &  x617 &  x680 &  x692 &  x701 &  x710 &  x713 &  x715 &  x764 &  x767 &  x773 &  x778 &  x788 &  x799 &  x821 &  x833 &  x839 &  x844 &  x850 &  x896 &  x908 &  x914 &  x950 &  x956 &  x962 &  x977 &  x989 &  x1034 &  x1052 &  x1085 &  x1100 &  x1121 &  x1124;
assign c7279 =  x73 &  x140 &  x256 &  x509 &  x632 &  x770 & ~x120 & ~x636 & ~x1104;
assign c7281 =  x589 &  x994 & ~x3;
assign c7283 =  x328 &  x784 &  x823 & ~x78 & ~x117 & ~x714 & ~x1035;
assign c7285 =  x430 &  x560 &  x563 &  x757 &  x884 & ~x51 & ~x90 & ~x399 & ~x474 & ~x513 & ~x552 & ~x558 & ~x675;
assign c7287 =  x667 &  x706 &  x940 & ~x3 & ~x198 & ~x318;
assign c7291 =  x42 &  x592 &  x718 & ~x52;
assign c7293 =  x358 &  x433 &  x949 & ~x303;
assign c7295 =  x76 &  x221 &  x280 &  x319 &  x338 &  x467 &  x683 &  x716 &  x746 &  x752 &  x779 &  x1010 &  x1127 & ~x516 & ~x903 & ~x1125;
assign c7297 =  x784 &  x940 & ~x118;
assign c7299 =  x134 &  x235 &  x272 &  x273 &  x521 &  x572 &  x611 &  x650 &  x743 &  x959 &  x1081 & ~x90 & ~x91 & ~x207 & ~x588;

endmodule