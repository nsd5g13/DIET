module tm( x0,x1,x2,x3,x4,x5,x6,x7,x8,x9,x10,x11,x12,x13,x14,x15,x16,x17,x18,x19,x20,x21,x22,x23,x24,x25,x26,x27,x28,x29,x30,x31,x32,x33,x34,x35,x36,x37,x38,x39,x40,x41,x42,x43,x44,x45,x46,x47,x48,x49,x50,x51,x52,x53,x54,x55,x56,x57,x58,x59,x60,x61,x62,x63,x64,x65,x66,x67,x68,x69,x70,x71,x72,x73,x74,x75,x76,x77,x78,x79,x80,x81,x82,x83,x84,x85,x86,x87,x88,x89,x90,x91,x92,x93,x94,x95,x96,x97,x98,x99,x100,x101,x102,x103,x104,x105,x106,x107,x108,x109,x110,x111,x112,x113,x114,x115,x116,x117,x118,x119,x120,x121,x122,x123,x124,x125,x126,x127,x128,x129,x130,x131,x132,x133,x134,x135,x136,x137,x138,x139,x140,x141,x142,x143,x144,x145,x146,x147,x148,x149,x150,x151,x152,x153,x154,x155,x156,x157,x158,x159,x160,x161,x162,x163,x164,x165,x166,x167,x168,x169,x170,x171,x172,x173,x174,x175,x176,x177,x178,x179,x180,x181,x182,x183,x184,x185,x186,x187,x188,x189,x190,x191,x192,x193,x194,x195,x196,x197,x198,x199,x200,x201,x202,x203,x204,x205,x206,x207,x208,x209,x210,x211,x212,x213,x214,x215,x216,x217,x218,x219,x220,x221,x222,x223,x224,x225,x226,x227,x228,x229,x230,x231,x232,x233,x234,x235,x236,x237,x238,x239,x240,x241,x242,x243,x244,x245,x246,x247,x248,x249,x250,x251,x252,x253,x254,x255,x256,x257,x258,x259,x260,x261,x262,x263,x264,x265,x266,x267,x268,x269,x270,x271,x272,x273,x274,x275,x276,x277,x278,x279,x280,x281,x282,x283,x284,x285,x286,x287,x288,x289,x290,x291,x292,x293,x294,x295,x296,x297,x298,x299,x300,x301,x302,x303,x304,x305,x306,x307,x308,x309,x310,x311,x312,x313,x314,x315,x316,x317,x318,x319,x320,x321,x322,x323,x324,x325,x326,x327,x328,x329,x330,x331,x332,x333,x334,x335,x336,x337,x338,x339,x340,x341,x342,x343,x344,x345,x346,x347,x348,x349,x350,x351,x352,x353,x354,x355,x356,x357,x358,x359,x360,x361,x362,x363,x364,x365,x366,x367,x368,x369,x370,x371,x372,x373,x374,x375,x376,x377,x378,x379,x380,x381,x382,x383,x384,x385,x386,x387,x388,x389,x390,x391,x392,x393,x394,x395,x396,x397,x398,x399,x400,x401,x402,x403,x404,x405,x406,x407,x408,x409,x410,x411,x412,x413,x414,x415,x416,x417,x418,x419,x420,x421,x422,x423,x424,x425,x426,x427,x428,x429,x430,x431,x432,x433,x434,x435,x436,x437,x438,x439,x440,x441,x442,x443,x444,x445,x446,x447,x448,x449,x450,x451,x452,x453,x454,x455,x456,x457,x458,x459,x460,x461,x462,x463,x464,x465,x466,x467,x468,x469,x470,x471,x472,x473,x474,x475,x476,x477,x478,x479,x480,x481,x482,x483,x484,x485,x486,x487,x488,x489,x490,x491,x492,x493,x494,x495,x496,x497,x498,x499,x500,x501,x502,x503,x504,x505,x506,x507,x508,x509,x510,x511,x512,x513,x514,x515,x516,x517,x518,x519,x520,x521,x522,x523,x524,x525,x526,x527,x528,x529,x530,x531,x532,x533,x534,x535,x536,x537,x538,x539,x540,x541,x542,x543,x544,x545,x546,x547,x548,x549,x550,x551,x552,x553,x554,x555,x556,x557,x558,x559,x560,x561,x562,x563,x564,x565,x566,x567,x568,x569,x570,x571,x572,x573,x574,x575,x576,x577,x578,x579,x580,x581,x582,x583,x584,x585,x586,x587,x588,x589,x590,x591,x592,x593,x594,x595,x596,x597,x598,x599,x600,x601,x602,x603,x604,x605,x606,x607,x608,x609,x610,x611,x612,x613,x614,x615,x616,x617,x618,x619,x620,x621,x622,x623,x624,x625,x626,x627,x628,x629,x630,x631,x632,x633,x634,x635,x636,x637,x638,x639,x640,x641,x642,x643,x644,x645,x646,x647,x648,x649,x650,x651,x652,x653,x654,x655,x656,x657,x658,x659,x660,x661,x662,x663,x664,x665,x666,x667,x668,x669,x670,x671,x672,x673,x674,x675,x676,x677,x678,x679,x680,x681,x682,x683,x684,x685,x686,x687,x688,x689,x690,x691,x692,x693,x694,x695,x696,x697,x698,x699,x700,x701,x702,x703,x704,x705,x706,x707,x708,x709,x710,x711,x712,x713,x714,x715,x716,x717,x718,x719,x720,x721,x722,x723,x724,x725,x726,x727,x728,x729,x730,x731,x732,x733,x734,x735,x736,x737,x738,x739,x740,x741,x742,x743,x744,x745,x746,x747,x748,x749,x750,x751,x752,x753,x754,x755,x756,x757,x758,x759,x760,x761,x762,x763,x764,x765,x766,x767,x768,x769,x770,x771,x772,x773,x774,x775,x776,x777,x778,x779,x780,x781,x782,x783,x784,x785,x786,x787,x788,x789,x790,x791,x792,x793,x794,x795,x796,x797,x798,x799,x800,x801,x802,x803,x804,x805,x806,x807,x808,x809,x810,x811,x812,x813,x814,x815,x816,x817,x818,x819,x820,x821,x822,x823,x824,x825,x826,x827,x828,x829,x830,x831,x832,x833,x834,x835,x836,x837,x838,x839,x840,x841,x842,x843,x844,x845,x846,x847,x848,x849,x850,x851,x852,x853,x854,x855,x856,x857,x858,x859,x860,x861,x862,x863,x864,x865,x866,x867,x868,x869,x870,x871,x872,x873,x874,x875,x876,x877,x878,x879,x880,x881,x882,x883,x884,x885,x886,x887,x888,x889,x890,x891,x892,x893,x894,x895,x896,x897,x898,x899,x900,x901,x902,x903,x904,x905,x906,x907,x908,x909,x910,x911,x912,x913,x914,x915,x916,x917,x918,x919,x920,x921,x922,x923,x924,x925,x926,x927,x928,x929,x930,x931,x932,x933,x934,x935,x936,x937,x938,x939,x940,x941,x942,x943,x944,x945,x946,x947,x948,x949,x950,x951,x952,x953,x954,x955,x956,x957,x958,x959,x960,x961,x962,x963,x964,x965,x966,x967,x968,x969,x970,x971,x972,x973,x974,x975,x976,x977,x978,x979,x980,x981,x982,x983,x984,x985,x986,x987,x988,x989,x990,x991,x992,x993,x994,x995,x996,x997,x998,x999,x1000,x1001,x1002,x1003,x1004,x1005,x1006,x1007,x1008,x1009,x1010,x1011,x1012,x1013,x1014,x1015,x1016,x1017,x1018,x1019,x1020,x1021,x1022,x1023,x1024,x1025,x1026,x1027,x1028,x1029,x1030,x1031,x1032,x1033,x1034,x1035,x1036,x1037,x1038,x1039,x1040,x1041,x1042,x1043,x1044,x1045,x1046,x1047,x1048,x1049,x1050,x1051,x1052,x1053,x1054,x1055,x1056,x1057,x1058,x1059,x1060,x1061,x1062,x1063,x1064,x1065,x1066,x1067,x1068,x1069,x1070,x1071,x1072,x1073,x1074,x1075,x1076,x1077,x1078,x1079,x1080,x1081,x1082,x1083,x1084,x1085,x1086,x1087,x1088,x1089,x1090,x1091,x1092,x1093,x1094,x1095,x1096,x1097,x1098,x1099,x1100,x1101,x1102,x1103,x1104,x1105,x1106,x1107,x1108,x1109,x1110,x1111,x1112,x1113,x1114,x1115,x1116,x1117,x1118,x1119,x1120,x1121,x1122,x1123,x1124,x1125,x1126,x1127,x1128,x1129,x1130,c0219,c1253,c5138,c4199,c10,c0130,c6133,c7113,c3121,c6236,c0182,c4187,c650,c41,c7299,c5289,c0298,c5161,c698,c3284,c454,c4250,c737,c58,c332,c134,c4181,c468,c1279,c032,c7220,c6164,c0185,c348,c0217,c2171,c5288,c21,c4198,c145,c378,c358,c399,c55,c116,c4221,c7159,c270,c7133,c1165,c3279,c578,c4269,c4151,c6285,c3189,c492,c2142,c1299,c7161,c686,c7285,c247,c7176,c0214,c7125,c3162,c4170,c2274,c1297,c7116,c3133,c721,c15,c4243,c5235,c0104,c722,c370,c572,c5222,c532,c1150,c5199,c038,c335,c513,c123,c5230,c651,c6124,c147,c050,c6225,c3228,c3215,c4291,c6202,c2293,c210,c1184,c276,c4185,c2165,c3273,c214,c3122,c6186,c0200,c2117,c6138,c7251,c2280,c0238,c1124,c7289,c039,c057,c2109,c5112,c3288,c4176,c3207,c6221,c23,c798,c7157,c2249,c33,c3219,c556,c7249,c5187,c5272,c4147,c7164,c5197,c13,c0294,c7150,c125,c3244,c021,c727,c0276,c2262,c158,c1132,c2284,c1209,c4165,c6166,c3221,c498,c0113,c146,c460,c5225,c2224,c2244,c1206,c6156,c6281,c740,c1180,c597,c2217,c222,c1200,c6110,c0146,c4188,c739,c1264,c1123,c345,c539,c4222,c3270,c632,c7278,c196,c6289,c5170,c6226,c3124,c1273,c777,c6299,c220,c5265,c7221,c218,c0132,c5105,c0189,c6102,c7257,c3182,c494,c379,c7224,c6224,c052,c0179,c133,c7228,c769,c475,c575,c5132,c212,c096,c176,c664,c0291,c1213,c6198,c687,c0259,c1160,c3136,c1278,c618,c1274,c3267,c4200,c4173,c2164,c248,c7281,c234,c2172,c794,c411,c699,c5278,c3138,c2273,c779,c09,c3141,c1283,c476,c483,c1269,c7219,c7296,c1291,c2237,c173,c4201,c464,c245,c4215,c4264,c4274,c2139,c4161,c7202,c751,c0117,c7162,c3106,c184,c5143,c510,c3283,c59,c3179,c1227,c3140,c6119,c4276,c3195,c6290,c3161,c4137,c4116,c6120,c6151,c7141,c180,c1252,c5208,c0203,c782,c012,c2182,c2207,c19,c393,c536,c7290,c251,c3236,c0241,c5211,c4225,c0224,c770,c0153,c5109,c6175,c1192,c5104,c1151,c3127,c199,c0122,c4156,c6271,c768,c431,c2166,c7256,c5145,c0293,c3298,c7172,c2196,c14,c5209,c7232,c7269,c0116,c111,c5251,c718,c0147,c6167,c322,c5231,c4183,c3278,c6170,c74,c4229,c1282,c5136,c1186,c2153,c619,c6297,c5174,c3252,c1163,c450,c3134,c5244,c4235,c5139,c6114,c6192,c1289,c5134,c0149,c7143,c37,c0204,c6172,c5146,c7112,c17,c0143,c070,c663,c3282,c0159,c3276,c479,c5121,c2180,c221,c7124,c7265,c274,c1233,c645,c642,c1140,c5293,c261,c5290,c238,c7233,c4263,c3254,c48,c3253,c7155,c2113,c452,c489,c581,c331,c3105,c294,c4267,c5178,c7167,c5218,c5204,c0234,c3172,c242,c5198,c516,c535,c4298,c680,c2185,c372,c377,c0161,c0262,c669,c4106,c0281,c361,c3251,c0295,c1219,c4233,c398,c5295,c0180,c0134,c6275,c2108,c5229,c6242,c2211,c2299,c416,c570,c7139,c2140,c5297,c3110,c3292,c47,c195,c4211,c71,c5245,c098,c423,c2122,c693,c0198,c7110,c4287,c4252,c235,c7207,c6288,c066,c433,c1183,c4209,c1137,c758,c254,c4132,c4139,c5129,c0272,c0243,c4281,c2227,c1194,c6274,c0120,c5264,c3203,c1272,c6130,c4133,c5206,c76,c692,c088,c3148,c7166,c353,c3143,c1136,c00,c3116,c3152,c7208,c040,c112,c3209,c6195,c22,c2186,c3234,c4149,c3243,c5276,c3197,c312,c323,c589,c5151,c7126,c1158,c0154,c2214,c477,c3232,c463,c5113,c5281,c3206,c0229,c7200,c4193,c4128,c6181,c5268,c2110,c387,c1131,c3131,c140,c042,c065,c480,c3247,c491,c7226,c121,c4142,c7185,c7227,c5182,c1107,c5190,c4114,c4195,c0183,c048,c075,c0158,c314,c627,c7122,c4240,c493,c3125,c6251,c641,c6270,c229,c4277,c397,c0136,c7171,c243,c1142,c1118,c4294,c5115,c6207,c6272,c559,c32,c3132,c1152,c657,c689,c6105,c6174,c1189,c3220,c2193,c316,c2124,c149,c1268,c3275,c2145,c634,c3107,c067,c2132,c453,c177,c1281,c5216,c7198,c533,c7206,c1134,c0196,c519,c045,c6171,c2102,c120,c5262,c428,c5186,c1292,c2163,c4120,c5176,c1256,c557,c0226,c778,c0218,c3216,c7252,c0285,c3184,c4270,c2136,c2178,c172,c78,c339,c2160,c246,c5116,c156,c0274,c7115,c435,c036,c7111,c0115,c2295,c781,c2255,c4228,c3103,c4191,c3272,c4121,c329,c5131,c451,c613,c3249,c0275,c797,c750,c2159,c4248,c5158,c390,c0249,c3150,c4282,c2148,c164,c6142,c053,c1277,c290,c5202,c371,c5128,c161,c6122,c2288,c5255,c671,c5155,c1280,c6250,c1231,c2278,c2257,c4205,c5201,c61,c6239,c4148,c3169,c6222,c4157,c4126,c759,c2246,c2215,c6121,c6169,c1254,c3277,c2183,c1104,c010,c4158,c4101,c5296,c3144,c138,c673,c3155,c6134,c3257,c4146,c0118,c5210,c1246,c26,c1122,c1290,c4164,c5181,c1110,c4179,c130,c0223,c414,c612,c670,c0192,c0145,c4135,c2233,c5154,c7214,c7240,c5184,c320,c328,c3214,c1237,c7277,c497,c1135,c631,c041,c730,c4265,c4254,c2285,c2112,c394,c082,c5253,c6205,c34,c4175,c3237,c644,c1211,c3293,c0142,c6232,c2268,c044,c6152,c090,c5233,c3229,c0282,c469,c6162,c7298,c7268,c2167,c637,c776,c3218,c594,c1262,c3146,c2222,c3111,c2188,c5141,c352,c7271,c4143,c656,c6103,c6154,c616,c3199,c6223,c3290,c061,c117,c7130,c461,c4238,c0232,c4256,c6267,c6111,c1170,c175,c1263,c6257,c324,c337,c6140,c262,c2208,c167,c0267,c2168,c343,c7294,c2232,c118,c646,c6287,c756,c719,c7118,c771,c0206,c019,c183,c565,c0252,c255,c2204,c1169,c6282,c062,c1275,c2298,c4289,c258,c0209,c30,c580,c1109,c2128,c554,c2118,c2245,c3296,c0127,c3289,c7107,c5196,c5246,c2212,c0207,c2270,c056,c4154,c659,c7182,c2236,c035,c0254,c2252,c4266,c0169,c5126,c5277,c313,c1224,c5111,c0106,c1127,c295,c4241,c185,c1156,c1255,c0257,c5147,c667,c160,c4226,c647,c577,c064,c598,c6125,c2281,c7146,c0155,c696,c60,c544,c5167,c579,c1121,c5150,c68,c7108,c0255,c521,c5207,c793,c4192,c2158,c364,c374,c789,c6254,c3212,c3266,c2105,c5120,c2169,c472,c7201,c2195,c588,c3178,c260,c1129,c5217,c7135,c0278,c1216,c3118,c355,c439,c485,c1113,c351,c283,c0220,c2272,c51,c2170,c165,c655,c382,c749,c2239,c3168,c094,c287,c3213,c5127,c2251,c0227,c6245,c6199,c587,c7204,c2275,c7194,c6163,c6244,c3281,c1190,c043,c0190,c2152,c4118,c5172,c7272,c5180,c4214,c148,c6279,c0260,c457,c590,c53,c2101,c2265,c4283,c63,c5152,c783,c5169,c267,c2175,c0213,c092,c2242,c289,c31,c735,c5254,c3258,c1159,c2123,c660,c764,c2241,c4141,c6217,c444,c2216,c526,c7180,c745,c4236,c4131,c690,c6136,c427,c6296,c788,c169,c319,c3194,c5287,c599,c6208,c6231,c368,c4104,c6213,c380,c4258,c4224,c6190,c432,c5189,c6249,c1167,c253,c7273,c5292,c4145,c2297,c2261,c4136,c078,c1220,c0253,c7203,c3104,c2210,c349,c5135,c0231,c4177,c5164,c1146,c5142,c1222,c3204,c014,c1271,c731,c7129,c7173,c279,c189,c2125,c4174,c6259,c241,c06,c27,c1196,c5248,c3262,c3126,c4124,c49,c3294,c216,c1210,c760,c2225,c293,c7237,c0290,c2229,c540,c7222,c263,c266,c4134,c5194,c4100,c6144,c7276,c3246,c020,c350,c638,c6161,c5103,c3139,c4286,c058,c676,c4261,c197,c7218,c5234,c2279,c159,c142,c211,c1130,c5215,c3291,c6182,c3271,c675,c4260,c357,c7242,c3217,c2276,c4212,c0222,c0279,c6113,c333,c115,c186,c5291,c2129,c7261,c512,c3129,c013,c44,c1203,c5259,c7120,c213,c016,c514,c233,c0288,c5221,c4245,c317,c3286,c1173,c7184,c4140,c1266,c561,c055,c1119,c2127,c746,c1221,c086,c5108,c1197,c697,c6212,c1177,c7297,c079,c5157,c574,c7103,c7142,c5117,c3239,c2219,c4255,c1181,c4272,c3142,c6132,c6178,c4259,c0184,c192,c3259,c4249,c026,c534,c029,c487,c467,c0172,c528,c5160,c5193,c1101,c16,c518,c7128,c0150,c4117,c0195,c366,c4206,c5122,c0193,c6216,c1285,c0248,c7286,c7134,c280,c1125,c7245,c3156,c4246,c720,c1248,c7239,c1164,c520,c7193,c73,c3187,c3223,c269,c0233,c129,c470,c3108,c7179,c6139,c5185,c6280,c6183,c679,c0266,c6284,c141,c2291,c499,c7248,c7149,c135,c5271,c3287,c0139,c2116,c473,c592,c6234,c0121,c678,c7190,c1153,c227,c5279,c6135,c6292,c1260,c7205,c1114,c1174,c6241,c3240,c028,c1182,c4244,c7199,c419,c711,c424,c0162,c3114,c5227,c567,c2226,c347,c542,c69,c38,c0131,c591,c430,c547,c3163,c1191,c658,c02,c537,c3145,c373,c5294,c1241,c43,c356,c2200,c5166,c1187,c0191,c4189,c7105,c684,c7192,c0100,c6118,c0160,c063,c2107,c4232,c6180,c6230,c3166,c2181,c6235,c1247,c4115,c7160,c224,c6108,c2202,c5162,c555,c6187,c635,c1166,c3268,c1204,c0168,c5130,c1175,c6298,c2256,c0268,c456,c443,c2162,c465,c7152,c298,c155,c2157,c4251,c7136,c278,c5195,c0215,c6127,c3147,c7260,c0221,c6277,c346,c426,c6184,c775,c6252,c4297,c344,c236,c7241,c1240,c1257,c264,c07,c6240,c7186,c1111,c639,c018,c0171,c7209,c7195,c083,c6165,c1128,c273,c0107,c630,c5156,c2177,c4210,c2290,c363,c2254,c2104,c7145,c0299,c1139,c0271,c1235,c6238,c7254,c4122,c3160,c478,c7284,c330,c5205,c6233,c6168,c7183,c5102,c170,c3113,c0277,c1228,c568,c677,c2235,c2263,c0124,c437,c0283,c194,c3211,c5137,c04,c562,c0188,c7274,c369,c45,c2179,c5214,c2135,c0105,c097,c4182,c714,c0244,c0289,c383,c6262,c790,c755,c2203,c2267,c2120,c4295,c023,c3256,c228,c66,c7175,c442,c027,c113,c5191,c4163,c4180,c531,c011,c5213,c736,c7197,c1223,c672,c0126,c665,c05,c5260,c515,c1145,c1226,c5123,c386,c4194,c448,c0211,c5168,c7102,c7127,c179,c522,c034,c7267,c2134,c3153,c458,c3198,c2260,c5153,c136,c2282,c0135,c7283,c03,c1218,c18,c734,c4196,c1296,c35,c087,c6137,c3205,c488,c6157,c4253,c1176,c3175,c4296,c649,c1229,c1249,c4123,c5243,c743,c2199,c384,c3181,c546,c767,c742,c2191,c6256,c585,c2144,c418,c282,c694,c2190,c633,c5285,c1154,c1232,c1178,c2286,c4125,c7138,c7247,c6291,c766,c2121,c4105,c215,c126,c12,c5163,c1293,c01,c682,c037,c2155,c2151,c3123,c4150,c780,c2223,c774,c524,c420,c4219,c2130,c6265,c051,c2154,c5223,c0119,c5149,c6126,c1242,c3261,c6158,c3130,c0264,c681,c527,c0141,c0245,c5220,c413,c4280,c3185,c5179,c069,c6220,c7119,c272,c6286,c318,c5110,c297,c77,c6188,c447,c7295,c2194,c2289,c0181,c7106,c747,c1225,c4160,c4102,c754,c325,c410,c4271,c563,c310,c292,c5107,c391,c2221,c2228,c3264,c0280,c7181,c1198,c362,c7264,c017,c446,c5269,c7163,c7191,c7211,c360,c0235,c1276,c611,c1138,c1162,c2259,c388,c733,c122,c3248,c3280,c5133,c4208,c490,c661,c5118,c5250,c713,c2131,c3233,c1207,c2213,c6143,c025,c151,c582,c2106,c662,c412,c226,c3235,c2253,c5175,c4113,c6117,c2150,c0174,c288,c4217,c0216,c6293,c2198,c7187,c2292,c7258,c7244,c367,c4103,c5258,c342,c3226,c030,c5299,c786,c093,c3241,c2143,c054,c3157,c0173,c1270,c541,c392,c417,c4223,c4129,c1243,c1149,c796,c2137,c0284,c3188,c359,c4184,c163,c7238,c610,c0250,c75,c1251,c7189,c6148,c0197,c1141,c389,c787,c7140,c077,c1143,c471,c321,c4172,c586,c7196,c7156,c326,c4292,c6260,c2138,c7177,c7293,c571,c0242,c29,c3117,c614,c1298,c6100,c7234,c668,c7292,c7231,c334,c6123,c4293,c7131,c6261,c5114,c621,c2220,c6215,c573,c0102,c2243,c4239,c5274,c2111,c5256,c265,c2271,c3274,c748,c6264,c2205,c7223,c395,c08,c230,c2209,c652,c6219,c1265,c0144,c6258,c3255,c2147,c3208,c7235,c2296,c4213,c2192,c1295,c1157,c710,c1245,c6294,c728,c2234,c6278,c7154,c422,c762,c250,c5242,c0205,c3102,c150,c726,c4216,c2250,c0133,c0225,c0194,c5200,c685,c1168,c57,c4144,c7151,c4290,c6200,c4220,c67,c0128,c791,c3119,c271,c4186,c772,c5280,c4108,c7153,c550,c6263,c2231,c0265,c3186,c5203,c256,c2115,c132,c523,c595,c2247,c538,c1205,c268,c0186,c1188,c3183,c4110,c285,c1287,c3158,c6218,c191,c336,c1133,c3128,c6201,c7212,c1171,c7148,c28,c484,c763,c198,c1199,c2201,c4169,c6155,c085,c529,c5183,c6191,c144,c4153,c4207,c315,c049,c1115,c640,c552,c3196,c3202,c239,c4130,c1117,c4167,c46,c3170,c059,c429,c455,c2189,c421,c1103,c4197,c3180,c084,c72,c7280,c1155,c1147,c636,c3149,c6283,c0263,c0286,c1267,c7217,c0156,c744,c5282,c626,c081,c4285,c2126,c4166,c0163,c6147,c286,c7109,c275,c259,c593,c1244,c4111,c7243,c2266,c154,c0103,c629,c6116,c291,c4138,c4262,c0137,c143,c2218,c7137,c3238,c0261,c653,c3176,c0246,c1215,c6149,c0175,c723,c459,c6128,c0247,c3200,c7270,c0292,c396,c5263,c2173,c5257,c3174,c56,c139,c643,c5275,c7114,c666,c622,c225,c223,c0140,c244,c0151,c0129,c6150,c3224,c095,c162,c217,c257,c4152,c2114,c080,c0273,c64,c65,c2206,c617,c7123,c4204,c3231,c7169,c5247,c5232,c6115,c6246,c738,c4288,c1250,c157,c178,c3227,c6253,c3109,c732,c434,c0256,c1105,c376,c40,c1106,c0152,c4268,c6197,c6145,c2161,c1208,c5270,c7250,c1238,c7275,c3230,c1185,c2294,c2184,c1236,c4119,c249,c152,c5119,c2248,c340,c4218,c237,c482,c1148,c281,c076,c7216,c7262,c6196,c0258,c3151,c0166,c3177,c481,c511,c3173,c071,c7132,c7253,c015,c4178,c153,c4190,c39,c3101,c42,c7282,c716,c3159,c0114,c4227,c7213,c0287,c2187,c2197,c625,c1161,c252,c5286,c628,c70,c127,c3193,c089,c338,c495,c5237,c137,c4112,c2174,c5159,c6189,c7101,c7255,c2103,c438,c1172,c6101,c219,c1144,c717,c6276,c545,c6185,c0239,c5144,c0228,c7168,c099,c576,c7230,c1212,c6176,c232,c425,c2156,c0178,c171,c548,c0240,c5228,c240,c3137,c1116,c4275,c7165,c3171,c0201,c3201,c046,c20,c1179,c6210,c784,c327,c4155,c564,c3297,c0110,c566,c2283,c525,c6209,c5224,c7174,c0208,c1234,c7291,c0167,c2240,c6173,c068,c799,c7147,c354,c445,c168,c381,c4247,c5284,c4203,c6237,c757,c174,c25,c5100,c091,c741,c0297,c3295,c6160,c1230,c6273,c5298,c0125,c7100,c0199,c50,c073,c1202,c5148,c436,c0270,c1126,c440,c4278,c5226,c128,c773,c6269,c551,c3260,c6107,c7144,c6131,c0165,c284,c3222,c6268,c193,c7225,c553,c0202,c4234,c4231,c5236,c4273,c24,c7266,c3269,c0236,c474,c277,c5252,c623,c688,c299,c0138,c2238,c5266,c119,c7158,c5238,c031,c3263,c3245,c5283,c3100,c7121,c0157,c5171,c52,c0108,c4299,c569,c1214,c110,c795,c2141,c2119,c5261,c3299,c4242,c7288,c725,c6193,c0230,c0269,c2269,c2230,c7236,c3120,c0296,c3115,c0212,c1284,c5240,c6104,c311,c0177,c3135,c4162,c674,c441,c5192,c4284,c5273,c4237,c648,c615,c0170,c6203,c166,c2146,c724,c5239,c365,c4109,c3112,c683,c131,c624,c0187,c6141,c462,c5101,c596,c2133,c5249,c4230,c296,c6255,c0109,c584,c3242,c2277,c187,c729,c415,c7117,c3165,c341,c785,c62,c1102,c6153,c654,c715,c36,c4107,c072,c4171,c792,c0111,c1261,c2100,c1193,c5173,c1120,c691,c6227,c765,c6248,c060,c695,c3190,c4257,c188,c1286,c047,c560,c496,c6228,c7178,c3164,c7259,c1258,c6214,c0210,c4159,c5140,c6109,c6243,c517,c022,c3167,c6179,c6211,c4279,c5241,c6159,c182,c753,c449,c0251,c1195,c181,c7229,c486,c0123,c5125,c7263,c2287,c1201,c3210,c3192,c0112,c033,c3225,c5124,c79,c0148,c1259,c54,c6204,c7104,c0164,c0176,c3154,c6112,c231,c7246,c0237,c7188,c7287,c583,c190,c1288,c6106,c7279,c0101,c620,c6177,c466,c1217,c7215,c4127,c024,c6266,c530,c4168,c712,c6295,c7170,c3265,c6129,c6206,c761,c1112,c5219,c549,c1239,c6247,c114,c543,c3285,c1108,c3191,c558,c7210,c752,c6229,c074,c4202,c5106,c5177,c11,c375,c5188,c1294,c2258,c2176,c2264,c6146,c2149,c5165,c124,c1100,c5212,c5267,c6194,c3250,c385 );

input x0;
input x1;
input x2;
input x3;
input x4;
input x5;
input x6;
input x7;
input x8;
input x9;
input x10;
input x11;
input x12;
input x13;
input x14;
input x15;
input x16;
input x17;
input x18;
input x19;
input x20;
input x21;
input x22;
input x23;
input x24;
input x25;
input x26;
input x27;
input x28;
input x29;
input x30;
input x31;
input x32;
input x33;
input x34;
input x35;
input x36;
input x37;
input x38;
input x39;
input x40;
input x41;
input x42;
input x43;
input x44;
input x45;
input x46;
input x47;
input x48;
input x49;
input x50;
input x51;
input x52;
input x53;
input x54;
input x55;
input x56;
input x57;
input x58;
input x59;
input x60;
input x61;
input x62;
input x63;
input x64;
input x65;
input x66;
input x67;
input x68;
input x69;
input x70;
input x71;
input x72;
input x73;
input x74;
input x75;
input x76;
input x77;
input x78;
input x79;
input x80;
input x81;
input x82;
input x83;
input x84;
input x85;
input x86;
input x87;
input x88;
input x89;
input x90;
input x91;
input x92;
input x93;
input x94;
input x95;
input x96;
input x97;
input x98;
input x99;
input x100;
input x101;
input x102;
input x103;
input x104;
input x105;
input x106;
input x107;
input x108;
input x109;
input x110;
input x111;
input x112;
input x113;
input x114;
input x115;
input x116;
input x117;
input x118;
input x119;
input x120;
input x121;
input x122;
input x123;
input x124;
input x125;
input x126;
input x127;
input x128;
input x129;
input x130;
input x131;
input x132;
input x133;
input x134;
input x135;
input x136;
input x137;
input x138;
input x139;
input x140;
input x141;
input x142;
input x143;
input x144;
input x145;
input x146;
input x147;
input x148;
input x149;
input x150;
input x151;
input x152;
input x153;
input x154;
input x155;
input x156;
input x157;
input x158;
input x159;
input x160;
input x161;
input x162;
input x163;
input x164;
input x165;
input x166;
input x167;
input x168;
input x169;
input x170;
input x171;
input x172;
input x173;
input x174;
input x175;
input x176;
input x177;
input x178;
input x179;
input x180;
input x181;
input x182;
input x183;
input x184;
input x185;
input x186;
input x187;
input x188;
input x189;
input x190;
input x191;
input x192;
input x193;
input x194;
input x195;
input x196;
input x197;
input x198;
input x199;
input x200;
input x201;
input x202;
input x203;
input x204;
input x205;
input x206;
input x207;
input x208;
input x209;
input x210;
input x211;
input x212;
input x213;
input x214;
input x215;
input x216;
input x217;
input x218;
input x219;
input x220;
input x221;
input x222;
input x223;
input x224;
input x225;
input x226;
input x227;
input x228;
input x229;
input x230;
input x231;
input x232;
input x233;
input x234;
input x235;
input x236;
input x237;
input x238;
input x239;
input x240;
input x241;
input x242;
input x243;
input x244;
input x245;
input x246;
input x247;
input x248;
input x249;
input x250;
input x251;
input x252;
input x253;
input x254;
input x255;
input x256;
input x257;
input x258;
input x259;
input x260;
input x261;
input x262;
input x263;
input x264;
input x265;
input x266;
input x267;
input x268;
input x269;
input x270;
input x271;
input x272;
input x273;
input x274;
input x275;
input x276;
input x277;
input x278;
input x279;
input x280;
input x281;
input x282;
input x283;
input x284;
input x285;
input x286;
input x287;
input x288;
input x289;
input x290;
input x291;
input x292;
input x293;
input x294;
input x295;
input x296;
input x297;
input x298;
input x299;
input x300;
input x301;
input x302;
input x303;
input x304;
input x305;
input x306;
input x307;
input x308;
input x309;
input x310;
input x311;
input x312;
input x313;
input x314;
input x315;
input x316;
input x317;
input x318;
input x319;
input x320;
input x321;
input x322;
input x323;
input x324;
input x325;
input x326;
input x327;
input x328;
input x329;
input x330;
input x331;
input x332;
input x333;
input x334;
input x335;
input x336;
input x337;
input x338;
input x339;
input x340;
input x341;
input x342;
input x343;
input x344;
input x345;
input x346;
input x347;
input x348;
input x349;
input x350;
input x351;
input x352;
input x353;
input x354;
input x355;
input x356;
input x357;
input x358;
input x359;
input x360;
input x361;
input x362;
input x363;
input x364;
input x365;
input x366;
input x367;
input x368;
input x369;
input x370;
input x371;
input x372;
input x373;
input x374;
input x375;
input x376;
input x377;
input x378;
input x379;
input x380;
input x381;
input x382;
input x383;
input x384;
input x385;
input x386;
input x387;
input x388;
input x389;
input x390;
input x391;
input x392;
input x393;
input x394;
input x395;
input x396;
input x397;
input x398;
input x399;
input x400;
input x401;
input x402;
input x403;
input x404;
input x405;
input x406;
input x407;
input x408;
input x409;
input x410;
input x411;
input x412;
input x413;
input x414;
input x415;
input x416;
input x417;
input x418;
input x419;
input x420;
input x421;
input x422;
input x423;
input x424;
input x425;
input x426;
input x427;
input x428;
input x429;
input x430;
input x431;
input x432;
input x433;
input x434;
input x435;
input x436;
input x437;
input x438;
input x439;
input x440;
input x441;
input x442;
input x443;
input x444;
input x445;
input x446;
input x447;
input x448;
input x449;
input x450;
input x451;
input x452;
input x453;
input x454;
input x455;
input x456;
input x457;
input x458;
input x459;
input x460;
input x461;
input x462;
input x463;
input x464;
input x465;
input x466;
input x467;
input x468;
input x469;
input x470;
input x471;
input x472;
input x473;
input x474;
input x475;
input x476;
input x477;
input x478;
input x479;
input x480;
input x481;
input x482;
input x483;
input x484;
input x485;
input x486;
input x487;
input x488;
input x489;
input x490;
input x491;
input x492;
input x493;
input x494;
input x495;
input x496;
input x497;
input x498;
input x499;
input x500;
input x501;
input x502;
input x503;
input x504;
input x505;
input x506;
input x507;
input x508;
input x509;
input x510;
input x511;
input x512;
input x513;
input x514;
input x515;
input x516;
input x517;
input x518;
input x519;
input x520;
input x521;
input x522;
input x523;
input x524;
input x525;
input x526;
input x527;
input x528;
input x529;
input x530;
input x531;
input x532;
input x533;
input x534;
input x535;
input x536;
input x537;
input x538;
input x539;
input x540;
input x541;
input x542;
input x543;
input x544;
input x545;
input x546;
input x547;
input x548;
input x549;
input x550;
input x551;
input x552;
input x553;
input x554;
input x555;
input x556;
input x557;
input x558;
input x559;
input x560;
input x561;
input x562;
input x563;
input x564;
input x565;
input x566;
input x567;
input x568;
input x569;
input x570;
input x571;
input x572;
input x573;
input x574;
input x575;
input x576;
input x577;
input x578;
input x579;
input x580;
input x581;
input x582;
input x583;
input x584;
input x585;
input x586;
input x587;
input x588;
input x589;
input x590;
input x591;
input x592;
input x593;
input x594;
input x595;
input x596;
input x597;
input x598;
input x599;
input x600;
input x601;
input x602;
input x603;
input x604;
input x605;
input x606;
input x607;
input x608;
input x609;
input x610;
input x611;
input x612;
input x613;
input x614;
input x615;
input x616;
input x617;
input x618;
input x619;
input x620;
input x621;
input x622;
input x623;
input x624;
input x625;
input x626;
input x627;
input x628;
input x629;
input x630;
input x631;
input x632;
input x633;
input x634;
input x635;
input x636;
input x637;
input x638;
input x639;
input x640;
input x641;
input x642;
input x643;
input x644;
input x645;
input x646;
input x647;
input x648;
input x649;
input x650;
input x651;
input x652;
input x653;
input x654;
input x655;
input x656;
input x657;
input x658;
input x659;
input x660;
input x661;
input x662;
input x663;
input x664;
input x665;
input x666;
input x667;
input x668;
input x669;
input x670;
input x671;
input x672;
input x673;
input x674;
input x675;
input x676;
input x677;
input x678;
input x679;
input x680;
input x681;
input x682;
input x683;
input x684;
input x685;
input x686;
input x687;
input x688;
input x689;
input x690;
input x691;
input x692;
input x693;
input x694;
input x695;
input x696;
input x697;
input x698;
input x699;
input x700;
input x701;
input x702;
input x703;
input x704;
input x705;
input x706;
input x707;
input x708;
input x709;
input x710;
input x711;
input x712;
input x713;
input x714;
input x715;
input x716;
input x717;
input x718;
input x719;
input x720;
input x721;
input x722;
input x723;
input x724;
input x725;
input x726;
input x727;
input x728;
input x729;
input x730;
input x731;
input x732;
input x733;
input x734;
input x735;
input x736;
input x737;
input x738;
input x739;
input x740;
input x741;
input x742;
input x743;
input x744;
input x745;
input x746;
input x747;
input x748;
input x749;
input x750;
input x751;
input x752;
input x753;
input x754;
input x755;
input x756;
input x757;
input x758;
input x759;
input x760;
input x761;
input x762;
input x763;
input x764;
input x765;
input x766;
input x767;
input x768;
input x769;
input x770;
input x771;
input x772;
input x773;
input x774;
input x775;
input x776;
input x777;
input x778;
input x779;
input x780;
input x781;
input x782;
input x783;
input x784;
input x785;
input x786;
input x787;
input x788;
input x789;
input x790;
input x791;
input x792;
input x793;
input x794;
input x795;
input x796;
input x797;
input x798;
input x799;
input x800;
input x801;
input x802;
input x803;
input x804;
input x805;
input x806;
input x807;
input x808;
input x809;
input x810;
input x811;
input x812;
input x813;
input x814;
input x815;
input x816;
input x817;
input x818;
input x819;
input x820;
input x821;
input x822;
input x823;
input x824;
input x825;
input x826;
input x827;
input x828;
input x829;
input x830;
input x831;
input x832;
input x833;
input x834;
input x835;
input x836;
input x837;
input x838;
input x839;
input x840;
input x841;
input x842;
input x843;
input x844;
input x845;
input x846;
input x847;
input x848;
input x849;
input x850;
input x851;
input x852;
input x853;
input x854;
input x855;
input x856;
input x857;
input x858;
input x859;
input x860;
input x861;
input x862;
input x863;
input x864;
input x865;
input x866;
input x867;
input x868;
input x869;
input x870;
input x871;
input x872;
input x873;
input x874;
input x875;
input x876;
input x877;
input x878;
input x879;
input x880;
input x881;
input x882;
input x883;
input x884;
input x885;
input x886;
input x887;
input x888;
input x889;
input x890;
input x891;
input x892;
input x893;
input x894;
input x895;
input x896;
input x897;
input x898;
input x899;
input x900;
input x901;
input x902;
input x903;
input x904;
input x905;
input x906;
input x907;
input x908;
input x909;
input x910;
input x911;
input x912;
input x913;
input x914;
input x915;
input x916;
input x917;
input x918;
input x919;
input x920;
input x921;
input x922;
input x923;
input x924;
input x925;
input x926;
input x927;
input x928;
input x929;
input x930;
input x931;
input x932;
input x933;
input x934;
input x935;
input x936;
input x937;
input x938;
input x939;
input x940;
input x941;
input x942;
input x943;
input x944;
input x945;
input x946;
input x947;
input x948;
input x949;
input x950;
input x951;
input x952;
input x953;
input x954;
input x955;
input x956;
input x957;
input x958;
input x959;
input x960;
input x961;
input x962;
input x963;
input x964;
input x965;
input x966;
input x967;
input x968;
input x969;
input x970;
input x971;
input x972;
input x973;
input x974;
input x975;
input x976;
input x977;
input x978;
input x979;
input x980;
input x981;
input x982;
input x983;
input x984;
input x985;
input x986;
input x987;
input x988;
input x989;
input x990;
input x991;
input x992;
input x993;
input x994;
input x995;
input x996;
input x997;
input x998;
input x999;
input x1000;
input x1001;
input x1002;
input x1003;
input x1004;
input x1005;
input x1006;
input x1007;
input x1008;
input x1009;
input x1010;
input x1011;
input x1012;
input x1013;
input x1014;
input x1015;
input x1016;
input x1017;
input x1018;
input x1019;
input x1020;
input x1021;
input x1022;
input x1023;
input x1024;
input x1025;
input x1026;
input x1027;
input x1028;
input x1029;
input x1030;
input x1031;
input x1032;
input x1033;
input x1034;
input x1035;
input x1036;
input x1037;
input x1038;
input x1039;
input x1040;
input x1041;
input x1042;
input x1043;
input x1044;
input x1045;
input x1046;
input x1047;
input x1048;
input x1049;
input x1050;
input x1051;
input x1052;
input x1053;
input x1054;
input x1055;
input x1056;
input x1057;
input x1058;
input x1059;
input x1060;
input x1061;
input x1062;
input x1063;
input x1064;
input x1065;
input x1066;
input x1067;
input x1068;
input x1069;
input x1070;
input x1071;
input x1072;
input x1073;
input x1074;
input x1075;
input x1076;
input x1077;
input x1078;
input x1079;
input x1080;
input x1081;
input x1082;
input x1083;
input x1084;
input x1085;
input x1086;
input x1087;
input x1088;
input x1089;
input x1090;
input x1091;
input x1092;
input x1093;
input x1094;
input x1095;
input x1096;
input x1097;
input x1098;
input x1099;
input x1100;
input x1101;
input x1102;
input x1103;
input x1104;
input x1105;
input x1106;
input x1107;
input x1108;
input x1109;
input x1110;
input x1111;
input x1112;
input x1113;
input x1114;
input x1115;
input x1116;
input x1117;
input x1118;
input x1119;
input x1120;
input x1121;
input x1122;
input x1123;
input x1124;
input x1125;
input x1126;
input x1127;
input x1128;
input x1129;
input x1130;
output c0219;
output c1253;
output c5138;
output c4199;
output c10;
output c0130;
output c6133;
output c7113;
output c3121;
output c6236;
output c0182;
output c4187;
output c650;
output c41;
output c7299;
output c5289;
output c0298;
output c5161;
output c698;
output c3284;
output c454;
output c4250;
output c737;
output c58;
output c332;
output c134;
output c4181;
output c468;
output c1279;
output c032;
output c7220;
output c6164;
output c0185;
output c348;
output c0217;
output c2171;
output c5288;
output c21;
output c4198;
output c145;
output c378;
output c358;
output c399;
output c55;
output c116;
output c4221;
output c7159;
output c270;
output c7133;
output c1165;
output c3279;
output c578;
output c4269;
output c4151;
output c6285;
output c3189;
output c492;
output c2142;
output c1299;
output c7161;
output c686;
output c7285;
output c247;
output c7176;
output c0214;
output c7125;
output c3162;
output c4170;
output c2274;
output c1297;
output c7116;
output c3133;
output c721;
output c15;
output c4243;
output c5235;
output c0104;
output c722;
output c370;
output c572;
output c5222;
output c532;
output c1150;
output c5199;
output c038;
output c335;
output c513;
output c123;
output c5230;
output c651;
output c6124;
output c147;
output c050;
output c6225;
output c3228;
output c3215;
output c4291;
output c6202;
output c2293;
output c210;
output c1184;
output c276;
output c4185;
output c2165;
output c3273;
output c214;
output c3122;
output c6186;
output c0200;
output c2117;
output c6138;
output c7251;
output c2280;
output c0238;
output c1124;
output c7289;
output c039;
output c057;
output c2109;
output c5112;
output c3288;
output c4176;
output c3207;
output c6221;
output c23;
output c798;
output c7157;
output c2249;
output c33;
output c3219;
output c556;
output c7249;
output c5187;
output c5272;
output c4147;
output c7164;
output c5197;
output c13;
output c0294;
output c7150;
output c125;
output c3244;
output c021;
output c727;
output c0276;
output c2262;
output c158;
output c1132;
output c2284;
output c1209;
output c4165;
output c6166;
output c3221;
output c498;
output c0113;
output c146;
output c460;
output c5225;
output c2224;
output c2244;
output c1206;
output c6156;
output c6281;
output c740;
output c1180;
output c597;
output c2217;
output c222;
output c1200;
output c6110;
output c0146;
output c4188;
output c739;
output c1264;
output c1123;
output c345;
output c539;
output c4222;
output c3270;
output c632;
output c7278;
output c196;
output c6289;
output c5170;
output c6226;
output c3124;
output c1273;
output c777;
output c6299;
output c220;
output c5265;
output c7221;
output c218;
output c0132;
output c5105;
output c0189;
output c6102;
output c7257;
output c3182;
output c494;
output c379;
output c7224;
output c6224;
output c052;
output c0179;
output c133;
output c7228;
output c769;
output c475;
output c575;
output c5132;
output c212;
output c096;
output c176;
output c664;
output c0291;
output c1213;
output c6198;
output c687;
output c0259;
output c1160;
output c3136;
output c1278;
output c618;
output c1274;
output c3267;
output c4200;
output c4173;
output c2164;
output c248;
output c7281;
output c234;
output c2172;
output c794;
output c411;
output c699;
output c5278;
output c3138;
output c2273;
output c779;
output c09;
output c3141;
output c1283;
output c476;
output c483;
output c1269;
output c7219;
output c7296;
output c1291;
output c2237;
output c173;
output c4201;
output c464;
output c245;
output c4215;
output c4264;
output c4274;
output c2139;
output c4161;
output c7202;
output c751;
output c0117;
output c7162;
output c3106;
output c184;
output c5143;
output c510;
output c3283;
output c59;
output c3179;
output c1227;
output c3140;
output c6119;
output c4276;
output c3195;
output c6290;
output c3161;
output c4137;
output c4116;
output c6120;
output c6151;
output c7141;
output c180;
output c1252;
output c5208;
output c0203;
output c782;
output c012;
output c2182;
output c2207;
output c19;
output c393;
output c536;
output c7290;
output c251;
output c3236;
output c0241;
output c5211;
output c4225;
output c0224;
output c770;
output c0153;
output c5109;
output c6175;
output c1192;
output c5104;
output c1151;
output c3127;
output c199;
output c0122;
output c4156;
output c6271;
output c768;
output c431;
output c2166;
output c7256;
output c5145;
output c0293;
output c3298;
output c7172;
output c2196;
output c14;
output c5209;
output c7232;
output c7269;
output c0116;
output c111;
output c5251;
output c718;
output c0147;
output c6167;
output c322;
output c5231;
output c4183;
output c3278;
output c6170;
output c74;
output c4229;
output c1282;
output c5136;
output c1186;
output c2153;
output c619;
output c6297;
output c5174;
output c3252;
output c1163;
output c450;
output c3134;
output c5244;
output c4235;
output c5139;
output c6114;
output c6192;
output c1289;
output c5134;
output c0149;
output c7143;
output c37;
output c0204;
output c6172;
output c5146;
output c7112;
output c17;
output c0143;
output c070;
output c663;
output c3282;
output c0159;
output c3276;
output c479;
output c5121;
output c2180;
output c221;
output c7124;
output c7265;
output c274;
output c1233;
output c645;
output c642;
output c1140;
output c5293;
output c261;
output c5290;
output c238;
output c7233;
output c4263;
output c3254;
output c48;
output c3253;
output c7155;
output c2113;
output c452;
output c489;
output c581;
output c331;
output c3105;
output c294;
output c4267;
output c5178;
output c7167;
output c5218;
output c5204;
output c0234;
output c3172;
output c242;
output c5198;
output c516;
output c535;
output c4298;
output c680;
output c2185;
output c372;
output c377;
output c0161;
output c0262;
output c669;
output c4106;
output c0281;
output c361;
output c3251;
output c0295;
output c1219;
output c4233;
output c398;
output c5295;
output c0180;
output c0134;
output c6275;
output c2108;
output c5229;
output c6242;
output c2211;
output c2299;
output c416;
output c570;
output c7139;
output c2140;
output c5297;
output c3110;
output c3292;
output c47;
output c195;
output c4211;
output c71;
output c5245;
output c098;
output c423;
output c2122;
output c693;
output c0198;
output c7110;
output c4287;
output c4252;
output c235;
output c7207;
output c6288;
output c066;
output c433;
output c1183;
output c4209;
output c1137;
output c758;
output c254;
output c4132;
output c4139;
output c5129;
output c0272;
output c0243;
output c4281;
output c2227;
output c1194;
output c6274;
output c0120;
output c5264;
output c3203;
output c1272;
output c6130;
output c4133;
output c5206;
output c76;
output c692;
output c088;
output c3148;
output c7166;
output c353;
output c3143;
output c1136;
output c00;
output c3116;
output c3152;
output c7208;
output c040;
output c112;
output c3209;
output c6195;
output c22;
output c2186;
output c3234;
output c4149;
output c3243;
output c5276;
output c3197;
output c312;
output c323;
output c589;
output c5151;
output c7126;
output c1158;
output c0154;
output c2214;
output c477;
output c3232;
output c463;
output c5113;
output c5281;
output c3206;
output c0229;
output c7200;
output c4193;
output c4128;
output c6181;
output c5268;
output c2110;
output c387;
output c1131;
output c3131;
output c140;
output c042;
output c065;
output c480;
output c3247;
output c491;
output c7226;
output c121;
output c4142;
output c7185;
output c7227;
output c5182;
output c1107;
output c5190;
output c4114;
output c4195;
output c0183;
output c048;
output c075;
output c0158;
output c314;
output c627;
output c7122;
output c4240;
output c493;
output c3125;
output c6251;
output c641;
output c6270;
output c229;
output c4277;
output c397;
output c0136;
output c7171;
output c243;
output c1142;
output c1118;
output c4294;
output c5115;
output c6207;
output c6272;
output c559;
output c32;
output c3132;
output c1152;
output c657;
output c689;
output c6105;
output c6174;
output c1189;
output c3220;
output c2193;
output c316;
output c2124;
output c149;
output c1268;
output c3275;
output c2145;
output c634;
output c3107;
output c067;
output c2132;
output c453;
output c177;
output c1281;
output c5216;
output c7198;
output c533;
output c7206;
output c1134;
output c0196;
output c519;
output c045;
output c6171;
output c2102;
output c120;
output c5262;
output c428;
output c5186;
output c1292;
output c2163;
output c4120;
output c5176;
output c1256;
output c557;
output c0226;
output c778;
output c0218;
output c3216;
output c7252;
output c0285;
output c3184;
output c4270;
output c2136;
output c2178;
output c172;
output c78;
output c339;
output c2160;
output c246;
output c5116;
output c156;
output c0274;
output c7115;
output c435;
output c036;
output c7111;
output c0115;
output c2295;
output c781;
output c2255;
output c4228;
output c3103;
output c4191;
output c3272;
output c4121;
output c329;
output c5131;
output c451;
output c613;
output c3249;
output c0275;
output c797;
output c750;
output c2159;
output c4248;
output c5158;
output c390;
output c0249;
output c3150;
output c4282;
output c2148;
output c164;
output c6142;
output c053;
output c1277;
output c290;
output c5202;
output c371;
output c5128;
output c161;
output c6122;
output c2288;
output c5255;
output c671;
output c5155;
output c1280;
output c6250;
output c1231;
output c2278;
output c2257;
output c4205;
output c5201;
output c61;
output c6239;
output c4148;
output c3169;
output c6222;
output c4157;
output c4126;
output c759;
output c2246;
output c2215;
output c6121;
output c6169;
output c1254;
output c3277;
output c2183;
output c1104;
output c010;
output c4158;
output c4101;
output c5296;
output c3144;
output c138;
output c673;
output c3155;
output c6134;
output c3257;
output c4146;
output c0118;
output c5210;
output c1246;
output c26;
output c1122;
output c1290;
output c4164;
output c5181;
output c1110;
output c4179;
output c130;
output c0223;
output c414;
output c612;
output c670;
output c0192;
output c0145;
output c4135;
output c2233;
output c5154;
output c7214;
output c7240;
output c5184;
output c320;
output c328;
output c3214;
output c1237;
output c7277;
output c497;
output c1135;
output c631;
output c041;
output c730;
output c4265;
output c4254;
output c2285;
output c2112;
output c394;
output c082;
output c5253;
output c6205;
output c34;
output c4175;
output c3237;
output c644;
output c1211;
output c3293;
output c0142;
output c6232;
output c2268;
output c044;
output c6152;
output c090;
output c5233;
output c3229;
output c0282;
output c469;
output c6162;
output c7298;
output c7268;
output c2167;
output c637;
output c776;
output c3218;
output c594;
output c1262;
output c3146;
output c2222;
output c3111;
output c2188;
output c5141;
output c352;
output c7271;
output c4143;
output c656;
output c6103;
output c6154;
output c616;
output c3199;
output c6223;
output c3290;
output c061;
output c117;
output c7130;
output c461;
output c4238;
output c0232;
output c4256;
output c6267;
output c6111;
output c1170;
output c175;
output c1263;
output c6257;
output c324;
output c337;
output c6140;
output c262;
output c2208;
output c167;
output c0267;
output c2168;
output c343;
output c7294;
output c2232;
output c118;
output c646;
output c6287;
output c756;
output c719;
output c7118;
output c771;
output c0206;
output c019;
output c183;
output c565;
output c0252;
output c255;
output c2204;
output c1169;
output c6282;
output c062;
output c1275;
output c2298;
output c4289;
output c258;
output c0209;
output c30;
output c580;
output c1109;
output c2128;
output c554;
output c2118;
output c2245;
output c3296;
output c0127;
output c3289;
output c7107;
output c5196;
output c5246;
output c2212;
output c0207;
output c2270;
output c056;
output c4154;
output c659;
output c7182;
output c2236;
output c035;
output c0254;
output c2252;
output c4266;
output c0169;
output c5126;
output c5277;
output c313;
output c1224;
output c5111;
output c0106;
output c1127;
output c295;
output c4241;
output c185;
output c1156;
output c1255;
output c0257;
output c5147;
output c667;
output c160;
output c4226;
output c647;
output c577;
output c064;
output c598;
output c6125;
output c2281;
output c7146;
output c0155;
output c696;
output c60;
output c544;
output c5167;
output c579;
output c1121;
output c5150;
output c68;
output c7108;
output c0255;
output c521;
output c5207;
output c793;
output c4192;
output c2158;
output c364;
output c374;
output c789;
output c6254;
output c3212;
output c3266;
output c2105;
output c5120;
output c2169;
output c472;
output c7201;
output c2195;
output c588;
output c3178;
output c260;
output c1129;
output c5217;
output c7135;
output c0278;
output c1216;
output c3118;
output c355;
output c439;
output c485;
output c1113;
output c351;
output c283;
output c0220;
output c2272;
output c51;
output c2170;
output c165;
output c655;
output c382;
output c749;
output c2239;
output c3168;
output c094;
output c287;
output c3213;
output c5127;
output c2251;
output c0227;
output c6245;
output c6199;
output c587;
output c7204;
output c2275;
output c7194;
output c6163;
output c6244;
output c3281;
output c1190;
output c043;
output c0190;
output c2152;
output c4118;
output c5172;
output c7272;
output c5180;
output c4214;
output c148;
output c6279;
output c0260;
output c457;
output c590;
output c53;
output c2101;
output c2265;
output c4283;
output c63;
output c5152;
output c783;
output c5169;
output c267;
output c2175;
output c0213;
output c092;
output c2242;
output c289;
output c31;
output c735;
output c5254;
output c3258;
output c1159;
output c2123;
output c660;
output c764;
output c2241;
output c4141;
output c6217;
output c444;
output c2216;
output c526;
output c7180;
output c745;
output c4236;
output c4131;
output c690;
output c6136;
output c427;
output c6296;
output c788;
output c169;
output c319;
output c3194;
output c5287;
output c599;
output c6208;
output c6231;
output c368;
output c4104;
output c6213;
output c380;
output c4258;
output c4224;
output c6190;
output c432;
output c5189;
output c6249;
output c1167;
output c253;
output c7273;
output c5292;
output c4145;
output c2297;
output c2261;
output c4136;
output c078;
output c1220;
output c0253;
output c7203;
output c3104;
output c2210;
output c349;
output c5135;
output c0231;
output c4177;
output c5164;
output c1146;
output c5142;
output c1222;
output c3204;
output c014;
output c1271;
output c731;
output c7129;
output c7173;
output c279;
output c189;
output c2125;
output c4174;
output c6259;
output c241;
output c06;
output c27;
output c1196;
output c5248;
output c3262;
output c3126;
output c4124;
output c49;
output c3294;
output c216;
output c1210;
output c760;
output c2225;
output c293;
output c7237;
output c0290;
output c2229;
output c540;
output c7222;
output c263;
output c266;
output c4134;
output c5194;
output c4100;
output c6144;
output c7276;
output c3246;
output c020;
output c350;
output c638;
output c6161;
output c5103;
output c3139;
output c4286;
output c058;
output c676;
output c4261;
output c197;
output c7218;
output c5234;
output c2279;
output c159;
output c142;
output c211;
output c1130;
output c5215;
output c3291;
output c6182;
output c3271;
output c675;
output c4260;
output c357;
output c7242;
output c3217;
output c2276;
output c4212;
output c0222;
output c0279;
output c6113;
output c333;
output c115;
output c186;
output c5291;
output c2129;
output c7261;
output c512;
output c3129;
output c013;
output c44;
output c1203;
output c5259;
output c7120;
output c213;
output c016;
output c514;
output c233;
output c0288;
output c5221;
output c4245;
output c317;
output c3286;
output c1173;
output c7184;
output c4140;
output c1266;
output c561;
output c055;
output c1119;
output c2127;
output c746;
output c1221;
output c086;
output c5108;
output c1197;
output c697;
output c6212;
output c1177;
output c7297;
output c079;
output c5157;
output c574;
output c7103;
output c7142;
output c5117;
output c3239;
output c2219;
output c4255;
output c1181;
output c4272;
output c3142;
output c6132;
output c6178;
output c4259;
output c0184;
output c192;
output c3259;
output c4249;
output c026;
output c534;
output c029;
output c487;
output c467;
output c0172;
output c528;
output c5160;
output c5193;
output c1101;
output c16;
output c518;
output c7128;
output c0150;
output c4117;
output c0195;
output c366;
output c4206;
output c5122;
output c0193;
output c6216;
output c1285;
output c0248;
output c7286;
output c7134;
output c280;
output c1125;
output c7245;
output c3156;
output c4246;
output c720;
output c1248;
output c7239;
output c1164;
output c520;
output c7193;
output c73;
output c3187;
output c3223;
output c269;
output c0233;
output c129;
output c470;
output c3108;
output c7179;
output c6139;
output c5185;
output c6280;
output c6183;
output c679;
output c0266;
output c6284;
output c141;
output c2291;
output c499;
output c7248;
output c7149;
output c135;
output c5271;
output c3287;
output c0139;
output c2116;
output c473;
output c592;
output c6234;
output c0121;
output c678;
output c7190;
output c1153;
output c227;
output c5279;
output c6135;
output c6292;
output c1260;
output c7205;
output c1114;
output c1174;
output c6241;
output c3240;
output c028;
output c1182;
output c4244;
output c7199;
output c419;
output c711;
output c424;
output c0162;
output c3114;
output c5227;
output c567;
output c2226;
output c347;
output c542;
output c69;
output c38;
output c0131;
output c591;
output c430;
output c547;
output c3163;
output c1191;
output c658;
output c02;
output c537;
output c3145;
output c373;
output c5294;
output c1241;
output c43;
output c356;
output c2200;
output c5166;
output c1187;
output c0191;
output c4189;
output c7105;
output c684;
output c7192;
output c0100;
output c6118;
output c0160;
output c063;
output c2107;
output c4232;
output c6180;
output c6230;
output c3166;
output c2181;
output c6235;
output c1247;
output c4115;
output c7160;
output c224;
output c6108;
output c2202;
output c5162;
output c555;
output c6187;
output c635;
output c1166;
output c3268;
output c1204;
output c0168;
output c5130;
output c1175;
output c6298;
output c2256;
output c0268;
output c456;
output c443;
output c2162;
output c465;
output c7152;
output c298;
output c155;
output c2157;
output c4251;
output c7136;
output c278;
output c5195;
output c0215;
output c6127;
output c3147;
output c7260;
output c0221;
output c6277;
output c346;
output c426;
output c6184;
output c775;
output c6252;
output c4297;
output c344;
output c236;
output c7241;
output c1240;
output c1257;
output c264;
output c07;
output c6240;
output c7186;
output c1111;
output c639;
output c018;
output c0171;
output c7209;
output c7195;
output c083;
output c6165;
output c1128;
output c273;
output c0107;
output c630;
output c5156;
output c2177;
output c4210;
output c2290;
output c363;
output c2254;
output c2104;
output c7145;
output c0299;
output c1139;
output c0271;
output c1235;
output c6238;
output c7254;
output c4122;
output c3160;
output c478;
output c7284;
output c330;
output c5205;
output c6233;
output c6168;
output c7183;
output c5102;
output c170;
output c3113;
output c0277;
output c1228;
output c568;
output c677;
output c2235;
output c2263;
output c0124;
output c437;
output c0283;
output c194;
output c3211;
output c5137;
output c04;
output c562;
output c0188;
output c7274;
output c369;
output c45;
output c2179;
output c5214;
output c2135;
output c0105;
output c097;
output c4182;
output c714;
output c0244;
output c0289;
output c383;
output c6262;
output c790;
output c755;
output c2203;
output c2267;
output c2120;
output c4295;
output c023;
output c3256;
output c228;
output c66;
output c7175;
output c442;
output c027;
output c113;
output c5191;
output c4163;
output c4180;
output c531;
output c011;
output c5213;
output c736;
output c7197;
output c1223;
output c672;
output c0126;
output c665;
output c05;
output c5260;
output c515;
output c1145;
output c1226;
output c5123;
output c386;
output c4194;
output c448;
output c0211;
output c5168;
output c7102;
output c7127;
output c179;
output c522;
output c034;
output c7267;
output c2134;
output c3153;
output c458;
output c3198;
output c2260;
output c5153;
output c136;
output c2282;
output c0135;
output c7283;
output c03;
output c1218;
output c18;
output c734;
output c4196;
output c1296;
output c35;
output c087;
output c6137;
output c3205;
output c488;
output c6157;
output c4253;
output c1176;
output c3175;
output c4296;
output c649;
output c1229;
output c1249;
output c4123;
output c5243;
output c743;
output c2199;
output c384;
output c3181;
output c546;
output c767;
output c742;
output c2191;
output c6256;
output c585;
output c2144;
output c418;
output c282;
output c694;
output c2190;
output c633;
output c5285;
output c1154;
output c1232;
output c1178;
output c2286;
output c4125;
output c7138;
output c7247;
output c6291;
output c766;
output c2121;
output c4105;
output c215;
output c126;
output c12;
output c5163;
output c1293;
output c01;
output c682;
output c037;
output c2155;
output c2151;
output c3123;
output c4150;
output c780;
output c2223;
output c774;
output c524;
output c420;
output c4219;
output c2130;
output c6265;
output c051;
output c2154;
output c5223;
output c0119;
output c5149;
output c6126;
output c1242;
output c3261;
output c6158;
output c3130;
output c0264;
output c681;
output c527;
output c0141;
output c0245;
output c5220;
output c413;
output c4280;
output c3185;
output c5179;
output c069;
output c6220;
output c7119;
output c272;
output c6286;
output c318;
output c5110;
output c297;
output c77;
output c6188;
output c447;
output c7295;
output c2194;
output c2289;
output c0181;
output c7106;
output c747;
output c1225;
output c4160;
output c4102;
output c754;
output c325;
output c410;
output c4271;
output c563;
output c310;
output c292;
output c5107;
output c391;
output c2221;
output c2228;
output c3264;
output c0280;
output c7181;
output c1198;
output c362;
output c7264;
output c017;
output c446;
output c5269;
output c7163;
output c7191;
output c7211;
output c360;
output c0235;
output c1276;
output c611;
output c1138;
output c1162;
output c2259;
output c388;
output c733;
output c122;
output c3248;
output c3280;
output c5133;
output c4208;
output c490;
output c661;
output c5118;
output c5250;
output c713;
output c2131;
output c3233;
output c1207;
output c2213;
output c6143;
output c025;
output c151;
output c582;
output c2106;
output c662;
output c412;
output c226;
output c3235;
output c2253;
output c5175;
output c4113;
output c6117;
output c2150;
output c0174;
output c288;
output c4217;
output c0216;
output c6293;
output c2198;
output c7187;
output c2292;
output c7258;
output c7244;
output c367;
output c4103;
output c5258;
output c342;
output c3226;
output c030;
output c5299;
output c786;
output c093;
output c3241;
output c2143;
output c054;
output c3157;
output c0173;
output c1270;
output c541;
output c392;
output c417;
output c4223;
output c4129;
output c1243;
output c1149;
output c796;
output c2137;
output c0284;
output c3188;
output c359;
output c4184;
output c163;
output c7238;
output c610;
output c0250;
output c75;
output c1251;
output c7189;
output c6148;
output c0197;
output c1141;
output c389;
output c787;
output c7140;
output c077;
output c1143;
output c471;
output c321;
output c4172;
output c586;
output c7196;
output c7156;
output c326;
output c4292;
output c6260;
output c2138;
output c7177;
output c7293;
output c571;
output c0242;
output c29;
output c3117;
output c614;
output c1298;
output c6100;
output c7234;
output c668;
output c7292;
output c7231;
output c334;
output c6123;
output c4293;
output c7131;
output c6261;
output c5114;
output c621;
output c2220;
output c6215;
output c573;
output c0102;
output c2243;
output c4239;
output c5274;
output c2111;
output c5256;
output c265;
output c2271;
output c3274;
output c748;
output c6264;
output c2205;
output c7223;
output c395;
output c08;
output c230;
output c2209;
output c652;
output c6219;
output c1265;
output c0144;
output c6258;
output c3255;
output c2147;
output c3208;
output c7235;
output c2296;
output c4213;
output c2192;
output c1295;
output c1157;
output c710;
output c1245;
output c6294;
output c728;
output c2234;
output c6278;
output c7154;
output c422;
output c762;
output c250;
output c5242;
output c0205;
output c3102;
output c150;
output c726;
output c4216;
output c2250;
output c0133;
output c0225;
output c0194;
output c5200;
output c685;
output c1168;
output c57;
output c4144;
output c7151;
output c4290;
output c6200;
output c4220;
output c67;
output c0128;
output c791;
output c3119;
output c271;
output c4186;
output c772;
output c5280;
output c4108;
output c7153;
output c550;
output c6263;
output c2231;
output c0265;
output c3186;
output c5203;
output c256;
output c2115;
output c132;
output c523;
output c595;
output c2247;
output c538;
output c1205;
output c268;
output c0186;
output c1188;
output c3183;
output c4110;
output c285;
output c1287;
output c3158;
output c6218;
output c191;
output c336;
output c1133;
output c3128;
output c6201;
output c7212;
output c1171;
output c7148;
output c28;
output c484;
output c763;
output c198;
output c1199;
output c2201;
output c4169;
output c6155;
output c085;
output c529;
output c5183;
output c6191;
output c144;
output c4153;
output c4207;
output c315;
output c049;
output c1115;
output c640;
output c552;
output c3196;
output c3202;
output c239;
output c4130;
output c1117;
output c4167;
output c46;
output c3170;
output c059;
output c429;
output c455;
output c2189;
output c421;
output c1103;
output c4197;
output c3180;
output c084;
output c72;
output c7280;
output c1155;
output c1147;
output c636;
output c3149;
output c6283;
output c0263;
output c0286;
output c1267;
output c7217;
output c0156;
output c744;
output c5282;
output c626;
output c081;
output c4285;
output c2126;
output c4166;
output c0163;
output c6147;
output c286;
output c7109;
output c275;
output c259;
output c593;
output c1244;
output c4111;
output c7243;
output c2266;
output c154;
output c0103;
output c629;
output c6116;
output c291;
output c4138;
output c4262;
output c0137;
output c143;
output c2218;
output c7137;
output c3238;
output c0261;
output c653;
output c3176;
output c0246;
output c1215;
output c6149;
output c0175;
output c723;
output c459;
output c6128;
output c0247;
output c3200;
output c7270;
output c0292;
output c396;
output c5263;
output c2173;
output c5257;
output c3174;
output c56;
output c139;
output c643;
output c5275;
output c7114;
output c666;
output c622;
output c225;
output c223;
output c0140;
output c244;
output c0151;
output c0129;
output c6150;
output c3224;
output c095;
output c162;
output c217;
output c257;
output c4152;
output c2114;
output c080;
output c0273;
output c64;
output c65;
output c2206;
output c617;
output c7123;
output c4204;
output c3231;
output c7169;
output c5247;
output c5232;
output c6115;
output c6246;
output c738;
output c4288;
output c1250;
output c157;
output c178;
output c3227;
output c6253;
output c3109;
output c732;
output c434;
output c0256;
output c1105;
output c376;
output c40;
output c1106;
output c0152;
output c4268;
output c6197;
output c6145;
output c2161;
output c1208;
output c5270;
output c7250;
output c1238;
output c7275;
output c3230;
output c1185;
output c2294;
output c2184;
output c1236;
output c4119;
output c249;
output c152;
output c5119;
output c2248;
output c340;
output c4218;
output c237;
output c482;
output c1148;
output c281;
output c076;
output c7216;
output c7262;
output c6196;
output c0258;
output c3151;
output c0166;
output c3177;
output c481;
output c511;
output c3173;
output c071;
output c7132;
output c7253;
output c015;
output c4178;
output c153;
output c4190;
output c39;
output c3101;
output c42;
output c7282;
output c716;
output c3159;
output c0114;
output c4227;
output c7213;
output c0287;
output c2187;
output c2197;
output c625;
output c1161;
output c252;
output c5286;
output c628;
output c70;
output c127;
output c3193;
output c089;
output c338;
output c495;
output c5237;
output c137;
output c4112;
output c2174;
output c5159;
output c6189;
output c7101;
output c7255;
output c2103;
output c438;
output c1172;
output c6101;
output c219;
output c1144;
output c717;
output c6276;
output c545;
output c6185;
output c0239;
output c5144;
output c0228;
output c7168;
output c099;
output c576;
output c7230;
output c1212;
output c6176;
output c232;
output c425;
output c2156;
output c0178;
output c171;
output c548;
output c0240;
output c5228;
output c240;
output c3137;
output c1116;
output c4275;
output c7165;
output c3171;
output c0201;
output c3201;
output c046;
output c20;
output c1179;
output c6210;
output c784;
output c327;
output c4155;
output c564;
output c3297;
output c0110;
output c566;
output c2283;
output c525;
output c6209;
output c5224;
output c7174;
output c0208;
output c1234;
output c7291;
output c0167;
output c2240;
output c6173;
output c068;
output c799;
output c7147;
output c354;
output c445;
output c168;
output c381;
output c4247;
output c5284;
output c4203;
output c6237;
output c757;
output c174;
output c25;
output c5100;
output c091;
output c741;
output c0297;
output c3295;
output c6160;
output c1230;
output c6273;
output c5298;
output c0125;
output c7100;
output c0199;
output c50;
output c073;
output c1202;
output c5148;
output c436;
output c0270;
output c1126;
output c440;
output c4278;
output c5226;
output c128;
output c773;
output c6269;
output c551;
output c3260;
output c6107;
output c7144;
output c6131;
output c0165;
output c284;
output c3222;
output c6268;
output c193;
output c7225;
output c553;
output c0202;
output c4234;
output c4231;
output c5236;
output c4273;
output c24;
output c7266;
output c3269;
output c0236;
output c474;
output c277;
output c5252;
output c623;
output c688;
output c299;
output c0138;
output c2238;
output c5266;
output c119;
output c7158;
output c5238;
output c031;
output c3263;
output c3245;
output c5283;
output c3100;
output c7121;
output c0157;
output c5171;
output c52;
output c0108;
output c4299;
output c569;
output c1214;
output c110;
output c795;
output c2141;
output c2119;
output c5261;
output c3299;
output c4242;
output c7288;
output c725;
output c6193;
output c0230;
output c0269;
output c2269;
output c2230;
output c7236;
output c3120;
output c0296;
output c3115;
output c0212;
output c1284;
output c5240;
output c6104;
output c311;
output c0177;
output c3135;
output c4162;
output c674;
output c441;
output c5192;
output c4284;
output c5273;
output c4237;
output c648;
output c615;
output c0170;
output c6203;
output c166;
output c2146;
output c724;
output c5239;
output c365;
output c4109;
output c3112;
output c683;
output c131;
output c624;
output c0187;
output c6141;
output c462;
output c5101;
output c596;
output c2133;
output c5249;
output c4230;
output c296;
output c6255;
output c0109;
output c584;
output c3242;
output c2277;
output c187;
output c729;
output c415;
output c7117;
output c3165;
output c341;
output c785;
output c62;
output c1102;
output c6153;
output c654;
output c715;
output c36;
output c4107;
output c072;
output c4171;
output c792;
output c0111;
output c1261;
output c2100;
output c1193;
output c5173;
output c1120;
output c691;
output c6227;
output c765;
output c6248;
output c060;
output c695;
output c3190;
output c4257;
output c188;
output c1286;
output c047;
output c560;
output c496;
output c6228;
output c7178;
output c3164;
output c7259;
output c1258;
output c6214;
output c0210;
output c4159;
output c5140;
output c6109;
output c6243;
output c517;
output c022;
output c3167;
output c6179;
output c6211;
output c4279;
output c5241;
output c6159;
output c182;
output c753;
output c449;
output c0251;
output c1195;
output c181;
output c7229;
output c486;
output c0123;
output c5125;
output c7263;
output c2287;
output c1201;
output c3210;
output c3192;
output c0112;
output c033;
output c3225;
output c5124;
output c79;
output c0148;
output c1259;
output c54;
output c6204;
output c7104;
output c0164;
output c0176;
output c3154;
output c6112;
output c231;
output c7246;
output c0237;
output c7188;
output c7287;
output c583;
output c190;
output c1288;
output c6106;
output c7279;
output c0101;
output c620;
output c6177;
output c466;
output c1217;
output c7215;
output c4127;
output c024;
output c6266;
output c530;
output c4168;
output c712;
output c6295;
output c7170;
output c3265;
output c6129;
output c6206;
output c761;
output c1112;
output c5219;
output c549;
output c1239;
output c6247;
output c114;
output c543;
output c3285;
output c1108;
output c3191;
output c558;
output c7210;
output c752;
output c6229;
output c074;
output c4202;
output c5106;
output c5177;
output c11;
output c375;
output c5188;
output c1294;
output c2258;
output c2176;
output c2264;
output c6146;
output c2149;
output c5165;
output c124;
output c1100;
output c5212;
output c5267;
output c6194;
output c3250;
output c385;

assign c00 =  x134 &  x182 &  x206 &  x209 &  x234 &  x254 &  x273 &  x274 &  x312 &  x320 &  x430 &  x434 &  x536 &  x605 &  x767 &  x799 &  x838 &  x877 &  x941 &  x944 &  x995 &  x1076 &  x1082 & ~x213 & ~x219 & ~x240 & ~x258 & ~x280 & ~x319 & ~x357 & ~x480;
assign c02 =  x83 &  x149 &  x152 &  x155 &  x161 &  x170 &  x173 &  x176 &  x185 &  x188 &  x206 &  x230 &  x263 &  x275 &  x284 &  x290 &  x305 &  x311 &  x338 &  x356 &  x370 &  x395 &  x407 &  x416 &  x428 &  x442 &  x481 &  x485 &  x521 &  x524 &  x551 &  x554 &  x563 &  x572 &  x587 &  x605 &  x611 &  x635 &  x650 &  x653 &  x668 &  x703 &  x704 &  x719 &  x737 &  x742 &  x758 &  x781 &  x791 &  x820 &  x830 &  x833 &  x854 &  x859 &  x881 &  x898 &  x932 &  x938 &  x968 &  x976 &  x979 &  x998 &  x1004 &  x1015 &  x1017 &  x1049 &  x1052 &  x1056 &  x1057 &  x1063 &  x1064 &  x1076 &  x1095 &  x1115 & ~x237 & ~x276 & ~x354 & ~x393 & ~x432 & ~x471 & ~x648;
assign c04 =  x14 &  x41 &  x44 &  x56 &  x110 &  x127 &  x131 &  x165 &  x204 &  x205 &  x224 &  x244 &  x254 &  x299 &  x335 &  x383 &  x394 &  x407 &  x410 &  x428 &  x433 &  x434 &  x472 &  x476 &  x494 &  x515 &  x518 &  x542 &  x551 &  x578 &  x605 &  x614 &  x616 &  x655 &  x793 &  x812 &  x818 &  x832 &  x838 &  x871 &  x877 &  x881 &  x899 &  x910 &  x917 &  x935 &  x955 &  x1031 &  x1052 &  x1079 &  x1118 & ~x702 & ~x741 & ~x780 & ~x819;
assign c06 =  x471 &  x539 &  x605 &  x836 &  x848 &  x851 &  x878 &  x926 &  x944 &  x1115 & ~x201 & ~x220 & ~x240;
assign c08 =  x55 &  x74 &  x94 &  x271 &  x299 &  x421 &  x463 &  x484 &  x530 &  x598 &  x632 &  x638 &  x640 &  x689 &  x757 & ~x1059 & ~x1098;
assign c010 =  x8 &  x29 &  x46 &  x85 &  x122 &  x124 &  x130 &  x140 &  x169 &  x170 &  x176 &  x239 &  x257 &  x308 &  x338 &  x341 &  x356 &  x401 &  x440 &  x443 &  x500 &  x503 &  x647 &  x832 &  x871 &  x875 &  x923 &  x1022 &  x1046 &  x1064 & ~x183 & ~x300 & ~x339 & ~x396 & ~x768;
assign c012 =  x5 &  x29 &  x131 &  x134 &  x137 &  x149 &  x155 &  x161 &  x173 &  x200 &  x260 &  x284 &  x287 &  x299 &  x320 &  x322 &  x338 &  x356 &  x365 &  x380 &  x410 &  x430 &  x449 &  x468 &  x469 &  x482 &  x500 &  x536 &  x547 &  x551 &  x557 &  x569 &  x586 &  x589 &  x590 &  x625 &  x638 &  x650 &  x664 &  x692 &  x703 &  x719 &  x724 &  x742 &  x749 &  x758 &  x802 &  x841 &  x860 &  x862 &  x878 &  x880 &  x941 &  x983 &  x1004 &  x1043 &  x1061 &  x1064 &  x1106 & ~x474;
assign c014 =  x161 &  x206 &  x275 &  x394 &  x433 &  x510 &  x549 &  x588 &  x883 &  x910 &  x1061 &  x1106 & ~x33 & ~x66 & ~x105 & ~x138 & ~x741;
assign c016 =  x2 &  x29 &  x155 &  x209 &  x272 &  x335 &  x338 &  x428 &  x467 &  x506 &  x507 &  x515 &  x546 &  x547 &  x572 &  x586 &  x625 &  x664 &  x695 &  x703 &  x742 &  x745 &  x776 &  x781 &  x791 &  x845 &  x854 &  x878 &  x887 &  x914 &  x935 &  x959 &  x971 &  x974 &  x995 &  x1004 &  x1016 &  x1028 &  x1043 &  x1072 &  x1073 &  x1082 &  x1103 & ~x276 & ~x474 & ~x513 & ~x552;
assign c018 =  x53 &  x80 &  x155 &  x170 &  x215 &  x245 &  x296 &  x356 &  x433 &  x542 &  x626 &  x628 &  x737 &  x836 &  x877 &  x905 &  x916 &  x1043 &  x1049 & ~x123 & ~x135 & ~x162 & ~x174 & ~x201 & ~x241 & ~x258 & ~x280 & ~x297;
assign c020 =  x2 &  x5 &  x11 &  x20 &  x32 &  x41 &  x50 &  x86 &  x92 &  x137 &  x146 &  x155 &  x185 &  x203 &  x242 &  x263 &  x266 &  x284 &  x305 &  x312 &  x316 &  x326 &  x350 &  x351 &  x352 &  x355 &  x365 &  x380 &  x392 &  x394 &  x398 &  x429 &  x430 &  x431 &  x433 &  x449 &  x452 &  x470 &  x472 &  x485 &  x503 &  x508 &  x511 &  x512 &  x515 &  x550 &  x557 &  x563 &  x569 &  x586 &  x587 &  x605 &  x611 &  x617 &  x628 &  x653 &  x665 &  x683 &  x707 &  x722 &  x731 &  x737 &  x755 &  x767 &  x782 &  x845 &  x854 &  x857 &  x881 &  x884 &  x893 &  x926 &  x938 &  x941 &  x959 &  x968 &  x983 &  x995 &  x1001 &  x1064 &  x1076 &  x1082 &  x1094 &  x1118 & ~x297 & ~x357 & ~x358 & ~x396;
assign c022 =  x104 &  x161 &  x182 &  x200 &  x206 &  x218 &  x254 &  x275 &  x386 &  x425 &  x464 &  x481 &  x503 &  x515 &  x551 &  x560 &  x586 &  x596 &  x611 &  x624 &  x626 &  x629 &  x644 &  x674 &  x680 &  x742 &  x770 &  x820 &  x830 &  x859 &  x881 &  x893 &  x898 &  x901 &  x937 &  x979 &  x995 &  x1010 &  x1015 &  x1052 &  x1054 &  x1093 &  x1121 & ~x432 & ~x510 & ~x708 & ~x709 & ~x747 & ~x786 & ~x825 & ~x831 & ~x864;
assign c024 =  x74 &  x107 &  x131 &  x149 &  x152 &  x173 &  x203 &  x206 &  x215 &  x275 &  x326 &  x395 &  x430 &  x468 &  x507 &  x508 &  x530 &  x536 &  x546 &  x547 &  x569 &  x586 &  x625 &  x644 &  x650 &  x664 &  x703 &  x704 &  x742 &  x767 &  x776 &  x830 &  x878 &  x902 &  x908 &  x956 &  x971 &  x1004 &  x1070 &  x1082 &  x1085 & ~x276 & ~x315 & ~x408 & ~x447 & ~x453 & ~x474 & ~x513 & ~x552 & ~x591 & ~x675;
assign c026 =  x68 &  x149 &  x185 &  x194 &  x200 &  x203 &  x209 &  x275 &  x338 &  x356 &  x386 &  x389 &  x395 &  x407 &  x437 &  x488 &  x497 &  x518 &  x559 &  x598 &  x601 &  x671 &  x680 &  x692 &  x797 &  x860 &  x863 &  x893 &  x902 &  x929 &  x940 &  x944 &  x975 &  x976 &  x979 &  x995 &  x1014 &  x1015 &  x1055 &  x1093 &  x1118 &  x1121 & ~x198 & ~x237 & ~x276 & ~x354 & ~x393 & ~x432 & ~x510 & ~x588 & ~x708 & ~x747 & ~x909;
assign c028 =  x29 &  x161 &  x221 &  x234 &  x273 &  x312 &  x430 &  x467 &  x686 &  x1010 & ~x201 & ~x219 & ~x258 & ~x259 & ~x297 & ~x516 & ~x555 & ~x819;
assign c030 =  x194 &  x284 &  x392 &  x547 &  x557 &  x586 &  x625 &  x626 &  x627 &  x664 &  x666 &  x737 &  x758 &  x783 &  x822 &  x861 &  x881 &  x1049 & ~x474 & ~x495 & ~x513 & ~x552;
assign c032 =  x11 &  x20 &  x95 &  x104 &  x113 &  x125 &  x134 &  x149 &  x206 &  x293 &  x317 &  x326 &  x353 &  x377 &  x425 &  x446 &  x461 &  x500 &  x503 &  x518 &  x527 &  x536 &  x546 &  x557 &  x566 &  x572 &  x586 &  x587 &  x625 &  x653 &  x664 &  x686 &  x692 &  x703 &  x719 &  x742 &  x746 &  x767 &  x782 &  x797 &  x818 &  x824 &  x827 &  x854 &  x857 &  x859 &  x881 &  x893 &  x959 &  x976 &  x983 &  x986 &  x1007 &  x1019 &  x1037 &  x1049 &  x1067 &  x1094 &  x1114 &  x1115 & ~x198 & ~x237 & ~x276 & ~x315 & ~x354 & ~x393 & ~x432 & ~x471 & ~x474 & ~x498 & ~x513 & ~x552 & ~x630;
assign c034 =  x128 &  x134 &  x137 &  x154 &  x155 &  x173 &  x193 &  x206 &  x209 &  x257 &  x287 &  x305 &  x386 &  x425 &  x455 &  x458 &  x461 &  x491 &  x497 &  x503 &  x644 &  x650 &  x677 &  x689 &  x745 &  x758 &  x764 &  x797 &  x822 &  x823 &  x861 &  x890 &  x900 &  x905 &  x926 &  x944 &  x947 &  x998 &  x1064 & ~x66 & ~x222 & ~x235 & ~x306 & ~x573;
assign c036 =  x125 &  x155 &  x170 &  x208 &  x356 &  x505 &  x605 &  x627 &  x666 &  x706 &  x823 &  x844 &  x854 &  x883 &  x921 &  x922 &  x960 &  x1049 &  x1112;
assign c038 =  x11 &  x149 &  x161 &  x173 &  x282 &  x283 &  x322 &  x347 &  x355 &  x433 &  x434 &  x440 &  x550 &  x608 &  x881 &  x884 &  x910 &  x959 &  x1022 & ~x396 & ~x516 & ~x555;
assign c040 =  x5 &  x14 &  x49 &  x55 &  x68 &  x88 &  x94 &  x127 &  x131 &  x146 &  x165 &  x166 &  x173 &  x182 &  x205 &  x215 &  x251 &  x263 &  x275 &  x287 &  x293 &  x302 &  x335 &  x338 &  x347 &  x356 &  x389 &  x398 &  x419 &  x433 &  x446 &  x449 &  x461 &  x497 &  x511 &  x524 &  x527 &  x533 &  x557 &  x605 &  x611 &  x632 &  x644 &  x665 &  x689 &  x694 &  x716 &  x737 &  x749 &  x821 &  x830 &  x833 &  x874 &  x875 &  x881 &  x887 &  x905 &  x908 &  x962 &  x995 &  x1004 &  x1037 &  x1046 &  x1052 &  x1058 &  x1073 &  x1109 & ~x219;
assign c042 =  x8 &  x44 &  x62 &  x74 &  x104 &  x116 &  x125 &  x131 &  x154 &  x155 &  x179 &  x182 &  x192 &  x193 &  x206 &  x221 &  x231 &  x232 &  x254 &  x270 &  x271 &  x281 &  x314 &  x317 &  x326 &  x353 &  x362 &  x377 &  x380 &  x383 &  x398 &  x422 &  x428 &  x431 &  x446 &  x473 &  x497 &  x506 &  x509 &  x515 &  x521 &  x527 &  x530 &  x539 &  x581 &  x602 &  x620 &  x638 &  x701 &  x743 &  x776 &  x782 &  x800 &  x824 &  x827 &  x845 &  x872 &  x878 &  x890 &  x901 &  x902 &  x923 &  x968 &  x979 &  x995 &  x1010 &  x1025 &  x1052 &  x1058 &  x1064 &  x1070 &  x1073 &  x1082 &  x1100 &  x1112 &  x1118 & ~x534 & ~x969 & ~x1041;
assign c044 =  x11 &  x23 &  x44 &  x56 &  x95 &  x104 &  x122 &  x128 &  x152 &  x185 &  x212 &  x215 &  x236 &  x247 &  x263 &  x272 &  x286 &  x302 &  x325 &  x338 &  x356 &  x364 &  x380 &  x404 &  x407 &  x422 &  x428 &  x455 &  x461 &  x473 &  x497 &  x533 &  x545 &  x551 &  x569 &  x581 &  x587 &  x611 &  x614 &  x644 &  x653 &  x662 &  x680 &  x683 &  x689 &  x704 &  x737 &  x749 &  x773 &  x824 &  x832 &  x845 &  x854 &  x872 &  x875 &  x878 &  x905 &  x916 &  x932 &  x935 &  x955 &  x959 &  x994 &  x1028 &  x1037 &  x1046 &  x1082 & ~x252 & ~x369 & ~x408 & ~x474 & ~x513;
assign c046 =  x2 &  x20 &  x23 &  x38 &  x50 &  x74 &  x131 &  x140 &  x143 &  x149 &  x164 &  x200 &  x203 &  x221 &  x233 &  x236 &  x251 &  x263 &  x269 &  x272 &  x284 &  x287 &  x293 &  x320 &  x323 &  x332 &  x338 &  x350 &  x362 &  x368 &  x416 &  x419 &  x422 &  x473 &  x485 &  x500 &  x518 &  x521 &  x533 &  x551 &  x587 &  x590 &  x596 &  x611 &  x625 &  x629 &  x638 &  x644 &  x647 &  x664 &  x698 &  x701 &  x719 &  x722 &  x731 &  x734 &  x740 &  x742 &  x755 &  x758 &  x767 &  x773 &  x781 &  x809 &  x820 &  x830 &  x848 &  x859 &  x875 &  x890 &  x898 &  x899 &  x901 &  x937 &  x938 &  x941 &  x944 &  x950 &  x971 &  x976 &  x979 &  x995 &  x1010 &  x1015 &  x1018 &  x1019 &  x1049 &  x1052 &  x1054 &  x1057 &  x1070 &  x1076 &  x1127 & ~x315 & ~x354 & ~x393 & ~x432 & ~x471 & ~x549 & ~x630 & ~x669 & ~x670 & ~x708 & ~x709 & ~x747 & ~x748 & ~x786 & ~x787 & ~x825 & ~x831 & ~x864 & ~x870;
assign c048 =  x55 &  x541 & ~x96 & ~x102 & ~x123 & ~x162 & ~x213 & ~x216 & ~x240 & ~x255;
assign c050 =  x77 &  x86 &  x101 &  x149 &  x155 &  x170 &  x227 &  x236 &  x284 &  x356 &  x383 &  x386 &  x471 &  x479 &  x494 &  x500 &  x510 &  x512 &  x549 &  x588 &  x590 &  x605 &  x608 &  x611 &  x620 &  x627 &  x628 &  x644 &  x683 &  x692 &  x707 &  x716 &  x755 &  x767 &  x803 &  x823 &  x845 &  x869 &  x883 &  x908 &  x935 &  x1013 &  x1025 &  x1094 & ~x27 & ~x33 & ~x300 & ~x339 & ~x378 & ~x417 & ~x456 & ~x495;
assign c052 =  x98 &  x113 &  x236 &  x239 &  x251 &  x254 &  x311 &  x329 &  x356 &  x388 &  x392 &  x433 &  x434 &  x446 &  x503 &  x530 &  x554 &  x605 &  x611 &  x632 &  x644 &  x689 &  x695 &  x704 &  x844 &  x854 &  x881 &  x883 &  x922 &  x941 &  x965 &  x995 &  x1028 &  x1049 & ~x774 & ~x775 & ~x813 & ~x1041 & ~x1080;
assign c054 =  x155 &  x260 &  x416 &  x430 &  x551 &  x574 &  x586 &  x587 &  x613 &  x625 &  x652 &  x656 &  x664 &  x703 &  x742 &  x776 &  x788 &  x794 &  x881 &  x944 &  x955 &  x959 &  x994 &  x1064 &  x1072 & ~x297 & ~x1020;
assign c056 =  x56 &  x80 &  x104 &  x110 &  x143 &  x185 &  x218 &  x236 &  x242 &  x254 &  x299 &  x317 &  x329 &  x404 &  x410 &  x416 &  x419 &  x433 &  x437 &  x602 &  x611 &  x617 &  x623 &  x641 &  x644 &  x683 &  x689 &  x701 &  x746 &  x752 &  x782 &  x805 &  x844 &  x854 &  x862 &  x881 &  x883 &  x914 &  x922 &  x923 &  x947 &  x968 &  x974 &  x1000 & ~x33 & ~x72 & ~x339 & ~x378 & ~x417 & ~x456 & ~x1002 & ~x1041 & ~x1080 & ~x1119;
assign c058 =  x5 &  x20 &  x35 &  x59 &  x77 &  x86 &  x104 &  x119 &  x149 &  x155 &  x170 &  x176 &  x206 &  x209 &  x215 &  x233 &  x251 &  x260 &  x266 &  x275 &  x287 &  x299 &  x302 &  x305 &  x308 &  x311 &  x317 &  x332 &  x356 &  x365 &  x380 &  x407 &  x455 &  x461 &  x470 &  x488 &  x518 &  x521 &  x527 &  x533 &  x547 &  x560 &  x586 &  x589 &  x620 &  x629 &  x641 &  x644 &  x647 &  x653 &  x656 &  x701 &  x758 &  x776 &  x779 &  x783 &  x794 &  x812 &  x823 &  x854 &  x860 &  x862 &  x863 &  x869 &  x884 &  x896 &  x899 &  x901 &  x920 &  x929 &  x935 &  x940 &  x941 &  x944 &  x947 &  x953 &  x956 &  x968 &  x998 &  x1004 &  x1022 &  x1049 &  x1076 &  x1082 &  x1124 & ~x222 & ~x294 & ~x339 & ~x378 & ~x513 & ~x1041 & ~x1053 & ~x1080 & ~x1119;
assign c060 =  x161 &  x182 &  x266 &  x290 &  x323 &  x338 &  x512 &  x605 &  x641 &  x689 &  x815 &  x821 &  x884 &  x919 &  x979 &  x983 &  x997 &  x1022 &  x1064 &  x1069 &  x1109 &  x1127 & ~x6 & ~x45 & ~x84 & ~x1080;
assign c062 =  x26 &  x62 &  x131 &  x143 &  x263 &  x305 &  x320 &  x344 &  x356 &  x430 &  x468 &  x469 &  x497 &  x500 &  x508 &  x509 &  x542 &  x547 &  x551 &  x586 &  x605 &  x625 &  x638 &  x655 &  x664 &  x683 &  x698 &  x703 &  x719 &  x742 &  x745 &  x749 &  x773 &  x820 &  x824 &  x836 &  x851 &  x914 &  x968 &  x979 &  x983 &  x1013 &  x1018 &  x1055 &  x1115 & ~x435 & ~x474 & ~x513 & ~x552 & ~x636;
assign c064 =  x17 &  x32 &  x68 &  x74 &  x83 &  x86 &  x104 &  x119 &  x149 &  x161 &  x167 &  x221 &  x235 &  x251 &  x273 &  x274 &  x277 &  x293 &  x308 &  x329 &  x354 &  x365 &  x391 &  x393 &  x398 &  x407 &  x410 &  x416 &  x432 &  x433 &  x449 &  x471 &  x473 &  x510 &  x527 &  x590 &  x632 &  x689 &  x695 &  x707 &  x713 &  x719 &  x743 &  x752 &  x758 &  x760 &  x767 &  x770 &  x773 &  x794 &  x799 &  x800 &  x806 &  x830 &  x838 &  x857 &  x877 &  x893 &  x905 &  x917 &  x920 &  x929 &  x938 &  x944 &  x992 &  x1010 &  x1052 &  x1079 &  x1082 &  x1091 &  x1106 &  x1118 &  x1130 & ~x780;
assign c066 =  x1 &  x67 &  x73 &  x106 &  x112 &  x118 &  x134 &  x278 &  x328 &  x502 &  x625 &  x664 &  x703 &  x730 &  x781 &  x808 &  x859 &  x880 &  x918 &  x919 &  x925 &  x979 &  x1015 &  x1018 &  x1057;
assign c068 =  x35 &  x65 &  x68 &  x104 &  x107 &  x119 &  x125 &  x137 &  x143 &  x155 &  x161 &  x185 &  x200 &  x215 &  x233 &  x251 &  x254 &  x272 &  x284 &  x287 &  x290 &  x299 &  x350 &  x356 &  x359 &  x365 &  x368 &  x380 &  x383 &  x398 &  x413 &  x416 &  x430 &  x431 &  x443 &  x458 &  x468 &  x470 &  x485 &  x507 &  x508 &  x512 &  x521 &  x536 &  x547 &  x554 &  x569 &  x575 &  x586 &  x587 &  x602 &  x611 &  x614 &  x625 &  x647 &  x659 &  x664 &  x668 &  x680 &  x692 &  x698 &  x703 &  x710 &  x719 &  x725 &  x740 &  x742 &  x749 &  x758 &  x770 &  x781 &  x782 &  x818 &  x823 &  x833 &  x857 &  x862 &  x878 &  x905 &  x923 &  x941 &  x956 &  x971 &  x1004 &  x1007 &  x1013 &  x1061 &  x1076 &  x1082 &  x1088 &  x1124 &  x1130 & ~x474 & ~x513 & ~x552 & ~x591 & ~x675 & ~x1119;
assign c070 =  x101 &  x155 &  x203 &  x212 &  x220 &  x236 &  x245 &  x287 &  x299 &  x332 &  x365 &  x407 &  x422 &  x428 &  x449 &  x452 &  x554 &  x569 &  x653 &  x664 &  x665 &  x671 &  x674 &  x689 &  x703 &  x719 &  x728 &  x742 &  x779 &  x782 &  x788 &  x859 &  x861 &  x863 &  x872 &  x890 &  x898 &  x900 &  x932 &  x938 &  x939 &  x950 &  x976 &  x978 &  x979 &  x1004 &  x1010 &  x1015 &  x1017 &  x1056 &  x1057 &  x1058 &  x1082 &  x1103 & ~x312 & ~x354 & ~x393 & ~x495 & ~x648;
assign c072 =  x80 &  x472 &  x592 &  x629 &  x640 &  x671 &  x761 &  x944 &  x956 &  x1052 &  x1070 &  x1130 & ~x99 & ~x123 & ~x138 & ~x162 & ~x168 & ~x177 & ~x201 & ~x216 & ~x240;
assign c074 =  x44 &  x89 &  x125 &  x140 &  x146 &  x176 &  x266 &  x323 &  x360 &  x405 &  x458 &  x506 &  x566 &  x586 &  x625 &  x629 &  x664 &  x668 &  x671 &  x764 &  x845 &  x863 &  x880 &  x938 &  x956 &  x962 &  x977 &  x1106 &  x1112;
assign c076 =  x8 &  x11 &  x26 &  x32 &  x59 &  x74 &  x83 &  x101 &  x107 &  x116 &  x131 &  x134 &  x137 &  x176 &  x182 &  x188 &  x206 &  x215 &  x239 &  x242 &  x257 &  x260 &  x275 &  x287 &  x311 &  x320 &  x323 &  x326 &  x338 &  x344 &  x356 &  x392 &  x401 &  x419 &  x437 &  x449 &  x470 &  x497 &  x515 &  x554 &  x563 &  x569 &  x584 &  x586 &  x602 &  x605 &  x611 &  x617 &  x629 &  x638 &  x641 &  x644 &  x650 &  x653 &  x664 &  x689 &  x698 &  x703 &  x704 &  x706 &  x713 &  x716 &  x719 &  x725 &  x731 &  x737 &  x740 &  x742 &  x745 &  x755 &  x767 &  x773 &  x782 &  x783 &  x785 &  x809 &  x812 &  x815 &  x818 &  x820 &  x822 &  x823 &  x833 &  x836 &  x845 &  x859 &  x861 &  x862 &  x881 &  x884 &  x893 &  x896 &  x898 &  x900 &  x917 &  x926 &  x939 &  x941 &  x944 &  x956 &  x959 &  x976 &  x979 &  x1010 &  x1018 &  x1034 &  x1037 &  x1049 &  x1057 &  x1061 &  x1066 &  x1073 &  x1100 &  x1114 &  x1130;
assign c078 =  x8 &  x38 &  x74 &  x83 &  x86 &  x101 &  x104 &  x116 &  x125 &  x128 &  x131 &  x134 &  x140 &  x146 &  x152 &  x155 &  x161 &  x164 &  x173 &  x185 &  x200 &  x242 &  x266 &  x275 &  x284 &  x293 &  x299 &  x305 &  x323 &  x338 &  x350 &  x356 &  x380 &  x386 &  x392 &  x401 &  x404 &  x410 &  x419 &  x425 &  x428 &  x434 &  x443 &  x446 &  x449 &  x470 &  x479 &  x497 &  x500 &  x512 &  x518 &  x536 &  x548 &  x551 &  x557 &  x562 &  x569 &  x601 &  x611 &  x626 &  x644 &  x647 &  x650 &  x664 &  x665 &  x671 &  x674 &  x686 &  x701 &  x702 &  x703 &  x704 &  x707 &  x719 &  x728 &  x731 &  x740 &  x742 &  x758 &  x767 &  x773 &  x781 &  x785 &  x794 &  x812 &  x815 &  x820 &  x830 &  x833 &  x854 &  x859 &  x862 &  x898 &  x899 &  x900 &  x902 &  x914 &  x920 &  x932 &  x937 &  x939 &  x940 &  x950 &  x956 &  x962 &  x965 &  x968 &  x976 &  x978 &  x979 &  x980 &  x995 &  x1007 &  x1010 &  x1015 &  x1017 &  x1018 &  x1034 &  x1043 &  x1049 &  x1054 &  x1056 &  x1057 &  x1082 &  x1088 &  x1093 &  x1095 &  x1109 &  x1112 &  x1130 & ~x669 & ~x708 & ~x831;
assign c080 =  x5 &  x29 &  x74 &  x161 &  x164 &  x179 &  x215 &  x221 &  x251 &  x254 &  x263 &  x320 &  x347 &  x356 &  x392 &  x410 &  x425 &  x430 &  x437 &  x469 &  x485 &  x503 &  x530 &  x550 &  x554 &  x557 &  x569 &  x587 &  x590 &  x616 &  x626 &  x647 &  x686 &  x698 &  x737 &  x770 &  x824 &  x854 &  x860 &  x881 &  x896 &  x902 &  x914 &  x929 &  x941 &  x944 &  x968 &  x1055 &  x1082 &  x1115 & ~x135 & ~x294 & ~x396 & ~x855 & ~x933 & ~x972;
assign c082 =  x62 &  x65 &  x80 &  x156 &  x299 &  x338 &  x378 &  x593 &  x599 & ~x142 & ~x180 & ~x201 & ~x219 & ~x258;
assign c084 =  x117 &  x156 &  x173 &  x182 &  x195 &  x196 &  x215 &  x234 &  x269 &  x316 &  x433 &  x721 &  x737 &  x776 &  x799 &  x908 &  x1061 &  x1066 & ~x141 & ~x142 & ~x180 & ~x220 & ~x258;
assign c086 =  x2 &  x17 &  x47 &  x68 &  x98 &  x101 &  x110 &  x122 &  x131 &  x234 &  x235 &  x242 &  x251 &  x305 &  x335 &  x362 &  x368 &  x374 &  x472 &  x518 &  x602 &  x611 &  x635 &  x659 &  x692 &  x701 &  x746 &  x758 &  x761 &  x782 &  x794 &  x812 &  x818 &  x833 &  x857 &  x881 &  x902 &  x908 &  x986 &  x989 &  x1004 &  x1016 &  x1040 &  x1076 &  x1094 & ~x201 & ~x213 & ~x219 & ~x220 & ~x252 & ~x258 & ~x259 & ~x291 & ~x298 & ~x819;
assign c088 =  x79 &  x82 &  x117 &  x156 &  x179 &  x196 &  x206 &  x234 &  x317 &  x355 &  x371 &  x394 &  x433 &  x461 &  x518 &  x548 &  x598 &  x689 &  x719 &  x721 &  x799 &  x838 &  x877 &  x1004 & ~x141 & ~x142 & ~x180 & ~x219 & ~x258 & ~x324 & ~x819;
assign c090 =  x284 &  x374 &  x433 &  x472 &  x539 &  x638 &  x727 &  x758 &  x805 &  x832 &  x904 &  x926 &  x943 &  x982 &  x1021 & ~x138 & ~x702 & ~x852 & ~x930 & ~x969 & ~x1047;
assign c092 =  x8 &  x29 &  x41 &  x44 &  x47 &  x50 &  x56 &  x74 &  x77 &  x80 &  x86 &  x92 &  x95 &  x104 &  x119 &  x128 &  x131 &  x140 &  x146 &  x149 &  x155 &  x158 &  x170 &  x173 &  x182 &  x191 &  x194 &  x206 &  x221 &  x224 &  x230 &  x251 &  x254 &  x260 &  x263 &  x266 &  x275 &  x281 &  x284 &  x287 &  x293 &  x299 &  x305 &  x308 &  x320 &  x329 &  x332 &  x338 &  x341 &  x347 &  x356 &  x365 &  x368 &  x374 &  x377 &  x380 &  x392 &  x395 &  x425 &  x428 &  x437 &  x440 &  x443 &  x452 &  x455 &  x467 &  x482 &  x500 &  x503 &  x512 &  x515 &  x518 &  x530 &  x539 &  x545 &  x560 &  x590 &  x593 &  x611 &  x620 &  x625 &  x647 &  x650 &  x653 &  x664 &  x668 &  x671 &  x677 &  x683 &  x695 &  x703 &  x704 &  x710 &  x716 &  x731 &  x734 &  x737 &  x742 &  x743 &  x745 &  x758 &  x761 &  x767 &  x770 &  x773 &  x776 &  x785 &  x788 &  x794 &  x803 &  x806 &  x830 &  x833 &  x842 &  x857 &  x859 &  x860 &  x866 &  x869 &  x872 &  x881 &  x886 &  x890 &  x893 &  x898 &  x902 &  x911 &  x935 &  x937 &  x938 &  x939 &  x940 &  x941 &  x944 &  x956 &  x959 &  x965 &  x968 &  x976 &  x978 &  x979 &  x983 &  x995 &  x1007 &  x1015 &  x1017 &  x1018 &  x1025 &  x1031 &  x1034 &  x1043 &  x1049 &  x1055 &  x1057 &  x1061 &  x1070 &  x1076 &  x1085 &  x1088 &  x1094 &  x1096 &  x1106 &  x1109 &  x1115 &  x1130 & ~x474 & ~x513;
assign c094 =  x49 &  x157 &  x195 &  x238 &  x355 &  x421 &  x433 &  x605 &  x640 &  x739 &  x968 &  x1127 & ~x546;
assign c096 =  x8 &  x26 &  x86 &  x89 &  x98 &  x218 &  x263 &  x278 &  x317 &  x359 &  x742 &  x784 &  x851 &  x859 &  x861 &  x881 &  x898 &  x902 &  x939 &  x976 &  x978 &  x979 &  x1015 &  x1017 &  x1018 &  x1025 &  x1054 &  x1056 &  x1057 &  x1095 & ~x15 & ~x54 & ~x249 & ~x327;
assign c098 =  x17 &  x55 &  x134 &  x248 &  x281 &  x574 &  x640 &  x647 &  x719 &  x857 &  x877 &  x886 &  x924 &  x925 &  x964 &  x1063 &  x1087 &  x1102 & ~x6;
assign c0100 =  x5 &  x38 &  x164 &  x206 &  x275 &  x344 &  x497 &  x627 &  x628 &  x680 &  x682 &  x689 &  x798 &  x823 &  x838 &  x860 &  x877 &  x914 &  x916 &  x998 &  x1021 &  x1060;
assign c0102 =  x275 &  x445 &  x518 &  x769 &  x808 &  x859 &  x885 &  x886 &  x979 &  x1057 & ~x120 & ~x198 & ~x237 & ~x276 & ~x354;
assign c0104 =  x23 &  x71 &  x119 &  x137 &  x164 &  x251 &  x296 &  x299 &  x308 &  x319 &  x329 &  x488 &  x494 &  x515 &  x536 &  x547 &  x586 &  x625 &  x664 &  x674 &  x677 &  x725 &  x734 &  x742 &  x770 &  x820 &  x821 &  x859 &  x866 &  x872 &  x878 &  x884 &  x898 &  x944 &  x956 &  x979 &  x1015 &  x1018 &  x1022 &  x1057 &  x1061 &  x1093 &  x1096 &  x1112 & ~x354 & ~x393 & ~x432 & ~x513 & ~x552 & ~x567 & ~x591;
assign c0106 =  x73 &  x79 &  x92 &  x110 &  x146 &  x151 &  x167 &  x178 &  x217 &  x322 &  x338 &  x339 &  x340 &  x377 &  x419 &  x442 &  x502 &  x518 &  x524 &  x541 &  x551 &  x562 &  x574 &  x704 &  x734 &  x806 &  x919 &  x956 &  x976 &  x1025 &  x1048 &  x1052 &  x1057;
assign c0108 =  x11 &  x53 &  x80 &  x86 &  x89 &  x125 &  x134 &  x158 &  x170 &  x206 &  x224 &  x227 &  x233 &  x281 &  x284 &  x299 &  x344 &  x359 &  x368 &  x374 &  x416 &  x422 &  x440 &  x458 &  x476 &  x482 &  x512 &  x520 &  x559 &  x563 &  x569 &  x608 &  x629 &  x683 &  x686 &  x698 &  x701 &  x722 &  x776 &  x812 &  x854 &  x859 &  x893 &  x897 &  x898 &  x905 &  x911 &  x936 &  x940 &  x959 &  x975 &  x976 &  x979 &  x989 &  x1014 &  x1053 &  x1057 &  x1064 &  x1070 &  x1091 &  x1092 &  x1093 & ~x471 & ~x510 & ~x708 & ~x747 & ~x786 & ~x972;
assign c0110 =  x32 &  x215 &  x338 &  x368 &  x500 &  x586 &  x625 &  x626 &  x664 &  x703 &  x742 &  x764 &  x845 &  x859 &  x866 &  x898 &  x979 &  x1018 &  x1055 &  x1057 &  x1064 &  x1103 & ~x354 & ~x474 & ~x513 & ~x528 & ~x552 & ~x567 & ~x631 & ~x708 & ~x747;
assign c0112 =  x37 &  x91 &  x170 &  x521 &  x589 &  x716 &  x785 &  x800 &  x805 &  x811 &  x818 &  x832 &  x844 &  x871 &  x883 &  x910 &  x922 &  x961 &  x983 &  x1039 & ~x294 & ~x333;
assign c0114 =  x71 &  x78 &  x104 &  x117 &  x156 &  x194 &  x196 &  x218 &  x221 &  x234 &  x274 &  x320 &  x394 &  x433 &  x446 &  x530 &  x539 &  x650 &  x656 &  x659 &  x677 &  x716 &  x734 &  x760 &  x812 &  x839 &  x845 &  x872 &  x890 &  x902 &  x959 &  x968 &  x1022 &  x1073 &  x1112 & ~x102 & ~x135 & ~x141 & ~x142 & ~x162 & ~x180 & ~x181 & ~x201 & ~x258 & ~x297;
assign c0116 =  x203 &  x274 &  x299 &  x359 &  x374 &  x418 &  x425 &  x473 &  x541 &  x557 &  x559 &  x578 &  x584 &  x598 &  x635 &  x656 &  x662 &  x697 &  x698 &  x701 &  x757 &  x808 &  x836 &  x995 &  x1010 & ~x84 & ~x123 & ~x162 & ~x201 & ~x708 & ~x1059;
assign c0118 =  x65 &  x77 &  x92 &  x116 &  x152 &  x161 &  x239 &  x266 &  x305 &  x323 &  x386 &  x392 &  x398 &  x419 &  x446 &  x455 &  x485 &  x497 &  x500 &  x507 &  x508 &  x530 &  x546 &  x547 &  x585 &  x586 &  x608 &  x624 &  x625 &  x664 &  x671 &  x703 &  x730 &  x737 &  x742 &  x788 &  x797 &  x809 &  x836 &  x898 &  x899 &  x920 &  x932 &  x940 &  x941 &  x979 &  x986 &  x1001 &  x1007 &  x1013 &  x1022 &  x1028 &  x1034 &  x1091 &  x1118 &  x1121 & ~x474 & ~x513 & ~x552 & ~x591 & ~x672 & ~x675;
assign c0120 =  x77 &  x98 &  x104 &  x125 &  x203 &  x206 &  x272 &  x314 &  x332 &  x359 &  x362 &  x374 &  x464 &  x518 &  x530 &  x536 &  x569 &  x587 &  x593 &  x644 &  x650 &  x683 &  x704 &  x800 &  x803 &  x809 &  x833 &  x881 &  x896 &  x914 &  x929 &  x950 &  x986 &  x995 &  x1027 &  x1030 &  x1031 &  x1061 &  x1066 &  x1091 &  x1127 & ~x6 & ~x45 & ~x84 & ~x123 & ~x162 & ~x201 & ~x207 & ~x249 & ~x288;
assign c0122 =  x209 &  x440 &  x725 &  x822 &  x968 &  x979 &  x1052 &  x1130 & ~x33 & ~x177 & ~x216 & ~x294 & ~x300 & ~x339 & ~x474 & ~x489 & ~x495 & ~x1041;
assign c0124 =  x5 &  x43 &  x47 &  x62 &  x65 &  x68 &  x79 &  x80 &  x82 &  x98 &  x117 &  x137 &  x140 &  x149 &  x157 &  x160 &  x176 &  x182 &  x188 &  x194 &  x209 &  x233 &  x236 &  x245 &  x260 &  x316 &  x344 &  x355 &  x380 &  x393 &  x394 &  x395 &  x401 &  x421 &  x422 &  x443 &  x479 &  x530 &  x575 &  x587 &  x605 &  x626 &  x644 &  x659 &  x668 &  x677 &  x683 &  x701 &  x721 &  x725 &  x739 &  x752 &  x758 &  x779 &  x799 &  x818 &  x881 &  x896 &  x916 &  x938 &  x956 &  x977 &  x1034 &  x1064 &  x1121 &  x1130 & ~x546;
assign c0126 =  x8 &  x35 &  x59 &  x89 &  x92 &  x131 &  x134 &  x149 &  x152 &  x161 &  x176 &  x182 &  x188 &  x215 &  x224 &  x227 &  x233 &  x254 &  x260 &  x266 &  x272 &  x275 &  x293 &  x299 &  x326 &  x353 &  x374 &  x386 &  x392 &  x407 &  x425 &  x428 &  x440 &  x449 &  x469 &  x497 &  x507 &  x508 &  x527 &  x536 &  x546 &  x547 &  x551 &  x566 &  x585 &  x586 &  x587 &  x620 &  x624 &  x625 &  x629 &  x638 &  x653 &  x656 &  x662 &  x664 &  x674 &  x698 &  x703 &  x710 &  x713 &  x742 &  x745 &  x749 &  x764 &  x776 &  x781 &  x782 &  x794 &  x830 &  x854 &  x862 &  x878 &  x881 &  x938 &  x944 &  x998 &  x1010 &  x1028 &  x1043 &  x1076 &  x1106 & ~x447 & ~x453 & ~x474 & ~x513 & ~x552 & ~x591 & ~x708 & ~x747;
assign c0128 =  x182 &  x341 &  x428 &  x443 &  x445 &  x482 &  x485 &  x518 &  x520 &  x536 &  x559 &  x605 &  x611 &  x689 &  x710 &  x764 &  x769 &  x808 &  x956 &  x959 &  x1004 &  x1019 &  x1064 &  x1076 &  x1100 & ~x6 & ~x45 & ~x84 & ~x123 & ~x201 & ~x606 & ~x1083;
assign c0130 =  x56 &  x164 &  x170 &  x182 &  x185 &  x274 &  x316 &  x338 &  x356 &  x394 &  x452 &  x482 &  x566 &  x577 &  x656 &  x659 &  x694 &  x718 &  x728 &  x733 &  x778 &  x796 &  x798 &  x821 &  x838 &  x850 &  x851 &  x863 &  x876 &  x881 &  x889 &  x941 &  x947 &  x953 &  x955 &  x968 &  x995 &  x1006 &  x1027 &  x1043 &  x1049 &  x1066 & ~x702 & ~x741 & ~x780;
assign c0132 =  x52 &  x155 & ~x69 & ~x177 & ~x216 & ~x222 & ~x294 & ~x969 & ~x1002 & ~x1041;
assign c0134 =  x35 &  x89 &  x125 &  x149 &  x188 &  x206 &  x212 &  x227 &  x251 &  x266 &  x329 &  x338 &  x374 &  x419 &  x434 &  x443 &  x461 &  x482 &  x521 &  x524 &  x533 &  x547 &  x572 &  x581 &  x586 &  x617 &  x625 &  x650 &  x664 &  x703 &  x719 &  x731 &  x742 &  x770 &  x820 &  x824 &  x857 &  x859 &  x884 &  x898 &  x937 &  x940 &  x976 &  x979 &  x1010 &  x1016 &  x1031 &  x1040 & ~x474 & ~x487 & ~x513 & ~x552 & ~x591 & ~x630;
assign c0136 =  x17 &  x41 &  x74 &  x149 &  x182 &  x206 &  x215 &  x274 &  x275 &  x312 &  x352 &  x394 &  x433 &  x455 &  x469 &  x508 &  x511 &  x518 &  x547 &  x566 &  x569 &  x586 &  x596 &  x623 &  x692 &  x719 &  x838 &  x848 &  x854 &  x877 &  x916 &  x929 &  x955 &  x956 &  x968 &  x994 &  x1004 &  x1061 &  x1073 &  x1082 & ~x702 & ~x819;
assign c0138 =  x5 &  x23 &  x53 &  x59 &  x149 &  x152 &  x155 &  x161 &  x188 &  x206 &  x209 &  x251 &  x284 &  x380 &  x485 &  x488 &  x491 &  x509 &  x515 &  x518 &  x554 &  x560 &  x608 &  x611 &  x644 &  x671 &  x698 &  x705 &  x719 &  x737 &  x744 &  x746 &  x758 &  x783 &  x821 &  x823 &  x860 &  x877 &  x878 &  x908 &  x914 &  x915 &  x923 &  x941 &  x954 &  x955 &  x993 &  x994 &  x995 &  x1052 &  x1064 &  x1072;
assign c0140 =  x5 &  x149 &  x182 &  x299 &  x356 &  x430 &  x1073 & ~x138 & ~x177 & ~x216 & ~x436 & ~x475 & ~x480 & ~x513 & ~x555;
assign c0142 =  x74 &  x89 &  x131 &  x191 &  x245 &  x350 &  x425 &  x452 &  x548 &  x560 &  x664 &  x745 &  x746 &  x776 &  x785 &  x845 &  x848 &  x854 &  x859 &  x860 &  x861 &  x869 &  x893 &  x898 &  x902 &  x908 &  x939 &  x959 &  x968 &  x979 &  x986 &  x1015 &  x1037 &  x1056 &  x1057 &  x1070 &  x1094 & ~x642 & ~x643 & ~x708;
assign c0144 =  x28 &  x38 &  x55 &  x66 &  x105 &  x106 &  x107 &  x143 &  x144 &  x151 &  x182 &  x190 &  x230 &  x338 &  x386 &  x580 &  x586 &  x619 &  x659 &  x664 &  x820 &  x898 &  x959 &  x1015 &  x1048 &  x1093 & ~x237 & ~x276 & ~x354 & ~x393 & ~x471;
assign c0146 =  x38 &  x53 &  x74 &  x86 &  x176 &  x191 &  x197 &  x209 &  x221 &  x254 &  x263 &  x274 &  x290 &  x296 &  x302 &  x323 &  x371 &  x394 &  x430 &  x433 &  x455 &  x467 &  x472 &  x512 &  x539 &  x569 &  x581 &  x650 &  x668 &  x674 &  x689 &  x695 &  x701 &  x704 &  x731 &  x755 &  x770 &  x773 &  x794 &  x827 &  x851 &  x854 &  x878 &  x926 &  x941 &  x944 &  x1001 &  x1019 &  x1028 &  x1031 &  x1055 &  x1070 &  x1073 &  x1130 & ~x138 & ~x177 & ~x180 & ~x819 & ~x858 & ~x1020 & ~x1059 & ~x1098;
assign c0148 =  x43 &  x131 &  x224 &  x431 &  x505 &  x560 &  x592 &  x632 &  x637 &  x728 &  x748 &  x838 &  x992 &  x1031 &  x1064 & ~x63 & ~x102 & ~x141 & ~x210 & ~x249;
assign c0150 =  x73 &  x112 &  x265 &  x523 &  x559 &  x858 &  x897 &  x898 &  x936 &  x975 &  x1014 &  x1052 &  x1092 &  x1093 & ~x12 & ~x276 & ~x708;
assign c0152 =  x74 &  x89 &  x110 &  x117 &  x125 &  x155 &  x156 &  x157 &  x164 &  x182 &  x195 &  x203 &  x234 &  x266 &  x275 &  x281 &  x311 &  x350 &  x356 &  x380 &  x389 &  x392 &  x394 &  x407 &  x410 &  x433 &  x440 &  x472 &  x473 &  x500 &  x518 &  x526 &  x563 &  x566 &  x575 &  x584 &  x611 &  x640 &  x642 &  x650 &  x668 &  x681 &  x695 &  x709 &  x713 &  x737 &  x746 &  x748 &  x758 &  x779 &  x782 &  x791 &  x809 &  x812 &  x836 &  x851 &  x860 &  x875 &  x878 &  x890 &  x917 &  x944 &  x998 &  x1004 &  x1007 &  x1016 &  x1019 &  x1025 &  x1049;
assign c0154 =  x149 &  x182 &  x230 &  x247 &  x305 &  x325 &  x547 &  x586 &  x587 &  x625 &  x627 &  x628 &  x638 &  x668 &  x698 &  x703 &  x704 &  x719 &  x822 &  x861 &  x939 &  x944 &  x962 &  x1004 &  x1019 &  x1055 &  x1103 & ~x552;
assign c0156 =  x74 &  x89 &  x104 &  x131 &  x215 &  x232 &  x278 &  x293 &  x323 &  x326 &  x329 &  x359 &  x440 &  x503 &  x511 &  x560 &  x563 &  x590 &  x608 &  x629 &  x638 &  x680 &  x725 &  x772 &  x810 &  x812 &  x817 &  x821 &  x871 &  x884 &  x902 &  x1010 &  x1026 &  x1042 &  x1049 &  x1124;
assign c0158 =  x176 &  x196 &  x230 &  x234 &  x254 &  x311 &  x433 &  x476 &  x511 &  x563 &  x799 &  x1046 & ~x141 & ~x142 & ~x201 & ~x219 & ~x241 & ~x258 & ~x280;
assign c0160 =  x86 &  x392 &  x433 &  x458 &  x563 &  x588 &  x620 &  x627 &  x782 &  x793 &  x832 &  x871 &  x916 &  x944 &  x949 &  x955 &  x994 &  x1072 & ~x294;
assign c0162 =  x131 &  x134 &  x254 &  x392 &  x482 &  x557 &  x650 &  x664 &  x686 &  x703 &  x742 &  x745 &  x758 &  x820 &  x823 &  x859 &  x861 &  x898 &  x900 &  x901 &  x929 &  x939 &  x976 &  x978 &  x979 &  x1018 &  x1057 &  x1085 & ~x120 & ~x198 & ~x237 & ~x276 & ~x354 & ~x432 & ~x648 & ~x708 & ~x747 & ~x786 & ~x825;
assign c0164 =  x26 &  x59 &  x68 &  x176 &  x182 &  x218 &  x242 &  x308 &  x590 &  x608 &  x644 &  x656 &  x665 &  x893 &  x902 &  x1058 &  x1067 & ~x69 & ~x186 & ~x735 & ~x819 & ~x855 & ~x930 & ~x963 & ~x969 & ~x1002 & ~x1041 & ~x1080 & ~x1086 & ~x1125;
assign c0166 =  x8 &  x26 &  x29 &  x59 &  x62 &  x68 &  x113 &  x122 &  x125 &  x140 &  x143 &  x149 &  x152 &  x164 &  x191 &  x203 &  x212 &  x215 &  x218 &  x245 &  x254 &  x263 &  x299 &  x305 &  x362 &  x368 &  x392 &  x398 &  x410 &  x416 &  x422 &  x425 &  x428 &  x449 &  x458 &  x464 &  x476 &  x500 &  x512 &  x515 &  x533 &  x536 &  x563 &  x566 &  x575 &  x578 &  x585 &  x586 &  x596 &  x599 &  x605 &  x617 &  x624 &  x625 &  x662 &  x664 &  x671 &  x677 &  x692 &  x703 &  x707 &  x719 &  x731 &  x740 &  x743 &  x746 &  x758 &  x767 &  x788 &  x791 &  x800 &  x812 &  x848 &  x861 &  x866 &  x872 &  x890 &  x898 &  x900 &  x902 &  x908 &  x917 &  x929 &  x940 &  x950 &  x971 &  x979 &  x998 &  x1004 &  x1018 &  x1034 &  x1037 &  x1049 &  x1052 &  x1055 &  x1057 &  x1061 &  x1073 &  x1076 &  x1091 &  x1109 &  x1112 &  x1130 & ~x432 & ~x471;
assign c0168 =  x59 &  x71 &  x104 &  x149 &  x155 &  x182 &  x275 &  x284 &  x338 &  x356 &  x394 &  x433 &  x449 &  x452 &  x458 &  x554 &  x569 &  x587 &  x599 &  x644 &  x689 &  x704 &  x719 &  x737 &  x754 &  x758 &  x793 &  x803 &  x831 &  x832 &  x854 &  x870 &  x871 &  x881 &  x902 &  x920 &  x941 &  x944 &  x949 &  x968 &  x1027 &  x1064 &  x1073 &  x1105 &  x1130 & ~x336 & ~x375 & ~x453 & ~x858;
assign c0170 =  x20 &  x71 &  x221 &  x236 &  x284 &  x362 &  x374 &  x429 &  x449 &  x468 &  x563 &  x566 &  x586 &  x605 &  x664 &  x665 &  x703 &  x742 &  x749 &  x932 &  x1010 & ~x436 & ~x474 & ~x475 & ~x513 & ~x514 & ~x552 & ~x708;
assign c0172 =  x260 &  x507 &  x546 &  x586 &  x625 &  x664 &  x703 &  x730 &  x875 &  x989 &  x1091 & ~x453 & ~x474 & ~x513 & ~x514 & ~x552 & ~x553 & ~x708 & ~x747;
assign c0174 =  x2 &  x44 &  x50 &  x53 &  x68 &  x86 &  x98 &  x137 &  x155 &  x167 &  x173 &  x200 &  x206 &  x218 &  x260 &  x299 &  x305 &  x394 &  x430 &  x433 &  x497 &  x511 &  x554 &  x617 &  x644 &  x647 &  x674 &  x683 &  x706 &  x716 &  x719 &  x725 &  x740 &  x809 &  x812 &  x824 &  x854 &  x872 &  x941 &  x956 &  x959 &  x971 &  x1040 &  x1049 &  x1052 &  x1094 &  x1109 &  x1121 & ~x33 & ~x72 & ~x336 & ~x375 & ~x396 & ~x441 & ~x453 & ~x480 & ~x516;
assign c0176 =  x328 &  x356 &  x429 &  x452 &  x468 &  x469 &  x586 &  x587 &  x625 &  x664 &  x665 &  x703 &  x713 &  x737 &  x742 &  x761 &  x812 &  x1043 &  x1073 & ~x198 & ~x369 & ~x453 & ~x474 & ~x513 & ~x552 & ~x591;
assign c0178 =  x473 &  x494 &  x644 &  x664 &  x703 &  x859 &  x898 &  x979 &  x980 & ~x354 & ~x393 & ~x432 & ~x489 & ~x513 & ~x529 & ~x567 & ~x708;
assign c0180 =  x41 &  x122 &  x152 &  x161 &  x263 &  x275 &  x356 &  x413 &  x425 &  x473 &  x587 &  x588 &  x627 &  x628 &  x809 &  x811 &  x839 &  x848 &  x857 &  x890 &  x904 &  x943 &  x955 &  x968 &  x982 &  x1021 &  x1049 &  x1072 &  x1076 &  x1079 &  x1109 & ~x177 & ~x294 & ~x819;
assign c0182 =  x14 &  x17 &  x128 &  x173 &  x290 &  x311 &  x356 &  x371 &  x377 &  x400 &  x410 &  x439 &  x445 &  x479 &  x484 &  x523 &  x536 &  x541 &  x562 &  x575 &  x601 &  x625 &  x626 &  x650 &  x663 &  x664 &  x671 &  x689 &  x702 &  x707 &  x741 &  x742 &  x752 &  x782 &  x812 &  x819 &  x824 &  x848 &  x863 &  x881 &  x923 &  x936 &  x940 &  x950 &  x956 &  x959 &  x974 &  x1018 &  x1019 &  x1034 &  x1085 &  x1091 &  x1118 &  x1130 & ~x669;
assign c0184 =  x5 &  x52 &  x71 &  x91 &  x206 &  x251 &  x335 &  x389 &  x392 &  x395 &  x449 &  x470 &  x479 &  x485 &  x515 &  x554 &  x563 &  x589 &  x605 &  x629 &  x650 &  x710 &  x746 &  x767 &  x811 &  x850 &  x910 &  x949 &  x998 &  x1025 &  x1031 &  x1037 &  x1049 &  x1066 &  x1085 &  x1105 & ~x177 & ~x579 & ~x1086;
assign c0186 =  x82 &  x104 &  x137 &  x156 &  x164 &  x173 &  x185 &  x203 &  x221 &  x234 &  x251 &  x260 &  x274 &  x275 &  x299 &  x314 &  x332 &  x338 &  x344 &  x355 &  x356 &  x383 &  x386 &  x394 &  x431 &  x433 &  x443 &  x485 &  x503 &  x542 &  x569 &  x626 &  x629 &  x686 &  x689 &  x721 &  x746 &  x755 &  x758 &  x760 &  x791 &  x830 &  x833 &  x838 &  x854 &  x877 &  x878 &  x908 &  x947 &  x956 &  x965 &  x968 &  x1022 &  x1034 &  x1064 &  x1085 &  x1109 & ~x102 & ~x123 & ~x141 & ~x162 & ~x201 & ~x324 & ~x741 & ~x780 & ~x897;
assign c0188 =  x5 &  x32 &  x44 &  x83 &  x86 &  x122 &  x131 &  x143 &  x149 &  x191 &  x200 &  x245 &  x284 &  x287 &  x326 &  x332 &  x338 &  x344 &  x429 &  x430 &  x455 &  x468 &  x476 &  x479 &  x515 &  x518 &  x547 &  x586 &  x590 &  x608 &  x625 &  x629 &  x644 &  x647 &  x650 &  x659 &  x664 &  x683 &  x689 &  x698 &  x737 &  x742 &  x758 &  x761 &  x815 &  x827 &  x848 &  x923 &  x941 &  x944 &  x956 &  x968 &  x1049 &  x1073 &  x1130 & ~x237 & ~x276 & ~x315 & ~x453 & ~x474 & ~x513 & ~x552 & ~x591 & ~x594 & ~x675;
assign c0190 =  x182 &  x224 &  x338 &  x433 &  x797 &  x878 &  x1066 & ~x33 & ~x138 & ~x294 & ~x339 & ~x523;
assign c0192 =  x251 &  x356 &  x467 &  x491 &  x625 &  x664 &  x758 &  x788 &  x859 &  x1018 &  x1025 &  x1052 &  x1124 & ~x123 & ~x396 & ~x708 & ~x747 & ~x867 & ~x1011 & ~x1050 & ~x1089;
assign c0194 =  x2 &  x5 &  x17 &  x41 &  x50 &  x74 &  x101 &  x164 &  x233 &  x245 &  x278 &  x305 &  x326 &  x353 &  x365 &  x373 &  x383 &  x412 &  x425 &  x455 &  x485 &  x499 &  x514 &  x521 &  x533 &  x539 &  x542 &  x581 &  x590 &  x598 &  x632 &  x637 &  x653 &  x799 &  x805 &  x812 &  x838 &  x857 &  x875 &  x877 &  x878 &  x883 &  x887 &  x908 &  x917 &  x922 &  x932 &  x944 &  x959 &  x986 &  x989 &  x1010 &  x1013 &  x1016 &  x1019 &  x1049 &  x1061 &  x1076 &  x1109 &  x1121 & ~x768;
assign c0196 =  x149 &  x173 &  x377 &  x656 &  x755 &  x776 &  x821 &  x848 &  x908 &  x968 &  x1015 &  x1057 &  x1095 &  x1109 & ~x630 & ~x708 & ~x1012 & ~x1129;
assign c0198 =  x41 &  x65 &  x77 &  x152 &  x161 &  x164 &  x170 &  x206 &  x266 &  x275 &  x347 &  x356 &  x425 &  x428 &  x506 &  x628 &  x689 &  x707 &  x749 &  x830 &  x863 &  x875 &  x890 &  x911 &  x920 &  x998 &  x1019 &  x1109 &  x1118 &  x1127 & ~x27 & ~x339 & ~x534 & ~x555 & ~x696 & ~x697;
assign c0200 =  x2 &  x11 &  x44 &  x47 &  x56 &  x59 &  x77 &  x83 &  x98 &  x107 &  x125 &  x155 &  x161 &  x191 &  x194 &  x257 &  x260 &  x265 &  x281 &  x296 &  x299 &  x302 &  x323 &  x326 &  x344 &  x368 &  x392 &  x398 &  x401 &  x442 &  x461 &  x467 &  x470 &  x488 &  x509 &  x527 &  x542 &  x547 &  x554 &  x581 &  x586 &  x587 &  x596 &  x614 &  x617 &  x620 &  x625 &  x647 &  x653 &  x662 &  x664 &  x695 &  x722 &  x728 &  x731 &  x749 &  x791 &  x822 &  x823 &  x833 &  x845 &  x851 &  x872 &  x878 &  x887 &  x899 &  x902 &  x914 &  x920 &  x932 &  x935 &  x940 &  x950 &  x968 &  x979 &  x1001 &  x1022 &  x1031 &  x1049 &  x1091 &  x1118 & ~x198 & ~x237 & ~x354 & ~x393 & ~x432;
assign c0202 =  x17 &  x56 &  x74 &  x113 &  x221 &  x236 &  x242 &  x247 &  x254 &  x302 &  x325 &  x353 &  x364 &  x386 &  x431 &  x434 &  x442 &  x445 &  x449 &  x476 &  x481 &  x512 &  x562 &  x602 &  x664 &  x683 &  x686 &  x703 &  x742 &  x758 &  x769 &  x785 &  x794 &  x808 &  x820 &  x821 &  x881 &  x887 &  x898 &  x902 &  x953 &  x968 &  x971 &  x976 &  x1004 &  x1015 &  x1046 &  x1054 &  x1106 &  x1130 & ~x120 & ~x198 & ~x237 & ~x276 & ~x315 & ~x354 & ~x432 & ~x471;
assign c0204 =  x2 &  x5 &  x44 &  x62 &  x71 &  x89 &  x98 &  x104 &  x134 &  x137 &  x140 &  x143 &  x149 &  x173 &  x176 &  x188 &  x209 &  x215 &  x233 &  x263 &  x287 &  x320 &  x335 &  x383 &  x410 &  x416 &  x428 &  x515 &  x527 &  x536 &  x547 &  x560 &  x572 &  x581 &  x586 &  x587 &  x590 &  x593 &  x611 &  x625 &  x632 &  x641 &  x644 &  x650 &  x664 &  x665 &  x683 &  x695 &  x703 &  x713 &  x719 &  x725 &  x742 &  x758 &  x770 &  x781 &  x782 &  x820 &  x824 &  x839 &  x842 &  x848 &  x854 &  x859 &  x860 &  x866 &  x893 &  x898 &  x917 &  x929 &  x932 &  x937 &  x947 &  x959 &  x968 &  x976 &  x979 &  x983 &  x986 &  x1004 &  x1015 &  x1018 &  x1022 &  x1034 &  x1037 &  x1040 &  x1043 &  x1057 &  x1058 &  x1091 &  x1109 &  x1112 &  x1130 & ~x135 & ~x393 & ~x432 & ~x567 & ~x570 & ~x591 & ~x630 & ~x669 & ~x708 & ~x747 & ~x786;
assign c0206 =  x23 &  x29 &  x53 &  x56 &  x77 &  x83 &  x92 &  x146 &  x152 &  x182 &  x203 &  x206 &  x209 &  x218 &  x227 &  x263 &  x278 &  x284 &  x293 &  x299 &  x305 &  x326 &  x335 &  x338 &  x341 &  x365 &  x431 &  x437 &  x470 &  x515 &  x518 &  x521 &  x524 &  x542 &  x548 &  x586 &  x587 &  x589 &  x602 &  x608 &  x617 &  x625 &  x626 &  x632 &  x647 &  x650 &  x664 &  x689 &  x703 &  x705 &  x707 &  x719 &  x737 &  x744 &  x783 &  x822 &  x823 &  x854 &  x861 &  x881 &  x900 &  x938 &  x939 &  x941 &  x947 &  x959 &  x968 &  x979 &  x983 &  x988 &  x1018 &  x1043 &  x1049 &  x1055 &  x1057 &  x1072 &  x1076 &  x1082 & ~x795 & ~x834;
assign c0208 =  x104 &  x137 &  x140 &  x149 &  x158 &  x173 &  x185 &  x248 &  x263 &  x275 &  x281 &  x287 &  x290 &  x299 &  x314 &  x338 &  x344 &  x351 &  x365 &  x425 &  x430 &  x443 &  x455 &  x479 &  x542 &  x547 &  x586 &  x596 &  x614 &  x626 &  x628 &  x647 &  x650 &  x653 &  x665 &  x671 &  x677 &  x689 &  x698 &  x737 &  x758 &  x767 &  x812 &  x854 &  x881 &  x887 &  x941 &  x959 &  x968 &  x971 &  x989 &  x1055 &  x1076 & ~x291 & ~x330 & ~x369 & ~x375 & ~x435 & ~x474 & ~x513 & ~x516 & ~x552 & ~x555;
assign c0210 =  x74 &  x125 &  x128 &  x149 &  x161 &  x176 &  x194 &  x206 &  x227 &  x242 &  x245 &  x263 &  x278 &  x320 &  x323 &  x332 &  x353 &  x356 &  x394 &  x433 &  x443 &  x472 &  x515 &  x521 &  x542 &  x545 &  x548 &  x563 &  x628 &  x632 &  x659 &  x709 &  x719 &  x761 &  x767 &  x818 &  x832 &  x836 &  x857 &  x881 &  x884 &  x944 &  x980 &  x1043 &  x1070 &  x1085 &  x1121 & ~x138 & ~x741 & ~x819 & ~x930 & ~x963 & ~x969 & ~x1002 & ~x1008 & ~x1041 & ~x1047 & ~x1080;
assign c0212 =  x11 &  x26 &  x32 &  x47 &  x134 &  x149 &  x154 &  x155 &  x158 &  x182 &  x185 &  x193 &  x232 &  x233 &  x245 &  x265 &  x332 &  x338 &  x377 &  x419 &  x425 &  x461 &  x473 &  x500 &  x527 &  x566 &  x596 &  x602 &  x623 &  x625 &  x632 &  x650 &  x659 &  x664 &  x677 &  x683 &  x689 &  x704 &  x707 &  x710 &  x719 &  x742 &  x746 &  x781 &  x859 &  x881 &  x898 &  x902 &  x941 &  x944 &  x953 &  x956 &  x976 &  x979 &  x998 &  x1013 &  x1018 &  x1031 &  x1037 &  x1052 &  x1070 &  x1073 &  x1088 &  x1097 & ~x237 & ~x276 & ~x315 & ~x354 & ~x393 & ~x432 & ~x471 & ~x549 & ~x708 & ~x747 & ~x786 & ~x825 & ~x864 & ~x903 & ~x942;
assign c0214 =  x251 &  x260 &  x299 &  x338 &  x344 &  x380 &  x407 &  x419 &  x422 &  x428 &  x470 &  x479 &  x500 &  x518 &  x539 &  x557 &  x563 &  x575 &  x680 &  x794 &  x830 &  x845 &  x854 &  x857 &  x908 &  x916 &  x941 &  x944 &  x954 &  x955 &  x968 &  x983 &  x993 &  x994 &  x1004 &  x1039 &  x1049 &  x1072 &  x1073 &  x1082 &  x1109 & ~x6 & ~x138 & ~x177 & ~x561;
assign c0216 =  x17 &  x29 &  x35 &  x44 &  x59 &  x74 &  x86 &  x107 &  x116 &  x131 &  x134 &  x137 &  x152 &  x158 &  x161 &  x185 &  x200 &  x206 &  x209 &  x212 &  x218 &  x227 &  x245 &  x266 &  x284 &  x287 &  x320 &  x323 &  x332 &  x344 &  x356 &  x362 &  x401 &  x404 &  x443 &  x464 &  x500 &  x509 &  x515 &  x557 &  x581 &  x587 &  x602 &  x644 &  x671 &  x701 &  x704 &  x722 &  x745 &  x758 &  x767 &  x770 &  x783 &  x800 &  x809 &  x815 &  x822 &  x827 &  x854 &  x884 &  x893 &  x901 &  x914 &  x929 &  x971 &  x979 &  x995 &  x1007 &  x1022 &  x1055 &  x1061 &  x1130 & ~x54 & ~x93 & ~x138 & ~x144 & ~x177 & ~x222 & ~x306 & ~x339 & ~x495;
assign c0218 =  x104 &  x155 &  x206 &  x209 &  x274 &  x293 &  x302 &  x312 &  x344 &  x433 &  x437 &  x446 &  x467 &  x469 &  x698 &  x719 &  x832 &  x877 &  x916 &  x968 &  x995 &  x1115 & ~x336 & ~x375 & ~x516 & ~x555 & ~x819;
assign c0220 =  x232 &  x247 &  x299 &  x395 &  x629 &  x703 &  x710 &  x898 &  x900 &  x976 &  x978 &  x989 &  x1015 &  x1016 &  x1017 &  x1056 &  x1057 &  x1104;
assign c0222 =  x5 &  x26 &  x32 &  x41 &  x53 &  x56 &  x89 &  x98 &  x113 &  x116 &  x155 &  x170 &  x179 &  x188 &  x197 &  x206 &  x212 &  x245 &  x254 &  x260 &  x263 &  x275 &  x281 &  x287 &  x290 &  x299 &  x308 &  x323 &  x335 &  x347 &  x353 &  x356 &  x362 &  x365 &  x380 &  x382 &  x383 &  x386 &  x401 &  x419 &  x422 &  x425 &  x440 &  x446 &  x458 &  x470 &  x527 &  x539 &  x557 &  x566 &  x575 &  x587 &  x596 &  x599 &  x602 &  x605 &  x608 &  x614 &  x620 &  x623 &  x625 &  x626 &  x635 &  x641 &  x662 &  x664 &  x668 &  x680 &  x692 &  x698 &  x703 &  x707 &  x733 &  x734 &  x742 &  x749 &  x752 &  x772 &  x788 &  x794 &  x800 &  x806 &  x810 &  x815 &  x830 &  x845 &  x848 &  x857 &  x859 &  x860 &  x863 &  x884 &  x898 &  x911 &  x923 &  x929 &  x940 &  x944 &  x968 &  x976 &  x979 &  x983 &  x1015 &  x1018 &  x1043 &  x1057 &  x1058 &  x1073 &  x1096 &  x1100 &  x1103 &  x1112 &  x1121 &  x1127 &  x1130;
assign c0224 =  x11 &  x104 &  x128 &  x194 &  x212 &  x227 &  x293 &  x305 &  x323 &  x371 &  x403 &  x449 &  x455 &  x494 &  x500 &  x539 &  x572 &  x611 &  x650 &  x713 &  x770 &  x776 &  x820 &  x842 &  x854 &  x859 &  x878 &  x920 &  x950 &  x976 &  x979 &  x995 &  x1004 &  x1010 &  x1061 &  x1100 &  x1109 &  x1112 & ~x81 & ~x120 & ~x198 & ~x237 & ~x354 & ~x747 & ~x765 & ~x834 & ~x864 & ~x903 & ~x972 & ~x1077;
assign c0226 =  x38 &  x134 &  x320 &  x335 &  x386 &  x442 &  x445 &  x481 &  x539 &  x562 &  x593 &  x625 &  x664 &  x703 &  x725 &  x742 &  x781 &  x808 &  x859 &  x896 &  x898 &  x976 &  x979 &  x1015 &  x1018 &  x1049 &  x1052 &  x1057 &  x1093 &  x1096 & ~x237 & ~x276 & ~x471 & ~x708;
assign c0228 =  x2 &  x68 &  x85 &  x124 &  x137 &  x143 &  x173 &  x182 &  x197 &  x247 &  x266 &  x275 &  x284 &  x286 &  x305 &  x320 &  x338 &  x380 &  x428 &  x464 &  x554 &  x590 &  x596 &  x611 &  x627 &  x635 &  x641 &  x704 &  x722 &  x734 &  x758 &  x767 &  x832 &  x890 &  x953 &  x968 &  x1004 &  x1022 &  x1091 &  x1127 & ~x294 & ~x333 & ~x474 & ~x513;
assign c0230 =  x14 &  x85 &  x131 &  x182 &  x247 &  x269 &  x344 &  x403 &  x442 &  x445 &  x587 &  x590 &  x611 &  x650 &  x703 &  x704 &  x737 &  x739 &  x758 &  x859 &  x898 &  x959 &  x962 &  x976 &  x979 &  x1007 &  x1049 &  x1057 & ~x198 & ~x237 & ~x276 & ~x315 & ~x354 & ~x393 & ~x432;
assign c0232 =  x155 &  x173 &  x209 &  x281 &  x312 &  x323 &  x332 &  x351 &  x353 &  x395 &  x430 &  x452 &  x473 &  x500 &  x518 &  x547 &  x560 &  x566 &  x586 &  x587 &  x589 &  x596 &  x628 &  x629 &  x638 &  x644 &  x668 &  x683 &  x707 &  x722 &  x725 &  x767 &  x821 &  x854 &  x899 &  x980 &  x1052 &  x1121 & ~x279 & ~x357 & ~x397 & ~x436 & ~x474 & ~x480 & ~x591;
assign c0234 =  x1 &  x43 &  x55 &  x73 &  x112 &  x151 &  x392 &  x400 &  x439 &  x502 &  x518 &  x523 &  x541 &  x644 &  x662 &  x695 &  x812 &  x854 &  x997 &  x1043 &  x1091 & ~x45 & ~x51;
assign c0236 =  x17 &  x59 &  x140 &  x155 &  x197 &  x224 &  x266 &  x273 &  x312 &  x355 &  x389 &  x394 &  x401 &  x413 &  x425 &  x431 &  x472 &  x572 &  x668 &  x698 &  x785 &  x800 &  x911 &  x932 &  x944 &  x983 &  x995 &  x1019 &  x1028 &  x1121 & ~x123 & ~x162 & ~x201 & ~x213 & ~x258 & ~x280 & ~x319 & ~x702 & ~x780;
assign c0238 =  x146 &  x161 &  x185 &  x218 &  x269 &  x275 &  x313 &  x432 &  x471 &  x538 &  x550 &  x589 &  x635 &  x637 &  x838 &  x842 &  x887 &  x1012 & ~x258 & ~x297;
assign c0240 =  x179 &  x202 &  x241 &  x247 &  x292 &  x356 &  x403 &  x442 &  x481 &  x523 &  x562 &  x742 &  x767 &  x812 &  x861 &  x881 &  x898 &  x900 &  x937 &  x939 &  x1017 &  x1056 &  x1057 &  x1095;
assign c0242 =  x4 &  x43 &  x104 &  x140 &  x215 &  x293 &  x394 &  x422 &  x505 &  x509 &  x518 &  x569 &  x682 &  x767 &  x770 &  x812 &  x838 &  x876 &  x915 &  x916 &  x954 &  x955 &  x1007 &  x1016 &  x1046 &  x1066 & ~x819 & ~x858;
assign c0244 =  x197 &  x395 &  x461 &  x515 &  x635 &  x812 &  x1124 & ~x120 & ~x159 & ~x474 & ~x513 & ~x552 & ~x555 & ~x567 & ~x595 & ~x634;
assign c0246 =  x8 &  x23 &  x26 &  x32 &  x53 &  x83 &  x107 &  x110 &  x119 &  x128 &  x134 &  x137 &  x167 &  x182 &  x185 &  x191 &  x206 &  x236 &  x251 &  x272 &  x332 &  x347 &  x350 &  x353 &  x389 &  x452 &  x494 &  x500 &  x557 &  x566 &  x572 &  x647 &  x650 &  x686 &  x689 &  x713 &  x758 &  x797 &  x818 &  x821 &  x833 &  x902 &  x905 &  x940 &  x944 &  x1010 &  x1052 &  x1055 &  x1061 &  x1070 &  x1073 &  x1103 &  x1109 &  x1118 &  x1124 & ~x33 & ~x105 & ~x138 & ~x177 & ~x201 & ~x216 & ~x255 & ~x294 & ~x339 & ~x489 & ~x513 & ~x534 & ~x963 & ~x1002 & ~x1041 & ~x1080;
assign c0248 =  x20 &  x49 &  x55 &  x80 &  x88 &  x94 &  x110 &  x113 &  x119 &  x127 &  x131 &  x134 &  x143 &  x164 &  x166 &  x173 &  x188 &  x212 &  x221 &  x248 &  x284 &  x287 &  x341 &  x350 &  x356 &  x389 &  x410 &  x430 &  x446 &  x468 &  x470 &  x473 &  x476 &  x479 &  x482 &  x485 &  x521 &  x557 &  x569 &  x575 &  x586 &  x590 &  x608 &  x625 &  x632 &  x716 &  x737 &  x758 &  x776 &  x782 &  x785 &  x803 &  x815 &  x872 &  x881 &  x905 &  x920 &  x971 &  x980 &  x997 &  x1013 &  x1025 &  x1034 &  x1037 &  x1058 &  x1064 &  x1067 &  x1076 &  x1085 &  x1091 &  x1100 & ~x396 & ~x474 & ~x555;
assign c0250 =  x14 &  x32 &  x71 &  x80 &  x83 &  x104 &  x107 &  x125 &  x137 &  x143 &  x155 &  x209 &  x260 &  x266 &  x275 &  x284 &  x293 &  x299 &  x308 &  x320 &  x325 &  x380 &  x392 &  x395 &  x398 &  x419 &  x428 &  x431 &  x440 &  x443 &  x476 &  x488 &  x494 &  x500 &  x515 &  x518 &  x560 &  x569 &  x593 &  x605 &  x608 &  x620 &  x629 &  x635 &  x644 &  x653 &  x677 &  x680 &  x689 &  x713 &  x737 &  x742 &  x745 &  x749 &  x755 &  x758 &  x767 &  x770 &  x776 &  x782 &  x784 &  x791 &  x820 &  x824 &  x827 &  x830 &  x859 &  x860 &  x862 &  x881 &  x896 &  x898 &  x902 &  x914 &  x939 &  x940 &  x941 &  x944 &  x959 &  x974 &  x976 &  x978 &  x979 &  x995 &  x998 &  x1004 &  x1015 &  x1017 &  x1018 &  x1037 &  x1055 &  x1056 &  x1057 &  x1064 &  x1070 &  x1076 &  x1082 &  x1118 &  x1130 & ~x306 & ~x513 & ~x708;
assign c0252 =  x254 &  x320 &  x433 &  x896 & ~x6 & ~x30 & ~x69 & ~x123 & ~x280;
assign c0254 =  x17 &  x374 &  x446 &  x628 &  x955 & ~x319 & ~x358 & ~x397 & ~x480 & ~x741;
assign c0256 =  x92 &  x128 &  x161 &  x182 &  x265 &  x382 &  x442 &  x481 &  x664 &  x702 &  x741 &  x770 &  x780 &  x819 &  x820 &  x851 &  x858 &  x859 &  x872 &  x897 &  x898 &  x899 &  x936 &  x968 &  x976 &  x1015 &  x1076 & ~x393 & ~x432 & ~x471 & ~x588 & ~x747 & ~x786 & ~x825 & ~x903 & ~x909;
assign c0258 =  x56 &  x107 &  x134 &  x149 &  x173 &  x182 &  x191 &  x200 &  x206 &  x215 &  x251 &  x263 &  x265 &  x272 &  x284 &  x287 &  x344 &  x353 &  x356 &  x365 &  x380 &  x395 &  x442 &  x443 &  x481 &  x497 &  x500 &  x518 &  x536 &  x551 &  x554 &  x560 &  x562 &  x563 &  x601 &  x629 &  x650 &  x662 &  x664 &  x665 &  x668 &  x671 &  x683 &  x698 &  x703 &  x719 &  x722 &  x737 &  x742 &  x776 &  x781 &  x794 &  x797 &  x820 &  x830 &  x842 &  x848 &  x854 &  x857 &  x859 &  x860 &  x866 &  x878 &  x881 &  x896 &  x898 &  x914 &  x929 &  x941 &  x976 &  x983 &  x995 &  x1015 &  x1022 &  x1049 &  x1054 &  x1057 &  x1064 &  x1076 &  x1093 &  x1100 &  x1112 & ~x120 & ~x159 & ~x198 & ~x237 & ~x276 & ~x315 & ~x354 & ~x393 & ~x432 & ~x471 & ~x510 & ~x549 & ~x630 & ~x708 & ~x747 & ~x786;
assign c0260 =  x59 &  x77 &  x167 &  x394 &  x452 &  x455 &  x494 &  x518 &  x550 &  x587 &  x689 &  x695 &  x740 &  x850 &  x871 &  x910 &  x943 &  x944 &  x949 &  x1006 &  x1007 &  x1066 & ~x138 & ~x177 & ~x222 & ~x294;
assign c0262 =  x263 &  x500 &  x518 &  x671 &  x758 &  x770 &  x858 &  x859 &  x897 &  x898 &  x936 &  x953 &  x968 &  x975 &  x978 &  x983 &  x1013 &  x1015 &  x1017 &  x1043 &  x1054 &  x1056 &  x1057 &  x1095 & ~x747 & ~x865 & ~x903 & ~x942;
assign c0264 =  x91 &  x101 &  x134 &  x170 &  x247 &  x325 &  x386 &  x461 &  x581 &  x664 &  x698 &  x739 &  x758 &  x761 &  x881 &  x939 &  x986 &  x1058 &  x1082 &  x1115 &  x1118 & ~x354 & ~x393 & ~x630;
assign c0266 =  x312 &  x351 &  x356 &  x473 &  x518 &  x734 &  x854 &  x1001 &  x1049 & ~x258 & ~x297 & ~x396 & ~x474 & ~x477 & ~x480 & ~x516 & ~x555 & ~x780;
assign c0268 =  x182 &  x206 &  x394 &  x500 &  x1006 & ~x339 & ~x736 & ~x820 & ~x1119;
assign c0270 =  x2 &  x23 &  x29 &  x32 &  x65 &  x83 &  x113 &  x143 &  x161 &  x167 &  x182 &  x193 &  x209 &  x218 &  x232 &  x233 &  x263 &  x266 &  x272 &  x287 &  x323 &  x368 &  x446 &  x479 &  x548 &  x551 &  x569 &  x581 &  x593 &  x617 &  x623 &  x629 &  x632 &  x650 &  x658 &  x683 &  x697 &  x698 &  x704 &  x731 &  x734 &  x779 &  x832 &  x839 &  x851 &  x866 &  x880 &  x881 &  x910 &  x911 &  x914 &  x919 &  x932 &  x957 &  x959 &  x980 &  x997 &  x1037 &  x1043 &  x1046 &  x1048 &  x1085 &  x1118;
assign c0272 =  x8 &  x17 &  x34 &  x41 &  x73 &  x98 &  x112 &  x151 &  x161 &  x179 &  x247 &  x293 &  x320 &  x344 &  x364 &  x392 &  x403 &  x428 &  x440 &  x442 &  x452 &  x479 &  x481 &  x497 &  x533 &  x542 &  x580 &  x586 &  x608 &  x625 &  x664 &  x674 &  x677 &  x695 &  x707 &  x779 &  x785 &  x791 &  x794 &  x854 &  x884 &  x979 &  x983 &  x1013 &  x1043 &  x1049 &  x1064 & ~x120 & ~x159 & ~x198 & ~x237 & ~x276 & ~x315 & ~x432;
assign c0274 =  x10 &  x38 &  x56 &  x79 &  x92 &  x117 &  x149 &  x156 &  x195 &  x196 &  x221 &  x234 &  x254 &  x263 &  x326 &  x344 &  x356 &  x365 &  x422 &  x433 &  x488 &  x509 &  x515 &  x527 &  x530 &  x533 &  x539 &  x557 &  x569 &  x578 &  x599 &  x642 &  x662 &  x665 &  x681 &  x682 &  x722 &  x725 &  x787 &  x799 &  x818 &  x857 &  x860 &  x902 &  x962 &  x986 &  x1085 &  x1100 &  x1106 &  x1127 & ~x624;
assign c0276 =  x44 &  x47 &  x74 &  x86 &  x98 &  x104 &  x140 &  x149 &  x182 &  x209 &  x266 &  x380 &  x403 &  x442 &  x445 &  x455 &  x497 &  x500 &  x533 &  x562 &  x663 &  x702 &  x703 &  x758 &  x767 &  x770 &  x820 &  x830 &  x859 &  x898 &  x902 &  x914 &  x929 &  x939 &  x941 &  x978 &  x1015 &  x1017 &  x1037 &  x1054 &  x1056 &  x1057 &  x1064 &  x1073 &  x1076 &  x1082 &  x1097;
assign c0278 =  x29 &  x50 &  x155 &  x156 &  x157 &  x195 &  x234 &  x274 &  x350 &  x359 &  x389 &  x425 &  x695 &  x716 &  x767 &  x832 &  x851 &  x1043 &  x1103 & ~x102 & ~x141 & ~x142 & ~x180 & ~x181 & ~x219 & ~x258 & ~x1017 & ~x1083;
assign c0280 =  x134 &  x143 &  x149 &  x173 &  x175 &  x182 &  x232 &  x338 &  x392 &  x500 &  x569 &  x689 &  x704 &  x737 &  x767 & ~x12 & ~x105 & ~x150 & ~x177 & ~x300 & ~x456 & ~x495 & ~x534 & ~x1080;
assign c0282 =  x8 &  x65 &  x125 &  x156 &  x195 &  x230 &  x234 &  x275 &  x308 &  x394 &  x433 &  x473 &  x482 &  x511 &  x515 &  x689 &  x713 &  x779 &  x838 &  x877 &  x896 &  x902 &  x1019 &  x1094 & ~x138 & ~x180 & ~x201 & ~x279 & ~x363;
assign c0284 =  x8 &  x11 &  x20 &  x29 &  x71 &  x74 &  x107 &  x128 &  x176 &  x191 &  x194 &  x260 &  x266 &  x269 &  x284 &  x338 &  x356 &  x365 &  x374 &  x392 &  x398 &  x425 &  x439 &  x455 &  x469 &  x470 &  x500 &  x508 &  x512 &  x518 &  x536 &  x547 &  x584 &  x586 &  x614 &  x616 &  x623 &  x625 &  x629 &  x638 &  x664 &  x701 &  x703 &  x716 &  x742 &  x749 &  x752 &  x758 &  x764 &  x812 &  x848 &  x859 &  x884 &  x896 &  x898 &  x902 &  x914 &  x941 &  x944 &  x956 &  x965 &  x971 &  x979 &  x992 &  x998 &  x1061 &  x1070 &  x1103 &  x1112 &  x1127 & ~x393 & ~x453 & ~x474 & ~x513 & ~x552;
assign c0286 =  x5 &  x68 &  x86 &  x107 &  x137 &  x140 &  x155 &  x164 &  x185 &  x206 &  x224 &  x254 &  x266 &  x313 &  x314 &  x355 &  x371 &  x383 &  x425 &  x434 &  x455 &  x472 &  x473 &  x491 &  x515 &  x590 &  x611 &  x733 &  x748 &  x761 &  x772 &  x805 &  x811 &  x832 &  x839 &  x850 &  x863 &  x877 &  x881 &  x883 &  x890 &  x902 &  x914 &  x935 &  x941 &  x956 &  x959 &  x980 &  x983 &  x992 &  x998 &  x1004 &  x1028 &  x1046 &  x1064 &  x1076 &  x1082 &  x1097 & ~x6 & ~x27;
assign c0288 =  x113 &  x245 &  x265 &  x305 &  x572 &  x664 &  x703 &  x742 &  x820 &  x859 &  x898 &  x941 &  x979 &  x995 &  x1046 & ~x150 & ~x228 & ~x306 & ~x345 & ~x354 & ~x432 & ~x630 & ~x708 & ~x747 & ~x969 & ~x1008;
assign c0290 =  x167 &  x356 &  x428 &  x508 &  x586 &  x617 &  x651 &  x652 &  x664 &  x690 &  x691 &  x703 &  x704 &  x730 &  x742 &  x758 &  x769 &  x808 &  x809 &  x859 &  x898 &  x941 &  x959 &  x968 &  x1055 & ~x120 & ~x198 & ~x237 & ~x276;
assign c0292 =  x20 &  x503 &  x509 &  x609 &  x640 &  x655 &  x658 &  x694 &  x757 &  x796 &  x911 &  x1010 &  x1082 &  x1091 & ~x6;
assign c0294 =  x43 &  x230 &  x355 &  x587 &  x592 &  x631 &  x676 &  x770 &  x773 &  x968 &  x995 &  x1021 &  x1024 &  x1052 &  x1060 &  x1063 &  x1081;
assign c0296 =  x17 &  x131 &  x176 &  x274 &  x312 &  x335 &  x351 &  x469 &  x497 &  x500 &  x503 &  x515 &  x518 &  x547 &  x586 &  x625 &  x644 &  x704 &  x842 &  x854 &  x1085 & ~x120 & ~x297 & ~x357 & ~x358 & ~x396 & ~x480;
assign c0298 =  x95 &  x137 &  x170 &  x185 &  x215 &  x275 &  x290 &  x329 &  x338 &  x353 &  x356 &  x425 &  x428 &  x431 &  x515 &  x518 &  x546 &  x547 &  x585 &  x586 &  x602 &  x624 &  x625 &  x664 &  x703 &  x704 &  x713 &  x742 &  x746 &  x752 &  x758 &  x767 &  x770 &  x809 &  x820 &  x854 &  x859 &  x860 &  x869 &  x898 &  x932 &  x979 &  x995 &  x1103 &  x1130 & ~x432 & ~x471 & ~x474 & ~x513 & ~x552 & ~x591 & ~x630 & ~x631 & ~x708 & ~x747;
assign c01 =  x457 &  x521 & ~x660 & ~x877 & ~x915 & ~x1032 & ~x1104;
assign c03 =  x22 &  x623 & ~x810 & ~x949 & ~x993;
assign c05 =  x101 &  x203 &  x212 &  x310 &  x376 &  x578 &  x596 &  x698 &  x868 &  x907 &  x946 &  x1037 & ~x429 & ~x810 & ~x999;
assign c07 =  x152 &  x343 &  x346 &  x385 &  x424 &  x607 &  x628 &  x965 & ~x312 & ~x507;
assign c09 =  x457 &  x648 & ~x430;
assign c011 =  x8 &  x274 &  x583 &  x1078 & ~x304 & ~x666 & ~x750;
assign c013 =  x158 &  x206 &  x343 &  x371 &  x386 &  x671 &  x751 &  x782 &  x845 &  x851 & ~x9 & ~x204 & ~x243 & ~x321 & ~x1032;
assign c015 =  x64 &  x1117 & ~x702 & ~x783 & ~x1029 & ~x1035 & ~x1068;
assign c019 =  x314 &  x771 &  x848 &  x889 & ~x411 & ~x624 & ~x627 & ~x666 & ~x705;
assign c021 =  x98 &  x142 &  x181 &  x187 &  x448 & ~x921 & ~x1056;
assign c023 =  x74 &  x83 &  x103 &  x115 &  x164 &  x173 &  x197 &  x281 &  x299 &  x323 &  x343 &  x376 &  x446 &  x470 &  x503 &  x526 &  x539 &  x563 &  x565 &  x566 &  x604 &  x752 &  x875 &  x917 &  x1016 &  x1040 &  x1088 &  x1118 & ~x654 & ~x810;
assign c025 =  x182 &  x395 &  x686 &  x790 &  x974 &  x1061 & ~x111 & ~x312 & ~x429 & ~x717 & ~x954 & ~x1035 & ~x1113;
assign c027 =  x2 &  x5 &  x158 &  x170 &  x173 &  x212 &  x320 &  x347 &  x491 &  x581 &  x602 &  x605 &  x635 &  x689 &  x698 &  x725 &  x773 &  x866 &  x881 &  x911 &  x986 &  x1034 & ~x156 & ~x195 & ~x312 & ~x612 & ~x822 & ~x861;
assign c029 =  x359 &  x503 &  x555 &  x1103 & ~x420 & ~x1035;
assign c031 =  x744 & ~x273 & ~x312 & ~x321 & ~x777 & ~x811;
assign c033 =  x136 &  x478 &  x634 &  x673 &  x856 &  x1084 &  x1117 &  x1123 & ~x1014;
assign c035 =  x673 &  x867 & ~x654;
assign c037 =  x436 &  x983 & ~x520 & ~x598;
assign c039 =  x448 &  x1099 & ~x996 & ~x1114;
assign c041 =  x904 & ~x642 & ~x784;
assign c043 =  x8 &  x109 &  x122 &  x148 &  x214 &  x253 &  x365 &  x409 &  x581 &  x644 &  x1001 & ~x462 & ~x696 & ~x837;
assign c045 =  x280 &  x511 &  x548 &  x764 & ~x561 & ~x720 & ~x900;
assign c047 = ~x720 & ~x862;
assign c049 = ~x461;
assign c051 =  x22 &  x487 & ~x429 & ~x753 & ~x873 & ~x1074;
assign c053 =  x250 &  x454 &  x945 & ~x966 & ~x999;
assign c055 =  x903 & ~x654 & ~x720 & ~x840;
assign c057 =  x65 &  x104 &  x185 &  x329 &  x509 &  x646 &  x668 &  x895 &  x896 & ~x225 & ~x420 & ~x576 & ~x615;
assign c059 =  x631 &  x723 & ~x564 & ~x642;
assign c061 =  x280 &  x722 &  x869 &  x1127 & ~x520 & ~x798;
assign c063 =  x661 &  x700 & ~x381 & ~x420 & ~x663 & ~x705 & ~x750 & ~x1014;
assign c065 =  x304 &  x349 &  x365 &  x416 &  x506 &  x829 & ~x810 & ~x873 & ~x1032;
assign c067 = ~x760 & ~x918 & ~x978;
assign c069 =  x238 &  x245 &  x251 &  x299 &  x314 &  x353 &  x575 &  x581 &  x632 &  x662 &  x665 &  x689 &  x695 &  x736 &  x782 &  x833 &  x835 &  x938 &  x1049 &  x1064 & ~x474 & ~x705 & ~x706 & ~x744 & ~x822;
assign c071 =  x19 &  x331 &  x686 & ~x690 & ~x729 & ~x939;
assign c073 =  x101 &  x110 &  x200 &  x218 &  x631 &  x713 &  x1052 &  x1117 & ~x628;
assign c075 =  x829 & ~x132 & ~x273 & ~x390 & ~x429 & ~x850;
assign c077 =  x2 &  x65 &  x137 &  x167 &  x179 &  x194 &  x299 &  x356 &  x383 &  x392 &  x473 &  x497 &  x524 &  x646 &  x671 &  x692 &  x727 &  x734 &  x749 &  x809 &  x833 &  x895 &  x917 &  x971 &  x986 &  x995 &  x1003 &  x1012 &  x1018 &  x1043 &  x1052 &  x1057 & ~x270;
assign c079 =  x53 &  x239 &  x368 &  x371 &  x409 &  x833 &  x884 & ~x0 & ~x156 & ~x804 & ~x978;
assign c081 =  x928 & ~x9 & ~x285 & ~x831 & ~x951 & ~x1113;
assign c083 = ~x50;
assign c085 =  x611 & ~x922 & ~x1072 & ~x1113;
assign c087 =  x136 &  x493 &  x686 &  x728 &  x1126 & ~x810 & ~x960;
assign c089 =  x149 & ~x429 & ~x618 & ~x678 & ~x913 & ~x991 & ~x1074;
assign c091 =  x23 &  x50 &  x110 &  x347 &  x425 &  x572 &  x575 &  x604 &  x863 & ~x9 & ~x48 & ~x429 & ~x1074;
assign c093 = ~x598 & ~x652 & ~x691;
assign c095 =  x250 &  x358 &  x489 &  x490 &  x529 &  x606 &  x645 &  x646;
assign c097 =  x65 &  x223 &  x386 &  x536 &  x635 &  x818 &  x974 & ~x273 & ~x390 & ~x711 & ~x1066 & ~x1104;
assign c099 =  x136 &  x197 &  x476 &  x494 &  x785 &  x902 &  x1034 &  x1067 & ~x564 & ~x624 & ~x627 & ~x666;
assign c0101 =  x5 &  x700 &  x881 & ~x285 & ~x465 & ~x486 & ~x522 & ~x642;
assign c0103 = ~x416;
assign c0105 =  x59 &  x97 &  x136 &  x191 &  x211 &  x287 &  x290 &  x305 &  x869 &  x929 &  x1121 & ~x543 & ~x621 & ~x660 & ~x732 & ~x876;
assign c0107 =  x280 &  x474 & ~x885;
assign c0109 =  x589 & ~x156 & ~x717 & ~x759 & ~x996 & ~x1029 & ~x1032 & ~x1035;
assign c0111 =  x211 &  x250 &  x856 & ~x312 & ~x561 & ~x720;
assign c0113 =  x14 &  x110 &  x113 &  x233 &  x260 &  x436 &  x454 &  x476 &  x512 &  x689 &  x782 &  x824 &  x892 &  x896 &  x986 &  x1012 & ~x939;
assign c0115 =  x266 &  x281 & ~x922 & ~x999 & ~x1075;
assign c0117 = ~x462 & ~x537 & ~x822 & ~x978;
assign c0119 =  x682 & ~x739;
assign c0121 =  x236 &  x398 &  x517 &  x556 &  x595 &  x673 &  x1114 &  x1119 & ~x720 & ~x759;
assign c0123 = ~x911;
assign c0125 =  x158 &  x452 &  x788 & ~x144 & ~x585 & ~x589;
assign c0127 =  x68 &  x125 &  x179 &  x353 &  x365 &  x431 &  x553 &  x583 &  x688 &  x740 &  x839 &  x932 & ~x304 & ~x627 & ~x666;
assign c0129 = ~x318 & ~x609 & ~x628 & ~x667 & ~x705;
assign c0131 = ~x329;
assign c0133 =  x172 &  x255 &  x376 & ~x1095;
assign c0135 =  x607 &  x700 & ~x48 & ~x204 & ~x285;
assign c0137 = ~x609 & ~x745;
assign c0139 =  x16 & ~x730 & ~x1104;
assign c0141 = ~x248;
assign c0143 =  x275 &  x362 &  x544 &  x692 &  x928 &  x1019 &  x1123 & ~x525 & ~x624 & ~x666 & ~x705 & ~x711 & ~x750;
assign c0145 =  x490 &  x567 &  x657 & ~x609 & ~x783;
assign c0147 =  x65 &  x74 &  x98 &  x155 &  x1078 &  x1117 & ~x234 & ~x822 & ~x828 & ~x861 & ~x1023;
assign c0149 = ~x667 & ~x1053;
assign c0151 =  x11 &  x22 &  x65 &  x217 &  x290 &  x644 &  x911 &  x947 &  x983 &  x1115 &  x1120 &  x1127 & ~x309 & ~x348 & ~x651 & ~x678;
assign c0153 = ~x119;
assign c0155 = ~x584;
assign c0157 =  x1004 & ~x91 & ~x411 & ~x666 & ~x846 & ~x900;
assign c0159 = ~x290;
assign c0163 =  x206 &  x256 &  x458 &  x491 &  x947 &  x1022 & ~x285 & ~x481 & ~x558 & ~x564;
assign c0165 =  x229 &  x268 &  x326 &  x496 & ~x654 & ~x717 & ~x756 & ~x811;
assign c0167 =  x224 &  x353 &  x398 &  x485 &  x683 &  x821 &  x833 &  x1100 & ~x372 & ~x411 & ~x462 & ~x585 & ~x586 & ~x618 & ~x625 & ~x711 & ~x828 & ~x867;
assign c0169 =  x121 & ~x411 & ~x666 & ~x706 & ~x744 & ~x783;
assign c0171 =  x23 &  x92 &  x116 &  x254 &  x326 &  x407 &  x590 &  x602 &  x686 &  x806 &  x818 &  x857 &  x875 &  x908 &  x965 &  x1025 &  x1127 & ~x3 & ~x687 & ~x876 & ~x915 & ~x949 & ~x954 & ~x987 & ~x988 & ~x1027 & ~x1065 & ~x1066;
assign c0173 =  x187 &  x250 &  x415 &  x907 & ~x993 & ~x1032;
assign c0175 =  x89 &  x146 &  x782 &  x953 &  x1123 & ~x24 & ~x792 & ~x987 & ~x1032 & ~x1062;
assign c0177 =  x295 &  x346 &  x415 &  x454 &  x607 &  x727 &  x931 &  x952;
assign c0179 =  x493 &  x688 & ~x75 & ~x547 & ~x711 & ~x828;
assign c0181 =  x250 &  x868 & ~x429 & ~x468 & ~x717 & ~x756 & ~x771;
assign c0183 =  x159 &  x244 &  x962 & ~x627 & ~x628;
assign c0185 =  x442 &  x649 & ~x405 & ~x546 & ~x625 & ~x645;
assign c0187 = ~x364 & ~x442 & ~x564 & ~x753;
assign c0189 = ~x521;
assign c0191 =  x98 &  x855 &  x1117 & ~x744 & ~x822;
assign c0193 =  x163 & ~x231 & ~x285 & ~x705 & ~x1014;
assign c0195 =  x595 & ~x264 & ~x460 & ~x462;
assign c0197 = ~x863;
assign c0199 =  x182 &  x194 &  x277 &  x544 &  x583 &  x622 &  x677 &  x698 &  x1117 & ~x444 & ~x627 & ~x666 & ~x750;
assign c0201 =  x136 &  x409 & ~x921 & ~x1056;
assign c0203 =  x103 &  x181 &  x497 &  x595 &  x928 &  x1117 & ~x744;
assign c0205 = ~x312 & ~x940 & ~x979;
assign c0207 =  x376 &  x906 & ~x582 & ~x999;
assign c0209 =  x136 & ~x156 & ~x360 & ~x873 & ~x1104;
assign c0211 =  x142 &  x374 &  x496 &  x529 &  x731 &  x1022 & ~x654 & ~x1056;
assign c0213 =  x143 &  x203 &  x256 &  x343 &  x376 &  x415 &  x449 &  x454 &  x487 &  x515 &  x706 &  x745 &  x755 &  x875 &  x907 &  x946 &  x1055 & ~x810;
assign c0215 =  x256 &  x373 &  x457 &  x1050 & ~x9;
assign c0217 =  x136 &  x710 & ~x273 & ~x993 & ~x999 & ~x1113;
assign c0219 =  x243 &  x931 & ~x745;
assign c0221 = ~x156 & ~x684 & ~x685 & ~x723 & ~x729 & ~x900;
assign c0223 =  x44 &  x407 &  x700 &  x704 &  x788 &  x805 &  x817 &  x1084 & ~x246 & ~x309 & ~x525;
assign c0225 =  x32 &  x449 &  x511 &  x749 &  x914 &  x989 &  x1085 & ~x156 & ~x783 & ~x978 & ~x1023;
assign c0227 =  x1085 & ~x580 & ~x798 & ~x837;
assign c0229 =  x2 &  x80 &  x116 &  x245 &  x257 &  x266 &  x335 &  x470 &  x557 &  x797 &  x947 &  x956 & ~x204 & ~x261 & ~x381 & ~x420 & ~x483 & ~x783 & ~x828;
assign c0231 =  x17 &  x29 &  x71 &  x218 &  x848 &  x1019 &  x1079 &  x1082 &  x1112 &  x1118 & ~x39 & ~x312 & ~x804 & ~x978;
assign c0233 =  x248 &  x376 & ~x126 & ~x156 & ~x660 & ~x1005;
assign c0235 =  x14 & ~x642 & ~x978 & ~x979;
assign c0237 =  x775 &  x928 &  x1019 &  x1117 & ~x705 & ~x706 & ~x783;
assign c0239 =  x409 &  x608 &  x667 & ~x756 & ~x876 & ~x954 & ~x999 & ~x1074 & ~x1113;
assign c0241 = ~x78 & ~x285 & ~x612 & ~x900;
assign c0243 =  x250 &  x289 &  x302 &  x323 &  x409 &  x604 &  x611 &  x665 &  x761 &  x907 &  x1034 &  x1036 & ~x429 & ~x468;
assign c0245 =  x74 &  x137 &  x155 &  x194 &  x215 &  x272 &  x320 &  x323 &  x437 &  x473 &  x563 &  x583 &  x631 &  x632 &  x661 &  x707 &  x845 &  x848 &  x905 &  x923 &  x1022 &  x1037 &  x1045 & ~x261 & ~x624 & ~x666 & ~x705 & ~x783 & ~x822 & ~x936;
assign c0247 =  x294 &  x973 & ~x420 & ~x537;
assign c0249 =  x579 & ~x744;
assign c0251 = ~x720 & ~x726 & ~x940;
assign c0253 =  x1 &  x83 &  x100 &  x211 &  x227 &  x250 &  x343 &  x358 &  x646 &  x812 &  x862 &  x868 &  x905 &  x946 &  x971 &  x1061;
assign c0255 =  x5 &  x20 &  x23 &  x62 &  x116 &  x152 &  x170 &  x188 &  x230 &  x233 &  x250 &  x302 &  x338 &  x356 &  x386 &  x413 &  x443 &  x467 &  x473 &  x482 &  x506 &  x512 &  x518 &  x563 &  x566 &  x569 &  x572 &  x575 &  x596 &  x604 &  x623 &  x659 &  x671 &  x686 &  x698 &  x701 &  x704 &  x725 &  x731 &  x740 &  x773 &  x776 &  x821 &  x827 &  x866 &  x908 &  x917 &  x935 &  x938 &  x953 &  x959 &  x977 &  x983 &  x986 &  x998 &  x1001 &  x1025 &  x1028 &  x1043 &  x1046 &  x1061 &  x1064 &  x1070 &  x1103 &  x1112 &  x1115 & ~x312 & ~x351 & ~x504 & ~x543 & ~x621;
assign c0257 =  x262 &  x409 &  x539 &  x604 & ~x39 & ~x312 & ~x429;
assign c0259 =  x31 &  x595 & ~x742;
assign c0261 =  x22 &  x61 &  x131 &  x167 &  x253 &  x299 &  x331 &  x334 &  x607 &  x608 &  x643 &  x646 &  x727 &  x728 &  x737 &  x1018 &  x1079;
assign c0263 = ~x459 & ~x531 & ~x823 & ~x862;
assign c0265 =  x350 &  x419 &  x848 & ~x717 & ~x738 & ~x757 & ~x954 & ~x999;
assign c0267 = ~x753 & ~x835 & ~x991 & ~x1029 & ~x1032 & ~x1035;
assign c0269 =  x250 &  x385 &  x436 &  x475 &  x649 &  x784 & ~x696;
assign c0271 =  x110 &  x171 &  x217 &  x649 &  x763 & ~x1104 & ~x1122;
assign c0273 =  x103 &  x142 &  x292 &  x409 &  x473 &  x1036 &  x1075 & ~x939 & ~x978;
assign c0275 =  x661 &  x1123 & ~x420 & ~x703 & ~x783;
assign c0277 = ~x334 & ~x357 & ~x628;
assign c0279 =  x6 & ~x627 & ~x1014;
assign c0281 =  x89 &  x185 &  x203 &  x596 &  x704 &  x731 &  x928 &  x1043 &  x1049 & ~x249 & ~x381 & ~x642 & ~x666 & ~x705 & ~x744 & ~x783 & ~x822;
assign c0283 =  x595 &  x856 & ~x388 & ~x642;
assign c0285 =  x17 & ~x156 & ~x312 & ~x945 & ~x981 & ~x1035 & ~x1101;
assign c0287 =  x16 &  x177 &  x248 &  x256 &  x295 &  x371 &  x392 &  x422 &  x461 &  x614 &  x689 &  x716 &  x830 &  x892 &  x904 &  x926 &  x970 &  x1031 &  x1049 &  x1052 &  x1109 & ~x822;
assign c0289 =  x258 &  x411;
assign c0291 =  x422 & ~x433 & ~x585 & ~x777;
assign c0293 =  x7 &  x237 &  x752 &  x776 &  x893 & ~x171 & ~x627;
assign c0295 = ~x911;
assign c0297 = ~x320;
assign c0299 = ~x87 & ~x273 & ~x609 & ~x768 & ~x978;
assign c10 =  x50 &  x80 &  x83 &  x140 &  x155 &  x164 &  x197 &  x209 &  x224 &  x257 &  x266 &  x293 &  x296 &  x299 &  x335 &  x341 &  x362 &  x365 &  x376 &  x404 &  x415 &  x425 &  x428 &  x443 &  x524 &  x569 &  x578 &  x623 &  x706 &  x710 &  x755 &  x761 &  x788 &  x800 &  x803 &  x861 &  x881 &  x900 &  x923 &  x939 &  x950 &  x965 &  x978 &  x1001 &  x1013 &  x1016 &  x1018 &  x1055 &  x1057 &  x1061 &  x1082 &  x1094 & ~x312 & ~x477 & ~x630 & ~x759 & ~x798 & ~x951 & ~x990 & ~x1029;
assign c12 =  x17 &  x20 &  x23 &  x35 &  x53 &  x62 &  x71 &  x86 &  x89 &  x113 &  x131 &  x152 &  x164 &  x176 &  x185 &  x197 &  x200 &  x203 &  x215 &  x218 &  x278 &  x290 &  x311 &  x314 &  x317 &  x326 &  x335 &  x338 &  x362 &  x365 &  x383 &  x398 &  x422 &  x428 &  x440 &  x455 &  x470 &  x473 &  x476 &  x503 &  x515 &  x539 &  x542 &  x551 &  x554 &  x560 &  x563 &  x566 &  x578 &  x581 &  x596 &  x599 &  x632 &  x641 &  x644 &  x653 &  x656 &  x683 &  x701 &  x713 &  x746 &  x770 &  x776 &  x784 &  x785 &  x797 &  x803 &  x812 &  x827 &  x842 &  x851 &  x857 &  x887 &  x901 &  x902 &  x938 &  x962 &  x965 &  x974 &  x986 &  x989 &  x992 &  x995 &  x1016 &  x1025 &  x1040 &  x1046 &  x1058 &  x1064 &  x1073 &  x1079 &  x1085 &  x1106 & ~x138 & ~x234 & ~x237 & ~x276 & ~x315 & ~x660 & ~x699 & ~x700 & ~x738 & ~x777 & ~x855 & ~x951 & ~x990 & ~x1029 & ~x1050 & ~x1068;
assign c14 =  x19 &  x41 &  x68 &  x218 &  x272 &  x317 &  x356 &  x368 &  x394 &  x440 &  x491 &  x511 &  x551 &  x578 &  x669 &  x670 &  x671 &  x695 &  x709 &  x731 &  x787 &  x838 &  x851 &  x890 &  x950 &  x971 &  x1034 & ~x585 & ~x606 & ~x645 & ~x663 & ~x741 & ~x939;
assign c16 =  x98 &  x131 &  x161 &  x176 &  x197 &  x266 &  x305 &  x308 &  x337 &  x338 &  x343 &  x356 &  x371 &  x421 &  x464 &  x493 &  x532 &  x565 &  x604 &  x640 &  x671 &  x725 &  x796 &  x1037 &  x1055 &  x1091 &  x1096 & ~x471 & ~x588 & ~x627 & ~x666 & ~x1032 & ~x1065 & ~x1104;
assign c18 =  x35 &  x37 &  x47 &  x53 &  x68 &  x76 &  x131 &  x137 &  x140 &  x152 &  x197 &  x203 &  x218 &  x227 &  x239 &  x263 &  x278 &  x329 &  x331 &  x338 &  x365 &  x370 &  x383 &  x392 &  x410 &  x416 &  x437 &  x458 &  x494 &  x500 &  x518 &  x578 &  x596 &  x599 &  x608 &  x611 &  x629 &  x656 &  x668 &  x674 &  x728 &  x731 &  x734 &  x765 &  x766 &  x785 &  x791 &  x800 &  x805 &  x844 &  x848 &  x857 &  x860 &  x866 &  x893 &  x902 &  x914 &  x917 &  x920 &  x965 &  x974 &  x980 &  x1016 &  x1025 &  x1040 &  x1043 &  x1097 &  x1100 & ~x762 & ~x801;
assign c110 =  x20 &  x26 &  x35 &  x56 &  x77 &  x86 &  x89 &  x92 &  x200 &  x218 &  x236 &  x254 &  x275 &  x277 &  x293 &  x305 &  x316 &  x322 &  x404 &  x413 &  x443 &  x473 &  x488 &  x553 &  x566 &  x569 &  x578 &  x599 &  x614 &  x635 &  x641 &  x674 &  x692 &  x695 &  x698 &  x715 &  x728 &  x731 &  x771 &  x800 &  x806 &  x851 &  x878 &  x890 &  x893 &  x896 &  x920 &  x950 &  x956 &  x959 &  x971 &  x977 &  x1007 &  x1010 &  x1016 &  x1022 &  x1061 &  x1088 &  x1100 & ~x372 & ~x585 & ~x702;
assign c112 =  x14 &  x53 &  x62 &  x71 &  x74 &  x82 &  x86 &  x95 &  x101 &  x119 &  x137 &  x164 &  x167 &  x179 &  x185 &  x212 &  x218 &  x224 &  x230 &  x266 &  x277 &  x278 &  x284 &  x287 &  x293 &  x305 &  x316 &  x344 &  x380 &  x394 &  x407 &  x410 &  x419 &  x422 &  x428 &  x443 &  x467 &  x470 &  x472 &  x473 &  x503 &  x506 &  x511 &  x512 &  x518 &  x521 &  x527 &  x530 &  x557 &  x563 &  x584 &  x587 &  x593 &  x599 &  x611 &  x635 &  x638 &  x650 &  x698 &  x716 &  x722 &  x737 &  x743 &  x746 &  x749 &  x761 &  x778 &  x788 &  x791 &  x809 &  x836 &  x844 &  x845 &  x850 &  x854 &  x856 &  x860 &  x866 &  x877 &  x883 &  x890 &  x922 &  x928 &  x938 &  x953 &  x956 &  x961 &  x967 &  x968 &  x971 &  x989 &  x998 &  x1000 &  x1013 &  x1016 &  x1019 &  x1028 &  x1039 &  x1040 &  x1046 &  x1051 &  x1058 &  x1082 &  x1084 &  x1090 &  x1103 &  x1115 &  x1117 &  x1118 &  x1123 &  x1129 & ~x444 & ~x702 & ~x897 & ~x936;
assign c114 =  x52 &  x119 &  x164 &  x254 &  x281 &  x383 &  x407 &  x443 &  x455 &  x464 &  x469 &  x511 &  x578 &  x584 &  x628 &  x668 &  x716 &  x761 &  x767 &  x773 &  x785 &  x857 &  x865 &  x896 &  x950 &  x953 &  x998 &  x1016 &  x1073 & ~x420 & ~x459 & ~x498 & ~x840 & ~x879 & ~x918 & ~x936 & ~x951 & ~x957 & ~x990 & ~x996 & ~x1029 & ~x1035 & ~x1068 & ~x1092;
assign c116 =  x68 &  x107 &  x116 &  x122 &  x214 &  x253 &  x302 &  x337 &  x365 &  x382 &  x383 &  x415 &  x448 &  x487 &  x526 &  x584 &  x605 &  x746 &  x767 &  x785 &  x940 &  x950 &  x962 &  x1016 &  x1076 &  x1115 & ~x87 & ~x126 & ~x432 & ~x594 & ~x1029;
assign c118 =  x37 &  x76 &  x119 &  x146 &  x232 &  x253 &  x271 &  x292 &  x320 &  x331 &  x335 &  x337 &  x344 &  x353 &  x376 &  x386 &  x388 &  x415 &  x421 &  x422 &  x440 &  x443 &  x452 &  x494 &  x526 &  x536 &  x554 &  x557 &  x572 &  x578 &  x584 &  x599 &  x605 &  x632 &  x656 &  x758 &  x890 &  x923 &  x946 &  x985 &  x1018 &  x1024 &  x1063 &  x1094 & ~x915;
assign c120 =  x415 &  x488 &  x491 &  x532 &  x539 &  x551 &  x559 &  x578 &  x640 &  x716 &  x742 &  x781 &  x820 &  x1015 &  x1096 & ~x738 & ~x855 & ~x888 & ~x966 & ~x1005 & ~x1044;
assign c122 =  x5 &  x29 &  x119 &  x242 &  x251 &  x269 &  x314 &  x317 &  x338 &  x341 &  x403 &  x446 &  x467 &  x557 &  x596 &  x611 &  x665 &  x680 &  x698 &  x716 &  x728 &  x746 &  x773 &  x818 &  x914 &  x1018 &  x1070 &  x1097 &  x1106 & ~x243 & ~x432 & ~x510 & ~x732 & ~x834 & ~x849 & ~x874 & ~x912 & ~x915 & ~x951 & ~x990 & ~x993 & ~x1029 & ~x1068;
assign c124 =  x11 &  x17 &  x41 &  x59 &  x77 &  x200 &  x203 &  x227 &  x249 &  x272 &  x288 &  x317 &  x328 &  x350 &  x367 &  x413 &  x425 &  x443 &  x461 &  x485 &  x488 &  x491 &  x524 &  x575 &  x578 &  x590 &  x605 &  x611 &  x623 &  x629 &  x650 &  x677 &  x695 &  x784 &  x785 &  x803 &  x896 &  x929 &  x956 &  x971 &  x1010 &  x1019 &  x1046 &  x1055 & ~x240 & ~x357 & ~x474 & ~x777;
assign c126 =  x17 &  x20 &  x113 &  x116 &  x119 &  x128 &  x203 &  x227 &  x275 &  x286 &  x311 &  x320 &  x335 &  x376 &  x392 &  x415 &  x422 &  x443 &  x452 &  x518 &  x536 &  x545 &  x554 &  x578 &  x593 &  x602 &  x665 &  x692 &  x713 &  x737 &  x749 &  x752 &  x773 &  x776 &  x800 &  x845 &  x900 &  x938 &  x939 &  x950 &  x965 &  x974 &  x1010 &  x1018 &  x1037 &  x1040 &  x1043 &  x1064 &  x1088 &  x1091 & ~x195 & ~x429 & ~x528 & ~x606 & ~x645 & ~x762 & ~x801 & ~x840 & ~x918;
assign c128 =  x20 &  x44 &  x74 &  x86 &  x110 &  x113 &  x116 &  x119 &  x152 &  x203 &  x224 &  x254 &  x263 &  x287 &  x293 &  x317 &  x323 &  x356 &  x368 &  x389 &  x404 &  x419 &  x437 &  x440 &  x443 &  x473 &  x491 &  x506 &  x518 &  x527 &  x572 &  x575 &  x578 &  x596 &  x605 &  x617 &  x629 &  x641 &  x647 &  x671 &  x692 &  x698 &  x710 &  x728 &  x746 &  x749 &  x751 &  x752 &  x784 &  x790 &  x803 &  x826 &  x828 &  x829 &  x833 &  x851 &  x865 &  x867 &  x868 &  x899 &  x901 &  x907 &  x932 &  x965 &  x977 &  x995 &  x1007 &  x1070 &  x1073 &  x1082 &  x1094 &  x1100 & ~x273 & ~x795 & ~x834 & ~x873 & ~x876 & ~x960;
assign c130 =  x11 &  x14 &  x23 &  x38 &  x62 &  x86 &  x98 &  x125 &  x142 &  x181 &  x200 &  x203 &  x220 &  x224 &  x254 &  x275 &  x443 &  x509 &  x527 &  x560 &  x578 &  x596 &  x628 &  x641 &  x667 &  x680 &  x706 &  x745 &  x767 &  x770 &  x773 &  x865 &  x883 &  x890 &  x904 &  x922 &  x961 &  x962 &  x995 &  x1000 &  x1039 &  x1076 &  x1117 & ~x360 & ~x513 & ~x795;
assign c132 =  x5 &  x14 &  x29 &  x35 &  x41 &  x47 &  x62 &  x65 &  x92 &  x95 &  x98 &  x104 &  x107 &  x122 &  x131 &  x140 &  x149 &  x155 &  x158 &  x185 &  x191 &  x227 &  x239 &  x242 &  x254 &  x287 &  x293 &  x314 &  x317 &  x329 &  x341 &  x344 &  x350 &  x353 &  x359 &  x362 &  x368 &  x395 &  x398 &  x440 &  x443 &  x446 &  x472 &  x473 &  x476 &  x488 &  x491 &  x494 &  x511 &  x530 &  x533 &  x545 &  x563 &  x572 &  x578 &  x587 &  x589 &  x590 &  x605 &  x614 &  x617 &  x623 &  x632 &  x638 &  x647 &  x650 &  x656 &  x659 &  x665 &  x667 &  x674 &  x680 &  x686 &  x692 &  x698 &  x701 &  x704 &  x707 &  x713 &  x731 &  x734 &  x745 &  x746 &  x748 &  x785 &  x787 &  x788 &  x800 &  x818 &  x824 &  x825 &  x826 &  x830 &  x833 &  x836 &  x845 &  x854 &  x865 &  x866 &  x872 &  x875 &  x884 &  x890 &  x893 &  x902 &  x905 &  x923 &  x929 &  x943 &  x944 &  x962 &  x974 &  x980 &  x1022 &  x1028 &  x1040 &  x1061 &  x1073 &  x1082 &  x1091 &  x1094 &  x1103 &  x1112 &  x1127 &  x1130 & ~x858 & ~x897 & ~x1014 & ~x1029 & ~x1053 & ~x1062 & ~x1068 & ~x1092 & ~x1101;
assign c134 =  x1 &  x21 &  x22 &  x38 &  x40 &  x47 &  x50 &  x61 &  x73 &  x99 &  x113 &  x138 &  x145 &  x172 &  x178 &  x215 &  x217 &  x272 &  x308 &  x317 &  x331 &  x367 &  x406 &  x410 &  x485 &  x506 &  x518 &  x578 &  x605 &  x671 &  x707 &  x784 &  x803 &  x926 &  x1097 & ~x966;
assign c136 =  x16 &  x35 &  x38 &  x83 &  x94 &  x125 &  x151 &  x172 &  x184 &  x211 &  x214 &  x223 &  x224 &  x227 &  x236 &  x253 &  x254 &  x266 &  x278 &  x284 &  x311 &  x317 &  x326 &  x341 &  x383 &  x413 &  x416 &  x419 &  x437 &  x461 &  x491 &  x527 &  x536 &  x566 &  x575 &  x578 &  x596 &  x623 &  x677 &  x686 &  x698 &  x709 &  x767 &  x790 &  x794 &  x832 &  x854 &  x871 &  x910 &  x935 &  x956 &  x977 &  x1004 &  x1022 &  x1058 &  x1088 & ~x720;
assign c138 =  x128 &  x271 &  x376 &  x382 &  x389 &  x395 &  x415 &  x421 &  x487 &  x562 &  x596 &  x664 &  x706 &  x905 &  x939 &  x1018 &  x1022 & ~x390 & ~x660 & ~x915 & ~x954 & ~x993;
assign c140 =  x2 &  x14 &  x38 &  x44 &  x50 &  x68 &  x86 &  x104 &  x113 &  x125 &  x143 &  x146 &  x176 &  x185 &  x191 &  x200 &  x203 &  x209 &  x227 &  x242 &  x254 &  x259 &  x278 &  x293 &  x314 &  x317 &  x329 &  x341 &  x347 &  x356 &  x368 &  x383 &  x395 &  x404 &  x425 &  x434 &  x440 &  x443 &  x470 &  x479 &  x482 &  x494 &  x511 &  x527 &  x533 &  x563 &  x578 &  x584 &  x589 &  x590 &  x593 &  x596 &  x608 &  x628 &  x629 &  x632 &  x647 &  x659 &  x667 &  x668 &  x706 &  x709 &  x725 &  x731 &  x743 &  x745 &  x746 &  x747 &  x752 &  x776 &  x784 &  x786 &  x787 &  x826 &  x845 &  x860 &  x865 &  x866 &  x869 &  x899 &  x904 &  x920 &  x944 &  x950 &  x956 &  x974 &  x995 &  x998 &  x1010 &  x1037 &  x1046 &  x1049 &  x1079 &  x1085 &  x1103 &  x1106 &  x1121 &  x1130 & ~x660 & ~x795;
assign c142 =  x74 &  x199 &  x206 &  x277 &  x437 &  x475 &  x536 &  x553 &  x559 &  x578 &  x637 &  x676 &  x715 &  x716 &  x860 &  x917 & ~x99 & ~x177 & ~x216 & ~x333 & ~x462 & ~x501;
assign c144 =  x5 &  x62 &  x65 &  x74 &  x89 &  x170 &  x185 &  x203 &  x242 &  x329 &  x392 &  x395 &  x449 &  x521 &  x527 &  x631 &  x632 &  x731 &  x752 &  x761 &  x782 &  x809 &  x836 &  x842 &  x848 &  x878 &  x881 &  x968 &  x1049 &  x1058 & ~x303 & ~x384 & ~x423 & ~x501 & ~x579 & ~x705 & ~x969 & ~x1005 & ~x1050;
assign c146 =  x41 &  x44 &  x47 &  x80 &  x83 &  x143 &  x173 &  x176 &  x199 &  x209 &  x224 &  x238 &  x248 &  x275 &  x277 &  x284 &  x290 &  x316 &  x392 &  x394 &  x413 &  x437 &  x473 &  x479 &  x491 &  x511 &  x512 &  x517 &  x527 &  x539 &  x542 &  x553 &  x560 &  x596 &  x616 &  x623 &  x655 &  x665 &  x715 &  x725 &  x752 &  x772 &  x791 &  x818 &  x821 &  x871 &  x899 &  x908 &  x910 &  x932 &  x938 &  x950 &  x953 &  x965 &  x995 &  x1007 &  x1016 &  x1046 &  x1100 & ~x444 & ~x486 & ~x507 & ~x546 & ~x585 & ~x702 & ~x741;
assign c148 =  x8 &  x14 &  x56 &  x65 &  x74 &  x80 &  x89 &  x119 &  x146 &  x176 &  x179 &  x191 &  x215 &  x218 &  x227 &  x236 &  x260 &  x278 &  x284 &  x305 &  x308 &  x311 &  x317 &  x335 &  x338 &  x347 &  x359 &  x376 &  x389 &  x403 &  x442 &  x455 &  x470 &  x473 &  x482 &  x487 &  x494 &  x512 &  x526 &  x533 &  x536 &  x554 &  x565 &  x566 &  x575 &  x578 &  x581 &  x593 &  x604 &  x641 &  x643 &  x665 &  x668 &  x692 &  x695 &  x698 &  x710 &  x713 &  x758 &  x767 &  x773 &  x776 &  x785 &  x800 &  x818 &  x827 &  x851 &  x890 &  x899 &  x914 &  x935 &  x941 &  x950 &  x956 &  x974 &  x980 &  x995 &  x1007 &  x1016 &  x1025 &  x1055 &  x1079 &  x1085 &  x1094 &  x1118 & ~x549 & ~x660 & ~x888 & ~x927 & ~x960 & ~x966 & ~x1005 & ~x1044 & ~x1083;
assign c150 =  x38 &  x40 &  x77 &  x83 &  x128 &  x185 &  x191 &  x275 &  x302 &  x317 &  x401 &  x406 &  x413 &  x415 &  x425 &  x445 &  x449 &  x527 &  x578 &  x626 &  x640 &  x728 &  x758 &  x767 &  x780 &  x820 &  x908 &  x914 &  x956 &  x976 & ~x276 & ~x432 & ~x792 & ~x909 & ~x948 & ~x954 & ~x993 & ~x1032;
assign c152 =  x8 &  x56 &  x70 &  x86 &  x125 &  x182 &  x203 &  x215 &  x259 &  x281 &  x298 &  x331 &  x376 &  x381 &  x389 &  x392 &  x404 &  x406 &  x407 &  x415 &  x443 &  x445 &  x452 &  x473 &  x527 &  x560 &  x562 &  x584 &  x596 &  x599 &  x640 &  x644 &  x707 &  x746 &  x767 &  x851 &  x863 &  x866 &  x890 &  x896 &  x968 &  x974 &  x989 &  x1010 &  x1118 & ~x351 & ~x429 & ~x471;
assign c154 =  x17 &  x29 &  x35 &  x41 &  x44 &  x53 &  x95 &  x143 &  x146 &  x164 &  x227 &  x254 &  x314 &  x362 &  x365 &  x389 &  x394 &  x410 &  x419 &  x440 &  x443 &  x461 &  x548 &  x596 &  x650 &  x671 &  x683 &  x692 &  x695 &  x701 &  x709 &  x712 &  x716 &  x728 &  x734 &  x749 &  x751 &  x767 &  x776 &  x787 &  x803 &  x818 &  x826 &  x844 &  x865 &  x875 &  x877 &  x883 &  x890 &  x902 &  x917 &  x922 &  x950 &  x956 &  x961 &  x994 &  x1000 &  x1004 &  x1007 &  x1010 &  x1027 &  x1032 &  x1039 &  x1071 &  x1130 & ~x663 & ~x702 & ~x741;
assign c156 =  x23 &  x35 &  x56 &  x59 &  x65 &  x74 &  x82 &  x86 &  x92 &  x95 &  x101 &  x121 &  x125 &  x143 &  x152 &  x160 &  x164 &  x173 &  x191 &  x199 &  x218 &  x235 &  x263 &  x266 &  x272 &  x275 &  x277 &  x290 &  x293 &  x296 &  x299 &  x313 &  x316 &  x355 &  x359 &  x371 &  x389 &  x394 &  x398 &  x413 &  x416 &  x440 &  x446 &  x461 &  x467 &  x475 &  x512 &  x530 &  x536 &  x539 &  x553 &  x581 &  x587 &  x592 &  x593 &  x596 &  x599 &  x631 &  x632 &  x641 &  x655 &  x677 &  x692 &  x695 &  x701 &  x749 &  x766 &  x767 &  x772 &  x785 &  x794 &  x800 &  x808 &  x809 &  x815 &  x838 &  x842 &  x845 &  x863 &  x884 &  x902 &  x908 &  x929 &  x938 &  x944 &  x947 &  x953 &  x956 &  x989 &  x995 &  x1007 &  x1010 &  x1025 &  x1040 &  x1043 &  x1046 &  x1085 &  x1088 &  x1091 &  x1112 & ~x153 & ~x327 & ~x624 & ~x663 & ~x702 & ~x705 & ~x744;
assign c158 =  x23 &  x176 &  x260 &  x302 &  x374 &  x494 &  x517 &  x556 &  x559 &  x595 &  x596 &  x673 &  x734 &  x753 &  x833 &  x920 &  x922 &  x961 &  x1000 &  x1049 &  x1051 &  x1058 &  x1067 &  x1070 &  x1090 &  x1123 &  x1127 &  x1129 & ~x663 & ~x702;
assign c160 =  x5 &  x38 &  x56 &  x74 &  x77 &  x80 &  x92 &  x95 &  x98 &  x116 &  x131 &  x152 &  x167 &  x182 &  x188 &  x191 &  x203 &  x206 &  x212 &  x227 &  x239 &  x245 &  x278 &  x281 &  x299 &  x317 &  x320 &  x329 &  x338 &  x347 &  x368 &  x374 &  x398 &  x404 &  x413 &  x416 &  x425 &  x428 &  x431 &  x446 &  x452 &  x455 &  x458 &  x461 &  x464 &  x470 &  x482 &  x491 &  x542 &  x563 &  x569 &  x578 &  x581 &  x586 &  x590 &  x596 &  x605 &  x623 &  x632 &  x650 &  x653 &  x664 &  x665 &  x668 &  x673 &  x674 &  x692 &  x695 &  x706 &  x712 &  x713 &  x716 &  x728 &  x731 &  x737 &  x743 &  x746 &  x751 &  x758 &  x761 &  x764 &  x770 &  x782 &  x790 &  x803 &  x806 &  x815 &  x821 &  x828 &  x829 &  x830 &  x842 &  x862 &  x865 &  x866 &  x867 &  x868 &  x872 &  x878 &  x896 &  x899 &  x901 &  x904 &  x905 &  x906 &  x907 &  x914 &  x917 &  x941 &  x946 &  x950 &  x956 &  x959 &  x965 &  x968 &  x971 &  x974 &  x980 &  x985 &  x998 &  x1019 &  x1022 &  x1034 &  x1040 &  x1043 &  x1082 &  x1094 &  x1100 &  x1109 &  x1112 &  x1127 & ~x759 & ~x798 & ~x837;
assign c162 =  x38 &  x50 &  x245 &  x314 &  x316 &  x329 &  x341 &  x394 &  x452 &  x455 &  x474 &  x513 &  x552 &  x631 &  x659 &  x716 &  x787 &  x794 &  x836 &  x1037 & ~x264 & ~x522 & ~x546 & ~x585 & ~x703 & ~x742;
assign c164 =  x35 &  x56 &  x68 &  x71 &  x86 &  x113 &  x122 &  x131 &  x176 &  x179 &  x185 &  x236 &  x314 &  x317 &  x320 &  x332 &  x335 &  x338 &  x341 &  x362 &  x383 &  x392 &  x406 &  x413 &  x416 &  x445 &  x482 &  x485 &  x500 &  x524 &  x536 &  x566 &  x575 &  x578 &  x584 &  x586 &  x647 &  x665 &  x680 &  x683 &  x689 &  x692 &  x701 &  x734 &  x758 &  x784 &  x785 &  x794 &  x823 &  x827 &  x829 &  x830 &  x862 &  x868 &  x869 &  x890 &  x908 &  x917 &  x920 &  x923 &  x932 &  x941 &  x950 &  x956 &  x962 &  x965 &  x968 &  x977 &  x1007 &  x1010 &  x1043 &  x1067 &  x1070 &  x1091 &  x1094 & ~x474 & ~x576 & ~x615 & ~x616 & ~x654 & ~x655 & ~x694 & ~x732 & ~x771 & ~x795 & ~x834;
assign c166 =  x5 &  x20 &  x32 &  x38 &  x44 &  x59 &  x116 &  x125 &  x137 &  x161 &  x164 &  x170 &  x176 &  x191 &  x203 &  x239 &  x242 &  x272 &  x278 &  x302 &  x305 &  x320 &  x323 &  x359 &  x362 &  x365 &  x382 &  x428 &  x434 &  x440 &  x443 &  x448 &  x452 &  x464 &  x476 &  x479 &  x487 &  x494 &  x526 &  x542 &  x554 &  x565 &  x578 &  x581 &  x584 &  x614 &  x620 &  x623 &  x701 &  x704 &  x713 &  x716 &  x725 &  x737 &  x773 &  x818 &  x851 &  x884 &  x956 &  x1010 &  x1061 &  x1064 &  x1067 &  x1079 &  x1085 &  x1088 &  x1096 &  x1097 & ~x126 & ~x165 & ~x204 & ~x321 & ~x399 & ~x432 & ~x471 & ~x738 & ~x993 & ~x1032 & ~x1068;
assign c168 =  x38 &  x68 &  x86 &  x125 &  x131 &  x176 &  x224 &  x227 &  x248 &  x284 &  x317 &  x368 &  x389 &  x434 &  x443 &  x521 &  x545 &  x640 &  x698 &  x716 &  x728 &  x734 &  x752 &  x761 &  x797 &  x818 &  x857 &  x860 &  x950 &  x956 &  x974 &  x1022 &  x1052 & ~x42 & ~x81 & ~x120 & ~x237 & ~x432 & ~x471 & ~x510 & ~x588 & ~x666 & ~x705 & ~x738 & ~x954 & ~x987 & ~x993 & ~x1026 & ~x1032;
assign c170 =  x11 &  x22 &  x40 &  x50 &  x60 &  x79 &  x92 &  x134 &  x139 &  x151 &  x155 &  x177 &  x185 &  x194 &  x215 &  x227 &  x254 &  x275 &  x314 &  x320 &  x338 &  x359 &  x368 &  x389 &  x392 &  x443 &  x484 &  x491 &  x512 &  x521 &  x623 &  x632 &  x641 &  x689 &  x692 &  x698 &  x725 &  x731 &  x749 &  x776 &  x779 &  x872 &  x875 &  x905 &  x932 &  x959 &  x971 &  x983 &  x985 &  x989 &  x995 &  x998 &  x1010 &  x1016 &  x1043 &  x1079 &  x1097 &  x1109 & ~x12 & ~x246 & ~x660;
assign c172 =  x14 &  x17 &  x35 &  x62 &  x68 &  x164 &  x218 &  x224 &  x242 &  x263 &  x272 &  x278 &  x284 &  x293 &  x302 &  x317 &  x335 &  x338 &  x353 &  x359 &  x383 &  x395 &  x413 &  x443 &  x452 &  x473 &  x511 &  x521 &  x527 &  x539 &  x542 &  x554 &  x578 &  x581 &  x602 &  x611 &  x641 &  x665 &  x670 &  x671 &  x695 &  x698 &  x709 &  x728 &  x734 &  x746 &  x747 &  x748 &  x761 &  x776 &  x787 &  x803 &  x818 &  x826 &  x842 &  x860 &  x865 &  x896 &  x905 &  x920 &  x938 &  x956 &  x965 &  x974 &  x1022 &  x1031 &  x1037 &  x1039 &  x1040 &  x1043 &  x1058 &  x1064 &  x1073 &  x1091 &  x1106 & ~x420 & ~x459 & ~x460 & ~x498 & ~x819 & ~x897 & ~x951 & ~x1092;
assign c174 =  x38 &  x53 &  x55 &  x82 &  x121 &  x160 &  x164 &  x199 &  x277 &  x302 &  x314 &  x316 &  x394 &  x407 &  x413 &  x422 &  x536 &  x554 &  x578 &  x676 &  x692 &  x709 &  x715 &  x719 &  x748 &  x806 &  x836 &  x851 &  x866 &  x871 &  x910 &  x928 &  x932 &  x938 &  x956 &  x989 &  x1007 &  x1106 & ~x684 & ~x723;
assign c176 =  x1 &  x40 &  x212 &  x215 &  x224 &  x278 &  x317 &  x371 &  x443 &  x446 &  x506 &  x554 &  x578 &  x596 &  x671 &  x731 &  x734 &  x776 &  x833 &  x847 &  x896 & ~x6 & ~x45 & ~x84 & ~x123 & ~x141 & ~x180 & ~x240 & ~x456 & ~x495;
assign c178 =  x2 &  x8 &  x14 &  x20 &  x35 &  x56 &  x59 &  x62 &  x68 &  x71 &  x83 &  x86 &  x95 &  x119 &  x125 &  x146 &  x152 &  x170 &  x188 &  x194 &  x197 &  x200 &  x227 &  x230 &  x242 &  x251 &  x260 &  x275 &  x278 &  x302 &  x311 &  x314 &  x317 &  x332 &  x335 &  x356 &  x365 &  x374 &  x380 &  x392 &  x407 &  x428 &  x440 &  x443 &  x449 &  x455 &  x467 &  x485 &  x491 &  x494 &  x509 &  x511 &  x512 &  x518 &  x527 &  x542 &  x551 &  x554 &  x578 &  x586 &  x589 &  x596 &  x602 &  x605 &  x623 &  x628 &  x641 &  x653 &  x662 &  x665 &  x667 &  x668 &  x671 &  x674 &  x692 &  x698 &  x706 &  x716 &  x734 &  x737 &  x745 &  x761 &  x773 &  x785 &  x794 &  x839 &  x854 &  x866 &  x881 &  x896 &  x908 &  x917 &  x935 &  x950 &  x956 &  x959 &  x968 &  x974 &  x980 &  x983 &  x995 &  x1007 &  x1010 &  x1016 &  x1037 &  x1040 &  x1046 &  x1058 &  x1064 &  x1085 & ~x321 & ~x360 & ~x477 & ~x678 & ~x720 & ~x756 & ~x759 & ~x795 & ~x798 & ~x834 & ~x912 & ~x951 & ~x990;
assign c180 =  x14 &  x35 &  x41 &  x98 &  x119 &  x146 &  x203 &  x227 &  x251 &  x338 &  x350 &  x353 &  x371 &  x428 &  x455 &  x470 &  x488 &  x511 &  x542 &  x641 &  x707 &  x713 &  x731 &  x746 &  x764 &  x787 &  x791 &  x803 &  x839 &  x842 &  x866 &  x971 &  x1006 &  x1034 &  x1067 &  x1094 &  x1109 & ~x87 & ~x624 & ~x663 & ~x696 & ~x702 & ~x717 & ~x774 & ~x795 & ~x834 & ~x936 & ~x996 & ~x1029 & ~x1035 & ~x1074;
assign c182 =  x40 &  x41 &  x79 &  x113 &  x164 &  x176 &  x194 &  x215 &  x224 &  x407 &  x448 &  x481 &  x487 &  x494 &  x526 &  x527 &  x532 &  x554 &  x695 &  x752 &  x770 &  x773 &  x800 &  x806 &  x827 &  x929 &  x1007 &  x1025 &  x1031 &  x1037 &  x1100 & ~x90 & ~x129 & ~x168 & ~x207 & ~x471 & ~x549 & ~x588 & ~x627 & ~x1026 & ~x1032 & ~x1071 & ~x1104;
assign c184 =  x11 &  x20 &  x26 &  x41 &  x47 &  x62 &  x68 &  x80 &  x86 &  x98 &  x101 &  x113 &  x116 &  x119 &  x125 &  x128 &  x146 &  x152 &  x158 &  x164 &  x173 &  x176 &  x179 &  x182 &  x197 &  x200 &  x203 &  x206 &  x212 &  x227 &  x245 &  x257 &  x275 &  x284 &  x296 &  x302 &  x314 &  x317 &  x320 &  x338 &  x341 &  x344 &  x347 &  x353 &  x365 &  x383 &  x389 &  x392 &  x395 &  x398 &  x407 &  x413 &  x416 &  x428 &  x434 &  x437 &  x443 &  x470 &  x476 &  x479 &  x488 &  x491 &  x494 &  x509 &  x515 &  x518 &  x545 &  x554 &  x572 &  x578 &  x581 &  x584 &  x590 &  x593 &  x596 &  x602 &  x608 &  x611 &  x617 &  x635 &  x638 &  x644 &  x653 &  x656 &  x662 &  x668 &  x671 &  x695 &  x713 &  x716 &  x722 &  x725 &  x734 &  x745 &  x749 &  x752 &  x770 &  x779 &  x784 &  x785 &  x788 &  x794 &  x800 &  x812 &  x815 &  x818 &  x833 &  x845 &  x851 &  x854 &  x857 &  x863 &  x866 &  x872 &  x875 &  x890 &  x896 &  x902 &  x905 &  x911 &  x920 &  x935 &  x950 &  x956 &  x965 &  x980 &  x989 &  x995 &  x998 &  x1001 &  x1007 &  x1010 &  x1037 &  x1040 &  x1064 &  x1070 &  x1076 &  x1079 &  x1091 &  x1094 &  x1109 &  x1112 &  x1118 & ~x66 & ~x228 & ~x267 & ~x321 & ~x384 & ~x411 & ~x450 & ~x489 & ~x528 & ~x840 & ~x873 & ~x879 & ~x912 & ~x918 & ~x951 & ~x957 & ~x990 & ~x996 & ~x1029 & ~x1035 & ~x1068 & ~x1107;
assign c186 =  x132 &  x171 &  x829 &  x865 &  x945 &  x946 &  x1024 &  x1063;
assign c188 =  x11 &  x47 &  x50 &  x71 &  x146 &  x170 &  x182 &  x185 &  x194 &  x200 &  x203 &  x227 &  x239 &  x242 &  x245 &  x259 &  x263 &  x271 &  x275 &  x278 &  x284 &  x298 &  x305 &  x310 &  x317 &  x325 &  x326 &  x331 &  x337 &  x340 &  x404 &  x416 &  x440 &  x443 &  x445 &  x470 &  x479 &  x482 &  x484 &  x539 &  x584 &  x593 &  x596 &  x602 &  x605 &  x628 &  x656 &  x668 &  x706 &  x707 &  x734 &  x755 &  x776 &  x784 &  x797 &  x809 &  x818 &  x851 &  x863 &  x890 &  x896 &  x902 &  x904 &  x914 &  x938 &  x940 &  x946 &  x956 &  x962 &  x977 &  x980 &  x985 &  x1007 &  x1018 &  x1021 &  x1024 &  x1063 &  x1091 & ~x351;
assign c190 =  x32 &  x35 &  x107 &  x176 &  x245 &  x281 &  x338 &  x464 &  x467 &  x500 &  x520 &  x554 &  x559 &  x560 &  x584 &  x593 &  x637 &  x647 &  x677 &  x690 &  x692 &  x767 &  x769 &  x808 &  x827 &  x1067 &  x1106 &  x1112 & ~x840 & ~x888;
assign c192 =  x20 &  x38 &  x47 &  x86 &  x128 &  x191 &  x197 &  x206 &  x209 &  x233 &  x278 &  x284 &  x365 &  x371 &  x374 &  x383 &  x406 &  x413 &  x415 &  x434 &  x482 &  x632 &  x635 &  x644 &  x667 &  x707 &  x722 &  x746 &  x827 &  x845 &  x866 &  x875 &  x890 &  x938 &  x1018 &  x1043 &  x1049 &  x1070 &  x1091 &  x1118 & ~x273 & ~x321 & ~x477 & ~x654 & ~x732 & ~x733 & ~x771 & ~x915;
assign c194 =  x2 &  x11 &  x14 &  x20 &  x29 &  x35 &  x44 &  x47 &  x50 &  x56 &  x65 &  x68 &  x70 &  x80 &  x83 &  x86 &  x89 &  x101 &  x107 &  x110 &  x113 &  x115 &  x125 &  x134 &  x143 &  x146 &  x154 &  x155 &  x161 &  x164 &  x170 &  x182 &  x185 &  x194 &  x212 &  x233 &  x239 &  x242 &  x260 &  x263 &  x272 &  x278 &  x284 &  x287 &  x290 &  x293 &  x296 &  x302 &  x305 &  x308 &  x314 &  x317 &  x320 &  x326 &  x335 &  x338 &  x341 &  x344 &  x350 &  x353 &  x365 &  x368 &  x371 &  x374 &  x380 &  x383 &  x386 &  x398 &  x401 &  x407 &  x413 &  x416 &  x422 &  x437 &  x440 &  x443 &  x449 &  x461 &  x467 &  x470 &  x473 &  x488 &  x491 &  x494 &  x500 &  x503 &  x511 &  x512 &  x524 &  x527 &  x542 &  x551 &  x557 &  x560 &  x578 &  x581 &  x587 &  x596 &  x620 &  x623 &  x628 &  x629 &  x632 &  x638 &  x641 &  x647 &  x650 &  x653 &  x667 &  x668 &  x689 &  x692 &  x707 &  x715 &  x719 &  x728 &  x731 &  x734 &  x740 &  x748 &  x758 &  x770 &  x773 &  x776 &  x782 &  x787 &  x793 &  x818 &  x824 &  x827 &  x830 &  x832 &  x836 &  x845 &  x848 &  x851 &  x860 &  x863 &  x869 &  x870 &  x871 &  x875 &  x887 &  x890 &  x896 &  x902 &  x908 &  x910 &  x911 &  x920 &  x932 &  x941 &  x944 &  x947 &  x950 &  x953 &  x956 &  x959 &  x974 &  x980 &  x988 &  x995 &  x998 &  x1007 &  x1010 &  x1013 &  x1025 &  x1034 &  x1037 &  x1040 &  x1046 &  x1055 &  x1066 &  x1076 &  x1079 &  x1094 &  x1100 &  x1103 &  x1105 &  x1106 &  x1112 &  x1117 &  x1121 &  x1127 & ~x741;
assign c196 =  x17 &  x77 &  x79 &  x82 &  x83 &  x98 &  x118 &  x182 &  x196 &  x199 &  x206 &  x257 &  x299 &  x316 &  x344 &  x353 &  x394 &  x404 &  x446 &  x488 &  x511 &  x527 &  x530 &  x551 &  x554 &  x578 &  x614 &  x631 &  x635 &  x653 &  x707 &  x722 &  x734 &  x752 &  x815 &  x824 &  x854 &  x922 &  x950 &  x956 &  x980 &  x1034 &  x1067 & ~x186 & ~x291 & ~x303 & ~x546 & ~x585 & ~x663 & ~x858;
assign c198 =  x63 &  x191 &  x239 &  x287 &  x338 &  x362 &  x511 &  x527 &  x545 &  x578 &  x710 &  x731 &  x758 &  x815 &  x818 &  x826 &  x896 &  x922 &  x932 &  x988 &  x1000 &  x1006 &  x1039 &  x1046 &  x1085 &  x1117 &  x1123 &  x1129 & ~x897;
assign c1100 =  x11 &  x23 &  x32 &  x35 &  x56 &  x82 &  x86 &  x110 &  x121 &  x160 &  x199 &  x230 &  x235 &  x245 &  x260 &  x275 &  x277 &  x278 &  x302 &  x311 &  x314 &  x316 &  x322 &  x323 &  x332 &  x335 &  x386 &  x394 &  x413 &  x425 &  x428 &  x443 &  x446 &  x458 &  x464 &  x475 &  x476 &  x491 &  x497 &  x511 &  x527 &  x553 &  x554 &  x566 &  x578 &  x581 &  x592 &  x596 &  x623 &  x656 &  x670 &  x674 &  x692 &  x695 &  x698 &  x701 &  x716 &  x725 &  x770 &  x794 &  x797 &  x799 &  x827 &  x838 &  x866 &  x877 &  x878 &  x893 &  x896 &  x920 &  x935 &  x938 &  x971 &  x994 &  x1019 &  x1079 &  x1085 &  x1106 & ~x186 & ~x663 & ~x702 & ~x741;
assign c1102 =  x2 &  x50 &  x80 &  x110 &  x176 &  x181 &  x254 &  x263 &  x281 &  x335 &  x338 &  x353 &  x364 &  x410 &  x437 &  x440 &  x443 &  x479 &  x491 &  x520 &  x530 &  x553 &  x559 &  x565 &  x571 &  x581 &  x593 &  x596 &  x604 &  x605 &  x614 &  x632 &  x650 &  x676 &  x715 &  x716 &  x809 &  x881 &  x884 &  x929 &  x1004 &  x1043 &  x1049 &  x1055 &  x1061 &  x1097 & ~x705 & ~x1089;
assign c1104 =  x8 &  x32 &  x158 &  x316 &  x355 &  x407 &  x433 &  x474 &  x475 &  x513 &  x553 &  x569 &  x578 &  x587 &  x592 &  x626 &  x655 &  x683 &  x773 &  x851 &  x857 &  x920 &  x1022 &  x1109 & ~x264 & ~x507 & ~x585 & ~x663 & ~x664 & ~x702 & ~x705;
assign c1106 =  x11 &  x23 &  x41 &  x47 &  x68 &  x74 &  x86 &  x89 &  x104 &  x131 &  x143 &  x158 &  x173 &  x212 &  x215 &  x278 &  x284 &  x314 &  x344 &  x359 &  x362 &  x383 &  x395 &  x409 &  x446 &  x452 &  x455 &  x464 &  x473 &  x485 &  x491 &  x554 &  x572 &  x578 &  x590 &  x596 &  x629 &  x650 &  x665 &  x677 &  x695 &  x734 &  x737 &  x758 &  x764 &  x776 &  x815 &  x818 &  x845 &  x848 &  x881 &  x899 &  x929 &  x938 &  x940 &  x1067 &  x1103 &  x1124 & ~x3 & ~x42 & ~x159 & ~x198 & ~x237 & ~x354 & ~x393 & ~x528 & ~x654 & ~x694 & ~x732 & ~x733 & ~x771 & ~x772;
assign c1108 =  x2 &  x14 &  x26 &  x32 &  x53 &  x74 &  x80 &  x86 &  x104 &  x107 &  x121 &  x134 &  x158 &  x160 &  x176 &  x185 &  x188 &  x194 &  x199 &  x200 &  x209 &  x227 &  x236 &  x238 &  x239 &  x272 &  x277 &  x308 &  x311 &  x314 &  x316 &  x317 &  x338 &  x341 &  x365 &  x386 &  x394 &  x422 &  x425 &  x428 &  x443 &  x461 &  x467 &  x473 &  x509 &  x514 &  x527 &  x530 &  x553 &  x554 &  x566 &  x575 &  x578 &  x584 &  x592 &  x596 &  x602 &  x608 &  x617 &  x631 &  x670 &  x671 &  x674 &  x676 &  x677 &  x680 &  x686 &  x710 &  x715 &  x731 &  x734 &  x737 &  x740 &  x746 &  x749 &  x752 &  x764 &  x773 &  x788 &  x791 &  x800 &  x803 &  x809 &  x836 &  x851 &  x863 &  x866 &  x869 &  x887 &  x893 &  x908 &  x911 &  x935 &  x941 &  x950 &  x956 &  x959 &  x971 &  x989 &  x995 &  x1010 &  x1043 &  x1055 &  x1085 &  x1109 &  x1130 & ~x189 & ~x264 & ~x303 & ~x444 & ~x585 & ~x600 & ~x624 & ~x663 & ~x702 & ~x912 & ~x951;
assign c1110 =  x38 &  x50 &  x53 &  x89 &  x137 &  x203 &  x236 &  x266 &  x269 &  x272 &  x308 &  x317 &  x320 &  x323 &  x326 &  x377 &  x383 &  x413 &  x440 &  x460 &  x491 &  x506 &  x521 &  x532 &  x533 &  x572 &  x626 &  x640 &  x641 &  x668 &  x683 &  x692 &  x695 &  x749 &  x767 &  x773 &  x779 &  x785 &  x800 &  x821 &  x842 &  x866 &  x869 &  x893 &  x896 &  x914 &  x917 &  x923 &  x953 &  x956 &  x984 &  x992 &  x998 &  x1024 &  x1055 &  x1063 &  x1118 & ~x273 & ~x390 & ~x471 & ~x1005 & ~x1083;
assign c1112 =  x2 &  x65 &  x107 &  x128 &  x143 &  x227 &  x277 &  x293 &  x299 &  x314 &  x316 &  x317 &  x320 &  x332 &  x347 &  x365 &  x394 &  x413 &  x419 &  x431 &  x527 &  x548 &  x578 &  x629 &  x631 &  x641 &  x709 &  x782 &  x794 &  x811 &  x821 &  x838 &  x844 &  x877 &  x883 &  x908 &  x914 &  x950 &  x956 &  x1055 &  x1091 & ~x309 & ~x349 & ~x387 & ~x388 & ~x426 & ~x444 & ~x663 & ~x702 & ~x741 & ~x858;
assign c1114 =  x11 &  x56 &  x68 &  x152 &  x239 &  x248 &  x272 &  x299 &  x302 &  x320 &  x338 &  x382 &  x407 &  x410 &  x427 &  x449 &  x460 &  x464 &  x482 &  x497 &  x527 &  x565 &  x601 &  x604 &  x640 &  x674 &  x746 &  x784 &  x833 &  x860 &  x866 &  x920 &  x932 &  x939 &  x944 &  x959 &  x978 &  x1017 &  x1096 & ~x390 & ~x432 & ~x471 & ~x510 & ~x954 & ~x993 & ~x1032;
assign c1116 =  x2 &  x11 &  x14 &  x41 &  x47 &  x68 &  x74 &  x80 &  x86 &  x98 &  x131 &  x137 &  x152 &  x164 &  x182 &  x185 &  x188 &  x215 &  x224 &  x248 &  x251 &  x266 &  x299 &  x314 &  x335 &  x338 &  x359 &  x371 &  x392 &  x428 &  x440 &  x443 &  x449 &  x473 &  x512 &  x515 &  x527 &  x554 &  x578 &  x581 &  x596 &  x602 &  x640 &  x662 &  x668 &  x671 &  x674 &  x677 &  x713 &  x719 &  x731 &  x734 &  x749 &  x758 &  x767 &  x773 &  x779 &  x800 &  x824 &  x845 &  x851 &  x857 &  x860 &  x866 &  x890 &  x896 &  x911 &  x920 &  x950 &  x956 &  x968 &  x980 &  x1007 &  x1016 &  x1019 &  x1070 &  x1079 &  x1088 &  x1112 &  x1127 & ~x81 & ~x315 & ~x393 & ~x432 & ~x471 & ~x510 & ~x738 & ~x777 & ~x855 & ~x951 & ~x990 & ~x1029 & ~x1050 & ~x1068 & ~x1107;
assign c1118 =  x2 &  x20 &  x23 &  x41 &  x65 &  x68 &  x74 &  x80 &  x83 &  x86 &  x104 &  x110 &  x113 &  x125 &  x128 &  x131 &  x143 &  x152 &  x164 &  x176 &  x191 &  x227 &  x230 &  x242 &  x245 &  x254 &  x263 &  x275 &  x290 &  x305 &  x311 &  x320 &  x323 &  x326 &  x341 &  x350 &  x356 &  x365 &  x374 &  x383 &  x389 &  x395 &  x407 &  x419 &  x422 &  x428 &  x434 &  x443 &  x445 &  x446 &  x467 &  x470 &  x484 &  x500 &  x503 &  x506 &  x509 &  x533 &  x548 &  x566 &  x575 &  x578 &  x581 &  x584 &  x586 &  x593 &  x596 &  x611 &  x614 &  x623 &  x625 &  x644 &  x656 &  x662 &  x671 &  x683 &  x689 &  x692 &  x695 &  x698 &  x701 &  x707 &  x710 &  x716 &  x725 &  x734 &  x737 &  x749 &  x761 &  x770 &  x784 &  x785 &  x800 &  x818 &  x833 &  x836 &  x839 &  x842 &  x848 &  x851 &  x854 &  x860 &  x862 &  x868 &  x884 &  x901 &  x904 &  x905 &  x907 &  x908 &  x917 &  x920 &  x929 &  x938 &  x940 &  x947 &  x950 &  x956 &  x974 &  x980 &  x992 &  x998 &  x1010 &  x1025 &  x1085 &  x1088 &  x1091 &  x1094 &  x1097 &  x1103 &  x1106 &  x1118 &  x1121 & ~x654 & ~x693 & ~x717 & ~x720 & ~x732 & ~x771 & ~x795 & ~x798 & ~x834 & ~x837 & ~x873 & ~x876;
assign c1120 =  x2 &  x8 &  x17 &  x23 &  x56 &  x58 &  x71 &  x89 &  x113 &  x158 &  x164 &  x188 &  x209 &  x230 &  x236 &  x254 &  x275 &  x281 &  x316 &  x323 &  x326 &  x338 &  x347 &  x365 &  x371 &  x392 &  x413 &  x431 &  x434 &  x437 &  x449 &  x473 &  x482 &  x485 &  x491 &  x494 &  x503 &  x512 &  x553 &  x554 &  x572 &  x584 &  x587 &  x592 &  x593 &  x596 &  x631 &  x635 &  x641 &  x644 &  x659 &  x698 &  x704 &  x716 &  x728 &  x743 &  x752 &  x758 &  x764 &  x776 &  x791 &  x800 &  x803 &  x806 &  x827 &  x848 &  x857 &  x860 &  x893 &  x902 &  x911 &  x932 &  x935 &  x971 &  x992 &  x995 &  x1016 &  x1052 &  x1073 &  x1088 &  x1112 &  x1115 &  x1124 & ~x309 & ~x546 & ~x585 & ~x606 & ~x702 & ~x741 & ~x819 & ~x858 & ~x951 & ~x1029 & ~x1068 & ~x1107;
assign c1122 =  x11 &  x35 &  x62 &  x68 &  x86 &  x119 &  x131 &  x137 &  x152 &  x161 &  x167 &  x209 &  x227 &  x236 &  x254 &  x275 &  x278 &  x284 &  x302 &  x311 &  x323 &  x326 &  x335 &  x359 &  x365 &  x383 &  x395 &  x407 &  x413 &  x434 &  x440 &  x443 &  x467 &  x491 &  x506 &  x509 &  x527 &  x545 &  x551 &  x578 &  x584 &  x596 &  x602 &  x623 &  x625 &  x628 &  x644 &  x647 &  x706 &  x734 &  x745 &  x751 &  x758 &  x767 &  x770 &  x773 &  x784 &  x790 &  x794 &  x797 &  x829 &  x842 &  x851 &  x865 &  x881 &  x890 &  x904 &  x911 &  x920 &  x929 &  x950 &  x956 &  x965 &  x995 &  x1001 &  x1010 &  x1013 &  x1034 &  x1064 & ~x360 & ~x435 & ~x513 & ~x558 & ~x597 & ~x636 & ~x756 & ~x795;
assign c1124 =  x29 &  x50 &  x77 &  x161 &  x227 &  x254 &  x281 &  x296 &  x302 &  x314 &  x320 &  x332 &  x368 &  x386 &  x464 &  x491 &  x494 &  x506 &  x527 &  x584 &  x596 &  x602 &  x668 &  x674 &  x716 &  x785 &  x803 &  x812 &  x848 &  x851 &  x869 &  x901 &  x920 &  x932 &  x956 &  x965 &  x1004 &  x1028 &  x1049 &  x1058 & ~x276 & ~x390 & ~x432 & ~x510 & ~x732 & ~x811 & ~x849 & ~x850 & ~x888 & ~x913 & ~x927 & ~x951 & ~x952 & ~x966 & ~x990 & ~x1005;
assign c1126 =  x2 &  x8 &  x11 &  x14 &  x20 &  x41 &  x68 &  x82 &  x113 &  x125 &  x143 &  x152 &  x160 &  x167 &  x199 &  x200 &  x206 &  x212 &  x224 &  x227 &  x245 &  x248 &  x251 &  x272 &  x277 &  x302 &  x308 &  x314 &  x316 &  x320 &  x322 &  x323 &  x326 &  x335 &  x338 &  x341 &  x347 &  x361 &  x365 &  x371 &  x394 &  x413 &  x440 &  x464 &  x470 &  x473 &  x482 &  x491 &  x503 &  x514 &  x527 &  x536 &  x542 &  x545 &  x548 &  x551 &  x553 &  x569 &  x578 &  x584 &  x592 &  x596 &  x641 &  x659 &  x668 &  x670 &  x692 &  x707 &  x713 &  x716 &  x722 &  x758 &  x761 &  x769 &  x772 &  x773 &  x776 &  x785 &  x788 &  x791 &  x794 &  x800 &  x805 &  x808 &  x827 &  x830 &  x842 &  x845 &  x847 &  x851 &  x866 &  x872 &  x886 &  x893 &  x908 &  x914 &  x923 &  x950 &  x956 &  x989 &  x998 &  x1010 &  x1016 &  x1037 &  x1040 &  x1097 &  x1118 &  x1124 &  x1127 & ~x444 & ~x507 & ~x585 & ~x663 & ~x702 & ~x705;
assign c1128 =  x5 &  x56 &  x86 &  x91 &  x92 &  x98 &  x110 &  x119 &  x130 &  x167 &  x169 &  x197 &  x200 &  x208 &  x221 &  x242 &  x251 &  x257 &  x278 &  x284 &  x290 &  x317 &  x328 &  x332 &  x335 &  x362 &  x367 &  x368 &  x380 &  x422 &  x425 &  x440 &  x443 &  x452 &  x455 &  x470 &  x485 &  x491 &  x524 &  x527 &  x532 &  x545 &  x551 &  x554 &  x571 &  x578 &  x609 &  x610 &  x629 &  x641 &  x649 &  x668 &  x680 &  x683 &  x692 &  x698 &  x701 &  x704 &  x719 &  x731 &  x734 &  x743 &  x745 &  x749 &  x755 &  x800 &  x845 &  x860 &  x905 &  x908 &  x935 &  x941 &  x950 &  x956 &  x959 &  x974 &  x977 &  x1010 &  x1016 &  x1040 &  x1058 &  x1061 &  x1064 &  x1070 &  x1079 & ~x723;
assign c1130 =  x65 &  x80 &  x86 &  x92 &  x119 &  x134 &  x140 &  x164 &  x170 &  x197 &  x203 &  x269 &  x284 &  x302 &  x305 &  x317 &  x335 &  x338 &  x389 &  x443 &  x464 &  x476 &  x493 &  x503 &  x521 &  x527 &  x532 &  x596 &  x644 &  x656 &  x665 &  x670 &  x671 &  x704 &  x710 &  x728 &  x752 &  x755 &  x782 &  x896 &  x911 &  x914 &  x926 &  x932 &  x950 &  x1001 &  x1004 &  x1037 &  x1040 &  x1121 &  x1129 &  x1130 & ~x6 & ~x411 & ~x489 & ~x528 & ~x606 & ~x663 & ~x702 & ~x780 & ~x897 & ~x936 & ~x939;
assign c1132 =  x5 &  x38 &  x86 &  x152 &  x185 &  x200 &  x206 &  x212 &  x227 &  x236 &  x242 &  x278 &  x284 &  x314 &  x320 &  x383 &  x413 &  x437 &  x440 &  x443 &  x467 &  x485 &  x494 &  x506 &  x527 &  x539 &  x548 &  x557 &  x581 &  x596 &  x671 &  x695 &  x710 &  x713 &  x716 &  x740 &  x745 &  x761 &  x767 &  x773 &  x809 &  x851 &  x866 &  x881 &  x883 &  x941 &  x947 &  x950 &  x956 &  x989 &  x1040 &  x1043 &  x1045 &  x1058 &  x1064 &  x1094 &  x1106 &  x1118 & ~x417 & ~x456 & ~x457 & ~x495 & ~x496 & ~x534 & ~x558 & ~x597 & ~x600 & ~x612 & ~x636 & ~x936;
assign c1134 =  x86 &  x113 &  x292 &  x314 &  x370 &  x374 &  x383 &  x409 &  x448 &  x566 &  x641 &  x758 &  x893 &  x902 &  x1016 & ~x801 & ~x879 & ~x918 & ~x951 & ~x952 & ~x957 & ~x991 & ~x996 & ~x1030 & ~x1032 & ~x1068 & ~x1071 & ~x1074 & ~x1107;
assign c1136 =  x119 &  x121 &  x316 &  x320 &  x335 &  x394 &  x449 &  x461 &  x524 &  x592 &  x631 &  x694 &  x721 &  x761 &  x785 &  x788 &  x798 &  x838 &  x883 &  x905 &  x922 &  x1007 &  x1049 &  x1058 &  x1097 & ~x444 & ~x624 & ~x703 & ~x742 & ~x781 & ~x936;
assign c1138 =  x203 &  x277 &  x316 &  x322 &  x553 &  x591 &  x614 &  x677 &  x715 &  x857 & ~x309 & ~x489;
assign c1140 =  x83 &  x119 &  x125 &  x164 &  x220 &  x253 &  x292 &  x298 &  x325 &  x331 &  x337 &  x347 &  x364 &  x376 &  x382 &  x487 &  x506 &  x520 &  x527 &  x545 &  x578 &  x598 &  x637 &  x644 &  x671 &  x695 &  x715 &  x716 &  x734 &  x782 &  x974 &  x1007 &  x1010 &  x1018 & ~x315 & ~x1107;
assign c1142 =  x20 &  x29 &  x32 &  x68 &  x86 &  x224 &  x236 &  x296 &  x317 &  x341 &  x404 &  x443 &  x446 &  x467 &  x472 &  x485 &  x512 &  x527 &  x554 &  x578 &  x595 &  x673 &  x712 &  x728 &  x751 &  x787 &  x803 &  x865 &  x878 &  x896 &  x932 &  x941 &  x950 &  x974 &  x995 &  x1064 &  x1094 &  x1103 & ~x501 & ~x576 & ~x579 & ~x723 & ~x762 & ~x795 & ~x801 & ~x873;
assign c1144 =  x14 &  x20 &  x23 &  x35 &  x44 &  x82 &  x121 &  x160 &  x199 &  x224 &  x266 &  x272 &  x278 &  x293 &  x308 &  x311 &  x316 &  x323 &  x338 &  x341 &  x347 &  x353 &  x416 &  x464 &  x473 &  x475 &  x494 &  x509 &  x513 &  x527 &  x532 &  x542 &  x553 &  x571 &  x578 &  x584 &  x592 &  x623 &  x631 &  x659 &  x662 &  x665 &  x715 &  x725 &  x758 &  x785 &  x845 &  x863 &  x866 &  x890 &  x893 &  x896 &  x941 &  x947 &  x950 &  x956 &  x959 &  x962 &  x1007 &  x1010 &  x1016 & ~x366 & ~x405 & ~x663;
assign c1146 =  x53 &  x68 &  x206 &  x302 &  x374 &  x428 &  x437 &  x491 &  x511 &  x527 &  x550 &  x578 &  x628 &  x671 &  x701 &  x706 &  x728 &  x731 &  x758 &  x776 &  x782 &  x800 &  x818 &  x842 &  x865 &  x890 &  x917 &  x950 &  x1007 &  x1016 &  x1025 & ~x117 & ~x126 & ~x321 & ~x795 & ~x801 & ~x840 & ~x873 & ~x1014 & ~x1074 & ~x1092;
assign c1148 =  x2 &  x14 &  x80 &  x86 &  x212 &  x239 &  x278 &  x302 &  x308 &  x320 &  x389 &  x422 &  x443 &  x491 &  x527 &  x539 &  x542 &  x545 &  x572 &  x578 &  x584 &  x611 &  x667 &  x671 &  x716 &  x734 &  x745 &  x746 &  x752 &  x758 &  x767 &  x784 &  x794 &  x812 &  x845 &  x851 &  x860 &  x864 &  x865 &  x866 &  x903 &  x904 &  x908 &  x914 &  x941 &  x950 &  x956 &  x965 &  x977 &  x1010 &  x1021 & ~x321 & ~x621 & ~x756 & ~x801 & ~x834 & ~x840 & ~x918;
assign c1150 =  x14 &  x38 &  x47 &  x65 &  x71 &  x92 &  x104 &  x119 &  x134 &  x143 &  x167 &  x199 &  x254 &  x313 &  x316 &  x389 &  x410 &  x475 &  x491 &  x511 &  x515 &  x539 &  x545 &  x553 &  x556 &  x581 &  x584 &  x595 &  x596 &  x629 &  x631 &  x665 &  x674 &  x680 &  x686 &  x689 &  x716 &  x719 &  x725 &  x830 &  x896 &  x914 &  x920 &  x947 &  x950 &  x956 &  x959 &  x962 &  x971 &  x995 &  x1109 & ~x45 & ~x84 & ~x303 & ~x702;
assign c1152 =  x53 &  x74 &  x119 &  x131 &  x254 &  x278 &  x311 &  x316 &  x350 &  x383 &  x392 &  x428 &  x440 &  x443 &  x596 &  x631 &  x677 &  x701 &  x749 &  x776 &  x785 &  x803 &  x851 &  x890 &  x896 &  x938 &  x974 &  x1016 &  x1043 & ~x381 & ~x388 & ~x459 & ~x702 & ~x780 & ~x795 & ~x1101;
assign c1154 =  x11 &  x65 &  x86 &  x164 &  x302 &  x335 &  x410 &  x437 &  x475 &  x476 &  x500 &  x527 &  x553 &  x596 &  x631 &  x644 &  x668 &  x688 &  x709 &  x722 &  x725 &  x728 &  x766 &  x772 &  x773 &  x785 &  x800 &  x838 &  x844 &  x866 &  x883 &  x899 &  x920 &  x932 &  x953 &  x968 &  x989 &  x992 &  x1016 &  x1028 &  x1040 & ~x45 & ~x168 & ~x426 & ~x705 & ~x822;
assign c1156 =  x2 &  x56 &  x68 &  x122 &  x164 &  x185 &  x200 &  x215 &  x218 &  x224 &  x227 &  x254 &  x263 &  x389 &  x392 &  x401 &  x443 &  x485 &  x491 &  x506 &  x527 &  x578 &  x611 &  x614 &  x662 &  x680 &  x713 &  x716 &  x725 &  x731 &  x752 &  x797 &  x800 &  x842 &  x848 &  x851 &  x866 &  x896 &  x908 &  x920 &  x950 &  x956 &  x965 &  x1007 &  x1085 &  x1088 &  x1100 & ~x87 & ~x165 & ~x204 & ~x243 & ~x321 & ~x399 & ~x645 & ~x684 & ~x723 & ~x732 & ~x840 & ~x879 & ~x918 & ~x951 & ~x957 & ~x990 & ~x996 & ~x1029 & ~x1035 & ~x1068 & ~x1074 & ~x1107;
assign c1158 =  x38 &  x41 &  x44 &  x101 &  x197 &  x263 &  x311 &  x413 &  x416 &  x443 &  x454 &  x482 &  x532 &  x553 &  x559 &  x569 &  x578 &  x598 &  x631 &  x637 &  x648 &  x649 &  x674 &  x676 &  x746 &  x769 &  x808 &  x832 &  x845 &  x854 &  x881 &  x902 &  x908 &  x974 &  x998 & ~x723;
assign c1160 =  x38 &  x86 &  x116 &  x142 &  x146 &  x152 &  x259 &  x308 &  x335 &  x359 &  x437 &  x445 &  x473 &  x476 &  x484 &  x506 &  x542 &  x578 &  x584 &  x617 &  x641 &  x644 &  x662 &  x665 &  x674 &  x707 &  x773 &  x791 &  x851 &  x911 &  x959 &  x989 &  x1016 &  x1022 &  x1117 & ~x6 & ~x45 & ~x84 & ~x123 & ~x162 & ~x201 & ~x240 & ~x315 & ~x513 & ~x630 & ~x669;
assign c1162 =  x8 &  x11 &  x74 &  x89 &  x113 &  x152 &  x191 &  x206 &  x224 &  x239 &  x257 &  x269 &  x296 &  x359 &  x371 &  x407 &  x416 &  x485 &  x494 &  x497 &  x500 &  x506 &  x515 &  x518 &  x524 &  x527 &  x545 &  x578 &  x611 &  x623 &  x638 &  x641 &  x665 &  x667 &  x698 &  x706 &  x740 &  x745 &  x749 &  x784 &  x845 &  x869 &  x875 &  x905 &  x908 &  x911 &  x935 &  x947 &  x959 &  x965 &  x989 &  x1010 &  x1058 &  x1064 & ~x87 & ~x126 & ~x165 & ~x321 & ~x360 & ~x384 & ~x399 & ~x423 & ~x528 & ~x840 & ~x879 & ~x912 & ~x918 & ~x951 & ~x990 & ~x996 & ~x1029 & ~x1035 & ~x1068 & ~x1107;
assign c1164 =  x38 &  x73 &  x92 &  x106 &  x173 &  x200 &  x210 &  x227 &  x236 &  x249 &  x250 &  x293 &  x302 &  x316 &  x386 &  x389 &  x455 &  x488 &  x512 &  x524 &  x545 &  x592 &  x617 &  x620 &  x631 &  x686 &  x701 &  x740 &  x826 &  x865 &  x908;
assign c1166 =  x17 &  x41 &  x53 &  x113 &  x164 &  x185 &  x200 &  x203 &  x218 &  x224 &  x242 &  x251 &  x254 &  x350 &  x365 &  x371 &  x437 &  x488 &  x533 &  x623 &  x671 &  x692 &  x713 &  x728 &  x761 &  x773 &  x782 &  x784 &  x812 &  x890 &  x902 &  x905 &  x923 &  x940 &  x941 &  x1016 &  x1031 &  x1040 & ~x393 & ~x528 & ~x576 & ~x616 & ~x655 & ~x694 & ~x732 & ~x733 & ~x772 & ~x795 & ~x957;
assign c1168 =  x5 &  x22 &  x61 &  x106 &  x139 &  x263 &  x268 &  x302 &  x320 &  x328 &  x586 &  x680 &  x737 &  x829 &  x868 &  x881 &  x889 &  x899 &  x950 &  x1016 & ~x6 & ~x45 & ~x84 & ~x681;
assign c1170 =  x11 &  x47 &  x68 &  x131 &  x185 &  x197 &  x200 &  x203 &  x218 &  x227 &  x232 &  x242 &  x271 &  x293 &  x302 &  x308 &  x311 &  x317 &  x335 &  x383 &  x455 &  x521 &  x575 &  x584 &  x593 &  x644 &  x656 &  x668 &  x683 &  x692 &  x731 &  x734 &  x737 &  x794 &  x812 &  x829 &  x851 &  x866 &  x868 &  x907 &  x923 &  x938 &  x946 &  x953 &  x959 &  x995 &  x998 &  x1022 &  x1070 & ~x234 & ~x654 & ~x694 & ~x733 & ~x771 & ~x772 & ~x795 & ~x873 & ~x912 & ~x918 & ~x951;
assign c1172 =  x47 &  x53 &  x86 &  x197 &  x203 &  x224 &  x227 &  x275 &  x302 &  x311 &  x314 &  x329 &  x335 &  x353 &  x356 &  x383 &  x389 &  x416 &  x437 &  x443 &  x485 &  x488 &  x511 &  x539 &  x545 &  x554 &  x581 &  x605 &  x668 &  x671 &  x698 &  x713 &  x716 &  x731 &  x734 &  x737 &  x758 &  x761 &  x766 &  x773 &  x805 &  x844 &  x845 &  x851 &  x881 &  x896 &  x905 &  x908 &  x947 &  x950 &  x953 &  x956 &  x977 &  x989 &  x1007 &  x1010 &  x1016 &  x1064 &  x1076 &  x1097 &  x1115 & ~x372 & ~x450 & ~x451 & ~x456 & ~x489 & ~x495 & ~x528 & ~x612 & ~x651 & ~x780;
assign c1174 =  x23 &  x38 &  x74 &  x80 &  x142 &  x164 &  x197 &  x224 &  x242 &  x323 &  x335 &  x389 &  x422 &  x449 &  x472 &  x494 &  x511 &  x512 &  x527 &  x533 &  x550 &  x551 &  x590 &  x628 &  x673 &  x686 &  x695 &  x701 &  x712 &  x713 &  x737 &  x803 &  x809 &  x832 &  x839 &  x860 &  x871 &  x875 &  x887 &  x910 &  x917 &  x950 &  x1000 &  x1019 &  x1039 &  x1051 &  x1090 &  x1117 &  x1130 & ~x723 & ~x762 & ~x801;
assign c1176 =  x332 &  x382 &  x415 &  x532 &  x538 &  x559 &  x565 &  x572 &  x598 &  x604 &  x623 &  x640 &  x686 &  x752 &  x773 &  x896 &  x938 &  x950 &  x1096 & ~x351 & ~x432 & ~x471 & ~x510 & ~x888 & ~x927 & ~x1032;
assign c1178 =  x65 &  x316 &  x347 &  x511 &  x578 &  x687 &  x1000 &  x1007 &  x1051 & ~x48 & ~x600 & ~x723;
assign c1180 =  x41 &  x62 &  x119 &  x122 &  x152 &  x176 &  x191 &  x197 &  x209 &  x236 &  x242 &  x257 &  x275 &  x284 &  x302 &  x305 &  x341 &  x350 &  x356 &  x389 &  x392 &  x413 &  x422 &  x428 &  x443 &  x491 &  x494 &  x500 &  x509 &  x527 &  x539 &  x542 &  x554 &  x572 &  x584 &  x596 &  x599 &  x623 &  x641 &  x665 &  x668 &  x692 &  x695 &  x716 &  x719 &  x734 &  x749 &  x758 &  x761 &  x785 &  x800 &  x803 &  x851 &  x890 &  x908 &  x923 &  x950 &  x980 &  x989 &  x1031 &  x1064 &  x1088 & ~x141 & ~x180 & ~x198 & ~x276 & ~x315 & ~x399 & ~x513 & ~x654 & ~x954 & ~x1065 & ~x1104 & ~x1116;
assign c1182 =  x116 &  x239 &  x245 &  x254 &  x284 &  x311 &  x335 &  x338 &  x377 &  x394 &  x416 &  x511 &  x536 &  x554 &  x578 &  x605 &  x669 &  x670 &  x671 &  x673 &  x708 &  x709 &  x712 &  x716 &  x722 &  x725 &  x743 &  x746 &  x787 &  x800 &  x815 &  x836 &  x860 &  x883 &  x890 &  x899 &  x922 &  x929 &  x994 &  x1016 &  x1031 &  x1129 & ~x606 & ~x663 & ~x1092;
assign c1184 =  x40 &  x56 &  x65 &  x79 &  x86 &  x89 &  x104 &  x107 &  x146 &  x164 &  x235 &  x242 &  x266 &  x284 &  x313 &  x368 &  x377 &  x422 &  x482 &  x506 &  x545 &  x575 &  x578 &  x604 &  x605 &  x614 &  x617 &  x671 &  x674 &  x686 &  x743 &  x797 &  x818 &  x824 &  x830 &  x860 &  x881 &  x917 &  x938 &  x1016 &  x1061 &  x1064 &  x1109 & ~x6 & ~x45 & ~x46 & ~x84 & ~x123 & ~x705 & ~x792;
assign c1186 =  x38 &  x173 &  x185 &  x269 &  x277 &  x311 &  x317 &  x353 &  x362 &  x377 &  x461 &  x497 &  x509 &  x545 &  x599 &  x641 &  x653 &  x680 &  x700 &  x791 &  x797 &  x845 &  x914 &  x965 &  x983 &  x1001 &  x1022 &  x1043 &  x1076 &  x1109 &  x1124 & ~x420 & ~x756 & ~x1014 & ~x1024 & ~x1029;
assign c1188 =  x305 &  x485 &  x494 &  x542 &  x680 &  x784 &  x995 & ~x87 & ~x165 & ~x432 & ~x477 & ~x654 & ~x771 & ~x951 & ~x952 & ~x954 & ~x990 & ~x993 & ~x1029 & ~x1032 & ~x1068 & ~x1071;
assign c1190 =  x35 &  x53 &  x59 &  x74 &  x86 &  x121 &  x158 &  x160 &  x164 &  x191 &  x199 &  x224 &  x236 &  x238 &  x257 &  x272 &  x278 &  x316 &  x341 &  x350 &  x394 &  x413 &  x416 &  x433 &  x440 &  x443 &  x452 &  x455 &  x475 &  x497 &  x509 &  x513 &  x514 &  x542 &  x551 &  x553 &  x575 &  x592 &  x611 &  x617 &  x631 &  x641 &  x671 &  x676 &  x709 &  x715 &  x716 &  x728 &  x740 &  x746 &  x748 &  x749 &  x785 &  x787 &  x806 &  x809 &  x824 &  x833 &  x848 &  x911 &  x920 &  x926 &  x956 &  x1007 &  x1025 &  x1037 &  x1040 &  x1061 &  x1070 &  x1091 &  x1094 &  x1109 & ~x153 & ~x231 & ~x366 & ~x444 & ~x663 & ~x702;
assign c1192 =  x29 &  x68 &  x86 &  x115 &  x154 &  x164 &  x181 &  x218 &  x224 &  x253 &  x259 &  x292 &  x298 &  x304 &  x310 &  x317 &  x320 &  x335 &  x413 &  x437 &  x443 &  x445 &  x479 &  x484 &  x488 &  x542 &  x545 &  x596 &  x638 &  x668 &  x671 &  x728 &  x749 &  x773 &  x866 &  x905 &  x950 &  x956 &  x965 &  x974 &  x1007 &  x1010 &  x1076 &  x1085 & ~x81 & ~x120 & ~x315 & ~x474 & ~x480 & ~x513;
assign c1194 =  x116 &  x142 &  x181 &  x239 &  x278 &  x409 &  x448 &  x487 &  x526 &  x565 &  x578 &  x643 &  x677 &  x680 &  x716 &  x896 &  x1010 & ~x618 & ~x657 & ~x696 & ~x697 & ~x762 & ~x813;
assign c1196 =  x14 &  x47 &  x74 &  x95 &  x110 &  x176 &  x212 &  x251 &  x254 &  x269 &  x284 &  x365 &  x425 &  x428 &  x458 &  x524 &  x545 &  x548 &  x554 &  x572 &  x581 &  x677 &  x692 &  x731 &  x770 &  x812 &  x815 &  x827 &  x845 &  x859 &  x881 &  x896 &  x902 &  x905 &  x914 &  x950 &  x959 &  x985 &  x1001 &  x1007 &  x1013 &  x1018 &  x1024 &  x1040 &  x1058 &  x1063 &  x1088 &  x1096 & ~x660 & ~x699 & ~x700 & ~x723 & ~x738 & ~x954;
assign c1198 =  x1 &  x8 &  x40 &  x50 &  x79 &  x215 &  x227 &  x235 &  x287 &  x311 &  x335 &  x368 &  x374 &  x446 &  x452 &  x506 &  x515 &  x518 &  x545 &  x557 &  x563 &  x578 &  x590 &  x599 &  x605 &  x608 &  x632 &  x635 &  x650 &  x701 &  x791 &  x794 &  x830 &  x842 &  x884 &  x890 &  x917 &  x932 &  x962 &  x1001 &  x1007 &  x1112 & ~x114 & ~x141 & ~x162 & ~x180 & ~x207 & ~x213 & ~x246 & ~x432 & ~x471 & ~x510 & ~x588 & ~x627 & ~x705 & ~x1005 & ~x1032 & ~x1065 & ~x1071 & ~x1104;
assign c1200 =  x38 &  x47 &  x50 &  x86 &  x121 &  x160 &  x188 &  x199 &  x218 &  x224 &  x235 &  x277 &  x302 &  x316 &  x322 &  x353 &  x383 &  x394 &  x410 &  x518 &  x527 &  x578 &  x584 &  x635 &  x773 &  x785 &  x799 &  x836 &  x844 &  x881 &  x883 &  x887 &  x889 &  x922 &  x950 &  x961 &  x968 &  x974 &  x1000 &  x1010 & ~x153 & ~x486 & ~x702;
assign c1202 =  x56 &  x68 &  x83 &  x86 &  x92 &  x104 &  x140 &  x188 &  x203 &  x215 &  x218 &  x227 &  x239 &  x302 &  x316 &  x317 &  x350 &  x365 &  x368 &  x371 &  x374 &  x383 &  x389 &  x443 &  x473 &  x488 &  x497 &  x542 &  x548 &  x553 &  x560 &  x563 &  x575 &  x578 &  x592 &  x631 &  x641 &  x665 &  x677 &  x709 &  x740 &  x748 &  x749 &  x755 &  x767 &  x776 &  x787 &  x818 &  x857 &  x877 &  x878 &  x887 &  x920 &  x935 &  x938 &  x956 &  x980 &  x986 &  x995 &  x1007 &  x1010 &  x1037 &  x1052 &  x1094 &  x1118 & ~x342 & ~x420 & ~x459 & ~x460 & ~x498 & ~x663 & ~x702 & ~x951;
assign c1204 =  x8 &  x11 &  x23 &  x143 &  x158 &  x164 &  x200 &  x224 &  x233 &  x266 &  x269 &  x278 &  x308 &  x314 &  x353 &  x382 &  x383 &  x389 &  x398 &  x415 &  x440 &  x443 &  x464 &  x527 &  x563 &  x617 &  x640 &  x791 &  x812 &  x859 &  x863 &  x896 &  x908 &  x911 &  x932 &  x937 &  x940 &  x950 &  x953 &  x956 &  x965 &  x974 &  x1004 &  x1013 &  x1015 &  x1031 &  x1056 &  x1079 &  x1093 &  x1096 & ~x432 & ~x468 & ~x471 & ~x507 & ~x510 & ~x588 & ~x627 & ~x1032 & ~x1071 & ~x1110;
assign c1206 =  x1 &  x26 &  x172 &  x178 &  x181 &  x253 &  x340 &  x409 &  x484 &  x487 &  x578 &  x781 &  x907 &  x941 &  x985 & ~x315 & ~x660;
assign c1208 =  x2 &  x14 &  x32 &  x41 &  x94 &  x135 &  x136 &  x215 &  x218 &  x236 &  x278 &  x284 &  x302 &  x311 &  x433 &  x443 &  x592 &  x596 &  x611 &  x641 &  x709 &  x713 &  x715 &  x728 &  x734 &  x787 &  x800 &  x827 &  x842 &  x851 &  x881 &  x950 &  x1007 &  x1058 &  x1079 &  x1115 & ~x585 & ~x624 & ~x663 & ~x702 & ~x741;
assign c1210 =  x35 &  x41 &  x68 &  x86 &  x152 &  x181 &  x230 &  x259 &  x298 &  x317 &  x335 &  x338 &  x353 &  x356 &  x377 &  x409 &  x428 &  x437 &  x446 &  x448 &  x455 &  x470 &  x487 &  x524 &  x525 &  x526 &  x527 &  x539 &  x542 &  x554 &  x565 &  x578 &  x584 &  x593 &  x596 &  x605 &  x623 &  x641 &  x665 &  x671 &  x713 &  x728 &  x767 &  x773 &  x818 &  x860 &  x861 &  x866 &  x881 &  x900 &  x901 &  x908 &  x914 &  x920 &  x923 &  x938 &  x939 &  x968 &  x974 &  x995 &  x1016 &  x1018 &  x1037 &  x1043 &  x1055 &  x1097 &  x1106 & ~x117 & ~x189 & ~x274 & ~x276 & ~x313 & ~x351;
assign c1212 =  x29 &  x37 &  x50 &  x52 &  x74 &  x76 &  x91 &  x103 &  x115 &  x142 &  x154 &  x181 &  x248 &  x284 &  x317 &  x353 &  x365 &  x419 &  x422 &  x443 &  x485 &  x497 &  x506 &  x527 &  x551 &  x569 &  x578 &  x589 &  x628 &  x641 &  x653 &  x659 &  x668 &  x725 &  x731 &  x737 &  x803 &  x821 &  x866 &  x869 &  x883 &  x920 &  x956 &  x965 &  x992 &  x1028 &  x1088 &  x1090 &  x1117 &  x1127 &  x1130 & ~x951 & ~x996 & ~x1029;
assign c1214 =  x16 &  x35 &  x47 &  x56 &  x83 &  x113 &  x119 &  x172 &  x211 &  x254 &  x257 &  x296 &  x299 &  x304 &  x328 &  x338 &  x344 &  x353 &  x365 &  x367 &  x374 &  x406 &  x415 &  x445 &  x448 &  x484 &  x494 &  x509 &  x512 &  x523 &  x530 &  x554 &  x562 &  x565 &  x640 &  x641 &  x665 &  x671 &  x707 &  x716 &  x800 &  x851 &  x890 &  x905 &  x935 &  x956 &  x976 &  x1064 &  x1094 &  x1102 & ~x276 & ~x432 & ~x471 & ~x549 & ~x588 & ~x1032 & ~x1071 & ~x1110;
assign c1216 =  x1 &  x22 &  x38 &  x41 &  x53 &  x61 &  x128 &  x139 &  x145 &  x172 &  x178 &  x197 &  x205 &  x218 &  x227 &  x250 &  x256 &  x257 &  x263 &  x328 &  x335 &  x356 &  x365 &  x366 &  x367 &  x406 &  x422 &  x443 &  x445 &  x473 &  x484 &  x527 &  x551 &  x572 &  x578 &  x596 &  x608 &  x617 &  x689 &  x716 &  x719 &  x728 &  x734 &  x749 &  x752 &  x758 &  x767 &  x773 &  x827 &  x829 &  x860 &  x866 &  x884 &  x890 &  x944 &  x950 &  x953 &  x956 &  x965 &  x983 &  x1016 &  x1022 &  x1058 &  x1079 &  x1121 & ~x753;
assign c1218 =  x32 &  x35 &  x38 &  x68 &  x86 &  x89 &  x95 &  x113 &  x125 &  x179 &  x182 &  x191 &  x206 &  x214 &  x215 &  x218 &  x253 &  x272 &  x302 &  x304 &  x305 &  x314 &  x332 &  x335 &  x353 &  x356 &  x365 &  x383 &  x407 &  x413 &  x443 &  x488 &  x491 &  x494 &  x527 &  x536 &  x557 &  x575 &  x605 &  x614 &  x625 &  x644 &  x668 &  x695 &  x698 &  x713 &  x731 &  x737 &  x752 &  x758 &  x761 &  x764 &  x800 &  x851 &  x854 &  x878 &  x881 &  x950 &  x956 &  x959 &  x962 &  x965 &  x989 &  x1007 &  x1022 &  x1028 &  x1040 &  x1049 &  x1058 &  x1082 &  x1088 &  x1097 & ~x81 & ~x120 & ~x237 & ~x276 & ~x315 & ~x504 & ~x513 & ~x543 & ~x582 & ~x621 & ~x660 & ~x699 & ~x738;
assign c1220 =  x68 &  x80 &  x86 &  x119 &  x125 &  x161 &  x191 &  x224 &  x293 &  x314 &  x317 &  x320 &  x326 &  x335 &  x347 &  x355 &  x356 &  x365 &  x380 &  x383 &  x394 &  x437 &  x443 &  x491 &  x506 &  x511 &  x551 &  x575 &  x578 &  x581 &  x593 &  x623 &  x668 &  x671 &  x680 &  x716 &  x725 &  x728 &  x734 &  x737 &  x743 &  x748 &  x749 &  x761 &  x770 &  x787 &  x833 &  x860 &  x905 &  x908 &  x935 &  x941 &  x1007 &  x1016 &  x1058 &  x1064 &  x1079 &  x1091 &  x1112 & ~x420 & ~x459 & ~x460 & ~x498 & ~x501 & ~x537 & ~x618 & ~x657 & ~x702 & ~x741 & ~x951 & ~x990;
assign c1222 =  x1 &  x8 &  x11 &  x17 &  x20 &  x32 &  x35 &  x40 &  x53 &  x65 &  x74 &  x83 &  x128 &  x131 &  x140 &  x149 &  x152 &  x167 &  x173 &  x194 &  x200 &  x209 &  x212 &  x253 &  x254 &  x269 &  x281 &  x296 &  x304 &  x317 &  x326 &  x335 &  x338 &  x365 &  x367 &  x383 &  x386 &  x392 &  x413 &  x425 &  x428 &  x431 &  x440 &  x452 &  x458 &  x485 &  x494 &  x521 &  x533 &  x539 &  x578 &  x581 &  x587 &  x611 &  x617 &  x623 &  x635 &  x638 &  x641 &  x647 &  x650 &  x659 &  x665 &  x668 &  x677 &  x698 &  x706 &  x716 &  x740 &  x745 &  x752 &  x764 &  x767 &  x773 &  x782 &  x784 &  x806 &  x815 &  x824 &  x833 &  x845 &  x866 &  x884 &  x890 &  x947 &  x968 &  x974 &  x983 &  x998 &  x1010 &  x1016 &  x1019 &  x1025 &  x1076 &  x1079 &  x1085 &  x1115 &  x1121 & ~x360 & ~x474 & ~x513 & ~x720 & ~x738 & ~x759;
assign c1224 =  x236 &  x277 &  x473 &  x556 &  x592 &  x595 &  x631 &  x676 &  x680 &  x778 &  x1051 &  x1129 & ~x309 & ~x486 & ~x585 & ~x663;
assign c1226 =  x26 &  x41 &  x110 &  x119 &  x173 &  x188 &  x200 &  x203 &  x220 &  x254 &  x259 &  x272 &  x293 &  x298 &  x308 &  x337 &  x353 &  x365 &  x389 &  x416 &  x443 &  x476 &  x479 &  x506 &  x509 &  x527 &  x551 &  x563 &  x575 &  x578 &  x634 &  x668 &  x671 &  x673 &  x692 &  x707 &  x710 &  x712 &  x728 &  x749 &  x751 &  x767 &  x770 &  x785 &  x787 &  x790 &  x815 &  x832 &  x845 &  x890 &  x905 &  x917 &  x941 &  x977 &  x988 &  x1040 &  x1079 &  x1103 & ~x567 & ~x606 & ~x684 & ~x723;
assign c1228 =  x35 &  x68 &  x278 &  x353 &  x383 &  x413 &  x428 &  x437 &  x448 &  x455 &  x559 &  x601 &  x728 &  x734 &  x758 &  x806 &  x896 &  x920 &  x938 &  x980 &  x1056 &  x1064 & ~x849 & ~x888 & ~x927 & ~x951 & ~x966 & ~x1005 & ~x1029 & ~x1068;
assign c1230 =  x11 &  x38 &  x82 &  x119 &  x152 &  x188 &  x199 &  x224 &  x277 &  x316 &  x394 &  x404 &  x491 &  x506 &  x551 &  x592 &  x596 &  x616 &  x644 &  x686 &  x716 &  x769 &  x778 &  x785 &  x808 &  x877 &  x889 &  x922 &  x956 &  x1043 &  x1051 &  x1090 &  x1123 &  x1129 & ~x303 & ~x546 & ~x585 & ~x741;
assign c1232 =  x40 &  x79 &  x245 &  x305 &  x362 &  x527 &  x551 &  x634 &  x674 &  x706 &  x745 &  x767 &  x829 &  x898 &  x985 &  x1024 &  x1063 &  x1102 & ~x660 & ~x699 & ~x738 & ~x954;
assign c1234 =  x20 &  x29 &  x47 &  x53 &  x74 &  x86 &  x104 &  x107 &  x122 &  x197 &  x200 &  x227 &  x230 &  x233 &  x239 &  x275 &  x278 &  x281 &  x293 &  x311 &  x314 &  x317 &  x335 &  x338 &  x344 &  x347 &  x350 &  x356 &  x365 &  x371 &  x374 &  x407 &  x410 &  x413 &  x416 &  x428 &  x443 &  x452 &  x473 &  x491 &  x503 &  x509 &  x515 &  x518 &  x527 &  x548 &  x572 &  x578 &  x581 &  x602 &  x605 &  x611 &  x625 &  x641 &  x647 &  x656 &  x695 &  x704 &  x706 &  x710 &  x716 &  x728 &  x734 &  x745 &  x752 &  x755 &  x758 &  x764 &  x781 &  x782 &  x785 &  x818 &  x830 &  x833 &  x842 &  x862 &  x866 &  x872 &  x875 &  x896 &  x905 &  x908 &  x917 &  x920 &  x929 &  x935 &  x950 &  x956 &  x974 &  x1010 &  x1016 &  x1022 &  x1025 &  x1040 &  x1052 &  x1055 &  x1082 &  x1088 &  x1106 & ~x237 & ~x276 & ~x315 & ~x321 & ~x360 & ~x399 & ~x438 & ~x591 & ~x630 & ~x660 & ~x669 & ~x699 & ~x738 & ~x792;
assign c1236 =  x26 &  x29 &  x143 &  x203 &  x242 &  x248 &  x257 &  x301 &  x325 &  x340 &  x364 &  x446 &  x449 &  x520 &  x559 &  x563 &  x578 &  x584 &  x590 &  x623 &  x632 &  x637 &  x674 &  x676 &  x689 &  x715 &  x728 &  x734 &  x785 &  x787 &  x832 &  x845 &  x866 &  x884 &  x910 &  x917 &  x949 &  x950 &  x1010 &  x1052 &  x1070 &  x1124 & ~x528 & ~x657 & ~x696;
assign c1238 =  x74 &  x80 &  x89 &  x131 &  x167 &  x221 &  x278 &  x281 &  x284 &  x305 &  x422 &  x443 &  x445 &  x452 &  x473 &  x484 &  x503 &  x509 &  x548 &  x560 &  x578 &  x584 &  x665 &  x668 &  x674 &  x701 &  x704 &  x706 &  x707 &  x731 &  x734 &  x749 &  x755 &  x785 &  x791 &  x815 &  x827 &  x833 &  x851 &  x901 &  x908 &  x974 &  x980 &  x989 &  x995 &  x1040 &  x1043 &  x1046 &  x1070 &  x1079 &  x1088 &  x1094 & ~x87 & ~x126 & ~x390 & ~x438 & ~x477 & ~x555 & ~x738 & ~x954 & ~x990 & ~x993 & ~x1029;
assign c1240 =  x17 &  x20 &  x68 &  x86 &  x113 &  x119 &  x122 &  x128 &  x137 &  x173 &  x194 &  x242 &  x254 &  x320 &  x332 &  x335 &  x341 &  x383 &  x389 &  x472 &  x491 &  x503 &  x511 &  x527 &  x548 &  x550 &  x578 &  x587 &  x671 &  x683 &  x689 &  x695 &  x716 &  x743 &  x758 &  x818 &  x842 &  x851 &  x863 &  x887 &  x893 &  x917 &  x950 &  x956 &  x959 &  x974 &  x989 &  x1019 &  x1037 &  x1064 &  x1067 &  x1076 &  x1118 &  x1127 & ~x240 & ~x357 & ~x459 & ~x474 & ~x498 & ~x537 & ~x576 & ~x678 & ~x897 & ~x936 & ~x957 & ~x990 & ~x1029 & ~x1035 & ~x1068;
assign c1242 =  x2 &  x17 &  x56 &  x71 &  x89 &  x104 &  x107 &  x182 &  x200 &  x206 &  x221 &  x224 &  x239 &  x242 &  x254 &  x287 &  x293 &  x323 &  x338 &  x371 &  x374 &  x380 &  x401 &  x407 &  x419 &  x425 &  x428 &  x437 &  x443 &  x461 &  x467 &  x473 &  x485 &  x488 &  x494 &  x509 &  x512 &  x530 &  x542 &  x545 &  x551 &  x557 &  x563 &  x572 &  x575 &  x581 &  x584 &  x593 &  x599 &  x611 &  x617 &  x623 &  x638 &  x641 &  x653 &  x656 &  x671 &  x680 &  x692 &  x695 &  x698 &  x710 &  x716 &  x755 &  x758 &  x784 &  x791 &  x803 &  x809 &  x824 &  x827 &  x842 &  x851 &  x884 &  x902 &  x908 &  x938 &  x940 &  x946 &  x953 &  x956 &  x980 &  x985 &  x998 &  x1004 &  x1007 &  x1016 &  x1024 &  x1031 &  x1040 &  x1043 &  x1055 &  x1063 &  x1085 &  x1088 &  x1091 &  x1094 & ~x432 & ~x471 & ~x510 & ~x654 & ~x732 & ~x733 & ~x772 & ~x811 & ~x849 & ~x888 & ~x912 & ~x915 & ~x951;
assign c1244 =  x143 &  x146 &  x152 &  x191 &  x239 &  x254 &  x271 &  x293 &  x335 &  x359 &  x374 &  x443 &  x536 &  x572 &  x584 &  x644 &  x706 &  x767 &  x785 &  x881 &  x908 &  x944 &  x1004 &  x1016 &  x1018 &  x1058 & ~x87 & ~x126 & ~x165 & ~x321 & ~x351 & ~x477 & ~x594 & ~x912 & ~x951 & ~x990 & ~x1029 & ~x1068;
assign c1246 =  x14 &  x38 &  x91 &  x131 &  x154 &  x173 &  x181 &  x220 &  x227 &  x284 &  x293 &  x296 &  x317 &  x335 &  x344 &  x353 &  x383 &  x395 &  x422 &  x440 &  x443 &  x488 &  x506 &  x518 &  x545 &  x653 &  x656 &  x698 &  x701 &  x716 &  x728 &  x734 &  x749 &  x758 &  x767 &  x827 &  x863 &  x865 &  x887 &  x908 &  x950 &  x953 &  x956 &  x992 &  x1097 &  x1123 &  x1127 & ~x81 & ~x276 & ~x315 & ~x528 & ~x912 & ~x918 & ~x951;
assign c1248 =  x137 &  x185 &  x224 &  x323 &  x359 &  x415 &  x437 &  x503 &  x527 &  x596 &  x626 &  x674 &  x722 &  x743 &  x752 &  x866 &  x890 &  x896 &  x910 &  x953 &  x959 &  x988 &  x1000 &  x1039 &  x1045 &  x1097 &  x1123 & ~x450 & ~x490 & ~x528 & ~x567 & ~x606 & ~x834;
assign c1250 =  x8 &  x56 &  x131 &  x146 &  x152 &  x200 &  x209 &  x215 &  x224 &  x236 &  x251 &  x290 &  x317 &  x368 &  x371 &  x419 &  x422 &  x527 &  x545 &  x581 &  x604 &  x641 &  x671 &  x683 &  x707 &  x758 &  x848 &  x860 &  x861 &  x881 &  x884 &  x896 &  x900 &  x905 &  x923 &  x940 &  x947 &  x953 &  x956 &  x974 &  x992 &  x1007 &  x1010 &  x1055 &  x1058 &  x1085 &  x1094 & ~x852 & ~x855 & ~x894 & ~x912 & ~x934 & ~x951 & ~x990;
assign c1252 =  x2 &  x11 &  x14 &  x38 &  x59 &  x68 &  x83 &  x104 &  x146 &  x185 &  x197 &  x200 &  x227 &  x236 &  x239 &  x254 &  x278 &  x293 &  x302 &  x314 &  x350 &  x365 &  x389 &  x392 &  x413 &  x425 &  x428 &  x448 &  x458 &  x467 &  x527 &  x542 &  x548 &  x554 &  x578 &  x584 &  x605 &  x629 &  x644 &  x659 &  x662 &  x668 &  x671 &  x680 &  x692 &  x695 &  x698 &  x716 &  x731 &  x749 &  x782 &  x797 &  x800 &  x809 &  x812 &  x827 &  x845 &  x848 &  x851 &  x896 &  x905 &  x923 &  x938 &  x950 &  x953 &  x974 &  x989 &  x1007 &  x1010 &  x1061 &  x1064 &  x1070 &  x1088 & ~x48 & ~x87 & ~x117 & ~x126 & ~x216 & ~x255 & ~x333 & ~x411 & ~x489 & ~x918 & ~x951 & ~x957 & ~x990 & ~x996 & ~x1029 & ~x1035 & ~x1068 & ~x1074 & ~x1092 & ~x1107;
assign c1254 =  x68 &  x248 &  x269 &  x326 &  x497 &  x511 &  x623 &  x689 &  x844 &  x883 &  x922 &  x1031 & ~x177 & ~x333 & ~x334 & ~x372 & ~x411 & ~x663 & ~x702 & ~x990;
assign c1256 =  x2 &  x23 &  x38 &  x41 &  x44 &  x47 &  x53 &  x56 &  x77 &  x86 &  x89 &  x92 &  x101 &  x104 &  x110 &  x113 &  x122 &  x128 &  x134 &  x143 &  x146 &  x149 &  x152 &  x155 &  x158 &  x173 &  x176 &  x179 &  x182 &  x185 &  x191 &  x194 &  x197 &  x200 &  x206 &  x209 &  x212 &  x215 &  x218 &  x224 &  x227 &  x230 &  x233 &  x269 &  x275 &  x278 &  x287 &  x290 &  x293 &  x296 &  x299 &  x302 &  x305 &  x311 &  x314 &  x317 &  x320 &  x323 &  x329 &  x332 &  x335 &  x343 &  x347 &  x353 &  x365 &  x374 &  x377 &  x380 &  x382 &  x389 &  x392 &  x398 &  x407 &  x410 &  x413 &  x415 &  x421 &  x428 &  x434 &  x437 &  x442 &  x443 &  x446 &  x455 &  x460 &  x461 &  x467 &  x479 &  x482 &  x485 &  x488 &  x491 &  x494 &  x499 &  x500 &  x506 &  x509 &  x515 &  x521 &  x527 &  x530 &  x542 &  x545 &  x554 &  x563 &  x578 &  x581 &  x584 &  x590 &  x599 &  x602 &  x608 &  x611 &  x614 &  x617 &  x626 &  x629 &  x632 &  x638 &  x640 &  x656 &  x665 &  x668 &  x671 &  x677 &  x698 &  x707 &  x710 &  x722 &  x725 &  x728 &  x737 &  x749 &  x752 &  x755 &  x761 &  x764 &  x767 &  x776 &  x782 &  x785 &  x788 &  x791 &  x803 &  x806 &  x815 &  x820 &  x824 &  x827 &  x830 &  x851 &  x859 &  x863 &  x866 &  x875 &  x878 &  x881 &  x887 &  x890 &  x898 &  x901 &  x902 &  x905 &  x908 &  x917 &  x920 &  x923 &  x926 &  x929 &  x935 &  x937 &  x938 &  x940 &  x941 &  x950 &  x953 &  x956 &  x959 &  x965 &  x974 &  x976 &  x977 &  x979 &  x989 &  x995 &  x998 &  x1004 &  x1007 &  x1016 &  x1018 &  x1031 &  x1040 &  x1043 &  x1064 &  x1067 &  x1070 &  x1076 &  x1091 &  x1096 &  x1100 &  x1106 &  x1121 &  x1130 & ~x393 & ~x432 & ~x471 & ~x510 & ~x549 & ~x588 & ~x660 & ~x915 & ~x954 & ~x993 & ~x1032;
assign c1258 =  x68 &  x119 &  x140 &  x170 &  x176 &  x188 &  x227 &  x263 &  x314 &  x317 &  x350 &  x395 &  x422 &  x527 &  x554 &  x596 &  x605 &  x689 &  x716 &  x728 &  x800 &  x860 &  x881 &  x920 &  x940 &  x950 &  x956 &  x1010 &  x1018 &  x1099 & ~x81 & ~x237 & ~x555 & ~x855 & ~x894 & ~x933 & ~x972 & ~x973 & ~x1029 & ~x1068 & ~x1107;
assign c1260 =  x1 &  x22 &  x40 &  x164 &  x185 &  x197 &  x205 &  x284 &  x293 &  x320 &  x326 &  x335 &  x443 &  x485 &  x556 &  x584 &  x596 &  x697 &  x712 &  x716 &  x736 &  x751 &  x785 &  x787 &  x790 &  x800 &  x803 &  x829 &  x833 &  x851 &  x902 &  x946 &  x950 &  x962 &  x985 &  x1024 &  x1063 &  x1093 &  x1100 &  x1102 &  x1120;
assign c1262 =  x80 &  x83 &  x86 &  x143 &  x239 &  x304 &  x317 &  x320 &  x343 &  x344 &  x347 &  x383 &  x386 &  x407 &  x415 &  x443 &  x464 &  x487 &  x578 &  x581 &  x596 &  x638 &  x710 &  x713 &  x722 &  x728 &  x784 &  x794 &  x851 &  x950 &  x989 &  x1040 &  x1106 &  x1121 & ~x399 & ~x750 & ~x816 & ~x855 & ~x951 & ~x990 & ~x1029 & ~x1068;
assign c1264 =  x128 &  x176 &  x185 &  x197 &  x200 &  x206 &  x215 &  x218 &  x224 &  x251 &  x254 &  x320 &  x353 &  x359 &  x401 &  x491 &  x527 &  x553 &  x554 &  x559 &  x590 &  x593 &  x631 &  x674 &  x692 &  x709 &  x715 &  x716 &  x734 &  x748 &  x771 &  x787 &  x830 &  x848 &  x890 &  x896 &  x917 &  x950 &  x953 &  x962 &  x1013 &  x1031 &  x1079 & ~x99 & ~x606 & ~x645;
assign c1266 =  x20 &  x68 &  x107 &  x110 &  x125 &  x176 &  x182 &  x191 &  x194 &  x200 &  x206 &  x215 &  x236 &  x293 &  x302 &  x329 &  x332 &  x347 &  x353 &  x395 &  x422 &  x437 &  x443 &  x445 &  x509 &  x512 &  x527 &  x578 &  x653 &  x680 &  x698 &  x742 &  x749 &  x905 &  x920 &  x932 &  x962 &  x980 &  x995 &  x1022 &  x1046 &  x1085 &  x1091 & ~x87 & ~x165 & ~x198 & ~x204 & ~x276 & ~x282 & ~x315 & ~x393 & ~x432 & ~x732 & ~x733 & ~x738;
assign c1268 =  x23 &  x86 &  x122 &  x155 &  x176 &  x188 &  x269 &  x326 &  x329 &  x356 &  x470 &  x527 &  x536 &  x548 &  x575 &  x578 &  x587 &  x662 &  x670 &  x671 &  x677 &  x680 &  x692 &  x698 &  x713 &  x791 &  x812 &  x845 &  x1019 &  x1058 &  x1079 & ~x334 & ~x372 & ~x459 & ~x624 & ~x663 & ~x780 & ~x781 & ~x820 & ~x898 & ~x1008 & ~x1029;
assign c1270 =  x65 &  x68 &  x119 &  x122 &  x197 &  x212 &  x236 &  x238 &  x251 &  x257 &  x277 &  x316 &  x320 &  x341 &  x344 &  x394 &  x410 &  x419 &  x461 &  x485 &  x491 &  x494 &  x518 &  x530 &  x536 &  x556 &  x569 &  x595 &  x620 &  x623 &  x634 &  x637 &  x665 &  x676 &  x686 &  x700 &  x701 &  x704 &  x715 &  x740 &  x761 &  x845 &  x866 &  x871 &  x881 &  x883 &  x920 &  x934 &  x1067 &  x1084 &  x1090 &  x1097 &  x1127 &  x1129 & ~x303 & ~x819;
assign c1272 =  x2 &  x5 &  x11 &  x20 &  x26 &  x38 &  x56 &  x68 &  x86 &  x101 &  x113 &  x119 &  x146 &  x200 &  x203 &  x218 &  x227 &  x230 &  x236 &  x254 &  x257 &  x275 &  x284 &  x302 &  x308 &  x329 &  x335 &  x353 &  x359 &  x377 &  x383 &  x392 &  x395 &  x443 &  x449 &  x461 &  x470 &  x472 &  x476 &  x497 &  x509 &  x533 &  x554 &  x556 &  x584 &  x587 &  x593 &  x594 &  x595 &  x605 &  x614 &  x620 &  x623 &  x626 &  x634 &  x650 &  x671 &  x673 &  x698 &  x701 &  x707 &  x709 &  x712 &  x716 &  x728 &  x737 &  x748 &  x751 &  x767 &  x787 &  x790 &  x800 &  x839 &  x851 &  x857 &  x860 &  x875 &  x881 &  x890 &  x908 &  x911 &  x914 &  x920 &  x956 &  x974 &  x977 &  x989 &  x1007 &  x1043 &  x1046 &  x1052 &  x1064 &  x1100 &  x1109 &  x1124 & ~x348 & ~x645 & ~x684 & ~x723;
assign c1274 =  x19 &  x23 &  x32 &  x35 &  x38 &  x41 &  x47 &  x50 &  x56 &  x68 &  x86 &  x94 &  x107 &  x133 &  x134 &  x206 &  x218 &  x221 &  x227 &  x236 &  x266 &  x269 &  x275 &  x281 &  x284 &  x290 &  x293 &  x302 &  x317 &  x335 &  x362 &  x394 &  x434 &  x446 &  x482 &  x491 &  x503 &  x506 &  x509 &  x521 &  x554 &  x566 &  x578 &  x581 &  x590 &  x592 &  x596 &  x611 &  x617 &  x631 &  x641 &  x670 &  x677 &  x689 &  x701 &  x709 &  x716 &  x719 &  x725 &  x731 &  x734 &  x764 &  x767 &  x770 &  x787 &  x797 &  x800 &  x809 &  x826 &  x833 &  x845 &  x848 &  x851 &  x865 &  x884 &  x896 &  x904 &  x911 &  x917 &  x923 &  x926 &  x950 &  x980 &  x989 &  x1007 &  x1010 &  x1013 &  x1033 &  x1037 &  x1082 &  x1088 &  x1100 &  x1103 &  x1118 &  x1129 & ~x663 & ~x702 & ~x936 & ~x1017;
assign c1276 =  x199 &  x277 &  x316 &  x458 &  x474 &  x553 &  x592 &  x593 &  x631 &  x655 &  x709 &  x787 &  x844 &  x883 &  x994 & ~x528 & ~x546 & ~x702 & ~x741;
assign c1278 =  x5 &  x8 &  x11 &  x29 &  x35 &  x50 &  x53 &  x59 &  x89 &  x95 &  x122 &  x125 &  x131 &  x137 &  x143 &  x146 &  x161 &  x164 &  x179 &  x194 &  x218 &  x224 &  x236 &  x242 &  x254 &  x257 &  x293 &  x302 &  x311 &  x314 &  x316 &  x320 &  x326 &  x332 &  x335 &  x344 &  x355 &  x365 &  x377 &  x380 &  x394 &  x416 &  x431 &  x437 &  x443 &  x472 &  x479 &  x491 &  x497 &  x506 &  x518 &  x527 &  x542 &  x545 &  x569 &  x578 &  x584 &  x587 &  x593 &  x605 &  x629 &  x638 &  x641 &  x668 &  x670 &  x677 &  x689 &  x704 &  x707 &  x734 &  x749 &  x758 &  x761 &  x773 &  x785 &  x797 &  x803 &  x806 &  x818 &  x844 &  x848 &  x854 &  x857 &  x860 &  x863 &  x875 &  x883 &  x890 &  x902 &  x914 &  x920 &  x922 &  x923 &  x950 &  x959 &  x961 &  x962 &  x977 &  x989 &  x995 &  x998 &  x1001 &  x1040 &  x1049 &  x1076 &  x1094 &  x1106 & ~x99 & ~x342 & ~x420 & ~x585 & ~x600 & ~x663 & ~x702 & ~x780 & ~x990 & ~x1014 & ~x1029 & ~x1068 & ~x1107;
assign c1280 =  x47 &  x53 &  x131 &  x160 &  x164 &  x191 &  x206 &  x215 &  x248 &  x263 &  x275 &  x284 &  x308 &  x316 &  x317 &  x338 &  x359 &  x410 &  x416 &  x431 &  x434 &  x439 &  x527 &  x530 &  x536 &  x553 &  x590 &  x611 &  x617 &  x670 &  x671 &  x677 &  x692 &  x734 &  x749 &  x779 &  x833 &  x851 &  x869 &  x902 &  x917 &  x926 &  x932 &  x935 &  x950 &  x956 &  x977 &  x1013 &  x1025 &  x1034 &  x1058 & ~x309 & ~x486 & ~x585 & ~x663 & ~x742 & ~x781 & ~x820 & ~x897;
assign c1282 =  x1 &  x17 &  x29 &  x38 &  x41 &  x47 &  x107 &  x113 &  x119 &  x176 &  x200 &  x224 &  x236 &  x239 &  x245 &  x251 &  x311 &  x317 &  x326 &  x332 &  x353 &  x365 &  x371 &  x406 &  x413 &  x437 &  x440 &  x443 &  x452 &  x484 &  x491 &  x493 &  x499 &  x523 &  x532 &  x536 &  x538 &  x539 &  x542 &  x545 &  x559 &  x562 &  x571 &  x572 &  x578 &  x601 &  x629 &  x640 &  x641 &  x668 &  x671 &  x680 &  x689 &  x692 &  x698 &  x716 &  x728 &  x734 &  x740 &  x746 &  x749 &  x767 &  x773 &  x781 &  x788 &  x794 &  x803 &  x809 &  x819 &  x820 &  x827 &  x859 &  x866 &  x896 &  x897 &  x905 &  x920 &  x923 &  x926 &  x929 &  x935 &  x937 &  x950 &  x956 &  x965 &  x971 &  x1010 &  x1015 &  x1019 &  x1031 &  x1063 &  x1064 &  x1076 &  x1085 &  x1093 &  x1100 &  x1102 & ~x237 & ~x315 & ~x393 & ~x432 & ~x471 & ~x510 & ~x549 & ~x588 & ~x627;
assign c1284 =  x44 &  x47 &  x53 &  x83 &  x89 &  x101 &  x116 &  x143 &  x173 &  x191 &  x218 &  x233 &  x257 &  x278 &  x280 &  x290 &  x296 &  x314 &  x317 &  x323 &  x326 &  x329 &  x335 &  x353 &  x359 &  x365 &  x383 &  x386 &  x389 &  x395 &  x404 &  x407 &  x416 &  x475 &  x476 &  x482 &  x518 &  x520 &  x524 &  x527 &  x548 &  x553 &  x559 &  x572 &  x578 &  x592 &  x596 &  x597 &  x598 &  x631 &  x637 &  x656 &  x662 &  x665 &  x668 &  x670 &  x671 &  x676 &  x692 &  x701 &  x704 &  x715 &  x716 &  x728 &  x754 &  x767 &  x782 &  x785 &  x796 &  x803 &  x815 &  x824 &  x832 &  x857 &  x871 &  x910 &  x917 &  x920 &  x956 &  x974 &  x983 &  x989 &  x998 &  x1004 &  x1028 &  x1076 &  x1091 &  x1115 &  x1117 &  x1121;
assign c1286 =  x5 &  x23 &  x308 &  x329 &  x398 &  x431 &  x470 &  x473 &  x527 &  x551 &  x797 &  x854 &  x884 &  x1004 &  x1016 &  x1115 & ~x324 & ~x363 & ~x384 & ~x402 & ~x618 & ~x924 & ~x948 & ~x987 & ~x1026 & ~x1029 & ~x1050 & ~x1065 & ~x1068 & ~x1104 & ~x1107;
assign c1288 =  x20 &  x116 &  x128 &  x302 &  x322 &  x437 &  x506 &  x542 &  x556 &  x578 &  x595 &  x605 &  x620 &  x698 &  x715 &  x743 &  x799 &  x838 &  x877 &  x956 & ~x45 & ~x84 & ~x420 & ~x498 & ~x1017;
assign c1290 =  x14 &  x31 &  x53 &  x95 &  x152 &  x164 &  x169 &  x176 &  x224 &  x239 &  x257 &  x263 &  x272 &  x302 &  x304 &  x325 &  x382 &  x383 &  x395 &  x406 &  x431 &  x464 &  x479 &  x536 &  x545 &  x578 &  x581 &  x593 &  x596 &  x599 &  x620 &  x632 &  x656 &  x665 &  x668 &  x713 &  x731 &  x734 &  x767 &  x773 &  x904 &  x926 &  x938 &  x940 &  x946 &  x953 &  x968 &  x985 &  x995 &  x1007 &  x1010 &  x1018 &  x1028 &  x1058 &  x1064 &  x1106 &  x1109 & ~x276 & ~x315;
assign c1292 =  x2 &  x11 &  x14 &  x17 &  x35 &  x38 &  x44 &  x68 &  x71 &  x74 &  x77 &  x86 &  x101 &  x107 &  x134 &  x140 &  x152 &  x164 &  x173 &  x176 &  x215 &  x218 &  x230 &  x236 &  x245 &  x248 &  x254 &  x260 &  x263 &  x275 &  x278 &  x284 &  x299 &  x302 &  x317 &  x335 &  x338 &  x341 &  x344 &  x365 &  x371 &  x374 &  x392 &  x406 &  x413 &  x437 &  x440 &  x443 &  x445 &  x455 &  x473 &  x482 &  x485 &  x494 &  x509 &  x527 &  x551 &  x554 &  x572 &  x578 &  x584 &  x586 &  x589 &  x632 &  x641 &  x656 &  x659 &  x671 &  x683 &  x686 &  x692 &  x695 &  x698 &  x706 &  x710 &  x728 &  x731 &  x734 &  x745 &  x758 &  x767 &  x770 &  x776 &  x784 &  x800 &  x803 &  x818 &  x827 &  x851 &  x866 &  x872 &  x890 &  x896 &  x902 &  x920 &  x929 &  x956 &  x974 &  x995 &  x1004 &  x1007 &  x1028 &  x1067 &  x1079 &  x1088 &  x1124 & ~x234 & ~x474 & ~x576 & ~x615 & ~x616 & ~x654 & ~x655 & ~x678 & ~x693 & ~x694 & ~x732 & ~x795;
assign c1294 =  x47 &  x116 &  x164 &  x194 &  x218 &  x299 &  x302 &  x359 &  x386 &  x473 &  x527 &  x542 &  x560 &  x599 &  x728 &  x734 &  x767 &  x818 &  x866 &  x905 &  x914 &  x935 &  x938 &  x950 &  x974 &  x1022 &  x1025 &  x1049 &  x1076 & ~x690 & ~x729 & ~x738 & ~x753 & ~x793 & ~x816 & ~x948 & ~x1029 & ~x1050 & ~x1107;
assign c1296 =  x8 &  x11 &  x20 &  x41 &  x47 &  x71 &  x80 &  x86 &  x122 &  x134 &  x173 &  x176 &  x182 &  x191 &  x194 &  x200 &  x214 &  x218 &  x253 &  x269 &  x275 &  x278 &  x281 &  x284 &  x302 &  x311 &  x326 &  x328 &  x341 &  x347 &  x356 &  x365 &  x367 &  x389 &  x406 &  x437 &  x443 &  x445 &  x455 &  x473 &  x509 &  x512 &  x518 &  x527 &  x550 &  x560 &  x575 &  x578 &  x586 &  x593 &  x623 &  x625 &  x628 &  x644 &  x659 &  x668 &  x706 &  x716 &  x734 &  x749 &  x773 &  x784 &  x785 &  x827 &  x851 &  x866 &  x881 &  x890 &  x896 &  x899 &  x914 &  x950 &  x959 &  x1007 &  x1025 &  x1045 &  x1084 &  x1112 &  x1123 & ~x360 & ~x435 & ~x474 & ~x513;
assign c1298 =  x20 &  x26 &  x38 &  x41 &  x47 &  x50 &  x62 &  x68 &  x83 &  x86 &  x98 &  x122 &  x197 &  x221 &  x227 &  x248 &  x263 &  x284 &  x290 &  x311 &  x332 &  x335 &  x341 &  x356 &  x362 &  x365 &  x401 &  x413 &  x437 &  x472 &  x473 &  x485 &  x509 &  x511 &  x518 &  x521 &  x524 &  x560 &  x575 &  x592 &  x641 &  x670 &  x677 &  x698 &  x707 &  x709 &  x734 &  x749 &  x755 &  x761 &  x787 &  x788 &  x826 &  x839 &  x878 &  x884 &  x968 &  x1004 &  x1058 &  x1088 &  x1106 &  x1112 &  x1121 & ~x450 & ~x489 & ~x490 & ~x528 & ~x529 & ~x567 & ~x606 & ~x645 & ~x663 & ~x702;
assign c11 = ~x248;
assign c13 =  x8 &  x14 &  x41 &  x46 &  x104 &  x119 &  x185 &  x212 &  x227 &  x344 &  x359 &  x392 &  x395 &  x413 &  x544 &  x578 &  x668 &  x719 &  x755 &  x767 &  x785 &  x815 &  x818 &  x853 &  x863 &  x875 &  x890 &  x950 &  x995 &  x1013 &  x1037 &  x1040 &  x1064 &  x1087 &  x1114 &  x1124 &  x1126 & ~x345;
assign c15 =  x496 &  x691 & ~x676;
assign c17 = ~x980;
assign c19 =  x936 & ~x796 & ~x904;
assign c111 = ~x59;
assign c113 =  x168 & ~x249;
assign c115 =  x67 &  x622 &  x724 &  x730 &  x1048 &  x1092 & ~x933;
assign c117 = ~x54 & ~x183 & ~x982;
assign c119 = ~x135 & ~x1051 & ~x1060;
assign c121 = ~x16 & ~x55 & ~x786 & ~x885 & ~x945;
assign c123 = ~x401;
assign c125 =  x281 &  x428 &  x856 &  x928 &  x1039 & ~x93 & ~x147 & ~x240 & ~x1053;
assign c127 =  x385 &  x424 &  x529 &  x568 &  x574 &  x622 &  x830 &  x853 &  x1111;
assign c131 = ~x1018;
assign c133 =  x356 &  x379 &  x691 &  x742 &  x806;
assign c135 =  x6 &  x7 &  x77 &  x179 &  x383 &  x658 &  x685 &  x731 &  x814 &  x815 &  x830 &  x853 &  x956 &  x971 &  x1124;
assign c137 =  x679 &  x864;
assign c139 =  x467 &  x488 &  x857 & ~x174 & ~x747 & ~x981 & ~x1098 & ~x1119;
assign c141 =  x451 &  x588;
assign c143 =  x951 &  x1087 & ~x846;
assign c145 =  x46 &  x874 &  x1087 & ~x156;
assign c147 =  x373 &  x490 &  x588 &  x660;
assign c149 =  x346 &  x457 &  x644 &  x652 &  x1001 & ~x135 & ~x174 & ~x297 & ~x441;
assign c151 =  x257 &  x625 &  x717 &  x794 &  x845 &  x973 & ~x861;
assign c153 = ~x631;
assign c155 =  x7 &  x739 &  x999;
assign c157 = ~x602 & ~x791;
assign c159 =  x9 &  x23 &  x464 &  x533 &  x647 &  x889 &  x1066 &  x1105 & ~x906 & ~x945;
assign c161 =  x226 &  x652 & ~x486 & ~x564 & ~x708 & ~x747 & ~x1119;
assign c163 =  x574 &  x955 &  x1066 & ~x75 & ~x174 & ~x297 & ~x375 & ~x414 & ~x663;
assign c165 =  x87 &  x273 & ~x297;
assign c169 =  x441 &  x477;
assign c171 =  x161 &  x163 &  x358 &  x397 &  x627 & ~x708 & ~x747;
assign c173 =  x385 & ~x220 & ~x258 & ~x780 & ~x1080;
assign c175 = ~x569;
assign c177 =  x67 &  x505 &  x529 &  x544 &  x568 &  x574 &  x596 &  x661 &  x752 &  x812 &  x914 &  x962 &  x1028 &  x1030 &  x1087;
assign c179 =  x112 &  x261 &  x451 &  x622 &  x970 &  x1030;
assign c181 =  x707 & ~x39 & ~x93 & ~x171 & ~x288 & ~x484 & ~x945;
assign c183 = ~x95;
assign c185 =  x969 & ~x156 & ~x882;
assign c187 =  x480 &  x558 &  x789;
assign c189 = ~x523 & ~x672;
assign c191 =  x241 &  x853 & ~x531 & ~x570 & ~x708 & ~x726 & ~x1122;
assign c193 =  x126 &  x754 & ~x219 & ~x258 & ~x891;
assign c195 = ~x617;
assign c197 = ~x514 & ~x784;
assign c199 =  x412 &  x451 &  x529 &  x660;
assign c1101 =  x724 &  x999 & ~x132 & ~x930;
assign c1103 =  x679 &  x1104;
assign c1105 = ~x39 & ~x747 & ~x1057;
assign c1107 =  x358 & ~x316 & ~x714 & ~x945;
assign c1109 =  x27 &  x379 &  x723;
assign c1113 = ~x866;
assign c1115 =  x716 & ~x174 & ~x258 & ~x807;
assign c1117 = ~x377;
assign c1119 = ~x436 & ~x745;
assign c1121 =  x412 &  x840 & ~x78;
assign c1123 =  x204;
assign c1125 =  x1069 & ~x787;
assign c1127 =  x1107 & ~x1045;
assign c1129 = ~x436;
assign c1131 =  x46 &  x352 &  x682 &  x734 &  x999;
assign c1133 =  x477 &  x624;
assign c1135 =  x11 &  x350 &  x568 &  x575 &  x607 &  x632 &  x760 &  x892 &  x1007 &  x1018 &  x1094 & ~x687;
assign c1137 =  x466 &  x505 & ~x540 & ~x648 & ~x981 & ~x1122;
assign c1139 = ~x380;
assign c1143 =  x64 &  x97 &  x475 &  x965 &  x985 & ~x1020;
assign c1145 =  x202 &  x913 & ~x144 & ~x339 & ~x765;
assign c1147 =  x516 & ~x687;
assign c1149 =  x46 & ~x183 & ~x823;
assign c1151 = ~x224;
assign c1153 =  x234 & ~x93 & ~x511;
assign c1155 =  x457 &  x496 & ~x414 & ~x442 & ~x481;
assign c1157 = ~x712;
assign c1159 =  x148 &  x1048 & ~x885 & ~x1117;
assign c1161 = ~x122;
assign c1163 = ~x644;
assign c1165 =  x64 &  x319 &  x557 &  x839 &  x1115 & ~x609 & ~x648 & ~x828;
assign c1167 =  x358 &  x433 & ~x592;
assign c1169 =  x226 &  x229 &  x334 &  x358 &  x435 & ~x561 & ~x600;
assign c1171 =  x645 &  x723 &  x762 &  x895;
assign c1173 =  x202 &  x319 &  x1107 & ~x234;
assign c1175 =  x126 &  x165 &  x200 &  x244 &  x371 &  x613 &  x760 &  x869;
assign c1177 = ~x1046;
assign c1179 = ~x253 & ~x400;
assign c1181 =  x428 &  x466 &  x622 &  x892 &  x1008 &  x1030;
assign c1183 =  x319 &  x349 &  x784 & ~x1098;
assign c1185 = ~x358 & ~x666 & ~x784;
assign c1187 =  x64 &  x652 &  x965 &  x1034 & ~x687 & ~x789 & ~x828;
assign c1189 = ~x197;
assign c1191 =  x85 &  x299 &  x737 &  x874 &  x1067 &  x1127 & ~x183 & ~x339 & ~x1095;
assign c1193 =  x319 &  x397 &  x1087 & ~x787 & ~x826;
assign c1195 =  x757 &  x1012 & ~x39 & ~x339 & ~x378 & ~x414;
assign c1197 =  x28 &  x622 &  x951 &  x1030;
assign c1199 = ~x40 & ~x183 & ~x492 & ~x864;
assign c1201 =  x53 &  x86 &  x236 &  x352 &  x374 &  x410 &  x437 &  x524 &  x560 &  x688 &  x923 &  x983 &  x986 &  x1066 &  x1079 &  x1118 & ~x297 & ~x336 & ~x441;
assign c1203 =  x574 &  x723;
assign c1205 =  x46 & ~x765 & ~x864 & ~x889;
assign c1207 = ~x286 & ~x937;
assign c1209 =  x631 & ~x414 & ~x667;
assign c1211 =  x639 &  x1072 & ~x453;
assign c1213 =  x49 & ~x96 & ~x297 & ~x318 & ~x906;
assign c1215 =  x702 & ~x709 & ~x1122;
assign c1217 =  x749 &  x756 &  x912 &  x1048;
assign c1221 =  x338 &  x500 & ~x181 & ~x220 & ~x259 & ~x846 & ~x867;
assign c1223 =  x103 &  x936 & ~x796;
assign c1225 =  x530 &  x544 &  x705 &  x710 &  x856 &  x952 &  x1067;
assign c1227 =  x931 & ~x844 & ~x943;
assign c1229 = ~x796 & ~x982;
assign c1231 =  x343 &  x478 & ~x570 & ~x1000;
assign c1233 =  x12 & ~x1041;
assign c1237 =  x451 & ~x679;
assign c1239 =  x952 &  x982 & ~x183 & ~x687;
assign c1241 =  x679 & ~x436;
assign c1243 = ~x30 & ~x105 & ~x339 & ~x747 & ~x981;
assign c1245 =  x45 & ~x219 & ~x406;
assign c1247 = ~x253 & ~x604;
assign c1249 =  x97 &  x691 &  x780;
assign c1251 = ~x539;
assign c1253 =  x717 & ~x570 & ~x783;
assign c1255 =  x1077 & ~x261 & ~x330 & ~x369 & ~x453;
assign c1257 = ~x200;
assign c1259 =  x1077 & ~x39 & ~x223;
assign c1261 = ~x748 & ~x861;
assign c1263 =  x477 &  x858 & ~x610;
assign c1265 = ~x111 & ~x132 & ~x249 & ~x648 & ~x687 & ~x864 & ~x903 & ~x981;
assign c1267 =  x529 &  x622 &  x681 &  x1030;
assign c1269 =  x165 & ~x249;
assign c1271 = ~x251;
assign c1273 =  x13 &  x26 &  x505 &  x653 &  x952 & ~x183 & ~x222 & ~x249 & ~x300;
assign c1275 =  x7 &  x25 &  x163 &  x934 &  x991 & ~x747;
assign c1277 =  x257 &  x854 &  x893 &  x983 &  x1106 & ~x144 & ~x261 & ~x262 & ~x807 & ~x846 & ~x945 & ~x1041;
assign c1279 =  x5 &  x188 &  x226 &  x254 &  x518 &  x745 & ~x765 & ~x1078;
assign c1281 =  x358 &  x613 & ~x637 & ~x715;
assign c1283 =  x319 &  x422 &  x508 &  x857 & ~x93 & ~x105 & ~x453;
assign c1285 =  x502 & ~x297 & ~x376 & ~x930;
assign c1287 =  x48 &  x312 &  x1060 &  x1117;
assign c1289 =  x161 &  x418 &  x557 &  x632 &  x688 &  x782 &  x908 & ~x403 & ~x867;
assign c1291 =  x7 & ~x57 & ~x147 & ~x1080;
assign c1293 =  x451 &  x529 &  x534 &  x613 &  x622 &  x661;
assign c1295 =  x80 &  x86 &  x110 &  x298 &  x319 &  x524 &  x611 &  x671 &  x704 &  x713 &  x773 &  x803 &  x1058 &  x1085 & ~x330 & ~x399 & ~x903 & ~x981 & ~x1098;
assign c1297 =  x352 &  x1060 & ~x93 & ~x288 & ~x846 & ~x976;
assign c1299 =  x46 &  x371 &  x544 &  x574 &  x577 & ~x897 & ~x1023;
assign c20 =  x50 &  x325 &  x338 &  x359 &  x400 &  x428 &  x478 &  x638 &  x674 &  x758 &  x803 &  x833 &  x944 &  x974 &  x989 &  x992 &  x1022 &  x1034 &  x1085 & ~x600 & ~x639 & ~x825 & ~x1038 & ~x1119;
assign c22 =  x199 &  x277 &  x302 &  x632 &  x725 &  x1022 & ~x378 & ~x414 & ~x453 & ~x492 & ~x531 & ~x570 & ~x648 & ~x666 & ~x744 & ~x1014 & ~x1074;
assign c24 = ~x0 & ~x33 & ~x48 & ~x72 & ~x111 & ~x261 & ~x339 & ~x456 & ~x531 & ~x570 & ~x633 & ~x687 & ~x804 & ~x900;
assign c26 =  x2 &  x38 &  x110 &  x122 &  x139 &  x152 &  x158 &  x173 &  x191 &  x209 &  x217 &  x230 &  x233 &  x236 &  x290 &  x296 &  x302 &  x308 &  x323 &  x440 &  x451 &  x458 &  x461 &  x467 &  x488 &  x490 &  x533 &  x539 &  x545 &  x581 &  x586 &  x590 &  x607 &  x614 &  x629 &  x635 &  x644 &  x664 &  x695 &  x703 &  x719 &  x725 &  x742 &  x821 &  x839 &  x859 &  x892 &  x902 &  x911 &  x919 &  x947 &  x1007 &  x1015 &  x1034 &  x1058 &  x1070 &  x1076 &  x1091 &  x1094 &  x1121 & ~x888 & ~x927 & ~x942 & ~x981 & ~x1038 & ~x1056;
assign c28 =  x124 &  x233 &  x241 &  x389 &  x505 &  x601 &  x679 &  x874 &  x991 &  x1009 &  x1030 &  x1048 &  x1126 & ~x441;
assign c210 =  x14 &  x215 &  x345 &  x385 &  x419 &  x757 &  x941 &  x989 & ~x63 & ~x64 & ~x129 & ~x627 & ~x705;
assign c212 =  x29 &  x101 &  x110 &  x122 &  x266 &  x401 &  x431 &  x623 &  x667 &  x710 &  x866 &  x989 &  x1010 &  x1043 &  x1109 & ~x786 & ~x804 & ~x825 & ~x844 & ~x864 & ~x870 & ~x954 & ~x1020 & ~x1038 & ~x1089;
assign c214 =  x160 &  x200 &  x423 &  x424 &  x462 &  x501 &  x502 &  x601 &  x640 &  x658 &  x718 &  x719 &  x743 &  x757 &  x814 &  x835 &  x874 &  x913 &  x952 &  x991 &  x1100 &  x1106 & ~x627;
assign c216 =  x220 &  x347 &  x439 &  x500 &  x512 &  x524 &  x667 &  x989 &  x995 &  x1037 & ~x687 & ~x882 & ~x903 & ~x904 & ~x921 & ~x1038;
assign c218 =  x5 &  x11 &  x41 &  x43 &  x68 &  x80 &  x86 &  x104 &  x121 &  x128 &  x146 &  x160 &  x170 &  x173 &  x196 &  x199 &  x272 &  x290 &  x346 &  x353 &  x356 &  x434 &  x457 &  x497 &  x500 &  x502 &  x503 &  x524 &  x539 &  x542 &  x563 &  x572 &  x587 &  x601 &  x605 &  x614 &  x640 &  x668 &  x679 &  x689 &  x716 &  x725 &  x839 &  x845 &  x854 &  x926 &  x929 &  x938 &  x953 &  x989 &  x992 &  x1022 &  x1058 &  x1082 &  x1100 &  x1118 & ~x918 & ~x1035;
assign c220 =  x2 &  x23 &  x125 &  x182 &  x191 &  x206 &  x269 &  x278 &  x334 &  x362 &  x412 &  x490 &  x521 &  x566 &  x640 &  x704 &  x835 &  x841 &  x965 &  x1010 &  x1019 &  x1076 &  x1115 & ~x420 & ~x421 & ~x459 & ~x498;
assign c222 =  x101 &  x286 &  x332 &  x439 &  x725 &  x929 &  x1028 & ~x639 & ~x651 & ~x690 & ~x729 & ~x747 & ~x786 & ~x903 & ~x978;
assign c224 =  x41 &  x80 &  x113 &  x154 &  x170 &  x359 &  x380 &  x392 &  x526 &  x539 &  x563 &  x565 &  x647 &  x650 &  x662 &  x716 &  x721 &  x728 &  x773 &  x790 &  x796 &  x824 &  x866 &  x929 &  x1010 &  x1104 &  x1105;
assign c226 =  x81 &  x86 &  x120 &  x121 &  x159 &  x191 &  x218 &  x317 &  x386 &  x506 &  x518 &  x641 &  x674 &  x710 &  x770 &  x785 &  x824 &  x851 &  x869 &  x881 &  x884 &  x956 &  x989 &  x995 &  x1004 &  x1019 &  x1082 &  x1102 &  x1121 & ~x321 & ~x606 & ~x702;
assign c228 =  x416 &  x487 &  x553 &  x745 & ~x429 & ~x687 & ~x864 & ~x1017 & ~x1038;
assign c230 =  x26 &  x47 &  x65 &  x77 &  x92 &  x107 &  x143 &  x146 &  x209 &  x218 &  x266 &  x272 &  x277 &  x278 &  x281 &  x302 &  x305 &  x311 &  x329 &  x392 &  x407 &  x410 &  x422 &  x430 &  x469 &  x470 &  x515 &  x629 &  x640 &  x656 &  x683 &  x707 &  x776 &  x791 &  x875 &  x890 &  x908 &  x923 &  x962 &  x977 &  x980 &  x989 &  x1010 &  x1016 &  x1055 &  x1097 &  x1121 & ~x324 & ~x363 & ~x480 & ~x492 & ~x519 & ~x531 & ~x597 & ~x627 & ~x666 & ~x667 & ~x705 & ~x706 & ~x822;
assign c232 =  x11 &  x23 &  x29 &  x53 &  x56 &  x86 &  x95 &  x110 &  x155 &  x185 &  x209 &  x239 &  x299 &  x332 &  x344 &  x371 &  x463 &  x470 &  x502 &  x524 &  x533 &  x566 &  x569 &  x587 &  x596 &  x599 &  x605 &  x614 &  x620 &  x623 &  x668 &  x731 &  x740 &  x782 &  x788 &  x815 &  x824 &  x836 &  x854 &  x878 &  x920 &  x923 &  x950 &  x989 &  x995 &  x1058 &  x1100 & ~x246 & ~x279 & ~x285 & ~x336 & ~x357 & ~x363 & ~x414 & ~x550 & ~x588 & ~x589 & ~x627 & ~x666;
assign c234 =  x35 &  x47 &  x92 &  x134 &  x152 &  x203 &  x230 &  x350 &  x440 &  x493 &  x527 &  x553 &  x584 &  x587 &  x665 &  x713 &  x740 &  x745 &  x872 &  x917 &  x1001 &  x1040 &  x1094 &  x1124 & ~x312 & ~x391 & ~x429 & ~x430 & ~x469 & ~x508 & ~x546 & ~x729 & ~x807 & ~x885 & ~x1038;
assign c236 =  x26 &  x44 &  x425 &  x455 &  x503 &  x526 &  x565 &  x603 &  x604 &  x638 &  x643 &  x712 &  x728 &  x760 &  x821 &  x854 &  x908 &  x959 &  x989 &  x1049 & ~x1117;
assign c238 =  x100 &  x139 &  x178 &  x436 &  x782 &  x813 &  x991 & ~x519 & ~x687;
assign c240 =  x14 &  x451 &  x1048 &  x1063 &  x1069 &  x1093 &  x1102 &  x1108 & ~x1000 & ~x1038 & ~x1039;
assign c242 =  x181 &  x221 &  x439 &  x455 &  x478 &  x569 &  x620 &  x962 & ~x534 & ~x573 & ~x574 & ~x612 & ~x630 & ~x669 & ~x708;
assign c244 =  x46 &  x85 &  x155 &  x158 &  x269 &  x277 &  x299 &  x383 &  x494 &  x502 &  x517 &  x544 &  x620 &  x701 &  x707 &  x710 &  x758 &  x814 &  x851 &  x868 &  x896 &  x995 &  x1022 &  x1043 &  x1052 & ~x627 & ~x744;
assign c246 =  x710 & ~x414 & ~x453 & ~x492 & ~x555 & ~x570 & ~x609 & ~x610 & ~x630 & ~x648 & ~x687 & ~x786 & ~x804 & ~x843 & ~x861 & ~x882;
assign c248 =  x8 &  x29 &  x38 &  x77 &  x86 &  x101 &  x107 &  x110 &  x131 &  x155 &  x206 &  x212 &  x218 &  x224 &  x227 &  x233 &  x239 &  x254 &  x275 &  x281 &  x326 &  x335 &  x353 &  x356 &  x358 &  x392 &  x407 &  x416 &  x431 &  x464 &  x500 &  x533 &  x539 &  x557 &  x569 &  x575 &  x584 &  x602 &  x608 &  x650 &  x710 &  x764 &  x773 &  x797 &  x803 &  x830 &  x854 &  x893 &  x896 &  x902 &  x914 &  x932 &  x1010 &  x1034 &  x1052 &  x1076 &  x1097 & ~x234 & ~x558 & ~x636 & ~x648 & ~x675 & ~x687 & ~x726 & ~x753 & ~x786 & ~x792 & ~x804 & ~x843 & ~x882 & ~x903 & ~x1017 & ~x1056;
assign c250 =  x59 &  x140 &  x200 &  x236 &  x290 &  x335 &  x365 &  x401 &  x419 &  x434 &  x452 &  x473 &  x725 &  x923 &  x1010 &  x1067 &  x1073 &  x1085 & ~x72 & ~x111 & ~x306 & ~x495 & ~x534 & ~x570 & ~x612 & ~x648 & ~x687 & ~x717 & ~x726 & ~x747 & ~x786 & ~x825 & ~x864 & ~x978;
assign c252 =  x278 & ~x66 & ~x138 & ~x300 & ~x457 & ~x495 & ~x573 & ~x708 & ~x1089;
assign c254 =  x7 &  x32 &  x68 &  x74 &  x98 &  x107 &  x122 &  x160 &  x173 &  x224 &  x227 &  x230 &  x260 &  x277 &  x365 &  x407 &  x440 &  x446 &  x487 &  x488 &  x505 &  x526 &  x544 &  x565 &  x596 &  x626 &  x640 &  x656 &  x716 &  x722 &  x760 &  x764 &  x773 &  x814 &  x818 &  x835 &  x857 &  x869 &  x874 &  x913 &  x941 &  x994 &  x1022 &  x1033 &  x1088;
assign c256 =  x14 &  x122 &  x137 &  x683 &  x725 & ~x54 & ~x111 & ~x261 & ~x378 & ~x456 & ~x786 & ~x804 & ~x880 & ~x918 & ~x1035;
assign c258 =  x35 &  x68 &  x77 &  x83 &  x92 &  x101 &  x110 &  x122 &  x124 &  x149 &  x163 &  x182 &  x197 &  x218 &  x227 &  x233 &  x242 &  x248 &  x263 &  x277 &  x283 &  x316 &  x329 &  x398 &  x422 &  x434 &  x440 &  x446 &  x452 &  x482 &  x533 &  x544 &  x548 &  x587 &  x611 &  x640 &  x647 &  x679 &  x680 &  x710 &  x716 &  x719 &  x725 &  x740 &  x773 &  x779 &  x785 &  x796 &  x806 &  x812 &  x835 &  x845 &  x887 &  x923 &  x929 &  x977 &  x1007 &  x1010 &  x1037 &  x1046 &  x1052 &  x1070 &  x1106 & ~x117 & ~x627 & ~x666 & ~x705;
assign c260 =  x59 &  x95 &  x635 &  x1109 & ~x0 & ~x9 & ~x33 & ~x54 & ~x72 & ~x87 & ~x93 & ~x111 & ~x597 & ~x804 & ~x825 & ~x861 & ~x900;
assign c262 =  x32 &  x83 &  x143 &  x200 &  x275 &  x278 &  x281 &  x317 &  x396 &  x407 &  x464 &  x472 &  x521 &  x547 &  x563 &  x586 &  x614 &  x653 &  x689 &  x710 &  x758 &  x827 &  x851 &  x977 &  x1028 &  x1102 &  x1121 & ~x687 & ~x1038;
assign c264 =  x113 &  x271 &  x286 &  x486 &  x487 &  x745 &  x1108 & ~x429 & ~x430 & ~x546;
assign c266 =  x122 &  x286 &  x364 &  x370 &  x448 &  x526 &  x565 &  x604 &  x977 &  x1097 & ~x687 & ~x690 & ~x867 & ~x906 & ~x1038;
assign c268 =  x23 &  x56 &  x125 &  x134 &  x143 &  x152 &  x179 &  x182 &  x197 &  x221 &  x236 &  x248 &  x254 &  x269 &  x275 &  x293 &  x329 &  x352 &  x380 &  x413 &  x467 &  x470 &  x476 &  x530 &  x539 &  x554 &  x563 &  x584 &  x587 &  x601 &  x605 &  x611 &  x617 &  x620 &  x640 &  x644 &  x647 &  x671 &  x683 &  x695 &  x698 &  x731 &  x757 &  x758 &  x764 &  x796 &  x800 &  x812 &  x839 &  x842 &  x869 &  x914 &  x935 &  x950 &  x980 &  x1019 &  x1022 &  x1037 &  x1055 &  x1064 &  x1097 &  x1106 &  x1109 &  x1112 & ~x66 & ~x105 & ~x106 & ~x144 & ~x183 & ~x222 & ~x223 & ~x261 & ~x588 & ~x663;
assign c270 =  x42 &  x83 &  x179 &  x194 &  x329 &  x371 &  x419 &  x434 &  x458 &  x689 &  x782 &  x788 &  x874 &  x896 &  x932 &  x952 &  x968 &  x988 &  x991 &  x1073 &  x1097 &  x1108 & ~x27 & ~x468 & ~x606 & ~x645;
assign c272 =  x68 &  x83 &  x89 &  x98 &  x188 &  x215 &  x238 &  x278 &  x281 &  x293 &  x359 &  x377 &  x391 &  x404 &  x458 &  x464 &  x473 &  x491 &  x506 &  x548 &  x560 &  x632 &  x665 &  x689 &  x707 &  x752 &  x794 &  x815 &  x821 &  x869 &  x935 &  x971 &  x983 &  x1010 &  x1037 &  x1052 &  x1118 & ~x72 & ~x73 & ~x111 & ~x261 & ~x435 & ~x513 & ~x627 & ~x666 & ~x705 & ~x1014;
assign c274 =  x11 &  x101 &  x107 &  x122 &  x149 &  x194 &  x218 &  x461 &  x488 &  x494 &  x521 &  x536 &  x539 &  x608 &  x698 &  x710 &  x779 &  x893 &  x977 &  x998 &  x1022 &  x1076 &  x1097 &  x1106 & ~x54 & ~x729 & ~x807 & ~x810 & ~x850 & ~x885 & ~x888 & ~x999 & ~x1020 & ~x1038 & ~x1059;
assign c276 =  x430 &  x502 &  x503 &  x579 &  x605 &  x749 &  x908 &  x1115 & ~x531 & ~x669 & ~x744 & ~x745;
assign c278 =  x41 &  x47 &  x146 &  x200 &  x242 &  x305 &  x331 &  x341 &  x370 &  x435 &  x436 &  x472 &  x475 &  x478 &  x548 &  x662 &  x695 &  x791 &  x839 &  x878 &  x881 &  x1076 & ~x429 & ~x882 & ~x1038;
assign c280 =  x500 &  x572 &  x640 &  x756 &  x795 &  x874 &  x1066 &  x1069 &  x1102 & ~x744 & ~x804;
assign c282 =  x3 &  x42 &  x43 &  x164 &  x173 &  x185 &  x194 &  x345 &  x365 &  x404 &  x424 &  x491 &  x502 &  x548 &  x623 &  x692 &  x761 &  x764 &  x776 &  x848 &  x874 &  x977 & ~x627 & ~x666 & ~x705;
assign c284 =  x11 &  x640 &  x1043 & ~x456 & ~x496 & ~x534 & ~x573 & ~x846 & ~x861 & ~x885 & ~x924 & ~x1041 & ~x1080 & ~x1119;
assign c286 =  x8 &  x20 &  x38 &  x68 &  x104 &  x113 &  x155 &  x159 &  x160 &  x167 &  x188 &  x199 &  x200 &  x230 &  x238 &  x260 &  x314 &  x317 &  x320 &  x374 &  x398 &  x419 &  x500 &  x512 &  x545 &  x557 &  x563 &  x605 &  x635 &  x641 &  x656 &  x689 &  x722 &  x746 &  x806 &  x836 &  x860 &  x917 &  x947 &  x950 &  x953 &  x956 &  x977 &  x986 &  x1016 &  x1019 &  x1106 & ~x66 & ~x105 & ~x183 & ~x184 & ~x222 & ~x223 & ~x261 & ~x300 & ~x375 & ~x1119;
assign c288 =  x710 &  x771 &  x775 &  x796 &  x814 &  x835 &  x853 &  x874 &  x913 &  x1030 &  x1073 & ~x480 & ~x519 & ~x675;
assign c290 =  x14 &  x35 &  x185 &  x206 &  x287 &  x338 &  x494 &  x524 &  x599 &  x635 &  x680 &  x776 &  x796 &  x980 &  x983 & ~x402 & ~x442 & ~x481 & ~x519 & ~x531 & ~x558 & ~x570 & ~x627 & ~x666 & ~x744 & ~x823 & ~x862;
assign c292 =  x77 &  x341 &  x389 &  x476 &  x503 &  x521 &  x548 &  x680 &  x803 &  x965 & ~x103 & ~x627 & ~x646;
assign c294 =  x53 &  x56 &  x62 &  x86 &  x104 &  x107 &  x110 &  x119 &  x140 &  x194 &  x206 &  x230 &  x236 &  x238 &  x242 &  x266 &  x277 &  x290 &  x308 &  x317 &  x323 &  x329 &  x338 &  x347 &  x371 &  x389 &  x398 &  x401 &  x428 &  x434 &  x437 &  x449 &  x455 &  x458 &  x491 &  x503 &  x521 &  x536 &  x563 &  x566 &  x575 &  x596 &  x644 &  x650 &  x662 &  x665 &  x671 &  x686 &  x713 &  x755 &  x770 &  x773 &  x803 &  x815 &  x833 &  x860 &  x920 &  x926 &  x929 &  x959 &  x962 &  x968 &  x989 &  x998 &  x1001 &  x1004 &  x1097 &  x1103 &  x1115 & ~x300 & ~x414 & ~x453 & ~x492 & ~x516 & ~x531 & ~x552 & ~x627 & ~x666 & ~x705 & ~x744 & ~x804 & ~x1014;
assign c296 =  x46 &  x159 &  x277 &  x752 &  x1040 &  x1066 & ~x261 & ~x298;
assign c298 =  x13 &  x218 &  x279 &  x318 &  x319 &  x355 &  x470 &  x512 &  x641 &  x796 &  x814 &  x835 &  x874 &  x929 &  x991 &  x1030 &  x1069;
assign c2100 =  x7 &  x17 &  x46 &  x146 &  x182 &  x194 &  x218 &  x335 &  x464 &  x503 &  x554 &  x668 &  x884 &  x890 &  x920 &  x974 &  x977 &  x989 &  x1007 &  x1019 &  x1022 &  x1037 &  x1067 &  x1079 &  x1097 & ~x651 & ~x729 & ~x958 & ~x997 & ~x1002 & ~x1035 & ~x1038 & ~x1041;
assign c2102 =  x74 &  x80 &  x86 &  x101 &  x113 &  x122 &  x131 &  x152 &  x155 &  x158 &  x188 &  x194 &  x196 &  x206 &  x215 &  x224 &  x233 &  x236 &  x242 &  x248 &  x263 &  x281 &  x293 &  x299 &  x314 &  x329 &  x362 &  x407 &  x413 &  x449 &  x452 &  x485 &  x503 &  x517 &  x554 &  x556 &  x587 &  x590 &  x608 &  x623 &  x671 &  x713 &  x722 &  x725 &  x731 &  x797 &  x800 &  x806 &  x839 &  x896 &  x905 &  x926 &  x952 &  x962 &  x965 &  x971 &  x980 &  x986 &  x1007 &  x1022 &  x1031 &  x1040 &  x1064 &  x1073 &  x1085 &  x1088 &  x1100 &  x1106 &  x1115 &  x1127 & ~x279 & ~x297 & ~x336 & ~x435 & ~x549 & ~x550 & ~x588 & ~x627;
assign c2104 =  x164 &  x194 &  x220 &  x334 &  x437 &  x439 &  x470 &  x478 &  x490 &  x517 &  x521 &  x554 &  x645 &  x695 &  x737 &  x806 &  x841 &  x857 &  x880 &  x913 &  x926 &  x974 &  x1009 &  x1127;
assign c2106 =  x176 &  x202 &  x241 &  x314 &  x404 &  x446 &  x464 &  x548 &  x689 &  x893 &  x896 &  x977 &  x1073 &  x1130 & ~x492 & ~x570 & ~x648 & ~x675 & ~x687 & ~x747 & ~x792 & ~x804 & ~x843 & ~x900 & ~x921;
assign c2108 =  x53 &  x80 &  x86 &  x101 &  x122 &  x161 &  x214 &  x365 &  x439 &  x614 &  x623 &  x716 &  x734 &  x758 &  x866 &  x887 &  x893 &  x908 &  x1058 & ~x39 & ~x234 & ~x492 & ~x570 & ~x609 & ~x630 & ~x648 & ~x687 & ~x708 & ~x726 & ~x861;
assign c2110 =  x43 &  x80 &  x176 &  x196 &  x229 &  x236 &  x272 &  x275 &  x384 &  x385 &  x424 &  x463 &  x502 &  x503 &  x518 &  x623 &  x710 &  x764 &  x839 &  x896 &  x1043 &  x1106 & ~x93 & ~x627;
assign c2112 =  x385 &  x409 &  x424 &  x448 &  x466 &  x470 &  x487 &  x505 &  x526 &  x565 &  x601 &  x640 &  x796 & ~x261 & ~x378;
assign c2114 =  x547 &  x569 &  x814 &  x835 &  x952 &  x1030 &  x1069 & ~x403 & ~x519 & ~x627 & ~x666 & ~x706;
assign c2116 =  x13 &  x56 &  x101 &  x227 &  x233 &  x323 &  x347 &  x374 &  x401 &  x416 &  x464 &  x487 &  x490 &  x503 &  x515 &  x518 &  x520 &  x529 &  x575 &  x587 &  x641 &  x643 &  x656 &  x725 &  x767 &  x872 &  x923 &  x968 &  x980 &  x1004 & ~x222 & ~x261 & ~x546 & ~x690 & ~x729;
assign c2118 =  x101 &  x659 &  x716 &  x781 &  x814 &  x852 &  x853 &  x891 &  x892 &  x962 & ~x651 & ~x690 & ~x864 & ~x1017;
assign c2120 =  x14 &  x17 &  x29 &  x44 &  x83 &  x89 &  x92 &  x110 &  x116 &  x122 &  x128 &  x134 &  x143 &  x149 &  x155 &  x173 &  x182 &  x191 &  x233 &  x236 &  x245 &  x248 &  x254 &  x266 &  x281 &  x296 &  x317 &  x341 &  x344 &  x350 &  x355 &  x359 &  x362 &  x383 &  x392 &  x401 &  x407 &  x419 &  x446 &  x449 &  x458 &  x461 &  x476 &  x491 &  x503 &  x506 &  x509 &  x533 &  x551 &  x554 &  x569 &  x572 &  x578 &  x584 &  x587 &  x590 &  x596 &  x599 &  x614 &  x623 &  x629 &  x635 &  x638 &  x647 &  x662 &  x677 &  x683 &  x695 &  x698 &  x752 &  x761 &  x764 &  x776 &  x779 &  x794 &  x800 &  x803 &  x812 &  x818 &  x848 &  x851 &  x857 &  x860 &  x863 &  x893 &  x911 &  x923 &  x929 &  x947 &  x956 &  x962 &  x968 &  x971 &  x983 &  x1007 &  x1010 &  x1013 &  x1016 &  x1034 &  x1046 &  x1049 &  x1067 &  x1097 &  x1100 &  x1106 & ~x261 & ~x301 & ~x339 & ~x340 & ~x375 & ~x378 & ~x414 & ~x453 & ~x456 & ~x492 & ~x531 & ~x687 & ~x744;
assign c2122 =  x23 &  x38 &  x83 &  x104 &  x110 &  x124 &  x128 &  x131 &  x155 &  x163 &  x185 &  x201 &  x230 &  x281 &  x356 &  x374 &  x386 &  x446 &  x461 &  x521 &  x565 &  x614 &  x650 &  x658 &  x668 &  x725 &  x731 &  x740 &  x764 &  x809 &  x814 &  x827 &  x893 &  x968 &  x971 &  x1001 &  x1052 &  x1055 &  x1070 &  x1105;
assign c2124 =  x23 &  x26 &  x35 &  x41 &  x65 &  x80 &  x92 &  x110 &  x122 &  x131 &  x160 &  x188 &  x203 &  x235 &  x251 &  x275 &  x281 &  x287 &  x293 &  x317 &  x323 &  x335 &  x341 &  x350 &  x359 &  x371 &  x383 &  x386 &  x395 &  x422 &  x431 &  x448 &  x452 &  x466 &  x487 &  x494 &  x502 &  x503 &  x505 &  x526 &  x541 &  x545 &  x554 &  x565 &  x572 &  x604 &  x608 &  x632 &  x635 &  x643 &  x665 &  x680 &  x695 &  x707 &  x716 &  x722 &  x725 &  x743 &  x776 &  x779 &  x782 &  x797 &  x799 &  x842 &  x845 &  x854 &  x863 &  x875 &  x884 &  x914 &  x929 &  x941 &  x965 &  x977 &  x980 &  x989 &  x995 &  x1007 &  x1013 &  x1022 &  x1040 &  x1052 &  x1055 &  x1073 &  x1076 &  x1094 &  x1109 & ~x588 & ~x729;
assign c2126 =  x26 &  x53 &  x62 &  x101 &  x146 &  x188 &  x215 &  x239 &  x257 &  x281 &  x347 &  x359 &  x365 &  x385 &  x401 &  x404 &  x424 &  x428 &  x437 &  x487 &  x490 &  x520 &  x526 &  x533 &  x565 &  x587 &  x599 &  x635 &  x643 &  x673 &  x710 &  x712 &  x722 &  x749 &  x872 &  x923 &  x962 &  x983 &  x1010 &  x1043 &  x1049 &  x1121 &  x1127 &  x1130 & ~x429 & ~x906;
assign c2128 =  x68 &  x80 &  x92 &  x113 &  x125 &  x134 &  x158 &  x266 &  x293 &  x371 &  x389 &  x416 &  x431 &  x536 &  x569 &  x614 &  x620 &  x695 &  x710 &  x764 &  x857 &  x974 &  x1070 &  x1100 & ~x480 & ~x519 & ~x570 & ~x609 & ~x648 & ~x675 & ~x687 & ~x747 & ~x792 & ~x804 & ~x843 & ~x870 & ~x882 & ~x909 & ~x1011 & ~x1056 & ~x1089;
assign c2130 =  x113 &  x218 &  x239 &  x370 &  x403 &  x409 &  x415 &  x454 &  x487 &  x493 &  x526 &  x532 &  x560 &  x565 &  x980 &  x1034 &  x1048 & ~x282 & ~x321 & ~x429 & ~x546 & ~x585 & ~x729 & ~x807 & ~x846 & ~x885;
assign c2132 =  x8 &  x11 &  x44 &  x50 &  x116 &  x122 &  x137 &  x146 &  x158 &  x173 &  x185 &  x197 &  x202 &  x241 &  x316 &  x347 &  x394 &  x422 &  x452 &  x479 &  x508 &  x515 &  x521 &  x548 &  x554 &  x583 &  x596 &  x605 &  x622 &  x644 &  x661 &  x668 &  x710 &  x716 &  x728 &  x739 &  x746 &  x794 &  x860 &  x872 &  x896 &  x911 &  x917 &  x935 &  x947 &  x965 &  x977 &  x989 &  x995 &  x1031 &  x1064 &  x1076 &  x1094 &  x1106 & ~x234 & ~x534 & ~x573 & ~x744 & ~x783;
assign c2134 =  x409 &  x475 &  x587 &  x773 &  x908 &  x931 &  x1040 &  x1048 & ~x282 & ~x429 & ~x729 & ~x843 & ~x903 & ~x921 & ~x1038;
assign c2136 = ~x15 & ~x54 & ~x72 & ~x73 & ~x111 & ~x261 & ~x340 & ~x379 & ~x418 & ~x729;
assign c2138 =  x269 &  x541 &  x619 &  x695 &  x796 & ~x339 & ~x378 & ~x417 & ~x418 & ~x456 & ~x630 & ~x669 & ~x708;
assign c2140 =  x17 &  x44 &  x65 &  x68 &  x107 &  x155 &  x170 &  x200 &  x239 &  x260 &  x277 &  x283 &  x311 &  x314 &  x316 &  x353 &  x356 &  x395 &  x419 &  x452 &  x497 &  x527 &  x542 &  x584 &  x674 &  x704 &  x740 &  x806 &  x818 &  x872 &  x875 &  x914 &  x950 &  x959 &  x980 &  x1064 &  x1070 &  x1076 &  x1082 &  x1094 &  x1103 &  x1118 & ~x300 & ~x396 & ~x474 & ~x588 & ~x606 & ~x627 & ~x705 & ~x744 & ~x786;
assign c2142 =  x32 &  x122 &  x227 &  x407 &  x503 &  x521 &  x839 & ~x156 & ~x402 & ~x441 & ~x480 & ~x531 & ~x648 & ~x675 & ~x687 & ~x708 & ~x726 & ~x765 & ~x792 & ~x861 & ~x870 & ~x909;
assign c2144 =  x38 &  x47 &  x71 &  x80 &  x83 &  x92 &  x107 &  x110 &  x122 &  x140 &  x146 &  x170 &  x227 &  x233 &  x236 &  x260 &  x266 &  x272 &  x284 &  x299 &  x302 &  x341 &  x347 &  x365 &  x377 &  x401 &  x437 &  x439 &  x446 &  x512 &  x518 &  x521 &  x527 &  x560 &  x566 &  x608 &  x614 &  x623 &  x632 &  x671 &  x680 &  x725 &  x827 &  x866 &  x884 &  x896 &  x920 &  x923 &  x941 &  x944 &  x950 &  x956 &  x968 &  x985 &  x989 &  x1022 &  x1023 &  x1031 &  x1037 &  x1043 &  x1063 &  x1097 &  x1100 &  x1102 &  x1103 &  x1109 &  x1115 & ~x1038 & ~x1083 & ~x1084;
assign c2146 =  x5 &  x8 &  x32 &  x41 &  x50 &  x74 &  x80 &  x101 &  x107 &  x113 &  x116 &  x134 &  x170 &  x173 &  x185 &  x203 &  x218 &  x230 &  x233 &  x239 &  x245 &  x260 &  x272 &  x275 &  x283 &  x287 &  x293 &  x299 &  x305 &  x311 &  x316 &  x320 &  x338 &  x347 &  x350 &  x352 &  x353 &  x356 &  x386 &  x395 &  x430 &  x431 &  x446 &  x458 &  x470 &  x473 &  x476 &  x503 &  x506 &  x527 &  x547 &  x551 &  x554 &  x557 &  x578 &  x593 &  x596 &  x599 &  x601 &  x614 &  x625 &  x632 &  x640 &  x641 &  x650 &  x656 &  x659 &  x662 &  x671 &  x677 &  x689 &  x710 &  x719 &  x746 &  x761 &  x767 &  x779 &  x782 &  x818 &  x821 &  x836 &  x851 &  x878 &  x887 &  x920 &  x929 &  x938 &  x953 &  x956 &  x962 &  x971 &  x977 &  x980 &  x992 &  x998 &  x1004 &  x1010 &  x1028 &  x1046 &  x1064 &  x1073 &  x1079 &  x1085 &  x1088 &  x1106 &  x1109 &  x1115 &  x1130 & ~x231 & ~x324 & ~x363 & ~x402 & ~x441 & ~x480 & ~x519 & ~x705 & ~x744 & ~x822;
assign c2148 =  x32 &  x80 &  x104 &  x116 &  x128 &  x179 &  x191 &  x200 &  x227 &  x245 &  x251 &  x254 &  x275 &  x283 &  x296 &  x299 &  x302 &  x353 &  x368 &  x437 &  x587 &  x590 &  x596 &  x601 &  x623 &  x640 &  x650 &  x674 &  x749 &  x752 &  x760 &  x761 &  x767 &  x769 &  x782 &  x796 &  x799 &  x800 &  x821 &  x833 &  x838 &  x866 &  x868 &  x874 &  x893 &  x913 &  x917 &  x929 &  x938 &  x952 &  x974 &  x998 &  x1016 &  x1052 &  x1102 &  x1108 & ~x492 & ~x531;
assign c2150 =  x839 & ~x111 & ~x171 & ~x327 & ~x363 & ~x414 & ~x588 & ~x589 & ~x627;
assign c2152 =  x14 &  x20 &  x29 &  x38 &  x47 &  x92 &  x101 &  x104 &  x113 &  x122 &  x131 &  x158 &  x161 &  x176 &  x182 &  x188 &  x191 &  x206 &  x218 &  x221 &  x269 &  x320 &  x323 &  x326 &  x338 &  x358 &  x359 &  x380 &  x419 &  x428 &  x436 &  x439 &  x446 &  x479 &  x497 &  x509 &  x554 &  x563 &  x584 &  x626 &  x653 &  x662 &  x665 &  x674 &  x701 &  x716 &  x722 &  x728 &  x734 &  x746 &  x749 &  x755 &  x824 &  x857 &  x893 &  x923 &  x947 &  x962 &  x974 &  x980 &  x989 &  x1010 &  x1025 &  x1094 &  x1100 &  x1109 & ~x429 & ~x540 & ~x675 & ~x714 & ~x753 & ~x792 & ~x864 & ~x978 & ~x1026;
assign c2154 =  x277 &  x467 & ~x226 & ~x261 & ~x298 & ~x336 & ~x414 & ~x453 & ~x627 & ~x666;
assign c2156 =  x14 &  x101 &  x122 &  x176 &  x194 &  x218 &  x230 &  x233 &  x319 &  x335 &  x464 &  x503 &  x587 &  x625 &  x695 &  x839 &  x896 &  x962 &  x968 &  x1013 &  x1118 & ~x234 & ~x558 & ~x630 & ~x669 & ~x675 & ~x708 & ~x747 & ~x753 & ~x786 & ~x792 & ~x825 & ~x864 & ~x909 & ~x978;
assign c2158 =  x409 &  x485 &  x517 &  x1109 & ~x12 & ~x285 & ~x807 & ~x1017 & ~x1089;
assign c2160 =  x59 &  x233 &  x521 &  x695 &  x796 &  x835 &  x1106 & ~x453 & ~x492 & ~x495 & ~x516 & ~x531 & ~x633 & ~x648 & ~x687 & ~x804;
assign c2162 =  x1097 & ~x580 & ~x676 & ~x792;
assign c2164 =  x11 &  x14 &  x62 &  x68 &  x101 &  x104 &  x113 &  x125 &  x143 &  x155 &  x158 &  x163 &  x170 &  x200 &  x233 &  x240 &  x241 &  x244 &  x277 &  x281 &  x283 &  x284 &  x293 &  x299 &  x322 &  x326 &  x335 &  x341 &  x361 &  x371 &  x392 &  x401 &  x413 &  x428 &  x430 &  x431 &  x443 &  x494 &  x497 &  x503 &  x539 &  x545 &  x566 &  x587 &  x611 &  x623 &  x644 &  x650 &  x656 &  x659 &  x668 &  x686 &  x710 &  x713 &  x716 &  x728 &  x737 &  x800 &  x827 &  x839 &  x854 &  x890 &  x893 &  x902 &  x905 &  x929 &  x956 &  x974 &  x989 &  x1022 &  x1037 &  x1043 &  x1058 &  x1076 &  x1097 &  x1106 & ~x705 & ~x744 & ~x822 & ~x861;
assign c2166 =  x11 &  x23 &  x80 &  x113 &  x122 &  x170 &  x173 &  x209 &  x215 &  x233 &  x248 &  x254 &  x314 &  x331 &  x335 &  x373 &  x395 &  x403 &  x431 &  x442 &  x448 &  x475 &  x482 &  x487 &  x520 &  x526 &  x565 &  x590 &  x604 &  x607 &  x643 &  x644 &  x682 &  x695 &  x721 &  x725 &  x760 &  x830 &  x857 &  x893 &  x932 &  x1097 &  x1106 & ~x321 & ~x468;
assign c2168 =  x11 &  x119 &  x152 &  x361 &  x373 &  x412 &  x451 &  x607 &  x622 &  x661 &  x757 &  x763 &  x812 &  x1037 &  x1043 &  x1055 & ~x381 & ~x420 & ~x459 & ~x498;
assign c2170 =  x95 &  x164 &  x236 &  x257 &  x341 &  x581 &  x962 &  x1016 &  x1130 & ~x402 & ~x480 & ~x639 & ~x648 & ~x675 & ~x786 & ~x909 & ~x960 & ~x978 & ~x1017 & ~x1038 & ~x1056;
assign c2172 =  x11 &  x53 &  x88 &  x95 &  x128 &  x170 &  x299 &  x494 &  x503 &  x526 &  x542 &  x565 &  x695 &  x756 &  x796 &  x830 &  x896 &  x908 &  x929 &  x994 &  x1076 & ~x589 & ~x627 & ~x666 & ~x744;
assign c2174 =  x20 &  x44 &  x49 &  x83 &  x98 &  x104 &  x137 &  x149 &  x167 &  x176 &  x209 &  x272 &  x299 &  x347 &  x383 &  x464 &  x476 &  x494 &  x500 &  x545 &  x596 &  x614 &  x643 &  x659 &  x668 &  x677 &  x680 &  x682 &  x699 &  x700 &  x720 &  x721 &  x759 &  x764 &  x782 &  x798 &  x799 &  x838 &  x839 &  x875 &  x876 &  x877 &  x915 &  x944 &  x954 &  x994 &  x1097;
assign c2176 =  x23 &  x65 &  x316 &  x355 &  x422 &  x449 &  x494 &  x527 &  x533 &  x563 &  x569 &  x656 &  x716 &  x767 &  x812 &  x842 &  x902 &  x926 &  x929 &  x935 & ~x39 & ~x339 & ~x453 & ~x516 & ~x531 & ~x555 & ~x570 & ~x633 & ~x648 & ~x687 & ~x726 & ~x921;
assign c2178 =  x26 &  x46 &  x149 &  x151 &  x161 &  x229 &  x317 &  x347 &  x356 &  x409 &  x413 &  x416 &  x422 &  x448 &  x487 &  x521 &  x526 &  x541 &  x548 &  x565 &  x604 &  x643 &  x682 &  x695 &  x707 &  x760 &  x779 &  x797 &  x799 &  x838 &  x896 &  x985 &  x1013 &  x1100 &  x1130;
assign c2180 =  x23 &  x32 &  x47 &  x62 &  x80 &  x86 &  x92 &  x113 &  x146 &  x158 &  x161 &  x167 &  x185 &  x188 &  x194 &  x200 &  x218 &  x227 &  x236 &  x278 &  x290 &  x299 &  x314 &  x320 &  x341 &  x356 &  x364 &  x377 &  x434 &  x446 &  x470 &  x476 &  x509 &  x527 &  x569 &  x575 &  x578 &  x590 &  x596 &  x607 &  x668 &  x728 &  x734 &  x737 &  x743 &  x767 &  x773 &  x784 &  x833 &  x884 &  x893 &  x896 &  x923 &  x938 &  x947 &  x965 &  x977 &  x980 &  x983 &  x986 &  x1010 &  x1015 &  x1037 &  x1040 &  x1043 &  x1046 &  x1053 &  x1093 &  x1118 & ~x351 & ~x429 & ~x729 & ~x885 & ~x942 & ~x1038 & ~x1059;
assign c2182 =  x32 &  x395 &  x509 &  x518 &  x868 &  x899 &  x946 &  x952 &  x989 &  x991 &  x1062 &  x1069 &  x1082 &  x1093 &  x1101 &  x1102 & ~x675 & ~x978;
assign c2184 =  x2 &  x11 &  x14 &  x53 &  x71 &  x110 &  x121 &  x125 &  x140 &  x159 &  x160 &  x161 &  x170 &  x224 &  x233 &  x238 &  x242 &  x277 &  x299 &  x308 &  x344 &  x371 &  x377 &  x386 &  x401 &  x428 &  x443 &  x461 &  x464 &  x509 &  x512 &  x562 &  x593 &  x599 &  x605 &  x617 &  x629 &  x635 &  x638 &  x640 &  x641 &  x665 &  x671 &  x674 &  x683 &  x689 &  x692 &  x701 &  x710 &  x725 &  x740 &  x758 &  x782 &  x791 &  x845 &  x854 &  x878 &  x914 &  x956 &  x977 &  x1004 &  x1037 &  x1043 &  x1066 &  x1100 &  x1104 &  x1105 &  x1112 &  x1124 & ~x375 & ~x414;
assign c2186 =  x101 &  x113 &  x265 &  x308 &  x401 &  x536 &  x581 &  x677 &  x788 &  x878 &  x881 &  x1058 & ~x93 & ~x99 & ~x339 & ~x390 & ~x495 & ~x573 & ~x613 & ~x651 & ~x652 & ~x690 & ~x729 & ~x807 & ~x885 & ~x903;
assign c2188 =  x122 &  x263 &  x325 &  x371 &  x410 &  x478 &  x503 &  x536 &  x667 &  x800 &  x866 &  x962 & ~x273 & ~x429 & ~x807 & ~x846 & ~x882 & ~x885 & ~x924 & ~x1020 & ~x1038;
assign c2190 =  x394 &  x656 &  x818 &  x830 &  x941 &  x1013 &  x1016 &  x1019 & ~x156 & ~x492 & ~x531 & ~x570 & ~x571 & ~x633 & ~x648 & ~x744 & ~x882;
assign c2192 =  x2 &  x11 &  x14 &  x20 &  x23 &  x44 &  x83 &  x86 &  x98 &  x101 &  x104 &  x110 &  x113 &  x122 &  x131 &  x137 &  x146 &  x160 &  x176 &  x194 &  x197 &  x199 &  x203 &  x206 &  x212 &  x221 &  x224 &  x227 &  x233 &  x235 &  x257 &  x260 &  x272 &  x275 &  x278 &  x302 &  x311 &  x313 &  x329 &  x335 &  x347 &  x350 &  x352 &  x359 &  x371 &  x385 &  x392 &  x395 &  x407 &  x423 &  x424 &  x437 &  x446 &  x452 &  x455 &  x497 &  x500 &  x502 &  x503 &  x512 &  x518 &  x539 &  x541 &  x551 &  x554 &  x560 &  x566 &  x584 &  x587 &  x608 &  x614 &  x619 &  x623 &  x632 &  x638 &  x647 &  x656 &  x662 &  x671 &  x677 &  x707 &  x710 &  x713 &  x718 &  x725 &  x734 &  x749 &  x755 &  x757 &  x764 &  x770 &  x773 &  x812 &  x833 &  x839 &  x842 &  x845 &  x848 &  x851 &  x857 &  x866 &  x872 &  x887 &  x902 &  x923 &  x929 &  x962 &  x968 &  x974 &  x977 &  x992 &  x995 &  x1007 &  x1016 &  x1031 &  x1061 &  x1076 &  x1097 &  x1103 &  x1106 &  x1109 &  x1118 & ~x207 & ~x246 & ~x627 & ~x666 & ~x705 & ~x706 & ~x783 & ~x861;
assign c2194 =  x250 &  x373 &  x479 &  x716 &  x848 &  x968 &  x1048 &  x1093 &  x1097 & ~x18 & ~x687 & ~x882 & ~x921 & ~x1000 & ~x1038 & ~x1039 & ~x1077;
assign c2196 =  x14 &  x31 &  x80 &  x92 &  x142 &  x275 &  x319 &  x358 &  x395 &  x572 &  x635 &  x770 &  x814 &  x835 &  x845 &  x854 &  x872 &  x874 &  x892 &  x896 &  x913 &  x952 &  x974 &  x991 &  x1030 &  x1069 &  x1103 &  x1108 & ~x675 & ~x753;
assign c2198 =  x5 &  x8 &  x17 &  x31 &  x74 &  x77 &  x146 &  x158 &  x167 &  x181 &  x182 &  x187 &  x191 &  x194 &  x220 &  x266 &  x272 &  x290 &  x314 &  x332 &  x350 &  x413 &  x449 &  x455 &  x464 &  x488 &  x494 &  x548 &  x560 &  x614 &  x668 &  x698 &  x713 &  x728 &  x737 &  x743 &  x755 &  x764 &  x779 &  x806 &  x824 &  x845 &  x857 &  x1016 &  x1048 &  x1073 &  x1087 & ~x1020 & ~x1059 & ~x1060;
assign c2200 =  x8 &  x14 &  x17 &  x56 &  x89 &  x101 &  x122 &  x143 &  x155 &  x158 &  x200 &  x221 &  x236 &  x269 &  x272 &  x329 &  x338 &  x371 &  x380 &  x392 &  x416 &  x419 &  x422 &  x424 &  x446 &  x449 &  x455 &  x482 &  x566 &  x569 &  x587 &  x629 &  x640 &  x641 &  x644 &  x671 &  x734 &  x740 &  x755 &  x764 &  x836 &  x839 &  x851 &  x908 &  x914 &  x923 &  x947 &  x968 &  x986 &  x992 &  x1055 &  x1066 &  x1067 &  x1070 &  x1085 &  x1124 & ~x66 & ~x105 & ~x183 & ~x184 & ~x222 & ~x261 & ~x858 & ~x1074;
assign c2202 =  x551 &  x956 & ~x9 & ~x48 & ~x480 & ~x528 & ~x747 & ~x786 & ~x798 & ~x825 & ~x864 & ~x909 & ~x954 & ~x1017;
assign c2204 =  x53 &  x146 &  x236 &  x278 &  x302 &  x770 &  x785 &  x815 &  x989 &  x1109 & ~x249 & ~x327 & ~x366 & ~x456 & ~x534 & ~x570 & ~x687 & ~x766 & ~x804 & ~x1057;
assign c2206 =  x2 &  x119 &  x236 &  x335 &  x701 & ~x0 & ~x33 & ~x39 & ~x72 & ~x414 & ~x453 & ~x492 & ~x531 & ~x570 & ~x648 & ~x687 & ~x744 & ~x786 & ~x1035;
assign c2208 =  x44 &  x68 &  x80 &  x110 &  x113 &  x200 &  x238 &  x239 &  x251 &  x277 &  x368 &  x374 &  x419 &  x497 &  x502 &  x509 &  x521 &  x527 &  x602 &  x640 &  x674 &  x680 &  x691 &  x695 &  x716 &  x773 &  x791 &  x796 &  x812 &  x827 &  x835 &  x857 &  x860 &  x962 &  x1004 &  x1010 &  x1052 &  x1091 &  x1118 & ~x207 & ~x285 & ~x324 & ~x363 & ~x402 & ~x597 & ~x627 & ~x666 & ~x705 & ~x744;
assign c2210 =  x11 &  x44 &  x74 &  x116 &  x121 &  x127 &  x160 &  x212 &  x218 &  x274 &  x313 &  x356 &  x428 &  x443 &  x455 &  x464 &  x485 &  x548 &  x560 &  x566 &  x692 &  x695 &  x719 &  x728 &  x740 &  x746 &  x977 &  x986 &  x989 &  x994 &  x1016 &  x1037 &  x1058 &  x1067 &  x1072 &  x1118 & ~x187 & ~x226 & ~x279 & ~x588 & ~x627 & ~x666 & ~x705 & ~x744 & ~x783;
assign c2212 =  x230 &  x250 &  x362 &  x410 &  x464 &  x814 &  x856 &  x935 &  x952 &  x991 &  x1093 &  x1097 & ~x675 & ~x726 & ~x804 & ~x843 & ~x882;
assign c2214 =  x160 &  x834 &  x956 &  x1102 &  x1104;
assign c2216 =  x491 &  x839 & ~x39 & ~x268 & ~x301 & ~x492 & ~x786;
assign c2218 =  x74 &  x389 & ~x234 & ~x480 & ~x669 & ~x675 & ~x687 & ~x747 & ~x753 & ~x792 & ~x804 & ~x940;
assign c2220 =  x67 &  x178 &  x200 &  x217 &  x256 &  x314 &  x334 &  x407 &  x475 &  x548 &  x813 &  x852 &  x853 &  x952 &  x1009 &  x1087 &  x1093 &  x1109 & ~x675;
assign c2222 =  x77 &  x155 &  x164 &  x197 &  x206 &  x271 &  x479 &  x500 &  x539 &  x611 &  x631 &  x644 &  x668 &  x728 &  x760 &  x851 &  x872 &  x896 &  x944 &  x1106 & ~x351 & ~x510 & ~x586 & ~x624 & ~x625 & ~x885 & ~x924 & ~x1035 & ~x1041;
assign c2224 =  x80 &  x191 &  x211 &  x233 &  x250 &  x319 &  x436 &  x503 &  x554 &  x775 &  x813 &  x814 &  x852 &  x891 &  x931 &  x952 &  x956 &  x962 &  x980 &  x991 &  x1009 &  x1030 &  x1069 &  x1108 & ~x675;
assign c2226 =  x116 &  x137 &  x173 &  x218 &  x251 &  x281 &  x296 &  x299 &  x428 &  x475 &  x512 &  x521 &  x572 &  x716 &  x719 &  x745 &  x749 &  x833 &  x878 &  x896 &  x899 &  x1001 &  x1061 &  x1070 &  x1082 &  x1093 &  x1109 &  x1124 & ~x753 & ~x792 & ~x837 & ~x909 & ~x981 & ~x1096;
assign c2228 =  x38 &  x68 &  x113 &  x122 &  x146 &  x152 &  x166 &  x167 &  x170 &  x182 &  x191 &  x205 &  x212 &  x254 &  x263 &  x274 &  x275 &  x311 &  x314 &  x317 &  x320 &  x326 &  x341 &  x352 &  x374 &  x383 &  x398 &  x407 &  x416 &  x422 &  x428 &  x434 &  x449 &  x458 &  x464 &  x482 &  x506 &  x527 &  x530 &  x539 &  x548 &  x554 &  x569 &  x578 &  x584 &  x605 &  x620 &  x623 &  x629 &  x656 &  x665 &  x671 &  x692 &  x710 &  x713 &  x716 &  x788 &  x791 &  x830 &  x839 &  x854 &  x863 &  x878 &  x893 &  x899 &  x902 &  x944 &  x959 &  x962 &  x965 &  x983 &  x988 &  x989 &  x1010 &  x1019 &  x1028 &  x1031 &  x1034 &  x1066 &  x1070 &  x1076 &  x1082 &  x1105 & ~x375 & ~x414 & ~x435 & ~x588 & ~x627 & ~x628 & ~x666 & ~x667 & ~x705 & ~x706 & ~x744 & ~x936 & ~x975 & ~x1053;
assign c2230 =  x472 &  x548 &  x658 &  x668 &  x697 &  x814 &  x839 &  x893 & ~x516 & ~x531 & ~x570 & ~x648 & ~x687 & ~x786 & ~x954;
assign c2232 =  x5 &  x14 &  x47 &  x80 &  x83 &  x110 &  x134 &  x137 &  x197 &  x200 &  x227 &  x277 &  x281 &  x293 &  x404 &  x422 &  x431 &  x434 &  x455 &  x458 &  x479 &  x482 &  x512 &  x539 &  x557 &  x560 &  x569 &  x581 &  x584 &  x587 &  x605 &  x680 &  x695 &  x698 &  x728 &  x743 &  x773 &  x788 &  x830 &  x863 &  x878 &  x893 &  x905 &  x911 &  x914 &  x962 &  x968 &  x1019 &  x1037 &  x1067 &  x1088 &  x1094 &  x1100 &  x1124 &  x1127 &  x1130 & ~x363 & ~x402 & ~x453 & ~x480 & ~x492 & ~x531 & ~x570 & ~x633 & ~x648 & ~x687 & ~x804 & ~x843 & ~x882;
assign c2234 =  x11 &  x14 &  x29 &  x101 &  x104 &  x107 &  x146 &  x188 &  x266 &  x290 &  x296 &  x329 &  x335 &  x341 &  x344 &  x362 &  x383 &  x415 &  x419 &  x452 &  x455 &  x467 &  x488 &  x490 &  x500 &  x506 &  x575 &  x602 &  x607 &  x623 &  x635 &  x638 &  x671 &  x695 &  x749 &  x764 &  x812 &  x872 &  x914 &  x980 &  x1022 &  x1037 &  x1043 &  x1058 &  x1064 &  x1127 & ~x810 & ~x811 & ~x882 & ~x888 & ~x921 & ~x927 & ~x1038 & ~x1059 & ~x1098;
assign c2236 =  x32 &  x35 &  x128 &  x208 &  x323 &  x370 &  x404 &  x409 &  x448 &  x467 &  x476 &  x487 &  x500 &  x527 &  x593 &  x602 &  x667 &  x707 &  x851 &  x1031 &  x1048 & ~x321 & ~x429 & ~x468 & ~x546 & ~x882 & ~x1038;
assign c2238 =  x71 &  x77 &  x95 &  x104 &  x119 &  x137 &  x143 &  x155 &  x221 &  x224 &  x236 &  x269 &  x277 &  x299 &  x305 &  x332 &  x335 &  x341 &  x347 &  x352 &  x374 &  x410 &  x443 &  x467 &  x482 &  x497 &  x509 &  x524 &  x545 &  x587 &  x593 &  x635 &  x656 &  x659 &  x662 &  x680 &  x722 &  x740 &  x812 &  x821 &  x824 &  x827 &  x830 &  x848 &  x851 &  x854 &  x857 &  x866 &  x872 &  x875 &  x881 &  x926 &  x980 &  x989 &  x1034 &  x1061 &  x1073 &  x1076 &  x1100 & ~x363 & ~x402 & ~x403 & ~x435 & ~x480 & ~x519 & ~x525 & ~x597 & ~x666 & ~x705 & ~x744 & ~x753 & ~x783;
assign c2240 =  x125 &  x215 &  x233 &  x272 &  x278 &  x281 &  x338 &  x539 &  x605 &  x623 &  x665 &  x704 &  x947 &  x962 &  x986 & ~x27 & ~x39 & ~x66 & ~x156 & ~x261 & ~x300 & ~x378 & ~x453 & ~x492 & ~x531 & ~x633 & ~x804 & ~x861 & ~x939;
assign c2242 =  x8 &  x74 &  x113 &  x197 &  x200 &  x203 &  x212 &  x224 &  x236 &  x248 &  x257 &  x272 &  x278 &  x320 &  x334 &  x341 &  x344 &  x364 &  x373 &  x376 &  x377 &  x424 &  x452 &  x475 &  x478 &  x482 &  x517 &  x521 &  x556 &  x575 &  x595 &  x617 &  x659 &  x680 &  x692 &  x710 &  x809 &  x812 &  x863 &  x874 &  x878 &  x884 &  x908 &  x911 &  x931 &  x962 &  x1022 &  x1037 &  x1046 &  x1048 &  x1070 &  x1076 &  x1087 &  x1102 &  x1112 &  x1126 & ~x429;
assign c2244 =  x41 &  x119 &  x243 &  x283 &  x544 &  x601 &  x640 &  x653 &  x796 &  x835 &  x1105 & ~x420 & ~x456 & ~x459;
assign c2246 =  x5 &  x80 &  x113 &  x188 &  x200 &  x218 &  x238 &  x277 &  x323 &  x335 &  x341 &  x353 &  x584 &  x620 &  x638 &  x692 &  x896 &  x1040 &  x1058 &  x1073 & ~x246 & ~x285 & ~x286 & ~x324 & ~x325 & ~x363 & ~x402 & ~x414 & ~x474 & ~x480 & ~x519 & ~x627 & ~x666 & ~x667 & ~x706 & ~x744;
assign c2248 =  x44 &  x92 &  x116 &  x125 &  x128 &  x143 &  x191 &  x227 &  x254 &  x299 &  x310 &  x371 &  x377 &  x383 &  x398 &  x403 &  x446 &  x524 &  x530 &  x539 &  x569 &  x617 &  x626 &  x692 &  x695 &  x710 &  x716 &  x725 &  x758 &  x824 &  x833 &  x848 &  x893 &  x956 &  x962 &  x965 &  x989 &  x1076 &  x1115 &  x1121 & ~x39 & ~x79 & ~x118 & ~x156 & ~x183 & ~x339 & ~x417 & ~x495 & ~x534 & ~x573 & ~x729 & ~x807 & ~x885;
assign c2250 =  x122 &  x410 &  x677 &  x917 &  x989 & ~x27 & ~x66 & ~x72 & ~x78 & ~x111 & ~x339 & ~x807 & ~x846 & ~x885 & ~x886 & ~x924 & ~x925 & ~x999 & ~x1002 & ~x1038;
assign c2252 =  x26 &  x475 &  x509 &  x545 &  x575 &  x689 &  x698 &  x745 &  x776 &  x824 &  x947 &  x1007 &  x1009 &  x1093 & ~x429 & ~x882 & ~x903 & ~x1000 & ~x1038 & ~x1039 & ~x1078 & ~x1117;
assign c2254 =  x101 &  x116 &  x122 &  x155 &  x233 &  x260 &  x272 &  x308 &  x335 &  x365 &  x398 &  x467 &  x503 &  x539 &  x557 &  x566 &  x605 &  x623 &  x638 &  x683 &  x695 &  x710 &  x887 &  x902 &  x938 &  x962 &  x989 &  x1010 &  x1040 &  x1061 &  x1097 &  x1100 & ~x0 & ~x78 & ~x117 & ~x156 & ~x570 & ~x648 & ~x669 & ~x687 & ~x708 & ~x726 & ~x747 & ~x786 & ~x825 & ~x864 & ~x903 & ~x978 & ~x1035;
assign c2256 =  x5 &  x43 &  x56 &  x68 &  x92 &  x95 &  x110 &  x127 &  x134 &  x139 &  x173 &  x178 &  x185 &  x212 &  x233 &  x236 &  x272 &  x277 &  x290 &  x329 &  x365 &  x371 &  x374 &  x377 &  x395 &  x428 &  x458 &  x490 &  x494 &  x500 &  x503 &  x506 &  x521 &  x527 &  x548 &  x556 &  x560 &  x563 &  x587 &  x595 &  x599 &  x617 &  x620 &  x641 &  x671 &  x682 &  x683 &  x752 &  x770 &  x863 &  x869 &  x877 &  x896 &  x902 &  x952 &  x974 &  x991 &  x998 &  x1007 &  x1019 &  x1022 &  x1040 &  x1103 &  x1115;
assign c2258 =  x43 &  x46 &  x59 &  x65 &  x81 &  x85 &  x98 &  x120 &  x159 &  x160 &  x179 &  x194 &  x197 &  x199 &  x274 &  x275 &  x320 &  x335 &  x365 &  x371 &  x503 &  x539 &  x629 &  x650 &  x725 &  x896 &  x914 &  x1004 &  x1019 &  x1028 &  x1037 &  x1106 & ~x1074;
assign c2260 =  x3 &  x4 &  x11 &  x32 &  x43 &  x80 &  x98 &  x101 &  x116 &  x160 &  x164 &  x233 &  x257 &  x305 &  x308 &  x314 &  x380 &  x395 &  x506 &  x512 &  x536 &  x548 &  x578 &  x593 &  x599 &  x620 &  x632 &  x650 &  x695 &  x701 &  x716 &  x752 &  x794 &  x803 &  x845 &  x860 &  x878 &  x947 &  x962 &  x1046 &  x1067 &  x1088 &  x1106 &  x1109 & ~x57 & ~x96 & ~x135 & ~x174 & ~x291 & ~x321 & ~x330 & ~x429 & ~x468;
assign c2262 =  x352 &  x716 &  x788 &  x839 & ~x363 & ~x402 & ~x456 & ~x480 & ~x708 & ~x765 & ~x786 & ~x804 & ~x870 & ~x909;
assign c2264 =  x159 &  x160 &  x212 &  x654 &  x677 &  x1100 & ~x1035;
assign c2266 =  x8 &  x38 &  x113 &  x128 &  x191 &  x200 &  x209 &  x233 &  x254 &  x325 &  x331 &  x362 &  x364 &  x365 &  x370 &  x398 &  x409 &  x440 &  x485 &  x551 &  x581 &  x587 &  x629 &  x677 &  x686 &  x833 &  x841 &  x863 &  x905 &  x908 &  x911 &  x962 &  x1004 &  x1076 &  x1097 & ~x429 & ~x885 & ~x903 & ~x924 & ~x1038;
assign c2268 =  x32 &  x44 &  x101 &  x104 &  x140 &  x167 &  x188 &  x209 &  x239 &  x244 &  x245 &  x248 &  x269 &  x277 &  x293 &  x352 &  x374 &  x398 &  x404 &  x422 &  x425 &  x440 &  x452 &  x455 &  x482 &  x506 &  x509 &  x530 &  x536 &  x554 &  x569 &  x584 &  x599 &  x620 &  x623 &  x632 &  x641 &  x692 &  x704 &  x716 &  x755 &  x785 &  x839 &  x860 &  x872 &  x920 &  x968 &  x980 &  x1001 &  x1013 &  x1016 &  x1028 &  x1031 &  x1040 &  x1049 &  x1052 &  x1055 &  x1058 &  x1070 & ~x474 & ~x531 & ~x627 & ~x705 & ~x744 & ~x747 & ~x783 & ~x823 & ~x861 & ~x862;
assign c2270 =  x7 &  x35 &  x164 &  x209 &  x278 &  x299 &  x302 &  x329 &  x374 &  x424 &  x452 &  x542 &  x569 &  x640 &  x662 &  x671 &  x686 &  x691 &  x692 &  x713 &  x740 &  x776 &  x815 &  x854 &  x874 &  x896 &  x920 &  x926 &  x977 &  x986 &  x1001 &  x1007 &  x1016 &  x1052 &  x1079 &  x1112 &  x1121 &  x1128;
assign c2272 =  x29 &  x47 &  x65 &  x101 &  x146 &  x158 &  x209 &  x220 &  x227 &  x236 &  x263 &  x265 &  x281 &  x286 &  x325 &  x368 &  x436 &  x550 &  x581 &  x623 &  x629 &  x668 &  x716 &  x761 &  x763 &  x776 &  x802 &  x839 &  x841 &  x848 &  x896 &  x974 &  x989 & ~x882 & ~x921 & ~x1038;
assign c2274 =  x11 &  x120 &  x466 &  x875 &  x893 & ~x148 & ~x226 & ~x510;
assign c2276 =  x46 &  x85 &  x104 &  x116 &  x131 &  x146 &  x176 &  x193 &  x217 &  x487 &  x526 &  x551 &  x565 &  x621 &  x716 &  x734 &  x764 &  x827 &  x838 &  x911 &  x1031 &  x1097 & ~x744;
assign c2278 =  x14 &  x88 &  x487 &  x502 &  x526 &  x565 &  x623 & ~x279 & ~x336 & ~x414 & ~x588 & ~x729;
assign c2280 =  x104 &  x356 &  x433 &  x500 &  x854 &  x950 &  x1022 &  x1040 & ~x234 & ~x480 & ~x519 & ~x531 & ~x648 & ~x675 & ~x687 & ~x747 & ~x753 & ~x804 & ~x870;
assign c2282 =  x43 &  x100 &  x139 &  x160 &  x217 &  x412 &  x529 &  x586 & ~x12 & ~x330 & ~x498 & ~x882;
assign c2284 =  x113 &  x160 &  x176 &  x238 &  x273 &  x277 &  x283 &  x305 &  x320 &  x350 &  x352 &  x368 &  x434 &  x503 &  x623 &  x716 &  x719 &  x725 &  x752 &  x854 &  x955 &  x994 &  x1055 &  x1097 &  x1115 & ~x357 & ~x552 & ~x588 & ~x589 & ~x627 & ~x628 & ~x666 & ~x705 & ~x744 & ~x897;
assign c2286 =  x152 &  x311 &  x527 &  x584 &  x800 &  x821 &  x848 &  x974 & ~x648 & ~x675 & ~x687 & ~x688 & ~x727 & ~x747 & ~x753 & ~x792 & ~x804 & ~x864 & ~x978 & ~x1056 & ~x1110;
assign c2288 =  x146 &  x149 &  x257 &  x680 &  x737 &  x796 &  x814 &  x839 &  x874 &  x952 &  x1030 &  x1076 & ~x363 & ~x414 & ~x453 & ~x480 & ~x597 & ~x627 & ~x666 & ~x675 & ~x705 & ~x753 & ~x909 & ~x948;
assign c2290 =  x29 &  x47 &  x74 &  x113 &  x233 &  x245 &  x317 &  x344 &  x401 &  x419 &  x485 &  x488 &  x497 &  x554 &  x608 &  x611 &  x623 &  x710 &  x761 &  x785 &  x833 &  x893 &  x968 &  x970 &  x1007 &  x1009 &  x1085 & ~x651 & ~x690 & ~x691 & ~x726 & ~x729 & ~x864 & ~x1017 & ~x1056;
assign c2292 =  x83 &  x101 &  x110 &  x113 &  x122 &  x134 &  x161 &  x176 &  x179 &  x200 &  x218 &  x233 &  x236 &  x271 &  x272 &  x293 &  x302 &  x368 &  x371 &  x404 &  x428 &  x464 &  x473 &  x476 &  x488 &  x494 &  x533 &  x536 &  x548 &  x554 &  x569 &  x587 &  x596 &  x599 &  x608 &  x617 &  x635 &  x650 &  x668 &  x686 &  x728 &  x731 &  x760 &  x785 &  x791 &  x799 &  x809 &  x854 &  x857 &  x863 &  x890 &  x893 &  x914 &  x923 &  x941 &  x947 &  x962 &  x977 &  x989 &  x1007 &  x1010 &  x1022 &  x1028 &  x1040 &  x1076 &  x1088 &  x1097 &  x1106 & ~x433 & ~x468 & ~x472 & ~x867 & ~x906 & ~x984;
assign c2294 =  x100 &  x142 &  x295 &  x475 &  x626 &  x641 &  x952 &  x991 &  x1009 &  x1014 &  x1030 &  x1094 & ~x1026;
assign c2296 =  x107 &  x113 &  x122 &  x149 &  x212 &  x251 &  x275 &  x302 &  x319 &  x325 &  x332 &  x353 &  x439 &  x476 &  x478 &  x506 &  x586 &  x587 &  x614 &  x625 &  x626 &  x659 &  x677 &  x704 &  x716 &  x719 &  x731 &  x773 &  x854 &  x899 &  x908 &  x911 &  x935 &  x1010 &  x1031 &  x1067 &  x1076 &  x1085 &  x1097 &  x1112 &  x1124 &  x1127 & ~x612 & ~x651 & ~x690 & ~x786 & ~x825 & ~x864 & ~x903;
assign c2298 =  x17 &  x53 &  x101 &  x116 &  x143 &  x170 &  x212 &  x233 &  x251 &  x274 &  x281 &  x329 &  x335 &  x374 &  x398 &  x434 &  x440 &  x446 &  x449 &  x464 &  x491 &  x497 &  x551 &  x557 &  x569 &  x596 &  x629 &  x638 &  x683 &  x710 &  x725 &  x737 &  x794 &  x830 &  x860 &  x953 &  x956 &  x1058 &  x1067 & ~x246 & ~x247 & ~x285 & ~x286 & ~x363 & ~x435 & ~x510 & ~x550 & ~x589 & ~x628 & ~x705;
assign c21 =  x702 &  x939;
assign c23 =  x961 &  x1049 & ~x352 & ~x399 & ~x891;
assign c25 =  x137 &  x152 &  x338 &  x470 &  x599 &  x644 &  x731 &  x847 &  x886 &  x964 & ~x108 & ~x654 & ~x816 & ~x933 & ~x1032;
assign c27 =  x230 &  x313 &  x513 &  x653 & ~x486 & ~x780;
assign c29 =  x421 &  x741 & ~x856 & ~x1104;
assign c211 =  x19 &  x23 &  x64 &  x421 &  x431 &  x443 &  x460 &  x535 &  x562 &  x574 &  x716 &  x737 &  x857 &  x983 &  x1061 & ~x354;
assign c213 =  x901 &  x940 &  x979 &  x1057 & ~x69 & ~x75 & ~x102 & ~x108 & ~x141 & ~x192 & ~x303;
assign c215 =  x52 &  x662 &  x943 &  x1127 & ~x315 & ~x450 & ~x615;
assign c217 = ~x484 & ~x703 & ~x898;
assign c219 =  x23 &  x223 &  x260 &  x694 &  x727 &  x812 & ~x108 & ~x252 & ~x828;
assign c221 =  x59 &  x104 &  x377 &  x464 &  x533 &  x548 &  x587 &  x590 &  x722 &  x731 &  x740 &  x797 &  x863 &  x875 &  x887 &  x940 &  x965 &  x979 &  x1018 &  x1097 &  x1100 & ~x237 & ~x315 & ~x354 & ~x477 & ~x603;
assign c223 =  x37 &  x940 & ~x159 & ~x354 & ~x891;
assign c225 =  x19 &  x148 &  x421 &  x574 &  x797 &  x958 &  x997;
assign c227 =  x610 &  x811 &  x895 & ~x504;
assign c229 =  x140 &  x197 &  x245 &  x401 &  x521 &  x608 &  x781 &  x823 &  x833 &  x901 &  x920 &  x926 &  x940 &  x983 &  x1018 &  x1043 &  x1052 &  x1057 &  x1070 & ~x159 & ~x354 & ~x795 & ~x834 & ~x933;
assign c231 =  x994 &  x1006 & ~x930;
assign c233 =  x173 &  x687 &  x748 & ~x618;
assign c235 =  x1129 & ~x42 & ~x123 & ~x213 & ~x819;
assign c237 =  x125 &  x329 &  x422 &  x509 &  x551 &  x695 &  x704 &  x710 &  x803 &  x809 &  x836 &  x920 &  x922 &  x1073 &  x1078 & ~x30 & ~x255 & ~x345;
assign c239 =  x146 &  x901 &  x1018 & ~x42 & ~x277;
assign c241 =  x592 &  x844 & ~x409 & ~x624 & ~x663 & ~x702;
assign c243 =  x312 &  x709 & ~x487;
assign c245 =  x940 &  x1018 & ~x255 & ~x826 & ~x1125;
assign c247 =  x867 & ~x234 & ~x312 & ~x354 & ~x951;
assign c249 =  x235 &  x302 &  x323 &  x344 &  x347 &  x458 &  x513 &  x524 &  x552 &  x566 &  x574 &  x587 &  x613 &  x788 &  x830 &  x866 &  x872 &  x881 &  x968 &  x1037 &  x1094 & ~x783;
assign c251 =  x16 &  x421 &  x807 &  x1039;
assign c253 =  x585 &  x833 &  x865 &  x904 & ~x354;
assign c255 =  x674 &  x932 & ~x399 & ~x699 & ~x891 & ~x930 & ~x951 & ~x969 & ~x990;
assign c257 =  x41 &  x101 &  x122 &  x182 &  x328 &  x410 &  x445 &  x470 &  x585 &  x632 &  x671 &  x710 &  x716 &  x728 &  x902 &  x958 &  x998 & ~x615 & ~x693 & ~x777 & ~x816 & ~x855;
assign c259 =  x195 &  x398 &  x616 &  x938 & ~x84 & ~x408 & ~x624 & ~x741;
assign c261 =  x64 &  x130 &  x421 &  x656 &  x904 &  x958 & ~x621;
assign c263 =  x61 &  x73 &  x421 &  x535 &  x689 &  x958 &  x965 & ~x816 & ~x1077;
assign c265 =  x11 &  x41 &  x95 &  x236 &  x413 &  x611 &  x617 &  x653 &  x668 &  x671 &  x704 &  x716 &  x901 &  x940 &  x998 &  x1031 & ~x438 & ~x477 & ~x603 & ~x693;
assign c267 =  x534 &  x847 & ~x1023;
assign c269 =  x5 &  x35 &  x223 &  x287 &  x530 &  x686 &  x692 &  x779 &  x901 &  x940 &  x953 &  x998 &  x1018 &  x1057 &  x1058 & ~x30 & ~x108 & ~x933 & ~x942;
assign c271 = ~x117 & ~x795 & ~x1086;
assign c273 =  x332 &  x443 & ~x561 & ~x601 & ~x657 & ~x858;
assign c275 =  x574 &  x827 &  x1078 & ~x84 & ~x267 & ~x423;
assign c277 =  x29 &  x134 &  x152 &  x164 &  x245 &  x332 &  x343 &  x428 &  x797 &  x839 &  x1055 & ~x42 & ~x553 & ~x609;
assign c279 =  x20 &  x140 &  x155 &  x170 &  x182 &  x233 &  x491 &  x503 &  x515 &  x542 &  x593 &  x610 &  x655 &  x767 &  x803 &  x811 &  x833 &  x836 &  x881 &  x908 &  x920 &  x1073 &  x1078 &  x1127 & ~x6 & ~x45 & ~x84 & ~x162;
assign c281 =  x628 & ~x240 & ~x405 & ~x444 & ~x696 & ~x735 & ~x813 & ~x1086;
assign c283 =  x26 &  x98 &  x134 &  x383 &  x470 &  x665 &  x715 &  x770 &  x1079 & ~x177 & ~x267 & ~x360 & ~x384 & ~x399 & ~x423 & ~x699;
assign c285 =  x95 &  x338 &  x670 &  x724 &  x766 &  x787 &  x883 & ~x828 & ~x981;
assign c287 =  x784 &  x901 & ~x159 & ~x795 & ~x1008 & ~x1047 & ~x1086;
assign c289 =  x787 &  x865 & ~x411 & ~x466 & ~x504;
assign c291 =  x2 &  x28 &  x41 &  x55 &  x88 &  x127 &  x146 &  x242 &  x262 &  x353 &  x407 &  x421 &  x428 &  x439 &  x460 &  x491 &  x527 &  x686 &  x713 &  x737 &  x881 &  x896 &  x941 &  x1070 & ~x777 & ~x816 & ~x855 & ~x1050;
assign c293 =  x79 &  x677 &  x766 &  x883 &  x961 & ~x135 & ~x186 & ~x828;
assign c295 =  x817 & ~x225 & ~x412 & ~x462;
assign c297 =  x65 &  x1018 & ~x354 & ~x471 & ~x871 & ~x1107;
assign c299 =  x340 & ~x45 & ~x108 & ~x615 & ~x738 & ~x777 & ~x894 & ~x933;
assign c2101 =  x34 &  x38 &  x112 &  x116 &  x287 &  x341 &  x421 &  x436 &  x499 &  x515 &  x542 &  x596 &  x613 &  x668 &  x835 &  x869 &  x938 &  x947 & ~x1032;
assign c2103 =  x226 &  x263 &  x371 &  x467 &  x523 &  x524 &  x530 &  x533 &  x566 &  x569 &  x641 &  x653 &  x677 &  x713 &  x790 &  x845 &  x906 &  x907 &  x1037 &  x1049 &  x1070 &  x1115 & ~x915;
assign c2105 =  x10 &  x28 &  x61 &  x92 &  x140 &  x185 &  x188 &  x242 &  x335 &  x338 &  x485 &  x518 &  x530 &  x694 &  x824 &  x896 &  x944 &  x958 &  x965 &  x986 &  x997 &  x1039 &  x1078 & ~x582;
assign c2107 =  x54 &  x613 &  x766 & ~x789;
assign c2109 =  x25 &  x52 &  x169 &  x208 &  x292 & ~x267 & ~x294 & ~x816;
assign c2111 =  x530 &  x766 &  x811 &  x817 &  x889 &  x922 &  x929 & ~x252 & ~x408 & ~x750;
assign c2113 =  x14 & ~x217 & ~x1047 & ~x1102;
assign c2115 =  x143 &  x350 &  x368 &  x422 &  x574 &  x613 &  x857 &  x925 &  x962 &  x1022 &  x1109 & ~x45 & ~x84 & ~x123 & ~x201 & ~x1023 & ~x1104;
assign c2117 =  x1020 & ~x354 & ~x877;
assign c2119 =  x23 &  x62 &  x101 &  x113 &  x116 &  x179 &  x203 &  x230 &  x272 &  x786 &  x787 &  x865 &  x887 &  x904 &  x1106 & ~x411 & ~x486;
assign c2121 =  x40 &  x41 &  x200 &  x329 &  x335 &  x395 &  x470 &  x482 &  x535 &  x611 &  x616 &  x617 &  x635 &  x680 &  x770 &  x776 &  x821 &  x878 &  x962 &  x1004 &  x1013 &  x1022 & ~x45 & ~x84 & ~x123 & ~x816 & ~x1104;
assign c2123 =  x133 &  x901 & ~x333 & ~x775;
assign c2125 =  x37 &  x343 & ~x592;
assign c2127 =  x900 & ~x709;
assign c2129 =  x77 &  x230 &  x398 &  x523 &  x605 &  x741 &  x890 &  x1130 & ~x276 & ~x315 & ~x549 & ~x910;
assign c2131 =  x315 &  x766 & ~x123 & ~x162;
assign c2133 =  x355 &  x433 &  x754 &  x910 &  x949 & ~x303 & ~x444 & ~x1008;
assign c2135 =  x301 &  x441 & ~x837;
assign c2137 =  x516 &  x1060 & ~x189 & ~x267 & ~x462 & ~x489;
assign c2139 =  x393 &  x1033 & ~x582 & ~x618;
assign c2141 =  x61 &  x259 &  x523 &  x958 &  x1021;
assign c2143 =  x706 &  x829 &  x917 & ~x559 & ~x735;
assign c2145 =  x445 &  x901 &  x940 &  x979 &  x1019 &  x1057 & ~x159 & ~x354 & ~x486;
assign c2147 =  x685 & ~x84 & ~x253 & ~x516 & ~x819;
assign c2149 =  x25 &  x130 &  x208 &  x786 &  x787 &  x904 &  x971 &  x982 &  x1052;
assign c2151 =  x28 &  x73 &  x572 &  x766 &  x805 &  x844 &  x883 &  x958 &  x1000 & ~x426;
assign c2153 =  x351 &  x997 & ~x448 & ~x1116;
assign c2155 =  x101 &  x125 &  x392 &  x585 &  x671 &  x674 &  x803 &  x812 &  x899 &  x1031 & ~x354 & ~x471 & ~x474 & ~x771 & ~x870;
assign c2157 =  x112 &  x236 &  x259 &  x262 &  x307 &  x367 &  x421 &  x613 &  x758 &  x899 &  x956 & ~x738 & ~x777;
assign c2159 =  x29 &  x146 &  x191 &  x260 &  x320 &  x421 &  x458 &  x500 &  x506 &  x569 &  x644 &  x781 &  x887 &  x901 &  x935 &  x940 &  x965 &  x968 &  x979 &  x1013 &  x1018 &  x1043 &  x1057 &  x1070 & ~x915 & ~x1029;
assign c2161 =  x191 &  x290 &  x509 &  x571 &  x616 &  x655 &  x668 &  x836 &  x850 &  x869 &  x1118 & ~x6 & ~x84 & ~x162 & ~x186;
assign c2163 =  x73 &  x460 &  x839 &  x1074 &  x1080;
assign c2165 =  x670 &  x953 & ~x240 & ~x486 & ~x990 & ~x1068;
assign c2167 =  x38 &  x77 &  x131 &  x353 &  x359 &  x365 &  x374 &  x395 &  x401 &  x574 &  x632 &  x671 &  x686 &  x695 &  x752 &  x845 &  x869 &  x920 &  x926 &  x995 &  x1007 &  x1019 &  x1034 &  x1073 &  x1085 &  x1115 & ~x751 & ~x790 & ~x829 & ~x907 & ~x945;
assign c2169 =  x883 &  x922 &  x1006 & ~x123 & ~x162 & ~x180;
assign c2171 =  x616 &  x739 &  x787 &  x817 &  x922 &  x973 & ~x387;
assign c2173 =  x249 & ~x622;
assign c2175 =  x44 &  x176 &  x254 &  x296 &  x710 &  x747 &  x845 &  x1037 & ~x486 & ~x858 & ~x1017;
assign c2177 =  x25 &  x298 &  x337 &  x376 &  x949 & ~x333 & ~x813;
assign c2179 =  x234 &  x513 & ~x447;
assign c2181 =  x23 &  x227 &  x254 &  x422 &  x470 &  x938 & ~x799 & ~x838 & ~x877 & ~x960 & ~x1071;
assign c2183 =  x5 &  x158 &  x823 &  x829 &  x1096 & ~x693 & ~x777;
assign c2185 =  x726 &  x910 &  x1084 & ~x483 & ~x819 & ~x858;
assign c2187 =  x135 &  x378;
assign c2189 =  x23 &  x817 & ~x168 & ~x328 & ~x367 & ~x672;
assign c2191 =  x440 &  x620 &  x686 &  x884 &  x953 &  x983 &  x1012 & ~x240 & ~x397 & ~x423;
assign c2193 =  x518 &  x770 & ~x3 & ~x355 & ~x993 & ~x1029;
assign c2195 =  x17 &  x29 &  x61 &  x125 &  x421 &  x653 &  x787 &  x889 &  x958 & ~x789;
assign c2197 =  x73 &  x787 &  x925 & ~x486 & ~x522 & ~x819;
assign c2199 =  x164 &  x1039 & ~x42 & ~x108 & ~x177 & ~x930;
assign c2201 =  x200 &  x260 &  x302 &  x445 &  x515 &  x722 &  x861 &  x944 &  x1056 &  x1112;
assign c2203 =  x628 &  x706 &  x960 &  x1039 &  x1045 &  x1111;
assign c2205 =  x44 &  x50 &  x113 &  x137 &  x152 &  x179 &  x188 &  x218 &  x287 &  x326 &  x383 &  x482 &  x628 &  x719 &  x959 &  x980 &  x1028 &  x1046 &  x1103 &  x1121 & ~x120 & ~x522 & ~x561 & ~x657 & ~x819;
assign c2207 =  x128 &  x278 &  x461 &  x911 &  x1021 &  x1031 &  x1043 &  x1060 & ~x204 & ~x411 & ~x423 & ~x816;
assign c2209 =  x312 &  x739 & ~x84 & ~x175;
assign c2211 =  x406 &  x507 &  x925 & ~x354 & ~x693;
assign c2213 = ~x256 & ~x309 & ~x334 & ~x576;
assign c2215 =  x262 &  x301 &  x569 &  x572 &  x617 &  x820 &  x851 &  x890 &  x1052 &  x1076 &  x1109 & ~x69 & ~x108 & ~x219 & ~x738 & ~x777 & ~x933 & ~x999 & ~x1083;
assign c2217 = ~x974;
assign c2219 = ~x339 & ~x564 & ~x661 & ~x739 & ~x816;
assign c2221 =  x754 & ~x30 & ~x126 & ~x423;
assign c2223 =  x936 &  x1017 &  x1095 & ~x510;
assign c2225 =  x29 &  x341 &  x425 &  x473 &  x500 &  x509 &  x548 &  x563 &  x617 &  x784 &  x848 &  x899 &  x901 &  x905 &  x940 &  x1016 &  x1043 &  x1058 &  x1115 & ~x3 & ~x717 & ~x756 & ~x795 & ~x834 & ~x1047;
assign c2227 =  x939 & ~x598;
assign c2229 =  x460 &  x1017 &  x1095;
assign c2231 =  x28 &  x901 &  x940 & ~x102 & ~x360 & ~x486;
assign c2233 =  x53 &  x89 &  x161 &  x191 &  x260 &  x359 &  x446 &  x494 &  x524 &  x527 &  x551 &  x572 &  x641 &  x650 &  x668 &  x671 &  x701 &  x703 &  x704 &  x722 &  x761 &  x781 &  x830 &  x839 &  x869 &  x878 &  x917 &  x937 &  x982 &  x1019 &  x1020 &  x1021 &  x1028 &  x1046 &  x1052 &  x1079 &  x1088 & ~x276 & ~x993;
assign c2235 =  x510 &  x628 &  x791 & ~x477 & ~x657;
assign c2237 =  x753 & ~x774;
assign c2239 =  x340 &  x441 & ~x553;
assign c2241 =  x1057 &  x1096 & ~x120 & ~x159 & ~x354 & ~x793;
assign c2243 =  x53 &  x71 &  x122 &  x266 &  x341 &  x485 &  x527 &  x584 &  x590 &  x686 &  x731 &  x848 &  x865 &  x904 &  x1103 & ~x45 & ~x267 & ~x423 & ~x933;
assign c2245 =  x301 &  x326 &  x367 &  x980 & ~x475 & ~x514;
assign c2247 =  x22 &  x32 &  x61 &  x73 &  x134 &  x242 &  x287 &  x290 &  x305 &  x314 &  x337 &  x343 &  x371 &  x401 &  x421 &  x422 &  x460 &  x479 &  x527 &  x566 &  x572 &  x638 &  x647 &  x659 &  x662 &  x764 &  x776 &  x800 &  x809 &  x812 &  x827 &  x833 &  x851 &  x878 &  x905 &  x1021 &  x1028 &  x1060 &  x1091 &  x1099;
assign c2249 =  x317 &  x353 &  x394 &  x452 &  x589 &  x628 &  x1006 &  x1123 & ~x741;
assign c2251 =  x164 &  x437 &  x533 &  x610 &  x616 &  x650 &  x655 &  x878 & ~x6 & ~x69 & ~x522;
assign c2253 =  x786 & ~x682;
assign c2255 =  x19 &  x25 &  x169 &  x379 &  x519;
assign c2257 =  x2 &  x197 &  x353 &  x419 &  x550 &  x563 &  x628 &  x650 &  x656 &  x791 &  x830 &  x1034 &  x1058 &  x1076 &  x1127 & ~x522 & ~x561 & ~x657 & ~x813 & ~x852 & ~x1008 & ~x1047 & ~x1083;
assign c2259 =  x634 &  x787 &  x878 &  x908 & ~x267 & ~x423 & ~x660;
assign c2261 =  x724 &  x787 &  x805 &  x844 &  x883 &  x922 & ~x348 & ~x486;
assign c2263 =  x308 &  x355 &  x648 &  x687 &  x910 & ~x303;
assign c2265 =  x25 &  x427 &  x627 &  x659 &  x1058 & ~x762 & ~x852 & ~x1086;
assign c2267 =  x585 & ~x42 & ~x400;
assign c2269 =  x41 &  x343 &  x382 &  x434 &  x479 &  x515 &  x716 &  x901 &  x922 & ~x384 & ~x423;
assign c2271 =  x513 &  x552 & ~x408 & ~x447 & ~x819;
assign c2273 =  x940 &  x1017 &  x1057 & ~x237 & ~x471;
assign c2275 =  x14 &  x89 &  x239 &  x332 &  x349 &  x388 &  x398 &  x422 &  x425 &  x427 &  x587 &  x608 &  x689 &  x734 &  x890 &  x929 &  x937 &  x940 &  x978 &  x1017 &  x1056 &  x1057 &  x1079 &  x1095;
assign c2277 =  x134 &  x155 &  x182 &  x215 &  x293 &  x353 &  x812 &  x865 &  x904 &  x953 &  x982 &  x1021 &  x1060 & ~x42 & ~x759 & ~x876;
assign c2279 =  x47 &  x312 &  x560 &  x695 &  x1058 & ~x84 & ~x258 & ~x408 & ~x828 & ~x945 & ~x1062;
assign c2281 =  x98 & ~x384 & ~x462 & ~x699 & ~x930 & ~x951 & ~x1068;
assign c2283 =  x22 &  x167 &  x346 &  x373 &  x460 &  x506 &  x737 &  x932 &  x976 &  x997 &  x1035 &  x1036 &  x1073 &  x1074 &  x1080;
assign c2285 =  x628 &  x1021 &  x1073 & ~x42 & ~x774;
assign c2287 = ~x626;
assign c2289 =  x1033 &  x1045 & ~x283 & ~x858 & ~x1102;
assign c2291 =  x148 &  x1018 &  x1056 &  x1057 & ~x471;
assign c2293 =  x549 &  x627 & ~x724;
assign c2295 =  x900 & ~x709;
assign c2297 =  x301 &  x546 & ~x700 & ~x739;
assign c2299 =  x23 &  x143 &  x355 &  x628 &  x883 &  x910 &  x922 &  x949 &  x998 &  x1051 &  x1090 &  x1123;
assign c30 =  x11 &  x17 &  x47 &  x53 &  x68 &  x104 &  x122 &  x125 &  x128 &  x185 &  x187 &  x188 &  x221 &  x226 &  x227 &  x230 &  x236 &  x239 &  x257 &  x278 &  x281 &  x332 &  x350 &  x359 &  x365 &  x392 &  x398 &  x461 &  x481 &  x484 &  x506 &  x512 &  x519 &  x520 &  x527 &  x539 &  x542 &  x548 &  x554 &  x560 &  x581 &  x587 &  x595 &  x611 &  x634 &  x656 &  x674 &  x680 &  x749 &  x776 &  x806 &  x822 &  x824 &  x830 &  x851 &  x861 &  x884 &  x901 &  x908 &  x938 &  x940 &  x944 &  x959 &  x986 &  x998 &  x1018 &  x1040 &  x1057 &  x1070 &  x1082 &  x1085 &  x1115 &  x1118;
assign c32 =  x8 &  x38 &  x50 &  x68 &  x92 &  x125 &  x134 &  x179 &  x188 &  x236 &  x368 &  x389 &  x431 &  x434 &  x560 &  x611 &  x614 &  x670 &  x725 &  x764 &  x805 &  x827 &  x844 &  x968 &  x977 &  x983 &  x1025 &  x1085 &  x1124 &  x1130 & ~x105 & ~x144 & ~x300 & ~x339 & ~x735 & ~x852 & ~x858 & ~x969 & ~x1068 & ~x1098;
assign c34 =  x8 &  x38 &  x47 &  x98 &  x170 &  x233 &  x239 &  x275 &  x278 &  x296 &  x311 &  x341 &  x356 &  x383 &  x404 &  x419 &  x422 &  x428 &  x434 &  x443 &  x530 &  x533 &  x539 &  x545 &  x554 &  x560 &  x566 &  x575 &  x602 &  x623 &  x632 &  x647 &  x653 &  x686 &  x719 &  x755 &  x758 &  x764 &  x803 &  x806 &  x818 &  x827 &  x848 &  x872 &  x884 &  x914 &  x923 &  x929 &  x938 &  x941 &  x950 &  x962 &  x974 &  x977 &  x983 &  x1031 &  x1046 &  x1052 &  x1064 &  x1067 &  x1079 &  x1112 & ~x30 & ~x837 & ~x870 & ~x909 & ~x921 & ~x993 & ~x1026 & ~x1029 & ~x1032 & ~x1065 & ~x1074 & ~x1089 & ~x1104 & ~x1122;
assign c36 =  x2 &  x44 &  x62 &  x68 &  x164 &  x200 &  x304 &  x314 &  x338 &  x386 &  x442 &  x448 &  x481 &  x487 &  x494 &  x512 &  x536 &  x560 &  x607 &  x645 &  x701 &  x776 &  x782 &  x901 &  x920 &  x965 &  x983 &  x1018 &  x1019 & ~x576;
assign c38 =  x2 &  x8 &  x14 &  x17 &  x20 &  x47 &  x56 &  x68 &  x71 &  x86 &  x89 &  x92 &  x173 &  x179 &  x185 &  x188 &  x200 &  x208 &  x236 &  x244 &  x275 &  x277 &  x284 &  x293 &  x317 &  x323 &  x341 &  x344 &  x350 &  x353 &  x359 &  x365 &  x368 &  x386 &  x394 &  x407 &  x413 &  x431 &  x433 &  x443 &  x461 &  x472 &  x476 &  x497 &  x503 &  x530 &  x539 &  x545 &  x557 &  x608 &  x611 &  x626 &  x628 &  x638 &  x656 &  x667 &  x692 &  x701 &  x708 &  x734 &  x746 &  x752 &  x755 &  x767 &  x773 &  x776 &  x787 &  x791 &  x803 &  x812 &  x815 &  x818 &  x826 &  x827 &  x844 &  x899 &  x902 &  x904 &  x908 &  x914 &  x917 &  x923 &  x926 &  x929 &  x932 &  x941 &  x944 &  x956 &  x959 &  x962 &  x980 &  x983 &  x992 &  x998 &  x1010 &  x1027 &  x1028 &  x1034 &  x1040 &  x1076 &  x1082 &  x1085 &  x1097 &  x1100 &  x1103 &  x1127 & ~x975;
assign c310 =  x2 &  x5 &  x8 &  x11 &  x17 &  x38 &  x41 &  x47 &  x50 &  x56 &  x68 &  x71 &  x74 &  x95 &  x101 &  x104 &  x158 &  x161 &  x164 &  x197 &  x203 &  x215 &  x224 &  x233 &  x236 &  x245 &  x248 &  x257 &  x263 &  x265 &  x293 &  x296 &  x304 &  x323 &  x326 &  x343 &  x350 &  x356 &  x362 &  x365 &  x368 &  x374 &  x403 &  x407 &  x419 &  x434 &  x442 &  x446 &  x448 &  x454 &  x481 &  x487 &  x494 &  x500 &  x503 &  x521 &  x526 &  x533 &  x548 &  x569 &  x590 &  x605 &  x608 &  x611 &  x623 &  x629 &  x632 &  x638 &  x677 &  x686 &  x728 &  x734 &  x746 &  x752 &  x755 &  x758 &  x764 &  x773 &  x806 &  x821 &  x836 &  x848 &  x851 &  x860 &  x875 &  x898 &  x899 &  x901 &  x908 &  x941 &  x950 &  x962 &  x968 &  x976 &  x977 &  x980 &  x995 &  x1015 &  x1016 &  x1018 &  x1028 &  x1040 &  x1043 &  x1057 &  x1067 &  x1070 &  x1085 &  x1088 &  x1096 &  x1103 &  x1121 &  x1124 & ~x282 & ~x351 & ~x390 & ~x699 & ~x738 & ~x921;
assign c312 =  x8 &  x17 &  x23 &  x47 &  x56 &  x71 &  x86 &  x95 &  x104 &  x110 &  x143 &  x161 &  x188 &  x200 &  x208 &  x212 &  x236 &  x257 &  x275 &  x278 &  x284 &  x323 &  x335 &  x356 &  x365 &  x377 &  x398 &  x404 &  x410 &  x425 &  x431 &  x433 &  x434 &  x449 &  x479 &  x482 &  x494 &  x515 &  x518 &  x521 &  x548 &  x550 &  x551 &  x593 &  x602 &  x628 &  x653 &  x656 &  x695 &  x704 &  x709 &  x725 &  x743 &  x746 &  x747 &  x748 &  x751 &  x767 &  x776 &  x787 &  x790 &  x794 &  x826 &  x827 &  x848 &  x865 &  x866 &  x884 &  x926 &  x950 &  x959 &  x968 &  x980 &  x1010 &  x1061 &  x1082 &  x1085 & ~x0 & ~x39 & ~x840 & ~x918 & ~x957 & ~x1053;
assign c314 =  x5 &  x8 &  x17 &  x26 &  x32 &  x38 &  x41 &  x44 &  x47 &  x56 &  x65 &  x71 &  x77 &  x86 &  x89 &  x92 &  x101 &  x104 &  x110 &  x113 &  x128 &  x137 &  x140 &  x158 &  x164 &  x170 &  x182 &  x185 &  x188 &  x191 &  x197 &  x200 &  x221 &  x224 &  x236 &  x257 &  x275 &  x287 &  x314 &  x317 &  x320 &  x322 &  x341 &  x356 &  x365 &  x368 &  x380 &  x386 &  x392 &  x404 &  x407 &  x410 &  x431 &  x433 &  x434 &  x446 &  x464 &  x467 &  x472 &  x479 &  x494 &  x518 &  x542 &  x545 &  x548 &  x581 &  x590 &  x593 &  x628 &  x632 &  x653 &  x659 &  x683 &  x686 &  x710 &  x749 &  x752 &  x770 &  x776 &  x787 &  x788 &  x803 &  x809 &  x818 &  x826 &  x848 &  x854 &  x875 &  x887 &  x905 &  x908 &  x911 &  x917 &  x941 &  x956 &  x962 &  x968 &  x974 &  x980 &  x983 &  x1001 &  x1025 &  x1028 &  x1031 &  x1037 &  x1043 &  x1058 &  x1061 &  x1067 &  x1070 &  x1081 &  x1082 &  x1085 &  x1094 &  x1115 &  x1121 & ~x498 & ~x537 & ~x561 & ~x576 & ~x600 & ~x615 & ~x639;
assign c316 =  x8 &  x14 &  x23 &  x38 &  x44 &  x56 &  x62 &  x68 &  x83 &  x92 &  x95 &  x98 &  x104 &  x113 &  x140 &  x143 &  x149 &  x155 &  x173 &  x176 &  x185 &  x188 &  x194 &  x215 &  x233 &  x242 &  x257 &  x269 &  x278 &  x284 &  x296 &  x311 &  x314 &  x317 &  x320 &  x332 &  x335 &  x344 &  x350 &  x353 &  x356 &  x365 &  x377 &  x383 &  x395 &  x404 &  x422 &  x434 &  x437 &  x443 &  x473 &  x488 &  x491 &  x499 &  x539 &  x548 &  x566 &  x571 &  x572 &  x578 &  x587 &  x599 &  x611 &  x620 &  x629 &  x632 &  x635 &  x650 &  x656 &  x659 &  x668 &  x674 &  x680 &  x688 &  x692 &  x725 &  x728 &  x733 &  x740 &  x752 &  x755 &  x770 &  x773 &  x776 &  x788 &  x791 &  x800 &  x812 &  x839 &  x842 &  x845 &  x848 &  x863 &  x884 &  x908 &  x911 &  x914 &  x932 &  x944 &  x947 &  x953 &  x980 &  x983 &  x1004 &  x1010 &  x1013 &  x1040 &  x1046 &  x1055 &  x1061 &  x1070 &  x1085 &  x1088 &  x1097 &  x1115 &  x1130 & ~x696 & ~x735 & ~x1032 & ~x1072;
assign c318 =  x71 &  x431 &  x448 &  x481 &  x526 &  x565 &  x685 &  x749 &  x1018 &  x1057 &  x1096 & ~x810 & ~x834 & ~x873 & ~x912 & ~x951 & ~x993;
assign c320 =  x2 &  x5 &  x8 &  x11 &  x23 &  x26 &  x29 &  x38 &  x44 &  x56 &  x68 &  x80 &  x92 &  x101 &  x104 &  x110 &  x119 &  x128 &  x140 &  x155 &  x158 &  x161 &  x164 &  x173 &  x179 &  x188 &  x191 &  x200 &  x209 &  x227 &  x257 &  x269 &  x275 &  x284 &  x296 &  x326 &  x332 &  x344 &  x350 &  x353 &  x356 &  x359 &  x368 &  x380 &  x383 &  x398 &  x404 &  x407 &  x413 &  x431 &  x443 &  x455 &  x458 &  x461 &  x473 &  x479 &  x491 &  x494 &  x500 &  x509 &  x512 &  x524 &  x539 &  x548 &  x551 &  x554 &  x560 &  x569 &  x578 &  x584 &  x590 &  x602 &  x605 &  x608 &  x611 &  x632 &  x638 &  x650 &  x665 &  x686 &  x695 &  x701 &  x710 &  x731 &  x734 &  x746 &  x752 &  x758 &  x761 &  x767 &  x773 &  x776 &  x779 &  x788 &  x791 &  x809 &  x824 &  x827 &  x836 &  x845 &  x854 &  x869 &  x872 &  x881 &  x893 &  x896 &  x899 &  x901 &  x911 &  x923 &  x926 &  x932 &  x935 &  x944 &  x959 &  x965 &  x968 &  x977 &  x979 &  x980 &  x983 &  x986 &  x989 &  x998 &  x1001 &  x1028 &  x1031 &  x1040 &  x1043 &  x1046 &  x1070 &  x1079 &  x1088 &  x1091 &  x1100 &  x1103 & ~x39 & ~x618 & ~x657 & ~x696 & ~x697 & ~x735 & ~x804 & ~x870 & ~x909 & ~x969 & ~x1008;
assign c322 =  x35 &  x67 &  x68 &  x86 &  x92 &  x100 &  x140 &  x188 &  x217 &  x256 &  x263 &  x269 &  x287 &  x298 &  x323 &  x335 &  x368 &  x383 &  x386 &  x431 &  x484 &  x494 &  x557 &  x611 &  x656 &  x668 &  x704 &  x746 &  x774 &  x776 &  x803 &  x806 &  x848 &  x854 &  x875 &  x884 &  x898 &  x899 &  x908 &  x917 &  x976 &  x983 &  x985 &  x986 &  x995 &  x1052 &  x1082 &  x1085 &  x1097 &  x1103 &  x1130;
assign c324 =  x8 &  x26 &  x35 &  x56 &  x62 &  x71 &  x92 &  x101 &  x104 &  x107 &  x119 &  x128 &  x158 &  x185 &  x194 &  x215 &  x227 &  x236 &  x257 &  x305 &  x322 &  x329 &  x344 &  x368 &  x394 &  x395 &  x425 &  x431 &  x433 &  x446 &  x449 &  x472 &  x508 &  x509 &  x515 &  x536 &  x542 &  x545 &  x548 &  x550 &  x581 &  x596 &  x628 &  x644 &  x653 &  x656 &  x667 &  x686 &  x698 &  x701 &  x725 &  x745 &  x746 &  x752 &  x761 &  x787 &  x797 &  x803 &  x806 &  x824 &  x826 &  x830 &  x854 &  x884 &  x923 &  x929 &  x965 &  x992 &  x1031 &  x1055 &  x1061 &  x1073 &  x1082 &  x1085 &  x1115 & ~x417 & ~x492 & ~x765 & ~x804;
assign c326 =  x2 &  x8 &  x14 &  x17 &  x56 &  x68 &  x80 &  x86 &  x92 &  x101 &  x158 &  x161 &  x164 &  x194 &  x205 &  x206 &  x236 &  x238 &  x257 &  x275 &  x277 &  x281 &  x293 &  x323 &  x326 &  x338 &  x344 &  x353 &  x356 &  x368 &  x394 &  x404 &  x431 &  x433 &  x434 &  x440 &  x446 &  x472 &  x473 &  x479 &  x485 &  x494 &  x511 &  x533 &  x545 &  x548 &  x554 &  x638 &  x650 &  x656 &  x677 &  x680 &  x701 &  x725 &  x731 &  x746 &  x752 &  x755 &  x758 &  x761 &  x803 &  x806 &  x818 &  x848 &  x854 &  x872 &  x884 &  x935 &  x974 &  x977 &  x983 &  x1010 &  x1019 &  x1028 &  x1061 &  x1082 &  x1085 & ~x522 & ~x537 & ~x561 & ~x576 & ~x600 & ~x601 & ~x615 & ~x639;
assign c328 =  x86 &  x185 &  x188 &  x197 &  x257 &  x269 &  x403 &  x431 &  x439 &  x441 &  x446 &  x481 &  x521 &  x560 &  x590 &  x638 &  x755 &  x806 &  x812 &  x830 &  x848 &  x854 &  x862 &  x884 &  x903 &  x904 &  x932 &  x946 &  x962 &  x985 &  x1019 &  x1028 &  x1079 &  x1082;
assign c330 =  x5 &  x44 &  x67 &  x71 &  x92 &  x100 &  x104 &  x106 &  x143 &  x172 &  x254 &  x257 &  x263 &  x344 &  x412 &  x479 &  x481 &  x524 &  x533 &  x629 &  x653 &  x659 &  x712 &  x713 &  x746 &  x790 &  x806 &  x828 &  x829 &  x868 &  x905 &  x907 &  x983 &  x1013 &  x1048 &  x1081;
assign c332 =  x26 &  x35 &  x38 &  x56 &  x59 &  x65 &  x86 &  x104 &  x122 &  x164 &  x215 &  x269 &  x278 &  x314 &  x323 &  x326 &  x337 &  x341 &  x347 &  x368 &  x374 &  x419 &  x431 &  x451 &  x452 &  x481 &  x490 &  x497 &  x503 &  x551 &  x556 &  x578 &  x595 &  x602 &  x620 &  x623 &  x626 &  x629 &  x634 &  x653 &  x665 &  x710 &  x712 &  x770 &  x790 &  x791 &  x800 &  x827 &  x829 &  x857 &  x872 &  x884 &  x899 &  x907 &  x923 &  x941 &  x980 &  x986 &  x989 &  x992 &  x998 &  x1028 &  x1088 &  x1106 &  x1109 & ~x6 & ~x45 & ~x84 & ~x123 & ~x393;
assign c334 =  x8 &  x17 &  x50 &  x56 &  x68 &  x71 &  x80 &  x92 &  x101 &  x104 &  x137 &  x149 &  x188 &  x200 &  x257 &  x263 &  x272 &  x275 &  x290 &  x317 &  x325 &  x368 &  x374 &  x392 &  x395 &  x403 &  x419 &  x428 &  x431 &  x434 &  x461 &  x467 &  x479 &  x536 &  x545 &  x551 &  x554 &  x584 &  x638 &  x644 &  x656 &  x662 &  x713 &  x746 &  x752 &  x770 &  x773 &  x803 &  x848 &  x866 &  x878 &  x884 &  x899 &  x901 &  x908 &  x923 &  x944 &  x968 &  x974 &  x979 &  x983 &  x992 &  x1016 &  x1018 &  x1043 &  x1057 &  x1076 &  x1082 &  x1088 &  x1096 & ~x39 & ~x42 & ~x78 & ~x156 & ~x165 & ~x351 & ~x417 & ~x429 & ~x456 & ~x468 & ~x612 & ~x651;
assign c336 =  x394 &  x552 &  x611 &  x613 &  x631 &  x727 &  x752 &  x772 &  x803 &  x811 &  x908 &  x1027 & ~x462;
assign c338 =  x17 &  x68 &  x104 &  x149 &  x179 &  x191 &  x209 &  x236 &  x275 &  x299 &  x302 &  x317 &  x380 &  x392 &  x422 &  x434 &  x485 &  x494 &  x512 &  x521 &  x548 &  x584 &  x590 &  x713 &  x821 &  x830 &  x890 &  x953 &  x965 &  x974 &  x983 &  x1016 &  x1028 & ~x10 & ~x21 & ~x27 & ~x39 & ~x49 & ~x78 & ~x156 & ~x183 & ~x189 & ~x195 & ~x228 & ~x417 & ~x930 & ~x1074 & ~x1086;
assign c340 =  x25 &  x64 &  x74 &  x89 &  x155 &  x175 &  x179 &  x193 &  x200 &  x215 &  x260 &  x284 &  x285 &  x287 &  x298 &  x314 &  x368 &  x374 &  x394 &  x403 &  x416 &  x431 &  x433 &  x473 &  x478 &  x479 &  x488 &  x517 &  x548 &  x725 &  x752 &  x788 &  x830 &  x848 &  x860 &  x904 &  x932 &  x941 &  x943 &  x983 &  x986 &  x992 &  x1019 &  x1127;
assign c342 =  x13 &  x14 &  x44 &  x53 &  x92 &  x104 &  x236 &  x248 &  x257 &  x260 &  x263 &  x277 &  x284 &  x296 &  x305 &  x314 &  x356 &  x374 &  x377 &  x422 &  x433 &  x434 &  x437 &  x461 &  x479 &  x533 &  x563 &  x566 &  x584 &  x617 &  x626 &  x635 &  x641 &  x647 &  x662 &  x668 &  x716 &  x719 &  x737 &  x746 &  x755 &  x773 &  x797 &  x803 &  x806 &  x824 &  x842 &  x844 &  x884 &  x896 &  x917 &  x920 &  x926 &  x947 &  x974 &  x977 &  x989 &  x998 &  x1010 &  x1031 &  x1094 &  x1097 & ~x0 & ~x27 & ~x859 & ~x898 & ~x930 & ~x937 & ~x963 & ~x1053 & ~x1086;
assign c344 =  x17 &  x23 &  x62 &  x92 &  x125 &  x131 &  x136 &  x194 &  x215 &  x224 &  x233 &  x239 &  x242 &  x257 &  x272 &  x285 &  x302 &  x305 &  x314 &  x316 &  x323 &  x335 &  x355 &  x368 &  x394 &  x403 &  x433 &  x479 &  x482 &  x494 &  x533 &  x545 &  x548 &  x587 &  x628 &  x638 &  x656 &  x659 &  x686 &  x749 &  x758 &  x805 &  x818 &  x844 &  x845 &  x866 &  x878 &  x883 &  x887 &  x938 &  x962 &  x983 &  x1046 &  x1058 &  x1079 &  x1082 &  x1106 &  x1124 & ~x150;
assign c346 =  x11 &  x29 &  x47 &  x50 &  x56 &  x59 &  x68 &  x71 &  x86 &  x89 &  x98 &  x101 &  x122 &  x134 &  x182 &  x188 &  x194 &  x200 &  x203 &  x206 &  x209 &  x215 &  x224 &  x233 &  x257 &  x260 &  x269 &  x275 &  x302 &  x322 &  x323 &  x329 &  x356 &  x360 &  x361 &  x368 &  x374 &  x399 &  x400 &  x404 &  x413 &  x419 &  x422 &  x425 &  x438 &  x439 &  x455 &  x458 &  x478 &  x503 &  x512 &  x517 &  x524 &  x530 &  x533 &  x548 &  x556 &  x566 &  x569 &  x595 &  x605 &  x611 &  x629 &  x659 &  x665 &  x668 &  x673 &  x686 &  x701 &  x704 &  x752 &  x755 &  x764 &  x767 &  x791 &  x803 &  x818 &  x821 &  x827 &  x842 &  x848 &  x851 &  x869 &  x884 &  x902 &  x911 &  x920 &  x923 &  x929 &  x938 &  x968 &  x977 &  x986 &  x1004 &  x1010 &  x1028 &  x1040 &  x1043 &  x1046 &  x1052 &  x1070 &  x1091 &  x1097 &  x1106 &  x1130 & ~x162 & ~x240 & ~x1056 & ~x1095;
assign c348 =  x5 &  x8 &  x17 &  x38 &  x44 &  x56 &  x62 &  x68 &  x71 &  x74 &  x77 &  x89 &  x92 &  x95 &  x104 &  x137 &  x140 &  x158 &  x170 &  x176 &  x188 &  x194 &  x203 &  x215 &  x221 &  x257 &  x269 &  x275 &  x281 &  x347 &  x365 &  x368 &  x383 &  x407 &  x419 &  x434 &  x440 &  x443 &  x473 &  x494 &  x503 &  x506 &  x520 &  x533 &  x536 &  x542 &  x545 &  x548 &  x554 &  x556 &  x566 &  x595 &  x602 &  x605 &  x629 &  x632 &  x638 &  x656 &  x665 &  x689 &  x702 &  x752 &  x767 &  x773 &  x776 &  x794 &  x797 &  x806 &  x812 &  x815 &  x820 &  x827 &  x830 &  x839 &  x848 &  x860 &  x862 &  x884 &  x893 &  x899 &  x901 &  x908 &  x911 &  x923 &  x929 &  x962 &  x968 &  x974 &  x976 &  x979 &  x980 &  x992 &  x1015 &  x1018 &  x1028 &  x1057 &  x1058 &  x1070 &  x1082 &  x1088 &  x1091 &  x1096 &  x1100 &  x1103 & ~x669 & ~x687 & ~x708 & ~x726 & ~x747 & ~x834 & ~x873 & ~x912;
assign c350 =  x11 &  x104 &  x152 &  x170 &  x173 &  x236 &  x296 &  x386 &  x403 &  x434 &  x439 &  x441 &  x481 &  x527 &  x533 &  x539 &  x548 &  x602 &  x695 &  x698 &  x773 &  x803 &  x815 &  x878 &  x884 &  x901 &  x905 &  x917 &  x962 &  x1018 &  x1022 &  x1055 &  x1070 & ~x39 & ~x78 & ~x313 & ~x429 & ~x507 & ~x1053 & ~x1092;
assign c352 =  x2 &  x8 &  x17 &  x44 &  x50 &  x56 &  x59 &  x62 &  x89 &  x92 &  x95 &  x104 &  x107 &  x128 &  x137 &  x140 &  x188 &  x200 &  x209 &  x224 &  x227 &  x236 &  x251 &  x257 &  x269 &  x275 &  x278 &  x281 &  x284 &  x296 &  x299 &  x310 &  x323 &  x338 &  x341 &  x350 &  x362 &  x368 &  x383 &  x413 &  x416 &  x422 &  x434 &  x443 &  x448 &  x473 &  x481 &  x487 &  x490 &  x494 &  x500 &  x503 &  x518 &  x521 &  x529 &  x530 &  x533 &  x545 &  x557 &  x596 &  x598 &  x605 &  x611 &  x623 &  x629 &  x632 &  x637 &  x638 &  x656 &  x659 &  x722 &  x725 &  x740 &  x746 &  x752 &  x758 &  x773 &  x782 &  x803 &  x812 &  x815 &  x818 &  x823 &  x830 &  x836 &  x845 &  x848 &  x863 &  x866 &  x875 &  x884 &  x893 &  x898 &  x899 &  x902 &  x908 &  x929 &  x932 &  x937 &  x962 &  x968 &  x974 &  x979 &  x980 &  x983 &  x995 &  x1007 &  x1016 &  x1018 &  x1019 &  x1028 &  x1043 &  x1055 &  x1057 &  x1063 &  x1076 &  x1079 &  x1082 &  x1091 &  x1096 &  x1097 &  x1103 & ~x351 & ~x390 & ~x873 & ~x912 & ~x951;
assign c354 =  x5 &  x8 &  x14 &  x47 &  x50 &  x56 &  x59 &  x62 &  x71 &  x86 &  x89 &  x104 &  x140 &  x164 &  x185 &  x188 &  x194 &  x200 &  x203 &  x215 &  x224 &  x233 &  x236 &  x242 &  x275 &  x284 &  x296 &  x298 &  x332 &  x335 &  x337 &  x344 &  x356 &  x365 &  x368 &  x374 &  x400 &  x403 &  x406 &  x428 &  x431 &  x438 &  x439 &  x440 &  x442 &  x473 &  x478 &  x482 &  x494 &  x500 &  x517 &  x518 &  x521 &  x533 &  x545 &  x548 &  x563 &  x578 &  x620 &  x625 &  x632 &  x659 &  x680 &  x683 &  x703 &  x706 &  x722 &  x746 &  x752 &  x755 &  x785 &  x788 &  x803 &  x839 &  x848 &  x854 &  x875 &  x884 &  x901 &  x902 &  x904 &  x917 &  x929 &  x943 &  x962 &  x968 &  x983 &  x989 &  x992 &  x995 &  x1010 &  x1019 &  x1022 &  x1097 &  x1103 &  x1112 &  x1130 & ~x351;
assign c356 =  x61 &  x86 &  x88 &  x92 &  x217 &  x236 &  x322 &  x368 &  x451 &  x487 &  x488 &  x490 &  x545 &  x595 &  x602 &  x683 &  x772 &  x790 &  x803 &  x811 &  x868 &  x1013 &  x1082;
assign c358 =  x56 &  x62 &  x179 &  x215 &  x278 &  x394 &  x398 &  x437 &  x632 &  x638 &  x737 &  x788 &  x827 &  x902 &  x932 &  x998 &  x1049 &  x1088 &  x1094 &  x1109 &  x1127 & ~x30 & ~x69 & ~x639 & ~x792 & ~x870 & ~x915 & ~x945 & ~x984 & ~x1065 & ~x1089 & ~x1104;
assign c360 =  x5 &  x8 &  x86 &  x89 &  x92 &  x155 &  x164 &  x281 &  x320 &  x350 &  x362 &  x446 &  x460 &  x484 &  x536 &  x598 &  x637 &  x643 &  x656 &  x668 &  x682 &  x752 &  x776 &  x901 &  x947 &  x978 &  x983 &  x1007 &  x1015 &  x1017 &  x1018 &  x1056 &  x1057 &  x1093 &  x1095 &  x1096 & ~x399 & ~x468 & ~x546 & ~x1029 & ~x1068;
assign c362 =  x50 &  x56 &  x173 &  x188 &  x236 &  x254 &  x287 &  x326 &  x335 &  x386 &  x404 &  x422 &  x449 &  x464 &  x476 &  x494 &  x497 &  x506 &  x515 &  x551 &  x632 &  x634 &  x698 &  x776 &  x848 &  x851 &  x857 &  x939 &  x965 &  x1018 &  x1037 &  x1040 &  x1057 &  x1059 &  x1061 &  x1094 &  x1096 &  x1098 &  x1109 &  x1124 & ~x39 & ~x78 & ~x195 & ~x507;
assign c364 =  x40 &  x92 &  x157 &  x188 &  x224 &  x236 &  x392 &  x479 &  x485 &  x713 &  x731 &  x983 & ~x69 & ~x96 & ~x141 & ~x153 & ~x180 & ~x192 & ~x264 & ~x309 & ~x387 & ~x870 & ~x909 & ~x987 & ~x993 & ~x1032 & ~x1050 & ~x1065 & ~x1089 & ~x1116 & ~x1122;
assign c366 =  x5 &  x8 &  x11 &  x20 &  x38 &  x44 &  x56 &  x59 &  x71 &  x86 &  x98 &  x101 &  x104 &  x110 &  x113 &  x119 &  x128 &  x137 &  x143 &  x164 &  x187 &  x188 &  x194 &  x197 &  x200 &  x218 &  x221 &  x224 &  x226 &  x236 &  x257 &  x263 &  x265 &  x272 &  x275 &  x281 &  x290 &  x296 &  x299 &  x314 &  x326 &  x344 &  x350 &  x353 &  x356 &  x359 &  x362 &  x368 &  x380 &  x383 &  x389 &  x398 &  x403 &  x404 &  x413 &  x431 &  x434 &  x442 &  x470 &  x476 &  x479 &  x491 &  x494 &  x503 &  x509 &  x512 &  x515 &  x518 &  x521 &  x533 &  x536 &  x545 &  x547 &  x548 &  x554 &  x560 &  x586 &  x590 &  x623 &  x625 &  x632 &  x638 &  x656 &  x662 &  x677 &  x680 &  x703 &  x713 &  x731 &  x737 &  x743 &  x746 &  x752 &  x755 &  x770 &  x773 &  x779 &  x782 &  x803 &  x812 &  x824 &  x827 &  x830 &  x836 &  x845 &  x848 &  x854 &  x860 &  x862 &  x869 &  x893 &  x901 &  x911 &  x917 &  x929 &  x932 &  x941 &  x959 &  x962 &  x968 &  x974 &  x980 &  x983 &  x995 &  x998 &  x1010 &  x1040 &  x1070 &  x1082 &  x1085 &  x1097 &  x1130 & ~x351 & ~x552 & ~x553 & ~x591 & ~x592 & ~x792 & ~x834;
assign c368 =  x5 &  x8 &  x38 &  x86 &  x92 &  x101 &  x104 &  x116 &  x137 &  x158 &  x164 &  x168 &  x182 &  x205 &  x208 &  x257 &  x263 &  x272 &  x277 &  x281 &  x284 &  x287 &  x296 &  x320 &  x335 &  x356 &  x383 &  x422 &  x430 &  x431 &  x433 &  x461 &  x479 &  x511 &  x533 &  x545 &  x560 &  x590 &  x608 &  x638 &  x656 &  x659 &  x689 &  x701 &  x710 &  x746 &  x755 &  x772 &  x773 &  x803 &  x811 &  x818 &  x845 &  x848 &  x854 &  x872 &  x875 &  x884 &  x905 &  x917 &  x923 &  x944 &  x962 &  x968 &  x983 &  x1028 &  x1082 &  x1100 &  x1109 &  x1124 & ~x522 & ~x561 & ~x897;
assign c370 =  x2 &  x5 &  x8 &  x14 &  x17 &  x20 &  x38 &  x47 &  x59 &  x92 &  x173 &  x188 &  x205 &  x206 &  x238 &  x257 &  x260 &  x276 &  x277 &  x287 &  x332 &  x355 &  x368 &  x377 &  x404 &  x407 &  x433 &  x449 &  x472 &  x494 &  x536 &  x550 &  x569 &  x644 &  x677 &  x728 &  x752 &  x773 &  x794 &  x812 &  x833 &  x842 &  x935 &  x941 &  x983 &  x1067 &  x1076 &  x1082 &  x1124 & ~x105 & ~x537 & ~x813 & ~x969 & ~x1047 & ~x1086;
assign c372 =  x8 &  x47 &  x56 &  x68 &  x71 &  x101 &  x104 &  x125 &  x158 &  x164 &  x176 &  x188 &  x236 &  x263 &  x275 &  x277 &  x326 &  x329 &  x356 &  x365 &  x394 &  x395 &  x422 &  x431 &  x433 &  x434 &  x470 &  x472 &  x479 &  x482 &  x494 &  x539 &  x548 &  x554 &  x563 &  x569 &  x611 &  x623 &  x626 &  x635 &  x656 &  x668 &  x670 &  x671 &  x725 &  x740 &  x755 &  x791 &  x806 &  x848 &  x854 &  x896 &  x962 &  x968 &  x995 &  x1001 &  x1010 &  x1016 &  x1079 &  x1094 &  x1106 & ~x0 & ~x105 & ~x144 & ~x222 & ~x300 & ~x339 & ~x600 & ~x639 & ~x885 & ~x891 & ~x930 & ~x963 & ~x969 & ~x1002 & ~x1029 & ~x1068 & ~x1092 & ~x1107;
assign c374 =  x5 &  x23 &  x41 &  x56 &  x92 &  x95 &  x98 &  x101 &  x122 &  x131 &  x134 &  x152 &  x164 &  x170 &  x188 &  x203 &  x205 &  x212 &  x221 &  x233 &  x244 &  x245 &  x250 &  x251 &  x281 &  x320 &  x321 &  x322 &  x361 &  x365 &  x389 &  x401 &  x433 &  x437 &  x479 &  x482 &  x508 &  x545 &  x595 &  x628 &  x634 &  x644 &  x671 &  x673 &  x686 &  x704 &  x707 &  x712 &  x728 &  x749 &  x755 &  x782 &  x818 &  x821 &  x854 &  x875 &  x911 &  x932 &  x965 &  x977 &  x992 &  x1013 &  x1019 &  x1028 &  x1058 &  x1076 &  x1112;
assign c376 =  x8 &  x56 &  x71 &  x92 &  x116 &  x131 &  x194 &  x251 &  x431 &  x533 &  x545 &  x602 &  x677 &  x708 &  x826 &  x848 &  x863 &  x881 &  x884 &  x1061 & ~x39 & ~x300 & ~x339 & ~x522 & ~x561 & ~x600 & ~x840 & ~x936 & ~x1056 & ~x1095;
assign c378 =  x20 &  x44 &  x71 &  x86 &  x89 &  x104 &  x137 &  x140 &  x143 &  x194 &  x200 &  x215 &  x230 &  x233 &  x263 &  x275 &  x281 &  x284 &  x314 &  x323 &  x338 &  x343 &  x377 &  x380 &  x395 &  x410 &  x431 &  x442 &  x473 &  x488 &  x494 &  x500 &  x509 &  x517 &  x533 &  x545 &  x548 &  x551 &  x554 &  x555 &  x556 &  x557 &  x560 &  x566 &  x595 &  x605 &  x617 &  x629 &  x650 &  x677 &  x695 &  x698 &  x702 &  x725 &  x737 &  x740 &  x752 &  x761 &  x803 &  x806 &  x815 &  x818 &  x824 &  x848 &  x887 &  x890 &  x896 &  x899 &  x901 &  x908 &  x917 &  x923 &  x941 &  x947 &  x971 &  x974 &  x983 &  x992 &  x998 &  x1016 &  x1028 &  x1034 &  x1064 &  x1079 &  x1085 &  x1088 &  x1097 &  x1121 & ~x670;
assign c380 =  x13 &  x16 &  x20 &  x44 &  x49 &  x92 &  x101 &  x131 &  x140 &  x155 &  x164 &  x194 &  x221 &  x224 &  x269 &  x281 &  x365 &  x398 &  x413 &  x434 &  x515 &  x566 &  x595 &  x608 &  x613 &  x638 &  x661 &  x677 &  x710 &  x725 &  x778 &  x803 &  x811 &  x854 &  x902 &  x917 &  x980 &  x989 &  x992 &  x1031 &  x1040 &  x1043 &  x1088 &  x1091 &  x1115 &  x1123;
assign c382 =  x5 &  x17 &  x32 &  x35 &  x38 &  x50 &  x56 &  x62 &  x71 &  x74 &  x83 &  x86 &  x92 &  x101 &  x104 &  x119 &  x137 &  x140 &  x146 &  x149 &  x152 &  x155 &  x164 &  x167 &  x179 &  x182 &  x185 &  x188 &  x191 &  x221 &  x227 &  x233 &  x236 &  x248 &  x257 &  x269 &  x272 &  x275 &  x284 &  x290 &  x293 &  x296 &  x298 &  x302 &  x314 &  x317 &  x323 &  x332 &  x338 &  x353 &  x356 &  x359 &  x368 &  x374 &  x380 &  x383 &  x394 &  x398 &  x403 &  x404 &  x410 &  x425 &  x431 &  x433 &  x434 &  x437 &  x443 &  x470 &  x472 &  x473 &  x476 &  x479 &  x482 &  x485 &  x494 &  x503 &  x508 &  x511 &  x512 &  x521 &  x527 &  x539 &  x545 &  x548 &  x551 &  x557 &  x566 &  x572 &  x584 &  x599 &  x602 &  x605 &  x608 &  x611 &  x623 &  x628 &  x629 &  x632 &  x656 &  x659 &  x667 &  x680 &  x695 &  x701 &  x707 &  x710 &  x713 &  x719 &  x725 &  x743 &  x745 &  x746 &  x749 &  x752 &  x755 &  x764 &  x776 &  x779 &  x797 &  x803 &  x806 &  x809 &  x818 &  x824 &  x826 &  x830 &  x836 &  x845 &  x848 &  x854 &  x862 &  x866 &  x875 &  x884 &  x893 &  x896 &  x901 &  x904 &  x917 &  x941 &  x943 &  x944 &  x956 &  x968 &  x974 &  x980 &  x983 &  x992 &  x1007 &  x1010 &  x1013 &  x1016 &  x1022 &  x1028 &  x1031 &  x1034 &  x1055 &  x1061 &  x1070 &  x1076 &  x1082 &  x1091 &  x1094 &  x1097 &  x1103 &  x1112 &  x1121 &  x1124 &  x1130 & ~x117 & ~x156 & ~x195 & ~x273 & ~x639 & ~x678 & ~x717 & ~x756;
assign c384 =  x8 &  x14 &  x17 &  x53 &  x56 &  x71 &  x101 &  x104 &  x119 &  x137 &  x179 &  x188 &  x194 &  x215 &  x242 &  x356 &  x365 &  x368 &  x404 &  x433 &  x434 &  x482 &  x641 &  x650 &  x656 &  x662 &  x710 &  x746 &  x754 &  x790 &  x806 &  x818 &  x848 &  x854 &  x895 &  x911 &  x956 &  x962 &  x983 &  x995 &  x998 &  x1007 &  x1052 &  x1079 &  x1097 & ~x492 & ~x522 & ~x561 & ~x903 & ~x1098;
assign c386 =  x17 &  x159 &  x315 &  x393 &  x398 &  x432 &  x433 &  x472 &  x473 &  x545 &  x787 &  x805 &  x854 &  x983 &  x1019 &  x1091 & ~x717 & ~x781;
assign c388 =  x47 &  x50 &  x134 &  x155 &  x236 &  x263 &  x277 &  x302 &  x305 &  x316 &  x317 &  x323 &  x368 &  x394 &  x422 &  x428 &  x433 &  x506 &  x589 &  x596 &  x628 &  x632 &  x683 &  x686 &  x692 &  x695 &  x725 &  x1040 & ~x339 & ~x340 & ~x378 & ~x379 & ~x417 & ~x456 & ~x639 & ~x897 & ~x930 & ~x969 & ~x984 & ~x1068 & ~x1107;
assign c390 =  x17 &  x44 &  x92 &  x176 &  x188 &  x215 &  x266 &  x326 &  x361 &  x368 &  x439 &  x478 &  x494 &  x512 &  x517 &  x569 &  x574 &  x598 &  x668 &  x722 &  x725 &  x743 &  x772 &  x787 &  x803 &  x805 &  x826 &  x845 &  x875 &  x917 &  x1004 &  x1091 & ~x1017 & ~x1056 & ~x1095;
assign c392 =  x86 &  x236 &  x263 &  x275 &  x394 &  x404 &  x433 &  x479 &  x514 &  x533 &  x545 &  x548 &  x591 &  x605 &  x670 &  x688 &  x739 &  x746 &  x773 &  x779 &  x797 &  x803 &  x805 &  x811 &  x826 &  x830 &  x836 &  x850 &  x854 &  x865 &  x884 &  x904 &  x910 &  x917 &  x983 &  x1019 &  x1028 &  x1061 &  x1082 & ~x703 & ~x741 & ~x742 & ~x781 & ~x1095;
assign c394 =  x8 &  x11 &  x17 &  x20 &  x38 &  x41 &  x44 &  x53 &  x56 &  x71 &  x86 &  x95 &  x101 &  x104 &  x137 &  x155 &  x164 &  x206 &  x233 &  x236 &  x257 &  x266 &  x278 &  x326 &  x353 &  x368 &  x392 &  x398 &  x404 &  x431 &  x448 &  x455 &  x479 &  x482 &  x487 &  x494 &  x503 &  x521 &  x524 &  x533 &  x542 &  x545 &  x548 &  x566 &  x590 &  x593 &  x605 &  x629 &  x647 &  x656 &  x734 &  x737 &  x746 &  x752 &  x776 &  x797 &  x800 &  x815 &  x830 &  x848 &  x859 &  x860 &  x875 &  x884 &  x899 &  x900 &  x917 &  x939 &  x953 &  x962 &  x965 &  x974 &  x979 &  x983 &  x998 &  x1001 &  x1018 &  x1028 &  x1043 &  x1046 &  x1057 &  x1070 &  x1088 &  x1103 & ~x807 & ~x951 & ~x990 & ~x1008 & ~x1029 & ~x1032 & ~x1068 & ~x1071;
assign c396 =  x11 &  x53 &  x62 &  x104 &  x106 &  x215 &  x221 &  x281 &  x290 &  x320 &  x347 &  x362 &  x404 &  x407 &  x410 &  x437 &  x461 &  x497 &  x614 &  x638 &  x665 &  x680 &  x701 &  x713 &  x752 &  x761 &  x848 &  x923 &  x962 &  x974 &  x986 &  x989 &  x1025 &  x1061 & ~x69 & ~x225 & ~x603 & ~x792 & ~x837 & ~x948 & ~x954 & ~x987 & ~x993 & ~x1026 & ~x1089 & ~x1104 & ~x1116;
assign c398 =  x13 &  x40 &  x118 &  x195 &  x314 &  x315 &  x335 &  x433 &  x652 &  x812 &  x844 &  x848 &  x938 & ~x507;
assign c3100 =  x8 &  x17 &  x56 &  x86 &  x92 &  x104 &  x110 &  x146 &  x188 &  x227 &  x344 &  x356 &  x365 &  x368 &  x377 &  x383 &  x455 &  x467 &  x479 &  x481 &  x484 &  x493 &  x494 &  x503 &  x519 &  x536 &  x545 &  x556 &  x575 &  x595 &  x605 &  x611 &  x632 &  x634 &  x638 &  x653 &  x656 &  x686 &  x746 &  x752 &  x755 &  x776 &  x788 &  x803 &  x827 &  x848 &  x851 &  x854 &  x884 &  x890 &  x904 &  x907 &  x911 &  x917 &  x935 &  x941 &  x943 &  x944 &  x946 &  x959 &  x974 &  x983 &  x985 &  x1001 &  x1007 &  x1024 &  x1028 &  x1091 &  x1100 &  x1121 & ~x429;
assign c3102 =  x41 &  x56 &  x176 &  x236 &  x269 &  x302 &  x467 &  x478 &  x506 &  x515 &  x517 &  x548 &  x556 &  x604 &  x643 &  x665 &  x668 &  x682 &  x692 &  x698 &  x721 &  x737 &  x752 &  x803 &  x830 &  x923 &  x980 &  x1100 &  x1109 & ~x84 & ~x123 & ~x162 & ~x699 & ~x825 & ~x1098;
assign c3104 =  x5 &  x17 &  x38 &  x62 &  x65 &  x71 &  x89 &  x104 &  x119 &  x164 &  x188 &  x191 &  x233 &  x238 &  x251 &  x257 &  x274 &  x277 &  x316 &  x350 &  x374 &  x383 &  x394 &  x398 &  x419 &  x443 &  x476 &  x479 &  x482 &  x515 &  x527 &  x533 &  x542 &  x545 &  x548 &  x554 &  x557 &  x563 &  x578 &  x584 &  x593 &  x631 &  x635 &  x653 &  x695 &  x701 &  x707 &  x709 &  x713 &  x746 &  x755 &  x767 &  x773 &  x776 &  x782 &  x788 &  x803 &  x805 &  x812 &  x836 &  x854 &  x860 &  x875 &  x890 &  x893 &  x932 &  x968 &  x971 &  x973 &  x974 &  x986 &  x1007 &  x1028 &  x1079 &  x1082 &  x1097 &  x1103 &  x1127 &  x1130 & ~x27 & ~x366 & ~x367 & ~x405 & ~x406 & ~x585 & ~x625 & ~x664 & ~x705 & ~x742 & ~x897 & ~x936 & ~x1014 & ~x1053 & ~x1092;
assign c3106 =  x2 &  x8 &  x17 &  x23 &  x38 &  x41 &  x53 &  x56 &  x59 &  x62 &  x68 &  x71 &  x86 &  x92 &  x104 &  x110 &  x128 &  x155 &  x161 &  x164 &  x179 &  x185 &  x188 &  x194 &  x215 &  x221 &  x230 &  x233 &  x236 &  x251 &  x254 &  x260 &  x263 &  x266 &  x272 &  x278 &  x281 &  x290 &  x311 &  x326 &  x332 &  x347 &  x368 &  x374 &  x425 &  x434 &  x455 &  x470 &  x473 &  x478 &  x479 &  x482 &  x488 &  x503 &  x521 &  x524 &  x530 &  x536 &  x545 &  x548 &  x557 &  x560 &  x569 &  x584 &  x590 &  x602 &  x605 &  x632 &  x650 &  x656 &  x663 &  x674 &  x677 &  x680 &  x689 &  x692 &  x702 &  x703 &  x741 &  x746 &  x749 &  x752 &  x755 &  x761 &  x773 &  x785 &  x788 &  x803 &  x818 &  x833 &  x854 &  x863 &  x872 &  x875 &  x887 &  x893 &  x898 &  x899 &  x901 &  x908 &  x926 &  x940 &  x947 &  x959 &  x962 &  x968 &  x971 &  x974 &  x983 &  x989 &  x992 &  x1007 &  x1010 &  x1019 &  x1022 &  x1031 &  x1040 &  x1055 &  x1070 &  x1073 &  x1076 &  x1082 &  x1091 &  x1097 &  x1103 &  x1109 &  x1115 &  x1118 &  x1124 &  x1130 & ~x669 & ~x708 & ~x726 & ~x816 & ~x834 & ~x1104;
assign c3108 =  x17 &  x67 &  x71 &  x73 &  x80 &  x86 &  x92 &  x101 &  x104 &  x106 &  x110 &  x112 &  x128 &  x145 &  x155 &  x184 &  x206 &  x211 &  x223 &  x224 &  x236 &  x245 &  x248 &  x257 &  x266 &  x281 &  x287 &  x307 &  x332 &  x335 &  x344 &  x356 &  x365 &  x368 &  x403 &  x404 &  x443 &  x448 &  x479 &  x484 &  x494 &  x506 &  x509 &  x524 &  x542 &  x593 &  x614 &  x653 &  x665 &  x683 &  x755 &  x782 &  x785 &  x854 &  x868 &  x902 &  x907 &  x917 &  x946 &  x968 &  x971 &  x985 &  x1001 &  x1018 &  x1079 &  x1112 &  x1127 & ~x669 & ~x1104;
assign c3110 =  x8 &  x17 &  x170 &  x185 &  x209 &  x269 &  x275 &  x407 &  x460 &  x490 &  x529 &  x558 &  x595 &  x597 &  x598 &  x656 &  x677 &  x686 &  x734 &  x746 &  x755 &  x764 &  x803 &  x812 &  x818 &  x848 &  x854 &  x974 &  x985 &  x1018 &  x1019 &  x1057 &  x1067 &  x1130 & ~x429;
assign c3112 =  x8 &  x13 &  x26 &  x35 &  x68 &  x86 &  x89 &  x98 &  x140 &  x188 &  x203 &  x212 &  x227 &  x233 &  x236 &  x275 &  x277 &  x284 &  x313 &  x352 &  x368 &  x371 &  x394 &  x401 &  x425 &  x428 &  x431 &  x433 &  x434 &  x472 &  x488 &  x494 &  x503 &  x533 &  x545 &  x548 &  x563 &  x590 &  x656 &  x683 &  x727 &  x733 &  x739 &  x752 &  x755 &  x770 &  x772 &  x778 &  x787 &  x806 &  x811 &  x812 &  x817 &  x821 &  x824 &  x826 &  x830 &  x838 &  x844 &  x848 &  x850 &  x856 &  x877 &  x887 &  x895 &  x896 &  x910 &  x928 &  x934 &  x968 &  x973 &  x983 &  x994 &  x1028 &  x1034 &  x1055 & ~x522 & ~x561 & ~x585 & ~x600;
assign c3114 =  x2 &  x5 &  x8 &  x35 &  x38 &  x44 &  x47 &  x50 &  x56 &  x71 &  x77 &  x86 &  x89 &  x92 &  x104 &  x107 &  x110 &  x119 &  x128 &  x134 &  x137 &  x155 &  x161 &  x164 &  x176 &  x179 &  x185 &  x188 &  x200 &  x251 &  x257 &  x263 &  x275 &  x278 &  x281 &  x284 &  x296 &  x329 &  x344 &  x356 &  x371 &  x374 &  x404 &  x419 &  x422 &  x431 &  x434 &  x442 &  x473 &  x481 &  x482 &  x494 &  x500 &  x515 &  x519 &  x527 &  x533 &  x539 &  x545 &  x554 &  x557 &  x559 &  x572 &  x581 &  x590 &  x598 &  x605 &  x608 &  x611 &  x629 &  x632 &  x659 &  x667 &  x704 &  x725 &  x752 &  x758 &  x773 &  x776 &  x785 &  x797 &  x803 &  x812 &  x823 &  x830 &  x833 &  x862 &  x893 &  x899 &  x901 &  x907 &  x908 &  x917 &  x946 &  x962 &  x977 &  x992 &  x995 &  x1010 &  x1031 &  x1046 &  x1073 &  x1097 &  x1100 &  x1103 &  x1130 & ~x648 & ~x687 & ~x726 & ~x765;
assign c3116 =  x17 &  x86 &  x113 &  x170 &  x197 &  x233 &  x254 &  x286 &  x288 &  x296 &  x324 &  x355 &  x362 &  x363 &  x398 &  x403 &  x433 &  x442 &  x481 &  x482 &  x494 &  x521 &  x545 &  x551 &  x560 &  x569 &  x599 &  x605 &  x614 &  x650 &  x667 &  x746 &  x773 &  x779 &  x794 &  x818 &  x851 &  x893 &  x917 &  x962 &  x968 &  x974 &  x983 &  x1031 &  x1043 &  x1091 & ~x273;
assign c3118 =  x8 &  x17 &  x20 &  x44 &  x50 &  x56 &  x86 &  x89 &  x92 &  x101 &  x104 &  x137 &  x140 &  x143 &  x155 &  x164 &  x188 &  x191 &  x209 &  x236 &  x257 &  x281 &  x311 &  x323 &  x368 &  x410 &  x413 &  x434 &  x443 &  x448 &  x481 &  x487 &  x494 &  x519 &  x533 &  x545 &  x565 &  x584 &  x605 &  x628 &  x656 &  x667 &  x707 &  x752 &  x755 &  x822 &  x824 &  x854 &  x868 &  x872 &  x875 &  x935 &  x941 &  x974 &  x983 &  x1016 &  x1018 &  x1043 &  x1046 &  x1057 &  x1082 & ~x273;
assign c3120 =  x88 &  x433 &  x778 &  x844 &  x850 &  x856 &  x934 &  x1046 &  x1079 & ~x820 & ~x859 & ~x1095;
assign c3122 =  x2 &  x38 &  x104 &  x188 &  x257 &  x338 &  x368 &  x394 &  x419 &  x503 &  x545 &  x644 &  x826 &  x854 &  x884 &  x926 &  x962 &  x1049 &  x1130 & ~x66 & ~x228 & ~x339 & ~x522 & ~x561 & ~x600 & ~x601 & ~x639 & ~x834 & ~x879 & ~x912;
assign c3124 =  x17 &  x106 &  x184 &  x222 &  x223 &  x236 &  x257 &  x368 &  x539 &  x742 &  x746 &  x806 &  x848 &  x908 &  x917 & ~x699 & ~x993 & ~x1029;
assign c3126 =  x2 &  x17 &  x50 &  x104 &  x149 &  x155 &  x182 &  x188 &  x197 &  x269 &  x311 &  x317 &  x323 &  x331 &  x347 &  x374 &  x392 &  x404 &  x428 &  x467 &  x479 &  x482 &  x494 &  x503 &  x512 &  x533 &  x545 &  x550 &  x575 &  x590 &  x595 &  x596 &  x634 &  x635 &  x665 &  x680 &  x698 &  x713 &  x745 &  x746 &  x752 &  x767 &  x773 &  x776 &  x782 &  x800 &  x818 &  x839 &  x851 &  x854 &  x881 &  x896 &  x899 &  x935 &  x986 &  x1034 &  x1052 &  x1091 &  x1097 &  x1118 & ~x765 & ~x804 & ~x930 & ~x931 & ~x969 & ~x1008;
assign c3128 =  x11 &  x47 &  x101 &  x104 &  x209 &  x227 &  x242 &  x257 &  x356 &  x362 &  x368 &  x448 &  x451 &  x458 &  x464 &  x490 &  x521 &  x548 &  x560 &  x569 &  x595 &  x608 &  x629 &  x632 &  x638 &  x713 &  x725 &  x758 &  x773 &  x779 &  x788 &  x809 &  x815 &  x866 &  x900 &  x937 &  x939 &  x974 &  x978 &  x979 &  x1017 &  x1018 &  x1056 &  x1082 & ~x507 & ~x1107;
assign c3130 =  x11 &  x17 &  x25 &  x38 &  x86 &  x89 &  x92 &  x101 &  x110 &  x113 &  x188 &  x200 &  x224 &  x244 &  x257 &  x277 &  x350 &  x368 &  x389 &  x392 &  x394 &  x398 &  x404 &  x431 &  x433 &  x461 &  x494 &  x500 &  x511 &  x521 &  x533 &  x539 &  x554 &  x560 &  x605 &  x611 &  x614 &  x628 &  x641 &  x671 &  x677 &  x731 &  x746 &  x776 &  x826 &  x866 &  x893 &  x908 &  x947 &  x983 &  x1022 &  x1028 &  x1046 &  x1061 &  x1064 &  x1070 &  x1100 & ~x522 & ~x600 & ~x639 & ~x640 & ~x717;
assign c3132 =  x8 &  x38 &  x50 &  x53 &  x110 &  x125 &  x137 &  x155 &  x158 &  x164 &  x179 &  x188 &  x200 &  x206 &  x221 &  x224 &  x233 &  x236 &  x242 &  x263 &  x278 &  x290 &  x299 &  x338 &  x341 &  x347 &  x356 &  x368 &  x371 &  x416 &  x425 &  x434 &  x455 &  x461 &  x470 &  x494 &  x515 &  x533 &  x539 &  x545 &  x548 &  x554 &  x569 &  x589 &  x628 &  x638 &  x653 &  x656 &  x667 &  x677 &  x710 &  x719 &  x734 &  x745 &  x755 &  x776 &  x782 &  x785 &  x803 &  x821 &  x830 &  x836 &  x842 &  x851 &  x881 &  x901 &  x908 &  x911 &  x932 &  x941 &  x947 &  x962 &  x974 &  x983 &  x989 &  x1001 &  x1061 &  x1082 &  x1103 &  x1109 &  x1115 &  x1121 & ~x27 & ~x66 & ~x78 & ~x144 & ~x189 & ~x195 & ~x228 & ~x234 & ~x417 & ~x834 & ~x1047 & ~x1086 & ~x1104;
assign c3134 =  x17 &  x22 &  x35 &  x44 &  x47 &  x50 &  x56 &  x61 &  x68 &  x71 &  x74 &  x89 &  x92 &  x98 &  x99 &  x100 &  x101 &  x104 &  x107 &  x110 &  x116 &  x122 &  x137 &  x138 &  x139 &  x158 &  x161 &  x178 &  x188 &  x194 &  x200 &  x209 &  x217 &  x218 &  x221 &  x233 &  x236 &  x263 &  x269 &  x275 &  x278 &  x281 &  x290 &  x293 &  x296 &  x308 &  x314 &  x320 &  x350 &  x365 &  x368 &  x374 &  x377 &  x383 &  x395 &  x398 &  x419 &  x431 &  x443 &  x446 &  x461 &  x464 &  x467 &  x473 &  x479 &  x494 &  x497 &  x533 &  x548 &  x569 &  x572 &  x593 &  x596 &  x602 &  x605 &  x608 &  x611 &  x632 &  x638 &  x659 &  x668 &  x680 &  x686 &  x710 &  x713 &  x725 &  x734 &  x752 &  x758 &  x767 &  x773 &  x782 &  x794 &  x800 &  x803 &  x806 &  x809 &  x826 &  x827 &  x830 &  x839 &  x869 &  x884 &  x893 &  x908 &  x911 &  x917 &  x923 &  x929 &  x935 &  x941 &  x944 &  x950 &  x959 &  x962 &  x974 &  x977 &  x980 &  x986 &  x989 &  x992 &  x995 &  x1016 &  x1019 &  x1028 &  x1031 &  x1034 &  x1055 &  x1061 &  x1070 &  x1076 &  x1079 &  x1082 &  x1085 &  x1100 &  x1106 &  x1121 &  x1124 &  x1130 & ~x225 & ~x639;
assign c3136 =  x5 &  x8 &  x11 &  x17 &  x56 &  x71 &  x77 &  x86 &  x92 &  x95 &  x104 &  x128 &  x140 &  x158 &  x164 &  x173 &  x182 &  x215 &  x218 &  x236 &  x257 &  x266 &  x317 &  x322 &  x329 &  x341 &  x360 &  x361 &  x362 &  x389 &  x395 &  x399 &  x400 &  x431 &  x434 &  x438 &  x439 &  x449 &  x478 &  x479 &  x494 &  x517 &  x527 &  x542 &  x572 &  x584 &  x602 &  x611 &  x701 &  x713 &  x719 &  x746 &  x752 &  x755 &  x776 &  x785 &  x788 &  x800 &  x803 &  x827 &  x830 &  x833 &  x848 &  x854 &  x884 &  x893 &  x908 &  x944 &  x950 &  x968 &  x974 &  x980 &  x983 &  x1028 &  x1031 &  x1097 & ~x162 & ~x240 & ~x993;
assign c3138 =  x11 &  x44 &  x50 &  x71 &  x98 &  x176 &  x230 &  x236 &  x239 &  x285 &  x286 &  x395 &  x403 &  x404 &  x433 &  x437 &  x464 &  x479 &  x506 &  x518 &  x533 &  x539 &  x575 &  x635 &  x650 &  x656 &  x683 &  x731 &  x755 &  x767 &  x824 &  x833 &  x836 &  x863 &  x865 &  x866 &  x872 &  x904 &  x908 &  x943 &  x1037 &  x1070 & ~x0 & ~x39 & ~x78 & ~x144 & ~x150 & ~x897 & ~x936 & ~x1047 & ~x1125;
assign c3140 =  x13 &  x86 &  x88 &  x95 &  x215 &  x236 &  x239 &  x296 &  x316 &  x344 &  x368 &  x386 &  x394 &  x398 &  x413 &  x431 &  x433 &  x461 &  x478 &  x494 &  x530 &  x545 &  x560 &  x563 &  x590 &  x610 &  x653 &  x656 &  x661 &  x665 &  x688 &  x710 &  x733 &  x752 &  x754 &  x772 &  x794 &  x806 &  x824 &  x860 &  x884 &  x929 &  x983 &  x1007 & ~x141;
assign c3142 =  x8 &  x52 &  x74 &  x104 &  x164 &  x272 &  x278 &  x323 &  x338 &  x393 &  x432 &  x433 &  x434 &  x476 &  x494 &  x503 &  x530 &  x533 &  x536 &  x542 &  x569 &  x581 &  x593 &  x596 &  x602 &  x605 &  x656 &  x668 &  x719 &  x722 &  x746 &  x748 &  x803 &  x854 &  x856 &  x895 &  x904 &  x922 &  x929 &  x932 &  x938 &  x968 &  x1001 &  x1058 &  x1078 &  x1085 & ~x561 & ~x639 & ~x717 & ~x742 & ~x781 & ~x859 & ~x898 & ~x975;
assign c3144 =  x35 &  x38 &  x44 &  x59 &  x74 &  x101 &  x110 &  x121 &  x122 &  x134 &  x137 &  x140 &  x164 &  x224 &  x227 &  x236 &  x257 &  x281 &  x302 &  x314 &  x315 &  x316 &  x323 &  x329 &  x354 &  x356 &  x368 &  x392 &  x394 &  x398 &  x416 &  x431 &  x432 &  x433 &  x434 &  x443 &  x473 &  x491 &  x500 &  x503 &  x509 &  x536 &  x539 &  x545 &  x551 &  x569 &  x608 &  x611 &  x614 &  x638 &  x650 &  x656 &  x662 &  x674 &  x677 &  x698 &  x701 &  x713 &  x728 &  x737 &  x755 &  x761 &  x773 &  x785 &  x812 &  x815 &  x844 &  x854 &  x860 &  x875 &  x905 &  x926 &  x944 &  x968 &  x986 &  x995 &  x1028 &  x1043 &  x1046 &  x1085 &  x1094 &  x1115 & ~x105 & ~x144 & ~x279 & ~x702 & ~x1098;
assign c3146 =  x157 &  x196 &  x365 &  x389 &  x451 &  x478 &  x481 &  x517 &  x526 &  x533 &  x556 &  x565 &  x598 &  x604 &  x643 &  x1129 & ~x162;
assign c3148 =  x8 &  x17 &  x38 &  x44 &  x56 &  x71 &  x74 &  x89 &  x92 &  x104 &  x136 &  x137 &  x161 &  x188 &  x206 &  x215 &  x236 &  x251 &  x275 &  x308 &  x335 &  x338 &  x344 &  x355 &  x368 &  x425 &  x431 &  x433 &  x434 &  x479 &  x488 &  x494 &  x497 &  x511 &  x550 &  x566 &  x578 &  x628 &  x656 &  x659 &  x665 &  x725 &  x752 &  x755 &  x761 &  x803 &  x815 &  x818 &  x848 &  x866 &  x869 &  x884 &  x908 &  x917 &  x932 &  x938 &  x968 &  x974 &  x1025 &  x1028 &  x1037 &  x1082 &  x1130 & ~x0 & ~x600 & ~x639 & ~x717 & ~x756 & ~x819 & ~x834 & ~x840 & ~x891 & ~x897 & ~x912 & ~x930 & ~x957 & ~x969 & ~x990 & ~x1008 & ~x1023 & ~x1029 & ~x1047 & ~x1053 & ~x1062 & ~x1068 & ~x1086;
assign c3150 =  x5 &  x13 &  x17 &  x20 &  x32 &  x38 &  x77 &  x86 &  x89 &  x125 &  x158 &  x173 &  x209 &  x215 &  x239 &  x266 &  x277 &  x305 &  x316 &  x341 &  x344 &  x433 &  x434 &  x464 &  x494 &  x518 &  x569 &  x593 &  x602 &  x631 &  x635 &  x647 &  x701 &  x752 &  x764 &  x772 &  x773 &  x815 &  x836 &  x884 &  x956 &  x989 &  x1013 &  x1016 &  x1031 &  x1037 &  x1046 & ~x27 & ~x387 & ~x702 & ~x984 & ~x1056;
assign c3152 =  x47 &  x77 &  x86 &  x104 &  x188 &  x206 &  x236 &  x263 &  x275 &  x344 &  x353 &  x410 &  x443 &  x503 &  x517 &  x548 &  x554 &  x556 &  x557 &  x575 &  x595 &  x602 &  x611 &  x634 &  x686 &  x707 &  x746 &  x752 &  x803 &  x839 &  x848 &  x932 &  x962 &  x974 &  x983 &  x995 &  x1010 &  x1082 &  x1130 & ~x153 & ~x192 & ~x423 & ~x777 & ~x855 & ~x972 & ~x1050 & ~x1089 & ~x1104;
assign c3154 =  x23 &  x62 &  x167 &  x245 &  x356 &  x380 &  x419 &  x431 &  x434 &  x497 &  x709 &  x793 &  x803 &  x805 &  x806 &  x856 &  x929 &  x959 &  x968 &  x1004 &  x1070 & ~x328 & ~x444 & ~x547 & ~x586 & ~x625 & ~x703 & ~x1095;
assign c3156 =  x23 &  x50 &  x86 &  x101 &  x134 &  x205 &  x209 &  x260 &  x277 &  x347 &  x368 &  x374 &  x383 &  x410 &  x433 &  x472 &  x539 &  x545 &  x620 &  x656 &  x662 &  x709 &  x713 &  x722 &  x739 &  x844 &  x910 &  x977 &  x983 &  x989 &  x1016 &  x1043 &  x1055 & ~x105 & ~x522 & ~x585 & ~x663 & ~x741 & ~x781 & ~x840 & ~x859 & ~x1053;
assign c3158 =  x2 &  x5 &  x8 &  x11 &  x38 &  x41 &  x44 &  x47 &  x50 &  x62 &  x71 &  x80 &  x86 &  x101 &  x104 &  x107 &  x122 &  x137 &  x140 &  x155 &  x164 &  x167 &  x185 &  x188 &  x203 &  x209 &  x230 &  x236 &  x245 &  x254 &  x263 &  x266 &  x272 &  x278 &  x281 &  x284 &  x293 &  x296 &  x311 &  x320 &  x323 &  x344 &  x347 &  x359 &  x365 &  x374 &  x383 &  x386 &  x398 &  x419 &  x422 &  x431 &  x449 &  x452 &  x455 &  x494 &  x500 &  x512 &  x539 &  x545 &  x548 &  x569 &  x581 &  x590 &  x593 &  x599 &  x608 &  x617 &  x629 &  x638 &  x656 &  x662 &  x677 &  x686 &  x710 &  x746 &  x752 &  x755 &  x758 &  x761 &  x767 &  x773 &  x787 &  x794 &  x803 &  x818 &  x826 &  x830 &  x836 &  x839 &  x842 &  x854 &  x869 &  x875 &  x884 &  x893 &  x896 &  x908 &  x911 &  x917 &  x920 &  x923 &  x929 &  x932 &  x941 &  x959 &  x968 &  x974 &  x980 &  x995 &  x1010 &  x1016 &  x1019 &  x1028 &  x1046 &  x1070 &  x1085 &  x1088 &  x1091 &  x1097 &  x1103 &  x1109 &  x1121 &  x1127 &  x1130 & ~x69 & ~x984 & ~x1005 & ~x1065 & ~x1089 & ~x1104 & ~x1128;
assign c3160 =  x1 &  x2 &  x16 &  x44 &  x50 &  x55 &  x62 &  x68 &  x71 &  x118 &  x155 &  x200 &  x236 &  x386 &  x392 &  x431 &  x451 &  x478 &  x479 &  x494 &  x517 &  x569 &  x598 &  x656 &  x755 &  x818 &  x884 &  x941 &  x977 &  x1031 & ~x279 & ~x309;
assign c3162 =  x8 &  x13 &  x51 &  x56 &  x101 &  x188 &  x236 &  x323 &  x419 &  x533 &  x591 &  x805 &  x824 &  x826 &  x844 &  x884 &  x1010 &  x1021 & ~x423 & ~x507;
assign c3164 =  x22 &  x56 &  x61 &  x73 &  x100 &  x106 &  x133 &  x139 &  x158 &  x172 &  x178 &  x185 &  x194 &  x217 &  x245 &  x250 &  x272 &  x278 &  x281 &  x290 &  x334 &  x368 &  x412 &  x451 &  x458 &  x481 &  x491 &  x503 &  x530 &  x533 &  x536 &  x539 &  x542 &  x587 &  x595 &  x608 &  x656 &  x752 &  x755 &  x790 &  x803 &  x848 &  x884 &  x893 &  x898 &  x911 &  x917 &  x925 &  x964 &  x980 &  x986 &  x1016 &  x1019 &  x1028 &  x1040 &  x1046 &  x1082;
assign c3166 =  x8 &  x23 &  x47 &  x113 &  x185 &  x207 &  x257 &  x314 &  x344 &  x356 &  x395 &  x398 &  x407 &  x464 &  x482 &  x494 &  x518 &  x587 &  x593 &  x650 &  x656 &  x704 &  x707 &  x722 &  x746 &  x752 &  x755 &  x791 &  x806 &  x827 &  x836 &  x839 &  x854 &  x871 &  x884 &  x910 &  x911 &  x917 &  x941 &  x983 &  x1070 &  x1073 &  x1088 &  x1130 & ~x262 & ~x522 & ~x600 & ~x897;
assign c3168 =  x2 &  x8 &  x44 &  x47 &  x56 &  x62 &  x68 &  x71 &  x86 &  x92 &  x101 &  x104 &  x136 &  x140 &  x148 &  x175 &  x187 &  x188 &  x275 &  x284 &  x304 &  x323 &  x331 &  x350 &  x419 &  x441 &  x442 &  x479 &  x481 &  x494 &  x521 &  x533 &  x545 &  x638 &  x644 &  x656 &  x722 &  x749 &  x773 &  x818 &  x842 &  x848 &  x854 &  x862 &  x875 &  x890 &  x899 &  x901 &  x911 &  x917 &  x946 &  x959 &  x974 &  x983 &  x998 &  x1018 &  x1085 &  x1097 &  x1130 & ~x273 & ~x390;
assign c3170 =  x1 &  x5 &  x8 &  x16 &  x55 &  x56 &  x61 &  x62 &  x71 &  x100 &  x104 &  x118 &  x139 &  x155 &  x157 &  x178 &  x188 &  x215 &  x236 &  x257 &  x281 &  x284 &  x344 &  x368 &  x386 &  x422 &  x446 &  x533 &  x545 &  x607 &  x608 &  x712 &  x746 &  x758 &  x773 &  x776 &  x803 &  x806 &  x829 &  x884 &  x917 &  x923 &  x962 &  x974 &  x1046 &  x1091 & ~x45 & ~x84 & ~x123 & ~x213 & ~x837 & ~x993 & ~x1128;
assign c3172 =  x14 &  x17 &  x44 &  x47 &  x59 &  x65 &  x68 &  x71 &  x74 &  x80 &  x95 &  x104 &  x107 &  x116 &  x122 &  x146 &  x158 &  x161 &  x164 &  x179 &  x194 &  x200 &  x203 &  x221 &  x236 &  x257 &  x263 &  x275 &  x284 &  x290 &  x296 &  x299 &  x314 &  x316 &  x323 &  x332 &  x356 &  x368 &  x383 &  x404 &  x428 &  x430 &  x431 &  x433 &  x434 &  x440 &  x449 &  x458 &  x464 &  x472 &  x482 &  x485 &  x494 &  x503 &  x508 &  x509 &  x511 &  x518 &  x533 &  x536 &  x542 &  x548 &  x566 &  x569 &  x578 &  x586 &  x590 &  x599 &  x605 &  x611 &  x623 &  x625 &  x628 &  x629 &  x632 &  x638 &  x659 &  x665 &  x667 &  x680 &  x689 &  x734 &  x737 &  x745 &  x779 &  x800 &  x806 &  x809 &  x812 &  x818 &  x821 &  x824 &  x829 &  x833 &  x842 &  x845 &  x848 &  x854 &  x860 &  x866 &  x881 &  x890 &  x911 &  x917 &  x932 &  x944 &  x953 &  x968 &  x971 &  x974 &  x977 &  x992 &  x995 &  x1004 &  x1013 &  x1043 &  x1049 &  x1082 &  x1091 &  x1124 &  x1130 & ~x492 & ~x513 & ~x522 & ~x561 & ~x600 & ~x717 & ~x765;
assign c3174 =  x1 &  x8 &  x16 &  x55 &  x61 &  x71 &  x79 &  x92 &  x100 &  x118 &  x133 &  x137 &  x145 &  x157 &  x164 &  x172 &  x184 &  x185 &  x211 &  x217 &  x242 &  x250 &  x347 &  x368 &  x404 &  x434 &  x455 &  x479 &  x482 &  x494 &  x539 &  x607 &  x656 &  x752 &  x818 &  x851 &  x884 &  x917 &  x992 &  x1082 &  x1097 & ~x36 & ~x69 & ~x264 & ~x1089 & ~x1104 & ~x1122 & ~x1128;
assign c3176 =  x8 &  x17 &  x20 &  x29 &  x59 &  x71 &  x74 &  x77 &  x92 &  x125 &  x128 &  x137 &  x146 &  x158 &  x161 &  x188 &  x200 &  x203 &  x224 &  x230 &  x236 &  x245 &  x269 &  x278 &  x296 &  x305 &  x322 &  x324 &  x326 &  x329 &  x332 &  x338 &  x356 &  x359 &  x363 &  x365 &  x368 &  x374 &  x380 &  x383 &  x392 &  x394 &  x398 &  x403 &  x404 &  x425 &  x431 &  x433 &  x434 &  x437 &  x443 &  x446 &  x449 &  x464 &  x467 &  x470 &  x472 &  x473 &  x476 &  x479 &  x482 &  x500 &  x508 &  x511 &  x515 &  x533 &  x554 &  x560 &  x566 &  x584 &  x590 &  x608 &  x617 &  x620 &  x626 &  x629 &  x632 &  x638 &  x653 &  x656 &  x659 &  x667 &  x686 &  x692 &  x698 &  x701 &  x706 &  x710 &  x713 &  x746 &  x752 &  x755 &  x797 &  x818 &  x839 &  x848 &  x854 &  x857 &  x875 &  x881 &  x890 &  x893 &  x917 &  x929 &  x953 &  x959 &  x968 &  x980 &  x983 &  x986 &  x1004 &  x1007 &  x1016 &  x1064 &  x1070 &  x1091 &  x1109 & ~x417;
assign c3178 =  x44 &  x56 &  x71 &  x89 &  x92 &  x98 &  x116 &  x125 &  x137 &  x146 &  x155 &  x170 &  x194 &  x203 &  x209 &  x215 &  x236 &  x245 &  x251 &  x257 &  x275 &  x308 &  x332 &  x344 &  x350 &  x359 &  x386 &  x458 &  x467 &  x479 &  x494 &  x509 &  x521 &  x533 &  x536 &  x545 &  x584 &  x587 &  x626 &  x629 &  x632 &  x644 &  x650 &  x698 &  x701 &  x746 &  x752 &  x755 &  x785 &  x809 &  x812 &  x823 &  x830 &  x848 &  x854 &  x866 &  x884 &  x890 &  x901 &  x920 &  x929 &  x935 &  x943 &  x965 &  x974 &  x977 &  x981 &  x983 &  x1016 &  x1018 &  x1020 &  x1025 &  x1052 &  x1082 &  x1091 &  x1103 &  x1130 & ~x39 & ~x117 & ~x273 & ~x423 & ~x792 & ~x873 & ~x912;
assign c3180 =  x11 &  x17 &  x23 &  x89 &  x92 &  x107 &  x119 &  x125 &  x134 &  x161 &  x173 &  x212 &  x215 &  x238 &  x245 &  x251 &  x254 &  x257 &  x287 &  x290 &  x317 &  x356 &  x365 &  x368 &  x383 &  x394 &  x404 &  x419 &  x425 &  x472 &  x497 &  x512 &  x515 &  x539 &  x542 &  x605 &  x611 &  x632 &  x647 &  x653 &  x671 &  x674 &  x688 &  x715 &  x716 &  x727 &  x728 &  x752 &  x754 &  x755 &  x761 &  x770 &  x773 &  x787 &  x800 &  x805 &  x812 &  x863 &  x893 &  x899 &  x910 &  x917 &  x920 &  x950 &  x959 &  x986 &  x1010 &  x1013 &  x1043 &  x1127 &  x1130 & ~x105 & ~x639 & ~x717 & ~x969 & ~x1008 & ~x1086;
assign c3182 =  x17 &  x50 &  x53 &  x62 &  x68 &  x71 &  x86 &  x89 &  x92 &  x101 &  x128 &  x164 &  x188 &  x197 &  x200 &  x205 &  x211 &  x230 &  x236 &  x244 &  x250 &  x257 &  x259 &  x275 &  x296 &  x322 &  x328 &  x347 &  x361 &  x368 &  x374 &  x392 &  x394 &  x404 &  x407 &  x410 &  x431 &  x433 &  x434 &  x446 &  x469 &  x472 &  x473 &  x494 &  x503 &  x533 &  x628 &  x638 &  x659 &  x667 &  x692 &  x706 &  x728 &  x745 &  x746 &  x748 &  x755 &  x773 &  x787 &  x803 &  x815 &  x826 &  x848 &  x854 &  x862 &  x884 &  x893 &  x902 &  x917 &  x932 &  x941 &  x968 &  x983 &  x998 &  x1010 &  x1013 &  x1028 &  x1082;
assign c3184 =  x8 &  x17 &  x62 &  x104 &  x257 &  x368 &  x404 &  x413 &  x431 &  x434 &  x490 &  x533 &  x536 &  x551 &  x554 &  x556 &  x595 &  x632 &  x634 &  x653 &  x848 &  x890 &  x962 &  x983 &  x1001 &  x1028 & ~x207 & ~x954 & ~x993 & ~x1029 & ~x1032 & ~x1089;
assign c3186 =  x5 &  x17 &  x38 &  x53 &  x56 &  x86 &  x89 &  x101 &  x188 &  x200 &  x215 &  x248 &  x257 &  x296 &  x431 &  x500 &  x548 &  x560 &  x605 &  x629 &  x632 &  x659 &  x680 &  x725 &  x746 &  x764 &  x770 &  x806 &  x812 &  x848 &  x854 &  x898 &  x976 &  x983 &  x989 &  x992 &  x1015 &  x1016 &  x1018 &  x1019 &  x1031 &  x1057 &  x1079 &  x1093 &  x1096 &  x1097 & ~x954 & ~x987 & ~x993 & ~x1032 & ~x1072 & ~x1078 & ~x1111 & ~x1116 & ~x1122;
assign c3188 =  x1 &  x38 &  x79 &  x92 &  x104 &  x118 &  x157 &  x164 &  x188 &  x257 &  x323 &  x433 &  x527 &  x557 &  x656 &  x724 &  x746 &  x1082 & ~x69 & ~x588 & ~x870 & ~x909 & ~x948 & ~x987 & ~x1026 & ~x1065 & ~x1104;
assign c3190 =  x77 &  x92 &  x101 &  x113 &  x179 &  x230 &  x233 &  x236 &  x331 &  x350 &  x374 &  x398 &  x446 &  x448 &  x451 &  x481 &  x490 &  x494 &  x526 &  x529 &  x545 &  x568 &  x581 &  x598 &  x607 &  x620 &  x632 &  x637 &  x680 &  x746 &  x839 &  x851 &  x904 &  x946 &  x965 &  x979 &  x985 &  x1018 &  x1037 &  x1055 &  x1097 &  x1112;
assign c3192 =  x14 &  x20 &  x26 &  x38 &  x47 &  x50 &  x53 &  x62 &  x71 &  x86 &  x98 &  x101 &  x104 &  x107 &  x110 &  x140 &  x143 &  x155 &  x161 &  x164 &  x170 &  x173 &  x176 &  x182 &  x209 &  x227 &  x236 &  x239 &  x245 &  x254 &  x269 &  x278 &  x281 &  x284 &  x302 &  x308 &  x314 &  x326 &  x341 &  x344 &  x347 &  x359 &  x365 &  x371 &  x383 &  x407 &  x410 &  x428 &  x431 &  x433 &  x437 &  x443 &  x449 &  x461 &  x488 &  x497 &  x503 &  x515 &  x518 &  x533 &  x536 &  x539 &  x542 &  x550 &  x551 &  x557 &  x563 &  x566 &  x581 &  x587 &  x589 &  x590 &  x593 &  x596 &  x599 &  x602 &  x608 &  x614 &  x617 &  x620 &  x626 &  x628 &  x632 &  x641 &  x647 &  x656 &  x659 &  x671 &  x677 &  x689 &  x692 &  x695 &  x698 &  x701 &  x713 &  x722 &  x725 &  x731 &  x734 &  x740 &  x745 &  x746 &  x755 &  x758 &  x776 &  x779 &  x791 &  x794 &  x797 &  x800 &  x803 &  x809 &  x821 &  x854 &  x860 &  x862 &  x863 &  x872 &  x875 &  x878 &  x887 &  x899 &  x901 &  x908 &  x911 &  x920 &  x926 &  x929 &  x935 &  x953 &  x956 &  x968 &  x977 &  x992 &  x998 &  x1007 &  x1013 &  x1016 &  x1025 &  x1031 &  x1040 &  x1058 &  x1076 &  x1082 &  x1127 &  x1130 & ~x105 & ~x144 & ~x417 & ~x792 & ~x831 & ~x870 & ~x909 & ~x948 & ~x987 & ~x1026 & ~x1065 & ~x1104;
assign c3194 =  x17 &  x26 &  x32 &  x62 &  x71 &  x86 &  x89 &  x98 &  x125 &  x140 &  x155 &  x164 &  x182 &  x188 &  x197 &  x203 &  x212 &  x224 &  x236 &  x239 &  x263 &  x272 &  x290 &  x314 &  x344 &  x347 &  x350 &  x365 &  x368 &  x371 &  x383 &  x434 &  x440 &  x443 &  x460 &  x461 &  x464 &  x467 &  x470 &  x482 &  x494 &  x503 &  x512 &  x530 &  x533 &  x536 &  x545 &  x548 &  x554 &  x560 &  x566 &  x569 &  x575 &  x608 &  x611 &  x638 &  x656 &  x677 &  x680 &  x698 &  x728 &  x746 &  x749 &  x752 &  x770 &  x815 &  x824 &  x848 &  x861 &  x863 &  x866 &  x884 &  x899 &  x900 &  x901 &  x914 &  x929 &  x944 &  x947 &  x965 &  x968 &  x974 &  x979 &  x980 &  x986 &  x995 &  x998 &  x1010 &  x1031 &  x1037 &  x1043 &  x1046 &  x1055 &  x1057 &  x1060 &  x1067 &  x1073 &  x1082 &  x1091 &  x1100 &  x1103 &  x1127 &  x1130 & ~x243 & ~x333 & ~x390 & ~x468 & ~x951 & ~x957 & ~x990 & ~x1074 & ~x1113;
assign c3196 =  x38 &  x236 &  x257 &  x281 &  x326 &  x353 &  x362 &  x365 &  x386 &  x407 &  x425 &  x440 &  x529 &  x554 &  x584 &  x637 &  x644 &  x761 &  x803 &  x842 &  x846 &  x892 &  x899 &  x908 &  x923 &  x926 &  x935 &  x950 &  x962 &  x964 &  x983 &  x1016 &  x1040 & ~x1104;
assign c3198 =  x8 &  x11 &  x14 &  x38 &  x65 &  x74 &  x80 &  x89 &  x92 &  x98 &  x101 &  x104 &  x113 &  x140 &  x164 &  x182 &  x185 &  x188 &  x191 &  x200 &  x203 &  x215 &  x236 &  x248 &  x275 &  x278 &  x284 &  x296 &  x305 &  x308 &  x311 &  x314 &  x320 &  x323 &  x325 &  x331 &  x344 &  x356 &  x374 &  x398 &  x403 &  x404 &  x419 &  x422 &  x431 &  x434 &  x443 &  x445 &  x452 &  x455 &  x461 &  x473 &  x476 &  x479 &  x481 &  x484 &  x494 &  x497 &  x500 &  x503 &  x521 &  x536 &  x548 &  x554 &  x559 &  x569 &  x595 &  x605 &  x608 &  x628 &  x629 &  x632 &  x647 &  x650 &  x656 &  x667 &  x677 &  x686 &  x689 &  x701 &  x710 &  x713 &  x734 &  x746 &  x752 &  x764 &  x773 &  x776 &  x791 &  x803 &  x815 &  x818 &  x827 &  x839 &  x861 &  x875 &  x884 &  x900 &  x901 &  x908 &  x911 &  x923 &  x932 &  x939 &  x941 &  x962 &  x977 &  x978 &  x986 &  x995 &  x1018 &  x1028 &  x1046 &  x1057 &  x1061 &  x1070 &  x1076 &  x1088 &  x1091 &  x1096 &  x1097 &  x1115 &  x1124 &  x1130 & ~x273 & ~x351 & ~x390 & ~x468 & ~x507;
assign c3200 =  x5 &  x32 &  x38 &  x41 &  x59 &  x62 &  x68 &  x71 &  x86 &  x110 &  x113 &  x122 &  x128 &  x161 &  x185 &  x188 &  x194 &  x215 &  x227 &  x239 &  x281 &  x287 &  x335 &  x344 &  x356 &  x365 &  x371 &  x374 &  x377 &  x401 &  x413 &  x425 &  x479 &  x494 &  x503 &  x527 &  x563 &  x578 &  x590 &  x614 &  x662 &  x677 &  x686 &  x698 &  x710 &  x713 &  x719 &  x740 &  x743 &  x749 &  x797 &  x806 &  x830 &  x848 &  x851 &  x914 &  x923 &  x950 &  x971 &  x1046 &  x1079 &  x1082 &  x1088 &  x1106 &  x1109 &  x1115 & ~x30 & ~x69 & ~x804 & ~x834 & ~x873 & ~x912 & ~x913 & ~x951 & ~x952 & ~x990 & ~x991 & ~x993 & ~x1026 & ~x1029 & ~x1032;
assign c3202 =  x182 &  x184 &  x200 &  x203 &  x257 &  x307 &  x373 &  x404 &  x419 &  x481 &  x521 &  x533 &  x546 &  x566 &  x624 &  x625 &  x629 &  x703 &  x725 &  x830 &  x887 &  x908 &  x983 &  x1019 &  x1049 &  x1070 &  x1130 & ~x993 & ~x1104;
assign c3204 =  x8 &  x17 &  x92 &  x182 &  x236 &  x368 &  x404 &  x431 &  x479 &  x494 &  x518 &  x527 &  x590 &  x604 &  x686 &  x776 &  x815 &  x818 &  x823 &  x901 &  x939 &  x968 &  x978 &  x1017 &  x1018 &  x1088 &  x1096 &  x1121 & ~x321 & ~x429 & ~x468 & ~x507 & ~x651 & ~x1128;
assign c3206 =  x1 &  x17 &  x74 &  x86 &  x92 &  x143 &  x155 &  x164 &  x188 &  x236 &  x272 &  x275 &  x287 &  x296 &  x323 &  x350 &  x359 &  x377 &  x383 &  x386 &  x425 &  x431 &  x434 &  x461 &  x488 &  x491 &  x535 &  x554 &  x556 &  x574 &  x593 &  x595 &  x607 &  x613 &  x631 &  x656 &  x701 &  x704 &  x743 &  x752 &  x754 &  x764 &  x803 &  x806 &  x847 &  x872 &  x884 &  x908 &  x920 &  x946 &  x962 &  x985 &  x998 &  x1010 &  x1016 &  x1028 &  x1040 &  x1048 &  x1058 &  x1076 &  x1130 & ~x141;
assign c3208 =  x5 &  x17 &  x41 &  x47 &  x55 &  x71 &  x95 &  x137 &  x140 &  x157 &  x185 &  x200 &  x218 &  x236 &  x244 &  x248 &  x260 &  x266 &  x277 &  x281 &  x284 &  x287 &  x290 &  x316 &  x323 &  x338 &  x359 &  x368 &  x371 &  x386 &  x394 &  x404 &  x407 &  x419 &  x431 &  x433 &  x434 &  x464 &  x470 &  x476 &  x488 &  x503 &  x521 &  x527 &  x533 &  x554 &  x560 &  x575 &  x593 &  x626 &  x650 &  x656 &  x659 &  x674 &  x709 &  x716 &  x719 &  x727 &  x739 &  x746 &  x752 &  x755 &  x770 &  x778 &  x791 &  x817 &  x827 &  x833 &  x842 &  x845 &  x848 &  x851 &  x856 &  x872 &  x884 &  x905 &  x920 &  x929 &  x934 &  x941 &  x962 &  x965 &  x974 &  x989 &  x998 &  x1016 &  x1043 &  x1130 & ~x339 & ~x663;
assign c3210 =  x2 &  x5 &  x8 &  x17 &  x36 &  x37 &  x38 &  x44 &  x56 &  x92 &  x155 &  x184 &  x212 &  x236 &  x239 &  x257 &  x263 &  x305 &  x311 &  x343 &  x344 &  x368 &  x398 &  x413 &  x431 &  x434 &  x479 &  x484 &  x509 &  x530 &  x545 &  x605 &  x623 &  x629 &  x689 &  x698 &  x719 &  x746 &  x752 &  x803 &  x860 &  x884 &  x914 &  x917 &  x938 &  x944 &  x974 &  x983 &  x1010 &  x1052 &  x1082 &  x1094 &  x1100 &  x1115 & ~x162 & ~x198;
assign c3212 =  x20 &  x56 &  x59 &  x148 &  x173 &  x191 &  x203 &  x242 &  x257 &  x263 &  x331 &  x413 &  x416 &  x431 &  x455 &  x481 &  x494 &  x536 &  x545 &  x643 &  x662 &  x668 &  x677 &  x680 &  x682 &  x701 &  x746 &  x752 &  x761 &  x764 &  x803 &  x809 &  x818 &  x823 &  x862 &  x911 &  x917 &  x983 &  x1018 &  x1019 &  x1028 &  x1043 &  x1070 &  x1079 &  x1112 & ~x507 & ~x873 & ~x912 & ~x1074;
assign c3214 =  x17 &  x47 &  x53 &  x68 &  x92 &  x104 &  x164 &  x218 &  x230 &  x236 &  x257 &  x331 &  x374 &  x404 &  x431 &  x479 &  x500 &  x524 &  x533 &  x566 &  x605 &  x650 &  x656 &  x680 &  x752 &  x761 &  x797 &  x848 &  x854 &  x862 &  x899 &  x901 &  x917 &  x950 &  x980 &  x989 &  x998 &  x1016 &  x1028 &  x1061 &  x1070 &  x1082 &  x1091 & ~x0 & ~x39 & ~x60 & ~x117 & ~x150 & ~x165 & ~x195 & ~x957 & ~x1074 & ~x1092 & ~x1128;
assign c3216 =  x8 &  x23 &  x44 &  x71 &  x73 &  x98 &  x101 &  x107 &  x110 &  x131 &  x134 &  x145 &  x164 &  x184 &  x188 &  x194 &  x236 &  x245 &  x257 &  x269 &  x272 &  x290 &  x296 &  x299 &  x311 &  x320 &  x326 &  x368 &  x371 &  x386 &  x392 &  x403 &  x434 &  x442 &  x461 &  x473 &  x476 &  x479 &  x481 &  x521 &  x533 &  x554 &  x560 &  x587 &  x593 &  x602 &  x605 &  x626 &  x662 &  x698 &  x719 &  x731 &  x752 &  x755 &  x836 &  x857 &  x862 &  x863 &  x901 &  x953 &  x962 &  x968 &  x992 &  x995 &  x1007 &  x1028 &  x1031 &  x1037 &  x1043 &  x1082 &  x1121 & ~x648 & ~x649 & ~x687 & ~x726 & ~x765;
assign c3218 =  x5 &  x8 &  x11 &  x17 &  x20 &  x23 &  x32 &  x35 &  x38 &  x44 &  x47 &  x50 &  x56 &  x62 &  x68 &  x71 &  x80 &  x83 &  x86 &  x89 &  x92 &  x95 &  x101 &  x104 &  x107 &  x113 &  x122 &  x128 &  x134 &  x137 &  x140 &  x164 &  x182 &  x185 &  x188 &  x194 &  x197 &  x200 &  x203 &  x206 &  x209 &  x212 &  x221 &  x230 &  x236 &  x242 &  x251 &  x257 &  x260 &  x269 &  x281 &  x284 &  x290 &  x296 &  x305 &  x308 &  x321 &  x322 &  x323 &  x326 &  x332 &  x338 &  x341 &  x344 &  x347 &  x353 &  x359 &  x361 &  x362 &  x365 &  x368 &  x371 &  x383 &  x389 &  x395 &  x400 &  x401 &  x404 &  x416 &  x422 &  x428 &  x431 &  x433 &  x434 &  x443 &  x452 &  x461 &  x464 &  x467 &  x473 &  x479 &  x491 &  x497 &  x500 &  x503 &  x506 &  x508 &  x509 &  x518 &  x521 &  x524 &  x533 &  x545 &  x547 &  x551 &  x554 &  x560 &  x566 &  x569 &  x572 &  x584 &  x590 &  x593 &  x596 &  x599 &  x602 &  x608 &  x629 &  x641 &  x644 &  x647 &  x653 &  x659 &  x665 &  x667 &  x692 &  x698 &  x701 &  x713 &  x725 &  x743 &  x746 &  x752 &  x755 &  x758 &  x761 &  x773 &  x785 &  x803 &  x806 &  x815 &  x827 &  x845 &  x857 &  x860 &  x866 &  x869 &  x875 &  x878 &  x881 &  x884 &  x893 &  x899 &  x902 &  x904 &  x908 &  x911 &  x917 &  x929 &  x932 &  x943 &  x947 &  x953 &  x965 &  x968 &  x971 &  x983 &  x989 &  x992 &  x995 &  x998 &  x1010 &  x1016 &  x1021 &  x1022 &  x1031 &  x1040 &  x1043 &  x1046 &  x1049 &  x1058 &  x1070 &  x1073 &  x1076 &  x1082 &  x1091 &  x1103 &  x1109 &  x1118 &  x1121 &  x1130 & ~x273 & ~x492 & ~x639;
assign c3220 =  x2 &  x11 &  x17 &  x29 &  x47 &  x56 &  x71 &  x74 &  x77 &  x80 &  x92 &  x101 &  x104 &  x110 &  x137 &  x140 &  x155 &  x164 &  x188 &  x197 &  x200 &  x206 &  x215 &  x236 &  x257 &  x260 &  x263 &  x275 &  x281 &  x284 &  x296 &  x323 &  x344 &  x368 &  x371 &  x386 &  x389 &  x392 &  x422 &  x431 &  x434 &  x443 &  x448 &  x455 &  x458 &  x460 &  x464 &  x479 &  x485 &  x488 &  x494 &  x500 &  x521 &  x533 &  x539 &  x545 &  x554 &  x566 &  x569 &  x593 &  x602 &  x604 &  x605 &  x629 &  x632 &  x643 &  x644 &  x682 &  x710 &  x719 &  x721 &  x728 &  x746 &  x752 &  x755 &  x767 &  x776 &  x791 &  x800 &  x803 &  x806 &  x812 &  x821 &  x823 &  x827 &  x845 &  x848 &  x854 &  x872 &  x884 &  x893 &  x898 &  x899 &  x901 &  x923 &  x929 &  x932 &  x944 &  x962 &  x976 &  x983 &  x992 &  x995 &  x1010 &  x1015 &  x1018 &  x1034 &  x1040 &  x1046 &  x1057 &  x1082 &  x1085 &  x1088 &  x1093 &  x1096 &  x1115 &  x1130 & ~x651 & ~x825 & ~x873 & ~x912 & ~x1029;
assign c3222 =  x200 &  x236 &  x278 &  x383 &  x395 &  x443 &  x451 &  x476 &  x482 &  x500 &  x536 &  x542 &  x548 &  x629 &  x707 &  x725 &  x752 &  x842 &  x848 &  x887 &  x920 &  x929 &  x1018 &  x1057 &  x1093 &  x1096 & ~x69 & ~x699 & ~x993 & ~x1006;
assign c3224 =  x2 &  x5 &  x8 &  x17 &  x38 &  x44 &  x68 &  x74 &  x98 &  x128 &  x131 &  x164 &  x188 &  x209 &  x215 &  x236 &  x277 &  x281 &  x365 &  x368 &  x374 &  x383 &  x419 &  x422 &  x431 &  x434 &  x455 &  x479 &  x482 &  x494 &  x506 &  x512 &  x514 &  x533 &  x539 &  x545 &  x548 &  x554 &  x566 &  x590 &  x605 &  x608 &  x611 &  x631 &  x632 &  x638 &  x649 &  x656 &  x680 &  x686 &  x689 &  x709 &  x710 &  x727 &  x728 &  x734 &  x740 &  x746 &  x752 &  x755 &  x764 &  x766 &  x773 &  x805 &  x809 &  x827 &  x830 &  x836 &  x839 &  x848 &  x854 &  x860 &  x917 &  x941 &  x944 &  x962 &  x983 &  x992 &  x995 &  x1010 &  x1019 &  x1031 &  x1061 &  x1070 &  x1079 &  x1100 &  x1118 &  x1124 & ~x429 & ~x468 & ~x507 & ~x508 & ~x547 & ~x585 & ~x586 & ~x624 & ~x625 & ~x664 & ~x703 & ~x742 & ~x780 & ~x897 & ~x984;
assign c3226 =  x118 &  x157 &  x164 &  x236 &  x278 &  x323 &  x329 &  x356 &  x556 &  x595 &  x616 &  x626 &  x634 &  x944 &  x992 &  x1013 & ~x96 & ~x162 & ~x180 & ~x837 & ~x1089 & ~x1104;
assign c3228 =  x25 &  x61 &  x88 &  x100 &  x137 &  x244 &  x308 &  x478 &  x517 &  x545 &  x613 &  x689 &  x713 &  x772 &  x776 &  x884 &  x943 &  x961 &  x1045;
assign c3230 =  x100 &  x178 &  x194 &  x197 &  x205 &  x244 &  x275 &  x278 &  x317 &  x321 &  x322 &  x344 &  x407 &  x449 &  x508 &  x628 &  x632 &  x653 &  x656 &  x712 &  x836 &  x884 &  x1034 &  x1040 &  x1085 &  x1106 & ~x456;
assign c3232 =  x1 &  x2 &  x11 &  x20 &  x29 &  x38 &  x53 &  x62 &  x65 &  x68 &  x71 &  x101 &  x104 &  x113 &  x119 &  x128 &  x134 &  x146 &  x152 &  x182 &  x185 &  x191 &  x194 &  x200 &  x209 &  x215 &  x218 &  x236 &  x239 &  x242 &  x248 &  x251 &  x260 &  x263 &  x266 &  x272 &  x275 &  x277 &  x281 &  x287 &  x290 &  x293 &  x296 &  x302 &  x316 &  x317 &  x320 &  x326 &  x329 &  x332 &  x335 &  x341 &  x356 &  x368 &  x371 &  x374 &  x377 &  x394 &  x398 &  x404 &  x410 &  x428 &  x431 &  x433 &  x434 &  x449 &  x452 &  x473 &  x482 &  x494 &  x497 &  x506 &  x512 &  x524 &  x548 &  x551 &  x560 &  x566 &  x569 &  x575 &  x578 &  x596 &  x607 &  x635 &  x653 &  x659 &  x698 &  x719 &  x728 &  x746 &  x752 &  x755 &  x761 &  x776 &  x791 &  x797 &  x800 &  x812 &  x818 &  x824 &  x827 &  x830 &  x836 &  x845 &  x848 &  x854 &  x857 &  x875 &  x884 &  x890 &  x895 &  x899 &  x908 &  x911 &  x917 &  x929 &  x934 &  x941 &  x962 &  x965 &  x968 &  x977 &  x983 &  x992 &  x1004 &  x1028 &  x1046 &  x1052 &  x1061 &  x1064 &  x1076 &  x1085 &  x1091 &  x1103 &  x1112 &  x1118 & ~x69 & ~x870 & ~x909 & ~x987 & ~x1026 & ~x1065 & ~x1104;
assign c3234 =  x2 &  x8 &  x17 &  x41 &  x56 &  x68 &  x71 &  x74 &  x86 &  x89 &  x92 &  x101 &  x104 &  x110 &  x119 &  x128 &  x134 &  x137 &  x167 &  x197 &  x203 &  x221 &  x236 &  x250 &  x275 &  x288 &  x320 &  x323 &  x324 &  x325 &  x328 &  x335 &  x344 &  x365 &  x368 &  x419 &  x431 &  x433 &  x434 &  x455 &  x494 &  x521 &  x530 &  x545 &  x548 &  x554 &  x560 &  x563 &  x590 &  x596 &  x602 &  x628 &  x656 &  x659 &  x680 &  x701 &  x706 &  x752 &  x755 &  x770 &  x773 &  x776 &  x803 &  x806 &  x812 &  x845 &  x848 &  x854 &  x860 &  x869 &  x875 &  x899 &  x901 &  x908 &  x941 &  x968 &  x974 &  x983 &  x1019 &  x1028 &  x1040 &  x1061 &  x1067 &  x1103 &  x1121 & ~x273;
assign c3236 =  x269 &  x368 &  x416 &  x425 &  x513 &  x514 &  x584 &  x599 &  x641 &  x661 &  x754 &  x839 &  x884 &  x1067 & ~x367 & ~x664 & ~x742 & ~x1056;
assign c3238 =  x1 &  x8 &  x40 &  x50 &  x56 &  x71 &  x79 &  x86 &  x88 &  x92 &  x101 &  x110 &  x113 &  x118 &  x137 &  x143 &  x157 &  x164 &  x166 &  x176 &  x185 &  x188 &  x194 &  x205 &  x230 &  x233 &  x244 &  x245 &  x251 &  x257 &  x266 &  x275 &  x281 &  x296 &  x322 &  x323 &  x356 &  x359 &  x361 &  x362 &  x368 &  x380 &  x383 &  x400 &  x422 &  x425 &  x431 &  x433 &  x434 &  x438 &  x439 &  x440 &  x446 &  x472 &  x478 &  x479 &  x488 &  x494 &  x517 &  x521 &  x533 &  x542 &  x545 &  x548 &  x554 &  x556 &  x560 &  x575 &  x578 &  x595 &  x602 &  x608 &  x632 &  x638 &  x656 &  x668 &  x683 &  x695 &  x698 &  x713 &  x734 &  x746 &  x752 &  x764 &  x767 &  x788 &  x791 &  x803 &  x827 &  x845 &  x851 &  x863 &  x884 &  x914 &  x929 &  x959 &  x968 &  x974 &  x983 &  x986 &  x1010 &  x1019 &  x1028 &  x1073 &  x1082 & ~x84 & ~x123;
assign c3240 =  x236 &  x481 &  x605 &  x731 &  x806 &  x839 &  x868 &  x938 &  x945 &  x985 &  x1082 &  x1096 &  x1112 & ~x390 & ~x729 & ~x768 & ~x990;
assign c3242 =  x8 &  x13 &  x50 &  x81 &  x86 &  x120 &  x137 &  x200 &  x263 &  x277 &  x394 &  x433 &  x482 &  x521 &  x701 &  x761 &  x803 &  x805 &  x844 &  x848 &  x877 &  x887 &  x974 &  x1004 & ~x366 & ~x405 & ~x586 & ~x625 & ~x664 & ~x703 & ~x1092;
assign c3244 =  x2 &  x11 &  x71 &  x101 &  x155 &  x173 &  x215 &  x230 &  x281 &  x296 &  x374 &  x407 &  x433 &  x472 &  x494 &  x503 &  x533 &  x653 &  x656 &  x662 &  x680 &  x708 &  x709 &  x737 &  x746 &  x748 &  x778 &  x800 &  x857 &  x917 &  x1073 & ~x642 & ~x780 & ~x1104;
assign c3246 =  x116 &  x205 &  x272 &  x277 &  x323 &  x365 &  x404 &  x437 &  x470 &  x479 &  x563 &  x569 &  x611 &  x628 &  x830 &  x893 &  x959 &  x962 &  x1121 & ~x300 & ~x339 & ~x417 & ~x418 & ~x885 & ~x1029;
assign c3248 =  x16 &  x17 &  x29 &  x161 &  x188 &  x322 &  x438 &  x439 &  x478 &  x539 &  x745 &  x751 &  x828 &  x829 &  x907;
assign c3250 =  x1 &  x8 &  x17 &  x38 &  x44 &  x92 &  x101 &  x118 &  x157 &  x161 &  x164 &  x188 &  x236 &  x260 &  x323 &  x344 &  x383 &  x434 &  x494 &  x607 &  x656 &  x659 &  x685 &  x691 &  x746 &  x803 &  x808 &  x847 &  x854 &  x884 &  x956 &  x968 &  x983 &  x1046 &  x1100 & ~x84 & ~x96 & ~x123 & ~x837 & ~x1065 & ~x1089;
assign c3252 =  x80 &  x188 &  x199 &  x236 &  x368 &  x431 &  x433 &  x545 &  x752 &  x884 &  x935 &  x983 & ~x33 & ~x57 & ~x66 & ~x105 & ~x144 & ~x261 & ~x301 & ~x339 & ~x639;
assign c3254 =  x8 &  x13 &  x68 &  x88 &  x95 &  x98 &  x134 &  x157 &  x161 &  x164 &  x188 &  x196 &  x254 &  x277 &  x278 &  x296 &  x314 &  x335 &  x368 &  x422 &  x433 &  x434 &  x500 &  x533 &  x539 &  x551 &  x552 &  x587 &  x631 &  x632 &  x656 &  x665 &  x670 &  x746 &  x752 &  x773 &  x805 &  x815 &  x836 &  x850 &  x908 &  x910 &  x935 &  x974 &  x1040 &  x1079 &  x1082 &  x1097 & ~x507 & ~x780;
assign c3256 =  x5 &  x17 &  x23 &  x26 &  x29 &  x32 &  x41 &  x47 &  x53 &  x56 &  x65 &  x68 &  x98 &  x104 &  x113 &  x125 &  x134 &  x164 &  x173 &  x182 &  x188 &  x200 &  x203 &  x215 &  x233 &  x251 &  x257 &  x263 &  x272 &  x284 &  x290 &  x305 &  x317 &  x325 &  x332 &  x350 &  x356 &  x359 &  x364 &  x368 &  x374 &  x389 &  x401 &  x403 &  x425 &  x434 &  x442 &  x446 &  x448 &  x455 &  x467 &  x481 &  x482 &  x500 &  x503 &  x506 &  x518 &  x527 &  x533 &  x545 &  x548 &  x575 &  x581 &  x584 &  x587 &  x590 &  x596 &  x599 &  x602 &  x629 &  x638 &  x641 &  x650 &  x656 &  x671 &  x680 &  x689 &  x716 &  x722 &  x728 &  x731 &  x734 &  x740 &  x743 &  x746 &  x752 &  x755 &  x776 &  x797 &  x806 &  x812 &  x815 &  x827 &  x830 &  x839 &  x854 &  x860 &  x869 &  x875 &  x884 &  x901 &  x908 &  x911 &  x917 &  x920 &  x923 &  x932 &  x935 &  x940 &  x962 &  x968 &  x974 &  x979 &  x995 &  x998 &  x1007 &  x1010 &  x1016 &  x1018 &  x1019 &  x1031 &  x1037 &  x1043 &  x1049 &  x1058 &  x1082 &  x1094 &  x1103 &  x1112 &  x1115 &  x1124 & ~x351 & ~x592 & ~x630 & ~x631 & ~x870;
assign c3258 =  x8 &  x32 &  x47 &  x50 &  x53 &  x56 &  x62 &  x71 &  x74 &  x79 &  x80 &  x86 &  x101 &  x104 &  x107 &  x118 &  x121 &  x137 &  x157 &  x164 &  x170 &  x173 &  x185 &  x188 &  x191 &  x196 &  x199 &  x200 &  x209 &  x224 &  x238 &  x248 &  x257 &  x263 &  x269 &  x275 &  x277 &  x284 &  x314 &  x316 &  x323 &  x326 &  x362 &  x368 &  x371 &  x383 &  x389 &  x394 &  x404 &  x419 &  x422 &  x425 &  x431 &  x433 &  x434 &  x472 &  x473 &  x479 &  x491 &  x494 &  x500 &  x503 &  x506 &  x509 &  x514 &  x517 &  x521 &  x533 &  x545 &  x548 &  x556 &  x608 &  x632 &  x647 &  x656 &  x671 &  x680 &  x701 &  x725 &  x731 &  x746 &  x749 &  x752 &  x766 &  x776 &  x779 &  x782 &  x803 &  x805 &  x806 &  x812 &  x839 &  x844 &  x845 &  x854 &  x860 &  x884 &  x893 &  x905 &  x917 &  x929 &  x935 &  x947 &  x956 &  x961 &  x962 &  x977 &  x986 &  x995 &  x998 &  x1004 &  x1016 &  x1019 &  x1028 &  x1052 &  x1055 &  x1061 &  x1070 &  x1082 &  x1085 &  x1091 &  x1097 &  x1103 &  x1106 &  x1109 & ~x507 & ~x528;
assign c3260 =  x89 &  x314 &  x481 &  x533 &  x597 &  x598 &  x637 &  x656 &  x659 &  x706 &  x851 &  x917 &  x979 &  x1061 &  x1096 & ~x267 & ~x315 & ~x351 & ~x393 & ~x468 & ~x508;
assign c3262 =  x8 &  x17 &  x47 &  x50 &  x56 &  x62 &  x65 &  x68 &  x71 &  x83 &  x89 &  x92 &  x101 &  x104 &  x128 &  x134 &  x140 &  x161 &  x188 &  x209 &  x236 &  x257 &  x263 &  x275 &  x277 &  x281 &  x296 &  x314 &  x316 &  x317 &  x323 &  x326 &  x344 &  x350 &  x353 &  x368 &  x389 &  x392 &  x394 &  x395 &  x404 &  x407 &  x413 &  x433 &  x434 &  x452 &  x461 &  x472 &  x473 &  x494 &  x503 &  x508 &  x511 &  x539 &  x545 &  x548 &  x554 &  x566 &  x589 &  x590 &  x593 &  x608 &  x632 &  x659 &  x667 &  x686 &  x716 &  x722 &  x725 &  x743 &  x745 &  x746 &  x752 &  x755 &  x776 &  x779 &  x803 &  x818 &  x830 &  x848 &  x854 &  x857 &  x878 &  x884 &  x893 &  x901 &  x905 &  x917 &  x926 &  x929 &  x932 &  x965 &  x968 &  x977 &  x979 &  x983 &  x992 &  x998 &  x1010 &  x1018 &  x1028 &  x1061 &  x1088 &  x1097 &  x1103 &  x1106 &  x1130 & ~x600 & ~x639 & ~x717 & ~x792 & ~x834 & ~x870;
assign c3264 =  x38 &  x47 &  x68 &  x71 &  x104 &  x137 &  x155 &  x158 &  x164 &  x193 &  x194 &  x197 &  x200 &  x212 &  x215 &  x224 &  x226 &  x233 &  x245 &  x257 &  x278 &  x281 &  x287 &  x292 &  x296 &  x304 &  x310 &  x331 &  x340 &  x341 &  x344 &  x377 &  x403 &  x407 &  x416 &  x431 &  x434 &  x448 &  x479 &  x481 &  x515 &  x545 &  x548 &  x554 &  x584 &  x608 &  x638 &  x656 &  x662 &  x695 &  x701 &  x752 &  x773 &  x803 &  x806 &  x848 &  x851 &  x854 &  x857 &  x860 &  x862 &  x868 &  x884 &  x896 &  x901 &  x907 &  x944 &  x946 &  x962 &  x968 &  x980 &  x983 &  x986 &  x1018 &  x1028 &  x1061 &  x1079 &  x1084 &  x1085 &  x1118 &  x1123 &  x1130 & ~x468;
assign c3266 =  x20 &  x29 &  x47 &  x50 &  x53 &  x56 &  x89 &  x92 &  x98 &  x101 &  x104 &  x110 &  x137 &  x152 &  x155 &  x164 &  x167 &  x182 &  x185 &  x188 &  x191 &  x203 &  x215 &  x221 &  x227 &  x233 &  x236 &  x239 &  x242 &  x245 &  x254 &  x257 &  x263 &  x278 &  x290 &  x296 &  x305 &  x308 &  x335 &  x344 &  x368 &  x377 &  x392 &  x395 &  x431 &  x433 &  x437 &  x440 &  x446 &  x448 &  x455 &  x464 &  x467 &  x473 &  x479 &  x482 &  x488 &  x497 &  x500 &  x509 &  x511 &  x518 &  x530 &  x533 &  x545 &  x560 &  x569 &  x572 &  x589 &  x590 &  x608 &  x617 &  x620 &  x623 &  x632 &  x644 &  x647 &  x656 &  x671 &  x686 &  x704 &  x713 &  x728 &  x731 &  x743 &  x752 &  x755 &  x773 &  x779 &  x784 &  x785 &  x803 &  x806 &  x812 &  x821 &  x823 &  x833 &  x845 &  x854 &  x857 &  x860 &  x862 &  x872 &  x875 &  x881 &  x887 &  x896 &  x901 &  x908 &  x911 &  x968 &  x974 &  x983 &  x986 &  x989 &  x992 &  x995 &  x1001 &  x1007 &  x1037 &  x1040 &  x1043 &  x1061 &  x1064 &  x1082 &  x1085 &  x1097 & ~x78 & ~x117 & ~x195 & ~x234 & ~x273 & ~x639 & ~x648 & ~x678 & ~x687 & ~x717 & ~x726 & ~x765 & ~x804;
assign c3268 =  x14 &  x17 &  x38 &  x68 &  x71 &  x104 &  x119 &  x149 &  x182 &  x344 &  x350 &  x353 &  x359 &  x374 &  x386 &  x389 &  x407 &  x419 &  x431 &  x449 &  x454 &  x479 &  x481 &  x494 &  x506 &  x520 &  x545 &  x596 &  x602 &  x683 &  x698 &  x701 &  x749 &  x752 &  x833 &  x898 &  x901 &  x917 &  x923 &  x932 &  x937 &  x941 &  x947 &  x976 &  x977 &  x979 &  x983 &  x1018 &  x1040 &  x1043 &  x1057 &  x1079 &  x1082 &  x1096 & ~x45 & ~x123 & ~x162 & ~x237 & ~x240 & ~x804 & ~x834 & ~x873 & ~x912 & ~x951;
assign c3270 =  x1 &  x8 &  x40 &  x56 &  x61 &  x100 &  x104 &  x118 &  x157 &  x178 &  x188 &  x196 &  x217 &  x296 &  x356 &  x398 &  x431 &  x451 &  x490 &  x503 &  x529 &  x530 &  x533 &  x545 &  x568 &  x607 &  x632 &  x638 &  x656 &  x725 &  x734 &  x746 &  x752 &  x773 &  x776 &  x790 &  x812 &  x829 &  x875 &  x944 &  x968 &  x1016 &  x1031 &  x1061 &  x1082 & ~x147 & ~x240 & ~x303 & ~x342;
assign c3272 =  x5 &  x8 &  x17 &  x47 &  x50 &  x53 &  x56 &  x59 &  x65 &  x83 &  x86 &  x101 &  x107 &  x116 &  x128 &  x131 &  x149 &  x155 &  x185 &  x188 &  x200 &  x209 &  x212 &  x215 &  x230 &  x236 &  x257 &  x260 &  x263 &  x275 &  x281 &  x287 &  x292 &  x296 &  x305 &  x314 &  x347 &  x356 &  x368 &  x374 &  x398 &  x403 &  x407 &  x410 &  x422 &  x431 &  x442 &  x461 &  x467 &  x481 &  x488 &  x500 &  x503 &  x520 &  x539 &  x545 &  x548 &  x554 &  x557 &  x605 &  x632 &  x644 &  x650 &  x653 &  x659 &  x674 &  x692 &  x734 &  x740 &  x746 &  x752 &  x755 &  x767 &  x770 &  x782 &  x797 &  x803 &  x818 &  x823 &  x854 &  x862 &  x866 &  x875 &  x884 &  x896 &  x901 &  x920 &  x968 &  x983 &  x995 &  x1018 &  x1022 &  x1046 &  x1055 &  x1057 &  x1076 &  x1079 &  x1085 &  x1096 &  x1103 & ~x39 & ~x78 & ~x156 & ~x195 & ~x234 & ~x267 & ~x417 & ~x456 & ~x468 & ~x612 & ~x651;
assign c3274 =  x1 &  x38 &  x71 &  x188 &  x215 &  x317 &  x332 &  x437 &  x556 &  x746 &  x773 &  x803 &  x917 &  x962 &  x1013 &  x1082 &  x1103 & ~x31 & ~x69 & ~x102 & ~x108 & ~x816 & ~x954 & ~x993 & ~x1005 & ~x1032 & ~x1065 & ~x1089;
assign c3276 =  x5 &  x62 &  x86 &  x128 &  x146 &  x185 &  x200 &  x207 &  x215 &  x257 &  x296 &  x323 &  x368 &  x398 &  x433 &  x479 &  x494 &  x545 &  x557 &  x617 &  x628 &  x728 &  x748 &  x785 &  x825 &  x826 &  x829 &  x833 &  x836 &  x851 &  x854 &  x904 &  x968 &  x980 &  x1058 &  x1067 &  x1082 &  x1097 & ~x39 & ~x78;
assign c3278 =  x38 &  x41 &  x44 &  x68 &  x134 &  x347 &  x548 &  x560 &  x605 &  x677 &  x752 &  x767 &  x782 &  x830 &  x893 &  x902 &  x905 &  x935 &  x986 &  x1124 & ~x300 & ~x696 & ~x729 & ~x774 & ~x775 & ~x813 & ~x885 & ~x964 & ~x1029 & ~x1108;
assign c3280 =  x13 &  x71 &  x205 &  x209 &  x257 &  x313 &  x316 &  x344 &  x356 &  x368 &  x434 &  x472 &  x545 &  x554 &  x653 &  x656 &  x731 &  x733 &  x739 &  x752 &  x754 &  x772 &  x778 &  x803 &  x805 &  x811 &  x1082 &  x1123 & ~x507 & ~x585;
assign c3282 =  x17 &  x26 &  x56 &  x71 &  x86 &  x137 &  x140 &  x175 &  x182 &  x236 &  x296 &  x304 &  x331 &  x356 &  x362 &  x409 &  x419 &  x434 &  x479 &  x481 &  x512 &  x515 &  x533 &  x545 &  x556 &  x595 &  x602 &  x653 &  x656 &  x725 &  x755 &  x773 &  x815 &  x818 &  x854 &  x859 &  x860 &  x901 &  x908 &  x911 &  x979 &  x980 &  x1018 &  x1028 &  x1037 &  x1057 &  x1096 & ~x84 & ~x123;
assign c3284 =  x92 &  x98 &  x110 &  x128 &  x245 &  x290 &  x481 &  x519 &  x566 &  x632 &  x638 &  x641 &  x659 &  x713 &  x722 &  x724 &  x734 &  x762 &  x782 &  x862 &  x875 &  x932 &  x974 &  x986 &  x989 &  x1031 &  x1040 &  x1043 &  x1082 &  x1097 &  x1100 &  x1130 & ~x429;
assign c3286 =  x47 &  x68 &  x107 &  x131 &  x170 &  x230 &  x314 &  x353 &  x356 &  x431 &  x460 &  x481 &  x503 &  x506 &  x512 &  x521 &  x532 &  x559 &  x632 &  x637 &  x647 &  x770 &  x782 &  x854 &  x926 &  x968 &  x976 &  x978 &  x998 &  x1013 &  x1015 &  x1018 &  x1031 &  x1046 &  x1049 &  x1052 &  x1056 &  x1096 &  x1097 &  x1127 & ~x315 & ~x391 & ~x393 & ~x430 & ~x508 & ~x547 & ~x651;
assign c3288 =  x1 &  x16 &  x50 &  x56 &  x100 &  x196 &  x203 &  x224 &  x295 &  x334 &  x373 &  x404 &  x434 &  x451 &  x481 &  x494 &  x526 &  x529 &  x556 &  x595 &  x607 &  x632 &  x946 &  x985 &  x1048 &  x1081;
assign c3290 =  x17 &  x92 &  x155 &  x218 &  x233 &  x260 &  x316 &  x394 &  x425 &  x433 &  x461 &  x472 &  x507 &  x509 &  x625 &  x667 &  x803 &  x806 &  x812 &  x862 &  x914 &  x1010 &  x1130 & ~x522 & ~x837;
assign c3292 =  x56 &  x104 &  x170 &  x188 &  x194 &  x200 &  x206 &  x284 &  x290 &  x494 &  x623 &  x630 &  x668 &  x670 &  x710 &  x728 &  x773 &  x776 &  x791 &  x842 &  x929 &  x1004 &  x1043 & ~x240 & ~x444 & ~x547 & ~x586 & ~x625;
assign c3294 =  x17 &  x26 &  x56 &  x68 &  x89 &  x92 &  x98 &  x113 &  x128 &  x137 &  x143 &  x157 &  x164 &  x173 &  x188 &  x199 &  x227 &  x238 &  x242 &  x263 &  x269 &  x272 &  x275 &  x277 &  x313 &  x314 &  x341 &  x356 &  x374 &  x377 &  x404 &  x407 &  x413 &  x416 &  x422 &  x431 &  x433 &  x446 &  x461 &  x473 &  x500 &  x533 &  x551 &  x590 &  x598 &  x616 &  x620 &  x623 &  x631 &  x637 &  x638 &  x641 &  x656 &  x674 &  x688 &  x691 &  x709 &  x721 &  x724 &  x727 &  x733 &  x746 &  x749 &  x754 &  x755 &  x760 &  x766 &  x770 &  x772 &  x785 &  x787 &  x799 &  x803 &  x805 &  x811 &  x827 &  x839 &  x844 &  x848 &  x854 &  x869 &  x881 &  x899 &  x902 &  x923 &  x977 &  x992 &  x1022 &  x1058 &  x1067 &  x1076 &  x1103 &  x1121 &  x1124 & ~x483 & ~x744;
assign c3296 =  x17 &  x38 &  x62 &  x68 &  x80 &  x92 &  x104 &  x164 &  x236 &  x257 &  x275 &  x323 &  x356 &  x368 &  x404 &  x455 &  x488 &  x494 &  x503 &  x506 &  x545 &  x548 &  x629 &  x632 &  x746 &  x752 &  x755 &  x821 &  x829 &  x848 &  x854 &  x862 &  x868 &  x869 &  x884 &  x901 &  x907 &  x983 &  x986 &  x1091 &  x1103 &  x1121 & ~x765 & ~x768 & ~x804 & ~x813 & ~x834 & ~x852 & ~x879 & ~x918 & ~x957;
assign c3298 =  x5 &  x17 &  x25 &  x44 &  x56 &  x62 &  x64 &  x98 &  x137 &  x233 &  x277 &  x314 &  x317 &  x329 &  x356 &  x433 &  x434 &  x479 &  x569 &  x602 &  x638 &  x659 &  x686 &  x713 &  x779 &  x812 &  x848 &  x908 &  x983 &  x1019 &  x1115 & ~x228 & ~x229 & ~x267 & ~x405 & ~x600 & ~x912;
assign c31 = ~x610;
assign c33 =  x232 &  x348 & ~x534 & ~x558 & ~x789 & ~x1119;
assign c35 =  x160 &  x834 &  x1069 &  x1097 & ~x591;
assign c37 =  x874 &  x991 & ~x826 & ~x888;
assign c39 =  x163 &  x350 &  x549 &  x740 & ~x363 & ~x441;
assign c311 =  x155 &  x379 &  x627 &  x835 &  x958 &  x980;
assign c313 = ~x1028;
assign c315 =  x2 &  x792 &  x1090 & ~x126 & ~x490;
assign c317 =  x109 & ~x516 & ~x636 & ~x787;
assign c319 = ~x288 & ~x915 & ~x943;
assign c321 =  x1060 &  x1089 & ~x214;
assign c323 =  x142 &  x240 &  x279 &  x827 &  x1025 & ~x288 & ~x501;
assign c325 =  x547 & ~x12 & ~x901;
assign c327 =  x1065 & ~x253;
assign c329 =  x600 &  x1051 & ~x267 & ~x861;
assign c331 =  x46 &  x697 & ~x550;
assign c333 =  x511 & ~x277 & ~x441 & ~x558 & ~x789;
assign c335 = ~x324 & ~x330 & ~x388 & ~x421;
assign c337 =  x835 &  x1029 &  x1102 & ~x882 & ~x960;
assign c339 =  x115 & ~x321 & ~x441 & ~x636 & ~x714;
assign c341 =  x121 &  x639 & ~x693 & ~x705;
assign c343 =  x639 & ~x420 & ~x693;
assign c345 =  x26 &  x796 & ~x288 & ~x474 & ~x570 & ~x822;
assign c347 =  x70 & ~x360 & ~x828 & ~x906;
assign c349 = ~x281 & ~x680;
assign c351 = ~x1109;
assign c353 =  x562 & ~x258 & ~x318 & ~x357 & ~x628;
assign c355 =  x987 & ~x801;
assign c357 =  x163 & ~x291 & ~x330 & ~x369 & ~x402 & ~x447 & ~x480 & ~x897;
assign c359 =  x1063 &  x1092 & ~x1099;
assign c361 =  x913 &  x1062 & ~x960 & ~x1011;
assign c363 =  x169 &  x395 & ~x198 & ~x204 & ~x441 & ~x636 & ~x714;
assign c365 = ~x285 & ~x402 & ~x438 & ~x636 & ~x714 & ~x1119;
assign c367 =  x273 &  x482 &  x994 &  x1006 &  x1039 & ~x186 & ~x207;
assign c369 =  x325 & ~x288 & ~x477 & ~x555 & ~x672 & ~x801;
assign c371 = ~x545;
assign c373 =  x682 & ~x46 & ~x438 & ~x900;
assign c375 =  x372 &  x382 &  x553 &  x755 &  x1035;
assign c377 =  x163 &  x697 & ~x943;
assign c379 = ~x394 & ~x471 & ~x477 & ~x636;
assign c381 = ~x511 & ~x718 & ~x786;
assign c383 =  x76 &  x188 &  x190 &  x229 &  x272 &  x356 &  x397 &  x437 &  x527 &  x560 &  x590 &  x761 &  x794 & ~x441 & ~x480;
assign c385 =  x160 &  x601 &  x949 &  x1019 & ~x24 & ~x148 & ~x258;
assign c387 =  x208 &  x622 & ~x474;
assign c389 =  x330 &  x1092 & ~x943;
assign c391 = ~x377;
assign c393 =  x81 &  x601 &  x679 &  x812 & ~x60 & ~x498;
assign c395 =  x109 &  x154 & ~x210 & ~x369 & ~x480;
assign c397 =  x852 &  x969 &  x1047 &  x1092 &  x1120;
assign c399 = ~x35;
assign c3101 =  x832 & ~x90 & ~x490;
assign c3103 =  x163 &  x422 &  x596 &  x767 &  x1118 & ~x207 & ~x402 & ~x606 & ~x936;
assign c3105 = ~x54 & ~x267 & ~x543 & ~x550;
assign c3107 =  x725 &  x961 &  x1026 & ~x252 & ~x291 & ~x408 & ~x621;
assign c3109 = ~x362;
assign c3111 =  x241 & ~x394 & ~x720;
assign c3113 =  x70 &  x76 &  x730 & ~x210 & ~x306;
assign c3115 =  x1065 &  x1072 & ~x357;
assign c3117 =  x949 & ~x138 & ~x258 & ~x292;
assign c3119 =  x233 &  x483 &  x522 &  x553 &  x562 &  x601 &  x619 &  x630 &  x670;
assign c3121 =  x163 &  x190 &  x229 &  x301 &  x436 &  x991 &  x1087 &  x1126 & ~x441;
assign c3123 =  x7 & ~x591;
assign c3125 =  x510 & ~x321 & ~x481;
assign c3127 =  x76 &  x248 &  x305 &  x374 &  x719 &  x809 &  x986 &  x1003 &  x1006 & ~x441 & ~x480;
assign c3129 =  x437 &  x995 & ~x177 & ~x550 & ~x1101;
assign c3131 =  x19 & ~x9 & ~x901;
assign c3133 =  x29 &  x83 &  x163 &  x221 &  x379 &  x397 &  x719 &  x875 &  x998 &  x1091 & ~x159 & ~x480;
assign c3135 =  x460 &  x909 &  x1069 & ~x864;
assign c3137 = ~x438 & ~x472 & ~x675;
assign c3139 =  x28 &  x835 & ~x447 & ~x484;
assign c3141 =  x241 &  x358 &  x407 & ~x433 & ~x636 & ~x714;
assign c3143 =  x1105 & ~x12 & ~x70 & ~x822;
assign c3145 = ~x199 & ~x441 & ~x718;
assign c3147 =  x640 &  x1008 &  x1035 & ~x75;
assign c3149 = ~x276 & ~x756 & ~x943;
assign c3151 =  x164 &  x562 &  x631 &  x641 &  x697 & ~x357 & ~x628;
assign c3153 = ~x199 & ~x481;
assign c3155 =  x697 & ~x345 & ~x589;
assign c3157 =  x2 &  x263 &  x311 &  x575 &  x608 &  x719 &  x824 &  x842 &  x1033 &  x1073 &  x1103 &  x1105 & ~x207 & ~x285 & ~x324 & ~x357 & ~x858;
assign c3159 =  x163 &  x197 &  x936 &  x1069;
assign c3161 = ~x199 & ~x523;
assign c3163 =  x1075 & ~x718 & ~x864;
assign c3165 = ~x670 & ~x901 & ~x979;
assign c3167 = ~x857;
assign c3169 = ~x12 & ~x51 & ~x168 & ~x705 & ~x901 & ~x940;
assign c3171 =  x601 &  x991 & ~x436;
assign c3173 =  x640 & ~x475;
assign c3175 =  x20 &  x23 &  x62 &  x155 &  x160 &  x163 &  x170 &  x173 &  x179 &  x221 &  x241 &  x251 &  x368 &  x452 &  x461 &  x701 &  x719 &  x737 &  x743 &  x757 &  x779 &  x802 &  x812 &  x830 &  x835 &  x874 &  x881 &  x890 &  x935 &  x991 &  x998 &  x1055 &  x1069 &  x1103;
assign c3177 =  x824 &  x988 & ~x48 & ~x87 & ~x285 & ~x330 & ~x801;
assign c3179 = ~x12 & ~x207 & ~x265 & ~x304;
assign c3181 = ~x160;
assign c3183 =  x127 &  x436 &  x631 & ~x636 & ~x798;
assign c3185 =  x156 & ~x13 & ~x327;
assign c3187 =  x160 &  x834 &  x923 &  x991 &  x1069 &  x1108 & ~x591;
assign c3189 =  x19 &  x279 &  x397;
assign c3191 =  x31 & ~x270 & ~x1021;
assign c3193 =  x76 &  x190 &  x991 & ~x288 & ~x771;
assign c3195 =  x312 &  x915 & ~x207;
assign c3197 =  x167 &  x200 &  x416 &  x581 &  x647 &  x701 & ~x354 & ~x399 & ~x636 & ~x714 & ~x846 & ~x864 & ~x972;
assign c3199 =  x17 &  x84 &  x113 &  x269 &  x353 &  x389 &  x476 &  x545 &  x641 &  x689 &  x749 &  x758 &  x835 &  x857 &  x874 &  x913 &  x997;
assign c3201 =  x6 & ~x801 & ~x1123;
assign c3203 =  x241 &  x397 &  x936 &  x997 & ~x753;
assign c3205 = ~x90 & ~x703 & ~x801;
assign c3207 = ~x206;
assign c3209 =  x601 &  x1117 & ~x589 & ~x628;
assign c3211 =  x744 & ~x394 & ~x519;
assign c3213 =  x862 &  x922 & ~x126 & ~x403;
assign c3215 =  x798 & ~x52;
assign c3217 = ~x731;
assign c3219 = ~x242;
assign c3221 =  x89 &  x131 &  x629 &  x827 &  x869 &  x1049 & ~x87 & ~x207 & ~x213 & ~x285 & ~x369 & ~x402 & ~x663 & ~x819;
assign c3223 =  x382 &  x1053;
assign c3225 =  x190 &  x1126 & ~x288 & ~x516 & ~x693;
assign c3227 =  x156 & ~x138 & ~x187 & ~x213;
assign c3229 =  x127 &  x248 &  x290 &  x301 &  x461 &  x473 &  x650 &  x767 &  x926 & ~x555 & ~x753 & ~x772;
assign c3231 = ~x670 & ~x901;
assign c3233 =  x163 & ~x285 & ~x484;
assign c3235 =  x387 &  x1128;
assign c3237 =  x14 &  x98 &  x134 &  x163 &  x863 &  x944 &  x1034 & ~x168 & ~x207 & ~x246 & ~x285 & ~x441 & ~x480 & ~x978;
assign c3239 =  x991 & ~x771 & ~x789 & ~x805;
assign c3241 =  x160 &  x561 &  x600 & ~x414;
assign c3243 =  x31 &  x1128 & ~x246 & ~x435;
assign c3245 =  x56 &  x85 &  x269 &  x272 &  x350 &  x356 &  x383 &  x410 &  x449 &  x470 &  x730 &  x770 &  x776 &  x851 &  x905 &  x986 &  x1103 &  x1109 & ~x396 & ~x450 & ~x451 & ~x489;
assign c3247 = ~x51 & ~x171 & ~x901;
assign c3249 =  x156 &  x949 & ~x99 & ~x226;
assign c3251 =  x121 &  x819 &  x835 &  x1030 & ~x1038;
assign c3253 =  x700 & ~x556 & ~x801;
assign c3255 =  x202 & ~x693 & ~x1123;
assign c3257 =  x76 &  x190 &  x466 &  x1069 & ~x210 & ~x888;
assign c3259 =  x76 &  x424 &  x657 & ~x960;
assign c3261 =  x169 &  x356 &  x467 &  x780 &  x1053 & ~x234;
assign c3263 = ~x748 & ~x979;
assign c3265 =  x418 & ~x526 & ~x565;
assign c3267 =  x5 &  x575 &  x1079 &  x1097 &  x1117 & ~x474 & ~x525 & ~x750 & ~x867 & ~x1119;
assign c3269 = ~x20;
assign c3271 =  x76 &  x853 &  x949 &  x1104 &  x1105 & ~x138;
assign c3273 =  x466 &  x544 &  x580 & ~x754;
assign c3275 = ~x609 & ~x784;
assign c3277 =  x349 &  x466 & ~x595 & ~x750;
assign c3279 =  x34 &  x163 &  x397 & ~x480 & ~x753;
assign c3281 =  x19 &  x70 &  x163 &  x190 &  x505 & ~x450;
assign c3283 =  x31 &  x154 &  x908 &  x965 & ~x324 & ~x363 & ~x441 & ~x714;
assign c3285 =  x352 &  x1105 & ~x15 & ~x207 & ~x591 & ~x822;
assign c3287 =  x85 & ~x511 & ~x714 & ~x753;
assign c3289 =  x240 &  x336 &  x375 &  x697;
assign c3291 =  x123 &  x279 &  x727 & ~x606;
assign c3293 = ~x204 & ~x276 & ~x441 & ~x501 & ~x750 & ~x789;
assign c3295 =  x431 &  x835 &  x1090 &  x1105 & ~x210 & ~x474;
assign c3297 =  x471 &  x505 &  x763 &  x796;
assign c3299 =  x31 &  x163 & ~x285 & ~x801 & ~x1119;
assign c40 =  x3 &  x4 &  x40 &  x42 &  x43 &  x44 &  x47 &  x79 &  x80 &  x81 &  x82 &  x118 &  x120 &  x121 &  x143 &  x160 &  x161 &  x164 &  x170 &  x199 &  x200 &  x230 &  x233 &  x238 &  x260 &  x266 &  x284 &  x347 &  x350 &  x353 &  x371 &  x404 &  x449 &  x452 &  x470 &  x497 &  x503 &  x512 &  x542 &  x545 &  x548 &  x557 &  x566 &  x575 &  x581 &  x584 &  x587 &  x601 &  x617 &  x620 &  x626 &  x632 &  x640 &  x644 &  x671 &  x679 &  x689 &  x701 &  x704 &  x707 &  x718 &  x725 &  x731 &  x740 &  x754 &  x757 &  x806 &  x812 &  x908 &  x926 &  x973 &  x974 &  x1013 &  x1022 &  x1049 &  x1064 &  x1082 &  x1112 & ~x387 & ~x426;
assign c42 =  x469 &  x637 &  x679 &  x718 &  x796 &  x835 & ~x435 & ~x462 & ~x489 & ~x528 & ~x606;
assign c44 =  x68 &  x80 &  x89 &  x116 &  x119 &  x143 &  x152 &  x170 &  x179 &  x188 &  x206 &  x224 &  x245 &  x272 &  x278 &  x290 &  x293 &  x311 &  x326 &  x338 &  x350 &  x371 &  x401 &  x419 &  x422 &  x425 &  x428 &  x443 &  x458 &  x461 &  x464 &  x467 &  x476 &  x511 &  x512 &  x527 &  x530 &  x545 &  x547 &  x560 &  x566 &  x599 &  x611 &  x625 &  x659 &  x686 &  x698 &  x704 &  x707 &  x719 &  x734 &  x743 &  x752 &  x779 &  x905 &  x908 &  x911 &  x917 &  x923 &  x935 &  x980 &  x983 &  x998 &  x1028 &  x1034 &  x1040 &  x1049 &  x1055 &  x1058 &  x1067 &  x1070 &  x1088 &  x1106 &  x1115 & ~x477 & ~x576 & ~x615 & ~x654 & ~x669 & ~x670 & ~x708 & ~x732 & ~x771 & ~x810 & ~x822;
assign c46 =  x20 &  x64 &  x299 &  x329 &  x337 &  x505 &  x987 &  x1040 &  x1088 & ~x321 & ~x903;
assign c48 =  x17 &  x43 &  x82 &  x109 &  x121 &  x128 &  x143 &  x160 &  x176 &  x199 &  x209 &  x269 &  x299 &  x335 &  x371 &  x398 &  x407 &  x446 &  x461 &  x497 &  x539 &  x557 &  x560 &  x562 &  x584 &  x590 &  x601 &  x638 &  x679 &  x695 &  x718 &  x749 &  x796 &  x800 &  x835 &  x851 &  x874 &  x887 &  x941 &  x947 &  x983 &  x1043 &  x1084 &  x1091 &  x1103 &  x1124 & ~x630 & ~x822;
assign c410 =  x32 &  x74 &  x86 &  x107 &  x182 &  x227 &  x290 &  x362 &  x368 &  x395 &  x404 &  x428 &  x482 &  x485 &  x656 &  x677 &  x679 &  x680 &  x718 &  x740 &  x752 &  x757 &  x835 &  x845 &  x860 &  x863 &  x872 &  x908 &  x911 &  x923 &  x977 &  x1001 &  x1013 &  x1070 &  x1085 & ~x15 & ~x54 & ~x165 & ~x279 & ~x501 & ~x540 & ~x744 & ~x930;
assign c412 =  x158 &  x182 &  x220 &  x242 &  x347 &  x539 &  x647 &  x659 &  x680 &  x683 &  x725 &  x757 &  x796 &  x835 &  x874 &  x910 &  x913 &  x952 &  x991 &  x1010 &  x1030 &  x1058 &  x1069 &  x1108 &  x1114 &  x1120 & ~x849;
assign c414 =  x237 &  x245 &  x272 &  x276 &  x316 &  x329 &  x368 &  x506 &  x512 &  x517 &  x595 &  x752 &  x796 &  x797 &  x835 &  x953 &  x1067 & ~x397 & ~x861 & ~x1017;
assign c416 =  x26 &  x65 &  x68 &  x77 &  x80 &  x104 &  x113 &  x116 &  x122 &  x146 &  x191 &  x230 &  x233 &  x245 &  x251 &  x263 &  x269 &  x272 &  x299 &  x344 &  x380 &  x386 &  x395 &  x398 &  x434 &  x467 &  x500 &  x512 &  x515 &  x518 &  x560 &  x572 &  x575 &  x584 &  x593 &  x596 &  x626 &  x635 &  x656 &  x710 &  x740 &  x746 &  x785 &  x788 &  x791 &  x809 &  x812 &  x836 &  x854 &  x870 &  x887 &  x950 &  x959 &  x965 &  x983 &  x989 &  x1019 &  x1022 &  x1030 &  x1034 &  x1046 &  x1049 &  x1064 &  x1067 &  x1069 &  x1082 &  x1103 &  x1108 &  x1112 &  x1115 &  x1121 &  x1130 & ~x156 & ~x390 & ~x786;
assign c418 =  x59 &  x119 &  x124 &  x142 &  x202 &  x206 &  x215 &  x241 &  x332 &  x341 &  x359 &  x371 &  x419 &  x471 &  x510 &  x530 &  x554 &  x569 &  x599 &  x689 &  x827 &  x830 &  x851 &  x866 &  x998 &  x1004 &  x1010 &  x1022 &  x1052 &  x1079 &  x1109 & ~x117 & ~x345 & ~x384 & ~x747;
assign c420 =  x73 &  x74 &  x79 &  x118 &  x119 &  x295 &  x302 &  x334 &  x350 &  x373 &  x386 &  x409 &  x419 &  x428 &  x449 &  x458 &  x539 &  x710 &  x743 &  x770 &  x794 &  x905 &  x914 &  x938 &  x997 &  x998 &  x1061 &  x1085 & ~x129 & ~x777 & ~x816 & ~x855 & ~x894 & ~x933 & ~x1077 & ~x1116 & ~x1122;
assign c422 =  x8 &  x143 &  x319 &  x323 &  x359 &  x394 &  x433 &  x461 &  x508 &  x860 &  x983 & ~x426 & ~x438 & ~x439 & ~x738 & ~x777 & ~x1017;
assign c424 =  x5 &  x26 &  x92 &  x146 &  x241 &  x248 &  x326 &  x404 &  x431 &  x440 &  x449 &  x469 &  x472 &  x527 &  x598 &  x602 &  x611 &  x636 &  x637 &  x640 &  x653 &  x675 &  x679 &  x698 &  x718 &  x725 &  x728 &  x755 &  x827 &  x836 &  x845 &  x851 &  x914 &  x950 &  x1022 & ~x438 & ~x552;
assign c426 =  x120 &  x121 &  x140 &  x159 &  x160 &  x198 &  x199 &  x308 &  x335 &  x368 &  x389 &  x442 &  x695 &  x803 &  x821 &  x935 &  x1028 &  x1121 & ~x279 & ~x318 & ~x319 & ~x358 & ~x435 & ~x705;
assign c428 =  x701 &  x741 &  x820 & ~x786 & ~x855 & ~x864 & ~x1017 & ~x1056 & ~x1110;
assign c430 =  x14 &  x188 &  x191 &  x290 &  x329 &  x335 &  x377 &  x461 &  x536 &  x569 &  x581 &  x638 &  x664 &  x713 &  x742 &  x757 &  x796 &  x835 &  x871 &  x874 &  x907 &  x992 &  x1103 & ~x709 & ~x748 & ~x786 & ~x787 & ~x825;
assign c432 =  x206 &  x705 &  x862 &  x984 &  x985 & ~x468 & ~x865 & ~x903 & ~x904 & ~x943 & ~x982;
assign c434 =  x2 &  x35 &  x89 &  x224 &  x272 &  x326 &  x338 &  x371 &  x431 &  x434 &  x488 &  x491 &  x640 &  x725 &  x770 &  x773 &  x788 &  x818 &  x998 &  x1019 &  x1049 & ~x51 & ~x90 & ~x96 & ~x135 & ~x498 & ~x606 & ~x864 & ~x1059;
assign c436 =  x65 &  x215 &  x257 &  x314 &  x389 &  x467 &  x515 &  x524 &  x536 &  x563 &  x683 &  x755 &  x806 &  x809 &  x833 &  x845 &  x851 &  x917 &  x998 &  x1001 &  x1043 & ~x234 & ~x579 & ~x826 & ~x840 & ~x879 & ~x880 & ~x888 & ~x903 & ~x918 & ~x927 & ~x942 & ~x981;
assign c438 =  x98 &  x140 &  x209 &  x212 &  x230 &  x241 &  x254 &  x259 &  x280 &  x308 &  x329 &  x389 &  x395 &  x398 &  x401 &  x422 &  x449 &  x452 &  x471 &  x494 &  x497 &  x510 &  x599 &  x632 &  x677 &  x689 &  x722 &  x749 &  x761 &  x764 &  x881 &  x902 &  x920 &  x952 &  x991 &  x1031 &  x1100 & ~x345 & ~x384 & ~x423;
assign c440 =  x4 &  x6 &  x43 &  x81 &  x101 &  x118 &  x120 &  x159 &  x199 &  x314 &  x601 &  x836 &  x860 &  x1055 & ~x300;
assign c442 =  x8 &  x26 &  x38 &  x47 &  x77 &  x98 &  x113 &  x128 &  x134 &  x137 &  x140 &  x167 &  x170 &  x203 &  x224 &  x226 &  x227 &  x245 &  x254 &  x260 &  x263 &  x265 &  x269 &  x275 &  x278 &  x290 &  x304 &  x305 &  x317 &  x326 &  x341 &  x343 &  x347 &  x358 &  x359 &  x368 &  x380 &  x386 &  x389 &  x398 &  x404 &  x413 &  x416 &  x425 &  x431 &  x433 &  x446 &  x449 &  x471 &  x472 &  x476 &  x509 &  x524 &  x533 &  x539 &  x547 &  x550 &  x551 &  x575 &  x581 &  x586 &  x593 &  x629 &  x632 &  x650 &  x665 &  x674 &  x677 &  x692 &  x707 &  x716 &  x722 &  x725 &  x749 &  x755 &  x773 &  x785 &  x788 &  x800 &  x809 &  x833 &  x836 &  x842 &  x848 &  x857 &  x863 &  x869 &  x878 &  x881 &  x902 &  x917 &  x923 &  x926 &  x932 &  x935 &  x947 &  x953 &  x986 &  x992 &  x1001 &  x1007 &  x1022 &  x1034 &  x1040 &  x1046 &  x1052 &  x1061 &  x1070 &  x1076 &  x1079 &  x1082 &  x1100 &  x1109 &  x1115 & ~x444 & ~x670 & ~x978;
assign c444 =  x89 &  x142 &  x155 &  x175 &  x202 &  x221 &  x280 &  x356 &  x432 &  x471 &  x510 &  x602 &  x674 &  x839 &  x842 &  x872 &  x920 &  x926 &  x1046 &  x1085 & ~x438 & ~x516 & ~x591;
assign c446 =  x59 &  x86 &  x266 &  x374 &  x506 &  x588 &  x617 &  x767 &  x829 & ~x543 & ~x709 & ~x825 & ~x864;
assign c448 =  x14 &  x65 &  x83 &  x89 &  x95 &  x131 &  x140 &  x143 &  x170 &  x179 &  x209 &  x221 &  x242 &  x248 &  x266 &  x269 &  x278 &  x284 &  x296 &  x329 &  x332 &  x374 &  x377 &  x380 &  x404 &  x413 &  x431 &  x440 &  x461 &  x467 &  x470 &  x473 &  x476 &  x482 &  x494 &  x497 &  x509 &  x518 &  x539 &  x563 &  x569 &  x599 &  x611 &  x614 &  x686 &  x716 &  x728 &  x740 &  x782 &  x794 &  x809 &  x824 &  x833 &  x875 &  x896 &  x899 &  x911 &  x914 &  x941 &  x968 &  x974 &  x980 &  x983 &  x1034 &  x1043 &  x1052 &  x1064 &  x1067 &  x1097 &  x1121 & ~x447 & ~x606 & ~x618 & ~x838 & ~x877;
assign c450 =  x176 &  x203 &  x242 &  x299 &  x350 &  x458 &  x521 &  x578 &  x686 &  x773 &  x788 &  x820 &  x897 &  x1064 &  x1091 &  x1130 & ~x321 & ~x618 & ~x696 & ~x735 & ~x903 & ~x942 & ~x966 & ~x981 & ~x982;
assign c452 =  x1 &  x4 &  x20 &  x40 &  x43 &  x68 &  x79 &  x82 &  x104 &  x149 &  x218 &  x221 &  x257 &  x308 &  x314 &  x317 &  x320 &  x335 &  x338 &  x347 &  x353 &  x359 &  x383 &  x467 &  x515 &  x533 &  x545 &  x575 &  x578 &  x601 &  x617 &  x620 &  x635 &  x641 &  x647 &  x653 &  x674 &  x689 &  x701 &  x707 &  x710 &  x719 &  x722 &  x725 &  x737 &  x740 &  x755 &  x770 &  x809 &  x818 &  x827 &  x923 &  x947 &  x980 &  x992 &  x998 &  x1049 &  x1055 &  x1088 &  x1112 &  x1121 & ~x30 & ~x69 & ~x90 & ~x153 & ~x192 & ~x309 & ~x348 & ~x384 & ~x582 & ~x621;
assign c454 =  x365 &  x446 &  x503 &  x545 &  x668 &  x926 &  x1118 & ~x255 & ~x321 & ~x579 & ~x711 & ~x801 & ~x825 & ~x840 & ~x864 & ~x879 & ~x903 & ~x918 & ~x927 & ~x957 & ~x963 & ~x966 & ~x1005;
assign c456 =  x5 &  x11 &  x56 &  x68 &  x71 &  x77 &  x80 &  x89 &  x98 &  x122 &  x140 &  x143 &  x155 &  x161 &  x176 &  x197 &  x203 &  x218 &  x257 &  x260 &  x269 &  x287 &  x302 &  x308 &  x359 &  x374 &  x398 &  x425 &  x437 &  x440 &  x446 &  x464 &  x491 &  x503 &  x506 &  x515 &  x548 &  x550 &  x557 &  x572 &  x578 &  x581 &  x588 &  x599 &  x614 &  x617 &  x647 &  x659 &  x665 &  x692 &  x698 &  x704 &  x716 &  x719 &  x758 &  x782 &  x791 &  x793 &  x800 &  x806 &  x818 &  x827 &  x829 &  x833 &  x836 &  x839 &  x845 &  x869 &  x872 &  x881 &  x947 &  x959 &  x1016 &  x1028 &  x1052 &  x1058 &  x1070 &  x1076 &  x1079 &  x1100 &  x1124 &  x1130 & ~x351 & ~x669 & ~x684 & ~x709 & ~x723 & ~x762 & ~x786 & ~x801;
assign c458 =  x198 &  x218 &  x237 &  x350 &  x362 &  x476 &  x517 &  x551 &  x578 &  x641 &  x815 &  x893 &  x920 & ~x358 & ~x397 & ~x436 & ~x474 & ~x475;
assign c460 =  x311 &  x530 &  x702 &  x824 &  x1034 & ~x570 & ~x594 & ~x621 & ~x771 & ~x786 & ~x810 & ~x849 & ~x855 & ~x927;
assign c462 =  x4 &  x22 &  x28 &  x61 &  x85 &  x106 &  x137 &  x143 &  x161 &  x221 &  x229 &  x302 &  x376 &  x380 &  x383 &  x415 &  x500 &  x551 &  x566 &  x581 &  x608 &  x682 &  x704 &  x719 &  x728 &  x866 &  x878 &  x899 &  x929 &  x932 &  x956 &  x962 &  x1046 &  x1079 &  x1108;
assign c464 =  x112 &  x223 &  x469 &  x527 &  x679 &  x718 &  x796 &  x835 &  x913 &  x952 &  x1030 &  x1087 & ~x348 & ~x387 & ~x465 & ~x504 & ~x621;
assign c466 =  x23 &  x32 &  x35 &  x65 &  x86 &  x137 &  x140 &  x179 &  x248 &  x251 &  x260 &  x265 &  x287 &  x320 &  x347 &  x383 &  x386 &  x433 &  x440 &  x458 &  x476 &  x510 &  x518 &  x524 &  x542 &  x548 &  x551 &  x563 &  x572 &  x586 &  x596 &  x620 &  x632 &  x662 &  x671 &  x680 &  x731 &  x779 &  x782 &  x803 &  x830 &  x833 &  x842 &  x851 &  x929 &  x956 &  x980 &  x986 &  x1010 &  x1025 &  x1043 &  x1055 &  x1067 &  x1118 & ~x606 & ~x786 & ~x1017 & ~x1056;
assign c468 =  x41 &  x80 &  x197 &  x266 &  x275 &  x278 &  x281 &  x311 &  x316 &  x320 &  x341 &  x401 &  x437 &  x581 &  x815 &  x872 &  x914 &  x1049 & ~x321 & ~x411 & ~x450 & ~x474 & ~x489 & ~x513 & ~x514 & ~x528 & ~x591 & ~x939 & ~x1017 & ~x1056;
assign c470 =  x31 &  x37 &  x70 &  x76 &  x103 &  x109 &  x115 &  x131 &  x142 &  x154 &  x181 &  x193 &  x202 &  x212 &  x226 &  x241 &  x280 &  x284 &  x319 &  x443 &  x461 &  x472 &  x722 &  x731 &  x791 &  x833 &  x887 &  x896 &  x920 &  x935 &  x956 &  x1016 &  x1112 & ~x438 & ~x477;
assign c472 =  x20 &  x26 &  x35 &  x41 &  x56 &  x83 &  x86 &  x101 &  x107 &  x113 &  x119 &  x120 &  x121 &  x122 &  x128 &  x149 &  x160 &  x176 &  x179 &  x182 &  x185 &  x198 &  x199 &  x203 &  x209 &  x218 &  x230 &  x236 &  x239 &  x254 &  x257 &  x263 &  x266 &  x269 &  x277 &  x287 &  x290 &  x302 &  x308 &  x314 &  x320 &  x356 &  x359 &  x368 &  x371 &  x383 &  x392 &  x398 &  x404 &  x413 &  x422 &  x449 &  x455 &  x476 &  x479 &  x482 &  x494 &  x509 &  x515 &  x518 &  x548 &  x557 &  x569 &  x572 &  x575 &  x584 &  x599 &  x626 &  x632 &  x638 &  x644 &  x650 &  x653 &  x671 &  x683 &  x686 &  x698 &  x701 &  x704 &  x713 &  x716 &  x719 &  x728 &  x731 &  x734 &  x740 &  x758 &  x761 &  x764 &  x773 &  x779 &  x797 &  x803 &  x809 &  x815 &  x818 &  x824 &  x833 &  x875 &  x878 &  x884 &  x893 &  x908 &  x914 &  x917 &  x920 &  x926 &  x929 &  x935 &  x938 &  x956 &  x962 &  x965 &  x1004 &  x1019 &  x1037 &  x1046 &  x1052 &  x1055 &  x1064 &  x1079 &  x1082 &  x1088 &  x1097 &  x1106 &  x1130 & ~x192 & ~x204 & ~x280 & ~x319 & ~x396;
assign c474 =  x20 &  x65 &  x113 &  x120 &  x122 &  x159 &  x160 &  x196 &  x224 &  x227 &  x242 &  x281 &  x347 &  x404 &  x512 &  x563 &  x596 &  x599 &  x620 &  x689 &  x743 &  x749 &  x800 &  x953 &  x1019 &  x1043 &  x1082 &  x1127 &  x1130 & ~x166 & ~x318 & ~x357 & ~x358;
assign c476 =  x28 &  x250 &  x328 &  x538 &  x881 &  x952 &  x990 &  x991 &  x1030 &  x1108 & ~x852;
assign c478 =  x4 &  x40 &  x79 &  x118 &  x233 &  x235 &  x308 &  x335 &  x445 &  x476 &  x538 &  x562 &  x577 &  x601 &  x616 &  x640 &  x679 &  x682 &  x718 &  x721 &  x796 &  x935 & ~x72;
assign c480 =  x20 &  x164 &  x254 &  x263 &  x298 &  x389 &  x401 &  x407 &  x476 &  x557 &  x584 &  x617 &  x632 &  x647 &  x692 &  x704 &  x740 &  x742 &  x860 &  x887 &  x896 &  x968 &  x986 &  x989 &  x1007 &  x1016 &  x1037 &  x1112 & ~x633 & ~x654 & ~x669 & ~x732 & ~x747 & ~x771 & ~x786 & ~x810 & ~x849 & ~x855 & ~x888 & ~x927 & ~x1017 & ~x1056;
assign c482 =  x11 &  x467 &  x470 &  x475 &  x487 &  x499 &  x509 &  x514 &  x526 &  x538 &  x542 &  x565 &  x593 &  x632 &  x695 &  x901 &  x992 & ~x751 & ~x807 & ~x846;
assign c484 =  x1 &  x16 &  x40 &  x118 &  x119 &  x143 &  x155 &  x176 &  x203 &  x250 &  x367 &  x368 &  x406 &  x440 &  x458 &  x538 &  x577 &  x578 &  x640 &  x734 &  x785 &  x926 &  x1058 &  x1068 &  x1069 &  x1092 &  x1103 &  x1107 &  x1108 & ~x1020;
assign c486 =  x42 &  x43 &  x79 &  x81 &  x82 &  x83 &  x120 &  x121 &  x159 &  x160 &  x195 &  x237 &  x277 &  x467 &  x491 &  x575 &  x578 &  x601 &  x640 &  x679 &  x863 &  x884 &  x956 &  x995 &  x1055 &  x1118 & ~x357;
assign c488 =  x28 &  x29 &  x35 &  x41 &  x44 &  x56 &  x62 &  x73 &  x112 &  x128 &  x134 &  x143 &  x152 &  x184 &  x188 &  x224 &  x230 &  x260 &  x275 &  x284 &  x287 &  x293 &  x317 &  x368 &  x371 &  x380 &  x385 &  x386 &  x395 &  x401 &  x404 &  x415 &  x431 &  x443 &  x446 &  x467 &  x497 &  x524 &  x529 &  x542 &  x548 &  x557 &  x575 &  x581 &  x587 &  x602 &  x613 &  x614 &  x620 &  x641 &  x662 &  x668 &  x680 &  x683 &  x707 &  x716 &  x740 &  x743 &  x749 &  x752 &  x764 &  x791 &  x797 &  x806 &  x827 &  x833 &  x851 &  x860 &  x878 &  x898 &  x899 &  x911 &  x926 &  x932 &  x935 &  x944 &  x976 &  x991 &  x995 &  x1031 &  x1054 &  x1069 &  x1093 &  x1108 &  x1124 &  x1130 & ~x927;
assign c490 =  x5 &  x257 &  x266 &  x284 &  x376 &  x475 &  x521 &  x820 &  x893 &  x965 &  x985 & ~x786 & ~x855 & ~x894 & ~x933 & ~x1017 & ~x1077;
assign c492 =  x23 &  x71 &  x281 &  x518 &  x910 &  x948 & ~x787 & ~x801 & ~x825 & ~x826 & ~x840 & ~x864 & ~x903;
assign c494 =  x20 &  x29 &  x50 &  x70 &  x109 &  x143 &  x202 &  x226 &  x241 &  x272 &  x280 &  x320 &  x349 &  x358 &  x364 &  x377 &  x410 &  x431 &  x461 &  x497 &  x589 &  x602 &  x611 &  x627 &  x722 &  x742 &  x782 &  x920 &  x1058 &  x1100 & ~x468 & ~x594;
assign c496 =  x199 &  x237 &  x254 &  x276 &  x338 &  x517 &  x679 &  x718 &  x797 & ~x435 & ~x436;
assign c498 =  x71 &  x116 &  x128 &  x143 &  x692 &  x758 &  x773 &  x812 &  x827 &  x830 &  x871 &  x935 &  x995 &  x1073 &  x1088 & ~x24 & ~x90 & ~x309 & ~x348 & ~x420 & ~x589 & ~x628 & ~x667 & ~x1017 & ~x1095;
assign c4100 =  x82 &  x121 &  x160 &  x198 &  x257 &  x281 &  x313 &  x338 &  x368 &  x452 &  x515 &  x523 &  x536 &  x601 &  x640 &  x653 &  x679 &  x718 &  x749 &  x776 &  x796 &  x835 &  x836 &  x910 &  x917 &  x929 &  x932 &  x950 &  x955 &  x956 &  x986 &  x1007 &  x1039 &  x1055 &  x1106 & ~x501;
assign c4102 =  x8 &  x50 &  x59 &  x119 &  x176 &  x197 &  x200 &  x257 &  x368 &  x371 &  x431 &  x527 &  x545 &  x587 &  x593 &  x602 &  x611 &  x785 &  x812 &  x875 &  x932 &  x989 &  x1013 &  x1025 &  x1058 &  x1097 &  x1100 & ~x30 & ~x225 & ~x231 & ~x270 & ~x309 & ~x348 & ~x420 & ~x543 & ~x582 & ~x696 & ~x738 & ~x816 & ~x855 & ~x933 & ~x972 & ~x999 & ~x1077 & ~x1116;
assign c4104 =  x4 &  x118 &  x284 &  x599 &  x836 & ~x93 & ~x336 & ~x345 & ~x411 & ~x450 & ~x729;
assign c4106 =  x20 &  x278 &  x308 &  x355 &  x508 &  x545 &  x587 &  x665 &  x755 &  x796 &  x835 &  x874 &  x875 &  x913 &  x952 &  x991 &  x1103 &  x1130 & ~x360 & ~x399 & ~x534 & ~x573 & ~x699;
assign c4108 =  x29 &  x329 &  x358 &  x383 &  x434 &  x437 &  x485 &  x509 &  x596 &  x626 &  x635 &  x703 &  x716 &  x791 &  x793 &  x863 &  x875 &  x907 & ~x609 & ~x654 & ~x693 & ~x786 & ~x810 & ~x849 & ~x927;
assign c4110 =  x3 &  x4 &  x79 &  x82 &  x601 &  x640 &  x679 &  x718 &  x728 &  x835 &  x959 &  x973 & ~x33 & ~x132;
assign c4112 = ~x132 & ~x255 & ~x567 & ~x645 & ~x684 & ~x729 & ~x769 & ~x774 & ~x807 & ~x864 & ~x903 & ~x1086;
assign c4114 =  x20 &  x308 &  x458 &  x461 &  x557 &  x590 &  x611 &  x725 &  x923 & ~x270 & ~x321 & ~x322 & ~x435 & ~x474 & ~x475;
assign c4116 =  x1 &  x8 &  x22 &  x184 &  x212 &  x295 &  x658 &  x871 &  x1030 &  x1069 &  x1081 &  x1087 &  x1108 &  x1114 & ~x1056;
assign c4118 =  x149 &  x347 &  x471 &  x510 &  x796 &  x835 &  x952 &  x965 & ~x423 & ~x462 & ~x501 & ~x747;
assign c4120 =  x28 &  x40 &  x79 &  x757 &  x835 & ~x186 & ~x264 & ~x291 & ~x486 & ~x504 & ~x1017 & ~x1056;
assign c4122 =  x35 &  x95 &  x170 &  x206 &  x260 &  x290 &  x308 &  x326 &  x335 &  x350 &  x392 &  x413 &  x434 &  x467 &  x476 &  x497 &  x518 &  x548 &  x575 &  x590 &  x656 &  x671 &  x686 &  x689 &  x704 &  x707 &  x740 &  x742 &  x794 &  x818 &  x845 &  x869 &  x875 &  x917 &  x920 &  x989 &  x991 &  x1030 &  x1031 &  x1069 &  x1106 &  x1124 & ~x237 & ~x516 & ~x810 & ~x816 & ~x849 & ~x855 & ~x903 & ~x942 & ~x972 & ~x1050 & ~x1077 & ~x1089 & ~x1110;
assign c4124 =  x2 &  x16 &  x55 &  x73 &  x80 &  x94 &  x133 &  x151 &  x173 &  x211 &  x215 &  x250 &  x287 &  x290 &  x314 &  x371 &  x458 &  x530 &  x626 &  x950 &  x952 &  x991 &  x1049 &  x1103 & ~x693 & ~x774 & ~x777 & ~x1083;
assign c4126 =  x35 &  x131 &  x146 &  x449 &  x572 &  x584 &  x662 &  x692 &  x827 &  x1088 &  x1097 & ~x90 & ~x129 & ~x231 & ~x336 & ~x459 & ~x588 & ~x706 & ~x745 & ~x784 & ~x1062;
assign c4128 =  x38 &  x159 &  x176 &  x198 &  x199 &  x209 &  x237 &  x239 &  x316 &  x575 &  x587 &  x716 &  x718 &  x797 &  x835 &  x836 &  x992 &  x1100 & ~x210 & ~x397;
assign c4130 =  x118 &  x120 &  x121 &  x157 &  x159 &  x160 &  x198 &  x199 &  x335 &  x640 & ~x127 & ~x1035;
assign c4132 =  x11 &  x16 &  x26 &  x35 &  x122 &  x125 &  x143 &  x221 &  x248 &  x254 &  x358 &  x367 &  x376 &  x385 &  x415 &  x445 &  x448 &  x494 &  x514 &  x530 &  x538 &  x554 &  x581 &  x584 &  x601 &  x632 &  x647 &  x650 &  x662 &  x689 &  x740 &  x806 &  x836 &  x952 &  x991 &  x1010 &  x1030 &  x1043 &  x1063 &  x1102 &  x1108;
assign c4134 =  x8 &  x38 &  x182 &  x200 &  x221 &  x299 &  x329 &  x410 &  x425 &  x434 &  x458 &  x494 &  x617 &  x716 &  x848 &  x929 &  x938 &  x956 &  x959 &  x989 &  x1043 &  x1094 &  x1112 &  x1121 & ~x411 & ~x420 & ~x450 & ~x504 & ~x534 & ~x543 & ~x573 & ~x582 & ~x612 & ~x690 & ~x696 & ~x729 & ~x774;
assign c4136 =  x364 & ~x45 & ~x51 & ~x801 & ~x825 & ~x846 & ~x1017 & ~x1071 & ~x1077 & ~x1095 & ~x1116;
assign c4138 =  x4 &  x40 &  x601 & ~x90 & ~x447 & ~x486 & ~x504 & ~x768 & ~x888 & ~x927;
assign c4140 =  x8 &  x113 &  x116 &  x119 &  x137 &  x155 &  x167 &  x212 &  x227 &  x280 &  x281 &  x290 &  x319 &  x332 &  x338 &  x416 &  x419 &  x422 &  x472 &  x473 &  x476 &  x500 &  x511 &  x569 &  x581 &  x586 &  x623 &  x671 &  x680 &  x713 &  x719 &  x770 &  x854 &  x881 &  x929 &  x953 &  x974 &  x1079 &  x1094 &  x1100 &  x1118 &  x1127 & ~x195 & ~x399 & ~x477 & ~x504 & ~x516 & ~x543 & ~x591 & ~x1017;
assign c4142 =  x5 &  x8 &  x20 &  x38 &  x59 &  x65 &  x68 &  x71 &  x95 &  x134 &  x143 &  x149 &  x158 &  x173 &  x179 &  x185 &  x197 &  x212 &  x215 &  x236 &  x254 &  x281 &  x308 &  x320 &  x323 &  x335 &  x356 &  x386 &  x407 &  x410 &  x413 &  x431 &  x452 &  x458 &  x461 &  x476 &  x485 &  x494 &  x497 &  x518 &  x524 &  x527 &  x533 &  x542 &  x548 &  x572 &  x587 &  x596 &  x599 &  x611 &  x617 &  x623 &  x644 &  x647 &  x650 &  x671 &  x677 &  x686 &  x689 &  x698 &  x701 &  x722 &  x734 &  x740 &  x755 &  x758 &  x767 &  x770 &  x782 &  x791 &  x793 &  x794 &  x815 &  x821 &  x869 &  x878 &  x902 &  x908 &  x911 &  x920 &  x926 &  x944 &  x1016 &  x1028 &  x1037 &  x1040 &  x1043 &  x1046 &  x1055 &  x1061 &  x1067 &  x1070 &  x1091 &  x1097 &  x1103 &  x1106 &  x1121 &  x1127 & ~x426 & ~x438 & ~x465 & ~x504 & ~x528 & ~x534 & ~x567 & ~x573 & ~x699 & ~x738 & ~x777 & ~x816 & ~x855;
assign c4144 =  x38 &  x128 &  x142 &  x202 &  x241 &  x318 &  x653 &  x719 &  x929 &  x932 &  x977 & ~x273 & ~x478;
assign c4146 =  x31 &  x70 &  x109 &  x499 &  x538 & ~x321 & ~x573 & ~x891 & ~x1008 & ~x1009;
assign c4148 =  x2 &  x5 &  x8 &  x32 &  x116 &  x125 &  x128 &  x143 &  x182 &  x202 &  x206 &  x241 &  x280 &  x296 &  x319 &  x323 &  x329 &  x362 &  x365 &  x380 &  x419 &  x428 &  x437 &  x446 &  x455 &  x470 &  x512 &  x530 &  x542 &  x599 &  x614 &  x647 &  x659 &  x683 &  x689 &  x701 &  x716 &  x761 &  x767 &  x770 &  x779 &  x902 &  x907 &  x917 &  x950 &  x953 &  x983 &  x998 &  x1019 &  x1043 &  x1046 &  x1064 &  x1085 &  x1097 & ~x438 & ~x786 & ~x825 & ~x864 & ~x903 & ~x978 & ~x1017 & ~x1056 & ~x1095;
assign c4150 =  x142 &  x227 &  x413 &  x749 &  x1079 & ~x27 & ~x132 & ~x150 & ~x210 & ~x249 & ~x261 & ~x288 & ~x345 & ~x444 & ~x810 & ~x840 & ~x879;
assign c4152 =  x26 &  x182 &  x239 &  x494 &  x499 &  x533 &  x538 &  x578 &  x745 &  x752 &  x784 &  x819 &  x905 &  x932 &  x940 &  x1085 & ~x882 & ~x888 & ~x903 & ~x960;
assign c4154 =  x191 &  x212 &  x248 &  x251 &  x308 &  x326 &  x344 &  x380 &  x452 &  x623 &  x637 &  x653 &  x755 &  x796 &  x835 &  x913 &  x952 &  x1031 &  x1070 & ~x399 & ~x435 & ~x475 & ~x514 & ~x553;
assign c4156 =  x780 &  x907 & ~x543 & ~x582 & ~x621 & ~x786 & ~x810 & ~x849 & ~x855 & ~x864 & ~x894 & ~x933;
assign c4158 =  x2 &  x68 &  x116 &  x176 &  x200 &  x215 &  x221 &  x250 &  x275 &  x290 &  x319 &  x374 &  x422 &  x547 &  x566 &  x575 &  x718 &  x722 &  x757 &  x791 &  x796 &  x824 &  x835 &  x914 &  x923 &  x952 &  x991 &  x1030 &  x1037 &  x1049 &  x1069 &  x1103 &  x1108 &  x1126 & ~x1017 & ~x1056;
assign c4160 =  x202 &  x218 &  x319 &  x323 &  x952 &  x991 &  x1030 &  x1069 &  x1103 &  x1108 & ~x321 & ~x771 & ~x810 & ~x849 & ~x855 & ~x894 & ~x933;
assign c4162 =  x20 &  x487 &  x780 &  x985 & ~x786 & ~x787 & ~x825 & ~x826 & ~x864 & ~x865 & ~x903 & ~x904 & ~x942 & ~x981;
assign c4164 =  x4 &  x22 &  x40 &  x43 &  x47 &  x53 &  x79 &  x104 &  x131 &  x167 &  x203 &  x209 &  x242 &  x341 &  x350 &  x356 &  x359 &  x391 &  x407 &  x413 &  x416 &  x458 &  x484 &  x488 &  x530 &  x545 &  x560 &  x562 &  x578 &  x601 &  x617 &  x629 &  x632 &  x665 &  x679 &  x718 &  x731 &  x734 &  x757 &  x761 &  x796 &  x797 &  x835 &  x839 &  x857 &  x874 &  x884 &  x1016 &  x1019 &  x1061 &  x1103 & ~x24 & ~x348 & ~x381 & ~x387 & ~x822 & ~x1017;
assign c4166 =  x601 &  x640 &  x655 & ~x982 & ~x996 & ~x1060 & ~x1099;
assign c4168 =  x121 &  x160 &  x198 &  x199 &  x266 &  x601 &  x640 &  x679 &  x718 &  x796 &  x835 &  x959 &  x1004 &  x1046 & ~x54 & ~x99 & ~x336 & ~x705;
assign c4170 =  x20 &  x28 &  x32 &  x40 &  x79 &  x143 &  x149 &  x170 &  x197 &  x272 &  x314 &  x350 &  x380 &  x407 &  x440 &  x457 &  x479 &  x500 &  x538 &  x562 &  x601 &  x604 &  x613 &  x629 &  x652 &  x656 &  x658 &  x659 &  x691 &  x718 &  x743 &  x785 &  x796 &  x835 &  x869 &  x884 &  x965 &  x977 &  x1085 &  x1088 &  x1108 &  x1120;
assign c4172 =  x38 &  x41 &  x71 &  x74 &  x83 &  x119 &  x122 &  x146 &  x167 &  x179 &  x206 &  x212 &  x227 &  x247 &  x278 &  x287 &  x290 &  x296 &  x308 &  x329 &  x335 &  x368 &  x380 &  x383 &  x428 &  x431 &  x458 &  x461 &  x470 &  x476 &  x494 &  x503 &  x524 &  x542 &  x545 &  x557 &  x565 &  x587 &  x599 &  x604 &  x627 &  x632 &  x641 &  x647 &  x701 &  x716 &  x731 &  x734 &  x743 &  x749 &  x770 &  x773 &  x794 &  x800 &  x848 &  x893 &  x911 &  x926 &  x938 &  x965 &  x968 &  x974 &  x998 &  x1052 &  x1073 &  x1088 &  x1103 & ~x429 & ~x468 & ~x747 & ~x801;
assign c4174 =  x128 &  x146 &  x188 &  x221 &  x224 &  x238 &  x242 &  x305 &  x316 &  x509 &  x524 &  x536 &  x596 &  x598 &  x611 &  x620 &  x659 &  x695 &  x718 &  x734 &  x757 &  x764 &  x796 &  x835 &  x913 &  x926 &  x952 &  x974 &  x991 &  x1049 &  x1052 &  x1073 &  x1085 & ~x435 & ~x436 & ~x588 & ~x591 & ~x666;
assign c4176 =  x664 &  x986 & ~x423 & ~x501 & ~x579 & ~x618 & ~x696 & ~x762 & ~x786 & ~x801 & ~x840 & ~x924 & ~x963 & ~x966 & ~x1056;
assign c4178 =  x50 &  x83 &  x551 &  x716 &  x737 &  x860 &  x1079 & ~x21 & ~x60 & ~x216 & ~x288 & ~x618 & ~x735 & ~x801 & ~x807 & ~x840 & ~x841 & ~x879 & ~x918 & ~x924 & ~x963 & ~x1005 & ~x1080 & ~x1083;
assign c4180 = ~x51 & ~x288 & ~x576 & ~x577 & ~x615 & ~x861 & ~x1017 & ~x1056;
assign c4182 =  x8 &  x50 &  x86 &  x107 &  x223 &  x233 &  x257 &  x281 &  x425 &  x440 &  x446 &  x550 &  x716 &  x731 &  x908 &  x932 &  x991 &  x1030 &  x1088 & ~x429 & ~x594 & ~x633 & ~x732 & ~x771 & ~x810 & ~x849 & ~x888 & ~x966 & ~x1005;
assign c4184 =  x2 &  x17 &  x41 &  x101 &  x120 &  x121 &  x143 &  x146 &  x159 &  x160 &  x173 &  x196 &  x198 &  x199 &  x200 &  x230 &  x233 &  x235 &  x237 &  x299 &  x308 &  x316 &  x350 &  x355 &  x386 &  x410 &  x413 &  x461 &  x464 &  x476 &  x491 &  x517 &  x518 &  x545 &  x554 &  x557 &  x584 &  x590 &  x593 &  x608 &  x728 &  x836 &  x929 &  x935 &  x947 &  x956 &  x989 &  x1010 &  x1016 &  x1045 &  x1058 &  x1118 & ~x279 & ~x319 & ~x358;
assign c4186 =  x627 & ~x826 & ~x864 & ~x865 & ~x904 & ~x942;
assign c4188 =  x8 &  x70 &  x77 &  x101 &  x104 &  x109 &  x110 &  x131 &  x173 &  x191 &  x227 &  x230 &  x233 &  x248 &  x278 &  x296 &  x311 &  x317 &  x350 &  x356 &  x362 &  x407 &  x410 &  x416 &  x428 &  x455 &  x518 &  x527 &  x536 &  x539 &  x572 &  x668 &  x689 &  x704 &  x722 &  x725 &  x743 &  x827 &  x836 &  x932 &  x947 &  x977 &  x1031 &  x1043 &  x1046 &  x1063 &  x1088 &  x1091 &  x1130 & ~x321 & ~x696 & ~x735 & ~x774 & ~x903 & ~x942 & ~x943 & ~x981 & ~x982;
assign c4190 =  x97 &  x175 &  x184 &  x185 &  x206 &  x223 &  x323 &  x395 &  x421 &  x436 &  x500 &  x577 &  x691 &  x884 &  x991 &  x1007 &  x1030 &  x1069 &  x1073 &  x1102 &  x1108 & ~x273;
assign c4192 =  x98 &  x212 &  x428 &  x545 &  x572 &  x947 & ~x51 & ~x615 & ~x762 & ~x774 & ~x801 & ~x822 & ~x1017 & ~x1056 & ~x1057 & ~x1095;
assign c4194 =  x56 &  x65 &  x80 &  x83 &  x101 &  x188 &  x196 &  x359 &  x371 &  x401 &  x476 &  x482 &  x523 &  x527 &  x530 &  x601 &  x623 &  x640 &  x679 &  x718 &  x730 &  x746 &  x752 &  x757 &  x796 &  x832 &  x835 &  x844 &  x871 &  x929 &  x1039 &  x1070 & ~x345 & ~x384 & ~x666;
assign c4196 =  x65 &  x86 &  x257 &  x269 &  x332 &  x380 &  x952 &  x1067 &  x1069 & ~x15 & ~x60 & ~x309 & ~x327 & ~x423 & ~x645 & ~x684;
assign c4198 =  x1 &  x2 &  x4 &  x20 &  x40 &  x43 &  x50 &  x79 &  x82 &  x86 &  x95 &  x101 &  x118 &  x121 &  x143 &  x149 &  x158 &  x170 &  x196 &  x200 &  x203 &  x227 &  x275 &  x302 &  x308 &  x323 &  x326 &  x356 &  x371 &  x386 &  x410 &  x419 &  x455 &  x461 &  x485 &  x497 &  x518 &  x533 &  x538 &  x578 &  x587 &  x601 &  x617 &  x635 &  x638 &  x640 &  x650 &  x656 &  x679 &  x683 &  x692 &  x701 &  x718 &  x725 &  x746 &  x752 &  x755 &  x757 &  x767 &  x794 &  x796 &  x797 &  x800 &  x806 &  x815 &  x824 &  x827 &  x835 &  x845 &  x854 &  x857 &  x872 &  x905 &  x916 &  x923 &  x929 &  x941 &  x959 &  x977 &  x995 &  x1013 &  x1022 &  x1043 &  x1049 &  x1052 &  x1061 &  x1067 &  x1076 &  x1094 & ~x51 & ~x90 & ~x192 & ~x309 & ~x348 & ~x504;
assign c4200 =  x56 &  x158 &  x167 &  x182 &  x247 &  x248 &  x263 &  x331 &  x376 &  x397 &  x415 &  x421 &  x448 &  x461 &  x473 &  x499 &  x506 &  x514 &  x533 &  x538 &  x539 &  x545 &  x568 &  x577 &  x587 &  x623 &  x632 &  x638 &  x656 &  x677 &  x680 &  x836 &  x862 &  x901 &  x929 &  x980 &  x1037 &  x1043 &  x1046 &  x1049 &  x1054 &  x1061 &  x1067 &  x1085 &  x1124 &  x1127 & ~x750;
assign c4202 =  x5 &  x8 &  x11 &  x17 &  x26 &  x29 &  x41 &  x44 &  x50 &  x65 &  x74 &  x77 &  x86 &  x89 &  x92 &  x95 &  x107 &  x113 &  x128 &  x131 &  x140 &  x149 &  x161 &  x173 &  x176 &  x179 &  x185 &  x206 &  x212 &  x218 &  x221 &  x227 &  x239 &  x248 &  x257 &  x260 &  x263 &  x266 &  x272 &  x278 &  x284 &  x296 &  x299 &  x305 &  x311 &  x314 &  x323 &  x326 &  x329 &  x332 &  x335 &  x338 &  x344 &  x353 &  x356 &  x359 &  x371 &  x374 &  x377 &  x386 &  x394 &  x395 &  x401 &  x404 &  x413 &  x422 &  x431 &  x446 &  x455 &  x467 &  x470 &  x473 &  x488 &  x491 &  x494 &  x497 &  x500 &  x506 &  x508 &  x521 &  x524 &  x533 &  x536 &  x547 &  x554 &  x557 &  x560 &  x563 &  x566 &  x572 &  x575 &  x584 &  x587 &  x590 &  x599 &  x602 &  x608 &  x614 &  x617 &  x629 &  x632 &  x635 &  x637 &  x638 &  x650 &  x653 &  x659 &  x662 &  x668 &  x674 &  x675 &  x680 &  x695 &  x698 &  x704 &  x707 &  x715 &  x719 &  x728 &  x731 &  x737 &  x740 &  x746 &  x752 &  x755 &  x767 &  x770 &  x773 &  x785 &  x788 &  x818 &  x824 &  x827 &  x842 &  x845 &  x848 &  x851 &  x854 &  x857 &  x863 &  x869 &  x872 &  x878 &  x881 &  x884 &  x887 &  x890 &  x893 &  x899 &  x911 &  x914 &  x923 &  x926 &  x929 &  x935 &  x938 &  x941 &  x944 &  x947 &  x950 &  x953 &  x968 &  x977 &  x980 &  x983 &  x992 &  x995 &  x1004 &  x1007 &  x1016 &  x1028 &  x1034 &  x1040 &  x1043 &  x1046 &  x1067 &  x1070 &  x1082 &  x1088 &  x1094 &  x1103 &  x1115 &  x1118 & ~x438 & ~x534 & ~x552 & ~x573 & ~x591 & ~x615;
assign c4204 =  x65 &  x89 &  x98 &  x158 &  x278 &  x305 &  x323 &  x338 &  x350 &  x365 &  x371 &  x461 &  x488 &  x524 &  x542 &  x545 &  x557 &  x578 &  x602 &  x665 &  x719 &  x734 &  x812 &  x950 &  x1022 &  x1094 &  x1109 & ~x15 & ~x54 & ~x78 & ~x93 & ~x132 & ~x150 & ~x171 & ~x189 & ~x228 & ~x249 & ~x288 & ~x321 & ~x378 & ~x495 & ~x534 & ~x540 & ~x573 & ~x678 & ~x774 & ~x813;
assign c4206 =  x2 &  x25 &  x64 &  x70 &  x109 &  x212 &  x233 &  x311 &  x350 &  x419 &  x476 &  x647 &  x752 &  x815 &  x836 &  x845 &  x890 &  x1052 &  x1085 & ~x78 & ~x111 & ~x411 & ~x450 & ~x534 & ~x723 & ~x762 & ~x801 & ~x1008;
assign c4208 =  x44 &  x788 &  x859 &  x866 &  x872 &  x901 &  x987 &  x1079 &  x1103 & ~x826 & ~x865 & ~x903 & ~x942 & ~x943 & ~x981;
assign c4210 =  x70 &  x237 &  x276 &  x545 &  x634 &  x668 & ~x189 & ~x210 & ~x1017;
assign c4212 =  x2 &  x8 &  x11 &  x29 &  x44 &  x47 &  x65 &  x71 &  x74 &  x104 &  x110 &  x113 &  x119 &  x146 &  x152 &  x155 &  x158 &  x176 &  x182 &  x188 &  x212 &  x227 &  x257 &  x272 &  x278 &  x290 &  x296 &  x302 &  x308 &  x329 &  x350 &  x371 &  x380 &  x410 &  x413 &  x440 &  x491 &  x494 &  x512 &  x518 &  x521 &  x551 &  x605 &  x623 &  x626 &  x644 &  x668 &  x671 &  x689 &  x701 &  x718 &  x737 &  x740 &  x776 &  x785 &  x791 &  x854 &  x878 &  x902 &  x932 &  x938 &  x998 &  x1001 &  x1028 &  x1067 &  x1070 &  x1094 &  x1100 &  x1106 &  x1121 & ~x15 & ~x33 & ~x51 & ~x225 & ~x384 & ~x423 & ~x426 & ~x930;
assign c4214 =  x20 &  x86 &  x89 &  x116 &  x125 &  x131 &  x164 &  x170 &  x182 &  x194 &  x224 &  x227 &  x233 &  x239 &  x248 &  x278 &  x287 &  x308 &  x332 &  x344 &  x350 &  x359 &  x398 &  x401 &  x431 &  x458 &  x470 &  x512 &  x539 &  x550 &  x569 &  x578 &  x608 &  x625 &  x656 &  x671 &  x677 &  x719 &  x737 &  x770 &  x785 &  x788 &  x815 &  x820 &  x867 &  x875 &  x893 &  x905 &  x907 &  x935 &  x956 &  x986 &  x989 &  x1067 &  x1070 &  x1073 &  x1103 &  x1115 &  x1121 & ~x748 & ~x786 & ~x787 & ~x825 & ~x826;
assign c4216 =  x22 &  x28 &  x61 &  x82 &  x184 &  x295 &  x640 &  x679 &  x718 &  x796 &  x835 &  x952 &  x1016 &  x1052 & ~x63 & ~x582 & ~x816;
assign c4218 =  x25 &  x38 &  x64 &  x68 &  x70 &  x77 &  x143 &  x158 &  x167 &  x170 &  x203 &  x284 &  x290 &  x315 &  x316 &  x398 &  x443 &  x497 &  x545 &  x578 &  x587 &  x593 &  x595 &  x626 &  x634 &  x638 &  x650 &  x656 &  x677 &  x695 &  x719 &  x725 &  x749 &  x757 &  x836 &  x874 &  x887 &  x902 &  x1064 &  x1121 & ~x189 & ~x435;
assign c4220 =  x29 &  x110 &  x176 &  x179 &  x182 &  x198 &  x199 &  x203 &  x238 &  x275 &  x350 &  x371 &  x380 &  x395 &  x407 &  x509 &  x560 &  x575 &  x593 &  x671 &  x761 &  x791 &  x875 &  x1034 &  x1103 &  x1109 &  x1127 & ~x15 & ~x33 & ~x54 & ~x72 & ~x93 & ~x435 & ~x666 & ~x930;
assign c4222 =  x29 &  x41 &  x50 &  x59 &  x83 &  x110 &  x167 &  x202 &  x230 &  x241 &  x242 &  x245 &  x263 &  x280 &  x320 &  x323 &  x368 &  x416 &  x446 &  x548 &  x566 &  x581 &  x674 &  x707 &  x751 &  x755 &  x790 &  x821 &  x851 &  x857 &  x914 &  x950 &  x968 &  x977 &  x980 &  x1031 &  x1079 & ~x708 & ~x783 & ~x978 & ~x1017 & ~x1032 & ~x1056 & ~x1071 & ~x1077 & ~x1095 & ~x1110;
assign c4224 =  x326 &  x413 &  x446 &  x494 &  x509 &  x520 &  x562 &  x587 &  x596 &  x601 &  x640 &  x689 &  x743 &  x779 &  x854 &  x973 &  x1013 &  x1019 &  x1039 &  x1073 &  x1094 & ~x411 & ~x435 & ~x978 & ~x1056 & ~x1095;
assign c4226 =  x112 &  x250 &  x415 &  x836 &  x985 &  x1024 &  x1030 & ~x786 & ~x972 & ~x1044;
assign c4228 =  x43 &  x80 &  x82 &  x121 &  x146 &  x160 &  x188 &  x199 &  x212 &  x230 &  x263 &  x308 &  x347 &  x506 &  x601 &  x611 &  x659 &  x679 &  x718 &  x757 &  x776 &  x788 &  x796 &  x835 &  x869 &  x896 &  x910 &  x935 &  x950 &  x967 &  x980 &  x1039 &  x1045 &  x1078 &  x1084 &  x1097 &  x1117 & ~x462 & ~x474;
assign c4230 =  x4 &  x43 &  x53 &  x68 &  x79 &  x82 &  x118 &  x329 &  x335 &  x458 &  x596 &  x601 &  x614 &  x679 &  x718 &  x743 &  x796 &  x832 &  x835 &  x1061 & ~x51 & ~x90 & ~x102 & ~x108 & ~x147 & ~x186 & ~x348 & ~x387;
assign c4232 =  x11 &  x56 &  x59 &  x77 &  x92 &  x98 &  x113 &  x116 &  x119 &  x122 &  x128 &  x140 &  x143 &  x155 &  x164 &  x185 &  x191 &  x197 &  x227 &  x245 &  x248 &  x263 &  x284 &  x319 &  x329 &  x374 &  x455 &  x458 &  x476 &  x491 &  x497 &  x506 &  x510 &  x518 &  x551 &  x602 &  x614 &  x662 &  x665 &  x667 &  x671 &  x695 &  x713 &  x737 &  x746 &  x752 &  x755 &  x785 &  x794 &  x800 &  x829 &  x860 &  x866 &  x884 &  x932 &  x938 &  x944 &  x959 &  x962 &  x974 &  x977 &  x1004 &  x1028 &  x1031 &  x1043 &  x1049 &  x1061 &  x1088 &  x1100 &  x1112 &  x1127 & ~x645 & ~x669 & ~x684 & ~x708 & ~x723 & ~x747;
assign c4234 =  x74 &  x107 &  x110 &  x122 &  x194 &  x265 &  x301 &  x356 &  x371 &  x376 &  x389 &  x397 &  x415 &  x436 &  x464 &  x470 &  x479 &  x491 &  x542 &  x554 &  x566 &  x608 &  x614 &  x620 &  x628 &  x710 &  x716 &  x725 &  x776 &  x815 &  x824 &  x832 &  x845 &  x890 &  x905 &  x944 &  x962 &  x992 &  x998 &  x1010 &  x1064 &  x1073 &  x1094 &  x1103 & ~x594 & ~x595 & ~x633;
assign c4236 =  x22 &  x28 &  x73 &  x92 &  x101 &  x112 &  x133 &  x139 &  x140 &  x167 &  x172 &  x184 &  x223 &  x229 &  x250 &  x266 &  x346 &  x496 &  x518 &  x569 &  x710 &  x718 &  x731 &  x742 &  x796 &  x820 &  x830 &  x835 &  x913 &  x989 &  x1103 & ~x738 & ~x777;
assign c4238 =  x98 &  x113 &  x203 &  x284 &  x347 &  x380 &  x476 &  x497 &  x551 &  x575 &  x577 &  x599 &  x605 &  x626 &  x638 &  x683 &  x698 &  x764 &  x780 &  x782 &  x785 &  x854 &  x898 &  x899 &  x913 &  x914 &  x941 &  x947 &  x983 &  x992 &  x1016 &  x1043 &  x1052 &  x1054 &  x1102 & ~x855 & ~x864 & ~x1059;
assign c4240 =  x62 &  x74 &  x80 &  x113 &  x125 &  x128 &  x158 &  x191 &  x224 &  x227 &  x238 &  x239 &  x276 &  x278 &  x293 &  x302 &  x308 &  x315 &  x320 &  x329 &  x377 &  x389 &  x419 &  x422 &  x428 &  x469 &  x470 &  x497 &  x509 &  x524 &  x542 &  x545 &  x566 &  x581 &  x587 &  x653 &  x668 &  x680 &  x683 &  x707 &  x779 &  x827 &  x830 &  x851 &  x866 &  x893 &  x896 &  x935 &  x941 &  x944 &  x968 &  x971 &  x977 &  x1001 &  x1019 &  x1064 &  x1079 &  x1124 & ~x78 & ~x189 & ~x228 & ~x435 & ~x474 & ~x475 & ~x513 & ~x591 & ~x783 & ~x822;
assign c4242 =  x101 &  x113 &  x188 &  x247 &  x266 &  x272 &  x314 &  x371 &  x410 &  x422 &  x482 &  x494 &  x515 &  x587 &  x638 &  x758 &  x770 &  x890 &  x896 &  x923 &  x944 &  x1022 &  x1058 &  x1064 &  x1076 &  x1079 &  x1103 & ~x60 & ~x99 & ~x216 & ~x255 & ~x288 & ~x501 & ~x540 & ~x579 & ~x672 & ~x840 & ~x918 & ~x924 & ~x927 & ~x963 & ~x966;
assign c4244 =  x2 &  x281 &  x329 &  x476 &  x508 &  x557 &  x734 &  x1046 &  x1073 &  x1085 & ~x321 & ~x411 & ~x450 & ~x474 & ~x475 & ~x489 & ~x514 & ~x528 & ~x567 & ~x978 & ~x1017 & ~x1056 & ~x1095;
assign c4246 =  x7 &  x23 &  x101 &  x131 &  x194 &  x278 &  x290 &  x335 &  x341 &  x359 &  x380 &  x416 &  x431 &  x440 &  x446 &  x470 &  x517 &  x523 &  x601 &  x617 &  x623 &  x640 &  x644 &  x668 &  x679 &  x689 &  x718 &  x743 &  x758 &  x812 &  x857 &  x911 &  x935 &  x949 &  x953 &  x1016 &  x1046 &  x1064 &  x1065 &  x1097 &  x1100 &  x1105 & ~x435;
assign c4248 =  x140 &  x260 &  x335 &  x706 &  x770 &  x867 &  x868 &  x908 &  x941 &  x946 &  x1109 & ~x723 & ~x786 & ~x787 & ~x825 & ~x826 & ~x864 & ~x903;
assign c4250 =  x125 &  x136 &  x175 &  x193 &  x226 &  x280 &  x323 &  x383 &  x410 &  x449 &  x471 &  x677 &  x679 &  x718 &  x796 &  x835 &  x874;
assign c4252 =  x198 &  x237 &  x517 &  x718 &  x1039 &  x1078 & ~x319 & ~x358 & ~x397;
assign c4254 =  x383 & ~x15 & ~x54 & ~x93 & ~x204 & ~x210 & ~x249 & ~x288 & ~x327 & ~x411 & ~x459 & ~x498 & ~x1017 & ~x1023 & ~x1056 & ~x1062 & ~x1095;
assign c4256 =  x155 &  x199 &  x237 &  x314 &  x383 &  x464 &  x521 &  x595 &  x601 &  x634 &  x640 &  x679 &  x728 &  x757 &  x796 &  x835 & ~x210 & ~x435;
assign c4258 =  x2 &  x11 &  x59 &  x134 &  x302 &  x308 &  x316 &  x467 &  x503 &  x634 &  x672 &  x785 &  x1070 &  x1103 & ~x435 & ~x474 & ~x475 & ~x514 & ~x528 & ~x567;
assign c4260 =  x121 &  x160 &  x199 &  x335 &  x406 &  x562 &  x601 &  x602 &  x640 &  x679 &  x689 &  x718 &  x973 &  x1084 & ~x306 & ~x345 & ~x384 & ~x423;
assign c4262 =  x37 &  x65 &  x68 &  x110 &  x134 &  x215 &  x371 &  x377 &  x470 &  x557 &  x635 &  x692 &  x752 &  x818 &  x835 &  x874 &  x913 &  x917 &  x956 &  x991 &  x1030 &  x1037 & ~x360 & ~x774 & ~x855 & ~x894 & ~x933;
assign c4264 =  x41 &  x71 &  x221 &  x233 &  x245 &  x314 &  x329 &  x395 &  x401 &  x413 &  x443 &  x446 &  x449 &  x476 &  x536 &  x538 &  x569 &  x701 &  x740 &  x797 &  x842 &  x863 &  x869 &  x905 &  x914 &  x1037 &  x1054 &  x1067 &  x1070 &  x1115 & ~x729 & ~x852 & ~x903 & ~x942 & ~x981 & ~x996 & ~x1020;
assign c4266 =  x80 &  x83 &  x98 &  x119 &  x125 &  x260 &  x287 &  x311 &  x347 &  x469 &  x470 &  x476 &  x488 &  x503 &  x508 &  x548 &  x554 &  x634 &  x637 &  x650 &  x672 &  x713 &  x743 &  x791 &  x796 &  x803 &  x812 &  x821 &  x824 &  x835 &  x836 &  x881 &  x890 &  x1013 &  x1061 &  x1103 &  x1112 & ~x411 & ~x450 & ~x489;
assign c4268 =  x14 &  x25 &  x26 &  x53 &  x64 &  x89 &  x103 &  x181 &  x212 &  x220 &  x236 &  x239 &  x265 &  x272 &  x275 &  x323 &  x350 &  x368 &  x394 &  x395 &  x410 &  x428 &  x461 &  x503 &  x509 &  x518 &  x542 &  x545 &  x563 &  x689 &  x695 &  x812 &  x893 &  x926 &  x952 &  x983 &  x991 &  x1030 &  x1031 &  x1034 &  x1037 &  x1052 & ~x78 & ~x321 & ~x477;
assign c4270 =  x82 &  x121 &  x160 &  x198 &  x237 &  x517 &  x835 & ~x319 & ~x358 & ~x397 & ~x435;
assign c4272 =  x8 &  x14 &  x23 &  x38 &  x43 &  x68 &  x82 &  x107 &  x110 &  x116 &  x125 &  x143 &  x160 &  x167 &  x170 &  x197 &  x199 &  x221 &  x224 &  x233 &  x248 &  x251 &  x263 &  x284 &  x287 &  x290 &  x335 &  x347 &  x352 &  x353 &  x383 &  x386 &  x389 &  x437 &  x443 &  x446 &  x458 &  x467 &  x482 &  x500 &  x503 &  x515 &  x519 &  x530 &  x536 &  x539 &  x569 &  x581 &  x614 &  x635 &  x641 &  x668 &  x677 &  x679 &  x695 &  x707 &  x716 &  x740 &  x752 &  x776 &  x812 &  x830 &  x842 &  x860 &  x869 &  x887 &  x911 &  x914 &  x917 &  x935 &  x953 &  x962 &  x977 &  x992 &  x1010 &  x1039 &  x1052 &  x1078 &  x1091 &  x1094 &  x1124 &  x1127 & ~x435;
assign c4274 =  x29 &  x86 &  x233 &  x332 &  x425 &  x487 &  x553 &  x577 &  x604 &  x605 &  x680 &  x705 &  x959 &  x1043 & ~x888 & ~x927 & ~x942 & ~x966 & ~x981;
assign c4276 =  x199 &  x287 &  x311 &  x315 &  x316 &  x410 &  x458 &  x566 &  x595 &  x601 &  x679 &  x718 &  x757 &  x796 &  x803 &  x835 &  x917 &  x1031 & ~x435 & ~x475 & ~x552;
assign c4278 =  x28 &  x65 &  x145 &  x913 &  x1022 &  x1108 & ~x90 & ~x108 & ~x738 & ~x933 & ~x1044 & ~x1077 & ~x1110;
assign c4280 =  x85 &  x121 &  x123 &  x124 &  x159 &  x160 &  x198 &  x199 &  x237 &  x276 &  x290 &  x315 &  x374 &  x386 &  x479 &  x842 &  x866 &  x953 &  x1121 & ~x228;
assign c4282 =  x95 &  x101 &  x104 &  x350 &  x497 &  x604 &  x679 &  x718 &  x757 &  x793 &  x796 &  x800 &  x967 & ~x384 & ~x387 & ~x423 & ~x426 & ~x462;
assign c4284 =  x2 &  x3 &  x4 &  x11 &  x35 &  x40 &  x42 &  x43 &  x44 &  x50 &  x53 &  x79 &  x81 &  x82 &  x89 &  x92 &  x101 &  x107 &  x116 &  x118 &  x120 &  x121 &  x122 &  x125 &  x128 &  x146 &  x155 &  x159 &  x160 &  x167 &  x176 &  x179 &  x185 &  x194 &  x199 &  x203 &  x206 &  x212 &  x215 &  x233 &  x257 &  x263 &  x266 &  x269 &  x272 &  x281 &  x284 &  x290 &  x293 &  x299 &  x302 &  x311 &  x323 &  x332 &  x350 &  x359 &  x362 &  x374 &  x377 &  x380 &  x383 &  x386 &  x389 &  x395 &  x410 &  x419 &  x428 &  x443 &  x446 &  x467 &  x473 &  x479 &  x482 &  x485 &  x497 &  x500 &  x512 &  x524 &  x545 &  x554 &  x563 &  x572 &  x578 &  x581 &  x587 &  x596 &  x599 &  x601 &  x605 &  x608 &  x623 &  x626 &  x640 &  x641 &  x647 &  x659 &  x671 &  x686 &  x692 &  x698 &  x716 &  x719 &  x725 &  x746 &  x770 &  x779 &  x782 &  x785 &  x791 &  x794 &  x800 &  x803 &  x812 &  x815 &  x818 &  x824 &  x845 &  x857 &  x872 &  x887 &  x896 &  x902 &  x905 &  x911 &  x920 &  x941 &  x968 &  x974 &  x989 &  x992 &  x995 &  x1001 &  x1025 &  x1031 &  x1046 &  x1049 &  x1058 &  x1064 &  x1067 &  x1085 &  x1097 &  x1100 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 & ~x9 & ~x48 & ~x60 & ~x780 & ~x858;
assign c4286 =  x353 &  x475 &  x568 &  x952 &  x990 &  x991 &  x1030 & ~x891 & ~x930 & ~x1020;
assign c4288 =  x23 &  x113 &  x194 &  x260 &  x263 &  x305 &  x371 &  x395 &  x557 &  x575 &  x680 &  x1127 & ~x723 & ~x762 & ~x786 & ~x801 & ~x825 & ~x840 & ~x879 & ~x885 & ~x924 & ~x963 & ~x1008 & ~x1056 & ~x1071 & ~x1095 & ~x1116;
assign c4290 =  x25 &  x64 &  x237 &  x276 &  x355 &  x679 &  x718 & ~x435 & ~x436 & ~x475;
assign c4292 =  x233 &  x371 &  x392 &  x473 &  x485 &  x572 &  x695 &  x701 &  x785 &  x1001 &  x1052 &  x1103 & ~x654 & ~x669 & ~x708 & ~x810 & ~x825 & ~x849 & ~x855 & ~x999 & ~x1017 & ~x1056 & ~x1095;
assign c4294 =  x319 &  x335 &  x359 &  x524 &  x796 &  x835 &  x913 &  x1103 &  x1112 & ~x525 & ~x738 & ~x777 & ~x778 & ~x816 & ~x1017 & ~x1056;
assign c4296 =  x149 &  x179 &  x188 &  x198 &  x199 &  x237 &  x257 &  x835 & ~x216 & ~x397;
assign c4298 =  x38 &  x120 &  x159 &  x167 &  x198 &  x199 &  x218 &  x238 &  x257 &  x260 &  x266 &  x344 &  x350 &  x377 &  x452 &  x557 &  x689 &  x764 &  x815 &  x827 &  x884 &  x1067 & ~x93 & ~x319 & ~x426 & ~x435;
assign c41 =  x152 &  x749 &  x1004 & ~x297 & ~x375 & ~x402 & ~x483 & ~x597 & ~x636 & ~x702 & ~x780;
assign c43 =  x410 &  x593 &  x631 &  x688 &  x766 &  x773 &  x793 &  x805 &  x844 &  x848 &  x1031 &  x1046 & ~x264 & ~x303 & ~x328;
assign c45 =  x161 &  x282 &  x321 &  x399 & ~x117;
assign c47 =  x110 &  x167 &  x388 &  x458 &  x466 &  x596 &  x656 &  x665 &  x701 &  x749 &  x863 &  x935 &  x962 & ~x555 & ~x747 & ~x909 & ~x990 & ~x1068 & ~x1107;
assign c49 =  x214 &  x781 &  x978 &  x1056 & ~x6;
assign c411 = ~x471 & ~x949;
assign c413 =  x403 &  x605 &  x775 &  x976 & ~x312 & ~x792 & ~x870 & ~x987;
assign c415 =  x248 &  x253 &  x1093 & ~x126 & ~x687 & ~x714 & ~x831;
assign c417 =  x62 &  x548 &  x607 &  x688 &  x722 & ~x246 & ~x363 & ~x516 & ~x555 & ~x780;
assign c419 =  x130 &  x283 &  x321 &  x893 & ~x9 & ~x39;
assign c421 =  x20 &  x158 &  x364 &  x377 &  x395 &  x585 &  x663 &  x1085 & ~x354 & ~x471;
assign c423 =  x10 &  x11 &  x122 &  x188 &  x191 &  x233 &  x283 &  x547 &  x575 &  x680 &  x719 &  x959 & ~x714 & ~x753 & ~x831 & ~x870 & ~x948 & ~x987;
assign c425 =  x110 &  x321 &  x429 & ~x117;
assign c427 =  x529 & ~x123 & ~x162 & ~x246 & ~x906 & ~x1107;
assign c429 =  x188 &  x283 &  x317 &  x321 &  x360 &  x361 &  x400 &  x430 &  x464 &  x956 &  x1004 & ~x81 & ~x120;
assign c431 =  x156 & ~x162 & ~x286 & ~x325 & ~x364 & ~x780;
assign c433 =  x104 &  x191 &  x281 &  x416 &  x449 &  x617 &  x749 &  x823 &  x842 &  x911 &  x1018 &  x1022 &  x1028 &  x1057 & ~x756 & ~x795 & ~x831 & ~x834 & ~x873;
assign c435 =  x597 &  x751 & ~x391;
assign c437 =  x649 &  x709 &  x727 &  x817 &  x850 & ~x480 & ~x600;
assign c439 =  x340 &  x403 &  x594 &  x673 & ~x354 & ~x393 & ~x432 & ~x909 & ~x1026;
assign c441 =  x10 &  x49 &  x88 &  x127 &  x273 &  x488 &  x713 &  x947 & ~x516 & ~x585 & ~x780;
assign c443 =  x325 &  x370 &  x376 &  x403 &  x409 &  x555 &  x820 &  x1013;
assign c445 = ~x531 & ~x714 & ~x720 & ~x871;
assign c447 = ~x1066 & ~x1084 & ~x1105;
assign c449 =  x53 &  x89 &  x164 &  x227 &  x242 &  x263 &  x268 &  x287 &  x338 &  x362 &  x409 &  x412 &  x427 &  x451 &  x466 &  x476 &  x490 &  x529 &  x548 &  x593 &  x673 &  x716 &  x751 &  x773 &  x827 &  x848 &  x899 &  x905 &  x907 &  x959 &  x979 &  x1018 &  x1031 &  x1085 &  x1088;
assign c451 =  x38 &  x77 &  x101 &  x212 &  x494 &  x500 &  x632 &  x677 &  x761 &  x842 &  x872 &  x884 &  x899 &  x944 &  x1007 &  x1060 & ~x3 & ~x42 & ~x81 & ~x120 & ~x237 & ~x354 & ~x393 & ~x432 & ~x471 & ~x549;
assign c453 =  x113 &  x382 &  x674 &  x929 & ~x393 & ~x471 & ~x726 & ~x909 & ~x988 & ~x1065 & ~x1105;
assign c455 =  x62 &  x83 &  x100 &  x221 &  x502 &  x518 &  x556 &  x668 &  x673 &  x740 &  x965 &  x1034 &  x1046 &  x1079 & ~x354 & ~x432 & ~x837 & ~x876;
assign c457 =  x236 &  x380 &  x751 &  x1046 & ~x3 & ~x42 & ~x159 & ~x237 & ~x354 & ~x471 & ~x510 & ~x726;
assign c459 =  x5 &  x74 &  x80 &  x128 &  x170 &  x176 &  x206 &  x212 &  x215 &  x224 &  x242 &  x275 &  x287 &  x302 &  x320 &  x365 &  x422 &  x443 &  x482 &  x485 &  x494 &  x512 &  x518 &  x521 &  x563 &  x575 &  x617 &  x626 &  x680 &  x707 &  x716 &  x725 &  x773 &  x788 &  x791 &  x818 &  x875 &  x887 &  x935 &  x950 &  x979 &  x995 &  x1018 &  x1037 &  x1040 &  x1057 &  x1064 &  x1118 &  x1124 & ~x246 & ~x453 & ~x492 & ~x756 & ~x873;
assign c461 =  x624 & ~x234 & ~x471;
assign c463 =  x321 &  x399 &  x635 & ~x42 & ~x120;
assign c465 =  x625 &  x842 &  x1046 & ~x87 & ~x675 & ~x753 & ~x792 & ~x795 & ~x831 & ~x834;
assign c467 =  x271 &  x436 &  x806 &  x919 &  x1075 & ~x432 & ~x825 & ~x870;
assign c469 =  x631 & ~x364 & ~x483 & ~x519 & ~x780;
assign c471 =  x978 &  x1018 &  x1057 &  x1096 & ~x195 & ~x954 & ~x990;
assign c473 =  x89 &  x91 &  x431 &  x683 &  x898 &  x956 &  x1048 & ~x471 & ~x948 & ~x987;
assign c475 =  x2 &  x86 &  x232 &  x239 &  x263 &  x506 &  x536 &  x589 &  x632 &  x662 &  x749 &  x779 & ~x393 & ~x432 & ~x592;
assign c477 =  x204 &  x243 &  x322 &  x351 &  x390 &  x722 &  x983 &  x1058 & ~x81 & ~x357;
assign c479 =  x579 &  x618 & ~x3 & ~x531;
assign c481 =  x116 &  x137 &  x239 &  x248 &  x356 &  x674 &  x737 &  x742 &  x824 &  x902 &  x923 &  x1013 &  x1124 & ~x126 & ~x156 & ~x354 & ~x432 & ~x909 & ~x948 & ~x987 & ~x1026;
assign c483 =  x169 &  x283 &  x288 &  x327 &  x826 & ~x538;
assign c485 =  x427 &  x436 &  x1020 &  x1059;
assign c487 =  x514 &  x877 &  x889 & ~x444 & ~x483 & ~x780;
assign c489 =  x13 &  x347 &  x669 &  x747 &  x786 &  x825 &  x904;
assign c491 =  x137 &  x338 &  x388 &  x413 &  x686 &  x692 &  x701 &  x749 &  x1043 &  x1082 &  x1091 & ~x354 & ~x393 & ~x432 & ~x471 & ~x510 & ~x588 & ~x954 & ~x990;
assign c493 =  x91 &  x450 &  x805;
assign c495 =  x10 &  x205 &  x383 &  x502 &  x583 &  x775 &  x805 &  x970 &  x1009 & ~x330;
assign c497 =  x266 &  x452 &  x533 &  x581 &  x725 &  x797 &  x800 &  x1001 &  x1106 &  x1124 & ~x276 & ~x354 & ~x393 & ~x753 & ~x759 & ~x792 & ~x798 & ~x831 & ~x837 & ~x870 & ~x909 & ~x948;
assign c499 =  x766 &  x883 & ~x562 & ~x624;
assign c4101 =  x260 &  x341 &  x354 &  x591 &  x611 &  x1100 & ~x585;
assign c4103 =  x49 &  x88 &  x127 &  x234 &  x273 &  x740 &  x779 &  x824 & ~x585 & ~x780;
assign c4105 =  x32 &  x74 &  x77 &  x110 &  x128 &  x131 &  x155 &  x161 &  x200 &  x254 &  x260 &  x272 &  x281 &  x287 &  x305 &  x335 &  x338 &  x365 &  x401 &  x422 &  x449 &  x464 &  x482 &  x491 &  x497 &  x578 &  x581 &  x583 &  x605 &  x611 &  x617 &  x641 &  x647 &  x671 &  x674 &  x680 &  x686 &  x695 &  x698 &  x709 &  x716 &  x782 &  x785 &  x787 &  x803 &  x812 &  x815 &  x817 &  x839 &  x842 &  x848 &  x854 &  x887 &  x916 &  x923 &  x956 &  x959 &  x977 &  x980 &  x995 &  x1004 &  x1073 &  x1076 &  x1088 &  x1106 &  x1112 &  x1118 & ~x444 & ~x483 & ~x585 & ~x663 & ~x780 & ~x858;
assign c4107 =  x68 &  x71 &  x227 &  x338 &  x398 &  x1033 & ~x639 & ~x675 & ~x678 & ~x756 & ~x780;
assign c4109 =  x98 &  x188 &  x191 &  x302 &  x313 &  x326 &  x542 &  x608 &  x680 &  x688 &  x799 &  x805 &  x844 &  x917 &  x1066 &  x1090 & ~x402 & ~x441 & ~x780;
assign c4111 =  x455 &  x497 &  x629 &  x701 &  x926 & ~x354 & ~x792 & ~x831 & ~x870 & ~x871 & ~x909 & ~x948 & ~x1026 & ~x1065 & ~x1104;
assign c4113 =  x688 &  x709 & ~x523;
assign c4115 =  x547 &  x586 & ~x639 & ~x718 & ~x757;
assign c4117 =  x226 &  x251 &  x379 &  x515 &  x635 &  x728 &  x904 & ~x354 & ~x471 & ~x798;
assign c4119 =  x628 &  x703 & ~x87 & ~x675 & ~x714 & ~x795 & ~x831 & ~x870;
assign c4121 =  x50 &  x56 &  x65 &  x194 &  x197 &  x203 &  x218 &  x242 &  x254 &  x272 &  x296 &  x317 &  x383 &  x388 &  x398 &  x407 &  x427 &  x467 &  x473 &  x563 &  x578 &  x596 &  x635 &  x647 &  x673 &  x710 &  x751 &  x764 &  x812 &  x821 &  x833 &  x836 &  x848 &  x872 &  x875 &  x926 &  x935 &  x947 &  x968 &  x976 &  x1009 &  x1010 &  x1015 &  x1019 &  x1034 &  x1048 &  x1055 &  x1091 &  x1130 & ~x393 & ~x432 & ~x471 & ~x510 & ~x738;
assign c4123 =  x388 &  x451 &  x673 &  x1021 &  x1060 & ~x912;
assign c4125 =  x176 &  x302 &  x410 &  x462 &  x463 &  x502 &  x540 &  x580 &  x788 &  x1127 & ~x516 & ~x1041;
assign c4127 =  x736 &  x774 &  x775 &  x1008 & ~x870;
assign c4129 =  x51 &  x130 &  x814 & ~x828 & ~x945;
assign c4131 =  x775 &  x787 & ~x562;
assign c4133 =  x670 &  x877 &  x883 & ~x523;
assign c4135 =  x202 & ~x571 & ~x714 & ~x792 & ~x870;
assign c4137 =  x116 &  x146 &  x176 &  x188 &  x233 &  x263 &  x278 &  x433 &  x553 &  x592 &  x608 &  x631 &  x638 &  x670 &  x704 &  x709 &  x748 &  x767 &  x776 &  x787 &  x791 &  x794 &  x863 &  x905 &  x932 &  x955 &  x968 &  x1001 &  x1033 &  x1091 &  x1100 & ~x483 & ~x663 & ~x702 & ~x741 & ~x780 & ~x819;
assign c4139 =  x10 &  x65 &  x87 &  x126 &  x659 &  x800 &  x911 & ~x252 & ~x369 & ~x705;
assign c4141 =  x131 &  x239 &  x494 &  x536 &  x546 &  x896 &  x1004 &  x1127 & ~x237 & ~x354 & ~x393 & ~x828;
assign c4143 =  x783 &  x864 &  x903 &  x1027;
assign c4145 =  x44 &  x56 &  x77 &  x80 &  x88 &  x127 &  x166 &  x188 &  x234 &  x269 &  x273 &  x371 &  x410 &  x431 &  x434 &  x551 &  x614 &  x662 &  x680 &  x749 &  x803 &  x839 &  x869 &  x875 &  x902 &  x953 &  x968 &  x998 &  x1019 &  x1034 &  x1055 &  x1073 &  x1094 &  x1118 & ~x624 & ~x663 & ~x702 & ~x741 & ~x780 & ~x783 & ~x819;
assign c4147 =  x751 & ~x351 & ~x393 & ~x876 & ~x990;
assign c4149 =  x10 &  x88 &  x188 &  x502 &  x544 &  x583 &  x607 &  x700 &  x727 &  x808 &  x892 &  x968;
assign c4151 =  x100 &  x317 &  x572 &  x605 &  x614 &  x653 &  x814 &  x866 &  x881 &  x892 &  x953 &  x998 &  x1025 &  x1034 & ~x354 & ~x393 & ~x432 & ~x471 & ~x831;
assign c4153 =  x104 &  x131 &  x155 &  x194 &  x224 &  x391 &  x659 &  x716 &  x839 &  x860 &  x1090 &  x1111 & ~x480 & ~x597 & ~x675 & ~x714;
assign c4155 =  x223 &  x534 & ~x909 & ~x987;
assign c4157 =  x2 &  x56 &  x83 &  x92 &  x137 &  x164 &  x178 &  x197 &  x233 &  x236 &  x242 &  x248 &  x263 &  x284 &  x302 &  x332 &  x416 &  x470 &  x494 &  x500 &  x518 &  x656 &  x664 &  x671 &  x686 &  x689 &  x716 &  x722 &  x734 &  x740 &  x755 &  x758 &  x803 &  x854 &  x878 &  x890 &  x926 &  x938 &  x959 &  x976 &  x986 &  x1015 &  x1043 &  x1046 &  x1124 & ~x648 & ~x675 & ~x687 & ~x753 & ~x792 & ~x831 & ~x870 & ~x909 & ~x948 & ~x987 & ~x1026;
assign c4159 =  x128 &  x583 &  x649 &  x688 &  x691 &  x727 &  x805 &  x854 &  x883 &  x1066 & ~x330 & ~x555 & ~x741;
assign c4161 =  x290 &  x536 &  x781 &  x841 & ~x393 & ~x954 & ~x990;
assign c4163 =  x91 &  x746 &  x791 &  x848 & ~x675 & ~x753 & ~x831 & ~x909;
assign c4165 =  x23 &  x71 &  x104 &  x137 &  x152 &  x167 &  x212 &  x308 &  x329 &  x359 &  x497 &  x587 &  x620 &  x656 &  x665 &  x671 &  x758 &  x787 &  x800 &  x812 &  x826 &  x830 &  x851 &  x893 &  x904 &  x908 &  x923 &  x929 &  x938 &  x943 &  x986 &  x989 &  x1004 &  x1022 &  x1025 &  x1027 &  x1031 &  x1066 &  x1073 & ~x600 & ~x639 & ~x756 & ~x858;
assign c4167 = ~x714 & ~x793 & ~x949;
assign c4169 =  x386 &  x713 &  x904 & ~x237 & ~x393 & ~x471 & ~x954;
assign c4171 =  x91 &  x169 &  x325 &  x386 &  x440 &  x452 &  x497 &  x683 &  x704 &  x775 &  x803 &  x814 &  x845 &  x929 &  x958 &  x1094 & ~x828 & ~x867;
assign c4173 =  x391 &  x962 & ~x442 & ~x636 & ~x780 & ~x819;
assign c4175 =  x52 &  x152 &  x620 &  x629 &  x791 & ~x432 & ~x433 & ~x510 & ~x771;
assign c4177 =  x101 &  x167 &  x257 &  x302 &  x503 &  x590 &  x629 &  x677 &  x731 &  x779 &  x794 &  x811 &  x845 &  x1027 &  x1066 &  x1091 &  x1094 & ~x600 & ~x639 & ~x756 & ~x780;
assign c4179 =  x391 &  x592 & ~x84 & ~x144 & ~x969 & ~x1125;
assign c4181 =  x329 &  x361 &  x400 & ~x36 & ~x561 & ~x639 & ~x702 & ~x936;
assign c4183 =  x335 &  x532 &  x596 &  x731 &  x764 &  x934 &  x1058 & ~x480 & ~x820 & ~x975;
assign c4185 =  x8 &  x41 &  x53 &  x65 &  x74 &  x149 &  x191 &  x224 &  x296 &  x332 &  x338 &  x356 &  x362 &  x440 &  x458 &  x511 &  x512 &  x532 &  x539 &  x572 &  x578 &  x649 &  x688 &  x707 &  x716 &  x743 &  x755 &  x767 &  x842 &  x860 &  x863 &  x877 &  x911 &  x935 &  x962 &  x1013 &  x1019 &  x1027 &  x1028 &  x1055 &  x1064 &  x1067 &  x1091 &  x1097 & ~x561 & ~x600 & ~x741 & ~x780 & ~x819;
assign c4187 =  x194 &  x822 &  x861 &  x979 &  x982 &  x1057 &  x1096;
assign c4189 =  x173 &  x398 &  x437 &  x593 &  x902 &  x1042 &  x1124 & ~x237 & ~x714 & ~x753 & ~x792 & ~x831 & ~x870 & ~x909 & ~x987 & ~x1026;
assign c4191 =  x778 &  x787 &  x817 &  x895 &  x934 &  x935 &  x1111 & ~x561 & ~x600 & ~x639;
assign c4193 =  x206 &  x688 &  x694 & ~x445 & ~x483 & ~x484;
assign c4195 =  x347 &  x362 &  x827 &  x920 &  x956 &  x980 & ~x81 & ~x237 & ~x570 & ~x648 & ~x687 & ~x720 & ~x828 & ~x867 & ~x906;
assign c4197 =  x556 &  x852 &  x930 &  x1014;
assign c4199 =  x83 &  x260 &  x518 &  x677 &  x783 &  x865 &  x904 &  x1025 & ~x87;
assign c4201 =  x751 & ~x835;
assign c4203 =  x532 &  x895 & ~x57 & ~x136 & ~x402;
assign c4205 =  x392 &  x536 &  x544 &  x583 &  x622 &  x661 &  x776 &  x779 &  x817 &  x856 &  x877 &  x895 &  x914 & ~x522 & ~x561 & ~x906 & ~x984;
assign c4207 =  x239 &  x392 &  x403 &  x404 &  x569 &  x989 &  x1015 & ~x687 & ~x831 & ~x909 & ~x1105;
assign c4209 =  x13 &  x130 &  x512 &  x1031 & ~x675 & ~x831 & ~x909 & ~x1065;
assign c4211 =  x77 &  x166 &  x205 &  x283 &  x322 &  x390 &  x429 &  x548 &  x1085 & ~x453 & ~x492;
assign c4213 = ~x636 & ~x675 & ~x754 & ~x871 & ~x910;
assign c4215 =  x155 &  x205 &  x272 &  x305 &  x353 &  x686 &  x725 &  x736 &  x808 &  x836 &  x880 &  x886 &  x932 &  x950 &  x1016 &  x1042 & ~x792;
assign c4217 =  x783 &  x822 &  x982 & ~x912;
assign c4221 =  x23 &  x65 &  x77 &  x80 &  x164 &  x191 &  x260 &  x389 &  x395 &  x431 &  x434 &  x449 &  x518 &  x587 &  x599 &  x617 &  x632 &  x644 &  x755 &  x860 &  x890 &  x895 &  x929 &  x934 &  x1040 & ~x3 & ~x81 & ~x159 & ~x354 & ~x432 & ~x471;
assign c4223 =  x460 & ~x471 & ~x792 & ~x871 & ~x1104;
assign c4225 =  x379 &  x419 &  x516 &  x555 &  x749 &  x1106 & ~x237;
assign c4227 =  x575 &  x1031 & ~x246 & ~x325 & ~x480 & ~x507 & ~x519 & ~x585 & ~x858 & ~x939;
assign c4229 =  x472 &  x850 &  x856 & ~x600 & ~x639 & ~x1101;
assign c4231 = ~x41;
assign c4233 =  x298 & ~x471 & ~x510 & ~x909 & ~x1027 & ~x1105;
assign c4235 =  x509 &  x578 &  x593 &  x839 &  x953 & ~x246 & ~x325 & ~x402 & ~x480 & ~x507 & ~x780 & ~x861;
assign c4237 =  x532 &  x605 &  x917 &  x955 &  x1070 & ~x402 & ~x702 & ~x703 & ~x742 & ~x780 & ~x781;
assign c4239 =  x609 & ~x976;
assign c4241 =  x477 &  x516 &  x585 & ~x354 & ~x591;
assign c4243 =  x232 &  x908 &  x1111 & ~x718;
assign c4245 =  x91 &  x607 &  x631 &  x684 &  x723 &  x801;
assign c4247 =  x32 &  x49 &  x340 &  x686 &  x779 &  x1112 & ~x354 & ~x393 & ~x792 & ~x948 & ~x1026 & ~x1065;
assign c4249 =  x80 &  x146 &  x149 &  x152 &  x248 &  x356 &  x377 &  x428 &  x490 &  x512 &  x607 &  x635 &  x646 &  x685 &  x701 &  x723 &  x790 &  x869 &  x884 &  x1037 &  x1121 & ~x144 & ~x183;
assign c4251 =  x632 &  x1121 & ~x510 & ~x832 & ~x871 & ~x1026 & ~x1065;
assign c4253 =  x10 &  x83 &  x88 &  x119 &  x196 &  x278 &  x353 &  x410 &  x413 &  x440 &  x500 &  x737 &  x788 &  x914 &  x1022 &  x1073 &  x1091 &  x1094 & ~x84 & ~x123 & ~x124 & ~x702 & ~x780;
assign c4255 =  x10 &  x322 & ~x18 & ~x369 & ~x990;
assign c4257 =  x476 &  x688 &  x727 &  x776 &  x1111 & ~x562;
assign c4259 =  x152 &  x462 &  x540 &  x751 &  x790 & ~x714;
assign c4261 =  x206 &  x322 & ~x123 & ~x714 & ~x792;
assign c4263 =  x10 &  x425 &  x428 &  x587 &  x680 &  x727 &  x782 &  x805 &  x850 &  x904 &  x943 &  x950 &  x982 &  x1066 & ~x84 & ~x123;
assign c4265 =  x10 &  x485 & ~x246 & ~x433;
assign c4267 =  x50 &  x77 &  x107 &  x125 &  x281 &  x311 &  x344 &  x350 &  x368 &  x449 &  x452 &  x476 &  x584 &  x586 &  x794 &  x845 &  x848 &  x863 &  x890 &  x902 &  x1003 &  x1040 &  x1042 &  x1112 & ~x237 & ~x714 & ~x792 & ~x798 & ~x837;
assign c4269 = ~x537 & ~x796;
assign c4271 =  x65 &  x127 &  x166 &  x173 &  x205 &  x244 &  x273 &  x482 &  x575 &  x620 &  x650 &  x908 &  x977 & ~x624 & ~x663 & ~x666 & ~x741 & ~x744 & ~x780 & ~x819 & ~x939;
assign c4273 =  x903 &  x1105;
assign c4275 =  x51 &  x1027 & ~x123 & ~x180 & ~x585;
assign c4277 =  x51 &  x736 &  x1039 & ~x633 & ~x975;
assign c4279 =  x388 &  x398 &  x427 &  x457 &  x529 &  x673 &  x712 &  x751 & ~x798;
assign c4281 =  x266 &  x269 &  x736 &  x764 &  x814 &  x956 & ~x714 & ~x792 & ~x871 & ~x948;
assign c4283 =  x221 &  x236 &  x238 &  x248 &  x283 &  x311 &  x391 &  x394 &  x422 &  x509 &  x605 &  x653 &  x662 &  x683 &  x713 &  x818 &  x866 &  x905 &  x962 &  x1004 &  x1070 & ~x366 & ~x405 & ~x406 & ~x483 & ~x522 & ~x702 & ~x780 & ~x819 & ~x900;
assign c4285 =  x233 &  x644 &  x692 &  x820 &  x1056 & ~x870 & ~x987 & ~x1107;
assign c4287 =  x331 &  x332 &  x451 &  x477 &  x841 & ~x537;
assign c4289 =  x110 &  x130 &  x169 &  x383 &  x686 &  x692 &  x899 &  x995 &  x1022 &  x1100 & ~x531 & ~x636 & ~x675 & ~x753 & ~x831;
assign c4291 =  x492 &  x844 &  x865 &  x943;
assign c4293 =  x278 &  x422 &  x553 &  x669 &  x755 &  x826 &  x833 &  x889 &  x926 &  x1028 &  x1067 &  x1112 & ~x483;
assign c4295 =  x544 & ~x325 & ~x756 & ~x780;
assign c4297 =  x86 &  x755 &  x783 &  x904 &  x982 &  x1018;
assign c4299 =  x1111 & ~x718 & ~x757 & ~x897;
assign c50 =  x2 &  x41 &  x71 &  x74 &  x77 &  x89 &  x107 &  x116 &  x176 &  x188 &  x263 &  x272 &  x281 &  x344 &  x389 &  x461 &  x500 &  x530 &  x563 &  x566 &  x638 &  x656 &  x680 &  x683 &  x686 &  x734 &  x746 &  x749 &  x781 &  x797 &  x833 &  x845 &  x893 &  x917 &  x923 &  x950 &  x1001 &  x1079 &  x1091 & ~x48 & ~x87 & ~x126 & ~x433 & ~x472 & ~x597 & ~x615 & ~x654 & ~x693 & ~x714 & ~x756 & ~x834;
assign c52 =  x32 &  x80 &  x155 &  x197 &  x323 &  x332 &  x338 &  x479 &  x530 &  x542 &  x584 &  x587 &  x632 &  x683 &  x688 &  x779 &  x785 &  x872 &  x971 &  x974 &  x1115 & ~x4 & ~x12 & ~x108 & ~x213 & ~x246 & ~x285 & ~x324;
assign c54 =  x86 &  x134 &  x239 &  x245 &  x281 &  x287 &  x314 &  x353 &  x389 &  x404 &  x446 &  x536 &  x587 &  x599 &  x623 &  x644 &  x662 &  x704 &  x761 &  x788 &  x854 &  x890 &  x896 &  x911 &  x916 &  x926 &  x944 &  x959 &  x994 &  x1004 &  x1034 &  x1076 & ~x12 & ~x42 & ~x43 & ~x82 & ~x91 & ~x129 & ~x246;
assign c56 =  x1 &  x40 &  x44 &  x47 &  x68 &  x155 &  x157 &  x266 &  x335 &  x389 &  x461 &  x503 &  x641 &  x650 &  x665 &  x671 &  x692 &  x734 &  x752 &  x821 &  x872 &  x908 &  x917 &  x1007 &  x1016 &  x1115 & ~x4 & ~x213 & ~x324 & ~x363;
assign c58 =  x8 &  x11 &  x23 &  x32 &  x47 &  x59 &  x92 &  x98 &  x101 &  x152 &  x155 &  x158 &  x161 &  x167 &  x182 &  x212 &  x221 &  x224 &  x230 &  x233 &  x245 &  x248 &  x257 &  x266 &  x323 &  x353 &  x383 &  x386 &  x392 &  x410 &  x449 &  x455 &  x467 &  x485 &  x494 &  x497 &  x503 &  x506 &  x515 &  x521 &  x523 &  x542 &  x551 &  x563 &  x569 &  x572 &  x574 &  x587 &  x590 &  x593 &  x599 &  x632 &  x635 &  x641 &  x703 &  x719 &  x725 &  x742 &  x752 &  x764 &  x791 &  x797 &  x803 &  x809 &  x815 &  x836 &  x845 &  x851 &  x859 &  x866 &  x881 &  x887 &  x896 &  x911 &  x947 &  x968 &  x974 &  x980 &  x992 &  x1001 &  x1016 &  x1028 &  x1037 &  x1043 &  x1052 &  x1055 &  x1057 &  x1058 &  x1067 &  x1073 &  x1076 &  x1079 &  x1082 &  x1112 &  x1115 &  x1121 &  x1127 & ~x432 & ~x433 & ~x472 & ~x511 & ~x621 & ~x675 & ~x714 & ~x831;
assign c510 =  x14 &  x32 &  x128 &  x170 &  x191 &  x194 &  x218 &  x239 &  x251 &  x280 &  x320 &  x332 &  x362 &  x368 &  x377 &  x395 &  x397 &  x445 &  x452 &  x475 &  x484 &  x514 &  x523 &  x557 &  x562 &  x599 &  x617 &  x632 &  x671 &  x674 &  x815 &  x869 &  x923 &  x932 &  x998 &  x1018 &  x1022 &  x1025 &  x1031 &  x1054 &  x1055 &  x1070 &  x1091 &  x1124 & ~x237 & ~x525 & ~x714 & ~x753 & ~x792 & ~x831 & ~x870 & ~x909 & ~x948 & ~x987 & ~x1026;
assign c512 =  x8 &  x14 &  x38 &  x77 &  x80 &  x101 &  x152 &  x164 &  x167 &  x206 &  x212 &  x239 &  x298 &  x347 &  x350 &  x380 &  x397 &  x475 &  x513 &  x514 &  x518 &  x552 &  x554 &  x592 &  x602 &  x613 &  x631 &  x632 &  x635 &  x647 &  x683 &  x731 &  x743 &  x746 &  x788 &  x794 &  x809 &  x842 &  x869 &  x875 &  x974 &  x1057 &  x1064 &  x1070 &  x1082 &  x1094 & ~x777 & ~x816 & ~x876;
assign c514 =  x53 &  x59 &  x98 &  x116 &  x179 &  x202 &  x344 &  x353 &  x365 &  x413 &  x467 &  x575 &  x584 &  x593 &  x677 &  x680 &  x704 &  x713 &  x761 &  x773 &  x863 &  x869 &  x890 &  x902 &  x1019 &  x1097 & ~x108 & ~x207 & ~x246 & ~x489 & ~x501 & ~x561 & ~x600 & ~x663 & ~x852 & ~x1029;
assign c516 =  x5 &  x8 &  x14 &  x32 &  x44 &  x50 &  x53 &  x77 &  x113 &  x122 &  x134 &  x140 &  x143 &  x155 &  x176 &  x200 &  x206 &  x230 &  x245 &  x275 &  x284 &  x287 &  x299 &  x305 &  x317 &  x332 &  x344 &  x353 &  x359 &  x368 &  x374 &  x380 &  x383 &  x389 &  x407 &  x416 &  x428 &  x434 &  x461 &  x476 &  x479 &  x485 &  x488 &  x524 &  x527 &  x551 &  x563 &  x566 &  x575 &  x584 &  x587 &  x593 &  x596 &  x599 &  x602 &  x614 &  x620 &  x629 &  x668 &  x671 &  x674 &  x680 &  x695 &  x710 &  x734 &  x737 &  x743 &  x770 &  x785 &  x791 &  x797 &  x800 &  x815 &  x824 &  x827 &  x833 &  x836 &  x845 &  x866 &  x893 &  x908 &  x920 &  x926 &  x929 &  x935 &  x941 &  x950 &  x974 &  x983 &  x989 &  x1001 &  x1019 &  x1034 &  x1040 &  x1043 &  x1049 &  x1064 &  x1085 &  x1088 &  x1097 &  x1103 &  x1112 & ~x160 & ~x237 & ~x324 & ~x363 & ~x603 & ~x678 & ~x696 & ~x717 & ~x735 & ~x756 & ~x774 & ~x789;
assign c518 =  x50 &  x56 &  x77 &  x95 &  x119 &  x164 &  x182 &  x266 &  x278 &  x290 &  x296 &  x311 &  x356 &  x359 &  x377 &  x404 &  x446 &  x461 &  x467 &  x527 &  x530 &  x536 &  x539 &  x599 &  x617 &  x623 &  x632 &  x644 &  x653 &  x704 &  x707 &  x752 &  x758 &  x809 &  x824 &  x899 &  x923 &  x1004 &  x1028 &  x1076 &  x1094 & ~x198 & ~x199 & ~x207 & ~x238 & ~x246 & ~x324 & ~x363 & ~x364 & ~x402 & ~x480 & ~x519 & ~x1029 & ~x1092;
assign c520 =  x29 &  x68 &  x172 &  x182 &  x209 &  x227 &  x233 &  x418 &  x514 &  x523 &  x562 &  x602 &  x646 &  x647 &  x652 &  x685 &  x724 &  x780 &  x892 &  x931 &  x953 &  x1010 &  x1018 &  x1057;
assign c522 =  x17 &  x38 &  x50 &  x53 &  x68 &  x74 &  x77 &  x80 &  x113 &  x140 &  x161 &  x176 &  x218 &  x239 &  x242 &  x287 &  x290 &  x305 &  x398 &  x407 &  x425 &  x446 &  x455 &  x458 &  x464 &  x473 &  x485 &  x494 &  x503 &  x509 &  x530 &  x542 &  x551 &  x557 &  x563 &  x575 &  x611 &  x641 &  x653 &  x656 &  x686 &  x689 &  x695 &  x704 &  x746 &  x773 &  x812 &  x823 &  x854 &  x878 &  x881 &  x900 &  x914 &  x977 &  x980 &  x986 &  x1013 &  x1046 &  x1049 &  x1052 &  x1058 &  x1112 &  x1115 &  x1127 &  x1130 & ~x234 & ~x273 & ~x550 & ~x621 & ~x714 & ~x831 & ~x874 & ~x951 & ~x952 & ~x1029;
assign c524 =  x34 &  x379 &  x568 &  x661 &  x817 &  x841 &  x898 &  x934 &  x969 &  x1051 &  x1075;
assign c526 =  x20 &  x167 &  x233 &  x290 &  x329 &  x341 &  x374 &  x410 &  x419 &  x473 &  x485 &  x488 &  x554 &  x599 &  x617 &  x656 &  x740 &  x746 &  x782 &  x785 &  x800 &  x1018 &  x1046 & ~x199 & ~x237 & ~x238 & ~x297 & ~x483 & ~x561 & ~x600 & ~x789;
assign c528 =  x32 &  x131 &  x176 &  x182 &  x227 &  x263 &  x269 &  x302 &  x350 &  x416 &  x464 &  x545 &  x571 &  x583 &  x610 &  x649 &  x668 &  x683 &  x707 &  x715 &  x754 &  x832 &  x842 &  x845 &  x871 &  x887 &  x944 &  x989 &  x1016 &  x1028 &  x1109 & ~x42 & ~x174 & ~x213 & ~x219 & ~x252;
assign c530 =  x125 &  x257 &  x293 &  x548 &  x704 & ~x82 & ~x121 & ~x160 & ~x199 & ~x246 & ~x285 & ~x324 & ~x325 & ~x364 & ~x441 & ~x600;
assign c532 =  x11 &  x26 &  x35 &  x62 &  x74 &  x98 &  x104 &  x110 &  x118 &  x146 &  x167 &  x206 &  x239 &  x251 &  x275 &  x281 &  x305 &  x312 &  x314 &  x317 &  x389 &  x407 &  x443 &  x458 &  x461 &  x476 &  x488 &  x506 &  x512 &  x527 &  x539 &  x545 &  x548 &  x563 &  x575 &  x578 &  x584 &  x587 &  x593 &  x611 &  x665 &  x680 &  x704 &  x722 &  x773 &  x791 &  x800 &  x806 &  x833 &  x848 &  x851 &  x902 &  x929 &  x965 &  x983 &  x998 &  x1004 &  x1010 &  x1028 &  x1034 &  x1049 &  x1052 &  x1103 &  x1106 & ~x81 & ~x82 & ~x121 & ~x207 & ~x633 & ~x819;
assign c534 =  x11 &  x14 &  x20 &  x32 &  x44 &  x47 &  x59 &  x62 &  x71 &  x80 &  x89 &  x95 &  x110 &  x125 &  x134 &  x137 &  x155 &  x157 &  x170 &  x179 &  x191 &  x200 &  x227 &  x230 &  x239 &  x257 &  x263 &  x281 &  x290 &  x305 &  x323 &  x326 &  x329 &  x347 &  x350 &  x356 &  x359 &  x374 &  x383 &  x416 &  x449 &  x482 &  x509 &  x524 &  x584 &  x608 &  x611 &  x632 &  x659 &  x692 &  x710 &  x722 &  x734 &  x740 &  x746 &  x749 &  x752 &  x755 &  x773 &  x776 &  x788 &  x833 &  x842 &  x854 &  x857 &  x863 &  x881 &  x905 &  x916 &  x923 &  x959 &  x962 &  x968 &  x974 &  x994 &  x1004 &  x1019 &  x1033 &  x1040 &  x1049 &  x1055 &  x1082 &  x1091 &  x1112 & ~x82 & ~x180 & ~x231 & ~x246 & ~x270 & ~x444;
assign c536 =  x47 &  x191 &  x224 &  x365 &  x395 &  x418 &  x422 &  x457 &  x475 &  x503 &  x514 &  x553 &  x560 &  x592 &  x671 &  x677 &  x695 &  x725 &  x737 &  x779 &  x839 &  x878 &  x962 &  x968 &  x1043 &  x1049 & ~x87 & ~x165 & ~x558 & ~x864 & ~x903 & ~x1029;
assign c538 =  x5 &  x8 &  x23 &  x26 &  x41 &  x47 &  x53 &  x59 &  x65 &  x77 &  x98 &  x128 &  x137 &  x142 &  x152 &  x167 &  x170 &  x188 &  x191 &  x194 &  x206 &  x209 &  x212 &  x218 &  x221 &  x230 &  x233 &  x236 &  x254 &  x259 &  x269 &  x284 &  x287 &  x290 &  x296 &  x298 &  x302 &  x308 &  x323 &  x326 &  x329 &  x350 &  x356 &  x367 &  x371 &  x373 &  x376 &  x398 &  x422 &  x436 &  x443 &  x449 &  x452 &  x455 &  x458 &  x467 &  x475 &  x476 &  x485 &  x488 &  x490 &  x494 &  x514 &  x518 &  x521 &  x536 &  x560 &  x563 &  x566 &  x568 &  x587 &  x593 &  x596 &  x607 &  x611 &  x629 &  x646 &  x647 &  x650 &  x653 &  x659 &  x677 &  x680 &  x683 &  x692 &  x698 &  x704 &  x710 &  x713 &  x716 &  x725 &  x743 &  x749 &  x752 &  x782 &  x785 &  x791 &  x800 &  x803 &  x812 &  x815 &  x824 &  x827 &  x842 &  x857 &  x860 &  x863 &  x866 &  x875 &  x878 &  x886 &  x890 &  x893 &  x905 &  x917 &  x920 &  x932 &  x934 &  x935 &  x938 &  x940 &  x947 &  x950 &  x962 &  x964 &  x971 &  x980 &  x983 &  x992 &  x995 &  x1001 &  x1010 &  x1019 &  x1028 &  x1031 &  x1037 &  x1043 &  x1049 &  x1055 &  x1067 &  x1082 &  x1112 &  x1121 &  x1130 & ~x393 & ~x432 & ~x471;
assign c540 =  x20 &  x50 &  x80 &  x125 &  x143 &  x152 &  x158 &  x164 &  x209 &  x215 &  x236 &  x329 &  x359 &  x371 &  x374 &  x392 &  x419 &  x425 &  x446 &  x455 &  x461 &  x467 &  x473 &  x476 &  x515 &  x545 &  x572 &  x575 &  x581 &  x584 &  x587 &  x593 &  x611 &  x620 &  x632 &  x647 &  x656 &  x668 &  x698 &  x713 &  x719 &  x746 &  x767 &  x791 &  x800 &  x824 &  x827 &  x830 &  x836 &  x839 &  x845 &  x858 &  x859 &  x872 &  x875 &  x890 &  x897 &  x902 &  x917 &  x944 &  x950 &  x962 &  x1017 &  x1025 &  x1031 &  x1049 &  x1055 &  x1061 &  x1064 &  x1079 &  x1085 &  x1096 & ~x432 & ~x589 & ~x628 & ~x714 & ~x792 & ~x831 & ~x870 & ~x909 & ~x948 & ~x1029;
assign c542 =  x10 &  x16 &  x22 &  x61 &  x178 &  x257 &  x260 &  x295 &  x334 &  x353 &  x373 &  x412 &  x490 &  x505 &  x568 &  x584 &  x593 &  x622 &  x638 &  x677 &  x731 &  x773 &  x880 &  x886 &  x914 &  x919 &  x1018 &  x1036 &  x1081 &  x1120 & ~x558;
assign c544 =  x19 &  x20 &  x97 &  x161 &  x163 &  x202 &  x260 &  x263 &  x266 &  x368 &  x383 &  x397 &  x422 &  x476 &  x542 &  x547 &  x551 &  x854 &  x878 &  x895 &  x1033 & ~x198 & ~x678;
assign c546 =  x8 &  x83 &  x119 &  x134 &  x140 &  x143 &  x191 &  x230 &  x242 &  x254 &  x319 &  x329 &  x332 &  x358 &  x380 &  x383 &  x389 &  x398 &  x446 &  x458 &  x461 &  x475 &  x476 &  x491 &  x506 &  x509 &  x515 &  x523 &  x545 &  x566 &  x578 &  x611 &  x614 &  x629 &  x659 &  x689 &  x692 &  x728 &  x800 &  x857 &  x860 &  x872 &  x875 &  x887 &  x893 &  x901 &  x934 &  x965 &  x968 &  x1001 &  x1013 &  x1025 &  x1040 &  x1091 &  x1118 &  x1124 & ~x432 & ~x433 & ~x471 & ~x537 & ~x576 & ~x615 & ~x636 & ~x654 & ~x675 & ~x693 & ~x714 & ~x870;
assign c548 =  x302 &  x404 &  x431 &  x593 &  x608 &  x713 &  x759 &  x791 &  x872 &  x905 &  x1033 &  x1112 &  x1121 & ~x192 & ~x207 & ~x231 & ~x246 & ~x1041;
assign c550 =  x65 &  x68 &  x134 &  x155 &  x188 &  x206 &  x239 &  x272 &  x296 &  x332 &  x338 &  x359 &  x506 &  x514 &  x518 &  x553 &  x575 &  x641 &  x689 &  x800 &  x819 &  x836 &  x878 &  x917 &  x940 &  x950 &  x968 &  x986 &  x1007 &  x1018 &  x1052 &  x1057 &  x1079 &  x1096 &  x1121 & ~x550 & ~x589 & ~x660 & ~x714 & ~x870 & ~x909;
assign c552 =  x29 &  x32 &  x77 &  x80 &  x167 &  x176 &  x185 &  x200 &  x209 &  x233 &  x235 &  x245 &  x260 &  x263 &  x296 &  x305 &  x377 &  x395 &  x428 &  x467 &  x548 &  x698 &  x704 &  x716 &  x725 &  x737 &  x740 &  x755 &  x794 &  x809 &  x815 &  x827 &  x842 &  x866 &  x869 &  x875 &  x950 &  x974 &  x1001 &  x1013 &  x1022 &  x1079 &  x1103 &  x1112 & ~x42 & ~x82 & ~x180 & ~x213 & ~x219 & ~x252 & ~x258 & ~x291 & ~x292 & ~x324 & ~x331 & ~x363 & ~x369 & ~x370;
assign c554 =  x386 &  x530 &  x794 &  x978 & ~x549 & ~x550 & ~x589 & ~x714 & ~x870 & ~x913 & ~x952;
assign c556 =  x53 &  x194 &  x302 &  x338 &  x383 &  x392 &  x395 &  x446 &  x515 &  x566 &  x800 &  x872 &  x910 &  x949 &  x994 &  x1027 &  x1066 & ~x12 & ~x51 & ~x52 & ~x91 & ~x129 & ~x168 & ~x207 & ~x246 & ~x405;
assign c558 =  x35 &  x77 &  x125 &  x176 &  x211 &  x245 &  x250 &  x263 &  x311 &  x446 &  x452 &  x547 &  x593 &  x649 &  x755 &  x761 &  x766 &  x923 &  x992 &  x1025 &  x1097 &  x1127 & ~x199 & ~x238 & ~x277 & ~x420 & ~x441 & ~x480 & ~x519 & ~x600;
assign c560 =  x8 &  x83 &  x158 &  x188 &  x227 &  x239 &  x251 &  x278 &  x302 &  x305 &  x332 &  x353 &  x389 &  x398 &  x410 &  x482 &  x506 &  x509 &  x550 &  x554 &  x563 &  x572 &  x575 &  x587 &  x602 &  x605 &  x610 &  x629 &  x632 &  x656 &  x661 &  x688 &  x695 &  x700 &  x704 &  x707 &  x725 &  x773 &  x785 &  x812 &  x857 &  x920 &  x968 &  x971 &  x986 &  x988 &  x1031 &  x1033 &  x1039 &  x1040 &  x1066 &  x1070 &  x1088 &  x1117 & ~x519 & ~x600 & ~x750 & ~x789;
assign c562 =  x23 &  x47 &  x77 &  x80 &  x83 &  x86 &  x89 &  x131 &  x176 &  x188 &  x194 &  x200 &  x272 &  x275 &  x326 &  x392 &  x401 &  x406 &  x422 &  x431 &  x443 &  x445 &  x449 &  x455 &  x484 &  x497 &  x509 &  x521 &  x523 &  x536 &  x551 &  x566 &  x578 &  x605 &  x611 &  x638 &  x644 &  x668 &  x683 &  x701 &  x707 &  x716 &  x725 &  x740 &  x742 &  x761 &  x764 &  x791 &  x797 &  x821 &  x869 &  x884 &  x893 &  x935 &  x940 &  x947 &  x971 &  x983 &  x992 &  x998 &  x1004 &  x1016 &  x1061 &  x1073 &  x1109 &  x1124 &  x1127 & ~x472 & ~x576 & ~x615 & ~x654 & ~x675 & ~x693 & ~x756 & ~x796 & ~x834;
assign c564 =  x110 &  x167 &  x239 &  x245 &  x326 &  x344 &  x356 &  x431 &  x490 &  x562 &  x568 &  x574 &  x599 &  x601 &  x607 &  x671 &  x710 &  x724 &  x743 &  x809 &  x830 &  x858 &  x898 &  x899 &  x1014 &  x1061 & ~x714 & ~x831 & ~x909 & ~x910 & ~x988;
assign c566 =  x17 &  x275 &  x395 &  x467 &  x470 &  x488 &  x527 &  x766 &  x905 &  x994 &  x1010 &  x1033 &  x1066 &  x1078 &  x1117 & ~x246 & ~x285 & ~x324 & ~x519 & ~x525 & ~x558 & ~x750 & ~x789 & ~x828 & ~x867 & ~x906;
assign c568 =  x16 &  x35 &  x40 &  x61 &  x62 &  x85 &  x164 &  x178 &  x200 &  x260 &  x380 &  x398 &  x457 &  x467 &  x491 &  x557 &  x583 &  x584 &  x701 &  x719 &  x758 &  x769 &  x782 &  x788 &  x791 &  x808 &  x817 &  x821 &  x824 &  x826 &  x827 &  x880 &  x934 &  x1055 &  x1106;
assign c570 =  x547 &  x588 &  x627 & ~x277 & ~x316 & ~x525 & ~x600 & ~x603 & ~x642;
assign c572 =  x2 &  x95 &  x182 &  x254 &  x317 &  x350 &  x473 &  x484 &  x506 &  x523 &  x530 &  x542 &  x562 &  x568 &  x600 &  x607 &  x716 &  x758 &  x773 &  x780 &  x794 &  x820 &  x859 &  x881 &  x940 &  x1019 &  x1076 &  x1088 &  x1103 & ~x354 & ~x432 & ~x550 & ~x589 & ~x693 & ~x714 & ~x831;
assign c574 =  x98 &  x146 &  x155 &  x206 &  x422 &  x587 &  x665 &  x749 &  x878 &  x890 & ~x324 & ~x639 & ~x679 & ~x718 & ~x835 & ~x874 & ~x913 & ~x930 & ~x951 & ~x990 & ~x1029 & ~x1125;
assign c576 =  x179 &  x224 &  x248 &  x410 &  x491 &  x691 &  x859 &  x1052 &  x1056 &  x1095 & ~x399 & ~x982;
assign c578 =  x40 &  x61 &  x80 &  x148 &  x178 &  x239 &  x373 &  x392 &  x412 &  x457 &  x460 &  x490 &  x515 &  x523 &  x596 &  x607 &  x698 &  x815 &  x842 &  x853 &  x899 &  x1076 & ~x393 & ~x714 & ~x753 & ~x831 & ~x870 & ~x909;
assign c580 =  x37 &  x152 &  x202 &  x263 &  x607 &  x622 &  x646 &  x649 &  x655 &  x754 &  x934 &  x938 &  x944 &  x983 &  x1007 & ~x672;
assign c582 =  x11 &  x50 &  x65 &  x74 &  x95 &  x98 &  x101 &  x116 &  x137 &  x146 &  x152 &  x179 &  x191 &  x218 &  x278 &  x302 &  x314 &  x338 &  x341 &  x353 &  x356 &  x365 &  x368 &  x377 &  x386 &  x431 &  x452 &  x455 &  x469 &  x482 &  x491 &  x509 &  x533 &  x547 &  x554 &  x581 &  x602 &  x608 &  x614 &  x620 &  x623 &  x629 &  x644 &  x647 &  x662 &  x668 &  x671 &  x677 &  x710 &  x722 &  x728 &  x737 &  x743 &  x761 &  x770 &  x784 &  x815 &  x833 &  x863 &  x872 &  x878 &  x881 &  x895 &  x911 &  x914 &  x923 &  x934 &  x947 &  x950 &  x965 &  x971 &  x977 &  x986 &  x1025 &  x1028 &  x1031 &  x1067 &  x1076 &  x1118 &  x1121 &  x1124 &  x1127 &  x1130 & ~x277 & ~x316 & ~x336 & ~x355 & ~x393 & ~x678;
assign c584 =  x61 &  x211 &  x334 &  x373 &  x460 &  x562 &  x646 &  x724 &  x853 &  x892 & ~x621 & ~x699 & ~x714 & ~x831 & ~x909;
assign c586 =  x26 &  x152 &  x206 &  x341 &  x347 &  x418 &  x431 &  x479 &  x494 &  x508 &  x509 &  x625 &  x638 &  x665 &  x744 &  x761 &  x959 &  x1079 & ~x355 & ~x394 & ~x678 & ~x681 & ~x759 & ~x795;
assign c588 =  x23 &  x34 &  x47 &  x77 &  x100 &  x110 &  x137 &  x146 &  x229 &  x256 &  x267 &  x295 &  x306 &  x307 &  x334 &  x380 &  x395 &  x407 &  x419 &  x422 &  x545 &  x548 &  x554 &  x599 &  x632 &  x649 &  x655 &  x692 &  x694 &  x772 &  x815 &  x821 &  x845 &  x887 &  x914 &  x935 &  x956 &  x959 &  x962 &  x1036 &  x1052 &  x1057 &  x1070 &  x1075 &  x1091 &  x1096 &  x1120 &  x1130;
assign c590 =  x157 &  x184 &  x202 &  x535 &  x568 &  x574 &  x607 &  x646 &  x652 &  x655 &  x694 &  x724 &  x763 &  x802 &  x880 &  x892 &  x1036;
assign c592 =  x11 &  x74 &  x134 &  x185 &  x212 &  x254 &  x257 &  x266 &  x362 &  x395 &  x482 &  x484 &  x512 &  x514 &  x553 &  x562 &  x566 &  x572 &  x581 &  x599 &  x611 &  x674 &  x770 &  x782 &  x819 &  x848 &  x858 &  x897 &  x941 &  x1019 &  x1054 & ~x273 & ~x315 & ~x589 & ~x627 & ~x714 & ~x870 & ~x909 & ~x910 & ~x987;
assign c594 =  x20 &  x71 &  x86 &  x179 &  x203 &  x215 &  x227 &  x320 &  x323 &  x359 &  x389 &  x419 &  x449 &  x458 &  x539 &  x578 &  x613 &  x644 &  x652 &  x701 &  x716 &  x719 &  x776 &  x788 &  x878 &  x975 &  x977 &  x986 &  x1056 &  x1057 &  x1076 &  x1093 &  x1095 &  x1096 &  x1127 &  x1130 & ~x667 & ~x987 & ~x1026 & ~x1029;
assign c596 =  x10 &  x34 &  x229 &  x383 &  x412 &  x451 &  x490 &  x622 &  x657 &  x691 &  x743 &  x769 &  x814 &  x853 &  x892 &  x1120;
assign c598 =  x95 &  x104 &  x197 &  x215 &  x239 &  x280 &  x326 &  x475 &  x553 &  x607 &  x815 &  x818 &  x897 &  x1004 &  x1018 &  x1057 & ~x312 & ~x589 & ~x621 & ~x699 & ~x738;
assign c5100 =  x11 &  x14 &  x32 &  x56 &  x59 &  x80 &  x83 &  x107 &  x116 &  x137 &  x140 &  x146 &  x152 &  x161 &  x167 &  x170 &  x182 &  x188 &  x194 &  x206 &  x212 &  x242 &  x245 &  x248 &  x254 &  x275 &  x284 &  x293 &  x296 &  x332 &  x335 &  x344 &  x353 &  x359 &  x386 &  x389 &  x395 &  x404 &  x410 &  x416 &  x434 &  x461 &  x476 &  x485 &  x488 &  x494 &  x508 &  x512 &  x518 &  x521 &  x530 &  x533 &  x548 &  x560 &  x569 &  x587 &  x590 &  x602 &  x605 &  x620 &  x629 &  x635 &  x644 &  x662 &  x665 &  x680 &  x689 &  x692 &  x698 &  x704 &  x710 &  x722 &  x725 &  x740 &  x764 &  x770 &  x782 &  x785 &  x794 &  x797 &  x806 &  x812 &  x818 &  x824 &  x851 &  x869 &  x890 &  x893 &  x905 &  x914 &  x923 &  x938 &  x944 &  x947 &  x950 &  x977 &  x983 &  x986 &  x989 &  x995 &  x998 &  x1004 &  x1007 &  x1022 &  x1031 &  x1040 &  x1043 &  x1049 &  x1064 &  x1082 &  x1088 &  x1097 &  x1118 & ~x237 & ~x277 & ~x309 & ~x315 & ~x316 & ~x348 & ~x349 & ~x354 & ~x388 & ~x426 & ~x427 & ~x465 & ~x486 & ~x525 & ~x564;
assign c5102 =  x56 &  x425 &  x483 &  x484 &  x522 &  x562 &  x940 & ~x550 & ~x714 & ~x831 & ~x912 & ~x951 & ~x952;
assign c5104 =  x32 &  x40 &  x47 &  x110 &  x118 &  x157 &  x196 &  x215 &  x274 &  x383 &  x452 &  x479 &  x571 &  x583 &  x610 &  x649 &  x668 &  x688 &  x764 &  x779 &  x815 &  x869 &  x872 &  x928 &  x977 &  x1040 &  x1043 &  x1049 &  x1064 & ~x42 & ~x405 & ~x585 & ~x624 & ~x663 & ~x780 & ~x897;
assign c5106 =  x83 &  x101 &  x182 &  x329 &  x362 &  x395 &  x476 &  x488 &  x503 &  x536 &  x566 &  x659 &  x731 &  x895 &  x929 &  x935 &  x940 &  x941 &  x980 &  x1004 &  x1094 &  x1115 & ~x480 & ~x558 & ~x675 & ~x714 & ~x720 & ~x834 & ~x837 & ~x874 & ~x912 & ~x913 & ~x951 & ~x1107;
assign c5108 =  x332 &  x503 &  x773 &  x830 &  x1028 & ~x400 & ~x438 & ~x672 & ~x831 & ~x832 & ~x903 & ~x909 & ~x942;
assign c5110 =  x176 &  x383 &  x476 &  x524 &  x743 &  x947 &  x1016 &  x1121 & ~x81 & ~x82 & ~x121 & ~x246 & ~x252 & ~x285 & ~x291 & ~x292 & ~x324 & ~x370 & ~x447 & ~x639;
assign c5112 =  x475 &  x514 &  x523 &  x901 & ~x433 & ~x511 & ~x525 & ~x714 & ~x792 & ~x831 & ~x834;
assign c5114 =  x29 &  x40 &  x155 &  x157 &  x182 &  x245 &  x278 &  x296 &  x341 &  x352 &  x391 &  x432 &  x455 &  x506 &  x542 &  x566 &  x575 &  x620 &  x656 &  x794 &  x833 &  x863 &  x878 &  x896 &  x935 &  x968 &  x986 &  x989 &  x1004 &  x1109 &  x1127 & ~x180 & ~x207 & ~x444 & ~x600 & ~x672;
assign c5116 =  x44 &  x47 &  x110 &  x149 &  x263 &  x293 &  x299 &  x302 &  x326 &  x329 &  x338 &  x386 &  x452 &  x467 &  x514 &  x515 &  x523 &  x553 &  x562 &  x572 &  x584 &  x592 &  x601 &  x605 &  x623 &  x632 &  x674 &  x701 &  x704 &  x824 &  x878 &  x898 &  x917 &  x962 &  x1007 &  x1096 & ~x792 & ~x831 & ~x912 & ~x913 & ~x951 & ~x952;
assign c5118 =  x17 &  x32 &  x89 &  x188 &  x257 &  x323 &  x389 &  x450 &  x451 &  x479 &  x490 &  x563 &  x568 &  x577 &  x581 &  x616 &  x655 &  x662 &  x671 &  x698 &  x719 &  x725 &  x761 &  x769 &  x797 &  x808 &  x962 &  x974 &  x986 &  x1022 &  x1040 &  x1055 &  x1070 & ~x633 & ~x789 & ~x828;
assign c5120 =  x14 &  x47 &  x77 &  x86 &  x104 &  x119 &  x128 &  x155 &  x236 &  x248 &  x263 &  x296 &  x314 &  x332 &  x443 &  x488 &  x491 &  x566 &  x578 &  x641 &  x644 &  x650 &  x707 &  x773 &  x809 &  x854 &  x863 &  x872 &  x881 &  x920 &  x926 &  x947 &  x965 &  x989 &  x1028 &  x1058 &  x1088 &  x1121 & ~x160 & ~x199 & ~x237 & ~x285 & ~x324 & ~x363 & ~x402 & ~x564 & ~x678 & ~x681 & ~x696 & ~x717 & ~x720 & ~x735 & ~x774;
assign c5122 = ~x4 & ~x129 & ~x169 & ~x208 & ~x213 & ~x246 & ~x285 & ~x324 & ~x813;
assign c5124 =  x19 &  x158 &  x211 &  x288 &  x585 &  x812 & ~x597 & ~x714;
assign c5126 =  x19 &  x29 &  x143 &  x341 &  x407 &  x428 &  x515 &  x530 &  x817 &  x869 &  x917 &  x1040 &  x1106 & ~x237 & ~x316 & ~x519 & ~x525 & ~x558 & ~x564 & ~x597 & ~x603 & ~x678;
assign c5128 =  x35 &  x71 &  x110 &  x137 &  x146 &  x182 &  x280 &  x284 &  x299 &  x329 &  x332 &  x384 &  x440 &  x491 &  x686 &  x725 &  x782 &  x791 &  x884 &  x896 &  x1019 &  x1049 &  x1067 &  x1079 &  x1097 &  x1130 & ~x276 & ~x486 & ~x525 & ~x603 & ~x642 & ~x681 & ~x714 & ~x753 & ~x837;
assign c5130 =  x53 &  x68 &  x157 &  x272 &  x432 &  x471 &  x533 &  x569 &  x593 &  x755 &  x797 &  x914 &  x968 &  x1037 & ~x180 & ~x367 & ~x406 & ~x445 & ~x523 & ~x633;
assign c5132 =  x150 &  x195 &  x383 &  x700 &  x958 &  x986 &  x994 &  x1120 &  x1126;
assign c5134 =  x155 & ~x199 & ~x238 & ~x246 & ~x285 & ~x324 & ~x403 & ~x442 & ~x480 & ~x519 & ~x717;
assign c5136 =  x8 &  x50 &  x224 &  x533 &  x542 &  x610 &  x803 &  x917 & ~x43 & ~x174 & ~x186 & ~x213 & ~x214 & ~x246 & ~x252 & ~x253 & ~x292 & ~x324;
assign c5138 =  x170 &  x185 &  x217 &  x332 &  x341 &  x368 &  x398 &  x497 &  x610 &  x644 &  x649 &  x764 &  x766 &  x815 &  x842 &  x884 &  x934 &  x944 & ~x96 & ~x213 & ~x214 & ~x252 & ~x253 & ~x324;
assign c5140 =  x173 &  x503 & ~x108 & ~x213 & ~x324 & ~x327 & ~x639 & ~x852 & ~x858 & ~x891 & ~x930 & ~x969 & ~x1035 & ~x1047 & ~x1074 & ~x1086 & ~x1107 & ~x1125;
assign c5142 =  x116 &  x158 &  x206 &  x319 &  x380 &  x623 &  x649 &  x656 &  x688 &  x727 &  x731 &  x766 &  x811 &  x1070 & ~x252 & ~x291 & ~x292 & ~x447 & ~x486 & ~x525 & ~x597;
assign c5144 =  x136 &  x392 &  x781 &  x809 &  x901 &  x1057 &  x1096 & ~x394 & ~x433 & ~x472 & ~x558 & ~x714 & ~x753 & ~x792 & ~x831;
assign c5146 =  x5 &  x11 &  x26 &  x35 &  x104 &  x134 &  x203 &  x290 &  x404 &  x416 &  x419 &  x446 &  x500 &  x572 &  x617 &  x632 &  x647 &  x656 &  x686 &  x695 &  x761 &  x782 &  x881 &  x926 &  x938 &  x1064 &  x1121 & ~x87 & ~x165 & ~x166 & ~x205 & ~x243 & ~x244 & ~x324 & ~x438 & ~x555 & ~x672 & ~x711 & ~x864 & ~x867 & ~x906 & ~x984;
assign c5148 =  x89 &  x125 &  x236 &  x287 &  x320 &  x443 &  x452 &  x455 &  x583 &  x608 &  x610 &  x622 &  x661 &  x662 &  x743 &  x773 &  x959 &  x974 &  x1037 & ~x207 & ~x246 & ~x285 & ~x324 & ~x325 & ~x364 & ~x402 & ~x600;
assign c5150 =  x77 &  x134 &  x248 &  x610 &  x622 &  x649 &  x731 &  x793 &  x799 &  x842 &  x857 &  x883 &  x922 &  x1040 &  x1067 &  x1070 & ~x81 & ~x108 & ~x147 & ~x186 & ~x633 & ~x672 & ~x711 & ~x789;
assign c5152 =  x19 &  x58 &  x98 &  x136 &  x614 &  x1070 & ~x316 & ~x324 & ~x525 & ~x681 & ~x720 & ~x759;
assign c5154 =  x40 &  x41 &  x98 &  x157 &  x182 &  x206 &  x227 &  x254 &  x472 &  x545 &  x821 &  x974 & ~x4 & ~x186 & ~x246 & ~x366;
assign c5156 =  x58 &  x85 &  x97 &  x103 &  x124 &  x163 &  x173 &  x241 &  x280 &  x319 &  x353 &  x365 &  x367 &  x389 &  x407 &  x445 &  x484 &  x584 &  x605 &  x620 &  x770 &  x815 &  x830 &  x878 &  x934 &  x1034 & ~x558;
assign c5158 =  x11 &  x34 &  x72 &  x157 &  x215 &  x218 &  x236 &  x251 &  x302 &  x460 &  x470 &  x566 &  x649 &  x746 &  x759 &  x772 &  x785 &  x793 &  x955 &  x992 &  x994 &  x995 &  x1033 &  x1091 &  x1100 &  x1118 &  x1121;
assign c5160 =  x20 &  x44 &  x65 &  x137 &  x143 &  x152 &  x171 &  x172 &  x194 &  x210 &  x221 &  x249 &  x250 &  x266 &  x272 &  x311 &  x327 &  x341 &  x398 &  x431 &  x457 &  x467 &  x470 &  x490 &  x491 &  x496 &  x515 &  x568 &  x584 &  x590 &  x599 &  x607 &  x646 &  x656 &  x671 &  x680 &  x710 &  x746 &  x755 &  x769 &  x776 &  x788 &  x815 &  x824 &  x841 &  x860 &  x890 &  x923 &  x929 &  x977 &  x997 &  x1001 &  x1070 &  x1085 &  x1115 & ~x315;
assign c5162 =  x68 &  x629 &  x803 &  x901 &  x1019 & ~x472 & ~x621 & ~x660 & ~x699 & ~x798 & ~x835 & ~x837 & ~x874 & ~x913 & ~x951 & ~x952;
assign c5164 =  x23 &  x26 &  x46 &  x47 &  x53 &  x59 &  x62 &  x85 &  x98 &  x158 &  x203 &  x209 &  x221 &  x230 &  x233 &  x281 &  x290 &  x299 &  x302 &  x362 &  x365 &  x377 &  x380 &  x389 &  x461 &  x473 &  x497 &  x500 &  x512 &  x515 &  x521 &  x581 &  x593 &  x614 &  x644 &  x647 &  x659 &  x671 &  x674 &  x725 &  x737 &  x743 &  x770 &  x800 &  x803 &  x809 &  x815 &  x817 &  x827 &  x833 &  x871 &  x878 &  x890 &  x910 &  x944 &  x949 &  x962 &  x988 &  x1025 &  x1027 &  x1055 &  x1066 &  x1079 &  x1085 &  x1097 &  x1100 &  x1105 & ~x36 & ~x525 & ~x678 & ~x696;
assign c5166 =  x16 &  x61 &  x148 &  x178 &  x295 &  x334 &  x373 &  x397 &  x451 &  x475 &  x490 &  x523 &  x841 & ~x393 & ~x714 & ~x792;
assign c5168 =  x61 &  x211 &  x547 &  x586 &  x1070 & ~x237 & ~x442 & ~x481 & ~x519 & ~x520 & ~x559 & ~x598 & ~x714 & ~x753;
assign c5170 =  x5 &  x41 &  x58 &  x68 &  x71 &  x104 &  x113 &  x137 &  x143 &  x148 &  x170 &  x233 &  x242 &  x263 &  x266 &  x272 &  x314 &  x365 &  x368 &  x374 &  x377 &  x464 &  x473 &  x476 &  x521 &  x539 &  x581 &  x647 &  x707 &  x710 &  x776 &  x782 &  x788 &  x791 &  x803 &  x815 &  x860 &  x901 &  x929 &  x944 &  x959 &  x986 &  x1049 &  x1064 &  x1067 &  x1076 &  x1088 &  x1103 &  x1115 &  x1118 & ~x472 & ~x558 & ~x576 & ~x615 & ~x831 & ~x870;
assign c5172 =  x514 & ~x126 & ~x394 & ~x433 & ~x519 & ~x637 & ~x714 & ~x834;
assign c5174 =  x22 &  x34 &  x40 &  x61 &  x89 &  x209 &  x218 &  x266 &  x293 &  x296 &  x334 &  x353 &  x373 &  x473 &  x485 &  x551 &  x590 &  x596 &  x649 &  x650 &  x655 &  x694 &  x719 &  x749 &  x763 &  x806 &  x818 &  x853 &  x854 &  x872 &  x962 & ~x36 & ~x558 & ~x597 & ~x948 & ~x987;
assign c5176 =  x611 & ~x12 & ~x52 & ~x91 & ~x129 & ~x147 & ~x186 & ~x246 & ~x328 & ~x367 & ~x406;
assign c5178 =  x11 &  x29 &  x38 &  x47 &  x89 &  x107 &  x125 &  x146 &  x152 &  x158 &  x173 &  x176 &  x194 &  x197 &  x203 &  x215 &  x236 &  x266 &  x275 &  x347 &  x350 &  x362 &  x392 &  x395 &  x401 &  x443 &  x455 &  x470 &  x473 &  x475 &  x488 &  x494 &  x503 &  x514 &  x523 &  x527 &  x547 &  x551 &  x578 &  x584 &  x608 &  x623 &  x656 &  x677 &  x680 &  x686 &  x689 &  x695 &  x698 &  x701 &  x702 &  x703 &  x710 &  x758 &  x767 &  x773 &  x776 &  x782 &  x785 &  x788 &  x803 &  x809 &  x812 &  x833 &  x857 &  x860 &  x863 &  x875 &  x893 &  x914 &  x917 &  x929 &  x940 &  x962 &  x965 &  x980 &  x992 &  x1001 &  x1016 &  x1019 &  x1022 &  x1037 &  x1061 &  x1070 &  x1073 & ~x354 & ~x393 & ~x433 & ~x471 & ~x472 & ~x675 & ~x714 & ~x753 & ~x756 & ~x792 & ~x795 & ~x831 & ~x870 & ~x873;
assign c5180 =  x2 &  x17 &  x695 &  x974 &  x1018 &  x1056 &  x1057 &  x1095 &  x1096 & ~x399 & ~x628 & ~x667 & ~x870 & ~x987 & ~x1026 & ~x1027 & ~x1029 & ~x1065 & ~x1068;
assign c5182 =  x26 &  x41 &  x62 &  x116 &  x134 &  x140 &  x356 &  x368 &  x404 &  x410 &  x434 &  x551 &  x557 &  x584 &  x638 &  x653 &  x683 &  x818 &  x821 &  x839 &  x860 &  x890 &  x911 &  x932 &  x1031 &  x1058 &  x1070 &  x1073 &  x1076 &  x1100 &  x1109 & ~x199 & ~x238 & ~x246 & ~x285 & ~x324 & ~x441 & ~x442 & ~x480 & ~x481 & ~x519 & ~x990 & ~x1029;
assign c5184 =  x8 &  x59 &  x149 &  x152 &  x155 &  x164 &  x170 &  x242 &  x245 &  x248 &  x296 &  x305 &  x311 &  x320 &  x356 &  x362 &  x389 &  x425 &  x446 &  x461 &  x467 &  x470 &  x482 &  x506 &  x545 &  x566 &  x572 &  x605 &  x614 &  x644 &  x659 &  x713 &  x752 &  x803 &  x809 &  x860 &  x905 &  x923 &  x965 &  x974 &  x986 &  x992 &  x998 &  x1010 &  x1017 &  x1018 &  x1019 &  x1025 &  x1056 & ~x312 & ~x621 & ~x628 & ~x870 & ~x909 & ~x987 & ~x1029 & ~x1068;
assign c5186 =  x76 &  x143 &  x280 &  x340 &  x350 &  x379 &  x397 &  x418 &  x503 &  x674 &  x878 &  x928 &  x1084 &  x1106 & ~x393 & ~x480 & ~x519 & ~x525 & ~x558;
assign c5188 =  x71 &  x197 &  x293 &  x383 &  x386 &  x436 &  x475 &  x484 &  x490 &  x514 &  x523 &  x553 &  x568 &  x602 &  x773 &  x901 &  x905 &  x979 &  x1091 & ~x603 & ~x681 & ~x714 & ~x792 & ~x831 & ~x870 & ~x909 & ~x912;
assign c5190 =  x32 &  x68 &  x296 &  x299 &  x395 &  x524 &  x584 &  x622 &  x680 &  x878 &  x989 &  x1010 & ~x82 & ~x186 & ~x192 & ~x246 & ~x546 & ~x819;
assign c5192 =  x16 &  x229 &  x267 &  x437 &  x452 &  x467 &  x505 &  x622 &  x623 &  x659 &  x661 &  x763 &  x817 &  x934 & ~x399;
assign c5194 =  x8 &  x22 &  x35 &  x47 &  x61 &  x94 &  x100 &  x107 &  x148 &  x164 &  x230 &  x239 &  x248 &  x296 &  x299 &  x326 &  x365 &  x397 &  x406 &  x418 &  x436 &  x457 &  x475 &  x484 &  x514 &  x521 &  x568 &  x578 &  x607 &  x632 &  x641 &  x646 &  x652 &  x656 &  x691 &  x769 &  x782 &  x803 &  x847 &  x887 &  x932 &  x974 &  x1049 &  x1121;
assign c5196 =  x29 &  x32 &  x176 &  x202 &  x212 &  x227 &  x272 &  x329 &  x365 &  x368 &  x383 &  x410 &  x440 &  x452 &  x475 &  x503 &  x514 &  x523 &  x536 &  x547 &  x611 &  x745 &  x784 &  x806 &  x839 &  x854 &  x862 &  x887 &  x929 &  x940 &  x995 &  x1013 &  x1100 &  x1121 & ~x394 & ~x433 & ~x675 & ~x714 & ~x795 & ~x834;
assign c5198 =  x29 &  x47 &  x80 &  x116 &  x125 &  x131 &  x149 &  x158 &  x164 &  x209 &  x224 &  x311 &  x344 &  x398 &  x404 &  x407 &  x422 &  x428 &  x437 &  x461 &  x473 &  x515 &  x539 &  x554 &  x566 &  x578 &  x614 &  x641 &  x668 &  x713 &  x734 &  x744 &  x745 &  x749 &  x791 &  x797 &  x815 &  x869 &  x878 &  x917 &  x989 &  x1007 &  x1025 &  x1040 &  x1043 &  x1076 &  x1079 &  x1097 &  x1112 &  x1115 & ~x198 & ~x237 & ~x316 & ~x324 & ~x363 & ~x480 & ~x519 & ~x597 & ~x675 & ~x678 & ~x714 & ~x720 & ~x756 & ~x834;
assign c5200 =  x86 &  x455 &  x458 &  x530 &  x971 & ~x48 & ~x525 & ~x837 & ~x846 & ~x874 & ~x885 & ~x913 & ~x952 & ~x990 & ~x991 & ~x1029 & ~x1068;
assign c5202 =  x155 &  x212 &  x488 &  x581 &  x620 &  x1040 &  x1130 & ~x9 & ~x238 & ~x277 & ~x316 & ~x453 & ~x465 & ~x525 & ~x718;
assign c5204 =  x119 &  x161 &  x173 &  x191 &  x209 &  x272 &  x313 &  x338 &  x368 &  x371 &  x377 &  x386 &  x407 &  x419 &  x446 &  x464 &  x494 &  x563 &  x602 &  x632 &  x677 &  x680 &  x686 &  x764 &  x773 &  x788 &  x818 &  x827 &  x875 &  x908 &  x917 &  x1004 &  x1040 &  x1043 &  x1049 &  x1064 &  x1070 &  x1106 &  x1124 & ~x3 & ~x4 & ~x42 & ~x186 & ~x253 & ~x405 & ~x780;
assign c5206 =  x32 &  x40 &  x47 &  x86 &  x146 &  x152 &  x254 &  x257 &  x296 &  x312 &  x326 &  x332 &  x350 &  x452 &  x539 &  x613 &  x680 &  x872 &  x995 &  x1067 & ~x82 & ~x180 & ~x363;
assign c5208 =  x206 &  x257 &  x434 &  x523 &  x553 &  x605 &  x625 &  x703 &  x722 &  x818 &  x863 &  x890 &  x901 &  x1040 &  x1096 & ~x519 & ~x558 & ~x621 & ~x714 & ~x792 & ~x831 & ~x837 & ~x870 & ~x909;
assign c5210 =  x40 &  x94 &  x98 &  x229 &  x410 &  x535 &  x763 &  x767 &  x781 &  x808 &  x1009 &  x1130 & ~x36 & ~x789 & ~x906;
assign c5212 =  x29 &  x56 &  x68 &  x80 &  x89 &  x97 &  x113 &  x115 &  x155 &  x206 &  x239 &  x245 &  x248 &  x266 &  x293 &  x359 &  x377 &  x464 &  x530 &  x553 &  x572 &  x578 &  x617 &  x716 &  x725 &  x746 &  x761 &  x803 &  x821 &  x861 &  x872 &  x893 &  x940 &  x941 &  x1034 &  x1070 & ~x354 & ~x432 & ~x433 & ~x472 & ~x510 & ~x714 & ~x876;
assign c5214 =  x65 &  x296 &  x461 &  x553 &  x631 &  x832 &  x866 &  x875 &  x953 &  x1004 &  x1060 &  x1070 &  x1088 & ~x207 & ~x246 & ~x852 & ~x879 & ~x918 & ~x969 & ~x1035 & ~x1047;
assign c5216 =  x92 &  x95 &  x104 &  x157 &  x179 &  x185 &  x196 &  x284 &  x437 &  x470 &  x610 &  x649 &  x671 &  x677 &  x752 &  x776 &  x821 &  x871 &  x883 &  x922 &  x950 &  x982 &  x1060 &  x1070 & ~x108 & ~x147 & ~x186 & ~x225 & ~x483 & ~x633;
assign c5218 =  x19 &  x29 &  x37 &  x56 &  x58 &  x97 &  x101 &  x116 &  x245 &  x251 &  x269 &  x341 &  x368 &  x407 &  x455 &  x599 &  x605 &  x611 &  x745 &  x791 &  x809 &  x827 &  x833 &  x854 &  x989 &  x1046 &  x1070 & ~x276 & ~x316 & ~x355 & ~x525 & ~x603 & ~x681 & ~x720 & ~x759;
assign c5220 =  x109 &  x209 &  x523 &  x614 &  x1076 & ~x433 & ~x486 & ~x675 & ~x714 & ~x718 & ~x753 & ~x757 & ~x792 & ~x795 & ~x796 & ~x835;
assign c5222 =  x26 &  x32 &  x74 &  x79 &  x107 &  x119 &  x157 &  x170 &  x200 &  x206 &  x224 &  x235 &  x257 &  x312 &  x401 &  x500 &  x638 &  x1031 &  x1070 &  x1097 & ~x82 & ~x324 & ~x402 & ~x711 & ~x750 & ~x789;
assign c5224 =  x155 &  x275 &  x352 &  x547 &  x584 &  x632 &  x818 &  x1025 & ~x199 & ~x238 & ~x277 & ~x480 & ~x519 & ~x525 & ~x558 & ~x561 & ~x600 & ~x678;
assign c5226 =  x32 &  x62 &  x80 &  x101 &  x155 &  x182 &  x197 &  x215 &  x224 &  x242 &  x274 &  x311 &  x314 &  x334 &  x401 &  x407 &  x425 &  x509 &  x512 &  x521 &  x536 &  x545 &  x566 &  x638 &  x662 &  x689 &  x725 &  x749 &  x766 &  x871 &  x875 &  x878 &  x889 &  x902 &  x911 &  x949 &  x983 &  x988 &  x1016 &  x1027 &  x1066 &  x1078 &  x1084 &  x1088 &  x1109 &  x1111 &  x1117 & ~x246 & ~x324 & ~x561 & ~x600 & ~x858;
assign c5228 =  x46 &  x163 &  x202 &  x211 &  x250 &  x280 &  x289 &  x475 &  x514 &  x617 &  x826 &  x953 & ~x441 & ~x480 & ~x525;
assign c5230 =  x17 &  x26 &  x29 &  x62 &  x74 &  x80 &  x86 &  x116 &  x131 &  x206 &  x212 &  x236 &  x245 &  x263 &  x266 &  x311 &  x314 &  x323 &  x335 &  x346 &  x383 &  x389 &  x416 &  x452 &  x488 &  x491 &  x500 &  x512 &  x530 &  x536 &  x539 &  x547 &  x560 &  x575 &  x596 &  x608 &  x617 &  x620 &  x626 &  x653 &  x662 &  x680 &  x686 &  x725 &  x743 &  x746 &  x764 &  x766 &  x788 &  x797 &  x800 &  x803 &  x805 &  x812 &  x818 &  x836 &  x839 &  x844 &  x845 &  x863 &  x881 &  x890 &  x896 &  x902 &  x911 &  x923 &  x929 &  x980 &  x989 &  x995 &  x1004 &  x1007 &  x1031 &  x1034 &  x1046 &  x1106 & ~x237 & ~x276 & ~x316 & ~x486 & ~x525 & ~x600 & ~x603 & ~x642 & ~x678 & ~x681;
assign c5232 =  x242 &  x530 &  x566 &  x575 &  x581 &  x587 &  x610 &  x632 &  x710 &  x815 &  x818 &  x917 &  x1004 & ~x82 & ~x121 & ~x252 & ~x265 & ~x303 & ~x447;
assign c5234 =  x32 &  x40 &  x41 &  x59 &  x86 &  x92 &  x107 &  x125 &  x158 &  x206 &  x257 &  x273 &  x314 &  x354 &  x394 &  x440 &  x467 &  x482 &  x485 &  x641 &  x644 &  x677 &  x689 &  x695 &  x740 &  x749 &  x773 &  x806 &  x839 &  x869 &  x929 &  x974 &  x1115 & ~x42 & ~x246 & ~x546;
assign c5236 =  x143 &  x206 &  x235 &  x389 & ~x199 & ~x238 & ~x277 & ~x483 & ~x523 & ~x558 & ~x562 & ~x678;
assign c5238 =  x83 &  x752 &  x1127 & ~x439 & ~x555 & ~x633 & ~x672 & ~x864 & ~x870 & ~x903 & ~x910;
assign c5240 =  x8 &  x26 &  x29 &  x134 &  x389 &  x647 &  x863 &  x1022 &  x1040 &  x1127 & ~x316 & ~x355 & ~x393 & ~x442 & ~x480 & ~x519 & ~x718 & ~x757;
assign c5242 =  x936 &  x975 &  x1017 &  x1095 & ~x399 & ~x471 & ~x667 & ~x987 & ~x1026 & ~x1029;
assign c5244 =  x2 &  x17 &  x23 &  x26 &  x29 &  x83 &  x116 &  x125 &  x143 &  x161 &  x173 &  x182 &  x284 &  x299 &  x326 &  x338 &  x341 &  x413 &  x518 &  x536 &  x641 &  x662 &  x727 &  x743 &  x764 &  x770 &  x788 &  x797 &  x818 &  x1010 &  x1052 &  x1103 & ~x82 & ~x246 & ~x600 & ~x820 & ~x859 & ~x990 & ~x1047 & ~x1086;
assign c5246 =  x11 &  x17 &  x32 &  x44 &  x50 &  x71 &  x89 &  x101 &  x116 &  x122 &  x125 &  x131 &  x134 &  x137 &  x143 &  x158 &  x167 &  x206 &  x209 &  x212 &  x236 &  x239 &  x263 &  x293 &  x338 &  x353 &  x362 &  x365 &  x422 &  x428 &  x464 &  x479 &  x482 &  x494 &  x509 &  x512 &  x545 &  x554 &  x557 &  x569 &  x590 &  x599 &  x611 &  x614 &  x629 &  x635 &  x649 &  x665 &  x677 &  x680 &  x683 &  x707 &  x710 &  x737 &  x740 &  x743 &  x746 &  x758 &  x764 &  x766 &  x767 &  x770 &  x779 &  x782 &  x791 &  x827 &  x842 &  x854 &  x863 &  x866 &  x869 &  x896 &  x917 &  x920 &  x932 &  x949 &  x955 &  x956 &  x965 &  x971 &  x983 &  x988 &  x989 &  x994 &  x1004 &  x1031 &  x1034 &  x1049 &  x1058 &  x1066 &  x1091 &  x1103 &  x1106 &  x1121 & ~x246 & ~x285 & ~x324 & ~x519 & ~x558 & ~x597 & ~x678 & ~x789 & ~x828 & ~x867;
assign c5248 =  x23 &  x40 &  x44 &  x47 &  x50 &  x74 &  x104 &  x209 &  x230 &  x308 &  x341 &  x377 &  x419 &  x527 &  x581 &  x599 &  x680 &  x725 &  x802 &  x833 &  x989 &  x998 &  x1007 &  x1031 &  x1064 &  x1070 &  x1091 &  x1112 & ~x24 & ~x63 & ~x64 & ~x102 & ~x246 & ~x285 & ~x555 & ~x600 & ~x633 & ~x672 & ~x828;
assign c5250 =  x29 &  x35 &  x202 &  x254 &  x266 &  x326 &  x440 &  x484 &  x625 &  x692 &  x703 &  x710 &  x1037 &  x1055 &  x1067 &  x1115 & ~x433 & ~x480 & ~x519 & ~x675 & ~x720 & ~x756 & ~x759 & ~x796 & ~x798 & ~x873;
assign c5252 =  x23 &  x44 &  x107 &  x143 &  x149 &  x197 &  x206 &  x209 &  x257 &  x263 &  x305 &  x334 &  x338 &  x398 &  x440 &  x443 &  x446 &  x451 &  x460 &  x518 &  x548 &  x568 &  x574 &  x607 &  x618 &  x626 &  x632 &  x638 &  x671 &  x692 &  x724 &  x742 &  x767 &  x781 &  x809 &  x820 &  x842 &  x859 &  x887 &  x898 &  x953 &  x968 &  x992 &  x1016 &  x1052 &  x1057 &  x1096 &  x1100 & ~x831 & ~x870 & ~x909 & ~x948;
assign c5254 =  x368 &  x389 &  x626 &  x731 & ~x316 & ~x480 & ~x519 & ~x520 & ~x525 & ~x676 & ~x714;
assign c5256 =  x2 &  x13 &  x109 &  x158 &  x182 &  x275 &  x278 &  x314 &  x377 &  x389 &  x407 &  x422 &  x440 &  x461 &  x548 &  x551 &  x572 &  x581 &  x593 &  x596 &  x602 &  x632 &  x692 &  x703 &  x731 &  x744 &  x749 &  x755 &  x758 &  x785 &  x803 &  x809 &  x860 &  x872 &  x956 &  x965 &  x992 &  x1007 &  x1016 &  x1034 &  x1037 &  x1076 &  x1094 &  x1112 &  x1118 & ~x117 & ~x156 & ~x678 & ~x718 & ~x756 & ~x757 & ~x759 & ~x795 & ~x796 & ~x835;
assign c5258 =  x23 &  x47 &  x167 &  x170 &  x181 &  x197 &  x203 &  x257 &  x260 &  x299 &  x359 &  x380 &  x392 &  x397 &  x401 &  x436 &  x475 &  x490 &  x523 &  x553 &  x562 &  x568 &  x579 &  x815 &  x830 &  x854 &  x887 &  x923 &  x1018 &  x1031 &  x1067 &  x1076 &  x1079 &  x1130 & ~x621;
assign c5260 =  x2 &  x8 &  x29 &  x95 &  x146 &  x155 &  x161 &  x182 &  x203 &  x224 &  x251 &  x326 &  x344 &  x365 &  x386 &  x404 &  x511 &  x530 &  x560 &  x593 &  x722 &  x740 &  x767 &  x878 &  x884 &  x917 &  x938 &  x947 &  x977 &  x995 &  x1007 &  x1019 &  x1076 &  x1078 &  x1106 & ~x160 & ~x199 & ~x207 & ~x238 & ~x246 & ~x324 & ~x402 & ~x561 & ~x600 & ~x1047 & ~x1086;
assign c5262 =  x40 &  x71 &  x72 &  x178 &  x191 &  x206 &  x397 &  x475 &  x617 &  x649 &  x688 &  x826 &  x836 &  x895 &  x914 &  x916 &  x934 &  x955 &  x994 &  x1043 &  x1066;
assign c5264 =  x2 &  x5 &  x11 &  x32 &  x44 &  x104 &  x122 &  x158 &  x182 &  x224 &  x230 &  x236 &  x245 &  x251 &  x293 &  x320 &  x329 &  x380 &  x389 &  x416 &  x440 &  x461 &  x506 &  x530 &  x566 &  x590 &  x644 &  x647 &  x662 &  x668 &  x716 &  x725 &  x785 &  x815 &  x818 &  x821 &  x824 &  x845 &  x890 &  x896 &  x908 &  x916 &  x932 &  x955 &  x968 &  x994 &  x1001 &  x1025 &  x1028 &  x1079 &  x1085 &  x1091 &  x1094 &  x1097 &  x1118 & ~x42 & ~x82 & ~x90 & ~x91 & ~x121 & ~x129 & ~x246;
assign c5266 =  x40 &  x47 &  x79 &  x86 &  x116 &  x137 &  x157 &  x206 &  x239 &  x260 &  x284 &  x350 &  x352 &  x389 &  x473 &  x509 &  x530 &  x536 &  x560 &  x566 &  x578 &  x581 &  x587 &  x593 &  x608 &  x626 &  x629 &  x638 &  x761 &  x773 &  x793 &  x821 &  x848 &  x863 &  x866 &  x878 &  x884 &  x890 &  x935 &  x950 &  x953 &  x1013 &  x1043 &  x1046 &  x1064 &  x1085 & ~x12 & ~x108 & ~x147 & ~x186 & ~x246 & ~x291 & ~x444 & ~x483 & ~x633 & ~x672 & ~x828;
assign c5268 =  x858 &  x897 &  x936 &  x1017 &  x1056 &  x1095 &  x1096 & ~x667 & ~x777 & ~x987;
assign c5270 =  x20 &  x32 &  x83 &  x116 &  x284 &  x296 &  x338 &  x350 &  x362 &  x413 &  x416 &  x419 &  x443 &  x446 &  x479 &  x513 &  x514 &  x515 &  x548 &  x553 &  x575 &  x605 &  x626 &  x644 &  x692 &  x701 &  x707 &  x776 &  x779 &  x785 &  x872 &  x920 &  x938 &  x968 &  x971 &  x1018 &  x1088 &  x1094 & ~x87 & ~x510 & ~x589;
assign c5272 =  x32 &  x266 &  x916 &  x917 &  x955 &  x994 &  x1032 &  x1033 &  x1071 &  x1111 & ~x297 & ~x639 & ~x678 & ~x828 & ~x885 & ~x906;
assign c5274 =  x155 &  x194 &  x206 &  x475 &  x553 &  x592 &  x631 &  x773 &  x819 &  x858 &  x896 &  x926 &  x932 &  x939 & ~x550 & ~x589 & ~x628;
assign c5276 =  x17 &  x26 &  x143 &  x155 &  x197 &  x233 &  x275 &  x284 &  x311 &  x352 &  x380 &  x416 &  x422 &  x443 &  x581 &  x626 &  x656 &  x701 &  x707 &  x770 &  x815 &  x842 &  x869 &  x872 &  x875 &  x902 &  x905 &  x917 &  x956 &  x1013 &  x1025 &  x1040 &  x1046 &  x1070 &  x1109 &  x1130 & ~x24 & ~x63 & ~x102 & ~x219 & ~x220 & ~x258 & ~x483 & ~x484 & ~x789 & ~x828 & ~x885;
assign c5278 =  x53 &  x86 &  x224 &  x395 &  x397 &  x406 &  x470 &  x524 &  x848 &  x953 &  x1118 &  x1124 & ~x355 & ~x519 & ~x558 & ~x559 & ~x598 & ~x637 & ~x676 & ~x714 & ~x753 & ~x831;
assign c5280 =  x16 &  x32 &  x40 &  x55 &  x59 &  x80 &  x83 &  x94 &  x118 &  x128 &  x133 &  x149 &  x155 &  x157 &  x158 &  x182 &  x194 &  x215 &  x221 &  x235 &  x266 &  x293 &  x312 &  x344 &  x352 &  x362 &  x401 &  x446 &  x458 &  x524 &  x560 &  x596 &  x608 &  x623 &  x635 &  x641 &  x644 &  x649 &  x653 &  x656 &  x659 &  x671 &  x688 &  x689 &  x695 &  x701 &  x704 &  x734 &  x746 &  x752 &  x770 &  x776 &  x788 &  x824 &  x845 &  x887 &  x917 &  x1007 &  x1016 &  x1019 &  x1088 &  x1094 &  x1100 &  x1112 & ~x82 & ~x252;
assign c5282 =  x125 &  x547 &  x557 &  x659 &  x815 &  x1013 & ~x9 & ~x48 & ~x238 & ~x277 & ~x316 & ~x621 & ~x846 & ~x885 & ~x1002;
assign c5284 =  x5 &  x17 &  x29 &  x92 &  x155 &  x188 &  x233 &  x248 &  x413 &  x419 &  x425 &  x503 &  x518 &  x575 &  x611 &  x620 &  x689 &  x803 &  x830 &  x854 &  x869 &  x893 &  x998 &  x1001 &  x1025 &  x1028 &  x1033 &  x1070 &  x1103 &  x1124 & ~x160 & ~x207 & ~x246 & ~x285 & ~x324 & ~x363 & ~x402 & ~x561 & ~x562 & ~x600 & ~x696 & ~x780;
assign c5286 =  x428 & ~x4 & ~x169 & ~x208 & ~x246 & ~x247 & ~x285 & ~x286 & ~x324 & ~x325 & ~x480 & ~x519;
assign c5288 =  x16 &  x110 &  x118 &  x157 &  x311 &  x607 &  x646 &  x724 &  x763 &  x815 & ~x247 & ~x285 & ~x286 & ~x324 & ~x325 & ~x402 & ~x403 & ~x519;
assign c5290 =  x16 &  x34 &  x71 &  x72 &  x98 &  x313 &  x356 &  x466 &  x490 &  x503 &  x527 &  x568 &  x607 &  x622 &  x685 &  x724 &  x769 &  x797 &  x800 &  x808 &  x841 &  x853 &  x872 &  x878 &  x880 &  x1018 &  x1028 &  x1057 &  x1087 &  x1120;
assign c5292 =  x28 &  x32 &  x34 &  x40 &  x44 &  x61 &  x100 &  x143 &  x182 &  x194 &  x206 &  x395 &  x404 &  x410 &  x422 &  x509 &  x524 &  x614 &  x632 &  x650 &  x655 &  x659 &  x731 &  x770 &  x810 &  x893 &  x916 &  x917 &  x955 &  x968 &  x974 &  x994 &  x1043 &  x1052 &  x1060 &  x1106 &  x1112 &  x1120;
assign c5294 =  x158 &  x188 &  x206 &  x257 &  x380 &  x437 &  x512 &  x518 &  x536 &  x551 &  x569 &  x770 &  x779 &  x878 &  x901 &  x974 &  x998 & ~x315 & ~x316 & ~x324 & ~x402 & ~x480 & ~x486 & ~x519 & ~x558 & ~x564 & ~x642 & ~x681 & ~x714 & ~x720 & ~x753 & ~x792 & ~x837;
assign c5296 =  x19 &  x50 &  x58 &  x74 &  x85 &  x86 &  x92 &  x97 &  x149 &  x161 &  x202 &  x215 &  x230 &  x241 &  x263 &  x272 &  x319 &  x326 &  x347 &  x362 &  x383 &  x389 &  x401 &  x470 &  x530 &  x547 &  x581 &  x584 &  x608 &  x665 &  x698 &  x766 &  x869 &  x887 &  x896 &  x1049 &  x1082 &  x1106 & ~x316;
assign c5298 =  x38 &  x125 &  x176 &  x245 &  x266 &  x269 &  x296 &  x305 &  x359 &  x437 &  x497 &  x653 &  x764 &  x782 &  x857 &  x901 &  x939 &  x947 &  x978 &  x1004 &  x1007 &  x1017 &  x1031 &  x1034 &  x1052 &  x1056 &  x1057 &  x1096 &  x1097 & ~x429 & ~x511 & ~x550 & ~x714 & ~x792 & ~x831 & ~x909 & ~x948 & ~x1029 & ~x1068;
assign c51 =  x427 &  x487 & ~x240 & ~x708 & ~x786 & ~x1071;
assign c53 =  x220 &  x226 &  x469 & ~x195 & ~x435 & ~x513 & ~x514;
assign c55 =  x472 &  x991 & ~x111 & ~x249 & ~x723;
assign c57 = ~x426 & ~x570 & ~x823 & ~x901 & ~x939 & ~x978 & ~x1095;
assign c59 =  x43 &  x71 &  x82 &  x160 &  x199 &  x242 &  x311 &  x332 &  x335 &  x344 &  x467 &  x563 &  x721 &  x722 &  x760 &  x854 &  x1061 & ~x309 & ~x936;
assign c511 = ~x630 & ~x709 & ~x927;
assign c513 =  x26 &  x68 &  x166 &  x168 &  x205 &  x208 &  x277 &  x896 &  x1094 & ~x0;
assign c515 =  x43 &  x82 &  x121 &  x160 &  x199 &  x238 &  x277 &  x311 &  x539 &  x542 &  x614 &  x713 &  x815 &  x1025 &  x1040 &  x1043 &  x1045 & ~x303 & ~x900;
assign c517 =  x161 &  x167 &  x188 &  x238 &  x548 &  x584 &  x811 & ~x72 & ~x111 & ~x939 & ~x978 & ~x1017 & ~x1056 & ~x1095;
assign c519 =  x31 &  x720 &  x911 & ~x105 & ~x333;
assign c521 =  x481 &  x492 & ~x312 & ~x670 & ~x1050;
assign c523 =  x190 &  x283 &  x463 &  x1063 & ~x273 & ~x921;
assign c525 =  x104 &  x155 &  x167 &  x316 &  x335 &  x560 &  x608 &  x725 &  x752 &  x830 &  x1007 &  x1046 & ~x78 & ~x93 & ~x111 & ~x897 & ~x936 & ~x1092 & ~x1101;
assign c527 =  x67 &  x247 &  x253 &  x259 &  x280 &  x587 &  x1106 & ~x435 & ~x474 & ~x513 & ~x552;
assign c529 =  x4 &  x170 &  x238 &  x277 &  x446 &  x463 &  x533 &  x881 &  x1100 & ~x378;
assign c531 =  x108 & ~x334;
assign c533 =  x238 &  x551 & ~x27 & ~x54 & ~x150 & ~x240 & ~x279;
assign c535 =  x17 &  x44 &  x53 &  x223 &  x254 &  x290 &  x301 &  x304 &  x310 &  x364 &  x376 &  x388 &  x403 &  x427 &  x442 &  x448 &  x527 &  x623 &  x745 &  x1010 &  x1024 & ~x390;
assign c537 =  x82 &  x709 &  x748 &  x865 &  x1012 & ~x306;
assign c539 =  x370 &  x442 &  x478 &  x624 & ~x591;
assign c541 =  x370 &  x414 & ~x631;
assign c543 =  x364 &  x376 &  x442 &  x596 &  x706 &  x820 &  x1037 & ~x474 & ~x513 & ~x552 & ~x708;
assign c545 =  x208 & ~x687 & ~x901 & ~x1095;
assign c547 =  x78 &  x82 &  x117 &  x473 &  x718 &  x952 & ~x75 & ~x123 & ~x1098;
assign c549 =  x52 &  x238 &  x524 &  x656 &  x1049 & ~x72 & ~x144 & ~x939 & ~x978 & ~x1017;
assign c551 =  x4 &  x43 &  x82 &  x121 &  x155 &  x160 &  x167 &  x194 &  x199 &  x206 &  x215 &  x238 &  x266 &  x560 &  x683 &  x884 &  x1001 &  x1034 &  x1045 &  x1094 &  x1121 & ~x69 & ~x375 & ~x666;
assign c553 =  x106 &  x182 &  x632 &  x872 & ~x306 & ~x495 & ~x513 & ~x552 & ~x630;
assign c555 =  x184 &  x789 & ~x594;
assign c557 =  x403 &  x442 &  x493 &  x526 &  x706 &  x809 & ~x882 & ~x960 & ~x1077 & ~x1116;
assign c559 =  x77 &  x382 &  x421 &  x493 &  x575 &  x1067 & ~x312 & ~x390 & ~x618 & ~x843 & ~x960 & ~x1038 & ~x1116;
assign c561 =  x4 &  x595 &  x638 &  x721 &  x748 &  x998 & ~x123 & ~x162;
assign c563 =  x472 &  x752 & ~x79 & ~x267 & ~x333 & ~x1092;
assign c565 =  x271 &  x361 &  x913 &  x991 & ~x687;
assign c567 =  x68 &  x80 &  x121 &  x179 &  x199 &  x224 &  x238 &  x274 &  x277 &  x391 &  x404 &  x473 &  x542 &  x590 &  x674 &  x707 &  x713 &  x746 &  x755 &  x757 &  x782 &  x809 &  x824 &  x833 &  x944 &  x1007 &  x1055 &  x1064 & ~x453 & ~x666 & ~x900 & ~x939;
assign c569 =  x4 &  x5 &  x43 &  x56 &  x82 &  x121 &  x128 &  x137 &  x143 &  x160 &  x196 &  x199 &  x227 &  x238 &  x269 &  x275 &  x341 &  x356 &  x401 &  x425 &  x428 &  x455 &  x542 &  x608 &  x620 &  x629 &  x668 &  x670 &  x671 &  x701 &  x746 &  x770 &  x782 &  x836 &  x842 &  x851 &  x1001 &  x1028 &  x1100 & ~x897 & ~x1101;
assign c571 =  x20 &  x119 &  x170 &  x238 &  x277 &  x308 &  x332 &  x485 &  x719 &  x749 &  x902 &  x926 &  x1090 & ~x27 & ~x780 & ~x1014 & ~x1092;
assign c573 =  x4 &  x82 &  x199 &  x238 &  x361 &  x517 &  x530 &  x1018;
assign c575 =  x271 &  x283 &  x952 &  x991 & ~x84;
assign c577 =  x706 & ~x306 & ~x967 & ~x1005;
assign c579 =  x166 &  x169 &  x205 &  x244 &  x247 &  x1064 &  x1127 & ~x435 & ~x474 & ~x513 & ~x777;
assign c581 =  x386 &  x427 & ~x57 & ~x513 & ~x934 & ~x1011 & ~x1032;
assign c583 =  x796 &  x951 &  x1048 & ~x162 & ~x1077;
assign c585 =  x208 &  x247 &  x589 & ~x345 & ~x849 & ~x1092;
assign c587 =  x427 & ~x123 & ~x162 & ~x201 & ~x240 & ~x318 & ~x669 & ~x825 & ~x1032 & ~x1038 & ~x1044;
assign c589 =  x64 &  x107 &  x134 &  x175 &  x197 &  x338 &  x398 &  x433 &  x479 &  x617 &  x620 &  x713 &  x740 &  x785 &  x857 &  x863 &  x929 &  x983 &  x1043 & ~x40 & ~x79 & ~x189 & ~x858;
assign c591 =  x121 &  x234 &  x718 &  x757 & ~x241;
assign c593 =  x314 &  x364 &  x370 &  x403 &  x419 &  x421 &  x667 &  x1016 & ~x843 & ~x882 & ~x921 & ~x1044;
assign c595 =  x68 &  x215 &  x292 &  x364 &  x428 &  x628 &  x686 &  x740 & ~x384 & ~x456 & ~x495 & ~x1092;
assign c597 =  x82 &  x159 &  x173 &  x199 &  x488 &  x560 &  x593 &  x659 &  x1082 & ~x294 & ~x858;
assign c599 =  x17 &  x307 &  x757 &  x938 & ~x30 & ~x582 & ~x939 & ~x1017 & ~x1056 & ~x1083 & ~x1095;
assign c5101 =  x151 &  x364 &  x385 &  x403 &  x425 &  x526 &  x598 &  x848 &  x893 &  x1102 & ~x507 & ~x1050;
assign c5103 =  x292 &  x297 &  x336 &  x364 &  x667 &  x1024;
assign c5105 =  x442 & ~x120 & ~x669 & ~x708 & ~x786 & ~x921;
assign c5107 =  x259 &  x265 &  x511 &  x906;
assign c5109 =  x154 &  x193 &  x355 & ~x117 & ~x534 & ~x978;
assign c5111 =  x714 & ~x771 & ~x1020;
assign c5113 =  x43 &  x82 &  x89 &  x101 &  x104 &  x118 &  x121 &  x160 &  x188 &  x199 &  x212 &  x224 &  x235 &  x239 &  x251 &  x272 &  x296 &  x311 &  x314 &  x338 &  x350 &  x380 &  x404 &  x407 &  x443 &  x473 &  x494 &  x506 &  x524 &  x533 &  x566 &  x593 &  x734 &  x773 &  x821 &  x827 &  x850 &  x854 &  x881 &  x889 &  x959 &  x967 &  x998 &  x1006 &  x1007 &  x1045 &  x1049 &  x1079 &  x1121 & ~x666 & ~x900;
assign c5115 =  x409 &  x493 &  x783 & ~x391 & ~x540;
assign c5117 =  x487 &  x667 & ~x456 & ~x534 & ~x573 & ~x1077 & ~x1116;
assign c5119 =  x337 &  x403 &  x425 &  x624 & ~x474 & ~x513;
assign c5121 =  x226 &  x265 &  x299 &  x314 &  x335 &  x364 &  x403 &  x458 &  x628 &  x629 &  x683 &  x722 &  x1088 & ~x313;
assign c5123 =  x559 & ~x391 & ~x1005;
assign c5125 =  x376 &  x493 & ~x79 & ~x306;
assign c5127 =  x523 &  x796 & ~x993 & ~x1018 & ~x1057;
assign c5129 =  x82 &  x238 &  x718 &  x1024 &  x1042 &  x1102 &  x1114 & ~x303;
assign c5131 =  x4 &  x199 & ~x588 & ~x1017 & ~x1032;
assign c5133 =  x421 &  x448 &  x520 &  x784 & ~x618 & ~x768;
assign c5135 =  x421 &  x667 & ~x30 & ~x507 & ~x804 & ~x921 & ~x1005 & ~x1038;
assign c5137 =  x258 &  x511 & ~x40;
assign c5139 = ~x6 & ~x33 & ~x144 & ~x249 & ~x684 & ~x900 & ~x1056 & ~x1095;
assign c5141 =  x181 &  x511 &  x632 &  x828 & ~x273;
assign c5143 =  x292 &  x409 &  x414 &  x453 &  x493 &  x674 &  x725 &  x953 & ~x747;
assign c5145 =  x4 &  x11 &  x82 &  x121 &  x137 &  x160 &  x161 &  x199 &  x287 &  x352 &  x682 &  x721 &  x734 &  x883 &  x905 &  x980 &  x1115 &  x1129 & ~x663 & ~x936;
assign c5147 = ~x993 & ~x1038 & ~x1057;
assign c5149 =  x59 &  x82 &  x95 &  x238 &  x458 & ~x33 & ~x1017;
assign c5151 =  x358 &  x388 &  x487 & ~x274 & ~x277;
assign c5153 =  x331 &  x564 &  x667 &  x745;
assign c5155 =  x181 &  x624 & ~x345 & ~x553 & ~x670;
assign c5157 =  x40 &  x166 &  x388 &  x419 &  x911 &  x952 &  x1076 &  x1109 & ~x6 & ~x396;
assign c5159 =  x43 &  x82 &  x159 &  x199 &  x238 & ~x333;
assign c5161 =  x427 & ~x669 & ~x786 & ~x825 & ~x1129;
assign c5163 =  x478 &  x760 & ~x54 & ~x358;
assign c5165 =  x5 &  x41 &  x56 &  x74 &  x82 &  x113 &  x134 &  x140 &  x160 &  x199 &  x215 &  x235 &  x238 &  x284 &  x353 &  x365 &  x416 &  x449 &  x470 &  x515 &  x566 &  x593 &  x596 &  x740 &  x748 &  x767 &  x887 &  x956 &  x962 &  x965 &  x983 &  x1025 &  x1055 &  x1079 &  x1085 &  x1097 &  x1121 &  x1127 & ~x303 & ~x897;
assign c5167 =  x20 &  x32 &  x64 &  x124 &  x137 &  x143 &  x155 &  x161 &  x170 &  x176 &  x203 &  x206 &  x218 &  x227 &  x277 &  x278 &  x293 &  x316 &  x329 &  x335 &  x371 &  x380 &  x383 &  x394 &  x433 &  x503 &  x506 &  x512 &  x542 &  x575 &  x587 &  x590 &  x626 &  x644 &  x668 &  x680 &  x722 &  x728 &  x740 &  x743 &  x767 &  x773 &  x803 &  x818 &  x830 &  x839 &  x878 &  x887 &  x893 &  x935 &  x938 &  x971 &  x974 &  x1004 &  x1013 &  x1019 &  x1028 &  x1049 &  x1052 &  x1064 &  x1085 &  x1112 &  x1118 &  x1130 & ~x117 & ~x435;
assign c5169 =  x127 &  x155 &  x347 &  x424 &  x425 &  x463 &  x500 &  x506 &  x569 &  x623 &  x647 &  x757 &  x758 &  x818 &  x1001 &  x1025 & ~x30 & ~x1083 & ~x1095 & ~x1110;
assign c5171 =  x4 &  x155 &  x874 & ~x358;
assign c5173 =  x364 &  x442 &  x487 &  x595 &  x820 &  x862 &  x893 & ~x618;
assign c5175 =  x4 &  x26 &  x43 &  x98 &  x119 &  x121 &  x125 &  x160 &  x199 &  x206 &  x230 &  x233 &  x236 &  x238 &  x277 &  x365 &  x374 &  x443 &  x503 &  x533 &  x587 &  x593 &  x644 &  x659 &  x739 &  x860 &  x869 &  x917 &  x992 &  x1001 & ~x303 & ~x897;
assign c5177 =  x233 &  x237 & ~x72 & ~x858 & ~x1092;
assign c5179 =  x376 &  x403 &  x442 &  x448 &  x559 &  x667 &  x745 &  x809 & ~x915 & ~x1032;
assign c5181 =  x4 &  x41 &  x82 &  x121 &  x199 &  x721 &  x733 &  x739 &  x760 &  x767 &  x799 &  x838 &  x905 &  x1045 & ~x1053;
assign c5183 =  x507 & ~x306 & ~x435 & ~x474 & ~x513;
assign c5185 =  x17 &  x52 &  x65 &  x317 &  x433 &  x476 &  x533 &  x709 &  x893 &  x920 &  x1001 &  x1007 &  x1046 &  x1049 &  x1091 & ~x228 & ~x897 & ~x1062 & ~x1101;
assign c5187 =  x107 &  x161 &  x206 &  x208 &  x233 &  x247 &  x292 &  x341 &  x422 &  x440 &  x482 &  x506 &  x545 &  x557 &  x653 &  x665 &  x761 &  x764 &  x872 &  x971 &  x980 &  x989 &  x995 &  x1034 &  x1067 &  x1085 &  x1097 &  x1115 &  x1118 & ~x81 & ~x381 & ~x939 & ~x1095;
assign c5189 = ~x33 & ~x249 & ~x411 & ~x534 & ~x594 & ~x1056 & ~x1095;
assign c5191 =  x82 &  x121 &  x160 &  x238 &  x539 &  x721 &  x733 &  x856 & ~x975 & ~x1062;
assign c5193 =  x112 &  x223 &  x262 &  x385 &  x403 &  x706 &  x1063 & ~x312 & ~x1071 & ~x1110;
assign c5195 =  x304 &  x310 &  x343 &  x349 &  x1069 & ~x84 & ~x474 & ~x894;
assign c5197 =  x38 &  x82 &  x143 &  x679 &  x757 &  x796 & ~x705 & ~x900 & ~x939 & ~x1017 & ~x1098;
assign c5199 =  x82 &  x185 &  x199 &  x739 &  x838 & ~x588 & ~x939 & ~x978;
assign c5201 =  x77 &  x125 &  x164 &  x191 &  x208 &  x230 &  x242 &  x310 &  x461 &  x542 &  x605 &  x677 &  x707 &  x835 &  x874 &  x884 &  x992 &  x1013 &  x1025 &  x1061 &  x1073 &  x1076 & ~x978 & ~x1017;
assign c5203 =  x145 &  x343 &  x364 &  x442 &  x487 &  x520 &  x598 &  x1024 & ~x282;
assign c5205 = ~x228 & ~x927 & ~x960 & ~x969 & ~x999 & ~x1038 & ~x1050 & ~x1083;
assign c5207 =  x531 &  x570 &  x745 & ~x430 & ~x540;
assign c5209 =  x4 &  x199 &  x238 &  x248 &  x355 &  x433 &  x511 &  x590 &  x641 &  x677 &  x866 &  x1010 &  x1061 & ~x669;
assign c5211 =  x223 &  x262 &  x346 &  x370 &  x463 &  x520 &  x598 &  x946 & ~x1083;
assign c5213 =  x26 &  x32 &  x278 &  x284 &  x344 &  x353 &  x395 &  x512 &  x527 &  x991 &  x1016 &  x1029 &  x1030 &  x1061 &  x1076 & ~x804 & ~x915 & ~x921 & ~x960 & ~x999 & ~x1038 & ~x1077;
assign c5215 =  x226 &  x403 &  x487 &  x493 &  x742 & ~x618;
assign c5217 =  x41 &  x59 &  x65 &  x68 &  x71 &  x77 &  x82 &  x83 &  x119 &  x121 &  x128 &  x160 &  x167 &  x203 &  x209 &  x233 &  x239 &  x245 &  x266 &  x293 &  x296 &  x314 &  x350 &  x353 &  x362 &  x383 &  x407 &  x422 &  x437 &  x443 &  x458 &  x494 &  x518 &  x521 &  x533 &  x563 &  x644 &  x647 &  x662 &  x698 &  x740 &  x743 &  x773 &  x800 &  x812 &  x818 &  x875 &  x926 &  x935 &  x953 &  x971 &  x1013 &  x1025 &  x1037 &  x1040 &  x1064 &  x1079 &  x1112 & ~x435 & ~x459 & ~x474 & ~x513 & ~x1011;
assign c5219 =  x913 & ~x688 & ~x822;
assign c5221 =  x262 &  x263 &  x290 &  x874 &  x913 &  x917 &  x1048 &  x1112 &  x1118 & ~x531 & ~x648 & ~x900 & ~x939 & ~x978 & ~x1017 & ~x1095;
assign c5223 =  x121 & ~x382 & ~x978;
assign c5225 =  x183 & ~x240 & ~x282 & ~x474;
assign c5227 =  x343 &  x349 &  x376 &  x517 &  x556 &  x635 &  x779 &  x842 & ~x606;
assign c5229 =  x29 &  x98 &  x283 &  x785 &  x813 &  x986 &  x1007 & ~x687 & ~x978;
assign c5231 =  x52 &  x954 & ~x138 & ~x177 & ~x411;
assign c5233 =  x226 & ~x313 & ~x450 & ~x684 & ~x927;
assign c5235 =  x625 & ~x234 & ~x333 & ~x384 & ~x552 & ~x708;
assign c5237 =  x238 &  x391 &  x472 & ~x543 & ~x544 & ~x583;
assign c5239 =  x11 &  x640 &  x718 &  x757 &  x796 &  x1094 & ~x570 & ~x687 & ~x900 & ~x939 & ~x978 & ~x1056 & ~x1095;
assign c5241 =  x112 &  x223 &  x335 &  x364 &  x403 &  x442 &  x478 &  x481 &  x524 &  x784 &  x959 & ~x390 & ~x1011;
assign c5243 =  x52 &  x86 &  x316 &  x452 &  x865 &  x911 &  x1045 &  x1123 & ~x267;
assign c5245 =  x88 &  x166 &  x205 &  x259 &  x442 &  x755 &  x820 & ~x474;
assign c5247 =  x62 &  x65 &  x251 &  x253 &  x254 &  x350 &  x368 &  x386 &  x472 &  x511 &  x521 &  x595 &  x634 &  x800 &  x815 &  x1085 & ~x204;
assign c5249 =  x140 &  x605 &  x863 &  x1082 & ~x60 & ~x93 & ~x99 & ~x132 & ~x171 & ~x345 & ~x435 & ~x513 & ~x519 & ~x756;
assign c5251 =  x5 &  x35 &  x41 &  x50 &  x65 &  x128 &  x134 &  x179 &  x193 &  x230 &  x233 &  x236 &  x239 &  x247 &  x253 &  x286 &  x344 &  x359 &  x404 &  x431 &  x472 &  x506 &  x509 &  x511 &  x515 &  x539 &  x629 &  x656 &  x659 &  x737 &  x851 &  x956 &  x1001 &  x1007 &  x1025 &  x1100 &  x1108;
assign c5253 = ~x72 & ~x823 & ~x862 & ~x1095;
assign c5255 =  x74 &  x170 &  x179 &  x281 &  x697 &  x718 &  x755 &  x830 &  x971 & ~x706 & ~x745 & ~x784 & ~x978 & ~x1095;
assign c5257 =  x317 &  x364 &  x524 &  x628 &  x783 & ~x261 & ~x339 & ~x378;
assign c5259 =  x77 &  x167 &  x608 &  x617 &  x653 &  x706 &  x1024 &  x1063 &  x1091 & ~x352 & ~x540;
assign c5261 =  x82 &  x110 &  x121 &  x371 &  x506 &  x626 &  x629 & ~x202 & ~x333 & ~x372;
assign c5263 =  x8 &  x80 &  x113 &  x134 &  x136 &  x169 &  x175 &  x181 &  x215 &  x218 &  x275 &  x472 &  x569 &  x581 &  x587 &  x623 &  x629 &  x632 &  x638 &  x692 &  x758 &  x761 &  x806 &  x818 &  x857 &  x872 &  x890 &  x911 &  x950 &  x1031 &  x1061 &  x1082 & ~x78 & ~x117 & ~x234 & ~x1092;
assign c5265 =  x89 &  x173 &  x674 & ~x123 & ~x177 & ~x216 & ~x217 & ~x627 & ~x666 & ~x822 & ~x939;
assign c5267 =  x43 &  x238 &  x796 &  x835 &  x874 & ~x1092;
assign c5269 =  x370 & ~x456 & ~x612 & ~x651 & ~x652 & ~x691 & ~x924;
assign c5271 =  x65 &  x82 &  x238 &  x689 &  x991 &  x1000 &  x1030 &  x1114 & ~x309;
assign c5273 =  x388 &  x487 &  x565 & ~x430 & ~x469 & ~x547 & ~x873;
assign c5275 =  x874 & ~x687 & ~x765 & ~x1095;
assign c5277 = ~x216 & ~x267 & ~x417 & ~x435 & ~x561 & ~x1081;
assign c5279 =  x112 &  x346 &  x427 &  x481 &  x559 &  x598 &  x1063 & ~x390 & ~x1005;
assign c5281 =  x292 &  x299 &  x364 &  x638 &  x668 &  x875 &  x959 &  x965 &  x974 & ~x384 & ~x1095;
assign c5283 =  x559 &  x570 &  x822 & ~x117;
assign c5285 =  x349 &  x1069 &  x1108 &  x1124 & ~x1032 & ~x1077;
assign c5287 =  x322 &  x463 &  x598 &  x697 &  x796 & ~x123;
assign c5289 =  x2 &  x5 &  x77 &  x82 &  x121 &  x160 &  x199 &  x344 &  x542 &  x590 &  x757 &  x796 &  x835 &  x878 &  x889 &  x935 &  x1043 &  x1085 &  x1088 & ~x141 & ~x330 & ~x369;
assign c5291 =  x265 &  x913 &  x991 & ~x492 & ~x687 & ~x1017 & ~x1056 & ~x1095;
assign c5293 =  x35 &  x95 &  x199 &  x206 &  x227 &  x332 &  x419 &  x527 &  x542 &  x554 &  x584 &  x689 &  x731 &  x998 &  x1106 & ~x543 & ~x582 & ~x939 & ~x1053;
assign c5295 =  x193 &  x226 &  x232 &  x262 &  x265 &  x349 &  x364 &  x667 &  x854 &  x1024 &  x1063 &  x1064 & ~x120;
assign c5297 =  x175 &  x316 &  x1124 & ~x78 & ~x118;
assign c5299 =  x32 &  x47 &  x50 &  x68 &  x71 &  x77 &  x137 &  x149 &  x155 &  x170 &  x197 &  x209 &  x257 &  x263 &  x275 &  x277 &  x281 &  x287 &  x296 &  x316 &  x317 &  x329 &  x341 &  x356 &  x359 &  x398 &  x430 &  x434 &  x443 &  x446 &  x449 &  x458 &  x469 &  x470 &  x485 &  x506 &  x509 &  x530 &  x539 &  x551 &  x575 &  x590 &  x596 &  x611 &  x644 &  x659 &  x662 &  x677 &  x758 &  x800 &  x809 &  x815 &  x842 &  x881 &  x884 &  x887 &  x899 &  x902 &  x938 &  x947 &  x956 &  x962 &  x968 &  x986 &  x1007 &  x1010 &  x1034 &  x1058 &  x1073 &  x1088 &  x1097 &  x1109 &  x1127 & ~x156 & ~x474 & ~x513;
assign c60 =  x2 &  x11 &  x23 &  x26 &  x35 &  x47 &  x68 &  x74 &  x77 &  x89 &  x101 &  x110 &  x131 &  x137 &  x149 &  x152 &  x176 &  x194 &  x197 &  x209 &  x242 &  x269 &  x284 &  x290 &  x293 &  x296 &  x299 &  x302 &  x308 &  x326 &  x329 &  x374 &  x380 &  x386 &  x389 &  x395 &  x398 &  x401 &  x404 &  x416 &  x419 &  x434 &  x446 &  x449 &  x464 &  x473 &  x476 &  x482 &  x491 &  x500 &  x506 &  x509 &  x515 &  x536 &  x539 &  x542 &  x551 &  x563 &  x566 &  x569 &  x572 &  x581 &  x602 &  x623 &  x644 &  x656 &  x659 &  x677 &  x680 &  x683 &  x695 &  x698 &  x707 &  x716 &  x722 &  x731 &  x746 &  x749 &  x758 &  x764 &  x767 &  x785 &  x803 &  x812 &  x818 &  x821 &  x830 &  x833 &  x848 &  x851 &  x860 &  x866 &  x869 &  x881 &  x890 &  x893 &  x899 &  x902 &  x932 &  x944 &  x974 &  x977 &  x983 &  x986 &  x989 &  x998 &  x1001 &  x1013 &  x1016 &  x1022 &  x1049 &  x1064 &  x1079 &  x1085 &  x1091 &  x1103 &  x1106 & ~x399 & ~x480 & ~x520 & ~x552 & ~x558 & ~x559 & ~x591 & ~x597 & ~x627 & ~x885;
assign c62 =  x32 &  x77 &  x101 &  x278 &  x284 &  x353 &  x374 &  x397 &  x398 &  x415 &  x431 &  x454 &  x466 &  x482 &  x491 &  x493 &  x532 &  x536 &  x563 &  x571 &  x650 &  x667 &  x706 &  x722 &  x737 &  x745 &  x784 &  x823 &  x839 &  x845 &  x860 &  x862 &  x878 &  x940 &  x962 &  x979 &  x992 &  x1055 &  x1057 &  x1079 & ~x273 & ~x312 & ~x718 & ~x756;
assign c64 =  x56 &  x80 &  x89 &  x92 &  x98 &  x106 &  x122 &  x146 &  x167 &  x176 &  x179 &  x197 &  x239 &  x257 &  x269 &  x380 &  x395 &  x398 &  x411 &  x419 &  x451 &  x482 &  x560 &  x563 &  x566 &  x569 &  x587 &  x593 &  x707 &  x728 &  x746 &  x770 &  x779 &  x809 &  x823 &  x881 &  x886 &  x899 &  x901 &  x902 &  x920 &  x940 &  x941 &  x953 &  x998 &  x1046 &  x1079 &  x1085 &  x1127 & ~x444;
assign c66 =  x14 &  x32 &  x35 &  x47 &  x83 &  x89 &  x101 &  x116 &  x128 &  x164 &  x176 &  x203 &  x230 &  x239 &  x251 &  x278 &  x284 &  x287 &  x302 &  x308 &  x326 &  x337 &  x347 &  x350 &  x368 &  x374 &  x376 &  x380 &  x388 &  x395 &  x413 &  x415 &  x416 &  x427 &  x431 &  x454 &  x458 &  x466 &  x482 &  x493 &  x518 &  x532 &  x536 &  x548 &  x551 &  x563 &  x566 &  x571 &  x575 &  x587 &  x610 &  x623 &  x641 &  x649 &  x650 &  x674 &  x680 &  x688 &  x692 &  x706 &  x713 &  x725 &  x734 &  x743 &  x745 &  x746 &  x764 &  x770 &  x788 &  x823 &  x827 &  x830 &  x848 &  x851 &  x860 &  x866 &  x902 &  x908 &  x923 &  x929 &  x947 &  x953 &  x968 &  x977 &  x979 &  x980 &  x989 &  x998 &  x1016 &  x1019 &  x1022 &  x1043 &  x1064 &  x1079 & ~x312 & ~x678 & ~x714 & ~x717;
assign c68 =  x65 &  x178 &  x217 &  x256 &  x268 &  x287 &  x295 &  x361 &  x400 &  x439 &  x532 &  x571 &  x587 &  x610 &  x724 &  x755 &  x801 &  x802 &  x829 &  x841 &  x879 &  x880;
assign c610 =  x83 &  x101 &  x140 &  x149 &  x167 &  x197 &  x284 &  x431 &  x466 &  x491 &  x503 &  x526 &  x538 &  x545 &  x566 &  x587 &  x605 &  x644 &  x677 &  x722 &  x764 &  x848 &  x866 &  x869 &  x884 &  x968 &  x995 &  x998 &  x1094 &  x1121 &  x1124 & ~x321 & ~x438 & ~x468 & ~x516 & ~x555 & ~x633 & ~x756 & ~x792 & ~x831 & ~x987;
assign c612 =  x14 &  x23 &  x44 &  x56 &  x65 &  x83 &  x89 &  x140 &  x149 &  x176 &  x194 &  x209 &  x221 &  x236 &  x242 &  x248 &  x257 &  x263 &  x269 &  x275 &  x284 &  x287 &  x317 &  x344 &  x359 &  x395 &  x404 &  x413 &  x434 &  x446 &  x464 &  x476 &  x479 &  x488 &  x491 &  x497 &  x500 &  x518 &  x521 &  x551 &  x563 &  x566 &  x569 &  x581 &  x587 &  x590 &  x611 &  x620 &  x632 &  x650 &  x653 &  x680 &  x688 &  x698 &  x716 &  x722 &  x734 &  x782 &  x799 &  x803 &  x824 &  x833 &  x838 &  x854 &  x866 &  x877 &  x878 &  x884 &  x893 &  x908 &  x923 &  x938 &  x950 &  x956 &  x968 &  x971 &  x973 &  x980 &  x986 &  x992 &  x998 &  x1016 &  x1022 &  x1025 &  x1031 &  x1040 &  x1051 &  x1052 &  x1055 &  x1067 &  x1072 &  x1082 &  x1094 &  x1097 &  x1100 &  x1111 & ~x9 & ~x48 & ~x87 & ~x165 & ~x321 & ~x483;
assign c614 =  x22 &  x100 &  x118 &  x151 &  x190 &  x256 &  x268 &  x295 &  x301 &  x307 &  x346 &  x365 &  x419 &  x535 &  x572 &  x697 &  x769 &  x808 &  x841 &  x890 &  x968 &  x1079 & ~x24 & ~x408;
assign c616 =  x7 &  x35 &  x53 &  x76 &  x77 &  x89 &  x104 &  x110 &  x116 &  x149 &  x197 &  x224 &  x239 &  x257 &  x266 &  x278 &  x317 &  x347 &  x368 &  x395 &  x419 &  x437 &  x443 &  x464 &  x491 &  x497 &  x545 &  x563 &  x569 &  x584 &  x605 &  x611 &  x650 &  x653 &  x668 &  x698 &  x731 &  x737 &  x740 &  x743 &  x826 &  x830 &  x833 &  x845 &  x875 &  x881 &  x902 &  x920 &  x923 &  x929 &  x938 &  x943 &  x950 &  x955 &  x961 &  x986 &  x992 &  x1001 &  x1019 &  x1022 &  x1033 &  x1043 &  x1046 &  x1049 &  x1055 &  x1082 &  x1085 &  x1115 & ~x249 & ~x288 & ~x327 & ~x405 & ~x444 & ~x483 & ~x852 & ~x891 & ~x930;
assign c618 =  x77 &  x104 &  x110 &  x128 &  x142 &  x149 &  x152 &  x155 &  x271 &  x284 &  x302 &  x317 &  x383 &  x395 &  x437 &  x482 &  x491 &  x503 &  x551 &  x563 &  x566 &  x571 &  x587 &  x602 &  x688 &  x698 &  x710 &  x734 &  x743 &  x749 &  x760 &  x788 &  x799 &  x824 &  x863 &  x932 &  x947 &  x959 &  x983 &  x986 &  x1001 &  x1031 &  x1033 &  x1072 &  x1079 & ~x402 & ~x483 & ~x522 & ~x939;
assign c620 =  x23 &  x32 &  x35 &  x71 &  x83 &  x92 &  x110 &  x119 &  x122 &  x128 &  x137 &  x146 &  x167 &  x176 &  x218 &  x221 &  x269 &  x284 &  x287 &  x311 &  x350 &  x374 &  x398 &  x407 &  x431 &  x437 &  x452 &  x491 &  x515 &  x518 &  x536 &  x542 &  x551 &  x554 &  x563 &  x587 &  x593 &  x604 &  x643 &  x647 &  x650 &  x659 &  x688 &  x692 &  x694 &  x721 &  x722 &  x760 &  x770 &  x773 &  x785 &  x806 &  x838 &  x839 &  x866 &  x884 &  x902 &  x929 &  x944 &  x956 &  x959 &  x973 &  x995 &  x1001 &  x1028 &  x1040 &  x1046 &  x1064 &  x1079 &  x1088 &  x1118 &  x1124 & ~x285 & ~x321 & ~x360 & ~x399 & ~x402 & ~x438 & ~x441 & ~x477 & ~x516 & ~x555;
assign c622 =  x2 &  x11 &  x14 &  x23 &  x35 &  x38 &  x41 &  x44 &  x71 &  x77 &  x80 &  x83 &  x89 &  x95 &  x98 &  x110 &  x113 &  x125 &  x128 &  x137 &  x143 &  x146 &  x149 &  x152 &  x167 &  x170 &  x173 &  x188 &  x191 &  x203 &  x209 &  x215 &  x224 &  x227 &  x245 &  x251 &  x254 &  x269 &  x278 &  x281 &  x284 &  x290 &  x305 &  x308 &  x314 &  x326 &  x332 &  x347 &  x353 &  x359 &  x365 &  x368 &  x371 &  x377 &  x380 &  x383 &  x386 &  x389 &  x395 &  x422 &  x434 &  x437 &  x440 &  x449 &  x467 &  x473 &  x500 &  x506 &  x515 &  x521 &  x533 &  x536 &  x542 &  x545 &  x548 &  x554 &  x563 &  x578 &  x581 &  x584 &  x590 &  x593 &  x599 &  x608 &  x632 &  x635 &  x641 &  x644 &  x656 &  x659 &  x680 &  x689 &  x692 &  x698 &  x704 &  x740 &  x743 &  x746 &  x755 &  x758 &  x761 &  x764 &  x773 &  x782 &  x785 &  x791 &  x803 &  x809 &  x812 &  x815 &  x818 &  x833 &  x836 &  x845 &  x860 &  x869 &  x875 &  x884 &  x890 &  x893 &  x899 &  x905 &  x908 &  x920 &  x923 &  x941 &  x950 &  x956 &  x959 &  x962 &  x965 &  x968 &  x980 &  x986 &  x989 &  x992 &  x1007 &  x1013 &  x1025 &  x1031 &  x1034 &  x1043 &  x1046 &  x1049 &  x1058 &  x1070 &  x1079 &  x1082 &  x1085 &  x1091 &  x1100 &  x1103 &  x1106 &  x1109 &  x1112 &  x1121 &  x1124 & ~x399 & ~x438 & ~x516 & ~x637 & ~x675 & ~x678 & ~x714 & ~x717 & ~x753 & ~x756 & ~x792 & ~x831 & ~x870 & ~x909;
assign c624 =  x77 &  x101 &  x116 &  x137 &  x170 &  x262 &  x308 &  x326 &  x395 &  x419 &  x491 &  x493 &  x503 &  x532 &  x536 &  x560 &  x563 &  x569 &  x571 &  x587 &  x605 &  x610 &  x649 &  x653 &  x680 &  x688 &  x692 &  x731 &  x743 &  x752 &  x764 &  x788 &  x844 &  x845 &  x902 &  x920 &  x929 &  x959 &  x1001 &  x1019 &  x1051 &  x1055 &  x1064 &  x1078 &  x1079 &  x1100 & ~x162 & ~x240 & ~x318 & ~x369;
assign c626 =  x23 &  x32 &  x35 &  x50 &  x53 &  x86 &  x116 &  x128 &  x140 &  x149 &  x152 &  x158 &  x163 &  x164 &  x170 &  x194 &  x197 &  x202 &  x203 &  x227 &  x239 &  x241 &  x248 &  x257 &  x269 &  x284 &  x287 &  x302 &  x308 &  x311 &  x329 &  x353 &  x377 &  x389 &  x392 &  x395 &  x404 &  x431 &  x434 &  x449 &  x452 &  x479 &  x482 &  x485 &  x491 &  x494 &  x500 &  x503 &  x518 &  x575 &  x590 &  x602 &  x614 &  x632 &  x635 &  x644 &  x659 &  x677 &  x686 &  x689 &  x707 &  x716 &  x725 &  x728 &  x737 &  x743 &  x761 &  x764 &  x779 &  x788 &  x800 &  x809 &  x827 &  x839 &  x845 &  x860 &  x865 &  x866 &  x869 &  x872 &  x881 &  x893 &  x899 &  x904 &  x920 &  x944 &  x953 &  x977 &  x992 &  x995 &  x1001 &  x1022 &  x1031 &  x1034 &  x1040 &  x1043 &  x1049 &  x1055 &  x1064 &  x1079 &  x1100 &  x1109 &  x1112 &  x1130 & ~x213 & ~x246 & ~x285 & ~x402 & ~x441 & ~x480 & ~x597 & ~x666 & ~x978;
assign c628 =  x26 &  x55 &  x56 &  x100 &  x122 &  x134 &  x151 &  x155 &  x170 &  x172 &  x190 &  x217 &  x221 &  x229 &  x245 &  x256 &  x272 &  x344 &  x347 &  x350 &  x359 &  x368 &  x385 &  x392 &  x422 &  x446 &  x476 &  x479 &  x482 &  x491 &  x494 &  x500 &  x518 &  x536 &  x560 &  x571 &  x572 &  x587 &  x596 &  x608 &  x610 &  x659 &  x719 &  x769 &  x830 &  x841 &  x848 &  x863 &  x908 &  x932 &  x938 &  x956 &  x971 &  x1001 &  x1049 & ~x162 & ~x246 & ~x285 & ~x363 & ~x864;
assign c630 =  x100 &  x139 &  x191 &  x217 &  x256 &  x295 &  x302 &  x308 &  x334 &  x392 &  x398 &  x412 &  x451 &  x500 &  x536 &  x563 &  x688 &  x692 &  x719 &  x721 &  x725 &  x746 &  x760 &  x763 &  x799 &  x802 &  x841 &  x848 &  x853 &  x872 &  x902 &  x944 &  x947 &  x986 &  x1016 &  x1022 &  x1100 & ~x84 & ~x123 & ~x396 & ~x552;
assign c632 =  x8 &  x11 &  x14 &  x23 &  x26 &  x32 &  x47 &  x71 &  x74 &  x80 &  x83 &  x89 &  x101 &  x107 &  x110 &  x116 &  x122 &  x128 &  x137 &  x146 &  x173 &  x182 &  x197 &  x200 &  x209 &  x218 &  x230 &  x233 &  x236 &  x239 &  x242 &  x266 &  x269 &  x278 &  x281 &  x284 &  x290 &  x293 &  x299 &  x308 &  x314 &  x320 &  x338 &  x344 &  x368 &  x371 &  x380 &  x386 &  x389 &  x392 &  x398 &  x404 &  x413 &  x422 &  x440 &  x452 &  x461 &  x467 &  x482 &  x485 &  x503 &  x509 &  x518 &  x530 &  x533 &  x536 &  x539 &  x542 &  x548 &  x560 &  x563 &  x566 &  x575 &  x578 &  x587 &  x602 &  x614 &  x620 &  x623 &  x632 &  x635 &  x647 &  x650 &  x656 &  x659 &  x668 &  x677 &  x680 &  x686 &  x689 &  x692 &  x695 &  x698 &  x707 &  x710 &  x716 &  x719 &  x722 &  x725 &  x731 &  x734 &  x743 &  x746 &  x755 &  x764 &  x767 &  x788 &  x809 &  x812 &  x818 &  x827 &  x833 &  x845 &  x851 &  x863 &  x881 &  x887 &  x890 &  x896 &  x902 &  x911 &  x920 &  x923 &  x926 &  x932 &  x935 &  x944 &  x965 &  x980 &  x986 &  x992 &  x995 &  x1001 &  x1019 &  x1022 &  x1028 &  x1034 &  x1040 &  x1046 &  x1055 &  x1058 &  x1082 &  x1088 &  x1091 &  x1103 &  x1109 &  x1112 &  x1115 &  x1118 &  x1124 &  x1127 & ~x432 & ~x438 & ~x471 & ~x477 & ~x510 & ~x516 & ~x549 & ~x636 & ~x714 & ~x747 & ~x753 & ~x792 & ~x909 & ~x942 & ~x948 & ~x987 & ~x1020 & ~x1026 & ~x1059 & ~x1116;
assign c634 =  x17 &  x29 &  x32 &  x44 &  x83 &  x95 &  x98 &  x140 &  x161 &  x167 &  x176 &  x305 &  x308 &  x323 &  x344 &  x374 &  x383 &  x431 &  x458 &  x461 &  x473 &  x493 &  x497 &  x509 &  x524 &  x532 &  x571 &  x584 &  x605 &  x622 &  x646 &  x653 &  x656 &  x661 &  x665 &  x692 &  x694 &  x698 &  x707 &  x725 &  x767 &  x775 &  x800 &  x806 &  x814 &  x824 &  x851 &  x853 &  x902 &  x917 &  x953 &  x1001 &  x1016 &  x1031 &  x1040 &  x1055 &  x1085 &  x1088 &  x1130 & ~x432 & ~x438 & ~x477 & ~x510 & ~x516 & ~x549 & ~x555 & ~x588 & ~x594 & ~x627 & ~x633 & ~x672;
assign c636 =  x41 &  x100 &  x178 &  x205 &  x242 &  x256 &  x262 &  x295 &  x395 &  x412 &  x437 &  x451 &  x529 &  x607 &  x685 &  x724 &  x760 &  x775 &  x799 &  x802 &  x814 &  x848 &  x877 &  x947 &  x1001 &  x1051;
assign c638 =  x68 &  x95 &  x122 &  x194 &  x218 &  x221 &  x311 &  x521 &  x632 &  x638 &  x650 &  x668 &  x689 &  x776 &  x785 &  x830 &  x848 &  x851 &  x908 &  x917 &  x953 &  x1055 & ~x52 & ~x93 & ~x132 & ~x171 & ~x210 & ~x264 & ~x588 & ~x627 & ~x664 & ~x666;
assign c640 =  x14 &  x32 &  x53 &  x74 &  x77 &  x83 &  x92 &  x101 &  x122 &  x143 &  x164 &  x167 &  x173 &  x182 &  x188 &  x194 &  x197 &  x203 &  x221 &  x224 &  x230 &  x236 &  x242 &  x257 &  x269 &  x272 &  x284 &  x296 &  x299 &  x302 &  x308 &  x335 &  x353 &  x374 &  x377 &  x380 &  x386 &  x388 &  x392 &  x395 &  x407 &  x416 &  x427 &  x431 &  x452 &  x455 &  x461 &  x466 &  x473 &  x479 &  x482 &  x491 &  x497 &  x503 &  x505 &  x530 &  x536 &  x544 &  x551 &  x554 &  x557 &  x569 &  x575 &  x583 &  x587 &  x602 &  x620 &  x622 &  x626 &  x638 &  x644 &  x650 &  x661 &  x668 &  x677 &  x680 &  x692 &  x695 &  x698 &  x700 &  x707 &  x722 &  x725 &  x737 &  x739 &  x740 &  x743 &  x746 &  x761 &  x770 &  x778 &  x785 &  x788 &  x794 &  x800 &  x806 &  x809 &  x812 &  x827 &  x833 &  x839 &  x845 &  x848 &  x851 &  x862 &  x869 &  x875 &  x884 &  x901 &  x902 &  x905 &  x917 &  x929 &  x934 &  x940 &  x944 &  x947 &  x953 &  x962 &  x968 &  x986 &  x992 &  x995 &  x1016 &  x1022 &  x1034 &  x1040 &  x1046 &  x1055 &  x1064 &  x1076 &  x1079 &  x1088 &  x1091 &  x1103 &  x1127 & ~x0 & ~x39 & ~x78 & ~x117 & ~x234 & ~x273 & ~x405 & ~x1008;
assign c642 =  x23 &  x53 &  x146 &  x194 &  x248 &  x266 &  x284 &  x302 &  x322 &  x323 &  x335 &  x361 &  x368 &  x371 &  x422 &  x458 &  x461 &  x464 &  x476 &  x482 &  x512 &  x524 &  x527 &  x529 &  x532 &  x560 &  x568 &  x571 &  x584 &  x587 &  x596 &  x623 &  x685 &  x695 &  x721 &  x724 &  x725 &  x755 &  x760 &  x763 &  x767 &  x769 &  x770 &  x797 &  x814 &  x818 &  x833 &  x842 &  x853 &  x854 &  x869 &  x871 &  x874 &  x883 &  x886 &  x938 &  x949 &  x955 &  x980 &  x1001 &  x1027 &  x1124 & ~x549 & ~x588 & ~x627 & ~x744;
assign c644 =  x2 &  x23 &  x32 &  x44 &  x53 &  x56 &  x71 &  x77 &  x80 &  x83 &  x86 &  x89 &  x92 &  x101 &  x110 &  x116 &  x122 &  x128 &  x137 &  x149 &  x164 &  x167 &  x176 &  x194 &  x197 &  x203 &  x221 &  x227 &  x239 &  x242 &  x257 &  x269 &  x278 &  x284 &  x302 &  x308 &  x311 &  x326 &  x335 &  x347 &  x350 &  x371 &  x374 &  x380 &  x386 &  x388 &  x395 &  x398 &  x407 &  x416 &  x419 &  x431 &  x434 &  x437 &  x452 &  x461 &  x473 &  x479 &  x482 &  x485 &  x491 &  x494 &  x500 &  x503 &  x506 &  x515 &  x518 &  x536 &  x548 &  x554 &  x563 &  x566 &  x569 &  x575 &  x578 &  x584 &  x587 &  x590 &  x602 &  x605 &  x611 &  x620 &  x623 &  x632 &  x635 &  x646 &  x647 &  x650 &  x659 &  x668 &  x677 &  x680 &  x686 &  x692 &  x707 &  x722 &  x725 &  x728 &  x731 &  x737 &  x743 &  x749 &  x755 &  x761 &  x764 &  x770 &  x779 &  x785 &  x788 &  x800 &  x824 &  x830 &  x839 &  x845 &  x848 &  x851 &  x860 &  x866 &  x869 &  x881 &  x884 &  x893 &  x899 &  x905 &  x920 &  x923 &  x926 &  x929 &  x935 &  x944 &  x953 &  x959 &  x968 &  x986 &  x989 &  x992 &  x995 &  x998 &  x1001 &  x1004 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1040 &  x1043 &  x1049 &  x1055 &  x1064 &  x1079 &  x1082 &  x1085 &  x1097 &  x1103 &  x1115 &  x1124 &  x1127 &  x1130 & ~x234 & ~x273 & ~x312 & ~x366 & ~x444 & ~x483 & ~x522 & ~x525 & ~x561 & ~x564;
assign c646 =  x71 &  x77 &  x83 &  x146 &  x203 &  x209 &  x221 &  x239 &  x278 &  x284 &  x302 &  x326 &  x374 &  x395 &  x404 &  x419 &  x452 &  x482 &  x491 &  x500 &  x515 &  x518 &  x548 &  x563 &  x569 &  x587 &  x620 &  x668 &  x677 &  x680 &  x773 &  x779 &  x800 &  x824 &  x833 &  x848 &  x851 &  x902 &  x920 &  x929 &  x947 &  x968 &  x1001 &  x1016 &  x1022 &  x1028 &  x1031 &  x1043 &  x1055 &  x1079 &  x1088 &  x1097 &  x1103 &  x1106 & ~x132 & ~x162 & ~x171 & ~x249 & ~x288 & ~x324 & ~x363 & ~x396 & ~x402 & ~x435 & ~x441 & ~x480 & ~x597 & ~x636 & ~x795 & ~x834 & ~x900;
assign c648 =  x2 &  x23 &  x53 &  x65 &  x89 &  x101 &  x113 &  x125 &  x137 &  x155 &  x167 &  x185 &  x203 &  x209 &  x215 &  x218 &  x242 &  x257 &  x263 &  x284 &  x296 &  x299 &  x308 &  x320 &  x332 &  x356 &  x377 &  x386 &  x395 &  x416 &  x431 &  x449 &  x455 &  x466 &  x476 &  x491 &  x506 &  x544 &  x548 &  x551 &  x554 &  x572 &  x581 &  x596 &  x605 &  x608 &  x617 &  x622 &  x647 &  x677 &  x680 &  x686 &  x698 &  x710 &  x731 &  x761 &  x791 &  x824 &  x833 &  x839 &  x848 &  x863 &  x866 &  x896 &  x926 &  x956 &  x962 &  x965 &  x980 &  x998 &  x1007 &  x1016 &  x1022 &  x1034 &  x1049 &  x1070 &  x1073 &  x1079 &  x1103 &  x1112 &  x1118 & ~x3 & ~x39 & ~x60 & ~x93 & ~x132 & ~x171 & ~x210 & ~x327 & ~x366 & ~x483 & ~x522 & ~x561 & ~x756 & ~x834 & ~x873;
assign c650 =  x2 &  x11 &  x14 &  x23 &  x41 &  x44 &  x47 &  x53 &  x65 &  x77 &  x83 &  x89 &  x92 &  x101 &  x104 &  x110 &  x113 &  x119 &  x122 &  x125 &  x128 &  x149 &  x164 &  x166 &  x167 &  x176 &  x188 &  x194 &  x197 &  x203 &  x206 &  x209 &  x215 &  x224 &  x239 &  x248 &  x269 &  x284 &  x302 &  x308 &  x323 &  x326 &  x343 &  x350 &  x365 &  x371 &  x380 &  x382 &  x388 &  x389 &  x392 &  x395 &  x398 &  x404 &  x407 &  x419 &  x421 &  x425 &  x427 &  x428 &  x431 &  x434 &  x449 &  x461 &  x466 &  x476 &  x479 &  x482 &  x491 &  x494 &  x500 &  x503 &  x518 &  x533 &  x536 &  x557 &  x563 &  x566 &  x569 &  x581 &  x590 &  x602 &  x605 &  x620 &  x623 &  x644 &  x650 &  x659 &  x677 &  x680 &  x692 &  x707 &  x713 &  x719 &  x722 &  x725 &  x728 &  x743 &  x746 &  x764 &  x767 &  x770 &  x779 &  x794 &  x806 &  x809 &  x812 &  x824 &  x839 &  x845 &  x848 &  x851 &  x860 &  x866 &  x869 &  x881 &  x884 &  x899 &  x902 &  x911 &  x917 &  x920 &  x944 &  x947 &  x953 &  x959 &  x968 &  x971 &  x980 &  x983 &  x986 &  x992 &  x995 &  x1001 &  x1007 &  x1016 &  x1019 &  x1022 &  x1025 &  x1028 &  x1031 &  x1046 &  x1049 &  x1052 &  x1055 &  x1061 &  x1064 &  x1070 &  x1072 &  x1079 &  x1103 &  x1106 &  x1111 &  x1124 & ~x444 & ~x483 & ~x975;
assign c652 =  x2 &  x5 &  x26 &  x35 &  x47 &  x50 &  x77 &  x89 &  x101 &  x122 &  x125 &  x128 &  x131 &  x134 &  x149 &  x152 &  x155 &  x194 &  x197 &  x209 &  x212 &  x221 &  x224 &  x227 &  x242 &  x251 &  x257 &  x260 &  x272 &  x302 &  x326 &  x353 &  x374 &  x377 &  x395 &  x398 &  x410 &  x425 &  x431 &  x446 &  x455 &  x473 &  x479 &  x485 &  x500 &  x503 &  x518 &  x527 &  x530 &  x536 &  x551 &  x554 &  x560 &  x566 &  x575 &  x581 &  x587 &  x590 &  x599 &  x602 &  x605 &  x614 &  x617 &  x620 &  x623 &  x638 &  x644 &  x650 &  x659 &  x673 &  x674 &  x680 &  x689 &  x692 &  x707 &  x728 &  x734 &  x743 &  x746 &  x749 &  x758 &  x767 &  x770 &  x773 &  x779 &  x782 &  x785 &  x788 &  x800 &  x824 &  x827 &  x830 &  x839 &  x860 &  x866 &  x869 &  x893 &  x902 &  x917 &  x944 &  x962 &  x965 &  x968 &  x974 &  x986 &  x995 &  x1001 &  x1016 &  x1031 &  x1034 &  x1064 &  x1067 &  x1118 & ~x438 & ~x477 & ~x516 & ~x747 & ~x915 & ~x942 & ~x1080 & ~x1083 & ~x1122;
assign c654 =  x200 &  x412 &  x436 &  x466 &  x475 &  x493 &  x515 &  x529 &  x530 &  x532 &  x535 &  x554 &  x568 &  x602 &  x845 &  x869 &  x959 &  x962 &  x968 &  x998 & ~x471 & ~x510 & ~x549 & ~x717 & ~x771 & ~x792 & ~x849;
assign c656 =  x20 &  x65 &  x92 &  x101 &  x146 &  x170 &  x194 &  x209 &  x215 &  x227 &  x263 &  x284 &  x329 &  x355 &  x392 &  x395 &  x398 &  x407 &  x425 &  x431 &  x434 &  x452 &  x464 &  x479 &  x500 &  x503 &  x524 &  x572 &  x638 &  x674 &  x680 &  x692 &  x725 &  x755 &  x776 &  x779 &  x806 &  x838 &  x851 &  x866 &  x881 &  x884 &  x914 &  x929 &  x967 &  x986 &  x1022 &  x1043 &  x1055 &  x1103 & ~x9 & ~x48 & ~x87 & ~x210 & ~x249 & ~x288 & ~x363 & ~x366 & ~x402 & ~x441 & ~x480 & ~x522 & ~x702;
assign c658 =  x5 &  x14 &  x32 &  x38 &  x47 &  x50 &  x53 &  x56 &  x65 &  x71 &  x74 &  x80 &  x83 &  x86 &  x89 &  x98 &  x104 &  x116 &  x122 &  x134 &  x137 &  x146 &  x149 &  x152 &  x176 &  x194 &  x200 &  x203 &  x209 &  x227 &  x236 &  x239 &  x263 &  x266 &  x284 &  x290 &  x308 &  x326 &  x329 &  x347 &  x374 &  x389 &  x392 &  x410 &  x416 &  x422 &  x431 &  x434 &  x452 &  x458 &  x466 &  x488 &  x494 &  x506 &  x518 &  x524 &  x539 &  x548 &  x554 &  x557 &  x563 &  x569 &  x572 &  x599 &  x605 &  x608 &  x614 &  x617 &  x623 &  x632 &  x644 &  x659 &  x667 &  x668 &  x677 &  x686 &  x692 &  x698 &  x706 &  x713 &  x719 &  x725 &  x731 &  x737 &  x740 &  x743 &  x755 &  x779 &  x785 &  x788 &  x794 &  x809 &  x821 &  x827 &  x830 &  x839 &  x845 &  x860 &  x869 &  x881 &  x884 &  x902 &  x920 &  x926 &  x935 &  x959 &  x965 &  x974 &  x979 &  x980 &  x986 &  x1001 &  x1016 &  x1022 &  x1034 &  x1040 &  x1046 &  x1049 &  x1055 &  x1058 &  x1061 &  x1067 &  x1076 &  x1079 &  x1085 &  x1091 &  x1097 &  x1112 &  x1118 &  x1127 & ~x312 & ~x393 & ~x597 & ~x636 & ~x675 & ~x714 & ~x732 & ~x771 & ~x810 & ~x831 & ~x870;
assign c660 =  x5 &  x8 &  x11 &  x20 &  x22 &  x32 &  x34 &  x41 &  x77 &  x80 &  x89 &  x101 &  x110 &  x112 &  x134 &  x139 &  x149 &  x176 &  x178 &  x194 &  x197 &  x203 &  x209 &  x217 &  x227 &  x239 &  x268 &  x284 &  x287 &  x295 &  x307 &  x308 &  x334 &  x337 &  x343 &  x346 &  x353 &  x376 &  x380 &  x385 &  x398 &  x401 &  x407 &  x415 &  x416 &  x419 &  x424 &  x463 &  x491 &  x493 &  x503 &  x532 &  x557 &  x566 &  x569 &  x571 &  x580 &  x590 &  x610 &  x619 &  x635 &  x641 &  x644 &  x650 &  x658 &  x677 &  x688 &  x692 &  x743 &  x770 &  x800 &  x809 &  x824 &  x830 &  x836 &  x839 &  x845 &  x848 &  x853 &  x860 &  x866 &  x881 &  x884 &  x892 &  x893 &  x899 &  x919 &  x920 &  x931 &  x944 &  x947 &  x958 &  x959 &  x965 &  x968 &  x980 &  x986 &  x992 &  x995 &  x997 &  x998 &  x1013 &  x1016 &  x1022 &  x1028 &  x1036 &  x1043 &  x1049 &  x1055 &  x1064 &  x1082 &  x1085 &  x1088 &  x1094 &  x1103 &  x1106 &  x1130;
assign c662 =  x73 &  x83 &  x89 &  x122 &  x268 &  x277 &  x284 &  x307 &  x347 &  x374 &  x386 &  x491 &  x503 &  x677 &  x769 &  x793 &  x871 &  x877 &  x931 &  x959 &  x988 &  x1049 &  x1130 & ~x324 & ~x480;
assign c664 =  x101 &  x128 &  x161 &  x182 &  x221 &  x284 &  x302 &  x386 &  x461 &  x470 &  x494 &  x542 &  x692 &  x707 &  x716 &  x722 &  x755 &  x779 &  x803 &  x836 &  x845 &  x848 &  x959 &  x1001 &  x1028 &  x1079 &  x1103 & ~x366 & ~x405 & ~x480 & ~x520 & ~x549 & ~x588 & ~x627 & ~x828;
assign c666 =  x8 &  x14 &  x17 &  x23 &  x41 &  x68 &  x77 &  x80 &  x83 &  x92 &  x95 &  x101 &  x107 &  x113 &  x146 &  x164 &  x176 &  x197 &  x202 &  x203 &  x209 &  x218 &  x221 &  x230 &  x242 &  x269 &  x278 &  x284 &  x293 &  x302 &  x308 &  x317 &  x350 &  x371 &  x392 &  x395 &  x404 &  x407 &  x419 &  x440 &  x455 &  x461 &  x464 &  x479 &  x482 &  x485 &  x491 &  x494 &  x503 &  x518 &  x536 &  x548 &  x551 &  x557 &  x563 &  x569 &  x578 &  x584 &  x587 &  x632 &  x635 &  x638 &  x647 &  x659 &  x668 &  x674 &  x680 &  x686 &  x692 &  x725 &  x728 &  x731 &  x734 &  x737 &  x740 &  x743 &  x770 &  x773 &  x785 &  x788 &  x800 &  x809 &  x818 &  x824 &  x830 &  x833 &  x839 &  x848 &  x866 &  x869 &  x881 &  x884 &  x899 &  x902 &  x905 &  x908 &  x926 &  x932 &  x934 &  x953 &  x956 &  x962 &  x968 &  x977 &  x983 &  x986 &  x998 &  x1022 &  x1028 &  x1031 &  x1043 &  x1049 &  x1055 &  x1064 &  x1085 &  x1088 &  x1091 &  x1109 &  x1124 &  x1130 & ~x60 & ~x78 & ~x99 & ~x126 & ~x165 & ~x196 & ~x210 & ~x249 & ~x255 & ~x288 & ~x294 & ~x327 & ~x444 & ~x483;
assign c668 =  x77 &  x83 &  x188 &  x256 &  x295 &  x379 &  x418 &  x496 &  x587 &  x800 &  x886 &  x992 &  x1007 & ~x474 & ~x480 & ~x513 & ~x552 & ~x597 & ~x1017;
assign c670 =  x10 &  x32 &  x49 &  x68 &  x77 &  x83 &  x88 &  x89 &  x95 &  x116 &  x127 &  x137 &  x164 &  x166 &  x167 &  x173 &  x176 &  x191 &  x194 &  x209 &  x221 &  x227 &  x239 &  x281 &  x284 &  x296 &  x302 &  x310 &  x326 &  x347 &  x350 &  x356 &  x374 &  x386 &  x388 &  x389 &  x395 &  x398 &  x401 &  x404 &  x407 &  x413 &  x419 &  x437 &  x452 &  x466 &  x470 &  x479 &  x485 &  x506 &  x509 &  x518 &  x524 &  x551 &  x557 &  x563 &  x566 &  x569 &  x587 &  x590 &  x593 &  x602 &  x614 &  x620 &  x623 &  x632 &  x644 &  x650 &  x659 &  x677 &  x680 &  x689 &  x707 &  x722 &  x728 &  x731 &  x743 &  x761 &  x764 &  x788 &  x800 &  x824 &  x827 &  x833 &  x839 &  x848 &  x860 &  x863 &  x866 &  x872 &  x884 &  x908 &  x920 &  x926 &  x944 &  x947 &  x968 &  x977 &  x980 &  x986 &  x995 &  x998 &  x1016 &  x1022 &  x1031 &  x1046 &  x1052 &  x1055 &  x1076 &  x1079 &  x1088 &  x1091 &  x1097 &  x1124 & ~x312 & ~x360 & ~x399 & ~x438 & ~x678 & ~x714 & ~x717;
assign c672 =  x14 &  x29 &  x65 &  x68 &  x83 &  x101 &  x110 &  x128 &  x191 &  x197 &  x203 &  x221 &  x227 &  x257 &  x284 &  x290 &  x292 &  x299 &  x302 &  x311 &  x341 &  x347 &  x374 &  x380 &  x392 &  x395 &  x398 &  x407 &  x419 &  x422 &  x425 &  x437 &  x473 &  x476 &  x482 &  x529 &  x536 &  x545 &  x568 &  x569 &  x578 &  x587 &  x590 &  x608 &  x619 &  x623 &  x644 &  x650 &  x671 &  x680 &  x692 &  x706 &  x719 &  x722 &  x728 &  x740 &  x743 &  x745 &  x758 &  x764 &  x788 &  x818 &  x836 &  x848 &  x860 &  x866 &  x881 &  x893 &  x902 &  x920 &  x950 &  x953 &  x979 &  x1016 &  x1022 &  x1031 &  x1043 &  x1067 &  x1088 &  x1097 &  x1127 &  x1130 & ~x393 & ~x399 & ~x438 & ~x717 & ~x756;
assign c674 =  x14 &  x23 &  x59 &  x77 &  x83 &  x101 &  x110 &  x116 &  x122 &  x137 &  x149 &  x161 &  x176 &  x194 &  x209 &  x242 &  x257 &  x287 &  x296 &  x353 &  x356 &  x401 &  x407 &  x419 &  x437 &  x455 &  x479 &  x503 &  x518 &  x536 &  x554 &  x557 &  x566 &  x587 &  x602 &  x604 &  x605 &  x608 &  x610 &  x611 &  x614 &  x643 &  x671 &  x677 &  x692 &  x701 &  x710 &  x722 &  x725 &  x728 &  x734 &  x743 &  x752 &  x764 &  x773 &  x785 &  x794 &  x809 &  x854 &  x884 &  x908 &  x920 &  x941 &  x947 &  x953 &  x965 &  x971 &  x983 &  x995 &  x998 &  x1001 &  x1022 &  x1040 &  x1046 &  x1049 &  x1073 &  x1079 &  x1097 &  x1103 & ~x12 & ~x246 & ~x285 & ~x303 & ~x342 & ~x363 & ~x364 & ~x366 & ~x402 & ~x441 & ~x480 & ~x663;
assign c676 =  x262 &  x301 &  x340 &  x410 &  x415 &  x427 &  x460 &  x493 &  x496 &  x532 &  x535 &  x602 &  x607 &  x646 &  x650 &  x685 &  x724 &  x800 &  x802 &  x812 &  x832 &  x863 &  x866 &  x886 &  x899 &  x1001 &  x1022 &  x1027 &  x1075 &  x1114;
assign c678 =  x22 &  x53 &  x56 &  x61 &  x83 &  x95 &  x98 &  x100 &  x101 &  x107 &  x134 &  x139 &  x151 &  x152 &  x155 &  x160 &  x167 &  x190 &  x191 &  x212 &  x215 &  x224 &  x229 &  x260 &  x268 &  x281 &  x293 &  x307 &  x308 &  x320 &  x344 &  x350 &  x359 &  x374 &  x392 &  x425 &  x436 &  x446 &  x455 &  x491 &  x515 &  x532 &  x535 &  x545 &  x569 &  x571 &  x610 &  x617 &  x649 &  x680 &  x688 &  x701 &  x716 &  x725 &  x730 &  x740 &  x743 &  x746 &  x752 &  x763 &  x769 &  x802 &  x808 &  x809 &  x815 &  x818 &  x841 &  x845 &  x848 &  x851 &  x880 &  x884 &  x886 &  x919 &  x935 &  x958 &  x974 &  x977 &  x986 &  x989 &  x997 &  x998 &  x1001 &  x1040 &  x1049 &  x1055 &  x1058 &  x1075 &  x1082 &  x1100 &  x1124;
assign c680 =  x5 &  x50 &  x59 &  x74 &  x116 &  x143 &  x146 &  x188 &  x284 &  x323 &  x341 &  x386 &  x395 &  x464 &  x479 &  x506 &  x521 &  x536 &  x569 &  x587 &  x593 &  x599 &  x622 &  x659 &  x661 &  x710 &  x728 &  x761 &  x791 &  x812 &  x824 &  x833 &  x836 &  x875 &  x884 &  x890 &  x941 &  x1010 &  x1055 &  x1070 & ~x0 & ~x3 & ~x222 & ~x249 & ~x288 & ~x327 & ~x483 & ~x549 & ~x588;
assign c682 =  x23 &  x26 &  x101 &  x110 &  x122 &  x143 &  x146 &  x170 &  x221 &  x230 &  x239 &  x278 &  x284 &  x299 &  x308 &  x311 &  x317 &  x350 &  x353 &  x362 &  x368 &  x380 &  x386 &  x389 &  x431 &  x434 &  x437 &  x451 &  x455 &  x479 &  x485 &  x497 &  x518 &  x529 &  x551 &  x563 &  x568 &  x569 &  x575 &  x605 &  x606 &  x623 &  x626 &  x644 &  x646 &  x650 &  x665 &  x677 &  x680 &  x685 &  x692 &  x728 &  x731 &  x734 &  x737 &  x743 &  x746 &  x779 &  x788 &  x800 &  x818 &  x824 &  x830 &  x836 &  x851 &  x857 &  x860 &  x866 &  x869 &  x877 &  x884 &  x889 &  x899 &  x920 &  x926 &  x932 &  x956 &  x959 &  x961 &  x968 &  x986 &  x994 &  x1016 &  x1027 &  x1028 &  x1033 &  x1064 &  x1066 &  x1067 &  x1072 &  x1085 &  x1097 &  x1109 &  x1111 &  x1117 &  x1124 & ~x135;
assign c684 =  x43 &  x82 &  x121 &  x122 &  x146 &  x160 &  x166 &  x221 &  x277 &  x392 &  x482 &  x661 &  x713 &  x743 &  x761 &  x830 &  x877 &  x881 &  x947 & ~x132 & ~x174 & ~x213 & ~x249 & ~x468;
assign c686 =  x14 &  x35 &  x56 &  x74 &  x80 &  x83 &  x92 &  x119 &  x128 &  x131 &  x155 &  x164 &  x176 &  x179 &  x185 &  x203 &  x209 &  x221 &  x224 &  x230 &  x239 &  x242 &  x257 &  x284 &  x290 &  x308 &  x341 &  x344 &  x356 &  x370 &  x383 &  x395 &  x398 &  x404 &  x413 &  x419 &  x427 &  x434 &  x437 &  x479 &  x485 &  x494 &  x500 &  x518 &  x524 &  x529 &  x568 &  x584 &  x593 &  x602 &  x620 &  x623 &  x641 &  x647 &  x667 &  x680 &  x686 &  x706 &  x707 &  x713 &  x734 &  x745 &  x758 &  x785 &  x800 &  x803 &  x823 &  x833 &  x842 &  x845 &  x862 &  x881 &  x890 &  x899 &  x901 &  x905 &  x908 &  x911 &  x923 &  x938 &  x944 &  x947 &  x953 &  x956 &  x959 &  x979 &  x1001 &  x1016 &  x1018 &  x1022 &  x1043 &  x1046 &  x1055 &  x1085 &  x1091 &  x1112 &  x1127 & ~x483 & ~x597 & ~x636;
assign c688 =  x23 &  x41 &  x62 &  x77 &  x80 &  x128 &  x146 &  x155 &  x161 &  x164 &  x176 &  x179 &  x191 &  x200 &  x218 &  x233 &  x236 &  x254 &  x263 &  x287 &  x299 &  x326 &  x335 &  x347 &  x356 &  x377 &  x380 &  x389 &  x392 &  x410 &  x467 &  x479 &  x485 &  x497 &  x500 &  x503 &  x512 &  x527 &  x533 &  x536 &  x548 &  x560 &  x563 &  x566 &  x584 &  x587 &  x605 &  x620 &  x623 &  x632 &  x635 &  x647 &  x650 &  x653 &  x659 &  x668 &  x671 &  x680 &  x689 &  x698 &  x701 &  x704 &  x719 &  x725 &  x731 &  x734 &  x737 &  x749 &  x761 &  x776 &  x779 &  x782 &  x788 &  x797 &  x800 &  x827 &  x839 &  x857 &  x866 &  x884 &  x887 &  x890 &  x893 &  x896 &  x908 &  x911 &  x923 &  x932 &  x935 &  x938 &  x941 &  x944 &  x953 &  x980 &  x986 &  x998 &  x1001 &  x1013 &  x1031 &  x1040 &  x1055 &  x1061 &  x1064 &  x1079 &  x1088 & ~x321 & ~x519 & ~x561 & ~x564 & ~x600 & ~x603 & ~x639 & ~x642 & ~x714 & ~x831 & ~x870 & ~x909 & ~x948 & ~x987 & ~x993 & ~x1026 & ~x1032 & ~x1065;
assign c690 =  x8 &  x11 &  x17 &  x29 &  x83 &  x95 &  x176 &  x284 &  x302 &  x332 &  x347 &  x350 &  x374 &  x386 &  x434 &  x455 &  x473 &  x491 &  x518 &  x530 &  x611 &  x668 &  x677 &  x770 &  x800 &  x833 &  x839 &  x845 &  x866 &  x875 &  x899 &  x926 &  x941 &  x968 &  x1001 &  x1022 &  x1031 &  x1097 &  x1127 & ~x132 & ~x150 & ~x171 & ~x210 & ~x288 & ~x666 & ~x717 & ~x795 & ~x834 & ~x867 & ~x873 & ~x906 & ~x945 & ~x984 & ~x1062 & ~x1080 & ~x1101 & ~x1119;
assign c692 =  x2 &  x23 &  x32 &  x53 &  x76 &  x77 &  x83 &  x89 &  x92 &  x101 &  x119 &  x128 &  x131 &  x140 &  x157 &  x158 &  x164 &  x173 &  x203 &  x230 &  x236 &  x242 &  x248 &  x260 &  x263 &  x266 &  x269 &  x275 &  x277 &  x278 &  x281 &  x296 &  x302 &  x326 &  x332 &  x344 &  x350 &  x374 &  x380 &  x392 &  x395 &  x398 &  x413 &  x485 &  x491 &  x494 &  x503 &  x515 &  x518 &  x532 &  x536 &  x548 &  x566 &  x569 &  x571 &  x578 &  x584 &  x587 &  x605 &  x610 &  x620 &  x649 &  x659 &  x671 &  x677 &  x680 &  x686 &  x688 &  x689 &  x695 &  x710 &  x743 &  x746 &  x749 &  x764 &  x776 &  x779 &  x785 &  x791 &  x800 &  x803 &  x851 &  x881 &  x887 &  x902 &  x905 &  x911 &  x914 &  x923 &  x926 &  x929 &  x932 &  x944 &  x947 &  x983 &  x986 &  x989 &  x992 &  x1001 &  x1016 &  x1022 &  x1025 &  x1028 &  x1031 &  x1043 &  x1085 &  x1097 &  x1100 &  x1106 &  x1124 &  x1127 & ~x423 & ~x462 & ~x468 & ~x501 & ~x510 & ~x546 & ~x549 & ~x588;
assign c694 =  x14 &  x77 &  x83 &  x89 &  x92 &  x101 &  x110 &  x152 &  x167 &  x203 &  x209 &  x239 &  x242 &  x269 &  x284 &  x302 &  x317 &  x326 &  x335 &  x350 &  x371 &  x374 &  x392 &  x395 &  x407 &  x431 &  x434 &  x482 &  x485 &  x491 &  x503 &  x518 &  x590 &  x635 &  x644 &  x653 &  x659 &  x680 &  x692 &  x698 &  x701 &  x707 &  x713 &  x722 &  x743 &  x746 &  x764 &  x770 &  x800 &  x824 &  x839 &  x848 &  x862 &  x866 &  x899 &  x901 &  x944 &  x947 &  x953 &  x959 &  x968 &  x980 &  x995 &  x1001 &  x1022 &  x1031 &  x1049 &  x1055 &  x1097 &  x1103 &  x1106 & ~x105 & ~x144 & ~x222 & ~x441 & ~x480 & ~x481 & ~x513 & ~x519 & ~x520 & ~x558 & ~x559 & ~x597 & ~x636;
assign c696 =  x8 &  x77 &  x95 &  x100 &  x110 &  x151 &  x178 &  x229 &  x295 &  x329 &  x347 &  x359 &  x395 &  x419 &  x428 &  x434 &  x451 &  x530 &  x568 &  x607 &  x619 &  x620 &  x707 &  x722 &  x734 &  x763 &  x770 &  x802 &  x848 &  x872 &  x880 &  x893 &  x919 &  x983 &  x1036 &  x1075 &  x1121 &  x1130 & ~x321 & ~x732 & ~x825;
assign c698 =  x197 &  x347 &  x356 &  x421 &  x460 &  x537 &  x575 &  x848 &  x854 &  x968 &  x986 &  x1018 &  x1069 &  x1129 & ~x549 & ~x753 & ~x792 & ~x831;
assign c6100 =  x2 &  x32 &  x86 &  x89 &  x92 &  x101 &  x110 &  x119 &  x137 &  x152 &  x164 &  x166 &  x170 &  x176 &  x182 &  x188 &  x194 &  x197 &  x205 &  x209 &  x221 &  x257 &  x269 &  x281 &  x284 &  x293 &  x305 &  x308 &  x326 &  x335 &  x362 &  x371 &  x374 &  x386 &  x388 &  x389 &  x395 &  x397 &  x404 &  x407 &  x415 &  x419 &  x427 &  x431 &  x452 &  x454 &  x466 &  x482 &  x491 &  x503 &  x515 &  x518 &  x521 &  x536 &  x548 &  x566 &  x569 &  x587 &  x590 &  x650 &  x659 &  x668 &  x674 &  x680 &  x698 &  x710 &  x722 &  x728 &  x749 &  x752 &  x764 &  x800 &  x806 &  x824 &  x839 &  x845 &  x848 &  x851 &  x860 &  x866 &  x899 &  x920 &  x947 &  x953 &  x956 &  x959 &  x989 &  x992 &  x998 &  x1016 &  x1022 &  x1034 &  x1040 &  x1055 &  x1079 &  x1088 &  x1097 &  x1106 & ~x391 & ~x399 & ~x429 & ~x430 & ~x438 & ~x468 & ~x477 & ~x678;
assign c6102 =  x35 &  x101 &  x110 &  x254 &  x404 &  x419 &  x436 &  x500 &  x536 &  x566 &  x620 &  x635 &  x644 &  x656 &  x680 &  x749 &  x800 &  x839 &  x848 &  x860 &  x1031 & ~x132 & ~x171 & ~x249 & ~x288 & ~x327 & ~x438 & ~x516 & ~x711 & ~x756 & ~x828 & ~x906 & ~x945 & ~x1023;
assign c6104 =  x77 &  x140 &  x176 &  x194 &  x203 &  x368 &  x377 &  x548 &  x650 &  x680 &  x746 &  x800 &  x929 &  x1028 &  x1055 &  x1109 & ~x396 & ~x435 & ~x438 & ~x627 & ~x666 & ~x708 & ~x825 & ~x903 & ~x942 & ~x981 & ~x982 & ~x1020 & ~x1026 & ~x1059 & ~x1065 & ~x1116;
assign c6106 =  x5 &  x32 &  x41 &  x53 &  x74 &  x77 &  x122 &  x221 &  x239 &  x257 &  x269 &  x344 &  x347 &  x407 &  x467 &  x482 &  x500 &  x536 &  x539 &  x569 &  x590 &  x605 &  x632 &  x635 &  x677 &  x707 &  x722 &  x746 &  x752 &  x779 &  x799 &  x824 &  x827 &  x848 &  x866 &  x899 &  x902 &  x908 &  x914 &  x947 &  x1001 &  x1022 &  x1034 &  x1055 & ~x210 & ~x249 & ~x324 & ~x363 & ~x364 & ~x396 & ~x402 & ~x435 & ~x441 & ~x474 & ~x480;
assign c6108 =  x14 &  x32 &  x35 &  x56 &  x77 &  x92 &  x167 &  x356 &  x386 &  x389 &  x413 &  x416 &  x506 &  x518 &  x563 &  x599 &  x731 &  x758 &  x818 &  x845 &  x862 &  x908 &  x920 &  x944 &  x986 &  x995 &  x1001 &  x1037 &  x1058 &  x1106 &  x1118 & ~x87 & ~x132 & ~x321 & ~x441 & ~x483 & ~x522 & ~x561 & ~x597 & ~x600 & ~x639 & ~x642;
assign c6110 =  x86 &  x101 &  x103 &  x116 &  x142 &  x205 &  x230 &  x278 &  x284 &  x308 &  x337 &  x353 &  x376 &  x377 &  x392 &  x425 &  x453 &  x454 &  x485 &  x493 &  x515 &  x532 &  x535 &  x536 &  x569 &  x574 &  x587 &  x668 &  x713 &  x749 &  x770 &  x785 &  x881 &  x889 &  x968 &  x1001 &  x1006 &  x1022 &  x1039;
assign c6112 =  x269 &  x677 &  x692 &  x764 &  x905 &  x934 &  x967 &  x980 & ~x132 & ~x211 & ~x249 & ~x250 & ~x285 & ~x289 & ~x328 & ~x828 & ~x906 & ~x945;
assign c6114 =  x32 &  x92 &  x164 &  x167 &  x221 &  x230 &  x242 &  x317 &  x347 &  x395 &  x398 &  x413 &  x503 &  x515 &  x539 &  x590 &  x605 &  x647 &  x764 &  x797 &  x830 &  x863 &  x866 &  x890 &  x899 &  x995 & ~x276 & ~x285 & ~x324 & ~x363 & ~x402 & ~x441 & ~x480 & ~x519 & ~x558 & ~x597 & ~x714 & ~x753 & ~x831 & ~x870 & ~x909 & ~x927 & ~x948 & ~x949 & ~x987 & ~x1026 & ~x1065;
assign c6116 =  x100 &  x184 &  x229 &  x296 &  x307 &  x340 &  x379 &  x388 &  x535 &  x620 &  x673 &  x752 &  x790 &  x844 &  x989 &  x1007 &  x1111 & ~x393 & ~x432;
assign c6118 =  x14 &  x41 &  x47 &  x77 &  x110 &  x119 &  x152 &  x176 &  x215 &  x221 &  x239 &  x257 &  x326 &  x368 &  x371 &  x374 &  x380 &  x392 &  x395 &  x425 &  x458 &  x479 &  x482 &  x485 &  x491 &  x518 &  x548 &  x557 &  x587 &  x590 &  x593 &  x599 &  x602 &  x611 &  x617 &  x623 &  x659 &  x701 &  x719 &  x746 &  x797 &  x800 &  x830 &  x833 &  x877 &  x884 &  x902 &  x926 &  x959 &  x968 &  x983 &  x986 &  x998 &  x1001 &  x1055 &  x1064 &  x1088 &  x1097 & ~x93 & ~x132 & ~x171 & ~x210 & ~x249 & ~x255 & ~x288 & ~x327 & ~x333 & ~x859 & ~x937 & ~x939 & ~x1017;
assign c6120 =  x4 &  x26 &  x32 &  x35 &  x43 &  x89 &  x110 &  x152 &  x164 &  x176 &  x197 &  x257 &  x269 &  x284 &  x308 &  x311 &  x326 &  x335 &  x359 &  x377 &  x383 &  x395 &  x398 &  x452 &  x491 &  x500 &  x536 &  x563 &  x569 &  x575 &  x587 &  x590 &  x605 &  x617 &  x623 &  x650 &  x680 &  x686 &  x698 &  x707 &  x713 &  x734 &  x737 &  x740 &  x761 &  x791 &  x797 &  x806 &  x830 &  x848 &  x875 &  x881 &  x884 &  x920 &  x947 &  x956 &  x995 &  x998 &  x1001 &  x1022 &  x1064 &  x1070 &  x1127 & ~x540 & ~x666 & ~x942 & ~x981 & ~x1020 & ~x1044 & ~x1080 & ~x1089 & ~x1119;
assign c6122 =  x2 &  x8 &  x29 &  x44 &  x65 &  x71 &  x77 &  x80 &  x89 &  x92 &  x110 &  x116 &  x128 &  x194 &  x197 &  x203 &  x209 &  x215 &  x221 &  x227 &  x230 &  x233 &  x242 &  x245 &  x260 &  x272 &  x278 &  x284 &  x290 &  x302 &  x308 &  x326 &  x335 &  x350 &  x371 &  x374 &  x386 &  x388 &  x392 &  x395 &  x398 &  x404 &  x407 &  x434 &  x455 &  x485 &  x500 &  x515 &  x518 &  x530 &  x533 &  x536 &  x551 &  x563 &  x566 &  x569 &  x575 &  x590 &  x602 &  x628 &  x632 &  x644 &  x647 &  x650 &  x653 &  x659 &  x667 &  x692 &  x695 &  x698 &  x701 &  x707 &  x719 &  x737 &  x743 &  x749 &  x785 &  x809 &  x815 &  x824 &  x833 &  x845 &  x860 &  x869 &  x887 &  x893 &  x902 &  x920 &  x929 &  x944 &  x953 &  x959 &  x980 &  x995 &  x1001 &  x1019 &  x1031 &  x1043 &  x1079 &  x1088 &  x1121 & ~x273 & ~x363 & ~x402 & ~x441 & ~x444 & ~x480 & ~x483 & ~x519 & ~x522 & ~x561 & ~x597 & ~x603 & ~x636;
assign c6124 =  x8 &  x14 &  x29 &  x32 &  x83 &  x110 &  x122 &  x125 &  x137 &  x149 &  x152 &  x164 &  x203 &  x221 &  x263 &  x266 &  x269 &  x272 &  x278 &  x302 &  x308 &  x316 &  x317 &  x323 &  x338 &  x344 &  x347 &  x355 &  x359 &  x374 &  x395 &  x404 &  x437 &  x446 &  x449 &  x455 &  x458 &  x467 &  x482 &  x494 &  x509 &  x518 &  x536 &  x548 &  x581 &  x590 &  x593 &  x602 &  x614 &  x620 &  x623 &  x632 &  x638 &  x647 &  x653 &  x659 &  x674 &  x686 &  x692 &  x719 &  x722 &  x725 &  x731 &  x734 &  x737 &  x740 &  x743 &  x770 &  x779 &  x785 &  x809 &  x827 &  x830 &  x832 &  x839 &  x845 &  x866 &  x871 &  x875 &  x878 &  x889 &  x893 &  x896 &  x899 &  x902 &  x904 &  x905 &  x908 &  x910 &  x917 &  x920 &  x922 &  x926 &  x932 &  x947 &  x949 &  x953 &  x959 &  x961 &  x962 &  x967 &  x968 &  x980 &  x983 &  x988 &  x992 &  x998 &  x1027 &  x1033 &  x1037 &  x1045 &  x1046 &  x1058 &  x1064 &  x1066 &  x1072 &  x1076 &  x1079 &  x1085 &  x1091 &  x1097 &  x1100 &  x1115 &  x1124 &  x1127 & ~x93 & ~x249 & ~x285 & ~x288 & ~x324 & ~x369 & ~x405;
assign c6126 =  x14 &  x23 &  x32 &  x35 &  x53 &  x83 &  x86 &  x110 &  x122 &  x128 &  x131 &  x137 &  x140 &  x152 &  x164 &  x167 &  x197 &  x209 &  x218 &  x239 &  x242 &  x272 &  x278 &  x296 &  x302 &  x308 &  x323 &  x326 &  x347 &  x350 &  x374 &  x395 &  x398 &  x410 &  x419 &  x425 &  x428 &  x431 &  x461 &  x464 &  x482 &  x503 &  x527 &  x548 &  x551 &  x563 &  x566 &  x587 &  x611 &  x647 &  x692 &  x707 &  x710 &  x716 &  x725 &  x728 &  x731 &  x734 &  x740 &  x743 &  x761 &  x770 &  x785 &  x788 &  x809 &  x818 &  x833 &  x839 &  x845 &  x848 &  x869 &  x881 &  x884 &  x899 &  x902 &  x905 &  x923 &  x935 &  x947 &  x956 &  x959 &  x962 &  x968 &  x989 &  x992 &  x995 &  x998 &  x1016 &  x1019 &  x1022 &  x1028 &  x1031 &  x1040 &  x1049 &  x1079 &  x1085 &  x1097 &  x1118 &  x1121 &  x1124 & ~x165 & ~x273 & ~x312 & ~x321 & ~x405 & ~x522 & ~x561 & ~x597 & ~x600 & ~x639 & ~x640 & ~x678 & ~x717 & ~x756 & ~x1119;
assign c6128 =  x5 &  x14 &  x23 &  x26 &  x32 &  x35 &  x47 &  x56 &  x71 &  x77 &  x83 &  x89 &  x92 &  x95 &  x101 &  x113 &  x116 &  x122 &  x128 &  x137 &  x149 &  x152 &  x155 &  x164 &  x188 &  x194 &  x197 &  x203 &  x209 &  x221 &  x230 &  x242 &  x269 &  x278 &  x302 &  x305 &  x317 &  x323 &  x329 &  x350 &  x371 &  x392 &  x397 &  x404 &  x434 &  x466 &  x473 &  x479 &  x482 &  x491 &  x497 &  x500 &  x527 &  x530 &  x533 &  x551 &  x575 &  x584 &  x587 &  x590 &  x602 &  x605 &  x638 &  x644 &  x647 &  x653 &  x686 &  x692 &  x698 &  x707 &  x713 &  x731 &  x734 &  x746 &  x764 &  x779 &  x784 &  x788 &  x797 &  x806 &  x823 &  x827 &  x830 &  x833 &  x836 &  x839 &  x845 &  x862 &  x866 &  x869 &  x881 &  x884 &  x899 &  x901 &  x902 &  x908 &  x926 &  x929 &  x935 &  x940 &  x947 &  x962 &  x968 &  x979 &  x989 &  x1001 &  x1004 &  x1016 &  x1028 &  x1031 &  x1034 &  x1037 &  x1057 &  x1064 &  x1085 &  x1097 &  x1127 & ~x321 & ~x399 & ~x405 & ~x429 & ~x438 & ~x477 & ~x516 & ~x555 & ~x594 & ~x633 & ~x792 & ~x951;
assign c6130 =  x14 &  x32 &  x53 &  x77 &  x83 &  x110 &  x128 &  x176 &  x239 &  x269 &  x284 &  x347 &  x374 &  x389 &  x395 &  x398 &  x419 &  x452 &  x455 &  x482 &  x485 &  x503 &  x518 &  x536 &  x602 &  x623 &  x650 &  x677 &  x692 &  x707 &  x722 &  x725 &  x743 &  x761 &  x779 &  x788 &  x812 &  x824 &  x830 &  x839 &  x848 &  x866 &  x887 &  x920 &  x947 &  x968 &  x992 &  x1022 &  x1043 &  x1049 &  x1055 &  x1097 &  x1103 & ~x462 & ~x501 & ~x540 & ~x541 & ~x580 & ~x619 & ~x633 & ~x657 & ~x789 & ~x906;
assign c6132 =  x20 &  x68 &  x74 &  x77 &  x86 &  x89 &  x149 &  x176 &  x239 &  x296 &  x302 &  x308 &  x323 &  x326 &  x368 &  x380 &  x419 &  x425 &  x466 &  x494 &  x524 &  x536 &  x563 &  x572 &  x575 &  x587 &  x602 &  x620 &  x623 &  x647 &  x650 &  x656 &  x671 &  x767 &  x800 &  x821 &  x851 &  x860 &  x884 &  x899 &  x920 &  x944 &  x962 &  x977 &  x1043 &  x1046 &  x1079 &  x1091 &  x1109 & ~x93 & ~x132 & ~x171 & ~x411 & ~x438 & ~x510 & ~x522 & ~x561 & ~x756 & ~x834 & ~x873 & ~x963 & ~x1119;
assign c6134 =  x8 &  x14 &  x32 &  x53 &  x65 &  x92 &  x95 &  x101 &  x103 &  x116 &  x142 &  x149 &  x194 &  x197 &  x200 &  x209 &  x218 &  x227 &  x230 &  x239 &  x242 &  x275 &  x284 &  x298 &  x323 &  x332 &  x337 &  x338 &  x341 &  x374 &  x376 &  x395 &  x398 &  x413 &  x415 &  x419 &  x425 &  x443 &  x452 &  x479 &  x500 &  x503 &  x518 &  x536 &  x545 &  x548 &  x563 &  x566 &  x569 &  x602 &  x608 &  x629 &  x632 &  x671 &  x692 &  x707 &  x713 &  x725 &  x728 &  x770 &  x779 &  x788 &  x800 &  x821 &  x824 &  x833 &  x839 &  x851 &  x866 &  x881 &  x884 &  x953 &  x1016 &  x1022 &  x1043 &  x1079 &  x1097 &  x1103 & ~x483 & ~x522 & ~x523 & ~x561 & ~x562 & ~x600 & ~x601 & ~x603 & ~x639 & ~x642;
assign c6136 =  x22 &  x28 &  x50 &  x89 &  x145 &  x152 &  x308 &  x361 &  x419 &  x421 &  x437 &  x439 &  x476 &  x535 &  x574 &  x673 &  x695 &  x730 &  x751 &  x769 &  x790 &  x824 &  x845 &  x869 &  x880 &  x886 &  x907 &  x946 &  x1097 & ~x471;
assign c6138 =  x5 &  x8 &  x11 &  x14 &  x23 &  x47 &  x56 &  x62 &  x86 &  x122 &  x125 &  x152 &  x164 &  x194 &  x197 &  x218 &  x221 &  x269 &  x287 &  x302 &  x311 &  x314 &  x317 &  x323 &  x326 &  x344 &  x347 &  x350 &  x371 &  x386 &  x395 &  x401 &  x419 &  x421 &  x422 &  x440 &  x443 &  x449 &  x461 &  x466 &  x479 &  x482 &  x491 &  x506 &  x527 &  x530 &  x533 &  x542 &  x545 &  x551 &  x557 &  x565 &  x572 &  x575 &  x578 &  x590 &  x605 &  x608 &  x611 &  x616 &  x622 &  x637 &  x638 &  x641 &  x643 &  x646 &  x668 &  x680 &  x707 &  x746 &  x758 &  x767 &  x779 &  x794 &  x802 &  x806 &  x821 &  x830 &  x848 &  x851 &  x869 &  x881 &  x884 &  x887 &  x902 &  x938 &  x959 &  x962 &  x968 &  x983 &  x986 &  x989 &  x995 &  x1004 &  x1016 &  x1019 &  x1043 &  x1055 &  x1079 &  x1115 &  x1118 & ~x471 & ~x510 & ~x549 & ~x588 & ~x627 & ~x628;
assign c6140 =  x2 &  x14 &  x32 &  x47 &  x56 &  x62 &  x77 &  x80 &  x83 &  x89 &  x122 &  x134 &  x137 &  x146 &  x170 &  x176 &  x194 &  x203 &  x209 &  x220 &  x239 &  x242 &  x266 &  x278 &  x284 &  x287 &  x290 &  x296 &  x299 &  x311 &  x326 &  x337 &  x343 &  x350 &  x353 &  x356 &  x365 &  x368 &  x376 &  x383 &  x388 &  x392 &  x395 &  x401 &  x407 &  x416 &  x419 &  x425 &  x431 &  x434 &  x455 &  x473 &  x476 &  x488 &  x494 &  x500 &  x503 &  x506 &  x512 &  x530 &  x533 &  x542 &  x545 &  x551 &  x560 &  x563 &  x572 &  x581 &  x584 &  x593 &  x599 &  x602 &  x605 &  x611 &  x614 &  x617 &  x623 &  x632 &  x647 &  x650 &  x677 &  x689 &  x692 &  x701 &  x713 &  x722 &  x734 &  x746 &  x770 &  x773 &  x779 &  x788 &  x791 &  x794 &  x809 &  x824 &  x842 &  x845 &  x854 &  x860 &  x866 &  x875 &  x881 &  x890 &  x901 &  x908 &  x914 &  x919 &  x926 &  x940 &  x958 &  x959 &  x968 &  x971 &  x980 &  x998 &  x1001 &  x1013 &  x1016 &  x1018 &  x1022 &  x1028 &  x1034 &  x1040 &  x1046 &  x1052 &  x1055 &  x1058 &  x1079 &  x1088 &  x1091 &  x1094 & ~x234 & ~x273 & ~x312 & ~x352 & ~x399 & ~x678;
assign c6142 =  x8 &  x11 &  x32 &  x38 &  x47 &  x74 &  x80 &  x83 &  x89 &  x92 &  x101 &  x119 &  x122 &  x143 &  x146 &  x149 &  x152 &  x209 &  x221 &  x227 &  x263 &  x284 &  x287 &  x308 &  x335 &  x374 &  x380 &  x392 &  x395 &  x404 &  x419 &  x434 &  x455 &  x461 &  x494 &  x503 &  x509 &  x515 &  x518 &  x524 &  x548 &  x563 &  x566 &  x608 &  x644 &  x647 &  x650 &  x659 &  x668 &  x692 &  x710 &  x722 &  x743 &  x746 &  x749 &  x785 &  x788 &  x800 &  x830 &  x845 &  x851 &  x856 &  x860 &  x899 &  x902 &  x923 &  x934 &  x944 &  x947 &  x953 &  x959 &  x968 &  x973 &  x980 &  x983 &  x995 &  x998 &  x1001 &  x1016 &  x1019 &  x1049 &  x1055 &  x1061 &  x1085 &  x1127 & ~x60 & ~x210 & ~x249 & ~x255 & ~x294 & ~x327 & ~x483 & ~x522 & ~x561 & ~x591 & ~x600 & ~x639 & ~x990;
assign c6144 =  x20 &  x89 &  x122 &  x131 &  x146 &  x149 &  x164 &  x170 &  x176 &  x194 &  x248 &  x329 &  x374 &  x398 &  x422 &  x425 &  x428 &  x515 &  x536 &  x542 &  x545 &  x563 &  x569 &  x590 &  x596 &  x602 &  x653 &  x719 &  x722 &  x764 &  x767 &  x770 &  x788 &  x839 &  x860 &  x863 &  x887 &  x902 &  x926 &  x947 &  x1052 &  x1103 & ~x3 & ~x93 & ~x132 & ~x171 & ~x210 & ~x222 & ~x249 & ~x285 & ~x327 & ~x402 & ~x480 & ~x483 & ~x522 & ~x561 & ~x702 & ~x897;
assign c6146 =  x35 &  x176 &  x197 &  x392 &  x449 &  x466 &  x515 &  x677 &  x710 &  x713 &  x731 &  x737 &  x758 &  x809 &  x851 &  x920 &  x940 &  x941 &  x986 &  x1091 & ~x430 & ~x522 & ~x792 & ~x795 & ~x796 & ~x831 & ~x834;
assign c6148 =  x291 &  x387 &  x622 &  x823 &  x929 & ~x312;
assign c6150 =  x14 &  x77 &  x101 &  x113 &  x140 &  x161 &  x191 &  x251 &  x275 &  x290 &  x356 &  x380 &  x383 &  x449 &  x479 &  x494 &  x506 &  x509 &  x557 &  x587 &  x635 &  x680 &  x686 &  x689 &  x716 &  x722 &  x746 &  x749 &  x764 &  x839 &  x866 &  x959 &  x979 &  x986 &  x998 &  x1004 &  x1064 & ~x165 & ~x195 & ~x210 & ~x249 & ~x288 & ~x327 & ~x405 & ~x444 & ~x480 & ~x483 & ~x522 & ~x561 & ~x562 & ~x600 & ~x601 & ~x678 & ~x717;
assign c6152 =  x23 &  x122 &  x131 &  x167 &  x197 &  x202 &  x257 &  x269 &  x353 &  x386 &  x388 &  x395 &  x407 &  x416 &  x454 &  x497 &  x512 &  x551 &  x557 &  x623 &  x722 &  x764 &  x845 &  x959 &  x1034 &  x1079 &  x1088 & ~x235 & ~x274 & ~x522 & ~x561 & ~x600 & ~x756 & ~x795 & ~x798;
assign c6154 =  x4 &  x26 &  x43 &  x62 &  x82 &  x83 &  x89 &  x100 &  x104 &  x110 &  x112 &  x128 &  x151 &  x173 &  x182 &  x194 &  x203 &  x209 &  x218 &  x266 &  x268 &  x284 &  x293 &  x314 &  x338 &  x353 &  x356 &  x359 &  x380 &  x392 &  x443 &  x455 &  x461 &  x464 &  x479 &  x482 &  x485 &  x491 &  x529 &  x530 &  x536 &  x563 &  x568 &  x584 &  x607 &  x611 &  x646 &  x653 &  x659 &  x662 &  x677 &  x685 &  x722 &  x724 &  x728 &  x763 &  x791 &  x802 &  x809 &  x836 &  x841 &  x893 &  x914 &  x929 &  x1043 &  x1055 &  x1075 &  x1079 &  x1103 &  x1127 & ~x360 & ~x399 & ~x438 & ~x477;
assign c6156 =  x11 &  x53 &  x68 &  x80 &  x83 &  x86 &  x119 &  x143 &  x152 &  x203 &  x269 &  x353 &  x380 &  x388 &  x395 &  x407 &  x427 &  x431 &  x437 &  x449 &  x466 &  x479 &  x491 &  x500 &  x506 &  x518 &  x527 &  x554 &  x575 &  x596 &  x620 &  x635 &  x650 &  x659 &  x662 &  x683 &  x686 &  x722 &  x725 &  x737 &  x746 &  x761 &  x806 &  x827 &  x851 &  x866 &  x908 &  x950 &  x953 &  x962 &  x980 &  x989 &  x1007 &  x1034 &  x1061 &  x1073 &  x1076 &  x1115 & ~x391 & ~x399 & ~x438 & ~x522 & ~x561 & ~x600 & ~x753 & ~x756 & ~x831;
assign c6158 =  x20 &  x41 &  x47 &  x53 &  x89 &  x92 &  x137 &  x140 &  x149 &  x152 &  x158 &  x164 &  x167 &  x188 &  x197 &  x203 &  x245 &  x272 &  x281 &  x284 &  x308 &  x371 &  x395 &  x428 &  x437 &  x476 &  x497 &  x551 &  x554 &  x563 &  x566 &  x572 &  x632 &  x656 &  x680 &  x713 &  x764 &  x767 &  x776 &  x779 &  x799 &  x824 &  x839 &  x848 &  x851 &  x860 &  x887 &  x917 &  x926 &  x973 &  x977 &  x998 &  x1016 &  x1027 &  x1043 &  x1064 & ~x9 & ~x48 & ~x171 & ~x210 & ~x402 & ~x702 & ~x750 & ~x789 & ~x828 & ~x897 & ~x906 & ~x945 & ~x1023;
assign c6160 =  x2 &  x11 &  x14 &  x32 &  x35 &  x53 &  x77 &  x83 &  x89 &  x92 &  x101 &  x113 &  x119 &  x122 &  x128 &  x134 &  x149 &  x152 &  x158 &  x161 &  x170 &  x173 &  x194 &  x197 &  x203 &  x209 &  x218 &  x221 &  x227 &  x230 &  x236 &  x239 &  x242 &  x263 &  x272 &  x281 &  x284 &  x287 &  x302 &  x308 &  x311 &  x323 &  x326 &  x338 &  x347 &  x359 &  x371 &  x374 &  x377 &  x380 &  x383 &  x386 &  x392 &  x395 &  x398 &  x407 &  x428 &  x431 &  x437 &  x449 &  x452 &  x473 &  x476 &  x479 &  x482 &  x488 &  x491 &  x497 &  x500 &  x503 &  x509 &  x515 &  x536 &  x548 &  x551 &  x563 &  x566 &  x569 &  x572 &  x578 &  x581 &  x584 &  x587 &  x590 &  x602 &  x620 &  x635 &  x638 &  x647 &  x650 &  x653 &  x677 &  x680 &  x692 &  x698 &  x707 &  x713 &  x719 &  x722 &  x725 &  x728 &  x731 &  x743 &  x746 &  x764 &  x770 &  x779 &  x785 &  x788 &  x791 &  x815 &  x824 &  x827 &  x830 &  x839 &  x848 &  x851 &  x854 &  x860 &  x866 &  x884 &  x887 &  x890 &  x896 &  x902 &  x905 &  x908 &  x911 &  x920 &  x929 &  x935 &  x944 &  x947 &  x959 &  x962 &  x968 &  x980 &  x986 &  x992 &  x995 &  x1001 &  x1006 &  x1016 &  x1019 &  x1022 &  x1028 &  x1043 &  x1049 &  x1055 &  x1061 &  x1064 &  x1079 &  x1094 &  x1097 &  x1106 &  x1121 & ~x48 & ~x87 & ~x213 & ~x249 & ~x288 & ~x327 & ~x366 & ~x405 & ~x408 & ~x444 & ~x459 & ~x483 & ~x498 & ~x522 & ~x663 & ~x702 & ~x741;
assign c6162 =  x14 &  x35 &  x53 &  x71 &  x77 &  x80 &  x89 &  x92 &  x110 &  x122 &  x128 &  x131 &  x134 &  x140 &  x143 &  x152 &  x155 &  x164 &  x176 &  x185 &  x194 &  x197 &  x206 &  x224 &  x242 &  x254 &  x260 &  x269 &  x272 &  x275 &  x278 &  x302 &  x326 &  x349 &  x350 &  x353 &  x374 &  x383 &  x388 &  x395 &  x413 &  x419 &  x427 &  x428 &  x446 &  x452 &  x464 &  x466 &  x467 &  x482 &  x485 &  x491 &  x494 &  x497 &  x505 &  x512 &  x518 &  x536 &  x539 &  x551 &  x563 &  x566 &  x569 &  x575 &  x587 &  x596 &  x602 &  x614 &  x623 &  x644 &  x650 &  x659 &  x665 &  x668 &  x674 &  x677 &  x680 &  x683 &  x692 &  x707 &  x710 &  x722 &  x725 &  x743 &  x746 &  x749 &  x752 &  x755 &  x764 &  x770 &  x782 &  x784 &  x788 &  x800 &  x823 &  x824 &  x827 &  x836 &  x839 &  x845 &  x851 &  x860 &  x863 &  x866 &  x869 &  x884 &  x899 &  x902 &  x920 &  x923 &  x929 &  x940 &  x944 &  x953 &  x959 &  x968 &  x979 &  x986 &  x995 &  x998 &  x1001 &  x1004 &  x1016 &  x1019 &  x1022 &  x1031 &  x1043 &  x1055 &  x1067 &  x1082 &  x1088 &  x1094 &  x1097 &  x1106 &  x1127 & ~x255 & ~x345 & ~x483 & ~x516 & ~x522 & ~x555 & ~x1101;
assign c6164 =  x8 &  x32 &  x77 &  x116 &  x137 &  x146 &  x152 &  x167 &  x194 &  x218 &  x230 &  x239 &  x254 &  x329 &  x355 &  x395 &  x398 &  x407 &  x431 &  x443 &  x500 &  x518 &  x587 &  x590 &  x622 &  x661 &  x734 &  x839 &  x854 &  x857 &  x881 &  x920 &  x932 &  x944 &  x989 &  x992 &  x995 &  x1007 &  x1013 &  x1028 &  x1031 &  x1034 &  x1043 &  x1046 &  x1052 &  x1088 & ~x54 & ~x93 & ~x132 & ~x171 & ~x210 & ~x438 & ~x516 & ~x546 & ~x547 & ~x555 & ~x585;
assign c6166 =  x83 &  x122 &  x176 &  x197 &  x335 &  x353 &  x452 &  x482 &  x518 &  x569 &  x754 &  x793 &  x809 &  x818 &  x832 &  x881 &  x889 &  x904 &  x905 &  x908 &  x910 &  x934 &  x943 &  x988 &  x1001 &  x1022 &  x1033 &  x1051 &  x1085 &  x1111 & ~x249 & ~x546 & ~x549 & ~x627 & ~x861;
assign c6168 =  x44 &  x119 &  x122 &  x128 &  x197 &  x269 &  x308 &  x343 &  x376 &  x395 &  x419 &  x421 &  x427 &  x431 &  x440 &  x452 &  x454 &  x455 &  x461 &  x464 &  x466 &  x479 &  x482 &  x493 &  x499 &  x500 &  x647 &  x650 &  x710 &  x764 &  x842 &  x848 &  x851 &  x869 &  x899 &  x902 &  x908 &  x923 &  x932 &  x950 &  x959 &  x968 &  x992 &  x1001 &  x1037 &  x1046 &  x1052 &  x1055 &  x1057 &  x1067 &  x1085 &  x1106 & ~x591 & ~x720 & ~x756;
assign c6170 =  x14 &  x35 &  x101 &  x110 &  x125 &  x128 &  x152 &  x176 &  x194 &  x215 &  x263 &  x287 &  x308 &  x317 &  x388 &  x392 &  x395 &  x466 &  x536 &  x569 &  x710 &  x737 &  x746 &  x779 &  x848 &  x860 &  x884 &  x953 &  x979 &  x1019 &  x1067 &  x1100 & ~x312 & ~x561 & ~x600 & ~x639 & ~x756 & ~x873 & ~x981;
assign c6172 =  x47 &  x83 &  x110 &  x164 &  x203 &  x239 &  x242 &  x302 &  x307 &  x326 &  x350 &  x374 &  x380 &  x401 &  x419 &  x425 &  x536 &  x553 &  x569 &  x587 &  x688 &  x707 &  x721 &  x754 &  x760 &  x764 &  x770 &  x779 &  x785 &  x799 &  x800 &  x830 &  x832 &  x839 &  x856 &  x860 &  x871 &  x877 &  x884 &  x893 &  x904 &  x934 &  x943 &  x944 &  x947 &  x955 &  x973 &  x989 &  x1016 &  x1061 &  x1127 & ~x441 & ~x480 & ~x519;
assign c6174 =  x11 &  x14 &  x23 &  x29 &  x35 &  x47 &  x53 &  x71 &  x77 &  x80 &  x83 &  x89 &  x92 &  x98 &  x101 &  x110 &  x113 &  x116 &  x122 &  x134 &  x140 &  x146 &  x149 &  x167 &  x173 &  x176 &  x185 &  x203 &  x209 &  x215 &  x218 &  x221 &  x224 &  x245 &  x266 &  x269 &  x281 &  x284 &  x299 &  x302 &  x308 &  x317 &  x326 &  x335 &  x338 &  x350 &  x395 &  x407 &  x416 &  x419 &  x425 &  x434 &  x437 &  x443 &  x446 &  x449 &  x455 &  x470 &  x482 &  x488 &  x491 &  x497 &  x500 &  x512 &  x518 &  x533 &  x539 &  x542 &  x545 &  x557 &  x569 &  x572 &  x578 &  x587 &  x593 &  x599 &  x605 &  x626 &  x629 &  x638 &  x641 &  x650 &  x659 &  x662 &  x683 &  x688 &  x707 &  x710 &  x725 &  x728 &  x743 &  x746 &  x758 &  x761 &  x764 &  x767 &  x779 &  x785 &  x788 &  x800 &  x806 &  x821 &  x824 &  x827 &  x830 &  x836 &  x842 &  x845 &  x851 &  x866 &  x875 &  x878 &  x881 &  x902 &  x908 &  x926 &  x938 &  x944 &  x950 &  x953 &  x959 &  x962 &  x965 &  x968 &  x992 &  x1001 &  x1010 &  x1016 &  x1019 &  x1022 &  x1028 &  x1037 &  x1049 &  x1058 &  x1082 &  x1085 &  x1091 &  x1097 &  x1100 &  x1103 & ~x78 & ~x126 & ~x165 & ~x210 & ~x249 & ~x288 & ~x327 & ~x366 & ~x405 & ~x420 & ~x444 & ~x459 & ~x483 & ~x522 & ~x561 & ~x672;
assign c6176 =  x29 &  x32 &  x65 &  x71 &  x89 &  x101 &  x112 &  x151 &  x161 &  x167 &  x203 &  x217 &  x229 &  x256 &  x268 &  x278 &  x307 &  x308 &  x373 &  x374 &  x380 &  x410 &  x412 &  x460 &  x461 &  x473 &  x500 &  x529 &  x584 &  x632 &  x634 &  x646 &  x647 &  x659 &  x685 &  x695 &  x724 &  x749 &  x790 &  x800 &  x806 &  x824 &  x829 &  x839 &  x880 &  x884 &  x887 &  x892 &  x902 &  x929 &  x958 &  x959 &  x986 &  x992 &  x997 &  x1036 &  x1055 &  x1097 &  x1102 &  x1108 &  x1118 &  x1124;
assign c6178 =  x77 &  x80 &  x122 &  x125 &  x176 &  x227 &  x230 &  x242 &  x308 &  x314 &  x377 &  x416 &  x452 &  x479 &  x503 &  x509 &  x518 &  x536 &  x575 &  x581 &  x587 &  x629 &  x635 &  x647 &  x650 &  x653 &  x701 &  x734 &  x743 &  x764 &  x821 &  x854 &  x872 &  x893 &  x908 &  x920 &  x929 &  x959 &  x986 &  x1082 &  x1100 & ~x402 & ~x441 & ~x480 & ~x483 & ~x520 & ~x552 & ~x559 & ~x561 & ~x597 & ~x598 & ~x783 & ~x819;
assign c6180 =  x176 &  x203 &  x221 &  x259 &  x398 &  x431 &  x500 &  x569 &  x602 &  x716 &  x776 &  x779 &  x824 &  x899 &  x995 &  x1127 & ~x222 & ~x261 & ~x306 & ~x345 & ~x462 & ~x501 & ~x696 & ~x720 & ~x735 & ~x736;
assign c6182 =  x1 &  x2 &  x32 &  x184 &  x266 &  x284 &  x308 &  x389 &  x692 &  x760 &  x764 &  x799 &  x806 &  x815 &  x863 &  x914 &  x940 &  x956 &  x965 &  x976 &  x986 &  x1052 & ~x441 & ~x480 & ~x825 & ~x1005;
assign c6184 =  x176 &  x269 &  x284 &  x338 &  x401 &  x413 &  x479 &  x491 &  x593 &  x611 &  x704 &  x719 &  x721 &  x785 &  x839 &  x863 &  x947 &  x992 &  x1028 &  x1031 & ~x9 & ~x162 & ~x246 & ~x285 & ~x324 & ~x438 & ~x516 & ~x555 & ~x633 & ~x666 & ~x861;
assign c6186 =  x308 &  x571 &  x610 &  x683 &  x823 & ~x627 & ~x714 & ~x792 & ~x831 & ~x870 & ~x927;
assign c6188 =  x2 &  x14 &  x53 &  x101 &  x110 &  x122 &  x142 &  x203 &  x239 &  x311 &  x337 &  x350 &  x356 &  x380 &  x386 &  x395 &  x407 &  x416 &  x491 &  x563 &  x587 &  x590 &  x610 &  x620 &  x647 &  x686 &  x698 &  x707 &  x743 &  x749 &  x761 &  x785 &  x800 &  x830 &  x848 &  x899 &  x947 &  x995 &  x1037 &  x1038 &  x1043 &  x1079 &  x1085 &  x1097 &  x1117 & ~x162 & ~x552;
assign c6190 =  x11 &  x23 &  x32 &  x47 &  x83 &  x89 &  x128 &  x149 &  x167 &  x179 &  x185 &  x194 &  x215 &  x224 &  x227 &  x242 &  x257 &  x260 &  x269 &  x278 &  x284 &  x287 &  x308 &  x314 &  x343 &  x371 &  x374 &  x383 &  x389 &  x395 &  x407 &  x413 &  x428 &  x431 &  x452 &  x466 &  x479 &  x488 &  x491 &  x494 &  x506 &  x524 &  x557 &  x569 &  x593 &  x611 &  x623 &  x638 &  x644 &  x650 &  x659 &  x686 &  x722 &  x728 &  x731 &  x743 &  x770 &  x794 &  x797 &  x809 &  x818 &  x839 &  x848 &  x854 &  x857 &  x860 &  x905 &  x908 &  x932 &  x941 &  x944 &  x947 &  x962 &  x974 &  x1001 &  x1037 &  x1061 &  x1064 &  x1079 &  x1082 &  x1115 & ~x39 & ~x60 & ~x216 & ~x234 & ~x255 & ~x274 & ~x294 & ~x312 & ~x313 & ~x321 & ~x360 & ~x444 & ~x483 & ~x756 & ~x969;
assign c6192 =  x23 &  x26 &  x56 &  x86 &  x101 &  x125 &  x131 &  x146 &  x152 &  x167 &  x179 &  x194 &  x197 &  x209 &  x221 &  x227 &  x236 &  x242 &  x278 &  x284 &  x299 &  x371 &  x374 &  x395 &  x404 &  x491 &  x503 &  x515 &  x557 &  x563 &  x566 &  x575 &  x587 &  x590 &  x602 &  x629 &  x635 &  x650 &  x659 &  x668 &  x677 &  x692 &  x698 &  x707 &  x710 &  x716 &  x731 &  x746 &  x755 &  x764 &  x767 &  x788 &  x800 &  x833 &  x848 &  x851 &  x860 &  x908 &  x947 &  x989 &  x1022 &  x1049 &  x1058 &  x1061 &  x1064 &  x1097 & ~x195 & ~x321 & ~x360 & ~x399 & ~x444 & ~x483 & ~x522 & ~x714 & ~x756 & ~x831 & ~x834 & ~x909 & ~x948 & ~x987 & ~x1026;
assign c6194 =  x14 &  x23 &  x35 &  x44 &  x53 &  x56 &  x77 &  x83 &  x92 &  x101 &  x116 &  x128 &  x140 &  x146 &  x176 &  x182 &  x185 &  x188 &  x197 &  x200 &  x242 &  x251 &  x272 &  x277 &  x290 &  x293 &  x316 &  x329 &  x335 &  x338 &  x350 &  x355 &  x365 &  x380 &  x386 &  x395 &  x407 &  x422 &  x437 &  x458 &  x461 &  x509 &  x542 &  x557 &  x566 &  x575 &  x602 &  x605 &  x617 &  x641 &  x725 &  x731 &  x788 &  x793 &  x800 &  x809 &  x821 &  x869 &  x871 &  x872 &  x905 &  x914 &  x920 &  x929 &  x941 &  x944 &  x953 &  x962 &  x1001 &  x1010 &  x1019 &  x1040 &  x1046 &  x1064 &  x1079 &  x1100 &  x1124 &  x1127 & ~x246 & ~x285 & ~x288 & ~x325 & ~x363 & ~x364 & ~x585 & ~x588 & ~x666 & ~x822;
assign c6196 =  x49 &  x71 &  x73 &  x74 &  x116 &  x260 &  x268 &  x308 &  x320 &  x380 &  x397 &  x421 &  x460 &  x491 &  x493 &  x499 &  x532 &  x536 &  x581 &  x605 &  x730 &  x743 &  x751 &  x769 &  x782 &  x803 &  x827 &  x829 &  x860 &  x880 &  x886 &  x902 &  x947 &  x968 &  x1049 &  x1055 &  x1085 &  x1112 & ~x432;
assign c6198 =  x14 &  x53 &  x71 &  x76 &  x77 &  x101 &  x154 &  x161 &  x167 &  x239 &  x284 &  x296 &  x314 &  x395 &  x479 &  x485 &  x530 &  x536 &  x569 &  x602 &  x626 &  x635 &  x674 &  x677 &  x695 &  x794 &  x806 &  x815 &  x833 &  x911 &  x935 &  x947 &  x968 &  x1004 &  x1019 &  x1022 & ~x183 & ~x210 & ~x222 & ~x249 & ~x288 & ~x327 & ~x363 & ~x364 & ~x367 & ~x402;
assign c6200 =  x32 &  x67 &  x77 &  x79 &  x92 &  x128 &  x152 &  x158 &  x205 &  x206 &  x251 &  x260 &  x262 &  x278 &  x284 &  x287 &  x317 &  x346 &  x400 &  x439 &  x455 &  x557 &  x620 &  x650 &  x659 &  x674 &  x677 &  x686 &  x707 &  x716 &  x719 &  x728 &  x730 &  x761 &  x769 &  x788 &  x791 &  x814 &  x827 &  x853 &  x863 &  x899 &  x941 &  x944 &  x947 &  x962 &  x986 &  x998 &  x1001 &  x1022 &  x1040 &  x1067 & ~x207 & ~x246 & ~x408 & ~x666 & ~x1122;
assign c6202 =  x14 &  x20 &  x29 &  x38 &  x53 &  x65 &  x77 &  x89 &  x92 &  x110 &  x116 &  x122 &  x128 &  x143 &  x149 &  x152 &  x164 &  x176 &  x182 &  x188 &  x194 &  x197 &  x209 &  x215 &  x218 &  x221 &  x242 &  x244 &  x266 &  x278 &  x284 &  x293 &  x302 &  x335 &  x344 &  x365 &  x368 &  x371 &  x373 &  x392 &  x395 &  x398 &  x407 &  x412 &  x416 &  x431 &  x439 &  x451 &  x460 &  x470 &  x473 &  x479 &  x489 &  x490 &  x491 &  x500 &  x506 &  x518 &  x521 &  x529 &  x536 &  x542 &  x548 &  x551 &  x557 &  x566 &  x568 &  x569 &  x584 &  x587 &  x590 &  x602 &  x605 &  x608 &  x617 &  x620 &  x623 &  x644 &  x649 &  x650 &  x677 &  x680 &  x683 &  x688 &  x692 &  x707 &  x710 &  x722 &  x743 &  x761 &  x767 &  x773 &  x788 &  x800 &  x824 &  x839 &  x842 &  x845 &  x866 &  x872 &  x878 &  x881 &  x884 &  x899 &  x905 &  x908 &  x920 &  x935 &  x941 &  x944 &  x959 &  x968 &  x980 &  x989 &  x992 &  x1001 &  x1016 &  x1022 &  x1028 &  x1043 &  x1049 &  x1055 &  x1064 &  x1073 &  x1079 &  x1082 &  x1085 &  x1088 &  x1103 &  x1106 &  x1118 &  x1127 & ~x972 & ~x1011;
assign c6204 =  x49 &  x67 &  x73 &  x88 &  x100 &  x112 &  x145 &  x166 &  x295 &  x301 &  x385 &  x395 &  x397 &  x436 &  x463 &  x524 &  x769 &  x802 &  x907 &  x919 &  x958 &  x983 &  x1024 &  x1075 &  x1109;
assign c6206 =  x14 &  x65 &  x146 &  x188 &  x194 &  x233 &  x251 &  x388 &  x413 &  x473 &  x491 &  x512 &  x560 &  x656 &  x719 &  x746 &  x749 &  x758 &  x794 &  x797 &  x800 &  x851 &  x878 &  x899 &  x938 &  x953 &  x998 &  x1106 & ~x84 & ~x240 & ~x435 & ~x474 & ~x483 & ~x513 & ~x552 & ~x561 & ~x669 & ~x825 & ~x903 & ~x942 & ~x981;
assign c6208 =  x29 &  x35 &  x47 &  x83 &  x89 &  x98 &  x116 &  x122 &  x125 &  x142 &  x155 &  x176 &  x197 &  x203 &  x206 &  x221 &  x269 &  x278 &  x284 &  x290 &  x293 &  x305 &  x326 &  x341 &  x344 &  x365 &  x374 &  x392 &  x395 &  x398 &  x401 &  x455 &  x479 &  x482 &  x491 &  x509 &  x512 &  x521 &  x542 &  x575 &  x584 &  x599 &  x629 &  x632 &  x638 &  x659 &  x661 &  x677 &  x680 &  x704 &  x707 &  x722 &  x734 &  x737 &  x740 &  x745 &  x761 &  x782 &  x784 &  x823 &  x845 &  x848 &  x862 &  x899 &  x901 &  x920 &  x940 &  x953 &  x968 &  x974 &  x979 &  x992 &  x1001 &  x1019 &  x1022 &  x1049 &  x1057 &  x1079 &  x1106 &  x1115 & ~x324 & ~x438 & ~x516 & ~x555 & ~x714 & ~x753 & ~x792;
assign c6210 =  x23 &  x50 &  x77 &  x83 &  x92 &  x227 &  x230 &  x257 &  x269 &  x281 &  x326 &  x329 &  x374 &  x380 &  x383 &  x395 &  x443 &  x452 &  x479 &  x482 &  x515 &  x518 &  x521 &  x530 &  x545 &  x551 &  x566 &  x632 &  x644 &  x668 &  x740 &  x743 &  x746 &  x764 &  x788 &  x812 &  x827 &  x857 &  x860 &  x866 &  x881 &  x899 &  x902 &  x908 &  x941 &  x947 &  x983 &  x992 &  x998 &  x1001 &  x1004 &  x1016 &  x1043 &  x1046 &  x1097 & ~x663 & ~x690 & ~x702 & ~x703 & ~x730 & ~x735 & ~x774;
assign c6212 =  x14 &  x29 &  x38 &  x41 &  x53 &  x56 &  x77 &  x80 &  x83 &  x89 &  x98 &  x101 &  x110 &  x128 &  x131 &  x146 &  x149 &  x152 &  x158 &  x164 &  x176 &  x179 &  x194 &  x197 &  x203 &  x215 &  x218 &  x227 &  x242 &  x266 &  x272 &  x296 &  x308 &  x326 &  x332 &  x356 &  x380 &  x383 &  x392 &  x395 &  x398 &  x407 &  x410 &  x419 &  x431 &  x455 &  x473 &  x479 &  x482 &  x491 &  x500 &  x503 &  x506 &  x515 &  x542 &  x545 &  x548 &  x566 &  x569 &  x578 &  x587 &  x590 &  x602 &  x610 &  x626 &  x635 &  x638 &  x644 &  x650 &  x656 &  x671 &  x688 &  x692 &  x698 &  x704 &  x707 &  x712 &  x713 &  x722 &  x728 &  x731 &  x746 &  x751 &  x758 &  x770 &  x773 &  x779 &  x788 &  x790 &  x800 &  x806 &  x824 &  x829 &  x833 &  x839 &  x851 &  x860 &  x866 &  x872 &  x881 &  x893 &  x902 &  x920 &  x923 &  x947 &  x953 &  x959 &  x961 &  x968 &  x977 &  x986 &  x989 &  x1000 &  x1001 &  x1010 &  x1019 &  x1022 &  x1028 &  x1031 &  x1055 &  x1064 &  x1067 &  x1079 &  x1091 &  x1097 &  x1103 &  x1106 &  x1109 &  x1118 & ~x285 & ~x324 & ~x363 & ~x402 & ~x441 & ~x480 & ~x519 & ~x663 & ~x705;
assign c6214 =  x2 &  x11 &  x14 &  x32 &  x38 &  x62 &  x74 &  x77 &  x80 &  x89 &  x110 &  x122 &  x128 &  x131 &  x146 &  x164 &  x167 &  x170 &  x176 &  x182 &  x194 &  x203 &  x209 &  x239 &  x269 &  x272 &  x284 &  x298 &  x308 &  x311 &  x329 &  x335 &  x337 &  x356 &  x361 &  x392 &  x395 &  x398 &  x407 &  x415 &  x419 &  x431 &  x437 &  x440 &  x446 &  x494 &  x503 &  x506 &  x512 &  x527 &  x536 &  x551 &  x563 &  x566 &  x569 &  x575 &  x587 &  x590 &  x605 &  x607 &  x608 &  x623 &  x632 &  x659 &  x662 &  x677 &  x680 &  x692 &  x713 &  x746 &  x749 &  x758 &  x761 &  x764 &  x770 &  x773 &  x779 &  x785 &  x794 &  x824 &  x827 &  x830 &  x839 &  x842 &  x851 &  x860 &  x869 &  x884 &  x887 &  x895 &  x896 &  x899 &  x902 &  x920 &  x934 &  x947 &  x959 &  x973 &  x977 &  x992 &  x1004 &  x1012 &  x1016 &  x1022 &  x1043 &  x1049 &  x1051 &  x1052 &  x1055 &  x1073 &  x1090 &  x1097 &  x1103 &  x1106 &  x1109 &  x1127 & ~x444 & ~x483 & ~x522 & ~x561;
assign c6216 =  x2 &  x13 &  x14 &  x20 &  x23 &  x26 &  x44 &  x74 &  x77 &  x80 &  x101 &  x103 &  x116 &  x122 &  x140 &  x142 &  x143 &  x164 &  x167 &  x173 &  x176 &  x181 &  x188 &  x197 &  x203 &  x221 &  x230 &  x242 &  x251 &  x257 &  x265 &  x278 &  x281 &  x284 &  x290 &  x298 &  x304 &  x308 &  x311 &  x320 &  x323 &  x326 &  x329 &  x332 &  x337 &  x341 &  x343 &  x344 &  x350 &  x359 &  x362 &  x368 &  x376 &  x386 &  x388 &  x392 &  x395 &  x398 &  x404 &  x419 &  x425 &  x427 &  x431 &  x443 &  x452 &  x455 &  x466 &  x467 &  x482 &  x485 &  x493 &  x503 &  x506 &  x524 &  x527 &  x530 &  x532 &  x536 &  x542 &  x557 &  x560 &  x563 &  x569 &  x572 &  x575 &  x578 &  x584 &  x587 &  x590 &  x596 &  x608 &  x611 &  x623 &  x632 &  x647 &  x653 &  x656 &  x662 &  x667 &  x671 &  x673 &  x674 &  x680 &  x698 &  x701 &  x704 &  x719 &  x749 &  x755 &  x758 &  x764 &  x773 &  x785 &  x800 &  x815 &  x824 &  x827 &  x839 &  x845 &  x851 &  x860 &  x866 &  x884 &  x887 &  x917 &  x920 &  x935 &  x941 &  x944 &  x950 &  x971 &  x980 &  x989 &  x995 &  x1001 &  x1016 &  x1019 &  x1037 &  x1040 &  x1043 &  x1046 &  x1055 &  x1058 &  x1064 &  x1079 &  x1088 &  x1097 &  x1106 & ~x273 & ~x312 & ~x639 & ~x678 & ~x717;
assign c6218 =  x14 &  x53 &  x76 &  x77 &  x128 &  x203 &  x212 &  x218 &  x290 &  x326 &  x395 &  x419 &  x458 &  x482 &  x494 &  x500 &  x563 &  x602 &  x605 &  x622 &  x661 &  x680 &  x688 &  x692 &  x704 &  x728 &  x746 &  x772 &  x779 &  x785 &  x830 &  x832 &  x844 &  x845 &  x848 &  x889 &  x968 &  x980 &  x1033 &  x1051 &  x1073 &  x1103 & ~x405 & ~x549 & ~x588 & ~x861;
assign c6220 =  x2 &  x35 &  x89 &  x101 &  x119 &  x122 &  x164 &  x194 &  x197 &  x203 &  x230 &  x278 &  x356 &  x359 &  x371 &  x374 &  x395 &  x434 &  x452 &  x482 &  x500 &  x503 &  x548 &  x551 &  x557 &  x560 &  x584 &  x623 &  x644 &  x647 &  x677 &  x680 &  x692 &  x698 &  x713 &  x722 &  x725 &  x737 &  x746 &  x806 &  x824 &  x881 &  x884 &  x968 &  x986 &  x998 &  x1022 &  x1031 &  x1034 &  x1043 &  x1079 &  x1124 &  x1127 & ~x0 & ~x60 & ~x78 & ~x132 & ~x210 & ~x249 & ~x288 & ~x327 & ~x405 & ~x444 & ~x483 & ~x672 & ~x750 & ~x789 & ~x807 & ~x828 & ~x936;
assign c6222 =  x4 &  x22 &  x40 &  x43 &  x44 &  x71 &  x73 &  x77 &  x82 &  x86 &  x100 &  x110 &  x112 &  x122 &  x131 &  x139 &  x146 &  x151 &  x160 &  x164 &  x197 &  x203 &  x224 &  x229 &  x248 &  x257 &  x268 &  x307 &  x346 &  x374 &  x377 &  x401 &  x422 &  x476 &  x494 &  x502 &  x524 &  x532 &  x536 &  x539 &  x551 &  x566 &  x581 &  x587 &  x590 &  x619 &  x623 &  x635 &  x638 &  x650 &  x671 &  x674 &  x695 &  x716 &  x719 &  x731 &  x758 &  x764 &  x785 &  x814 &  x845 &  x851 &  x853 &  x872 &  x875 &  x884 &  x890 &  x892 &  x899 &  x931 &  x947 &  x953 &  x956 &  x958 &  x959 &  x965 &  x977 &  x1004 &  x1019 &  x1028 &  x1031 &  x1064 &  x1079 &  x1091 &  x1097 &  x1106 & ~x471 & ~x510 & ~x549;
assign c6224 =  x76 &  x284 &  x569 &  x722 &  x889 &  x899 &  x920 &  x973 &  x998 & ~x210 & ~x327 & ~x483 & ~x627 & ~x1093;
assign c6226 =  x14 &  x32 &  x77 &  x185 &  x275 &  x284 &  x326 &  x337 &  x343 &  x374 &  x376 &  x419 &  x421 &  x427 &  x458 &  x460 &  x466 &  x491 &  x499 &  x503 &  x683 &  x692 &  x706 &  x761 &  x788 &  x833 &  x866 &  x920 &  x989 &  x992 &  x995 &  x1013 &  x1022 &  x1064 &  x1079 &  x1091 & ~x345 & ~x597 & ~x636 & ~x969;
assign c6228 =  x14 &  x17 &  x50 &  x62 &  x65 &  x74 &  x77 &  x122 &  x128 &  x170 &  x176 &  x191 &  x197 &  x227 &  x239 &  x281 &  x292 &  x308 &  x311 &  x317 &  x326 &  x337 &  x338 &  x350 &  x374 &  x386 &  x419 &  x461 &  x482 &  x515 &  x536 &  x557 &  x569 &  x587 &  x593 &  x620 &  x647 &  x650 &  x677 &  x725 &  x764 &  x784 &  x788 &  x800 &  x818 &  x830 &  x833 &  x845 &  x884 &  x893 &  x899 &  x944 &  x979 &  x992 &  x1001 &  x1018 &  x1055 &  x1057 &  x1064 &  x1085 &  x1088 &  x1091 &  x1118 &  x1127 & ~x399 & ~x600 & ~x639 & ~x714 & ~x903;
assign c6230 =  x22 &  x41 &  x59 &  x67 &  x80 &  x83 &  x139 &  x145 &  x164 &  x184 &  x190 &  x200 &  x217 &  x256 &  x301 &  x305 &  x346 &  x347 &  x401 &  x424 &  x476 &  x491 &  x503 &  x563 &  x587 &  x590 &  x619 &  x650 &  x680 &  x685 &  x724 &  x764 &  x769 &  x779 &  x800 &  x841 &  x947 &  x958 &  x974 &  x1022 &  x1079 & ~x285 & ~x402 & ~x1032 & ~x1065;
assign c6232 =  x17 &  x23 &  x26 &  x56 &  x68 &  x77 &  x86 &  x89 &  x101 &  x110 &  x119 &  x122 &  x128 &  x134 &  x137 &  x140 &  x152 &  x154 &  x164 &  x167 &  x170 &  x176 &  x179 &  x188 &  x197 &  x203 &  x215 &  x236 &  x254 &  x269 &  x275 &  x287 &  x308 &  x317 &  x347 &  x355 &  x368 &  x371 &  x392 &  x395 &  x404 &  x407 &  x413 &  x416 &  x425 &  x428 &  x431 &  x433 &  x455 &  x458 &  x464 &  x472 &  x479 &  x485 &  x491 &  x494 &  x503 &  x515 &  x518 &  x536 &  x545 &  x554 &  x563 &  x599 &  x611 &  x635 &  x647 &  x650 &  x668 &  x674 &  x677 &  x686 &  x689 &  x701 &  x721 &  x722 &  x728 &  x746 &  x755 &  x758 &  x760 &  x761 &  x785 &  x799 &  x800 &  x803 &  x806 &  x833 &  x851 &  x881 &  x884 &  x896 &  x902 &  x920 &  x929 &  x935 &  x944 &  x947 &  x968 &  x980 &  x983 &  x986 &  x989 &  x1001 &  x1007 &  x1028 &  x1040 &  x1046 &  x1055 &  x1079 &  x1085 &  x1097 &  x1106 &  x1121 &  x1130 & ~x285 & ~x324 & ~x363 & ~x364 & ~x366 & ~x402 & ~x405 & ~x441 & ~x444 & ~x480 & ~x663 & ~x666 & ~x702;
assign c6234 =  x8 &  x26 &  x32 &  x41 &  x47 &  x80 &  x83 &  x89 &  x92 &  x98 &  x110 &  x119 &  x128 &  x131 &  x143 &  x146 &  x149 &  x164 &  x176 &  x188 &  x191 &  x197 &  x203 &  x206 &  x239 &  x266 &  x269 &  x275 &  x278 &  x302 &  x311 &  x350 &  x353 &  x374 &  x380 &  x431 &  x434 &  x443 &  x449 &  x467 &  x482 &  x485 &  x488 &  x491 &  x521 &  x536 &  x539 &  x542 &  x557 &  x569 &  x572 &  x587 &  x589 &  x632 &  x644 &  x650 &  x659 &  x665 &  x668 &  x686 &  x707 &  x710 &  x713 &  x722 &  x745 &  x749 &  x764 &  x770 &  x784 &  x800 &  x806 &  x812 &  x824 &  x833 &  x848 &  x866 &  x869 &  x908 &  x917 &  x947 &  x959 &  x962 &  x968 &  x986 &  x995 &  x1001 &  x1025 &  x1028 &  x1055 &  x1061 &  x1079 &  x1091 &  x1103 &  x1109 &  x1121 & ~x321 & ~x405 & ~x484 & ~x513 & ~x522 & ~x552 & ~x561 & ~x600 & ~x639 & ~x640;
assign c6236 =  x11 &  x20 &  x38 &  x53 &  x71 &  x80 &  x89 &  x95 &  x104 &  x110 &  x116 &  x122 &  x137 &  x146 &  x149 &  x155 &  x164 &  x167 &  x179 &  x194 &  x203 &  x209 &  x218 &  x221 &  x259 &  x293 &  x308 &  x311 &  x329 &  x338 &  x343 &  x376 &  x377 &  x382 &  x386 &  x395 &  x398 &  x415 &  x419 &  x421 &  x422 &  x427 &  x437 &  x454 &  x460 &  x466 &  x473 &  x476 &  x482 &  x491 &  x493 &  x499 &  x506 &  x521 &  x524 &  x532 &  x544 &  x563 &  x569 &  x572 &  x583 &  x587 &  x596 &  x611 &  x622 &  x644 &  x647 &  x650 &  x659 &  x668 &  x671 &  x686 &  x689 &  x703 &  x719 &  x722 &  x737 &  x743 &  x745 &  x758 &  x782 &  x784 &  x791 &  x824 &  x833 &  x845 &  x866 &  x908 &  x920 &  x932 &  x959 &  x974 &  x980 &  x989 &  x1016 &  x1031 &  x1034 &  x1061 &  x1079 &  x1085 &  x1088 &  x1097 &  x1127 &  x1130 & ~x675 & ~x714 & ~x753 & ~x756 & ~x792 & ~x831;
assign c6238 =  x230 &  x287 &  x337 &  x503 &  x713 &  x728 &  x784 &  x800 &  x923 &  x979 &  x1057 & ~x399 & ~x438 & ~x600 & ~x639 & ~x714 & ~x756 & ~x942 & ~x948 & ~x981 & ~x987 & ~x1026;
assign c6240 =  x2 &  x7 &  x23 &  x46 &  x77 &  x221 &  x230 &  x242 &  x269 &  x326 &  x358 &  x359 &  x376 &  x388 &  x397 &  x398 &  x427 &  x466 &  x500 &  x518 &  x557 &  x728 &  x749 &  x827 &  x851 &  x901 &  x940 &  x986 &  x989 &  x992 & ~x0 & ~x117 & ~x234 & ~x273 & ~x522 & ~x561 & ~x600 & ~x639 & ~x678;
assign c6242 =  x17 &  x23 &  x170 &  x440 &  x512 &  x590 &  x661 &  x692 &  x698 &  x700 &  x800 &  x965 &  x1016 &  x1034 &  x1055 &  x1067 &  x1085 & ~x321 & ~x360 & ~x399 & ~x432 & ~x438 & ~x516 & ~x708 & ~x753 & ~x792 & ~x831 & ~x948 & ~x981 & ~x1026 & ~x1065;
assign c6244 =  x110 &  x143 &  x167 &  x197 &  x410 &  x416 &  x431 &  x518 &  x530 &  x551 &  x622 &  x641 &  x644 &  x661 &  x698 &  x740 &  x800 &  x809 &  x812 &  x899 &  x995 &  x1022 &  x1031 &  x1091 &  x1109 & ~x48 & ~x69 & ~x204 & ~x708 & ~x747 & ~x825 & ~x942 & ~x981 & ~x1059 & ~x1083;
assign c6246 =  x92 &  x98 &  x100 &  x101 &  x256 &  x449 &  x479 &  x509 &  x563 &  x610 &  x649 &  x650 &  x685 &  x707 &  x722 &  x730 &  x769 &  x791 &  x830 &  x932 &  x980 &  x986 & ~x84 & ~x162 & ~x201 & ~x285 & ~x441 & ~x588 & ~x666 & ~x747 & ~x825 & ~x942 & ~x1020;
assign c6248 =  x14 &  x23 &  x35 &  x47 &  x80 &  x110 &  x116 &  x128 &  x137 &  x152 &  x167 &  x233 &  x242 &  x269 &  x278 &  x287 &  x296 &  x302 &  x347 &  x350 &  x356 &  x371 &  x380 &  x386 &  x398 &  x407 &  x415 &  x452 &  x466 &  x479 &  x518 &  x532 &  x533 &  x542 &  x554 &  x575 &  x577 &  x602 &  x605 &  x622 &  x629 &  x644 &  x647 &  x668 &  x680 &  x692 &  x698 &  x710 &  x740 &  x761 &  x764 &  x788 &  x800 &  x823 &  x836 &  x845 &  x848 &  x860 &  x862 &  x866 &  x884 &  x893 &  x901 &  x902 &  x905 &  x929 &  x940 &  x944 &  x947 &  x953 &  x959 &  x968 &  x979 &  x980 &  x1001 &  x1016 &  x1019 &  x1028 &  x1057 &  x1079 &  x1127 & ~x393 & ~x429 & ~x432 & ~x471 & ~x510 & ~x549 & ~x753 & ~x756 & ~x792 & ~x795;
assign c6250 =  x11 &  x142 &  x143 &  x164 &  x179 &  x275 &  x336 &  x343 &  x376 &  x388 &  x500 &  x535 &  x851 &  x886 &  x901 &  x902 &  x907 &  x908 &  x940 &  x1100;
assign c6252 =  x83 &  x131 &  x239 &  x277 &  x308 &  x347 &  x350 &  x355 &  x386 &  x395 &  x398 &  x437 &  x449 &  x464 &  x470 &  x530 &  x539 &  x686 &  x689 &  x692 &  x695 &  x707 &  x721 &  x725 &  x731 &  x733 &  x754 &  x760 &  x764 &  x770 &  x772 &  x788 &  x793 &  x799 &  x809 &  x824 &  x830 &  x832 &  x871 &  x889 &  x920 &  x926 &  x968 &  x992 &  x1001 &  x1037 &  x1079 & ~x132 & ~x171 & ~x210 & ~x249 & ~x264 & ~x477 & ~x507 & ~x546 & ~x588 & ~x627;
assign c6254 =  x347 &  x680 &  x755 &  x782 & ~x321 & ~x360 & ~x399 & ~x441 & ~x591 & ~x597 & ~x714 & ~x747 & ~x753 & ~x792 & ~x831 & ~x942 & ~x981 & ~x1099;
assign c6256 =  x76 &  x80 &  x89 &  x116 &  x176 &  x215 &  x218 &  x227 &  x272 &  x277 &  x299 &  x353 &  x355 &  x395 &  x419 &  x440 &  x455 &  x479 &  x491 &  x605 &  x626 &  x649 &  x650 &  x688 &  x725 &  x731 &  x755 &  x824 &  x827 &  x842 &  x881 &  x908 &  x926 &  x929 &  x959 &  x1004 &  x1055 & ~x0 & ~x249 & ~x288 & ~x555 & ~x594 & ~x625;
assign c6258 =  x2 &  x11 &  x14 &  x23 &  x35 &  x56 &  x68 &  x83 &  x86 &  x92 &  x101 &  x113 &  x116 &  x137 &  x146 &  x149 &  x152 &  x167 &  x194 &  x197 &  x215 &  x239 &  x248 &  x257 &  x266 &  x332 &  x335 &  x350 &  x356 &  x359 &  x362 &  x377 &  x380 &  x386 &  x413 &  x419 &  x425 &  x431 &  x446 &  x452 &  x515 &  x521 &  x536 &  x539 &  x545 &  x548 &  x551 &  x563 &  x569 &  x572 &  x575 &  x578 &  x584 &  x590 &  x593 &  x611 &  x626 &  x632 &  x638 &  x662 &  x674 &  x704 &  x719 &  x734 &  x743 &  x746 &  x758 &  x764 &  x767 &  x770 &  x773 &  x800 &  x827 &  x842 &  x845 &  x848 &  x851 &  x857 &  x860 &  x863 &  x881 &  x884 &  x905 &  x920 &  x923 &  x929 &  x935 &  x944 &  x947 &  x953 &  x962 &  x968 &  x974 &  x992 &  x995 &  x998 &  x1001 &  x1016 &  x1019 &  x1031 &  x1046 &  x1058 &  x1064 &  x1085 &  x1091 &  x1097 &  x1106 &  x1109 &  x1112 & ~x198 & ~x327 & ~x522 & ~x558 & ~x597 & ~x636 & ~x714 & ~x753 & ~x756 & ~x792 & ~x795 & ~x831 & ~x834 & ~x870 & ~x909 & ~x942 & ~x948 & ~x987 & ~x1026;
assign c6260 =  x5 &  x8 &  x11 &  x32 &  x35 &  x38 &  x41 &  x53 &  x71 &  x77 &  x83 &  x92 &  x119 &  x140 &  x146 &  x149 &  x152 &  x164 &  x167 &  x176 &  x197 &  x200 &  x227 &  x269 &  x278 &  x293 &  x302 &  x308 &  x335 &  x347 &  x350 &  x374 &  x398 &  x404 &  x422 &  x431 &  x437 &  x500 &  x503 &  x536 &  x551 &  x554 &  x557 &  x563 &  x566 &  x590 &  x602 &  x607 &  x623 &  x632 &  x635 &  x644 &  x650 &  x668 &  x677 &  x692 &  x707 &  x710 &  x713 &  x722 &  x731 &  x734 &  x740 &  x746 &  x761 &  x788 &  x800 &  x809 &  x827 &  x830 &  x851 &  x856 &  x881 &  x887 &  x920 &  x935 &  x944 &  x956 &  x968 &  x971 &  x998 &  x1001 &  x1010 &  x1019 &  x1022 &  x1028 &  x1037 &  x1055 &  x1079 &  x1085 &  x1097 &  x1124 & ~x54 & ~x93 & ~x132 & ~x171 & ~x210 & ~x249 & ~x327 & ~x366 & ~x462 & ~x483 & ~x522 & ~x891 & ~x930 & ~x1086 & ~x1119 & ~x1125;
assign c6262 =  x14 &  x35 &  x110 &  x122 &  x142 &  x158 &  x167 &  x173 &  x227 &  x230 &  x232 &  x239 &  x308 &  x326 &  x332 &  x353 &  x395 &  x407 &  x440 &  x470 &  x503 &  x557 &  x569 &  x590 &  x650 &  x677 &  x686 &  x692 &  x694 &  x698 &  x707 &  x722 &  x733 &  x788 &  x806 &  x845 &  x851 &  x899 &  x920 &  x944 &  x947 &  x950 &  x962 &  x980 &  x986 &  x992 &  x995 &  x1016 &  x1049 &  x1079 &  x1085 &  x1127 & ~x480 & ~x481 & ~x519 & ~x525 & ~x597;
assign c6264 =  x2 &  x32 &  x35 &  x53 &  x56 &  x74 &  x77 &  x80 &  x83 &  x95 &  x98 &  x116 &  x122 &  x137 &  x143 &  x158 &  x161 &  x167 &  x176 &  x194 &  x197 &  x221 &  x224 &  x236 &  x245 &  x254 &  x269 &  x281 &  x287 &  x308 &  x311 &  x326 &  x329 &  x332 &  x335 &  x338 &  x350 &  x356 &  x359 &  x374 &  x380 &  x389 &  x404 &  x419 &  x425 &  x431 &  x437 &  x449 &  x458 &  x476 &  x485 &  x491 &  x509 &  x515 &  x518 &  x530 &  x536 &  x563 &  x566 &  x569 &  x572 &  x575 &  x581 &  x590 &  x602 &  x620 &  x638 &  x647 &  x677 &  x680 &  x689 &  x692 &  x695 &  x701 &  x704 &  x707 &  x710 &  x713 &  x719 &  x722 &  x737 &  x743 &  x770 &  x773 &  x779 &  x782 &  x785 &  x794 &  x809 &  x827 &  x839 &  x845 &  x851 &  x857 &  x866 &  x869 &  x878 &  x899 &  x914 &  x917 &  x920 &  x923 &  x926 &  x932 &  x947 &  x956 &  x962 &  x971 &  x977 &  x986 &  x1016 &  x1028 &  x1040 &  x1043 &  x1076 &  x1079 &  x1097 &  x1112 &  x1118 &  x1121 &  x1124 & ~x165 & ~x204 & ~x210 & ~x327 & ~x363 & ~x366 & ~x441 & ~x444 & ~x480 & ~x483 & ~x522 & ~x558 & ~x561 & ~x600 & ~x675 & ~x714 & ~x753 & ~x792 & ~x831 & ~x1080 & ~x1101 & ~x1119;
assign c6266 =  x29 &  x47 &  x53 &  x89 &  x140 &  x176 &  x221 &  x242 &  x257 &  x293 &  x326 &  x398 &  x431 &  x437 &  x449 &  x452 &  x485 &  x524 &  x532 &  x536 &  x571 &  x581 &  x602 &  x610 &  x638 &  x644 &  x665 &  x689 &  x707 &  x725 &  x770 &  x773 &  x800 &  x824 &  x833 &  x836 &  x839 &  x841 &  x848 &  x851 &  x860 &  x890 &  x899 &  x902 &  x959 &  x986 &  x1016 &  x1028 &  x1031 &  x1079 &  x1088 &  x1097 &  x1124 & ~x90 & ~x96 & ~x135 & ~x225 & ~x246 & ~x363 & ~x402 & ~x789 & ~x945 & ~x1020 & ~x1023 & ~x1059;
assign c6268 =  x11 &  x14 &  x20 &  x32 &  x38 &  x53 &  x68 &  x71 &  x92 &  x110 &  x119 &  x122 &  x128 &  x131 &  x155 &  x176 &  x197 &  x203 &  x224 &  x227 &  x230 &  x278 &  x302 &  x350 &  x380 &  x386 &  x394 &  x395 &  x419 &  x433 &  x434 &  x443 &  x452 &  x479 &  x482 &  x509 &  x515 &  x518 &  x536 &  x554 &  x569 &  x587 &  x620 &  x650 &  x665 &  x680 &  x710 &  x713 &  x746 &  x752 &  x758 &  x773 &  x785 &  x799 &  x812 &  x839 &  x845 &  x860 &  x884 &  x902 &  x908 &  x911 &  x941 &  x947 &  x968 &  x974 &  x997 &  x1004 &  x1022 &  x1088 &  x1097 &  x1106 & ~x48 & ~x171 & ~x288 & ~x402 & ~x408;
assign c6270 =  x35 &  x46 &  x98 &  x128 &  x164 &  x176 &  x227 &  x257 &  x308 &  x395 &  x431 &  x536 &  x620 &  x635 &  x680 &  x799 &  x809 &  x827 &  x833 &  x884 &  x904 &  x908 &  x943 &  x959 &  x994 &  x1022 &  x1027 &  x1072 &  x1079 &  x1106 &  x1111 & ~x78 & ~x210 & ~x249 & ~x406 & ~x522;
assign c6272 =  x11 &  x28 &  x32 &  x41 &  x47 &  x53 &  x56 &  x68 &  x77 &  x86 &  x100 &  x101 &  x122 &  x137 &  x139 &  x140 &  x149 &  x172 &  x176 &  x178 &  x179 &  x188 &  x191 &  x197 &  x209 &  x218 &  x269 &  x295 &  x296 &  x299 &  x301 &  x302 &  x308 &  x314 &  x326 &  x347 &  x350 &  x356 &  x371 &  x374 &  x380 &  x386 &  x392 &  x395 &  x404 &  x419 &  x422 &  x443 &  x449 &  x461 &  x479 &  x482 &  x491 &  x500 &  x503 &  x521 &  x524 &  x533 &  x536 &  x545 &  x569 &  x572 &  x581 &  x584 &  x587 &  x593 &  x602 &  x665 &  x677 &  x686 &  x692 &  x695 &  x704 &  x713 &  x722 &  x728 &  x740 &  x743 &  x746 &  x755 &  x758 &  x761 &  x764 &  x767 &  x770 &  x773 &  x785 &  x788 &  x800 &  x812 &  x839 &  x845 &  x848 &  x869 &  x880 &  x884 &  x887 &  x893 &  x902 &  x920 &  x923 &  x926 &  x932 &  x938 &  x947 &  x977 &  x980 &  x983 &  x992 &  x995 &  x998 &  x1001 &  x1013 &  x1016 &  x1019 &  x1022 &  x1028 &  x1034 &  x1055 &  x1061 &  x1085 &  x1088 &  x1097 &  x1103 &  x1106 &  x1127 & ~x312 & ~x483 & ~x522 & ~x561 & ~x600 & ~x639 & ~x642;
assign c6274 =  x8 &  x32 &  x50 &  x257 &  x284 &  x353 &  x455 &  x461 &  x532 &  x571 &  x610 &  x688 &  x689 &  x902 &  x947 &  x968 &  x1088 &  x1106 & ~x57 & ~x84 & ~x96 & ~x135 & ~x213 & ~x399 & ~x864 & ~x870 & ~x903 & ~x948 & ~x987 & ~x1059 & ~x1065 & ~x1116;
assign c6276 =  x8 &  x14 &  x23 &  x32 &  x71 &  x77 &  x83 &  x92 &  x110 &  x119 &  x134 &  x146 &  x152 &  x155 &  x158 &  x167 &  x194 &  x203 &  x215 &  x236 &  x239 &  x242 &  x248 &  x260 &  x266 &  x272 &  x275 &  x284 &  x308 &  x332 &  x337 &  x343 &  x353 &  x374 &  x376 &  x377 &  x380 &  x382 &  x388 &  x395 &  x415 &  x419 &  x421 &  x422 &  x427 &  x443 &  x452 &  x454 &  x460 &  x464 &  x466 &  x482 &  x491 &  x493 &  x499 &  x503 &  x532 &  x536 &  x539 &  x542 &  x569 &  x587 &  x590 &  x608 &  x622 &  x632 &  x650 &  x653 &  x680 &  x683 &  x692 &  x698 &  x706 &  x716 &  x725 &  x728 &  x731 &  x734 &  x737 &  x743 &  x745 &  x746 &  x755 &  x758 &  x761 &  x779 &  x784 &  x788 &  x803 &  x823 &  x836 &  x845 &  x862 &  x866 &  x881 &  x884 &  x893 &  x896 &  x923 &  x926 &  x935 &  x944 &  x947 &  x959 &  x962 &  x968 &  x971 &  x974 &  x977 &  x998 &  x1001 &  x1016 &  x1022 &  x1034 &  x1079 &  x1103 &  x1130 & ~x678 & ~x714 & ~x717 & ~x753 & ~x756;
assign c6278 =  x8 &  x14 &  x32 &  x47 &  x56 &  x83 &  x89 &  x101 &  x110 &  x116 &  x122 &  x140 &  x146 &  x149 &  x167 &  x179 &  x194 &  x197 &  x221 &  x224 &  x242 &  x260 &  x284 &  x287 &  x302 &  x326 &  x344 &  x350 &  x353 &  x356 &  x365 &  x368 &  x371 &  x380 &  x382 &  x386 &  x388 &  x392 &  x395 &  x398 &  x401 &  x419 &  x421 &  x422 &  x425 &  x460 &  x466 &  x473 &  x479 &  x488 &  x491 &  x494 &  x499 &  x503 &  x538 &  x548 &  x551 &  x563 &  x569 &  x590 &  x602 &  x632 &  x641 &  x644 &  x650 &  x659 &  x668 &  x674 &  x677 &  x689 &  x692 &  x716 &  x719 &  x722 &  x725 &  x731 &  x737 &  x740 &  x746 &  x749 &  x791 &  x794 &  x800 &  x815 &  x824 &  x827 &  x830 &  x833 &  x839 &  x848 &  x872 &  x878 &  x893 &  x899 &  x902 &  x917 &  x920 &  x929 &  x935 &  x941 &  x947 &  x962 &  x968 &  x971 &  x974 &  x983 &  x992 &  x1001 &  x1019 &  x1022 &  x1031 &  x1043 &  x1055 &  x1079 &  x1085 &  x1103 &  x1106 & ~x597 & ~x636 & ~x717 & ~x756 & ~x831 & ~x870 & ~x963;
assign c6280 =  x68 &  x98 &  x101 &  x110 &  x152 &  x185 &  x197 &  x230 &  x284 &  x287 &  x299 &  x326 &  x346 &  x371 &  x382 &  x385 &  x392 &  x395 &  x424 &  x428 &  x434 &  x451 &  x463 &  x491 &  x512 &  x542 &  x554 &  x569 &  x602 &  x611 &  x638 &  x650 &  x653 &  x698 &  x722 &  x740 &  x746 &  x752 &  x782 &  x806 &  x824 &  x842 &  x848 &  x860 &  x866 &  x875 &  x884 &  x899 &  x905 &  x944 &  x959 &  x977 &  x986 &  x1001 &  x1022 &  x1055 &  x1079 &  x1082 & ~x396 & ~x435 & ~x474 & ~x552 & ~x591 & ~x630 & ~x669 & ~x708 & ~x732 & ~x825 & ~x864;
assign c6282 =  x17 &  x65 &  x71 &  x83 &  x92 &  x194 &  x203 &  x218 &  x293 &  x296 &  x314 &  x341 &  x347 &  x368 &  x374 &  x395 &  x494 &  x518 &  x530 &  x560 &  x584 &  x635 &  x677 &  x719 &  x728 &  x770 &  x836 &  x839 &  x842 &  x845 &  x881 &  x884 &  x893 &  x896 &  x899 &  x992 &  x1022 &  x1034 &  x1055 &  x1058 &  x1076 &  x1097 &  x1103 & ~x99 & ~x117 & ~x132 & ~x138 & ~x144 & ~x171 & ~x177 & ~x183 & ~x210 & ~x216 & ~x249 & ~x255 & ~x294 & ~x327 & ~x483 & ~x522 & ~x561 & ~x600 & ~x639 & ~x678 & ~x834 & ~x945 & ~x951 & ~x984;
assign c6284 =  x8 &  x80 &  x128 &  x197 &  x299 &  x302 &  x380 &  x392 &  x398 &  x563 &  x568 &  x647 &  x649 &  x692 &  x722 &  x779 &  x830 &  x866 &  x887 &  x947 &  x959 &  x1106 & ~x132 & ~x171 & ~x345 & ~x483 & ~x522 & ~x795 & ~x834 & ~x873 & ~x942 & ~x951 & ~x1119;
assign c6286 =  x8 &  x62 &  x128 &  x139 &  x178 &  x194 &  x251 &  x257 &  x308 &  x322 &  x326 &  x356 &  x401 &  x431 &  x467 &  x536 &  x557 &  x566 &  x571 &  x602 &  x619 &  x647 &  x677 &  x685 &  x697 &  x713 &  x763 &  x801 &  x812 &  x814 &  x841 &  x878 &  x880 &  x1040 &  x1070 &  x1079 & ~x69;
assign c6288 =  x166 &  x199 &  x272 &  x277 &  x356 &  x371 &  x392 &  x428 &  x536 &  x590 &  x650 &  x760 &  x851 &  x884 &  x947 &  x998 &  x1019 &  x1022 &  x1031 &  x1097 & ~x132 & ~x210 & ~x213 & ~x471 & ~x546 & ~x549 & ~x627 & ~x666 & ~x861;
assign c6290 =  x203 &  x344 &  x355 &  x593 &  x596 &  x623 &  x725 &  x848 &  x944 &  x989 &  x1022 & ~x132 & ~x250 & ~x288 & ~x546 & ~x549 & ~x703 & ~x976 & ~x1092;
assign c6292 =  x50 &  x145 &  x161 &  x167 &  x197 &  x209 &  x260 &  x269 &  x302 &  x314 &  x326 &  x350 &  x425 &  x434 &  x443 &  x542 &  x659 &  x683 &  x725 &  x731 &  x760 &  x797 &  x799 &  x818 &  x848 &  x968 &  x980 &  x992 &  x1001 & ~x57 & ~x96 & ~x162 & ~x408 & ~x447 & ~x459 & ~x666 & ~x942;
assign c6294 =  x38 &  x119 &  x128 &  x176 &  x230 &  x263 &  x278 &  x347 &  x365 &  x377 &  x401 &  x404 &  x446 &  x455 &  x533 &  x587 &  x653 &  x659 &  x673 &  x677 &  x689 &  x722 &  x743 &  x782 &  x800 &  x893 &  x959 &  x962 &  x992 &  x995 &  x1031 &  x1064 &  x1079 &  x1106 & ~x96 & ~x207 & ~x252 & ~x543 & ~x552 & ~x831 & ~x864 & ~x927 & ~x1083;
assign c6296 =  x11 &  x20 &  x26 &  x29 &  x32 &  x38 &  x53 &  x58 &  x77 &  x80 &  x83 &  x89 &  x101 &  x110 &  x113 &  x119 &  x122 &  x125 &  x128 &  x149 &  x155 &  x176 &  x193 &  x194 &  x200 &  x203 &  x206 &  x209 &  x212 &  x232 &  x233 &  x239 &  x242 &  x251 &  x254 &  x260 &  x281 &  x284 &  x287 &  x308 &  x326 &  x338 &  x350 &  x355 &  x374 &  x386 &  x389 &  x394 &  x395 &  x398 &  x404 &  x407 &  x419 &  x433 &  x446 &  x452 &  x482 &  x485 &  x488 &  x491 &  x494 &  x500 &  x503 &  x506 &  x518 &  x548 &  x560 &  x563 &  x587 &  x590 &  x602 &  x605 &  x608 &  x620 &  x635 &  x650 &  x653 &  x659 &  x674 &  x680 &  x686 &  x689 &  x692 &  x695 &  x707 &  x722 &  x725 &  x728 &  x731 &  x746 &  x776 &  x779 &  x788 &  x799 &  x800 &  x809 &  x818 &  x821 &  x830 &  x839 &  x845 &  x848 &  x860 &  x863 &  x878 &  x884 &  x893 &  x896 &  x920 &  x947 &  x953 &  x956 &  x959 &  x968 &  x971 &  x980 &  x986 &  x1001 &  x1022 &  x1025 &  x1043 &  x1055 &  x1072 &  x1079 &  x1085 &  x1097 &  x1100 &  x1112 & ~x78 & ~x402 & ~x405 & ~x441 & ~x444 & ~x480 & ~x483 & ~x522 & ~x702;
assign c6298 =  x23 &  x32 &  x122 &  x176 &  x239 &  x338 &  x455 &  x491 &  x542 &  x590 &  x893 &  x952 &  x1073 & ~x69 & ~x321 & ~x480 & ~x597 & ~x636 & ~x693 & ~x870 & ~x948 & ~x987 & ~x1005 & ~x1044;
assign c61 =  x91 &  x204 &  x274 & ~x531;
assign c63 =  x304 &  x781 &  x859 & ~x777 & ~x817 & ~x960;
assign c65 = ~x688;
assign c67 =  x304 &  x481 & ~x246 & ~x960 & ~x1051 & ~x1111;
assign c69 =  x131 &  x282 & ~x231 & ~x492;
assign c611 =  x68 &  x146 &  x425 &  x445 &  x469 &  x484 &  x521 &  x664 &  x689 &  x704 &  x1080 &  x1097;
assign c613 =  x430 &  x547 &  x666 & ~x81;
assign c615 =  x94 &  x188 &  x195 &  x209 &  x234 & ~x180 & ~x858;
assign c617 =  x484 &  x562 &  x594 &  x601;
assign c619 =  x390 &  x547 & ~x297 & ~x475;
assign c621 =  x484 &  x666 & ~x654;
assign c623 =  x549 &  x744 & ~x1041;
assign c625 =  x109 &  x447 &  x511 &  x601;
assign c627 =  x469 &  x703 & ~x760;
assign c631 =  x274 &  x312 &  x469 & ~x231 & ~x258 & ~x978;
assign c633 =  x37 &  x587 &  x781 &  x859 & ~x699 & ~x804;
assign c635 =  x68 &  x128 &  x398 &  x425 &  x428 &  x511 &  x513 &  x549 &  x599 &  x689 &  x788 &  x989 &  x1067 &  x1088 & ~x390 & ~x429 & ~x546 & ~x1041;
assign c637 =  x352 &  x481 & ~x493;
assign c639 =  x198 &  x516;
assign c641 =  x25 &  x265 &  x1053 & ~x1000;
assign c643 =  x281 &  x563 &  x664 &  x742 &  x890 &  x1013 &  x1021 & ~x576 & ~x723;
assign c645 =  x3 &  x234 &  x592 & ~x220;
assign c647 =  x204 &  x391 & ~x298 & ~x1062;
assign c649 =  x325 &  x637 &  x945 & ~x960 & ~x996;
assign c651 = ~x466;
assign c653 =  x1122 & ~x688;
assign c655 =  x119 &  x187 &  x191 &  x304 &  x523 &  x593 &  x598 &  x956 &  x1070 & ~x648 & ~x660;
assign c657 =  x325 & ~x387 & ~x388 & ~x900;
assign c659 =  x37 &  x200 &  x664 &  x704 &  x770 &  x783 & ~x582 & ~x684;
assign c661 =  x469 & ~x387 & ~x694 & ~x837;
assign c663 =  x109 &  x430 &  x625 &  x664 & ~x495 & ~x837;
assign c665 = ~x670;
assign c667 =  x192 &  x208 &  x487 &  x831;
assign c669 =  x289 &  x367 &  x430 &  x469 & ~x382;
assign c671 =  x474 & ~x84 & ~x100 & ~x141 & ~x351;
assign c673 =  x220 &  x508 &  x663 &  x742 & ~x504;
assign c675 =  x562 &  x586 &  x650 &  x664 &  x710 &  x742 &  x869 &  x1034 &  x1106 & ~x576 & ~x918;
assign c677 = ~x844;
assign c679 =  x313 &  x589 &  x786 & ~x502;
assign c681 =  x17 &  x94 &  x117 &  x128 &  x195 &  x197 &  x234 &  x391 &  x578 &  x650 &  x748 &  x787 &  x794 &  x811 &  x944 &  x953 &  x1112 &  x1115;
assign c683 =  x175 &  x391 & ~x232;
assign c685 = ~x1000;
assign c687 =  x547 &  x742 &  x982 & ~x631;
assign c689 =  x108 &  x109 &  x147 &  x664 &  x703 &  x742;
assign c691 = ~x571 & ~x631;
assign c693 =  x274 &  x352 &  x549 & ~x781;
assign c695 =  x391 & ~x412 & ~x490;
assign c697 =  x204;
assign c699 =  x156 &  x234 &  x471;
assign c6101 = ~x457 & ~x681 & ~x1029;
assign c6103 = ~x415 & ~x901;
assign c6105 = ~x377 & ~x701;
assign c6107 =  x351 & ~x436;
assign c6109 =  x351 & ~x492 & ~x639 & ~x984;
assign c6111 =  x549 &  x744 & ~x465;
assign c6113 =  x523 &  x984;
assign c6115 =  x589 &  x597 &  x714 &  x753;
assign c6117 =  x403 &  x438 &  x442 & ~x573;
assign c6119 =  x109 &  x742 & ~x610;
assign c6121 =  x97 &  x214 &  x481 &  x541 &  x718 &  x1106 & ~x1047;
assign c6123 =  x663 & ~x291 & ~x991 & ~x1030;
assign c6125 =  x757 &  x897 &  x936 &  x1016 & ~x777;
assign c6127 =  x1 &  x234 &  x352 &  x974 & ~x220 & ~x258 & ~x858 & ~x975;
assign c6129 =  x313 &  x430 &  x883 & ~x295;
assign c6131 =  x1021 & ~x142 & ~x163;
assign c6133 =  x25 &  x167 &  x269 &  x347 &  x664 &  x703 &  x742 &  x859 & ~x537 & ~x576 & ~x837;
assign c6135 =  x265 &  x718 &  x936 & ~x787;
assign c6137 =  x549 &  x589 & ~x387 & ~x426 & ~x528;
assign c6139 =  x282 &  x289 &  x469;
assign c6141 = ~x492 & ~x567 & ~x649;
assign c6143 =  x44 &  x287 &  x305 &  x674 &  x742 &  x859 &  x986 &  x1004 &  x1076 & ~x1111 & ~x1113;
assign c6145 =  x80 &  x89 &  x152 &  x233 &  x296 &  x302 &  x356 &  x434 &  x584 &  x614 &  x719 &  x749 &  x797 &  x953 &  x995 &  x1031 &  x1043 &  x1061 &  x1103 & ~x219 & ~x231 & ~x297 & ~x337 & ~x378 & ~x780;
assign c6147 =  x70 &  x744 & ~x621 & ~x918;
assign c6149 =  x265 &  x936 & ~x777 & ~x846;
assign c6151 = ~x4 & ~x895 & ~x1077;
assign c6153 = ~x436;
assign c6155 =  x561 & ~x660;
assign c6157 =  x25 &  x274 &  x289 &  x383 &  x469 &  x797 &  x1007 & ~x342 & ~x381;
assign c6159 =  x70 &  x194 &  x224 &  x484 &  x523 &  x742 &  x859 & ~x648;
assign c6161 =  x481 &  x672 &  x859 & ~x27;
assign c6163 =  x35 &  x55 &  x68 &  x77 &  x92 &  x113 &  x218 &  x274 &  x275 &  x386 &  x431 &  x434 &  x461 &  x536 &  x563 &  x566 &  x611 &  x623 &  x680 &  x704 &  x707 &  x732 &  x734 &  x776 &  x830 &  x839 &  x851 &  x857 &  x860 &  x869 &  x923 &  x944 &  x986 &  x1058 &  x1121 & ~x147;
assign c6165 =  x79 &  x94 &  x234 &  x482 &  x700 & ~x975;
assign c6167 = ~x454 & ~x648 & ~x862 & ~x901;
assign c6169 =  x559 & ~x478 & ~x648;
assign c6171 =  x391 &  x403 & ~x379;
assign c6173 =  x78 &  x234 &  x274 &  x850 &  x929 &  x1025 & ~x102 & ~x103 & ~x180;
assign c6175 =  x79 &  x94 &  x156 &  x234 &  x1060;
assign c6177 =  x715 & ~x142 & ~x280;
assign c6179 =  x510 &  x589 &  x714;
assign c6181 =  x94 &  x234 &  x273 & ~x115;
assign c6183 =  x471 &  x589 &  x753 &  x870;
assign c6185 =  x187 &  x280 &  x403 &  x637 & ~x817;
assign c6187 =  x169 &  x945 & ~x958;
assign c6189 =  x196 &  x234 &  x273 & ~x70 & ~x103;
assign c6191 =  x78 &  x477;
assign c6193 =  x523 & ~x168 & ~x694;
assign c6195 =  x195 &  x235 & ~x36 & ~x717 & ~x780 & ~x984;
assign c6197 =  x541 &  x601 & ~x804 & ~x817;
assign c6199 =  x349 &  x640 &  x898 &  x1101 & ~x804;
assign c6201 =  x133 &  x274 & ~x723 & ~x1041 & ~x1068;
assign c6203 =  x25 &  x523 &  x547 &  x586 & ~x570 & ~x837;
assign c6205 =  x327 &  x391 & ~x421;
assign c6207 =  x549 &  x744 & ~x573;
assign c6209 =  x94 &  x234 &  x248 & ~x148 & ~x291;
assign c6211 =  x586 & ~x388;
assign c6213 =  x265 &  x533 &  x637 &  x704 &  x742 &  x761 &  x781 &  x859 &  x1130 & ~x762;
assign c6215 =  x858 &  x936 & ~x748;
assign c6217 =  x136 &  x483 &  x847;
assign c6219 =  x549 &  x666 &  x744 & ~x117;
assign c6221 =  x274 &  x630 & ~x567 & ~x684 & ~x1029 & ~x1068 & ~x1092;
assign c6223 =  x78 &  x235 &  x313 &  x771 &  x808;
assign c6227 =  x78 &  x194 &  x195 &  x235 &  x269 &  x274 &  x281 &  x313 &  x377 &  x509 &  x548 &  x592 &  x626 &  x668 &  x739 &  x845 &  x899 &  x998 &  x1064 &  x1106 &  x1121 & ~x180 & ~x666 & ~x783 & ~x822 & ~x858;
assign c6229 =  x481 &  x589 &  x859 &  x989 & ~x198 & ~x729;
assign c6231 =  x364 &  x703 & ~x727 & ~x787;
assign c6233 =  x232 &  x457 &  x562 &  x587 &  x604 &  x900 &  x939 & ~x654;
assign c6235 =  x481 &  x598 &  x632 &  x637 &  x676 &  x820 & ~x738 & ~x1035 & ~x1113;
assign c6237 =  x325 &  x481 &  x598 &  x637 & ~x685;
assign c6239 =  x594 &  x598 &  x679;
assign c6241 =  x241 & ~x778 & ~x918 & ~x960;
assign c6243 =  x321 &  x469 & ~x414;
assign c6245 =  x157 &  x471 &  x655 &  x1032;
assign c6247 =  x484 &  x547 &  x586 &  x744 &  x783 &  x1084;
assign c6249 =  x274 &  x430 &  x452 &  x616 & ~x192 & ~x232;
assign c6251 =  x351 & ~x271 & ~x436;
assign c6253 =  x52 &  x406 &  x483 &  x484 &  x496 &  x601 &  x617 &  x679 &  x737 &  x767 &  x1028 &  x1034;
assign c6255 =  x328 &  x430 & ~x343 & ~x378;
assign c6257 =  x561 & ~x291 & ~x727;
assign c6259 =  x55 &  x312 &  x430 & ~x154;
assign c6261 =  x483 &  x1050;
assign c6263 =  x525 & ~x733;
assign c6265 =  x331 &  x945 & ~x1036;
assign c6267 =  x265 &  x364 &  x403 & ~x427;
assign c6269 =  x29 &  x35 &  x50 &  x80 &  x97 &  x131 &  x188 &  x223 &  x248 &  x305 &  x338 &  x500 &  x601 &  x602 &  x701 &  x821 &  x859 &  x905 &  x998 & ~x918;
assign c6271 =  x481 & ~x532;
assign c6273 =  x265 &  x819 &  x897 & ~x661;
assign c6275 =  x265 &  x523 &  x562 &  x742 &  x897 &  x975 & ~x687;
assign c6277 =  x265 &  x592 &  x897 &  x975 & ~x960;
assign c6279 =  x2 &  x86 &  x89 &  x140 &  x146 &  x167 &  x282 &  x455 &  x469 &  x491 &  x508 &  x536 &  x542 &  x547 &  x563 &  x586 &  x625 &  x662 &  x680 &  x707 &  x839 &  x965 &  x1046 &  x1070 &  x1076;
assign c6281 =  x484 & ~x817 & ~x1035;
assign c6283 =  x313 &  x430 & ~x181 & ~x781;
assign c6285 =  x744 & ~x661 & ~x762;
assign c6287 =  x234 &  x391 & ~x114 & ~x180 & ~x262;
assign c6289 =  x147 &  x153 &  x364 &  x442 & ~x957;
assign c6291 =  x364 & ~x388;
assign c6293 =  x195 &  x196 &  x410 &  x434 &  x527 &  x739 & ~x36 & ~x76 & ~x219 & ~x1095;
assign c6295 =  x241 &  x469 & ~x387 & ~x553;
assign c6297 =  x70 &  x897 & ~x648;
assign c6299 = ~x492 & ~x498 & ~x504 & ~x688;
assign c70 =  x5 &  x8 &  x68 &  x257 &  x260 &  x389 &  x404 &  x407 &  x458 &  x521 &  x593 &  x689 &  x740 &  x827 &  x878 &  x890 & ~x387 & ~x426 & ~x673 & ~x712 & ~x751 & ~x765 & ~x828 & ~x829;
assign c72 =  x29 &  x53 &  x65 &  x74 &  x104 &  x125 &  x170 &  x182 &  x196 &  x212 &  x230 &  x239 &  x257 &  x274 &  x281 &  x287 &  x305 &  x312 &  x313 &  x326 &  x341 &  x351 &  x359 &  x362 &  x380 &  x395 &  x407 &  x413 &  x425 &  x431 &  x443 &  x446 &  x469 &  x479 &  x494 &  x518 &  x521 &  x533 &  x568 &  x572 &  x575 &  x581 &  x592 &  x626 &  x638 &  x641 &  x662 &  x671 &  x695 &  x731 &  x773 &  x782 &  x815 &  x818 &  x842 &  x866 &  x935 &  x959 &  x974 &  x995 &  x998 &  x1117 &  x1118 & ~x123 & ~x240;
assign c74 =  x91 &  x128 &  x131 &  x167 &  x282 &  x299 &  x569 &  x580 &  x635 &  x653 &  x658 &  x736 &  x775 &  x809 &  x842 &  x890 &  x1043 & ~x189 & ~x228;
assign c76 =  x2 &  x11 &  x20 &  x26 &  x32 &  x35 &  x80 &  x86 &  x131 &  x140 &  x164 &  x170 &  x173 &  x179 &  x194 &  x197 &  x200 &  x203 &  x209 &  x221 &  x242 &  x245 &  x248 &  x251 &  x260 &  x278 &  x281 &  x287 &  x290 &  x296 &  x350 &  x392 &  x399 &  x401 &  x404 &  x413 &  x419 &  x422 &  x434 &  x438 &  x439 &  x469 &  x470 &  x482 &  x500 &  x503 &  x507 &  x515 &  x524 &  x566 &  x569 &  x572 &  x586 &  x590 &  x593 &  x602 &  x605 &  x611 &  x617 &  x625 &  x632 &  x644 &  x650 &  x662 &  x680 &  x710 &  x716 &  x736 &  x737 &  x764 &  x779 &  x785 &  x809 &  x818 &  x821 &  x827 &  x836 &  x842 &  x854 &  x857 &  x869 &  x872 &  x890 &  x905 &  x920 &  x929 &  x938 &  x941 &  x944 &  x959 &  x965 &  x986 &  x998 &  x1004 &  x1016 &  x1019 &  x1040 &  x1043 &  x1046 &  x1064 &  x1082 &  x1094 &  x1100 & ~x396 & ~x426 & ~x435 & ~x465 & ~x474 & ~x744 & ~x783 & ~x784 & ~x822;
assign c78 =  x104 &  x107 &  x119 &  x185 &  x194 &  x278 &  x320 &  x352 &  x395 &  x419 &  x437 &  x446 &  x536 &  x575 &  x592 &  x596 &  x611 &  x631 &  x638 &  x669 &  x670 &  x708 &  x709 &  x710 &  x747 &  x752 &  x785 &  x818 &  x826 &  x848 &  x865 &  x899 &  x935 &  x959 &  x977 &  x1010 &  x1052 &  x1064 &  x1112 &  x1121 & ~x492 & ~x570 & ~x594 & ~x666 & ~x667 & ~x706 & ~x745 & ~x822 & ~x861;
assign c710 =  x29 &  x35 &  x47 &  x53 &  x83 &  x101 &  x107 &  x131 &  x134 &  x143 &  x146 &  x188 &  x194 &  x203 &  x209 &  x224 &  x245 &  x248 &  x260 &  x269 &  x281 &  x287 &  x311 &  x320 &  x323 &  x335 &  x347 &  x371 &  x377 &  x383 &  x404 &  x416 &  x419 &  x422 &  x467 &  x491 &  x518 &  x520 &  x605 &  x647 &  x656 &  x662 &  x680 &  x686 &  x695 &  x698 &  x734 &  x737 &  x770 &  x779 &  x788 &  x794 &  x797 &  x815 &  x821 &  x857 &  x869 &  x878 &  x890 &  x929 &  x941 &  x1073 &  x1079 &  x1115 & ~x33 & ~x66 & ~x72 & ~x111 & ~x126 & ~x150 & ~x189 & ~x228 & ~x267 & ~x306 & ~x567 & ~x606 & ~x726 & ~x765 & ~x940;
assign c712 =  x8 &  x82 &  x160 &  x172 &  x250 &  x350 &  x428 &  x434 &  x509 &  x601 &  x890 &  x892 &  x931 &  x970 &  x991 &  x1009 &  x1015 &  x1043 & ~x84 & ~x225 & ~x831 & ~x993;
assign c714 =  x41 &  x101 &  x176 &  x209 &  x239 &  x265 &  x286 &  x287 &  x380 &  x440 &  x524 &  x559 &  x581 &  x647 &  x674 &  x719 &  x752 &  x764 &  x779 &  x796 &  x826 &  x864 &  x874 &  x890 &  x903 &  x904 &  x942 &  x943 &  x1013 &  x1016 &  x1106;
assign c716 =  x11 &  x41 &  x49 &  x50 &  x56 &  x65 &  x86 &  x88 &  x157 &  x191 &  x197 &  x209 &  x235 &  x272 &  x335 &  x386 &  x440 &  x446 &  x496 &  x500 &  x503 &  x506 &  x530 &  x535 &  x553 &  x574 &  x590 &  x596 &  x638 &  x650 &  x695 &  x710 &  x734 &  x737 &  x812 &  x818 &  x821 &  x890 &  x911 &  x914 &  x929 &  x959 &  x983 &  x1001 &  x1016 &  x1037 &  x1046 &  x1049 &  x1061 &  x1073 &  x1088 &  x1121 & ~x162 & ~x163 & ~x180 & ~x201 & ~x219 & ~x258 & ~x393 & ~x433 & ~x472 & ~x511 & ~x549 & ~x550 & ~x589 & ~x627 & ~x666;
assign c718 =  x17 &  x26 &  x104 &  x131 &  x221 &  x226 &  x259 &  x260 &  x265 &  x281 &  x298 &  x349 &  x350 &  x376 &  x379 &  x380 &  x416 &  x418 &  x421 &  x457 &  x496 &  x520 &  x535 &  x557 &  x562 &  x638 &  x672 &  x689 &  x716 &  x752 &  x863 &  x890 &  x989 &  x992 &  x1004 & ~x156;
assign c720 =  x179 &  x286 &  x321 &  x324 &  x360 & ~x357 & ~x358 & ~x397 & ~x436 & ~x745;
assign c722 =  x209 &  x328 &  x451 &  x529 &  x535 &  x552 &  x562 &  x574 &  x592 &  x601 &  x640 &  x688 &  x725 &  x890 & ~x546;
assign c724 =  x20 &  x23 &  x47 &  x68 &  x71 &  x89 &  x152 &  x167 &  x194 &  x197 &  x221 &  x230 &  x244 &  x260 &  x266 &  x272 &  x278 &  x281 &  x290 &  x308 &  x314 &  x350 &  x371 &  x374 &  x383 &  x395 &  x398 &  x404 &  x473 &  x494 &  x506 &  x512 &  x536 &  x545 &  x580 &  x584 &  x626 &  x635 &  x653 &  x658 &  x668 &  x686 &  x697 &  x728 &  x736 &  x773 &  x775 &  x782 &  x788 &  x814 &  x833 &  x839 &  x872 &  x902 &  x932 &  x950 &  x956 &  x965 &  x971 &  x980 &  x992 &  x1004 &  x1082 &  x1097 &  x1112 &  x1124 & ~x357 & ~x358 & ~x397 & ~x435 & ~x531 & ~x706 & ~x745 & ~x783;
assign c726 =  x26 &  x35 &  x38 &  x41 &  x59 &  x62 &  x71 &  x86 &  x104 &  x110 &  x116 &  x128 &  x134 &  x137 &  x152 &  x164 &  x194 &  x206 &  x209 &  x239 &  x257 &  x260 &  x266 &  x269 &  x284 &  x290 &  x299 &  x305 &  x308 &  x320 &  x332 &  x344 &  x350 &  x356 &  x362 &  x368 &  x380 &  x386 &  x389 &  x392 &  x401 &  x416 &  x422 &  x428 &  x440 &  x469 &  x470 &  x512 &  x518 &  x524 &  x536 &  x548 &  x557 &  x569 &  x578 &  x584 &  x593 &  x602 &  x611 &  x631 &  x640 &  x641 &  x662 &  x669 &  x670 &  x686 &  x708 &  x709 &  x710 &  x713 &  x725 &  x747 &  x748 &  x758 &  x761 &  x776 &  x782 &  x787 &  x791 &  x797 &  x803 &  x809 &  x815 &  x821 &  x826 &  x827 &  x839 &  x854 &  x860 &  x865 &  x881 &  x884 &  x890 &  x902 &  x908 &  x914 &  x932 &  x935 &  x947 &  x950 &  x959 &  x986 &  x1007 &  x1010 &  x1019 &  x1028 &  x1031 &  x1037 &  x1049 &  x1067 &  x1070 &  x1079 &  x1088 &  x1094 &  x1124 & ~x705 & ~x745;
assign c728 =  x35 &  x44 &  x53 &  x59 &  x83 &  x130 &  x140 &  x143 &  x155 &  x158 &  x166 &  x224 &  x239 &  x245 &  x257 &  x263 &  x266 &  x272 &  x278 &  x293 &  x308 &  x365 &  x430 &  x449 &  x469 &  x488 &  x506 &  x509 &  x515 &  x530 &  x542 &  x562 &  x593 &  x600 &  x601 &  x631 &  x632 &  x640 &  x650 &  x656 &  x670 &  x679 &  x698 &  x701 &  x707 &  x709 &  x718 &  x728 &  x737 &  x833 &  x857 &  x860 &  x872 &  x896 &  x923 &  x941 &  x1001 &  x1055 &  x1085 &  x1100 &  x1109 & ~x240 & ~x279 & ~x666;
assign c730 =  x11 &  x29 &  x35 &  x41 &  x47 &  x74 &  x77 &  x98 &  x101 &  x116 &  x119 &  x131 &  x140 &  x164 &  x179 &  x197 &  x209 &  x281 &  x287 &  x292 &  x317 &  x353 &  x359 &  x370 &  x407 &  x416 &  x439 &  x440 &  x458 &  x461 &  x479 &  x480 &  x503 &  x509 &  x520 &  x524 &  x536 &  x554 &  x559 &  x566 &  x569 &  x572 &  x581 &  x586 &  x590 &  x602 &  x605 &  x620 &  x644 &  x662 &  x671 &  x683 &  x695 &  x710 &  x734 &  x742 &  x755 &  x781 &  x782 &  x791 &  x794 &  x797 &  x815 &  x842 &  x857 &  x869 &  x890 &  x898 &  x902 &  x935 &  x941 &  x970 &  x977 &  x983 &  x992 &  x1013 &  x1016 &  x1019 &  x1037 &  x1043 &  x1046 &  x1064 &  x1067 &  x1070 &  x1076 &  x1103 &  x1115 & ~x940 & ~x979;
assign c732 =  x26 &  x53 &  x74 &  x83 &  x107 &  x134 &  x137 &  x140 &  x146 &  x152 &  x155 &  x167 &  x170 &  x173 &  x209 &  x215 &  x221 &  x248 &  x275 &  x278 &  x293 &  x296 &  x308 &  x314 &  x323 &  x347 &  x383 &  x386 &  x416 &  x422 &  x431 &  x434 &  x467 &  x484 &  x500 &  x506 &  x515 &  x559 &  x562 &  x575 &  x578 &  x581 &  x590 &  x601 &  x640 &  x662 &  x677 &  x689 &  x710 &  x716 &  x725 &  x742 &  x743 &  x794 &  x797 &  x800 &  x809 &  x818 &  x830 &  x845 &  x859 &  x887 &  x897 &  x898 &  x920 &  x936 &  x937 &  x941 &  x975 &  x992 &  x1014 &  x1015 &  x1016 &  x1034 &  x1052 &  x1053 &  x1093 &  x1097 &  x1100 &  x1112 &  x1115 &  x1118 & ~x393 & ~x843 & ~x882 & ~x960 & ~x1089 & ~x1096;
assign c734 =  x9 &  x10 &  x14 &  x44 &  x47 &  x49 &  x59 &  x80 &  x101 &  x122 &  x156 &  x197 &  x230 &  x281 &  x329 &  x473 &  x479 &  x530 &  x548 &  x587 &  x652 &  x686 &  x689 &  x719 &  x803 &  x809 &  x863 &  x926 &  x980 &  x1019 &  x1031 &  x1118 & ~x298 & ~x433 & ~x666;
assign c736 =  x11 &  x26 &  x35 &  x59 &  x71 &  x74 &  x110 &  x125 &  x130 &  x140 &  x155 &  x166 &  x204 &  x239 &  x248 &  x251 &  x274 &  x275 &  x284 &  x317 &  x371 &  x383 &  x391 &  x467 &  x469 &  x473 &  x482 &  x491 &  x530 &  x562 &  x593 &  x617 &  x629 &  x683 &  x692 &  x725 &  x758 &  x782 &  x809 &  x821 &  x833 &  x851 &  x857 &  x863 &  x887 &  x905 &  x914 &  x953 &  x956 &  x959 &  x995 &  x1031 &  x1034 &  x1040 &  x1058 &  x1100 &  x1124 & ~x240 & ~x336 & ~x339 & ~x378 & ~x417;
assign c738 =  x179 &  x272 &  x308 &  x437 &  x440 &  x479 &  x581 &  x626 &  x653 &  x691 &  x695 &  x704 &  x730 &  x767 &  x782 &  x797 &  x800 &  x803 &  x821 &  x845 &  x872 &  x884 &  x935 &  x938 &  x941 &  x953 &  x959 &  x1028 &  x1043 &  x1076 &  x1109 &  x1118 & ~x486 & ~x603 & ~x642 & ~x681 & ~x711 & ~x744 & ~x790 & ~x829 & ~x906 & ~x945 & ~x1011 & ~x1023;
assign c740 =  x17 &  x59 &  x91 &  x107 &  x128 &  x131 &  x157 &  x167 &  x173 &  x194 &  x195 &  x197 &  x274 &  x338 &  x424 &  x491 &  x584 &  x692 &  x707 &  x737 &  x821 &  x1019 & ~x219 & ~x220 & ~x258 & ~x433 & ~x471;
assign c742 =  x83 &  x128 &  x131 &  x146 &  x206 &  x209 &  x227 &  x329 &  x350 &  x365 &  x409 &  x419 &  x448 &  x449 &  x515 &  x584 &  x602 &  x638 &  x644 &  x650 &  x686 &  x725 &  x755 &  x779 &  x782 &  x815 &  x820 &  x833 &  x859 &  x872 &  x881 &  x902 &  x905 &  x944 &  x950 &  x962 &  x970 &  x971 &  x1009 &  x1048 &  x1064 &  x1085 &  x1087 &  x1109 &  x1114 & ~x390 & ~x468 & ~x882 & ~x883 & ~x922 & ~x960 & ~x993;
assign c744 =  x26 &  x29 &  x47 &  x65 &  x77 &  x140 &  x185 &  x188 &  x191 &  x197 &  x200 &  x209 &  x224 &  x254 &  x260 &  x263 &  x278 &  x283 &  x287 &  x308 &  x320 &  x321 &  x352 &  x360 &  x361 &  x368 &  x398 &  x419 &  x422 &  x430 &  x437 &  x439 &  x446 &  x464 &  x469 &  x508 &  x509 &  x524 &  x542 &  x581 &  x590 &  x602 &  x635 &  x647 &  x650 &  x658 &  x697 &  x698 &  x710 &  x736 &  x737 &  x752 &  x764 &  x775 &  x782 &  x785 &  x788 &  x794 &  x797 &  x821 &  x872 &  x884 &  x890 &  x905 &  x923 &  x944 &  x1004 &  x1043 &  x1049 &  x1061 &  x1100 & ~x396 & ~x435 & ~x450 & ~x474 & ~x627 & ~x666 & ~x667 & ~x706 & ~x745 & ~x783 & ~x784;
assign c746 =  x2 &  x26 &  x35 &  x41 &  x47 &  x53 &  x56 &  x77 &  x86 &  x119 &  x128 &  x140 &  x146 &  x179 &  x191 &  x209 &  x233 &  x239 &  x245 &  x248 &  x260 &  x272 &  x278 &  x281 &  x320 &  x398 &  x416 &  x419 &  x422 &  x439 &  x442 &  x446 &  x458 &  x503 &  x509 &  x530 &  x554 &  x586 &  x605 &  x611 &  x644 &  x647 &  x664 &  x686 &  x698 &  x701 &  x703 &  x737 &  x758 &  x781 &  x782 &  x788 &  x791 &  x797 &  x809 &  x818 &  x821 &  x833 &  x848 &  x857 &  x890 &  x905 &  x911 &  x917 &  x929 &  x935 &  x941 &  x983 &  x986 &  x992 &  x1019 &  x1034 &  x1046 &  x1064 &  x1073 &  x1094 &  x1106 &  x1112 &  x1118 & ~x393 & ~x465 & ~x471 & ~x474 & ~x513 & ~x552 & ~x591 & ~x630 & ~x687 & ~x765 & ~x861 & ~x940 & ~x1026 & ~x1065 & ~x1104;
assign c748 =  x203 &  x221 &  x425 &  x439 &  x469 &  x507 &  x508 &  x515 &  x662 &  x779 &  x809 &  x875 &  x890 &  x1007 & ~x189 & ~x228 & ~x687 & ~x745 & ~x784;
assign c750 =  x56 &  x185 &  x209 &  x227 &  x242 &  x317 &  x320 &  x356 &  x449 &  x464 &  x602 &  x626 &  x638 &  x698 &  x878 &  x890 &  x905 &  x980 &  x992 &  x1019 &  x1043 &  x1088 &  x1099 &  x1118 & ~x327 & ~x501 & ~x606 & ~x805 & ~x844 & ~x882 & ~x883;
assign c752 =  x5 &  x23 &  x47 &  x68 &  x74 &  x77 &  x83 &  x89 &  x98 &  x131 &  x152 &  x176 &  x209 &  x215 &  x236 &  x242 &  x248 &  x275 &  x278 &  x293 &  x305 &  x308 &  x335 &  x344 &  x350 &  x428 &  x440 &  x443 &  x452 &  x458 &  x467 &  x473 &  x485 &  x524 &  x542 &  x548 &  x569 &  x584 &  x590 &  x602 &  x608 &  x641 &  x653 &  x662 &  x674 &  x698 &  x710 &  x719 &  x746 &  x758 &  x764 &  x773 &  x812 &  x863 &  x869 &  x890 &  x893 &  x896 &  x905 &  x914 &  x926 &  x929 &  x932 &  x935 &  x938 &  x959 &  x968 &  x971 &  x977 &  x983 &  x1028 &  x1043 &  x1052 &  x1058 &  x1064 &  x1087 &  x1100 &  x1115 &  x1124 & ~x390 & ~x432 & ~x468 & ~x549 & ~x882 & ~x915 & ~x921 & ~x922 & ~x954 & ~x960 & ~x961 & ~x993 & ~x994 & ~x999 & ~x1000 & ~x1033 & ~x1039 & ~x1072 & ~x1077 & ~x1078 & ~x1110 & ~x1111 & ~x1117 & ~x1128;
assign c754 =  x17 &  x23 &  x101 &  x128 &  x173 &  x263 &  x281 &  x383 &  x392 &  x422 &  x427 &  x523 &  x554 &  x634 &  x662 &  x710 &  x740 &  x764 &  x890 &  x941 &  x971 &  x1030 &  x1069 & ~x468 & ~x546 & ~x993 & ~x1033 & ~x1071 & ~x1072 & ~x1077 & ~x1110 & ~x1111 & ~x1117;
assign c756 =  x245 &  x254 &  x377 &  x446 &  x464 &  x470 &  x521 &  x620 &  x669 &  x670 &  x708 &  x747 &  x748 &  x980 &  x1061 & ~x177 & ~x667;
assign c758 =  x41 &  x131 &  x155 &  x194 &  x203 &  x209 &  x212 &  x224 &  x265 &  x335 &  x395 &  x422 &  x446 &  x491 &  x524 &  x581 &  x611 &  x650 &  x662 &  x672 &  x686 &  x710 &  x734 &  x737 &  x755 &  x782 &  x788 &  x821 &  x833 &  x890 &  x941 &  x959 &  x986 &  x1009 &  x1010 &  x1048 &  x1055 &  x1061 &  x1073 &  x1087 &  x1106 & ~x1062 & ~x1101 & ~x1116;
assign c760 =  x182 &  x329 &  x383 &  x596 &  x708 &  x709 &  x747 &  x748 &  x956 &  x1073 & ~x634;
assign c762 =  x35 &  x41 &  x56 &  x65 &  x83 &  x101 &  x140 &  x146 &  x188 &  x212 &  x220 &  x242 &  x245 &  x259 &  x263 &  x278 &  x284 &  x371 &  x398 &  x419 &  x440 &  x445 &  x449 &  x464 &  x482 &  x484 &  x487 &  x503 &  x518 &  x562 &  x575 &  x581 &  x584 &  x590 &  x611 &  x614 &  x635 &  x640 &  x644 &  x662 &  x716 &  x728 &  x758 &  x764 &  x779 &  x785 &  x797 &  x820 &  x821 &  x897 &  x905 &  x917 &  x931 &  x952 &  x959 &  x970 &  x975 &  x991 &  x1014 &  x1030 &  x1034 &  x1053 &  x1069 &  x1079 &  x1092 & ~x312 & ~x393;
assign c764 =  x26 &  x71 &  x86 &  x122 &  x125 &  x131 &  x152 &  x170 &  x179 &  x188 &  x191 &  x194 &  x245 &  x251 &  x284 &  x287 &  x293 &  x317 &  x323 &  x338 &  x347 &  x356 &  x377 &  x383 &  x404 &  x410 &  x422 &  x479 &  x509 &  x584 &  x602 &  x608 &  x617 &  x629 &  x635 &  x650 &  x653 &  x674 &  x677 &  x686 &  x701 &  x710 &  x764 &  x773 &  x785 &  x800 &  x803 &  x821 &  x833 &  x865 &  x904 &  x935 &  x943 &  x953 &  x982 &  x992 &  x1019 &  x1021 &  x1022 &  x1049 &  x1064 &  x1085 &  x1109 &  x1118 & ~x648 & ~x829 & ~x868 & ~x900 & ~x906 & ~x907 & ~x945 & ~x960 & ~x984 & ~x985 & ~x1023 & ~x1062;
assign c766 =  x77 &  x125 &  x131 &  x146 &  x209 &  x226 &  x260 &  x265 &  x287 &  x341 &  x434 &  x455 &  x500 &  x638 &  x647 &  x698 &  x707 &  x890 &  x929 &  x931 &  x941 &  x970 &  x1004 &  x1009 &  x1016 &  x1021 &  x1048 &  x1087 &  x1099 &  x1126 & ~x468 & ~x984 & ~x1023 & ~x1062 & ~x1101;
assign c768 =  x10 &  x17 &  x26 &  x41 &  x44 &  x47 &  x49 &  x77 &  x92 &  x107 &  x119 &  x121 &  x125 &  x131 &  x157 &  x167 &  x173 &  x176 &  x194 &  x209 &  x233 &  x239 &  x257 &  x284 &  x317 &  x350 &  x383 &  x404 &  x416 &  x464 &  x473 &  x484 &  x521 &  x523 &  x562 &  x572 &  x575 &  x584 &  x602 &  x611 &  x640 &  x650 &  x680 &  x686 &  x734 &  x737 &  x770 &  x776 &  x782 &  x806 &  x809 &  x845 &  x863 &  x887 &  x893 &  x917 &  x953 &  x959 &  x989 &  x998 &  x1052 &  x1061 &  x1121 & ~x84 & ~x162 & ~x219 & ~x258 & ~x369 & ~x408 & ~x433 & ~x510 & ~x549;
assign c770 =  x91 &  x128 &  x165 &  x166 &  x204 &  x205 &  x244 &  x365 &  x440 &  x580 &  x617 &  x662 &  x893 &  x914 &  x941 &  x950 &  x1100 & ~x258 & ~x589 & ~x627 & ~x628 & ~x667;
assign c772 =  x56 &  x86 &  x116 &  x131 &  x140 &  x179 &  x191 &  x197 &  x209 &  x224 &  x254 &  x257 &  x278 &  x281 &  x287 &  x329 &  x335 &  x377 &  x383 &  x398 &  x422 &  x491 &  x524 &  x572 &  x590 &  x611 &  x635 &  x644 &  x647 &  x662 &  x716 &  x742 &  x776 &  x794 &  x815 &  x857 &  x865 &  x869 &  x893 &  x904 &  x929 &  x935 &  x941 &  x943 &  x959 &  x982 &  x989 &  x1001 &  x1004 &  x1009 &  x1013 &  x1021 &  x1034 &  x1046 &  x1048 &  x1064 &  x1067 &  x1073 &  x1087 &  x1112 &  x1121 & ~x900 & ~x921 & ~x940 & ~x1018;
assign c774 =  x5 &  x29 &  x53 &  x56 &  x98 &  x107 &  x126 &  x127 &  x149 &  x165 &  x166 &  x196 &  x203 &  x205 &  x221 &  x248 &  x266 &  x302 &  x308 &  x332 &  x352 &  x362 &  x391 &  x392 &  x416 &  x455 &  x458 &  x464 &  x494 &  x563 &  x575 &  x587 &  x623 &  x674 &  x680 &  x719 &  x773 &  x785 &  x791 &  x806 &  x815 &  x857 &  x881 &  x905 &  x920 &  x956 &  x980 &  x1040 &  x1058 &  x1088 &  x1100 &  x1118 & ~x219 & ~x220 & ~x258 & ~x259 & ~x297 & ~x298 & ~x471 & ~x550 & ~x588 & ~x936;
assign c776 =  x88 &  x127 &  x166 &  x170 &  x194 &  x205 &  x317 &  x424 &  x444 &  x458 &  x602 &  x619 &  x658 &  x670 &  x710 &  x757 &  x821 &  x1006 &  x1049;
assign c778 =  x35 &  x91 &  x101 &  x104 &  x173 &  x275 &  x383 &  x395 &  x413 &  x482 &  x494 &  x635 &  x698 &  x709 &  x716 &  x731 &  x752 &  x761 &  x935 &  x992 & ~x744 & ~x777 & ~x856 & ~x933 & ~x960 & ~x972 & ~x1101;
assign c780 =  x49 &  x82 &  x121 &  x398 &  x572 &  x890 &  x928 &  x967 &  x1006 &  x1052 & ~x219 & ~x258 & ~x433 & ~x472 & ~x511 & ~x906;
assign c782 =  x41 &  x47 &  x95 &  x113 &  x122 &  x128 &  x131 &  x158 &  x173 &  x185 &  x194 &  x203 &  x209 &  x212 &  x218 &  x221 &  x239 &  x278 &  x311 &  x321 &  x322 &  x329 &  x332 &  x335 &  x359 &  x360 &  x364 &  x403 &  x434 &  x439 &  x440 &  x446 &  x467 &  x469 &  x509 &  x524 &  x581 &  x602 &  x611 &  x620 &  x623 &  x626 &  x632 &  x668 &  x680 &  x686 &  x707 &  x722 &  x725 &  x737 &  x773 &  x776 &  x779 &  x788 &  x794 &  x800 &  x815 &  x827 &  x830 &  x872 &  x890 &  x920 &  x929 &  x941 &  x959 &  x1013 &  x1040 &  x1055 &  x1064 & ~x357 & ~x450 & ~x666 & ~x706 & ~x745 & ~x822;
assign c784 =  x56 &  x83 &  x86 &  x101 &  x185 &  x188 &  x194 &  x197 &  x209 &  x227 &  x257 &  x284 &  x338 &  x359 &  x364 &  x365 &  x403 &  x422 &  x430 &  x467 &  x469 &  x479 &  x508 &  x557 &  x560 &  x569 &  x601 &  x605 &  x629 &  x635 &  x640 &  x650 &  x662 &  x679 &  x686 &  x695 &  x703 &  x716 &  x752 &  x755 &  x779 &  x782 &  x791 &  x802 &  x815 &  x835 &  x841 &  x842 &  x857 &  x874 &  x890 &  x902 &  x905 &  x917 &  x926 &  x958 &  x986 &  x1019 &  x1061 &  x1070 &  x1073 &  x1112 & ~x573 & ~x705;
assign c786 =  x13 &  x344 &  x574 &  x590 &  x592 &  x601 &  x740 &  x803 &  x836 &  x905 &  x1004 &  x1126 & ~x228 & ~x816;
assign c788 =  x32 &  x38 &  x77 &  x101 &  x131 &  x149 &  x158 &  x167 &  x179 &  x191 &  x209 &  x212 &  x221 &  x224 &  x226 &  x251 &  x257 &  x260 &  x272 &  x287 &  x296 &  x328 &  x362 &  x416 &  x419 &  x439 &  x446 &  x467 &  x477 &  x517 &  x569 &  x572 &  x584 &  x587 &  x635 &  x638 &  x647 &  x659 &  x662 &  x692 &  x716 &  x737 &  x752 &  x755 &  x758 &  x767 &  x781 &  x797 &  x842 &  x881 &  x890 &  x902 &  x929 &  x931 &  x932 &  x935 &  x944 &  x962 &  x970 &  x975 &  x983 &  x992 &  x1004 &  x1009 &  x1014 &  x1015 &  x1016 &  x1043 &  x1046 &  x1052 &  x1053 &  x1054 &  x1061 &  x1070 &  x1087 &  x1092 &  x1100 &  x1118 & ~x354;
assign c790 =  x126 &  x127 &  x165 &  x166 &  x234 &  x569 &  x575 &  x592 &  x983 &  x1006 &  x1013 & ~x589;
assign c792 =  x32 &  x35 &  x53 &  x56 &  x86 &  x92 &  x128 &  x179 &  x191 &  x194 &  x200 &  x203 &  x209 &  x215 &  x224 &  x226 &  x239 &  x265 &  x278 &  x287 &  x302 &  x317 &  x413 &  x440 &  x473 &  x527 &  x551 &  x569 &  x611 &  x617 &  x623 &  x632 &  x647 &  x725 &  x734 &  x755 &  x770 &  x788 &  x806 &  x821 &  x830 &  x860 &  x866 &  x872 &  x890 &  x893 &  x902 &  x905 &  x941 &  x956 &  x986 &  x1004 &  x1037 &  x1049 &  x1061 &  x1073 &  x1091 &  x1094 &  x1115 &  x1118 & ~x94 & ~x132 & ~x133 & ~x177 & ~x189 & ~x216 & ~x294 & ~x984 & ~x1023 & ~x1062 & ~x1101;
assign c794 =  x20 &  x35 &  x41 &  x53 &  x65 &  x77 &  x86 &  x101 &  x104 &  x119 &  x128 &  x131 &  x140 &  x179 &  x191 &  x203 &  x209 &  x212 &  x221 &  x224 &  x242 &  x260 &  x263 &  x278 &  x281 &  x320 &  x335 &  x338 &  x383 &  x398 &  x403 &  x434 &  x442 &  x467 &  x479 &  x491 &  x530 &  x545 &  x572 &  x602 &  x605 &  x611 &  x635 &  x647 &  x686 &  x698 &  x701 &  x710 &  x752 &  x764 &  x775 &  x779 &  x794 &  x821 &  x842 &  x872 &  x902 &  x913 &  x917 &  x929 &  x952 &  x953 &  x957 &  x958 &  x970 &  x983 &  x986 &  x991 &  x996 &  x1004 &  x1009 &  x1010 &  x1016 &  x1019 &  x1030 &  x1043 &  x1046 &  x1048 &  x1052 &  x1064 &  x1067 &  x1069 &  x1073 &  x1094 &  x1106 & ~x687 & ~x726 & ~x900 & ~x901 & ~x940;
assign c796 =  x26 &  x35 &  x41 &  x47 &  x53 &  x56 &  x101 &  x103 &  x148 &  x181 &  x187 &  x194 &  x197 &  x209 &  x226 &  x239 &  x257 &  x260 &  x265 &  x278 &  x302 &  x320 &  x386 &  x428 &  x442 &  x467 &  x470 &  x520 &  x611 &  x686 &  x695 &  x755 &  x764 &  x809 &  x815 &  x818 &  x872 &  x902 &  x908 &  x935 &  x941 &  x944 &  x959 &  x1043 &  x1070 &  x1118 & ~x234 & ~x423 & ~x823;
assign c798 =  x17 &  x35 &  x65 &  x77 &  x91 &  x101 &  x119 &  x179 &  x194 &  x197 &  x209 &  x239 &  x257 &  x290 &  x308 &  x335 &  x428 &  x434 &  x444 &  x445 &  x473 &  x479 &  x483 &  x522 &  x523 &  x561 &  x562 &  x596 &  x600 &  x601 &  x605 &  x626 &  x638 &  x639 &  x640 &  x644 &  x662 &  x678 &  x679 &  x695 &  x716 &  x717 &  x737 &  x752 &  x755 &  x757 &  x761 &  x794 &  x796 &  x800 &  x815 &  x824 &  x896 &  x902 &  x911 &  x926 &  x935 &  x941 &  x944 &  x983 &  x992 &  x1010 &  x1013 &  x1046 &  x1070 &  x1100 &  x1103 & ~x675 & ~x822;
assign c7100 =  x35 &  x56 &  x77 &  x128 &  x182 &  x197 &  x203 &  x209 &  x215 &  x239 &  x260 &  x281 &  x308 &  x350 &  x353 &  x359 &  x383 &  x389 &  x398 &  x413 &  x416 &  x434 &  x439 &  x473 &  x491 &  x539 &  x554 &  x557 &  x569 &  x586 &  x619 &  x638 &  x644 &  x647 &  x658 &  x665 &  x680 &  x686 &  x697 &  x707 &  x719 &  x722 &  x734 &  x736 &  x749 &  x752 &  x775 &  x781 &  x797 &  x820 &  x821 &  x836 &  x839 &  x842 &  x853 &  x892 &  x914 &  x919 &  x929 &  x931 &  x944 &  x958 &  x959 &  x970 &  x983 &  x986 &  x992 &  x1036 &  x1043 &  x1046 &  x1070 &  x1073 &  x1118 & ~x474 & ~x687 & ~x940;
assign c7102 =  x88 &  x116 &  x127 &  x128 &  x293 &  x383 &  x413 &  x416 &  x457 &  x475 &  x491 &  x496 &  x523 &  x535 &  x548 &  x562 &  x574 &  x601 &  x613 &  x640 &  x652 &  x869 &  x884 &  x911 &  x917 &  x986 &  x1118 & ~x33 & ~x177 & ~x258;
assign c7104 =  x32 &  x50 &  x125 &  x131 &  x172 &  x185 &  x250 &  x284 &  x314 &  x328 &  x335 &  x347 &  x398 &  x401 &  x422 &  x428 &  x434 &  x455 &  x562 &  x581 &  x590 &  x601 &  x608 &  x640 &  x644 &  x647 &  x679 &  x718 &  x749 &  x757 &  x788 &  x796 &  x800 &  x802 &  x835 &  x840 &  x841 &  x845 &  x874 &  x875 &  x880 &  x890 &  x892 &  x902 &  x931 &  x958 &  x959 &  x965 &  x991 &  x995 &  x997 &  x1043 &  x1046 &  x1052 &  x1064 &  x1088 &  x1121 & ~x396 & ~x783 & ~x861 & ~x900;
assign c7106 =  x26 &  x35 &  x56 &  x68 &  x77 &  x80 &  x86 &  x125 &  x134 &  x143 &  x155 &  x179 &  x209 &  x281 &  x350 &  x377 &  x383 &  x407 &  x410 &  x413 &  x473 &  x482 &  x497 &  x536 &  x545 &  x551 &  x593 &  x656 &  x734 &  x752 &  x755 &  x779 &  x781 &  x800 &  x815 &  x820 &  x848 &  x866 &  x872 &  x890 &  x917 &  x953 &  x976 &  x983 &  x986 &  x992 &  x1010 &  x1070 &  x1099 &  x1121 & ~x393 & ~x766 & ~x805 & ~x844 & ~x882 & ~x883 & ~x921 & ~x922 & ~x961 & ~x999 & ~x1000 & ~x1039 & ~x1057 & ~x1116;
assign c7108 =  x31 &  x35 &  x47 &  x56 &  x70 &  x83 &  x86 &  x104 &  x113 &  x149 &  x164 &  x179 &  x188 &  x194 &  x209 &  x254 &  x263 &  x278 &  x281 &  x287 &  x292 &  x320 &  x331 &  x335 &  x356 &  x383 &  x398 &  x409 &  x428 &  x440 &  x452 &  x467 &  x487 &  x494 &  x530 &  x554 &  x557 &  x566 &  x572 &  x594 &  x608 &  x633 &  x638 &  x650 &  x662 &  x707 &  x755 &  x764 &  x770 &  x779 &  x785 &  x824 &  x872 &  x881 &  x890 &  x905 &  x911 &  x935 &  x941 &  x968 &  x1070 &  x1073 & ~x762 & ~x1018;
assign c7110 =  x13 &  x89 &  x91 &  x101 &  x212 &  x266 &  x320 &  x335 &  x350 &  x395 &  x413 &  x416 &  x524 &  x569 &  x617 &  x758 &  x782 &  x788 &  x821 &  x851 &  x902 &  x929 &  x950 &  x1010 &  x1043 &  x1049 &  x1052 &  x1073 &  x1106 & ~x258 & ~x297 & ~x433 & ~x472 & ~x819;
assign c7112 =  x35 &  x52 &  x56 &  x91 &  x131 &  x188 &  x230 &  x335 &  x383 &  x467 &  x530 &  x562 &  x592 &  x631 &  x650 &  x737 &  x815 &  x833 &  x884 &  x941 & ~x99 & ~x201 & ~x511 & ~x550 & ~x589;
assign c7114 =  x26 &  x35 &  x86 &  x131 &  x146 &  x221 &  x224 &  x335 &  x359 &  x398 &  x482 &  x569 &  x572 &  x617 &  x626 &  x695 &  x725 &  x752 &  x779 &  x872 &  x874 &  x902 &  x911 &  x1043 &  x1054 &  x1064 &  x1087 &  x1106 & ~x354 & ~x501 & ~x513 & ~x540 & ~x567 & ~x579 & ~x798 & ~x837 & ~x915 & ~x987 & ~x993;
assign c7116 =  x35 &  x47 &  x52 &  x65 &  x83 &  x119 &  x128 &  x137 &  x160 &  x191 &  x194 &  x296 &  x353 &  x359 &  x392 &  x398 &  x413 &  x431 &  x461 &  x470 &  x500 &  x539 &  x553 &  x562 &  x575 &  x635 &  x710 &  x758 &  x815 &  x830 &  x902 &  x923 &  x929 &  x1004 &  x1064 &  x1106 &  x1130 & ~x258 & ~x511 & ~x549 & ~x550 & ~x589 & ~x628 & ~x667;
assign c7118 =  x13 &  x52 &  x53 &  x56 &  x77 &  x91 &  x104 &  x169 &  x209 &  x260 &  x263 &  x269 &  x308 &  x323 &  x365 &  x377 &  x416 &  x473 &  x491 &  x575 &  x587 &  x593 &  x605 &  x623 &  x650 &  x758 &  x794 &  x854 &  x890 &  x896 &  x914 &  x1034 &  x1043 &  x1049 &  x1079 & ~x240 & ~x258 & ~x279 & ~x297 & ~x336 & ~x628 & ~x667 & ~x1014;
assign c7120 =  x110 &  x323 &  x514 &  x553 &  x557 &  x574 &  x580 &  x640 &  x652 &  x680 &  x767 &  x887 &  x928 &  x967 &  x1006 &  x1084 &  x1109 &  x1111 & ~x219 & ~x258 & ~x369 & ~x408;
assign c7122 =  x35 &  x41 &  x56 &  x62 &  x83 &  x128 &  x131 &  x170 &  x179 &  x187 &  x209 &  x220 &  x226 &  x259 &  x263 &  x265 &  x269 &  x298 &  x341 &  x343 &  x350 &  x383 &  x398 &  x440 &  x442 &  x481 &  x491 &  x542 &  x559 &  x569 &  x590 &  x692 &  x710 &  x752 &  x785 &  x815 &  x842 &  x872 &  x929 &  x935 &  x941 &  x944 &  x959 &  x1004 &  x1073 &  x1100 &  x1118 & ~x510 & ~x630 & ~x940 & ~x979;
assign c7124 =  x35 &  x77 &  x83 &  x128 &  x131 &  x170 &  x233 &  x260 &  x265 &  x269 &  x292 &  x335 &  x341 &  x343 &  x350 &  x398 &  x409 &  x443 &  x460 &  x466 &  x487 &  x509 &  x542 &  x620 &  x641 &  x672 &  x686 &  x695 &  x711 &  x752 &  x764 &  x791 &  x806 &  x820 &  x842 &  x859 &  x869 &  x890 &  x898 &  x905 &  x941 &  x959 &  x962 &  x976 &  x995 &  x1028 &  x1043 &  x1054 &  x1064 &  x1127 &  x1130 & ~x390 & ~x468 & ~x546 & ~x960;
assign c7126 =  x191 &  x197 &  x221 &  x251 &  x260 &  x350 &  x467 &  x518 &  x562 &  x677 &  x716 &  x758 &  x796 &  x890 &  x941 &  x1031 &  x1064 & ~x21 & ~x99 & ~x138 & ~x144 & ~x177 & ~x216 & ~x468 & ~x472 & ~x511 & ~x846 & ~x885;
assign c7128 =  x35 &  x41 &  x59 &  x65 &  x92 &  x101 &  x116 &  x128 &  x131 &  x140 &  x179 &  x194 &  x203 &  x209 &  x212 &  x221 &  x224 &  x242 &  x257 &  x260 &  x263 &  x281 &  x287 &  x320 &  x335 &  x359 &  x383 &  x398 &  x434 &  x467 &  x491 &  x524 &  x536 &  x539 &  x548 &  x551 &  x569 &  x593 &  x662 &  x680 &  x686 &  x695 &  x710 &  x716 &  x725 &  x752 &  x755 &  x764 &  x781 &  x820 &  x854 &  x872 &  x884 &  x887 &  x890 &  x902 &  x905 &  x929 &  x941 &  x956 &  x958 &  x959 &  x968 &  x997 &  x1004 &  x1016 &  x1043 &  x1052 &  x1061 &  x1064 &  x1070 &  x1106 &  x1118 & ~x510 & ~x570 & ~x591 & ~x609 & ~x648 & ~x649 & ~x687 & ~x688 & ~x726 & ~x727 & ~x765 & ~x766 & ~x805 & ~x843 & ~x844 & ~x882 & ~x921 & ~x960 & ~x999;
assign c7130 =  x35 &  x41 &  x101 &  x131 &  x187 &  x194 &  x197 &  x209 &  x221 &  x224 &  x226 &  x233 &  x239 &  x242 &  x265 &  x278 &  x281 &  x377 &  x428 &  x455 &  x458 &  x516 &  x524 &  x542 &  x554 &  x569 &  x593 &  x602 &  x617 &  x664 &  x695 &  x701 &  x710 &  x725 &  x734 &  x737 &  x781 &  x791 &  x820 &  x821 &  x848 &  x859 &  x872 &  x890 &  x902 &  x920 &  x929 &  x935 &  x941 &  x959 &  x989 &  x1046 &  x1052 &  x1064 &  x1073 &  x1079 &  x1112 &  x1118 &  x1121 & ~x390 & ~x591 & ~x630 & ~x765 & ~x940 & ~x979;
assign c7132 =  x2 &  x5 &  x41 &  x50 &  x53 &  x56 &  x65 &  x71 &  x77 &  x101 &  x119 &  x131 &  x152 &  x179 &  x209 &  x218 &  x227 &  x245 &  x257 &  x260 &  x278 &  x305 &  x311 &  x329 &  x335 &  x347 &  x392 &  x398 &  x403 &  x410 &  x416 &  x418 &  x440 &  x443 &  x446 &  x449 &  x455 &  x457 &  x467 &  x518 &  x530 &  x536 &  x548 &  x554 &  x562 &  x602 &  x611 &  x620 &  x623 &  x650 &  x686 &  x695 &  x704 &  x710 &  x722 &  x761 &  x767 &  x791 &  x818 &  x821 &  x833 &  x845 &  x857 &  x875 &  x884 &  x902 &  x905 &  x913 &  x914 &  x917 &  x926 &  x929 &  x941 &  x944 &  x951 &  x958 &  x959 &  x965 &  x977 &  x989 &  x990 &  x991 &  x992 &  x998 &  x1030 &  x1052 &  x1070 &  x1079 &  x1091 & ~x837;
assign c7134 =  x41 &  x77 &  x83 &  x125 &  x140 &  x167 &  x179 &  x203 &  x248 &  x274 &  x275 &  x314 &  x391 &  x416 &  x422 &  x440 &  x479 &  x524 &  x530 &  x584 &  x592 &  x601 &  x630 &  x631 &  x640 &  x652 &  x670 &  x691 &  x701 &  x707 &  x709 &  x730 &  x752 &  x809 &  x833 &  x857 &  x941 &  x944 &  x1016 &  x1049 &  x1061 &  x1064 & ~x1107;
assign c7136 =  x4 &  x43 &  x121 &  x134 &  x148 &  x160 &  x179 &  x187 &  x224 &  x254 &  x298 &  x343 &  x434 &  x455 &  x482 &  x518 &  x520 &  x535 &  x542 &  x557 &  x559 &  x563 &  x574 &  x587 &  x593 &  x605 &  x613 &  x668 &  x677 &  x715 &  x770 &  x791 &  x887 &  x892 &  x902 &  x911 &  x947 &  x1037 &  x1048 &  x1052 &  x1069 &  x1070 &  x1085 &  x1087 &  x1094;
assign c7138 =  x10 &  x43 &  x82 &  x83 &  x121 &  x299 &  x314 &  x367 &  x424 &  x613 &  x944 &  x1009 &  x1030 &  x1103 & ~x45 & ~x258;
assign c7140 =  x209 &  x260 &  x287 &  x457 &  x512 &  x857 &  x1031 & ~x6 & ~x27 & ~x60 & ~x84 & ~x189 & ~x945 & ~x1023;
assign c7142 =  x35 &  x41 &  x116 &  x140 &  x148 &  x187 &  x194 &  x209 &  x221 &  x226 &  x239 &  x245 &  x257 &  x260 &  x265 &  x329 &  x335 &  x338 &  x343 &  x362 &  x395 &  x434 &  x439 &  x491 &  x509 &  x516 &  x559 &  x566 &  x569 &  x586 &  x629 &  x647 &  x662 &  x674 &  x695 &  x710 &  x737 &  x755 &  x764 &  x770 &  x781 &  x820 &  x890 &  x898 &  x902 &  x935 &  x937 &  x941 &  x1034 &  x1069 &  x1106;
assign c7144 =  x23 &  x82 &  x95 &  x116 &  x119 &  x121 &  x191 &  x239 &  x257 &  x320 &  x344 &  x350 &  x398 &  x467 &  x530 &  x545 &  x557 &  x590 &  x626 &  x644 &  x650 &  x686 &  x932 &  x935 &  x986 &  x1034 &  x1043 &  x1049 &  x1100 & ~x36 & ~x76 & ~x84 & ~x123 & ~x142 & ~x213 & ~x219 & ~x225 & ~x906 & ~x945;
assign c7146 =  x52 &  x91 &  x130 &  x208 &  x209 &  x230 &  x244 &  x283 &  x580 &  x605 &  x890 &  x929 &  x941 &  x1052 &  x1061 & ~x0 & ~x33 & ~x72 & ~x111 & ~x627 & ~x667 & ~x706 & ~x783;
assign c7148 =  x11 &  x107 &  x131 &  x137 &  x209 &  x273 &  x329 &  x352 &  x407 &  x410 &  x524 &  x590 &  x677 &  x698 &  x787 &  x803 &  x824 &  x842 &  x890 &  x902 &  x956 &  x974 &  x1025 &  x1034 &  x1055 &  x1118 & ~x201 & ~x202 & ~x240 & ~x241 & ~x297 & ~x375 & ~x376 & ~x589 & ~x627 & ~x628;
assign c7150 =  x26 &  x29 &  x35 &  x41 &  x47 &  x86 &  x101 &  x119 &  x155 &  x170 &  x173 &  x191 &  x194 &  x203 &  x209 &  x212 &  x221 &  x248 &  x254 &  x257 &  x266 &  x278 &  x281 &  x311 &  x314 &  x329 &  x335 &  x344 &  x350 &  x359 &  x398 &  x422 &  x440 &  x457 &  x473 &  x476 &  x479 &  x482 &  x491 &  x500 &  x503 &  x614 &  x617 &  x638 &  x686 &  x689 &  x692 &  x695 &  x710 &  x719 &  x737 &  x752 &  x755 &  x779 &  x782 &  x859 &  x872 &  x887 &  x890 &  x898 &  x899 &  x902 &  x905 &  x929 &  x935 &  x937 &  x941 &  x947 &  x970 &  x974 &  x976 &  x983 &  x992 &  x1004 &  x1015 &  x1034 &  x1043 &  x1052 &  x1064 &  x1070 &  x1097 &  x1106 & ~x837 & ~x844 & ~x882 & ~x883 & ~x954 & ~x955 & ~x960 & ~x993 & ~x994 & ~x999 & ~x1033 & ~x1050 & ~x1071;
assign c7152 =  x41 &  x70 &  x103 &  x104 &  x167 &  x383 &  x479 &  x593 &  x653 &  x680 &  x782 &  x785 &  x796 &  x809 &  x848 &  x863 &  x938 &  x953 &  x965 &  x971 &  x992 &  x1004 &  x1061 &  x1076 &  x1112 & ~x306 & ~x411 & ~x628 & ~x706 & ~x745;
assign c7154 =  x56 &  x59 &  x86 &  x209 &  x221 &  x260 &  x263 &  x367 &  x484 &  x497 &  x523 &  x562 &  x569 &  x601 &  x640 &  x719 &  x796 &  x800 &  x809 &  x904 &  x943 & ~x609 & ~x940 & ~x979 & ~x1011 & ~x1050 & ~x1089 & ~x1128;
assign c7156 =  x35 &  x41 &  x47 &  x53 &  x86 &  x101 &  x104 &  x128 &  x131 &  x140 &  x149 &  x188 &  x191 &  x194 &  x197 &  x209 &  x224 &  x239 &  x245 &  x254 &  x260 &  x263 &  x314 &  x335 &  x341 &  x359 &  x364 &  x383 &  x398 &  x403 &  x431 &  x439 &  x467 &  x482 &  x506 &  x509 &  x521 &  x524 &  x539 &  x557 &  x560 &  x563 &  x572 &  x581 &  x626 &  x638 &  x650 &  x662 &  x695 &  x710 &  x713 &  x746 &  x776 &  x781 &  x815 &  x820 &  x821 &  x878 &  x890 &  x902 &  x911 &  x929 &  x935 &  x992 &  x1004 &  x1043 &  x1046 &  x1049 &  x1052 &  x1067 &  x1118 & ~x591 & ~x642 & ~x681 & ~x687 & ~x720 & ~x765 & ~x843 & ~x882 & ~x900 & ~x940 & ~x979;
assign c7158 =  x17 &  x56 &  x68 &  x83 &  x119 &  x128 &  x131 &  x155 &  x179 &  x188 &  x191 &  x194 &  x200 &  x209 &  x212 &  x239 &  x275 &  x281 &  x284 &  x287 &  x290 &  x296 &  x341 &  x353 &  x359 &  x362 &  x365 &  x383 &  x398 &  x416 &  x422 &  x434 &  x440 &  x446 &  x464 &  x491 &  x494 &  x518 &  x521 &  x524 &  x548 &  x569 &  x575 &  x587 &  x593 &  x596 &  x602 &  x611 &  x620 &  x623 &  x632 &  x635 &  x650 &  x662 &  x664 &  x689 &  x695 &  x701 &  x710 &  x725 &  x752 &  x755 &  x764 &  x785 &  x788 &  x821 &  x864 &  x865 &  x872 &  x890 &  x893 &  x896 &  x903 &  x904 &  x905 &  x911 &  x929 &  x935 &  x943 &  x944 &  x959 &  x982 &  x1010 &  x1013 &  x1016 &  x1019 &  x1021 &  x1043 &  x1060 &  x1094 &  x1106 &  x1118 & ~x510 & ~x549 & ~x940;
assign c7160 =  x11 &  x23 &  x35 &  x38 &  x92 &  x104 &  x116 &  x134 &  x146 &  x149 &  x155 &  x179 &  x191 &  x197 &  x209 &  x221 &  x239 &  x242 &  x257 &  x278 &  x281 &  x287 &  x299 &  x308 &  x326 &  x332 &  x359 &  x371 &  x374 &  x377 &  x383 &  x389 &  x395 &  x398 &  x413 &  x416 &  x422 &  x443 &  x470 &  x473 &  x500 &  x530 &  x551 &  x554 &  x557 &  x590 &  x626 &  x644 &  x662 &  x683 &  x689 &  x695 &  x704 &  x734 &  x740 &  x746 &  x764 &  x788 &  x815 &  x872 &  x890 &  x896 &  x926 &  x941 &  x944 &  x959 &  x974 &  x983 &  x992 &  x1010 &  x1049 &  x1052 &  x1064 &  x1079 &  x1112 &  x1118 & ~x111 & ~x150 & ~x189 & ~x228 & ~x306 & ~x345 & ~x372 & ~x384 & ~x411 & ~x450 & ~x489 & ~x528 & ~x567 & ~x570 & ~x843 & ~x906 & ~x945 & ~x984 & ~x1023 & ~x1101;
assign c7162 =  x86 &  x137 &  x188 &  x203 &  x209 &  x278 &  x323 &  x398 &  x403 &  x422 &  x434 &  x482 &  x509 &  x545 &  x578 &  x629 &  x689 &  x701 &  x716 &  x770 &  x785 &  x944 &  x959 &  x962 &  x1004 &  x1016 &  x1052 &  x1118 & ~x351 & ~x777 & ~x816 & ~x817 & ~x856 & ~x933 & ~x972 & ~x1018 & ~x1071 & ~x1096 & ~x1110;
assign c7164 =  x10 &  x26 &  x50 &  x68 &  x78 &  x125 &  x128 &  x131 &  x137 &  x140 &  x149 &  x179 &  x182 &  x194 &  x206 &  x209 &  x233 &  x239 &  x248 &  x260 &  x269 &  x272 &  x275 &  x284 &  x311 &  x314 &  x328 &  x335 &  x338 &  x359 &  x365 &  x398 &  x416 &  x428 &  x434 &  x446 &  x449 &  x500 &  x539 &  x557 &  x584 &  x587 &  x599 &  x626 &  x635 &  x650 &  x665 &  x677 &  x680 &  x719 &  x721 &  x722 &  x725 &  x767 &  x773 &  x809 &  x812 &  x815 &  x830 &  x833 &  x869 &  x896 &  x902 &  x920 &  x935 &  x962 &  x983 &  x989 &  x1019 &  x1043 &  x1046 &  x1061 &  x1064 &  x1079 &  x1100 &  x1121 &  x1130 & ~x45 & ~x84 & ~x85 & ~x162 & ~x355 & ~x394 & ~x471;
assign c7166 =  x35 &  x68 &  x71 &  x77 &  x86 &  x92 &  x101 &  x116 &  x131 &  x173 &  x188 &  x194 &  x200 &  x203 &  x221 &  x227 &  x248 &  x284 &  x407 &  x446 &  x482 &  x503 &  x560 &  x575 &  x599 &  x602 &  x626 &  x635 &  x647 &  x665 &  x782 &  x794 &  x842 &  x869 &  x890 &  x896 &  x941 &  x944 &  x977 &  x989 &  x992 &  x1009 &  x1043 &  x1048 &  x1052 &  x1088 &  x1094 &  x1118 &  x1121 & ~x39 & ~x117 & ~x189 & ~x228 & ~x267 & ~x306 & ~x345 & ~x384 & ~x423 & ~x882 & ~x921 & ~x933 & ~x960 & ~x972 & ~x993 & ~x999 & ~x1038 & ~x1071 & ~x1110;
assign c7168 =  x25 &  x422 &  x736 &  x752 &  x797 &  x890 &  x944 &  x959 &  x1052 & ~x21 & ~x39 & ~x177 & ~x216 & ~x372 & ~x411 & ~x615 & ~x882;
assign c7170 =  x4 &  x35 &  x43 &  x121 &  x131 &  x140 &  x149 &  x160 &  x209 &  x211 &  x218 &  x230 &  x250 &  x323 &  x326 &  x398 &  x406 &  x476 &  x523 &  x527 &  x548 &  x554 &  x559 &  x562 &  x601 &  x620 &  x640 &  x647 &  x650 &  x662 &  x679 &  x710 &  x737 &  x757 &  x764 &  x796 &  x815 &  x830 &  x863 &  x872 &  x874 &  x890 &  x941 &  x962 &  x970 &  x976 &  x991 &  x1030 &  x1043 &  x1069 &  x1106 &  x1130 & ~x993;
assign c7172 =  x5 &  x8 &  x17 &  x35 &  x86 &  x101 &  x128 &  x131 &  x140 &  x149 &  x170 &  x194 &  x209 &  x215 &  x254 &  x260 &  x266 &  x275 &  x278 &  x281 &  x287 &  x302 &  x335 &  x347 &  x350 &  x371 &  x374 &  x383 &  x395 &  x413 &  x428 &  x434 &  x440 &  x449 &  x455 &  x467 &  x470 &  x497 &  x500 &  x503 &  x512 &  x518 &  x557 &  x587 &  x590 &  x593 &  x599 &  x605 &  x617 &  x620 &  x623 &  x635 &  x641 &  x650 &  x662 &  x695 &  x701 &  x710 &  x713 &  x734 &  x737 &  x748 &  x755 &  x770 &  x787 &  x800 &  x802 &  x803 &  x809 &  x815 &  x818 &  x825 &  x826 &  x830 &  x842 &  x854 &  x857 &  x865 &  x872 &  x884 &  x887 &  x890 &  x893 &  x902 &  x904 &  x905 &  x917 &  x929 &  x935 &  x941 &  x959 &  x962 &  x965 &  x977 &  x1019 &  x1043 &  x1058 &  x1061 &  x1064 &  x1073 &  x1076 &  x1091 &  x1106 &  x1112 &  x1118 &  x1121 &  x1127 & ~x783 & ~x822 & ~x888;
assign c7174 =  x2 &  x17 &  x26 &  x35 &  x41 &  x83 &  x91 &  x98 &  x104 &  x110 &  x113 &  x116 &  x130 &  x131 &  x158 &  x161 &  x167 &  x188 &  x209 &  x218 &  x245 &  x260 &  x272 &  x281 &  x305 &  x308 &  x311 &  x335 &  x341 &  x365 &  x377 &  x424 &  x428 &  x440 &  x443 &  x470 &  x497 &  x524 &  x527 &  x545 &  x551 &  x569 &  x584 &  x596 &  x614 &  x617 &  x647 &  x656 &  x662 &  x674 &  x683 &  x695 &  x704 &  x731 &  x740 &  x749 &  x764 &  x770 &  x779 &  x782 &  x791 &  x797 &  x821 &  x851 &  x857 &  x866 &  x881 &  x890 &  x896 &  x920 &  x926 &  x929 &  x941 &  x959 &  x977 &  x980 &  x992 &  x1007 &  x1016 &  x1046 &  x1052 &  x1061 &  x1109 &  x1112 & ~x144 & ~x627 & ~x628 & ~x667 & ~x706 & ~x745 & ~x783 & ~x900;
assign c7176 =  x239 &  x282 &  x383 &  x709 &  x748 &  x902 & ~x345 & ~x358 & ~x450 & ~x706;
assign c7178 =  x35 &  x53 &  x119 &  x197 &  x224 &  x257 &  x260 &  x275 &  x287 &  x308 &  x320 &  x335 &  x383 &  x395 &  x398 &  x434 &  x439 &  x524 &  x554 &  x557 &  x569 &  x581 &  x586 &  x590 &  x602 &  x635 &  x638 &  x686 &  x710 &  x716 &  x755 &  x782 &  x788 &  x815 &  x821 &  x842 &  x890 &  x902 &  x929 &  x941 &  x959 &  x1004 &  x1010 &  x1034 &  x1064 &  x1094 &  x1100 &  x1112 &  x1118 & ~x393 & ~x432 & ~x501 & ~x540 & ~x642 & ~x648 & ~x681 & ~x687 & ~x720 & ~x798 & ~x837 & ~x940;
assign c7180 =  x11 &  x35 &  x47 &  x49 &  x56 &  x83 &  x86 &  x88 &  x101 &  x119 &  x125 &  x127 &  x143 &  x155 &  x172 &  x185 &  x211 &  x212 &  x218 &  x239 &  x272 &  x284 &  x299 &  x308 &  x326 &  x328 &  x341 &  x391 &  x406 &  x425 &  x428 &  x467 &  x479 &  x484 &  x500 &  x509 &  x524 &  x548 &  x562 &  x563 &  x569 &  x599 &  x601 &  x640 &  x641 &  x662 &  x674 &  x698 &  x701 &  x707 &  x710 &  x713 &  x728 &  x752 &  x758 &  x779 &  x788 &  x796 &  x802 &  x821 &  x824 &  x866 &  x869 &  x874 &  x884 &  x902 &  x929 &  x937 &  x991 &  x998 &  x1001 &  x1004 &  x1016 &  x1028 &  x1034 &  x1052 &  x1067 &  x1073 &  x1115 &  x1130 & ~x6 & ~x45 & ~x85 & ~x123 & ~x162;
assign c7182 =  x11 &  x35 &  x41 &  x86 &  x125 &  x179 &  x508 &  x548 &  x620 &  x640 &  x695 &  x725 &  x747 &  x748 &  x755 &  x757 &  x764 &  x770 &  x785 &  x786 &  x787 &  x796 &  x825 &  x865 &  x890 &  x905 &  x929 &  x941 &  x986 & ~x744 & ~x745 & ~x784;
assign c7184 =  x11 &  x26 &  x47 &  x125 &  x131 &  x148 &  x185 &  x187 &  x209 &  x260 &  x281 &  x308 &  x329 &  x338 &  x359 &  x455 &  x461 &  x479 &  x515 &  x620 &  x635 &  x650 &  x662 &  x698 &  x710 &  x743 &  x758 &  x761 &  x775 &  x776 &  x813 &  x814 &  x852 &  x853 &  x863 &  x890 &  x891 &  x892 &  x905 &  x931 &  x941 &  x944 &  x962 &  x970 &  x1009 &  x1016 &  x1028 &  x1043 &  x1048 &  x1087 &  x1130 & ~x228;
assign c7186 =  x2 &  x5 &  x38 &  x77 &  x92 &  x98 &  x101 &  x107 &  x146 &  x167 &  x173 &  x179 &  x209 &  x226 &  x260 &  x263 &  x275 &  x278 &  x299 &  x311 &  x325 &  x347 &  x353 &  x395 &  x407 &  x419 &  x442 &  x452 &  x485 &  x500 &  x560 &  x569 &  x602 &  x608 &  x662 &  x710 &  x716 &  x725 &  x731 &  x764 &  x776 &  x851 &  x866 &  x881 &  x890 &  x902 &  x920 &  x929 &  x935 &  x941 &  x965 &  x971 &  x992 &  x1034 &  x1037 &  x1043 &  x1061 &  x1073 &  x1109 & ~x306 & ~x345 & ~x384 & ~x423 & ~x435 & ~x436 & ~x450 & ~x474 & ~x489;
assign c7188 =  x26 &  x87 &  x88 &  x101 &  x116 &  x125 &  x131 &  x134 &  x166 &  x197 &  x200 &  x209 &  x230 &  x239 &  x257 &  x263 &  x275 &  x290 &  x293 &  x314 &  x326 &  x335 &  x365 &  x383 &  x407 &  x422 &  x464 &  x470 &  x527 &  x557 &  x569 &  x620 &  x635 &  x640 &  x644 &  x647 &  x686 &  x695 &  x725 &  x782 &  x797 &  x809 &  x827 &  x833 &  x842 &  x854 &  x884 &  x893 &  x935 &  x941 &  x992 &  x1001 &  x1007 &  x1016 &  x1019 &  x1034 &  x1052 &  x1058 &  x1073 &  x1094 &  x1118 &  x1121 & ~x123 & ~x163 & ~x201 & ~x202 & ~x240 & ~x408 & ~x486 & ~x525 & ~x564 & ~x666;
assign c7190 =  x2 &  x14 &  x20 &  x23 &  x26 &  x29 &  x41 &  x53 &  x56 &  x65 &  x80 &  x86 &  x104 &  x116 &  x125 &  x128 &  x134 &  x140 &  x146 &  x170 &  x179 &  x188 &  x191 &  x194 &  x197 &  x209 &  x221 &  x230 &  x233 &  x239 &  x242 &  x260 &  x272 &  x287 &  x314 &  x317 &  x335 &  x347 &  x359 &  x365 &  x383 &  x389 &  x395 &  x403 &  x407 &  x410 &  x416 &  x422 &  x442 &  x446 &  x467 &  x482 &  x491 &  x500 &  x524 &  x539 &  x542 &  x554 &  x569 &  x581 &  x584 &  x602 &  x626 &  x635 &  x641 &  x644 &  x650 &  x653 &  x662 &  x668 &  x674 &  x701 &  x704 &  x731 &  x740 &  x752 &  x755 &  x764 &  x785 &  x796 &  x821 &  x835 &  x857 &  x866 &  x872 &  x881 &  x890 &  x905 &  x911 &  x929 &  x944 &  x959 &  x965 &  x992 &  x1004 &  x1016 &  x1019 &  x1043 &  x1052 &  x1088 &  x1094 & ~x471 & ~x687 & ~x726 & ~x765 & ~x805 & ~x843 & ~x882 & ~x900 & ~x921 & ~x940 & ~x1065 & ~x1104;
assign c7192 =  x32 &  x35 &  x41 &  x59 &  x119 &  x125 &  x128 &  x131 &  x200 &  x209 &  x248 &  x263 &  x266 &  x323 &  x325 &  x335 &  x383 &  x392 &  x419 &  x430 &  x449 &  x452 &  x473 &  x479 &  x491 &  x503 &  x515 &  x545 &  x629 &  x656 &  x695 &  x707 &  x749 &  x763 &  x773 &  x776 &  x779 &  x782 &  x791 &  x802 &  x818 &  x821 &  x824 &  x833 &  x841 &  x890 &  x923 &  x959 &  x992 &  x1016 &  x1052 &  x1064 &  x1070 &  x1091 &  x1100 & ~x396 & ~x397 & ~x435 & ~x436 & ~x667 & ~x706 & ~x745 & ~x784;
assign c7194 =  x2 &  x5 &  x20 &  x35 &  x41 &  x47 &  x56 &  x86 &  x92 &  x116 &  x131 &  x143 &  x158 &  x194 &  x203 &  x209 &  x248 &  x257 &  x260 &  x275 &  x287 &  x296 &  x305 &  x308 &  x311 &  x320 &  x329 &  x335 &  x341 &  x368 &  x410 &  x416 &  x428 &  x431 &  x434 &  x440 &  x491 &  x512 &  x545 &  x572 &  x578 &  x584 &  x587 &  x593 &  x605 &  x626 &  x633 &  x634 &  x647 &  x665 &  x672 &  x680 &  x686 &  x703 &  x719 &  x725 &  x781 &  x800 &  x815 &  x820 &  x842 &  x860 &  x872 &  x890 &  x902 &  x911 &  x938 &  x941 &  x944 &  x947 &  x983 &  x1010 &  x1013 &  x1025 &  x1046 &  x1048 &  x1052 &  x1058 &  x1064 &  x1070 &  x1106 &  x1118 &  x1121 & ~x510 & ~x627 & ~x684 & ~x723 & ~x762 & ~x1018 & ~x1057 & ~x1096;
assign c7196 =  x10 &  x17 &  x49 &  x82 &  x88 &  x157 &  x160 &  x221 &  x274 &  x359 &  x406 &  x424 &  x467 &  x485 &  x500 &  x523 &  x562 &  x590 &  x602 &  x611 &  x640 &  x689 &  x695 &  x737 &  x743 &  x755 &  x796 &  x797 &  x809 &  x881 &  x935 &  x1010 &  x1052 & ~x102 & ~x219 & ~x225 & ~x258 & ~x408;
assign c7198 =  x2 &  x11 &  x65 &  x71 &  x101 &  x107 &  x128 &  x131 &  x149 &  x179 &  x206 &  x212 &  x221 &  x233 &  x257 &  x299 &  x320 &  x341 &  x360 &  x400 &  x401 &  x416 &  x440 &  x455 &  x458 &  x461 &  x464 &  x468 &  x485 &  x488 &  x503 &  x508 &  x554 &  x575 &  x590 &  x596 &  x599 &  x605 &  x629 &  x635 &  x640 &  x641 &  x647 &  x662 &  x665 &  x695 &  x710 &  x718 &  x725 &  x734 &  x764 &  x794 &  x806 &  x812 &  x848 &  x854 &  x890 &  x905 &  x956 &  x962 &  x965 &  x971 &  x980 &  x995 &  x1019 &  x1043 &  x1052 &  x1061 &  x1070 &  x1091 &  x1100 &  x1124 & ~x357 & ~x387 & ~x396 & ~x783 & ~x784 & ~x822;
assign c7200 =  x23 &  x59 &  x65 &  x70 &  x116 &  x131 &  x134 &  x143 &  x149 &  x152 &  x253 &  x338 &  x341 &  x344 &  x383 &  x410 &  x469 &  x508 &  x512 &  x521 &  x533 &  x581 &  x587 &  x620 &  x638 &  x698 &  x707 &  x719 &  x755 &  x791 &  x809 &  x887 &  x893 &  x896 &  x917 &  x959 &  x1010 &  x1046 &  x1058 &  x1073 &  x1106 &  x1118 &  x1127 & ~x357 & ~x397 & ~x414 & ~x435 & ~x436 & ~x474 & ~x706 & ~x745;
assign c7202 =  x17 &  x29 &  x56 &  x59 &  x74 &  x91 &  x169 &  x212 &  x221 &  x254 &  x263 &  x302 &  x313 &  x338 &  x389 &  x470 &  x473 &  x497 &  x524 &  x541 &  x580 &  x584 &  x623 &  x632 &  x658 &  x692 &  x773 &  x893 &  x929 &  x1016 &  x1031 &  x1043 &  x1046 &  x1091 &  x1100 & ~x219 & ~x369 & ~x667 & ~x783 & ~x1062 & ~x1101;
assign c7204 =  x41 &  x47 &  x77 &  x112 &  x119 &  x122 &  x131 &  x143 &  x172 &  x209 &  x211 &  x250 &  x260 &  x275 &  x278 &  x298 &  x328 &  x337 &  x340 &  x373 &  x379 &  x385 &  x406 &  x416 &  x421 &  x434 &  x457 &  x499 &  x520 &  x523 &  x559 &  x562 &  x569 &  x601 &  x617 &  x650 &  x695 &  x710 &  x758 &  x859 &  x872 &  x884 &  x892 &  x898 &  x905 &  x926 &  x931 &  x941 &  x970 &  x1037 &  x1046 &  x1076 &  x1079 &  x1082 &  x1106 &  x1126;
assign c7206 =  x20 &  x41 &  x77 &  x86 &  x104 &  x131 &  x140 &  x155 &  x167 &  x185 &  x188 &  x191 &  x218 &  x224 &  x242 &  x275 &  x308 &  x332 &  x359 &  x361 &  x380 &  x395 &  x399 &  x413 &  x416 &  x425 &  x428 &  x438 &  x439 &  x443 &  x503 &  x515 &  x517 &  x524 &  x545 &  x554 &  x572 &  x581 &  x586 &  x590 &  x602 &  x605 &  x650 &  x662 &  x674 &  x686 &  x704 &  x716 &  x725 &  x737 &  x758 &  x785 &  x839 &  x872 &  x878 &  x890 &  x935 &  x941 &  x944 &  x965 &  x992 &  x1010 &  x1022 &  x1043 &  x1046 &  x1055 &  x1073 &  x1100 &  x1103 &  x1106 &  x1118 & ~x435 & ~x450 & ~x474 & ~x489 & ~x528 & ~x648 & ~x687 & ~x784 & ~x823;
assign c7208 =  x235 &  x335 &  x613 &  x691 & ~x201 & ~x232 & ~x271 & ~x550 & ~x589;
assign c7210 =  x49 &  x88 &  x121 &  x155 &  x170 &  x191 &  x274 &  x455 &  x545 &  x601 &  x656 &  x668 &  x737 &  x767 &  x782 &  x959 &  x1031 & ~x6 & ~x46 & ~x84 & ~x85 & ~x124 & ~x135 & ~x201 & ~x202 & ~x219 & ~x258 & ~x822;
assign c7212 =  x5 &  x26 &  x83 &  x143 &  x188 &  x221 &  x224 &  x243 &  x257 &  x272 &  x278 &  x290 &  x293 &  x419 &  x430 &  x440 &  x467 &  x476 &  x479 &  x533 &  x539 &  x554 &  x581 &  x584 &  x669 &  x670 &  x704 &  x709 &  x713 &  x728 &  x748 &  x755 &  x787 &  x809 &  x815 &  x833 &  x857 &  x896 &  x905 &  x971 &  x1001 &  x1010 &  x1016 &  x1043 &  x1052 &  x1073 &  x1082 &  x1118 & ~x667 & ~x706 & ~x745;
assign c7214 =  x244 &  x359 &  x390 &  x428 &  x429 &  x586 &  x593 &  x608 &  x671 &  x695 &  x749 &  x841 &  x929 &  x1001 &  x1103 & ~x318 & ~x357 & ~x358 & ~x397 & ~x435 & ~x666 & ~x667 & ~x706 & ~x745 & ~x784;
assign c7216 =  x25 &  x35 &  x47 &  x52 &  x53 &  x64 &  x86 &  x91 &  x103 &  x113 &  x130 &  x164 &  x169 &  x212 &  x224 &  x285 &  x286 &  x296 &  x389 &  x413 &  x440 &  x503 &  x551 &  x563 &  x601 &  x602 &  x629 &  x638 &  x640 &  x644 &  x677 &  x728 &  x755 &  x779 &  x842 &  x881 &  x890 &  x893 &  x938 &  x971 &  x1013 &  x1043 &  x1061 &  x1097 &  x1112 & ~x666 & ~x705 & ~x706 & ~x745 & ~x783 & ~x822;
assign c7218 =  x26 &  x56 &  x104 &  x116 &  x125 &  x128 &  x131 &  x209 &  x239 &  x245 &  x278 &  x341 &  x350 &  x458 &  x477 &  x480 &  x500 &  x554 &  x557 &  x581 &  x617 &  x644 &  x647 &  x701 &  x737 &  x874 &  x878 &  x890 &  x926 &  x944 &  x992 &  x998 &  x1046 &  x1052 &  x1058 &  x1112 & ~x592 & ~x630 & ~x940;
assign c7220 =  x26 &  x29 &  x53 &  x64 &  x65 &  x77 &  x103 &  x128 &  x181 &  x188 &  x197 &  x242 &  x257 &  x259 &  x323 &  x329 &  x340 &  x356 &  x373 &  x421 &  x460 &  x484 &  x487 &  x497 &  x499 &  x520 &  x523 &  x559 &  x716 &  x794 &  x820 &  x914 &  x929 &  x970 &  x976 &  x1004 &  x1009 &  x1015 &  x1052 &  x1058 &  x1094 &  x1112 & ~x1050;
assign c7222 =  x13 &  x17 &  x41 &  x131 &  x194 &  x209 &  x212 &  x281 &  x287 &  x314 &  x383 &  x428 &  x470 &  x491 &  x497 &  x509 &  x535 &  x545 &  x548 &  x569 &  x574 &  x575 &  x593 &  x602 &  x605 &  x692 &  x719 &  x815 &  x869 &  x884 &  x896 &  x917 &  x920 &  x1043 &  x1046 &  x1052 &  x1100 &  x1112 & ~x66 & ~x177 & ~x216 & ~x546 & ~x549 & ~x585 & ~x819;
assign c7224 =  x26 &  x29 &  x38 &  x86 &  x101 &  x140 &  x152 &  x155 &  x158 &  x173 &  x203 &  x220 &  x230 &  x251 &  x259 &  x263 &  x298 &  x304 &  x308 &  x407 &  x409 &  x415 &  x421 &  x434 &  x448 &  x457 &  x460 &  x476 &  x487 &  x497 &  x503 &  x520 &  x548 &  x559 &  x602 &  x620 &  x626 &  x677 &  x686 &  x710 &  x711 &  x722 &  x731 &  x751 &  x791 &  x794 &  x800 &  x812 &  x820 &  x860 &  x869 &  x932 &  x1007 &  x1015 &  x1022 &  x1031 &  x1034 &  x1054 &  x1064 &  x1073 & ~x273 & ~x468 & ~x507 & ~x999;
assign c7226 =  x161 &  x200 &  x209 &  x215 &  x244 &  x286 &  x469 &  x518 &  x580 &  x617 &  x658 &  x697 &  x707 &  x755 &  x770 &  x854 &  x872 &  x956 &  x1118 & ~x357 & ~x486 & ~x628 & ~x667 & ~x705 & ~x706 & ~x745 & ~x784 & ~x822;
assign c7228 =  x143 &  x152 &  x197 &  x203 &  x251 &  x265 &  x314 &  x413 &  x445 &  x484 &  x601 &  x661 &  x717 &  x756 &  x797 &  x833 &  x834 &  x873 &  x899 &  x951 &  x956 &  x1022;
assign c7230 =  x8 &  x26 &  x32 &  x74 &  x83 &  x116 &  x161 &  x164 &  x209 &  x230 &  x251 &  x263 &  x287 &  x290 &  x317 &  x326 &  x335 &  x344 &  x356 &  x359 &  x365 &  x380 &  x409 &  x515 &  x524 &  x527 &  x581 &  x632 &  x641 &  x644 &  x650 &  x674 &  x686 &  x698 &  x707 &  x725 &  x737 &  x755 &  x773 &  x797 &  x818 &  x848 &  x859 &  x890 &  x898 &  x914 &  x932 &  x937 &  x977 &  x1025 &  x1046 &  x1109 & ~x765 & ~x843 & ~x888 & ~x928 & ~x967 & ~x1006 & ~x1045 & ~x1057 & ~x1083 & ~x1084 & ~x1122;
assign c7232 =  x11 &  x26 &  x32 &  x35 &  x53 &  x59 &  x65 &  x83 &  x107 &  x119 &  x125 &  x128 &  x131 &  x149 &  x188 &  x203 &  x205 &  x209 &  x221 &  x239 &  x254 &  x278 &  x313 &  x341 &  x344 &  x350 &  x359 &  x383 &  x398 &  x422 &  x425 &  x428 &  x469 &  x503 &  x530 &  x541 &  x554 &  x560 &  x580 &  x581 &  x587 &  x605 &  x617 &  x619 &  x620 &  x632 &  x635 &  x638 &  x644 &  x653 &  x657 &  x658 &  x695 &  x696 &  x697 &  x701 &  x719 &  x731 &  x734 &  x735 &  x736 &  x752 &  x775 &  x827 &  x833 &  x841 &  x851 &  x863 &  x875 &  x892 &  x896 &  x905 &  x929 &  x931 &  x935 &  x941 &  x958 &  x986 &  x1019 &  x1046 &  x1064 &  x1070 &  x1073 &  x1121 &  x1124 & ~x369 & ~x408 & ~x447 & ~x486 & ~x822;
assign c7234 =  x41 &  x86 &  x93 &  x119 &  x125 &  x166 &  x205 &  x211 &  x239 &  x249 &  x257 &  x263 &  x265 &  x272 &  x284 &  x287 &  x323 &  x367 &  x407 &  x473 &  x497 &  x518 &  x584 &  x611 &  x626 &  x640 &  x650 &  x679 &  x680 &  x686 &  x791 &  x818 &  x857 &  x863 &  x875 &  x902 &  x1076 & ~x666 & ~x933;
assign c7236 =  x11 &  x41 &  x56 &  x65 &  x77 &  x86 &  x89 &  x104 &  x113 &  x119 &  x131 &  x172 &  x185 &  x203 &  x209 &  x211 &  x230 &  x245 &  x254 &  x260 &  x263 &  x278 &  x281 &  x284 &  x302 &  x311 &  x317 &  x320 &  x326 &  x335 &  x371 &  x377 &  x382 &  x383 &  x403 &  x413 &  x416 &  x419 &  x440 &  x442 &  x449 &  x455 &  x480 &  x481 &  x491 &  x497 &  x500 &  x518 &  x519 &  x530 &  x559 &  x566 &  x584 &  x590 &  x597 &  x605 &  x620 &  x623 &  x626 &  x638 &  x662 &  x689 &  x695 &  x752 &  x755 &  x779 &  x785 &  x796 &  x797 &  x812 &  x821 &  x824 &  x857 &  x872 &  x908 &  x911 &  x962 &  x971 &  x976 &  x992 &  x1015 &  x1034 &  x1052 &  x1054 &  x1061 &  x1067 &  x1069 &  x1100 &  x1108 &  x1112 &  x1118 &  x1121;
assign c7238 =  x11 &  x14 &  x17 &  x20 &  x26 &  x29 &  x35 &  x47 &  x53 &  x56 &  x65 &  x86 &  x101 &  x107 &  x125 &  x128 &  x131 &  x146 &  x155 &  x170 &  x173 &  x179 &  x185 &  x188 &  x194 &  x197 &  x200 &  x209 &  x212 &  x221 &  x224 &  x230 &  x239 &  x242 &  x248 &  x260 &  x278 &  x284 &  x293 &  x299 &  x314 &  x317 &  x335 &  x398 &  x407 &  x413 &  x415 &  x416 &  x419 &  x422 &  x431 &  x440 &  x443 &  x467 &  x479 &  x500 &  x506 &  x509 &  x554 &  x559 &  x569 &  x572 &  x605 &  x611 &  x620 &  x644 &  x647 &  x659 &  x662 &  x680 &  x686 &  x692 &  x695 &  x698 &  x707 &  x710 &  x716 &  x725 &  x752 &  x758 &  x776 &  x779 &  x781 &  x794 &  x797 &  x803 &  x814 &  x839 &  x842 &  x857 &  x872 &  x881 &  x890 &  x892 &  x914 &  x917 &  x931 &  x937 &  x952 &  x953 &  x970 &  x974 &  x976 &  x986 &  x991 &  x1007 &  x1015 &  x1019 &  x1030 &  x1034 &  x1043 &  x1049 &  x1052 &  x1054 &  x1055 &  x1067 &  x1069 &  x1073 &  x1094 &  x1106 &  x1118 & ~x117 & ~x195 & ~x273 & ~x882 & ~x921 & ~x960 & ~x1011;
assign c7240 =  x41 &  x101 &  x155 &  x259 &  x265 &  x296 &  x298 &  x338 &  x340 &  x343 &  x379 &  x383 &  x421 &  x457 &  x485 &  x500 &  x523 &  x559 &  x601 &  x611 &  x640 &  x650 &  x695 &  x734 &  x740 &  x874 &  x890 &  x897 &  x908 &  x941 &  x975 &  x991 &  x1014 &  x1029 &  x1030 &  x1043 &  x1052 &  x1053;
assign c7242 =  x65 &  x116 &  x140 &  x142 &  x148 &  x187 &  x209 &  x226 &  x253 &  x281 &  x286 &  x323 &  x365 &  x383 &  x416 &  x442 &  x464 &  x527 &  x551 &  x572 &  x601 &  x620 &  x640 &  x679 &  x686 &  x717 &  x718 &  x755 &  x756 &  x795 &  x796 &  x821 &  x872 &  x874 &  x890 &  x929 &  x944 &  x959 &  x983 &  x1064 &  x1070;
assign c7244 =  x47 &  x53 &  x56 &  x68 &  x164 &  x209 &  x224 &  x263 &  x281 &  x428 &  x434 &  x446 &  x479 &  x500 &  x533 &  x559 &  x569 &  x581 &  x602 &  x638 &  x680 &  x689 &  x695 &  x707 &  x725 &  x746 &  x781 &  x842 &  x854 &  x857 &  x859 &  x872 &  x887 &  x890 &  x941 &  x970 &  x1046 &  x1064 &  x1070 &  x1087 &  x1103 &  x1118 & ~x765 & ~x798 & ~x837 & ~x915 & ~x960 & ~x994 & ~x1033 & ~x1038 & ~x1072 & ~x1110 & ~x1111;
assign c7246 =  x205 &  x244 &  x260 &  x540 &  x735 &  x736 &  x1010 & ~x318 & ~x447 & ~x667 & ~x706;
assign c7248 =  x11 &  x35 &  x38 &  x41 &  x53 &  x59 &  x77 &  x101 &  x107 &  x131 &  x146 &  x149 &  x170 &  x176 &  x194 &  x200 &  x209 &  x221 &  x233 &  x239 &  x260 &  x278 &  x287 &  x292 &  x314 &  x320 &  x323 &  x335 &  x350 &  x359 &  x364 &  x370 &  x383 &  x389 &  x403 &  x407 &  x409 &  x410 &  x413 &  x422 &  x434 &  x439 &  x467 &  x477 &  x482 &  x494 &  x500 &  x516 &  x530 &  x545 &  x556 &  x569 &  x572 &  x575 &  x590 &  x617 &  x638 &  x644 &  x662 &  x686 &  x692 &  x695 &  x701 &  x707 &  x710 &  x725 &  x737 &  x764 &  x788 &  x794 &  x797 &  x812 &  x818 &  x833 &  x842 &  x854 &  x872 &  x884 &  x890 &  x896 &  x905 &  x911 &  x917 &  x929 &  x935 &  x941 &  x953 &  x956 &  x959 &  x965 &  x983 &  x1004 &  x1013 &  x1019 &  x1034 &  x1043 &  x1049 &  x1052 &  x1061 &  x1064 &  x1118 &  x1121 & ~x513 & ~x528 & ~x567 & ~x900 & ~x1026;
assign c7250 =  x91 &  x131 &  x320 &  x352 &  x527 &  x562 &  x581 &  x791 &  x857 &  x1043 & ~x258 & ~x298 & ~x337 & ~x511 & ~x741;
assign c7252 =  x19 &  x41 &  x44 &  x58 &  x65 &  x74 &  x91 &  x97 &  x101 &  x104 &  x107 &  x122 &  x130 &  x131 &  x169 &  x173 &  x185 &  x194 &  x208 &  x209 &  x212 &  x224 &  x230 &  x233 &  x236 &  x251 &  x260 &  x281 &  x284 &  x287 &  x293 &  x314 &  x325 &  x335 &  x350 &  x363 &  x364 &  x371 &  x403 &  x416 &  x428 &  x437 &  x467 &  x473 &  x518 &  x521 &  x530 &  x542 &  x545 &  x557 &  x569 &  x572 &  x602 &  x617 &  x638 &  x647 &  x695 &  x701 &  x707 &  x710 &  x716 &  x725 &  x737 &  x776 &  x782 &  x785 &  x791 &  x815 &  x824 &  x833 &  x842 &  x872 &  x890 &  x896 &  x926 &  x929 &  x935 &  x965 &  x977 &  x1031 &  x1043 &  x1052 &  x1061 &  x1067 &  x1073 &  x1082 &  x1094 &  x1100 &  x1106 & ~x0 & ~x39 & ~x117 & ~x156 & ~x450 & ~x861 & ~x940;
assign c7254 =  x20 &  x26 &  x41 &  x74 &  x83 &  x86 &  x101 &  x107 &  x125 &  x146 &  x149 &  x188 &  x191 &  x200 &  x209 &  x212 &  x224 &  x260 &  x281 &  x293 &  x302 &  x308 &  x335 &  x341 &  x413 &  x422 &  x428 &  x491 &  x503 &  x548 &  x557 &  x569 &  x572 &  x596 &  x605 &  x623 &  x626 &  x662 &  x686 &  x695 &  x698 &  x704 &  x707 &  x716 &  x725 &  x737 &  x755 &  x800 &  x818 &  x821 &  x833 &  x890 &  x905 &  x917 &  x935 &  x941 &  x962 &  x965 &  x1010 &  x1034 &  x1060 &  x1079 &  x1097 &  x1099 &  x1106 &  x1112 &  x1115 & ~x351 & ~x579 & ~x921 & ~x945 & ~x972 & ~x984 & ~x985 & ~x999 & ~x1023 & ~x1062 & ~x1101;
assign c7256 =  x20 &  x92 &  x125 &  x134 &  x215 &  x278 &  x326 &  x344 &  x359 &  x368 &  x401 &  x506 &  x512 &  x584 &  x601 &  x671 &  x677 &  x695 &  x716 &  x737 &  x776 &  x797 &  x842 &  x878 &  x938 &  x1007 &  x1037 &  x1046 & ~x96 & ~x99 & ~x439 & ~x492 & ~x624;
assign c7258 =  x29 &  x32 &  x53 &  x65 &  x68 &  x104 &  x107 &  x128 &  x170 &  x188 &  x197 &  x224 &  x260 &  x275 &  x304 &  x305 &  x308 &  x338 &  x343 &  x350 &  x359 &  x383 &  x388 &  x409 &  x427 &  x434 &  x467 &  x481 &  x509 &  x524 &  x548 &  x563 &  x572 &  x581 &  x594 &  x635 &  x641 &  x650 &  x662 &  x686 &  x698 &  x710 &  x725 &  x734 &  x752 &  x781 &  x782 &  x785 &  x821 &  x859 &  x872 &  x875 &  x896 &  x911 &  x941 &  x959 &  x1004 &  x1015 &  x1016 &  x1019 &  x1025 &  x1034 &  x1043 &  x1052 &  x1064 & ~x390 & ~x630 & ~x960;
assign c7260 =  x155 &  x167 &  x203 &  x209 &  x233 &  x239 &  x242 &  x317 &  x320 &  x323 &  x350 &  x442 &  x446 &  x473 &  x512 &  x554 &  x680 &  x692 &  x758 &  x764 &  x770 &  x791 &  x809 &  x821 &  x854 &  x866 &  x890 &  x902 &  x917 &  x941 &  x944 &  x953 &  x959 &  x965 &  x1013 &  x1118 & ~x0 & ~x39 & ~x78 & ~x117 & ~x177 & ~x189 & ~x210 & ~x228 & ~x249 & ~x267 & ~x306 & ~x423 & ~x513 & ~x528 & ~x798 & ~x837 & ~x921;
assign c7262 =  x26 &  x32 &  x35 &  x41 &  x44 &  x59 &  x86 &  x98 &  x101 &  x107 &  x119 &  x125 &  x128 &  x131 &  x149 &  x155 &  x170 &  x179 &  x182 &  x191 &  x194 &  x206 &  x209 &  x212 &  x218 &  x224 &  x233 &  x245 &  x248 &  x251 &  x254 &  x260 &  x275 &  x281 &  x284 &  x287 &  x293 &  x296 &  x302 &  x308 &  x320 &  x326 &  x335 &  x350 &  x353 &  x356 &  x377 &  x380 &  x383 &  x395 &  x407 &  x413 &  x416 &  x434 &  x440 &  x446 &  x449 &  x452 &  x455 &  x458 &  x467 &  x470 &  x476 &  x482 &  x491 &  x500 &  x515 &  x524 &  x530 &  x539 &  x548 &  x557 &  x569 &  x572 &  x575 &  x581 &  x590 &  x593 &  x602 &  x605 &  x620 &  x626 &  x635 &  x638 &  x641 &  x644 &  x647 &  x650 &  x662 &  x680 &  x686 &  x689 &  x692 &  x695 &  x701 &  x710 &  x725 &  x743 &  x746 &  x749 &  x752 &  x755 &  x758 &  x781 &  x782 &  x785 &  x788 &  x797 &  x800 &  x806 &  x815 &  x818 &  x820 &  x821 &  x833 &  x836 &  x851 &  x857 &  x858 &  x872 &  x884 &  x890 &  x896 &  x897 &  x902 &  x908 &  x911 &  x929 &  x937 &  x938 &  x941 &  x944 &  x962 &  x975 &  x983 &  x989 &  x991 &  x1010 &  x1014 &  x1015 &  x1016 &  x1019 &  x1030 &  x1043 &  x1046 &  x1049 &  x1052 &  x1053 &  x1054 &  x1055 &  x1061 &  x1069 &  x1070 &  x1073 &  x1092 &  x1100 &  x1106 &  x1112 &  x1115 &  x1118 &  x1121 &  x1124 &  x1127 & ~x846 & ~x882 & ~x921 & ~x960 & ~x999 & ~x1038 & ~x1056 & ~x1057 & ~x1083 & ~x1096 & ~x1122;
assign c7264 =  x10 &  x88 &  x121 &  x127 &  x209 &  x245 &  x284 &  x289 &  x293 &  x385 &  x457 &  x496 &  x613 &  x626 &  x652 &  x679 &  x695 &  x719 &  x721 &  x950 &  x1019 &  x1100 & ~x219 & ~x369 & ~x408;
assign c7266 =  x79 &  x86 &  x87 &  x88 &  x140 &  x152 &  x209 &  x533 &  x608 &  x809 &  x830 &  x875 &  x926 &  x941 &  x995 &  x1079 &  x1130 & ~x141 & ~x220 & ~x258 & ~x433 & ~x472 & ~x511 & ~x550;
assign c7268 =  x29 &  x35 &  x41 &  x50 &  x56 &  x80 &  x104 &  x134 &  x146 &  x179 &  x188 &  x191 &  x209 &  x224 &  x239 &  x245 &  x317 &  x395 &  x398 &  x422 &  x434 &  x443 &  x467 &  x497 &  x569 &  x602 &  x695 &  x707 &  x770 &  x781 &  x791 &  x872 &  x890 &  x892 &  x905 &  x929 &  x931 &  x941 &  x944 &  x956 &  x970 &  x992 &  x1008 &  x1009 &  x1010 &  x1013 &  x1047 &  x1048 &  x1049 &  x1070 &  x1073 &  x1087 &  x1100 &  x1106 &  x1126 & ~x432 & ~x882 & ~x883 & ~x921 & ~x960 & ~x999 & ~x1057 & ~x1077;
assign c7270 =  x20 &  x53 &  x56 &  x86 &  x146 &  x164 &  x170 &  x197 &  x209 &  x221 &  x244 &  x248 &  x257 &  x269 &  x323 &  x332 &  x365 &  x395 &  x406 &  x413 &  x416 &  x434 &  x461 &  x464 &  x470 &  x545 &  x551 &  x554 &  x587 &  x601 &  x626 &  x640 &  x670 &  x679 &  x692 &  x709 &  x718 &  x724 &  x752 &  x781 &  x796 &  x802 &  x809 &  x812 &  x824 &  x835 &  x841 &  x860 &  x872 &  x890 &  x902 &  x926 &  x929 &  x956 &  x968 &  x980 &  x983 &  x1031 &  x1049 &  x1064 &  x1073 &  x1085 &  x1094 &  x1097 &  x1103 &  x1121 & ~x357 & ~x745 & ~x822;
assign c7272 =  x104 &  x220 &  x259 &  x265 &  x520 &  x562 &  x615 &  x616 &  x644 &  x662 &  x694 &  x809 &  x827 &  x887 &  x935 &  x952 &  x991 &  x1043 &  x1052 &  x1069 &  x1118;
assign c7274 =  x8 &  x14 &  x29 &  x32 &  x41 &  x53 &  x71 &  x80 &  x86 &  x92 &  x107 &  x116 &  x119 &  x122 &  x140 &  x170 &  x173 &  x185 &  x191 &  x194 &  x197 &  x212 &  x244 &  x251 &  x263 &  x266 &  x272 &  x287 &  x290 &  x293 &  x299 &  x305 &  x329 &  x347 &  x352 &  x391 &  x392 &  x395 &  x410 &  x425 &  x430 &  x443 &  x469 &  x470 &  x482 &  x485 &  x488 &  x500 &  x542 &  x547 &  x551 &  x554 &  x569 &  x581 &  x584 &  x605 &  x614 &  x640 &  x641 &  x644 &  x656 &  x665 &  x670 &  x679 &  x686 &  x695 &  x698 &  x707 &  x719 &  x734 &  x755 &  x794 &  x796 &  x809 &  x812 &  x821 &  x851 &  x884 &  x890 &  x917 &  x947 &  x953 &  x956 &  x971 &  x974 &  x983 &  x986 &  x1001 &  x1010 &  x1034 &  x1037 &  x1046 &  x1052 &  x1055 &  x1061 &  x1064 &  x1070 &  x1078 &  x1079 &  x1085 &  x1088 &  x1100 &  x1127 & ~x375 & ~x414 & ~x564 & ~x627 & ~x628 & ~x667 & ~x705 & ~x706;
assign c7276 =  x56 &  x68 &  x71 &  x95 &  x194 &  x209 &  x226 &  x259 &  x265 &  x281 &  x298 &  x304 &  x314 &  x326 &  x337 &  x343 &  x350 &  x383 &  x409 &  x415 &  x421 &  x422 &  x470 &  x487 &  x527 &  x559 &  x569 &  x637 &  x650 &  x746 &  x761 &  x815 &  x830 &  x898 &  x941 &  x976 &  x1043 &  x1054 & ~x273 & ~x618 & ~x657 & ~x765 & ~x960;
assign c7278 =  x23 &  x29 &  x35 &  x56 &  x86 &  x149 &  x155 &  x173 &  x185 &  x191 &  x194 &  x209 &  x221 &  x239 &  x260 &  x275 &  x308 &  x323 &  x326 &  x341 &  x347 &  x350 &  x371 &  x377 &  x383 &  x398 &  x403 &  x442 &  x446 &  x470 &  x509 &  x520 &  x530 &  x551 &  x572 &  x584 &  x586 &  x590 &  x596 &  x617 &  x620 &  x623 &  x626 &  x638 &  x641 &  x644 &  x662 &  x664 &  x764 &  x779 &  x781 &  x782 &  x788 &  x791 &  x796 &  x809 &  x821 &  x830 &  x833 &  x842 &  x854 &  x872 &  x887 &  x890 &  x892 &  x898 &  x917 &  x920 &  x926 &  x929 &  x931 &  x937 &  x958 &  x959 &  x970 &  x971 &  x974 &  x992 &  x1004 &  x1009 &  x1016 &  x1019 &  x1043 &  x1046 &  x1049 &  x1054 &  x1067 &  x1112 &  x1124 &  x1130 & ~x237 & ~x393 & ~x687 & ~x940 & ~x1050;
assign c7280 =  x17 &  x127 &  x260 &  x281 &  x461 &  x470 &  x482 &  x483 &  x522 &  x523 &  x524 &  x561 &  x572 &  x629 &  x640 &  x686 &  x713 &  x796 &  x806 &  x824 &  x1037 & ~x219 & ~x258 & ~x298 & ~x744;
assign c7282 =  x13 &  x17 &  x56 &  x80 &  x104 &  x131 &  x146 &  x152 &  x167 &  x188 &  x194 &  x209 &  x235 &  x308 &  x329 &  x341 &  x377 &  x398 &  x416 &  x422 &  x428 &  x437 &  x467 &  x509 &  x524 &  x548 &  x557 &  x560 &  x620 &  x632 &  x638 &  x662 &  x686 &  x689 &  x695 &  x725 &  x770 &  x815 &  x827 &  x872 &  x890 &  x935 &  x944 &  x986 &  x1004 &  x1019 &  x1028 &  x1052 &  x1100 & ~x193 & ~x258 & ~x447 & ~x510 & ~x549 & ~x550 & ~x589 & ~x627;
assign c7284 =  x41 &  x89 &  x101 &  x131 &  x140 &  x146 &  x221 &  x257 &  x287 &  x487 &  x497 &  x572 &  x594 &  x605 &  x629 &  x633 &  x695 &  x710 &  x725 &  x794 &  x815 &  x842 &  x869 &  x890 &  x959 &  x976 &  x1052 &  x1073 & ~x798 & ~x799 & ~x838 & ~x954 & ~x993;
assign c7286 =  x8 &  x13 &  x29 &  x146 &  x160 &  x209 &  x230 &  x281 &  x335 &  x482 &  x535 &  x635 &  x716 &  x752 &  x815 &  x833 &  x1072 & ~x123 & ~x124 & ~x163;
assign c7288 =  x41 &  x49 &  x56 &  x101 &  x104 &  x113 &  x156 &  x188 &  x233 &  x248 &  x263 &  x278 &  x287 &  x302 &  x320 &  x383 &  x407 &  x449 &  x496 &  x535 &  x644 &  x734 &  x746 &  x752 &  x779 &  x857 &  x872 &  x875 &  x878 &  x902 &  x929 &  x1019 &  x1052 &  x1055 & ~x123 & ~x124 & ~x163 & ~x216 & ~x219 & ~x511;
assign c7290 =  x10 &  x14 &  x47 &  x88 &  x92 &  x95 &  x98 &  x119 &  x128 &  x131 &  x134 &  x143 &  x161 &  x173 &  x185 &  x191 &  x206 &  x209 &  x230 &  x260 &  x275 &  x293 &  x326 &  x335 &  x341 &  x353 &  x362 &  x368 &  x404 &  x410 &  x422 &  x428 &  x458 &  x461 &  x494 &  x500 &  x506 &  x527 &  x551 &  x569 &  x572 &  x611 &  x614 &  x626 &  x629 &  x662 &  x668 &  x691 &  x695 &  x701 &  x725 &  x749 &  x764 &  x773 &  x779 &  x788 &  x794 &  x797 &  x800 &  x803 &  x812 &  x836 &  x869 &  x890 &  x896 &  x902 &  x920 &  x932 &  x992 &  x1001 &  x1022 &  x1034 &  x1049 &  x1070 &  x1082 &  x1109 &  x1124 & ~x124 & ~x177 & ~x219 & ~x433 & ~x471 & ~x472;
assign c7292 =  x20 &  x23 &  x26 &  x41 &  x53 &  x59 &  x65 &  x74 &  x83 &  x86 &  x92 &  x95 &  x101 &  x116 &  x131 &  x149 &  x164 &  x179 &  x188 &  x194 &  x197 &  x203 &  x206 &  x209 &  x221 &  x224 &  x230 &  x233 &  x236 &  x239 &  x242 &  x245 &  x248 &  x254 &  x260 &  x263 &  x272 &  x278 &  x281 &  x284 &  x302 &  x317 &  x323 &  x335 &  x338 &  x341 &  x344 &  x350 &  x353 &  x359 &  x362 &  x365 &  x368 &  x374 &  x377 &  x380 &  x383 &  x389 &  x395 &  x398 &  x401 &  x413 &  x416 &  x419 &  x422 &  x428 &  x434 &  x440 &  x446 &  x449 &  x452 &  x488 &  x509 &  x524 &  x527 &  x530 &  x545 &  x548 &  x557 &  x560 &  x569 &  x572 &  x575 &  x587 &  x599 &  x602 &  x611 &  x617 &  x620 &  x629 &  x635 &  x638 &  x644 &  x650 &  x653 &  x686 &  x689 &  x695 &  x701 &  x710 &  x716 &  x725 &  x728 &  x740 &  x747 &  x748 &  x755 &  x758 &  x764 &  x770 &  x776 &  x779 &  x786 &  x787 &  x788 &  x797 &  x803 &  x809 &  x815 &  x821 &  x824 &  x825 &  x826 &  x842 &  x854 &  x865 &  x872 &  x878 &  x890 &  x893 &  x896 &  x902 &  x904 &  x911 &  x917 &  x920 &  x926 &  x929 &  x935 &  x941 &  x943 &  x950 &  x959 &  x962 &  x965 &  x971 &  x983 &  x1001 &  x1004 &  x1013 &  x1016 &  x1022 &  x1037 &  x1043 &  x1052 &  x1061 &  x1064 &  x1070 &  x1073 &  x1079 &  x1082 &  x1091 &  x1100 &  x1106 &  x1112 &  x1118 &  x1121 & ~x492 & ~x705 & ~x744 & ~x745 & ~x783 & ~x784 & ~x822 & ~x861 & ~x900;
assign c7294 =  x17 &  x20 &  x35 &  x47 &  x59 &  x68 &  x86 &  x128 &  x131 &  x140 &  x197 &  x209 &  x212 &  x221 &  x239 &  x245 &  x248 &  x260 &  x275 &  x281 &  x320 &  x335 &  x350 &  x383 &  x434 &  x438 &  x439 &  x440 &  x442 &  x478 &  x494 &  x508 &  x509 &  x517 &  x524 &  x557 &  x569 &  x581 &  x586 &  x593 &  x644 &  x650 &  x656 &  x662 &  x677 &  x695 &  x703 &  x731 &  x755 &  x758 &  x781 &  x821 &  x842 &  x866 &  x872 &  x890 &  x893 &  x911 &  x929 &  x935 &  x944 &  x980 &  x983 &  x1016 &  x1019 &  x1034 &  x1043 &  x1067 &  x1106 &  x1118 & ~x276 & ~x465 & ~x474 & ~x552 & ~x591 & ~x861 & ~x862 & ~x940 & ~x979;
assign c7296 =  x41 &  x53 &  x131 &  x140 &  x194 &  x205 &  x209 &  x212 &  x221 &  x236 &  x242 &  x278 &  x352 &  x359 &  x419 &  x428 &  x467 &  x469 &  x509 &  x635 &  x670 &  x708 &  x747 &  x748 &  x787 &  x826 &  x857 &  x865 &  x904 &  x929 &  x938 &  x941 &  x977 &  x1013 &  x1019 &  x1046 &  x1052 &  x1100 & ~x745;
assign c7298 =  x35 &  x41 &  x56 &  x77 &  x119 &  x179 &  x209 &  x212 &  x224 &  x260 &  x265 &  x287 &  x292 &  x320 &  x331 &  x350 &  x383 &  x422 &  x446 &  x467 &  x473 &  x509 &  x517 &  x524 &  x569 &  x581 &  x602 &  x620 &  x689 &  x779 &  x781 &  x836 &  x842 &  x857 &  x872 &  x890 &  x902 &  x935 &  x959 &  x983 &  x986 &  x1004 &  x1019 &  x1043 &  x1046 &  x1106 & ~x0 & ~x39 & ~x78 & ~x117 & ~x156 & ~x276 & ~x471 & ~x940 & ~x979 & ~x1057 & ~x1096;
assign c71 =  x472 &  x790 &  x832 & ~x600 & ~x741;
assign c73 =  x198 &  x1027 &  x1081;
assign c75 =  x585 &  x784 &  x862;
assign c77 =  x1057 & ~x313;
assign c79 =  x407 &  x674 &  x733 &  x769 &  x799 &  x916 &  x925 &  x1024 &  x1085 & ~x786 & ~x825 & ~x1056;
assign c711 =  x239 &  x278 &  x338 &  x380 &  x398 &  x605 &  x662 &  x940 &  x1013 &  x1055 &  x1057 &  x1096 & ~x87 & ~x165 & ~x243 & ~x282 & ~x321 & ~x870;
assign c713 =  x355 &  x532 &  x799 &  x934 & ~x1098;
assign c715 =  x26 &  x29 &  x101 &  x128 &  x136 &  x221 &  x371 &  x443 &  x656 &  x695 &  x784 &  x823 &  x854 &  x862 &  x901 &  x940 &  x979 &  x1073 &  x1082 &  x1088 &  x1091 & ~x237;
assign c717 =  x28 &  x780 &  x1018 & ~x3;
assign c719 =  x433 & ~x600 & ~x813 & ~x996 & ~x1014;
assign c721 =  x532 &  x897 &  x1057 &  x1102 & ~x825 & ~x909;
assign c723 =  x115 &  x861 &  x1096;
assign c725 =  x72 &  x133 &  x319 & ~x120 & ~x159 & ~x477 & ~x516 & ~x1020;
assign c727 =  x319 &  x472 & ~x403;
assign c729 =  x727 & ~x742;
assign c731 =  x176 &  x269 &  x397 &  x527 &  x908 &  x1070 &  x1102 & ~x621 & ~x711 & ~x747 & ~x825 & ~x855 & ~x864;
assign c733 =  x433 &  x449 &  x472 &  x511 &  x550 &  x587 &  x790 & ~x405 & ~x441 & ~x444;
assign c735 =  x22 &  x150 &  x151 &  x379 &  x397 & ~x558 & ~x726 & ~x1059;
assign c737 =  x355 &  x394 &  x676 &  x733 &  x778 &  x799 &  x838 &  x949 &  x961;
assign c739 =  x745 &  x823 &  x985 &  x1062 & ~x714;
assign c741 = ~x105 & ~x265 & ~x624;
assign c743 =  x124 & ~x645 & ~x963 & ~x1014;
assign c745 =  x76 &  x319 &  x511 & ~x477 & ~x1098;
assign c747 =  x355 & ~x291 & ~x483 & ~x561 & ~x735 & ~x930 & ~x1074;
assign c749 =  x471 &  x610 & ~x3;
assign c753 =  x76 &  x433 &  x1027 &  x1066 & ~x324;
assign c755 =  x14 &  x56 &  x74 &  x85 &  x124 &  x164 &  x215 &  x230 &  x236 &  x332 &  x341 &  x422 &  x434 &  x461 &  x488 &  x497 &  x530 &  x578 &  x586 &  x599 &  x605 &  x623 &  x713 &  x833 &  x860 &  x884 &  x893 &  x911 &  x917 &  x938 &  x941 &  x1070 &  x1073 &  x1094 & ~x246 & ~x285 & ~x324 & ~x441 & ~x1059 & ~x1098;
assign c757 =  x550 &  x949 & ~x1093;
assign c759 =  x232 &  x236 &  x290 &  x365 &  x397 &  x512 &  x668 &  x827 & ~x555 & ~x747 & ~x786 & ~x825 & ~x876 & ~x1098;
assign c761 = ~x347;
assign c763 =  x978 & ~x973;
assign c765 =  x368 &  x979 & ~x391 & ~x753 & ~x792;
assign c767 =  x225 & ~x520;
assign c769 =  x237 &  x988;
assign c771 =  x334 & ~x558 & ~x562 & ~x732;
assign c773 =  x472 &  x805 & ~x600 & ~x813;
assign c775 = ~x360 & ~x555 & ~x636 & ~x1098;
assign c777 =  x901 & ~x276 & ~x871 & ~x1005;
assign c779 =  x193 &  x310 & ~x105 & ~x261 & ~x516 & ~x555 & ~x1125;
assign c781 =  x237 & ~x367 & ~x444 & ~x862;
assign c783 =  x731 &  x1096 & ~x9 & ~x204 & ~x516 & ~x561 & ~x711;
assign c785 =  x271 &  x861 &  x1057;
assign c787 =  x28 &  x133 &  x262 &  x397 &  x410 &  x1102 & ~x621 & ~x672 & ~x825 & ~x1059 & ~x1116;
assign c789 =  x46 &  x829 & ~x363 & ~x1098 & ~x1125;
assign c791 =  x1024 & ~x562;
assign c793 =  x393 &  x550 &  x676 & ~x1095;
assign c797 =  x23 &  x173 &  x206 &  x293 &  x338 &  x452 &  x635 &  x665 &  x794 &  x901 &  x938 &  x940 &  x944 &  x947 &  x978 &  x992 &  x995 &  x1057 &  x1067 &  x1070 &  x1097 & ~x870;
assign c799 =  x73 &  x100 &  x745 &  x823 &  x862 &  x880 & ~x1098;
assign c7101 =  x7 &  x1096 & ~x325;
assign c7103 =  x433 & ~x403;
assign c7105 =  x115 &  x823 &  x900 &  x940 &  x1057 & ~x312 & ~x432;
assign c7107 =  x237 & ~x12 & ~x106 & ~x300;
assign c7109 =  x76 &  x511 & ~x519 & ~x963 & ~x1074 & ~x1113;
assign c7111 =  x139 &  x178 &  x901 &  x1102 & ~x3 & ~x114;
assign c7113 =  x586 &  x628 &  x823 & ~x427;
assign c7115 =  x34 &  x73 &  x80 &  x92 &  x170 &  x266 &  x359 &  x374 &  x509 &  x629 &  x710 &  x745 &  x784 &  x869 &  x902 &  x935 &  x947 & ~x636 & ~x1020;
assign c7117 =  x89 &  x155 &  x158 &  x206 &  x335 &  x704 &  x713 &  x741 &  x875 &  x881 &  x920 &  x940 &  x983 &  x1018 &  x1019 &  x1043 &  x1058 &  x1061 & ~x315;
assign c7119 =  x115 &  x706 &  x940 &  x979 &  x1066;
assign c7121 =  x585 & ~x520 & ~x826;
assign c7123 =  x28 &  x139 &  x223 &  x262 &  x347 &  x437 &  x494 &  x608 &  x784 &  x823 &  x914 &  x1018 &  x1081;
assign c7125 =  x16 &  x28 &  x68 &  x80 &  x109 &  x182 &  x245 &  x407 &  x518 &  x542 &  x635 &  x644 &  x745 &  x782 &  x784 &  x902 &  x908 &  x911 &  x917 &  x920 &  x923 &  x935 &  x968 &  x1001 &  x1018 &  x1064;
assign c7127 =  x823 &  x1023 & ~x873 & ~x876;
assign c7129 =  x227 &  x355 &  x532 &  x571 &  x715 &  x955 &  x973 & ~x1095;
assign c7131 =  x396 &  x472 &  x511 & ~x480;
assign c7133 =  x733 &  x799 &  x838 &  x1081 & ~x309 & ~x825;
assign c7135 =  x358 & ~x199 & ~x558 & ~x1099;
assign c7137 =  x489 & ~x523;
assign c7139 =  x780 &  x862 &  x1018 &  x1057 &  x1102;
assign c7141 =  x472 &  x511 &  x760 &  x799 & ~x459 & ~x1095;
assign c7143 =  x237 &  x559 &  x871 & ~x207 & ~x1047;
assign c7145 =  x115 &  x232 &  x823 &  x899 &  x1018 & ~x714;
assign c7147 =  x742 &  x745 &  x784 & ~x3 & ~x276 & ~x504 & ~x1020;
assign c7149 =  x72 &  x1057 & ~x3;
assign c7151 =  x355 &  x844 &  x1027 &  x1066 & ~x600 & ~x813;
assign c7153 =  x823 &  x862 &  x901 & ~x42 & ~x121 & ~x160;
assign c7155 =  x14 &  x217 &  x262 &  x338 &  x745 &  x758 &  x784 & ~x18 & ~x1020 & ~x1095;
assign c7157 =  x531 &  x888 & ~x742;
assign c7159 = ~x638;
assign c7161 =  x511 &  x1027 & ~x561 & ~x813 & ~x1053 & ~x1074;
assign c7163 =  x178 &  x302 &  x313 &  x419 &  x449 &  x461 &  x623 &  x659 &  x698 &  x740 &  x833 &  x907 &  x911 &  x946 &  x983 &  x1042 &  x1061 &  x1102 & ~x12 & ~x24 & ~x114 & ~x324;
assign c7165 =  x643 &  x655 &  x907 &  x1081 & ~x63 & ~x825;
assign c7167 =  x276 &  x556 & ~x168 & ~x261;
assign c7169 =  x822 & ~x234 & ~x849;
assign c7171 =  x394 &  x433 &  x799 & ~x781;
assign c7173 =  x355 &  x433 &  x593 &  x838 &  x844 &  x883 &  x895 &  x988 &  x994;
assign c7175 =  x73 &  x262 &  x862 & ~x24 & ~x348 & ~x1020;
assign c7177 =  x158 &  x229 &  x248 &  x702 &  x901 &  x940 &  x1130 & ~x849;
assign c7179 =  x44 &  x83 &  x122 &  x155 &  x185 &  x269 &  x298 &  x344 &  x365 &  x467 &  x512 &  x515 &  x602 &  x614 &  x745 &  x784 &  x818 &  x830 &  x842 &  x896 &  x911 &  x926 &  x940 &  x979 &  x1007 &  x1049 &  x1103 & ~x273 & ~x312 & ~x654;
assign c7181 =  x351 & ~x51 & ~x325;
assign c7183 =  x71 &  x317 &  x347 &  x497 &  x745 &  x784 &  x815 &  x823 &  x857 &  x862 &  x901 &  x940 &  x947 & ~x156 & ~x849 & ~x1047;
assign c7185 =  x237 &  x316 & ~x247 & ~x250;
assign c7187 =  x940 &  x978 &  x1096 &  x1097 & ~x390 & ~x870;
assign c7189 =  x502 & ~x9 & ~x87 & ~x261 & ~x669;
assign c7191 = ~x169 & ~x261 & ~x1053;
assign c7193 =  x472 & ~x4 & ~x360;
assign c7195 =  x355 &  x593 & ~x285 & ~x342 & ~x1014 & ~x1056;
assign c7197 =  x751 &  x844 &  x910 & ~x247 & ~x285;
assign c7199 =  x397 & ~x934 & ~x1068;
assign c7201 =  x85 &  x124 &  x217 &  x871 & ~x360 & ~x651;
assign c7203 =  x277 &  x739 &  x772 &  x778 &  x793 &  x799 &  x1040 & ~x1095;
assign c7205 = ~x524;
assign c7207 =  x277 &  x643 &  x655 &  x733 & ~x247;
assign c7209 =  x784 & ~x199 & ~x636 & ~x1059;
assign c7211 =  x634 & ~x51 & ~x897;
assign c7213 =  x472 & ~x402 & ~x561 & ~x936;
assign c7215 =  x28 &  x745 &  x955;
assign c7217 =  x139 &  x799 &  x1063 &  x1102 & ~x459 & ~x825 & ~x903;
assign c7219 =  x115 & ~x555 & ~x594 & ~x670 & ~x786;
assign c7221 =  x76 &  x232 &  x310 &  x901 & ~x477 & ~x672 & ~x789;
assign c7223 =  x784 &  x862 &  x945 & ~x714;
assign c7225 =  x124 &  x745 &  x1018 &  x1096 & ~x894;
assign c7227 = ~x364 & ~x405;
assign c7229 =  x472 &  x799 &  x805 &  x832 &  x838 &  x871 &  x889 &  x895;
assign c7231 =  x237 &  x799 & ~x625;
assign c7233 = ~x303;
assign c7235 = ~x360 & ~x810 & ~x928 & ~x1068;
assign c7237 =  x34 &  x124 &  x827 &  x1016 & ~x564 & ~x825 & ~x981;
assign c7239 = ~x313 & ~x952;
assign c7241 =  x511 &  x745 & ~x120 & ~x1113 & ~x1119;
assign c7243 = ~x170;
assign c7245 =  x73 &  x1075 & ~x12 & ~x24 & ~x51 & ~x75 & ~x207 & ~x477 & ~x1020;
assign c7247 =  x1018 &  x1024 & ~x753;
assign c7249 = ~x494;
assign c7251 =  x355 &  x675 &  x934 &  x1012 &  x1033 & ~x1053;
assign c7253 =  x119 &  x214 &  x319 & ~x750 & ~x864 & ~x903 & ~x904 & ~x942;
assign c7255 =  x355 &  x433 & ~x781;
assign c7257 =  x20 &  x544 &  x643 &  x769 &  x797 &  x985 &  x1042 &  x1081 & ~x207 & ~x246 & ~x285;
assign c7259 =  x298 & ~x243 & ~x559;
assign c7261 =  x472 & ~x403 & ~x897;
assign c7263 =  x315 &  x355 &  x636 & ~x1092;
assign c7265 =  x646 &  x877 &  x907 &  x1081 &  x1102 & ~x207 & ~x303;
assign c7267 =  x128 &  x571 &  x1018 &  x1081 & ~x114;
assign c7269 =  x315 &  x1012 & ~x703;
assign c7271 =  x95 &  x124 &  x217 &  x248 &  x278 &  x383 &  x416 &  x674 &  x677 &  x686 &  x692 &  x1061 &  x1112 & ~x282 & ~x321 & ~x867 & ~x942;
assign c7273 =  x900 & ~x870;
assign c7275 =  x59 &  x646 &  x663 &  x745 & ~x597;
assign c7277 =  x355 &  x433 &  x766 &  x778 &  x793 &  x805 &  x955;
assign c7279 =  x550 &  x706 &  x838 & ~x639 & ~x1059;
assign c7281 =  x550 &  x973 & ~x81 & ~x441;
assign c7283 =  x16 &  x34 &  x94 &  x139 &  x767 &  x784 &  x823 &  x986 & ~x636 & ~x714;
assign c7285 =  x806 &  x886 &  x985 & ~x321 & ~x444 & ~x477;
assign c7287 =  x542 &  x550 &  x790 & ~x717 & ~x780;
assign c7291 =  x907 & ~x247 & ~x1014;
assign c7293 =  x125 &  x173 &  x235 &  x461 &  x479 &  x655 &  x1079 &  x1102 & ~x63 & ~x90 & ~x162 & ~x303 & ~x669 & ~x825 & ~x903 & ~x981 & ~x1020 & ~x1098;
assign c7295 =  x271 &  x641 & ~x261 & ~x360 & ~x555 & ~x768 & ~x807;
assign c7297 =  x77 &  x85 &  x119 &  x124 &  x163 &  x175 &  x202 &  x215 &  x233 &  x275 &  x280 &  x319 &  x413 &  x488 &  x506 &  x788 &  x901 &  x940 &  x956 &  x980 &  x1025 &  x1057 &  x1096;
assign c7299 =  x139 &  x772 &  x1109 & ~x207 & ~x342 & ~x480 & ~x498;

endmodule