module tm( x0,x1,x2,x3,x4,x5,x6,x7,x8,x9,x10,x11,x12,x13,x14,x15,x16,x17,x18,x19,x20,x21,x22,x23,x24,x25,x26,x27,x28,x29,x30,x31,x32,x33,x34,x35,x36,x37,x38,x39,x40,x41,x42,x43,x44,x45,x46,x47,x48,x49,x50,x51,x52,x53,x54,x55,x56,x57,x58,x59,x60,x61,x62,x63,x64,x65,x66,x67,x68,x69,x70,x71,x72,x73,x74,x75,x76,x77,x78,x79,x80,x81,x82,x83,x84,x85,x86,x87,x88,x89,x90,x91,x92,x93,x94,x95,x96,x97,x98,x99,x100,x101,x102,x103,x104,x105,x106,x107,x108,x109,x110,x111,x112,x113,x114,x115,x116,x117,x118,x119,x120,x121,x122,x123,x124,x125,x126,x127,x128,x129,x130,x131,x132,x133,x134,x135,x136,x137,x138,x139,x140,x141,x142,x143,x144,x145,x146,x147,x148,x149,x150,x151,x152,x153,x154,x155,x156,x157,x158,x159,x160,x161,x162,x163,x164,x165,x166,x167,x168,x169,x170,x171,x172,x173,x174,x175,x176,x177,x178,x179,x180,x181,x182,x183,x184,x185,x186,x187,x188,x189,x190,x191,x192,x193,x194,x195,x196,x197,x198,x199,x200,x201,x202,x203,x204,x205,x206,x207,x208,x209,x210,x211,x212,x213,x214,x215,x216,x217,x218,x219,x220,x221,x222,x223,x224,x225,x226,x227,x228,x229,x230,x231,x232,x233,x234,x235,x236,x237,x238,x239,x240,x241,x242,x243,x244,x245,x246,x247,x248,x249,x250,x251,x252,x253,x254,x255,x256,x257,x258,x259,x260,x261,x262,x263,x264,x265,x266,x267,x268,x269,x270,x271,x272,x273,x274,x275,x276,x277,x278,x279,x280,x281,x282,x283,x284,x285,x286,x287,x288,x289,x290,x291,x292,x293,x294,x295,x296,x297,x298,x299,x300,x301,x302,x303,x304,x305,x306,x307,x308,x309,x310,x311,x312,x313,x314,x315,x316,x317,x318,x319,x320,x321,x322,x323,x324,x325,x326,x327,x328,x329,x330,x331,x332,x333,x334,x335,x336,x337,x338,x339,x340,x341,x342,x343,x344,x345,x346,x347,x348,x349,x350,x351,x352,x353,x354,x355,x356,x357,x358,x359,x360,x361,x362,x363,x364,x365,x366,x367,x368,x369,x370,x371,x372,x373,x374,x375,x376,x377,x378,x379,x380,x381,x382,x383,x384,x385,x386,x387,x388,x389,x390,x391,x392,x393,x394,x395,x396,x397,x398,x399,x400,x401,x402,x403,x404,x405,x406,x407,x408,x409,x410,x411,x412,x413,x414,x415,x416,x417,x418,x419,x420,x421,x422,x423,x424,x425,x426,x427,x428,x429,x430,x431,x432,x433,x434,x435,x436,x437,x438,x439,x440,x441,x442,x443,x444,x445,x446,x447,x448,x449,x450,x451,x452,x453,x454,x455,x456,x457,x458,x459,x460,x461,x462,x463,x464,x465,x466,x467,x468,x469,x470,x471,x472,x473,x474,x475,x476,x477,x478,x479,x480,x481,x482,x483,x484,x485,x486,x487,x488,x489,x490,x491,x492,x493,x494,x495,x496,x497,x498,x499,x500,x501,x502,x503,x504,x505,x506,x507,x508,x509,x510,x511,x512,x513,x514,x515,x516,x517,x518,x519,x520,x521,x522,x523,x524,x525,x526,x527,x528,x529,x530,x531,x532,x533,x534,x535,x536,x537,x538,x539,x540,x541,x542,x543,x544,x545,x546,x547,x548,x549,x550,x551,x552,x553,x554,x555,x556,x557,x558,x559,x560,x561,x562,x563,x564,x565,x566,x567,x568,x569,x570,x571,x572,x573,x574,x575,x576,x577,x578,x579,x580,x581,x582,x583,x584,x585,x586,x587,x588,x589,x590,x591,x592,x593,x594,x595,x596,x597,x598,x599,x600,x601,x602,x603,x604,x605,x606,x607,x608,x609,x610,x611,x612,x613,x614,x615,x616,x617,x618,x619,x620,x621,x622,x623,x624,x625,x626,x627,x628,x629,x630,x631,x632,x633,x634,x635,x636,x637,x638,x639,x640,x641,x642,x643,x644,x645,x646,x647,x648,x649,x650,x651,x652,x653,x654,x655,x656,x657,x658,x659,x660,x661,x662,x663,x664,x665,x666,x667,x668,x669,x670,x671,x672,x673,x674,x675,x676,x677,x678,x679,x680,x681,x682,x683,x684,x685,x686,x687,x688,x689,x690,x691,x692,x693,x694,x695,x696,x697,x698,x699,x700,x701,x702,x703,x704,x705,x706,x707,x708,x709,x710,x711,x712,x713,x714,x715,x716,x717,x718,x719,x720,x721,x722,x723,x724,x725,x726,x727,x728,x729,x730,x731,x732,x733,x734,x735,x736,x737,x738,x739,x740,x741,x742,x743,x744,x745,x746,x747,x748,x749,x750,x751,x752,x753,x754,x755,x756,x757,x758,x759,x760,x761,x762,x763,x764,x765,x766,x767,x768,x769,x770,x771,x772,x773,x774,x775,x776,x777,x778,x779,x780,x781,x782,x783,c3401,c1490,c5398,c7286,c439,c8240,c947,c4206,c2455,c152,c9300,c1113,c079,c3229,c8483,c969,c0269,c0366,c3285,c2162,c196,c3187,c8271,c136,c8471,c3480,c0371,c8104,c8242,c4330,c679,c6498,c5202,c5341,c473,c7454,c950,c6430,c6416,c6252,c298,c2366,c6422,c7102,c6294,c613,c753,c866,c0120,c8491,c7231,c195,c0334,c215,c1200,c2224,c54,c6353,c736,c7330,c1346,c4456,c8252,c3264,c137,c5319,c9241,c5363,c134,c6370,c7457,c4226,c5272,c7333,c8453,c1318,c371,c4183,c2298,c9210,c3391,c9196,c5484,c5451,c6327,c1498,c0381,c0415,c5339,c8468,c4460,c1411,c4110,c6113,c2313,c0324,c4348,c7345,c9322,c2426,c673,c9408,c4319,c4358,c9244,c3235,c4401,c531,c9165,c2367,c1465,c3299,c31,c6130,c3462,c773,c034,c8345,c5335,c7250,c7147,c8322,c2260,c4259,c2241,c395,c644,c1342,c8108,c6271,c5478,c619,c7285,c3303,c5224,c6278,c1316,c990,c3288,c6232,c479,c2218,c0491,c725,c6166,c6427,c4293,c1388,c6381,c970,c1353,c4222,c8245,c9329,c2108,c4404,c7464,c9164,c7271,c713,c1299,c4162,c7200,c5216,c5197,c8297,c3322,c9104,c284,c7223,c6142,c8109,c5294,c15,c655,c6339,c1275,c241,c636,c6249,c1420,c5191,c855,c1432,c7221,c1234,c3387,c676,c8436,c3461,c7213,c563,c1327,c3298,c5220,c4363,c2429,c1231,c3376,c3177,c8118,c3381,c6291,c211,c8329,c3443,c1466,c3331,c6434,c7182,c589,c7280,c3478,c7365,c6272,c364,c4291,c2267,c3195,c1469,c3252,c7337,c818,c3199,c0463,c0455,c917,c2114,c0123,c6264,c3435,c7245,c75,c9381,c3441,c4158,c1373,c7311,c0449,c3188,c7485,c1291,c6101,c1247,c3368,c6388,c2436,c2169,c143,c5252,c0487,c0256,c6236,c0435,c1340,c3448,c4414,c865,c8192,c6103,c3231,c7488,c2486,c3428,c3207,c6305,c233,c487,c8190,c0157,c9222,c9268,c8200,c3330,c0335,c6350,c5177,c2179,c5218,c3297,c2184,c3383,c7355,c0175,c5413,c1328,c5338,c5133,c992,c728,c0474,c89,c0447,c653,c7346,c711,c263,c914,c166,c7321,c7323,c7297,c7387,c8390,c9110,c942,c8466,c1106,c9371,c4114,c4221,c2322,c7450,c794,c0212,c4224,c553,c2269,c341,c8400,c2402,c3247,c0244,c4235,c76,c4495,c7113,c4230,c06,c8432,c9434,c9145,c7414,c161,c8125,c0254,c6100,c420,c7371,c8480,c640,c1268,c4428,c576,c6359,c458,c2462,c090,c3116,c5105,c690,c9308,c5258,c545,c0227,c462,c9201,c3417,c710,c443,c6231,c7139,c5350,c261,c1225,c0482,c5163,c9203,c3390,c2473,c6431,c789,c5382,c1241,c3260,c391,c0468,c081,c9160,c0428,c0265,c712,c5183,c8404,c2188,c6445,c2432,c859,c5389,c6367,c6243,c0287,c7194,c7195,c0398,c8127,c4246,c3342,c8235,c7201,c8144,c471,c3216,c6451,c556,c3238,c33,c2453,c0427,c2122,c9292,c8310,c5136,c0483,c8318,c7209,c933,c839,c862,c3282,c8462,c8237,c8317,c1453,c8267,c5275,c3453,c7149,c1159,c951,c6380,c3174,c2444,c3254,c6450,c2472,c9162,c8444,c8472,c7219,c8306,c3436,c3464,c1240,c2150,c6493,c4487,c3361,c4269,c6241,c4125,c8319,c9426,c287,c5357,c0253,c5390,c8187,c9346,c7421,c6134,c1473,c2204,c8386,c8259,c1398,c9126,c0306,c863,c1155,c6334,c237,c071,c62,c749,c7172,c7352,c431,c7498,c5140,c5443,c1153,c083,c040,c218,c9141,c7494,c5376,c0350,c5381,c9149,c0125,c6242,c2126,c3477,c4225,c7409,c2239,c0281,c8223,c1127,c6171,c4204,c8403,c1248,c1441,c212,c8183,c9199,c7295,c6131,c8156,c0189,c1306,c2450,c0264,c7165,c5166,c3371,c258,c5142,c1363,c9475,c6330,c4313,c91,c987,c6382,c3408,c8478,c9343,c850,c4106,c7445,c5474,c4413,c498,c6110,c7410,c4470,c7325,c1492,c068,c9299,c188,c025,c6136,c551,c7395,c1108,c423,c788,c3313,c2198,c8191,c9198,c8464,c9236,c61,c0387,c4100,c4177,c4129,c5115,c3122,c8388,c5119,c699,c5269,c482,c3409,c812,c3220,c9447,c784,c7444,c5471,c9364,c8314,c2401,c5238,c340,c3319,c9115,c1220,c6296,c0144,c0198,c1481,c2306,c2483,c0365,c9266,c8338,c0156,c2297,c4433,c9209,c046,c5212,c6155,c2248,c6220,c6146,c6317,c3492,c493,c573,c717,c2255,c9250,c076,c0304,c5372,c1372,c2328,c7456,c766,c0229,c5486,c4190,c0394,c9390,c8307,c5404,c1415,c0258,c4327,c8331,c348,c7292,c5309,c8206,c3159,c6248,c9180,c250,c6208,c3402,c7356,c339,c2112,c6384,c4290,c0214,c3283,c7117,c3400,c8397,c9288,c5113,c4402,c7307,c3148,c777,c6428,c7400,c1167,c0297,c623,c012,c2499,c9175,c3339,c6436,c7234,c321,c6293,c4390,c5491,c0465,c7279,c3194,c2156,c2430,c5282,c5380,c6214,c0312,c543,c0112,c396,c894,c3175,c4335,c9430,c8167,c5375,c0280,c021,c483,c0457,c6304,c1228,c7112,c5316,c6153,c6132,c0382,c199,c0385,c7125,c1475,c9176,c4176,c7141,c7226,c9304,c4196,c5345,c8325,c518,c1180,c2181,c8333,c6139,c5203,c650,c4112,c4325,c3263,c8258,c8262,c964,c9453,c1381,c7393,c9135,c3259,c4217,c189,c7495,c2186,c4374,c5296,c0400,c4130,c7187,c3241,c6473,c8399,c5280,c110,c1209,c635,c519,c5233,c6412,c1134,c612,c9310,c4286,c3485,c7374,c828,c2484,c4160,c3350,c617,c3149,c3218,c4298,c7466,c8121,c0218,c117,c289,c6140,c0126,c056,c3192,c3294,c2403,c4408,c674,c2476,c6224,c5353,c989,c3336,c4480,c4145,c5435,c0476,c7242,c547,c5368,c4139,c2318,c8215,c1238,c9182,c844,c4107,c4279,c1164,c194,c746,c8286,c7217,c3173,c3483,c0338,c891,c0127,c5449,c2394,c4387,c583,c1128,c834,c172,c2138,c760,c4321,c2201,c669,c4435,c4189,c0456,c4416,c0442,c6477,c3333,c835,c6141,c5208,c359,c5124,c610,c6483,c6230,c1282,c71,c525,c2203,c0135,c7150,c82,c848,c0110,c169,c1197,c7294,c9465,c4429,c4334,c0376,c8236,c447,c5165,c3459,c6240,c452,c2101,c3106,c9163,c0215,c5242,c125,c63,c765,c0163,c4193,c414,c4243,c114,c974,c4205,c3234,c22,c7233,c0369,c3410,c9116,c2194,c0409,c3332,c3171,c4257,c7246,c2358,c6297,c979,c3165,c3343,c4339,c7127,c0174,c572,c2331,c3181,c790,c8363,c575,c593,c0329,c366,c570,c4281,c6426,c1468,c4137,c167,c0310,c4120,c9237,c822,c0496,c080,c6184,c181,c3245,c5193,c6341,c7434,c825,c5460,c7403,c9290,c316,c6108,c5226,c4273,c6250,c9332,c956,c1349,c450,c171,c779,c6210,c1196,c976,c28,c8327,c982,c840,c0300,c1311,c6383,c7303,c2123,c5109,c7220,c6443,c3164,c7426,c2339,c5239,c3112,c1345,c1283,c5446,c7310,c665,c4352,c9356,c795,c2332,c4449,c8248,c9138,c8184,c8112,c9464,c6326,c0141,c07,c3270,c4212,c5384,c6345,c7357,c9369,c8175,c5118,c4295,c0116,c3365,c4307,c48,c7439,c0425,c2315,c0454,c8202,c9151,c2151,c4288,c1190,c6259,c9183,c6127,c7190,c8168,c780,c2434,c9384,c434,c4373,c6183,c3138,c160,c8186,c8456,c9234,c6352,c7477,c3424,c8394,c5402,c2288,c0453,c030,c2414,c4102,c4333,c1269,c4474,c2102,c857,c7133,c2423,c3243,c4447,c2235,c1243,c5123,c9276,c1150,c2246,c356,c9321,c577,c0140,c0313,c2498,c1211,c684,c1455,c0302,c3135,c2487,c3121,c888,c2145,c1274,c9494,c7342,c5168,c1338,c2304,c819,c1111,c4410,c1360,c5255,c4135,c9136,c3414,c4317,c5304,c6470,c7120,c3244,c1221,c7389,c1380,c072,c6129,c2404,c7230,c0199,c873,c5434,c2243,c911,c7399,c1483,c7467,c0275,c0337,c9233,c9281,c8197,c5205,c675,c7416,c1391,c3153,c846,c5321,c1460,c7351,c836,c3266,c381,c4371,c9121,c9311,c2211,c5122,c5217,c9345,c8169,c6338,c4260,c530,c9286,c8123,c14,c0498,c8298,c4418,c745,c149,c3219,c8342,c4364,c843,c8376,c3226,c5361,c3119,c2433,c7132,c775,c3262,c213,c3422,c7316,c7288,c3305,c4232,c5222,c3446,c9320,c9347,c6356,c4493,c0240,c177,c0402,c0160,c6209,c4454,c7218,c031,c2466,c3113,c0448,c9229,c6363,c8194,c0315,c6168,c6206,c6314,c0416,c3484,c6397,c754,c2431,c5179,c9471,c5388,c8225,c8229,c392,c4452,c6195,c5236,c7274,c427,c275,c8295,c4385,c418,c5427,c896,c9350,c5150,c5495,c4486,c4461,c629,c9359,c435,c3460,c1419,c2361,c925,c4415,c3102,c7479,c7180,c639,c3248,c5303,c469,c324,c1129,c662,c6275,c0327,c7106,c6467,c0401,c1174,c226,c2311,c932,c5181,c5129,c7465,c4328,c668,c0161,c68,c842,c049,c2289,c78,c7227,c5470,c5442,c8341,c496,c1255,c9108,c4168,c0311,c5359,c0115,c093,c7487,c9275,c9267,c5180,c8401,c2352,c279,c9440,c5106,c9212,c353,c95,c772,c9194,c3169,c8357,c1203,c7244,c4430,c1204,c6105,c3139,c9386,c5270,c9122,c2441,c569,c9442,c7343,c637,c8135,c5171,c6219,c743,c1384,c759,c098,c2442,c4383,c590,c3431,c0231,c7304,c3337,c4157,c1448,c2369,c468,c2277,c1280,c6286,c7305,c1343,c8359,c43,c6449,c7455,c84,c6119,c8181,c730,c4265,c7211,c3327,c8230,c4375,c8385,c5128,c1326,c889,c6182,c3452,c7140,c3329,c7257,c72,c8281,c692,c515,c7151,c955,c4432,c2368,c2425,c1216,c2301,c9134,c8178,c810,c5286,c560,c128,c4367,c1229,c6281,c8162,c8154,c3198,c6411,c3438,c3257,c2355,c7459,c4141,c6178,c2412,c0462,c9353,c387,c881,c7348,c8113,c2270,c9481,c3114,c3205,c1301,c3221,c1145,c3103,c9366,c0344,c5188,c440,c1329,c8365,c7329,c1287,c2159,c2262,c1371,c2274,c8343,c8373,c426,c582,c6116,c4331,c0220,c6179,c075,c2475,c4147,c5134,c7196,c1207,c7255,c6161,c1487,c0285,c4151,c6435,c5433,c315,c1339,c0249,c1140,c6458,c086,c1452,c5201,c2494,c111,c9449,c8459,c6223,c2175,c1124,c8351,c7484,c3454,c8347,c5457,c4411,c6292,c6124,c4136,c8448,c0323,c2464,c323,c5211,c2386,c0478,c0388,c7388,c0467,c5137,c5172,c8222,c1489,c9216,c0352,c2215,c9252,c9223,c9277,c268,c3228,c7162,c312,c9263,c2392,c4292,c592,c2164,c895,c9396,c965,c5189,c9291,c6313,c1114,c916,c1296,c085,c1232,c9309,c9407,c3240,c7447,c5110,c8411,c9107,c2193,c3306,c7283,c2479,c4266,c5302,c5424,c4194,c7490,c0472,c478,c9477,c3384,c1142,c7349,c633,c1257,c7225,c0331,c6306,c786,c36,c8176,c6322,c647,c9363,c3489,c3184,c052,c6320,c2439,c1364,c7273,c8257,c5408,c7236,c2185,c0274,c4166,c8484,c722,c9181,c354,c1401,c0164,c063,c8330,c2252,c5223,c475,c7458,c4301,c2146,c7469,c4372,c8410,c7378,c6174,c796,c4312,c9358,c0404,c7142,c059,c6181,c0370,c9451,c3321,c033,c4250,c752,c3267,c7193,c8247,c9178,c0348,c3211,c1271,c4494,c88,c4475,c0403,c0250,c628,c77,c3287,c9344,c4285,c7110,c5441,c4153,c8114,c3307,c2183,c5334,c9326,c2343,c3268,c9285,c1400,c4437,c4329,c6328,c16,c757,c131,c1183,c37,c4308,c884,c7446,c9226,c9114,c4417,c967,c4439,c6246,c2163,c3364,c7436,c0145,c3251,c7402,c5245,c5156,c7478,c245,c4150,c7468,c069,c5412,c17,c521,c257,c6390,c876,c5263,c4473,c0206,c9456,c1244,c0173,c2353,c8469,c4490,c6438,c56,c4116,c5248,c1480,c3326,c295,c1403,c817,c2259,c798,c599,c5432,c0192,c5186,c1166,c1252,c2417,c094,c7105,c1446,c0188,c6461,c0246,c1224,c6469,c2121,c689,c0417,c532,c42,c2247,c8221,c8250,c6347,c959,c2329,c9130,c6391,c9305,c998,c7100,c8292,c03,c4377,c0484,c5439,c1462,c5146,c078,c9379,c555,c296,c0405,c349,c3455,c574,c0266,c764,c4341,c5494,c7264,c9255,c0396,c7361,c9102,c347,c1214,c099,c1186,c1428,c4245,c5190,c1276,c2275,c7425,c8352,c6442,c2174,c7418,c6159,c1467,c34,c0392,c4214,c0397,c883,c813,c2314,c9156,c0113,c8487,c724,c8278,c755,c620,c7224,c731,c9186,c1109,c9211,c8253,c520,c0317,c0407,c3128,c6107,c5378,c962,c5315,c467,c4272,c8446,c9422,c45,c0309,c73,c548,c0142,c1152,c165,c3463,c2317,c7462,c5130,c0185,c0495,c552,c983,c7126,c2397,c3110,c0356,c8362,c8449,c6495,c7143,c1394,c5469,c8203,c491,c4237,c3272,c9144,c5452,c0460,c5237,c557,c7430,c112,c9323,c6454,c768,c7198,c8294,c4209,c2490,c1178,c1457,c792,c0339,c3362,c4173,c8336,c864,c2338,c2491,c984,c2154,c1437,c6394,c4247,c6118,c6480,c3423,c1181,c3232,c9499,c6419,c7101,c9485,c769,c5284,c3276,c122,c3214,c4197,c8101,c6269,c6408,c8498,c0393,c3356,c1350,c8420,c9303,c1223,c4202,c6463,c8243,c9306,c3354,c9242,c9120,c350,c9374,c8497,c5371,c838,c2229,c7207,c8289,c9432,c2292,c8296,c6488,c288,c8396,c3210,c7344,c9331,c0114,c4419,c0391,c3490,c2225,c1463,c8355,c8110,c3236,c9261,c373,c7491,c0191,c4356,c2419,c8208,c2468,c036,c3407,c791,c6482,c622,c1431,c961,c2197,c4315,c5173,c4398,c8427,c2155,c9433,c9296,c3233,c7214,c7319,c367,c264,c376,c4431,c645,c912,c7270,c4231,c060,c3355,c1456,c0284,c0421,c3166,c5182,c6409,c494,c3405,c9132,c8337,c3465,c4425,c524,c5214,c2172,c248,c7258,c1300,c8475,c2348,c977,c2460,c317,c6299,c4389,c8490,c4393,c7375,c0136,c6258,c4179,c8264,c8130,c2467,c4282,c824,c2461,c8389,c2321,c5403,c6444,c9395,c2384,c2233,c9490,c5445,c3386,c538,c915,c4164,c841,c1396,c9335,c041,c9105,c8321,c444,c6163,c8305,c9330,c0195,c0466,c2308,c0479,c6268,c5141,c6489,c0236,c937,c5326,c6122,c614,c1406,c9417,c1270,c0245,c7197,c9497,c8251,c413,c2242,c6192,c024,c2190,c4219,c0440,c0325,c5400,c3141,c762,c18,c5417,c0223,c8470,c1389,c0257,c529,c9123,c1488,c3304,c2228,c1491,c2111,c0117,c7204,c9462,c0438,c280,c3470,c641,c7239,c9167,c591,c7124,c0293,c5370,c018,c130,c1348,c9319,c4300,c671,c9169,c9450,c9314,c7266,c9192,c9455,c4472,c871,c2299,c6154,c1334,c0133,c4340,c1459,c285,c4304,c94,c718,c6282,c446,c7131,c5488,c5260,c5268,c6369,c3353,c140,c2359,c7496,c2128,c734,c8116,c9142,c1385,c2223,c930,c453,c7134,c5342,c0276,c4346,c6361,c089,c2438,c0434,c0259,c6287,c1298,c7160,c744,c2381,c1416,c5401,c0303,c7169,c6349,c2396,c8211,c9402,c3380,c6218,c0151,c3156,c8353,c7269,c3345,c7453,c8146,c7340,c3488,c3144,c6207,c7298,c8435,c5436,c0103,c9298,c5347,c0122,c2263,c9405,c973,c6111,c6490,c6355,c4233,c7390,c7287,c6298,c0341,c0459,c9348,c7372,c6439,c9370,c1193,c2363,c2496,c1235,c0295,c1254,c7184,c1279,c5479,c7115,c8131,c13,c93,c658,c6187,c0235,c1454,c9342,c7347,c6368,c497,c8474,c6216,c2178,c9385,c6485,c2210,c492,c1263,c8422,c338,c1286,c2236,c6312,c2360,c6365,c7384,c47,c6151,c170,c429,c7253,c2495,c9179,c0182,c0201,c2261,c3392,c8273,c0143,c9474,c9247,c3104,c921,c9172,c1239,c2349,c9297,c422,c0277,c0408,c2115,c9441,c2251,c0176,c9109,c2199,c019,c7415,c913,c3444,c1330,c2240,c118,c8102,c4403,c9283,c5354,c2165,c9428,c4143,c9340,c240,c1118,c3152,c6186,c4484,c972,c121,c2459,c4208,c3209,c4499,c379,c5259,c2157,c0321,c5145,c5311,c3147,c2207,c9131,c8285,c278,c5101,c1205,c682,c6188,c0159,c3255,c020,c6255,c6348,c774,c8372,c488,c4239,c7176,c244,c4174,c251,c397,c449,c861,c6309,c83,c0252,c5153,c7483,c5476,c4111,c2100,c7481,c3286,c815,c1277,c892,c4399,c1116,c135,c156,c6440,c8421,c4170,c657,c5421,c1461,c3109,c4322,c4388,c4421,c49,c0412,c0128,c0316,c523,c9452,c7206,c1387,c1177,c416,c9153,c1414,c4353,c9271,c2176,c991,c92,c5423,c1479,c9476,c8103,c382,c5349,c3183,c29,c9206,c1378,c8288,c6373,c85,c0205,c8374,c6266,c6396,c362,c1451,c2375,c5228,c5149,c8228,c1195,c8276,c351,c115,c8270,c380,c8492,c174,c477,c7205,c7135,c0389,c46,c1313,c9282,c084,c7407,c3499,c0450,c3341,c7386,c4443,c0147,c4234,c0158,c6245,c2173,c5366,c9398,c247,c0384,c3469,c0121,c8485,c8360,c0461,c3447,c829,c9378,c3379,c2217,c554,c4210,c2379,c1261,c8379,c9302,c5336,c8160,c0139,c331,c5116,c470,c6261,c6475,c634,c4444,c1450,c4103,c5132,c1139,c8106,c2427,c7431,c51,c7277,c273,c5210,c8179,c6325,c522,c0282,c9101,c7480,c8166,c9376,c2457,c3242,c981,c7364,c1314,c8234,c782,c142,c1315,c3334,c8308,c4351,c116,c512,c3456,c926,c3155,c9438,c3497,c6180,c045,c8152,c1312,c1310,c4228,c98,c9318,c1133,c6228,c6117,c7440,c1320,c7366,c6137,c9380,c5293,c5152,c0263,c8148,c5241,c191,c4192,c526,c7369,c2333,c5393,c3450,c9333,c7203,c4394,c6189,c495,c7276,c3352,c1262,c0213,c1425,c8290,c4113,c9461,c4284,c0262,c5249,c180,c1438,c90,c5346,c0497,c7417,c0202,c096,c327,c1176,c1141,c0330,c0445,c8473,c6260,c1210,c4146,c3143,c5144,c797,c0219,c335,c0154,c0107,c0314,c7103,c7383,c291,c0399,c6280,c6386,c3160,c86,c770,c6316,c2391,c8133,c1433,c9403,c4241,c1383,c6239,c8430,c3136,c9357,c827,c4203,c3290,c182,c8437,c0167,c5264,c0118,c5178,c954,c3389,c3275,c8226,c9187,c0357,c3273,c8241,c2202,c3300,c7397,c7210,c8188,c1405,c246,c3193,c4380,c480,c8476,c516,c8212,c4483,c451,c1148,c0299,c1256,c5215,c6360,c4381,c1355,c1302,c4491,c6378,c3158,c6413,c0261,c6125,c4109,c8440,c2330,c5231,c1100,c459,c2393,c9489,c9100,c1202,c6215,c4326,c9473,c9488,c5337,c9444,c0251,c9301,c1304,c6247,c4395,c0255,c8328,c3310,c9365,c2409,c0172,c2398,c2182,c3434,c3473,c8486,c1402,c113,c3363,c5147,c763,c26,c7332,c7111,c3279,c2395,c7476,c6476,c9189,c7123,c0486,c814,c4478,c6229,c3374,c533,c936,c4488,c9325,c179,c943,c5377,c4442,c4122,c8282,c1464,c3367,c6357,c0481,c7259,c5461,c4365,c6374,c1294,c7301,c5199,c0494,c7289,c9315,c852,c3280,c9328,c4223,c3118,c6465,c0152,c2279,c8443,c254,c4361,c1217,c3101,c7291,c3439,c157,c7472,c6263,c23,c3324,c3132,c1429,c425,c6289,c7119,c8304,c6170,c2416,c2144,c7166,c2148,c2280,c0228,c1259,c3397,c5374,c5428,c4355,c457,c9401,c7118,c0105,c6221,c0132,c3351,c1281,c1482,c0439,c3476,c3125,c232,c0180,c536,c4117,c5406,c3382,c5314,c2195,c3360,c8477,c4152,c793,c5462,c2287,c1290,c9257,c5289,c5104,c559,c8155,c0101,c0475,c360,c9334,c7473,c5437,c5121,c6418,c6167,c448,c8316,c616,c9117,c6484,c1123,c5473,c4349,c039,c60,c544,c9147,c3357,c042,c9217,c8377,c0243,c923,c6202,c3396,c4323,c5379,c8120,c2307,c466,c0278,c7254,c1417,c0187,c082,c5139,c8153,c928,c6112,c5170,c1362,c5362,c5243,c5312,c2106,c69,c5301,c0137,c3317,c8418,c4338,c3117,c3457,c7406,c3375,c9278,c952,c9478,c5383,c0270,c6417,c0138,c1147,c2265,c0222,c9260,c953,c8441,c1143,c6121,c1182,c1418,c8277,c7350,c2124,c1305,c8254,c0413,c09,c2281,c3246,c6407,c2372,c823,c1317,c3178,c236,c869,c293,c0414,c3182,c6128,c8143,c837,c5453,c2340,c6497,c9204,c9454,c0296,c6285,c0234,c3127,c1168,c8216,c2327,c9214,c8177,c5425,c4213,c428,c173,c7275,c9251,c6277,c162,c3284,c6244,c993,c1390,c1212,c6265,c8413,c4104,c4140,c5143,c931,c0319,c9129,c3189,c6303,c8164,c562,c8275,c740,c150,c5477,c3130,c0130,c061,c6420,c9316,c139,c4476,c8423,c652,c6145,c3150,c155,c517,c9177,c2220,c698,c2147,c4354,c1367,c1344,c6172,c4276,c5256,c7104,c8412,c878,c05,c0184,c9227,c0429,c4159,c2300,c6169,c0383,c7368,c5240,c811,c6106,c266,c087,c141,c4412,c8284,c7267,c4128,c6375,c0345,c9409,c558,c2271,c4267,c597,c9185,c1173,c945,c4236,c193,c374,c3421,c252,c6491,c7412,c8238,c8416,c272,c163,c5409,c070,c70,c816,c7128,c3308,c2488,c5490,c8244,c2411,c6425,c9368,c9436,c8147,c8132,c1191,c2341,c4132,c9492,c2166,c9360,c2129,c1470,c1249,c1377,c2320,c853,c7320,c858,c0423,c9191,c1242,c748,c9419,c5117,c7441,c6197,c8457,c3466,c7334,c7174,c2127,c3359,c5467,c3180,c490,c4485,c0349,c6288,c1478,c3170,c7442,c3176,c3498,c1309,c5221,c9197,c2481,c417,c4366,c5415,c1375,c546,c0492,c5297,c0360,c8279,c1272,c023,c621,c877,c066,c975,c2238,c7492,c997,c6185,c8332,c9256,c8182,c3215,c0436,c1352,c7261,c1332,c0237,c1267,c6432,c6198,c7154,c9399,c2276,c3320,c59,c5318,c7427,c3486,c65,c7168,c0165,c4127,c146,c0342,c79,c8163,c8415,c678,c5174,c8493,c186,c6196,c346,c5247,c4498,c9243,c1436,c2216,c4434,c6233,c527,c7130,c1101,c3265,c1499,c3271,c0390,c7252,c9337,c8218,c2406,c1265,c778,c7216,c3403,c3494,c0471,c9249,c4318,c941,c7404,c8366,c9139,c3393,c262,c3433,c6227,c5364,c1423,c1237,c626,c375,c0209,c4186,c7422,c899,c5246,c0343,c0374,c2370,c7475,c2400,c0488,c9460,c8439,c4489,c015,c2465,c5131,c9119,c2135,c4118,c4218,c3269,c9193,c6331,c3415,c5277,c5391,c1131,c8407,c4344,c6311,c2192,c7358,c1121,c9412,c1236,c3369,c1335,c017,c9170,c4172,c7474,c1495,c9388,c1412,c64,c5344,c3212,c0373,c2326,c994,c4263,c8405,c223,c4441,c5444,c7153,c9459,c3111,c6441,c9354,c99,c4481,c9472,c6123,c5164,c0441,c6144,c7413,c0432,c4242,c2383,c0232,c5169,c6403,c8198,c971,c2448,c4154,c890,c4178,c7370,c0333,c6447,c299,c411,c2107,c3411,c585,c377,c8488,c5176,c8256,c4459,c6211,c534,c4101,c8151,c0437,c2474,c5112,c4216,c6395,c9415,c5455,c0242,c8392,c5483,c2214,c2482,c4368,c3261,c6423,c7247,c2254,c0217,c249,c0153,c037,c4240,c7326,c1376,c2376,c3200,c5410,c9313,c6310,c733,c9414,c0326,c7336,c0368,c1336,c2334,c6323,c2250,c1104,c8224,c154,c7420,c783,c265,c7159,c8479,c5126,c4360,c259,c394,c7155,c2424,c6201,c0149,c2161,c8161,c3253,c0367,c7433,c2208,c7392,c3404,c6452,c8455,c8301,c6387,c9220,c21,c2385,c4271,c9225,c1445,c057,c9213,c412,c3419,c1130,c9352,c7470,c187,c5194,c0490,c6459,c8105,c129,c286,c1246,c2132,c8463,c1162,c0451,c8107,c9391,c25,c2415,c9289,c8438,c5498,c0109,c6114,c663,c8451,c1219,c833,c1427,c175,c011,c2258,c9159,c3312,c9140,c0129,c4138,c74,c4426,c8141,c2362,c849,c4405,c0419,c7186,c2291,c4119,c697,c924,c3378,c7449,c1110,c4370,c5250,c0207,c0272,c9143,c0328,c9400,c3203,c6270,c7443,c5229,c8335,c7185,c2196,c4131,c7235,c9137,c6372,c1189,c9221,c8299,c4108,c1333,c4144,c8122,c5482,c738,c5333,c219,c5485,c7114,c693,c0196,c1136,c0241,c3185,c9274,c1119,c0170,c5185,c7178,c6156,c0354,c695,c0186,c132,c168,c539,c4262,c3347,c0124,c5307,c9207,c7290,c5369,c3140,c1201,c445,c9125,c5405,c2452,c615,c9238,c729,c1160,c9200,c0418,c5291,c6494,c6267,c7138,c3451,c8136,c4169,c221,c410,c946,c880,c5175,c0221,c8313,c6204,c5279,c9418,c5151,c8128,c2237,c9284,c7158,c7122,c5138,c9253,c1393,c9270,c1472,c8207,c938,c0430,c8312,c9446,c00,c0267,c0322,c887,c5305,c4391,c9495,c1192,c239,c826,c944,c7499,c7164,c8433,c0420,c1397,c8280,c9362,c9427,c7152,c0433,c8195,c342,c7108,c856,c8467,c2445,c5135,c656,c5120,c7148,c7367,c2346,c489,c6222,c1486,c5200,c2446,c7362,c7222,c0362,c2283,c2104,c2109,c3377,c8367,c2447,c643,c0100,c8268,c073,c255,c333,c4467,c4397,c1366,c2312,c751,c1213,c7489,c3213,c8274,c4124,c1284,c2110,c8115,c2485,c8445,c5328,c9279,c5367,c9443,c4283,c4496,c028,c5285,c7373,c885,c935,c1494,c097,c4466,c9128,c6371,c9262,c787,c2336,c5426,c8419,c510,c5127,c9184,c0308,c5351,c8465,c0452,c5499,c2152,c910,c2105,c4492,c8170,c8499,c5308,c4400,c9486,c8300,c1253,c5298,c720,c4378,c6389,c511,c1245,c571,c5299,c96,c6321,c980,c7471,c1175,c5323,c2180,c7493,c7248,c238,c8157,c4436,c8447,c1382,c1138,c948,c750,c5324,c185,c8382,c1341,c158,c6401,c9155,c8324,c3338,c3301,c1188,c055,c1222,c5261,c985,c322,c292,c1426,c384,c7318,c383,c8145,c5317,c6377,c9146,c6376,c026,c5184,c2458,c5465,c566,c966,c785,c6343,c9467,c6333,c5234,c5266,c7278,c2295,c3274,c0131,c3230,c8460,c1439,c1324,c9484,c9111,c5219,c7181,c0226,c120,c1407,c587,c5114,c398,c9248,c053,c2470,c934,c0294,c2302,c1120,c4468,c4270,c3204,c6276,c2408,c436,c1289,c9382,c074,c4287,c1442,c0181,c649,c9273,c6148,c696,c6295,c3120,c3340,c9265,c963,c821,c3395,c7324,c4280,c320,c4195,c022,c2310,c04,c2469,c691,c3190,c9173,c0340,c2206,c7353,c735,c3154,c5454,c567,c9171,c9317,c190,c3427,c1374,c077,c1154,c3133,c24,c2149,c6499,c2428,c7137,c588,c7363,c0119,c138,c8269,c9157,c1386,c430,c5198,c6262,c6399,c922,c3131,c742,c1156,c8320,c4424,c1392,c3385,c8371,c0148,c8431,c7411,c4211,c5430,c6496,c1171,c3491,c4220,c4343,c0260,c334,c8201,c4336,c719,c5161,c5157,c8140,c7228,c8450,c3151,c1443,c7381,c3314,c7328,c5419,c8309,c6217,c5288,c3429,c1474,c0364,c5373,c3258,c088,c9377,c8111,c5329,c4453,c8302,c50,c044,c456,c0208,c4450,c7376,c2227,c6308,c7327,c5450,c9231,c231,c2471,c8291,c7161,c9389,c2177,c1137,c4386,c561,c5411,c3142,c3425,c8426,c0248,c4438,c6424,c7146,c6486,c0386,c767,c0320,c2380,c0426,c4187,c9416,c6446,c2118,c184,c9295,c1322,c3468,c4185,c6414,c0271,c9367,c2410,c3481,c694,c9493,c2492,c9232,c1413,c0239,c7429,c8171,c8129,c2443,c3325,c2364,c095,c271,c6162,c2117,c3163,c8378,c294,c549,c6437,c8489,c9205,c9287,c7183,c0200,c365,c8261,c3146,c3277,c358,c8185,c9483,c6143,c8496,c8227,c8232,c1358,c5306,c6468,c2290,c927,c2187,c2244,c8344,c4215,c715,c4134,c737,c9393,c0286,c683,c2278,c9406,c40,c6364,c4337,c4420,c2390,c6126,c0230,c651,c0178,c6462,c886,c7116,c2160,c7109,c4409,c8174,c7215,c3196,c9392,c7408,c0406,c872,c4440,c4446,c642,c9264,c2354,c9372,c9373,c7359,c1208,c0183,c5418,c133,c659,c1185,c0162,c5107,c5100,c4445,c0446,c7145,c4256,c464,c8204,c0289,c8381,c8193,c9133,c5287,c6324,c3426,c9258,c5310,c537,c0268,c1125,c3344,c3227,c2371,c378,c1163,c2249,c176,c5422,c8495,c1144,c6290,c97,c8454,c2205,c2454,c685,c0477,c7202,c4406,c0470,c5448,c3137,c0353,c918,c7460,c960,c4306,c7308,c4255,c1132,c8354,c9158,c9411,c81,c4244,c875,c6302,c4277,c39,c1308,c7435,c5155,c5204,c8414,c87,c9148,c9466,c8406,c3256,c310,c476,c336,c5416,c1194,c8334,c345,c6301,c5340,c5162,c0458,c8239,c7341,c0351,c681,c4121,c5492,c065,c415,c2120,c2344,c568,c832,c2222,c7315,c7121,c9336,c6274,c145,c7360,c6200,c3186,c4268,c8395,c8387,c968,c739,c5396,c6366,c3482,c253,c5356,c5273,c7377,c0410,c2357,c1303,c2477,c3278,c1149,c2143,c5196,c5274,c666,c0108,c6429,c6332,c7398,c8356,c6133,c2142,c1151,c9269,c8402,c3348,c5209,c3168,c7432,c4227,c5187,c5365,c6346,c3281,c01,c677,c939,c598,c5322,c6238,c4455,c4175,c3370,c2230,c2103,c0279,c6205,c9404,c5167,c421,c1251,c867,c067,c1435,c2141,c4200,c1112,c995,c6158,c2440,c8231,c8134,c035,c6257,c3394,c648,c6235,c66,c9161,c6336,c243,c4142,c9410,c0292,c820,c4345,c6318,c0473,c0155,c3373,c5360,c625,c9375,c6402,c047,c461,c2282,c1161,c747,c050,c092,c0493,c329,c0318,c3318,c2294,c313,c3145,c514,c3335,c7299,c1493,c8429,c0358,c2437,c8199,c4149,c7256,c7331,c596,c1476,c4161,c9435,c3398,c9152,c4422,c7191,c1359,c3328,c2319,c8384,c2221,c67,c5327,c7335,c1199,c8265,c3172,c9254,c7177,c4379,c830,c6199,c4302,c3358,c7272,c6406,c8139,c3296,c5487,c164,c474,c2356,c7241,c3222,c957,c2136,c0424,c8233,c1356,c1369,c234,c4427,c3202,c3129,c016,c062,c9235,c7385,c4314,c687,c1187,c7380,c4382,c3366,c41,c6212,c2418,c627,c4148,c5394,c2345,c7452,c442,c3289,c8323,c2449,c8393,c2256,c2342,c5108,c064,c7229,c6138,c6478,c6307,c6421,c586,c1126,c721,c3197,c460,c8370,c126,c210,c5271,c9361,c6479,c1146,c3420,c0355,c4342,c8255,c276,c3126,c274,c9230,c868,c1122,c4392,c5158,c52,c2200,c1477,c02,c6319,c7296,c7306,c6273,c1496,c0298,c3474,c4369,c229,c8172,c091,c8173,c6492,c7208,c3416,c3449,c9224,c4126,c9245,c6237,c4297,c5392,c6213,c0177,c2303,c4362,c9341,c58,c0379,c1117,c3249,c3162,c2134,c1444,c6283,c5431,c1440,c594,c5276,c486,c595,c9195,c385,c38,c632,c5192,c6147,c4191,c6379,c1421,c3239,c5463,c756,c9324,c2133,c5230,c4249,c667,c6160,c2219,c0134,c0307,c6173,c2137,c4359,c8340,c5459,c1285,c9124,c8283,c5292,c831,c8434,c3479,c1105,c9463,c9218,c147,c9168,c455,c4482,c8138,c0210,c3225,c014,c3372,c399,c1447,c242,c9113,c5358,c5283,c0288,c3323,c197,c433,c5290,c20,c277,c2189,c2377,c8180,c9293,c8346,c1399,c4309,c1273,c1395,c7423,c2420,c5493,c5480,c714,c1258,c920,c9470,c5159,c2268,c5352,c5257,c8266,c8189,c153,c5102,c2139,c119,c578,c0283,c727,c4182,c9338,c513,c5497,c1485,c7314,c2234,c5348,c3471,c7157,c949,c9349,c1410,c2435,c6176,c432,c4396,c5262,c8481,c9166,c879,c8350,c53,c1321,c1103,c7136,c1165,c8159,c32,c986,c4407,c7282,c3349,c5385,c7300,c4316,c7338,c3458,c8442,c7171,c8428,c7424,c3124,c661,c2273,c8452,c5265,c6455,c0106,c361,c4105,c2119,c1230,c4320,c9219,c7175,c1347,c290,c5254,c5160,c882,c1497,c3108,c6190,c5468,c4357,c4229,c2493,c7265,c454,c7382,c776,c4289,c5281,c8217,c9112,c2389,c8246,c6456,c9190,c0378,c4163,c4198,c4275,c4253,c3467,c224,c5447,c1264,c1102,c6464,c8260,c7461,c732,c2351,c618,c5458,c1172,c9174,c3418,c3399,c0216,c013,c6340,c5332,c4423,c540,c7396,c5300,c9394,c1206,c9448,c2296,c6102,c1449,c319,c0480,c485,c8494,c5464,c8326,c3191,c438,c0489,c761,c0171,c929,c1370,c7240,c441,c9103,c1471,c6254,c4376,c893,c260,c726,c4238,c1404,c686,c144,c611,c0363,c0111,c7163,c9429,c8311,c4261,c0375,c5244,c357,c3157,c5125,c9307,c44,c2293,c7173,c8287,c3107,c3115,c660,c7428,c624,c0168,c6253,c0204,c283,c1368,c5420,c1484,c9327,c2422,c7448,c8124,c3445,c7419,c8165,c9491,c6460,c481,c9294,c7486,c051,c3315,c9387,c9469,c6466,c484,c389,c0444,c225,c5475,c5489,c0485,c9458,c151,c7179,c3432,c370,c6351,c897,c8263,c1379,c564,c5251,c5148,c6400,c4252,c0211,c3413,c214,c235,c0233,c8210,c1227,c4311,c7284,c1430,c5456,c741,c4251,c330,c2116,c860,c6362,c029,c352,c8398,c127,c363,c6115,c0102,c7339,c3201,c8315,c9498,c368,c1179,c4199,c344,c2309,c7451,c1351,c5407,c3472,c0224,c9188,c124,c1250,c393,c7317,c1260,c5399,c148,c2382,c7238,c8213,c2399,c7438,c3105,c9240,c5343,c9208,c6225,c6487,c6474,c7281,c0332,c2286,c220,c1357,c0194,c2305,c1422,c8391,c1323,c8205,c8361,c6433,c5325,c1319,c6177,c8158,c6157,c6109,c297,c5213,c771,c9487,c8219,c1408,c4184,c8214,c854,c281,c217,c670,c328,c043,c2168,c424,c2387,c1107,c4465,c5232,c5225,c178,c3493,c9423,c638,c9425,c0431,c183,c5154,c2113,c269,c8364,c6251,c437,c6152,c2324,c390,c4133,c7107,c9445,c3224,c9482,c0377,c9383,c6165,c3250,c2405,c4477,c5438,c4171,c55,c0422,c9479,c9413,c1424,c5320,c3167,c4264,c4471,c2456,c6344,c9246,c6256,c7251,c7391,c8142,c7232,c1170,c35,c8383,c230,c2125,c6472,c2335,c6385,c12,c7237,c325,c6135,c9228,c1361,c9457,c1218,c6457,c2266,c5466,c579,c8150,c4463,c1325,c0499,c799,c8458,c0347,c2213,c542,c999,c6279,c2489,c465,c372,c7192,c7263,c654,c3291,c535,c631,c2378,c3179,c282,c7249,c0169,c0372,c256,c8119,c5111,c6175,c2497,c1293,c4254,c6203,c2463,c2347,c4201,c8272,c9154,c3475,c8303,c80,c326,c3412,c9118,c0193,c4458,c1157,c940,c7302,c851,c318,c7309,c343,c7167,c4347,c1233,c1295,c4462,c8126,c8293,c1292,c5195,c584,c4296,c6234,c5386,c8149,c4324,c1215,c8425,c2413,c5103,c9355,c048,c337,c7188,c8220,c4167,c6392,c4155,c5397,c8409,c5235,c6150,c5395,c1337,c7156,c3495,c6410,c4384,c0104,c2421,c4479,c8349,c8196,c5278,c0469,c9397,c7322,c2478,c4469,c2170,c3437,c2153,c3496,c8375,c6335,c6315,c9127,c5414,c996,c781,c0190,c9106,c7401,c0359,c2245,c4248,c4299,c672,c6194,c6120,c227,c1307,c4451,c9280,c3442,c3217,c027,c2325,c723,c5227,c6337,c3223,c845,c4115,c2264,c4332,c3237,c0247,c1226,c6104,c9468,c550,c5429,c054,c7129,c4464,c6415,c192,c010,c388,c9215,c159,c7463,c5331,c2374,c9239,c419,c267,c032,c4448,c4497,c0146,c0291,c038,c0305,c9259,c9496,c3206,c664,c8368,c0395,c10,c3311,c7170,c3487,c688,c6284,c0346,c8369,c2131,c6191,c1365,c2285,c2316,c216,c6342,c9421,c2284,c7394,c499,c4180,c0464,c0273,c2337,c08,c270,c2253,c2158,c4207,c8348,c2209,c3208,c5295,c0150,c3316,c4181,c11,c7482,c988,c0179,c2407,c332,c6404,c4305,c8482,c6453,c7379,c898,c870,c5355,c1115,c5387,c0443,c3295,c0197,c7437,c2130,c3134,c0203,c6398,c6300,c9150,c0411,c2323,c2257,c1158,c2140,c7354,c472,c7262,c7260,c2272,c3100,c9351,c9431,c3406,c57,c7243,c0301,c8358,c6149,c8117,c6164,c1184,c3440,c7144,c758,c7497,c978,c580,c7293,c8408,c314,c2167,c9437,c4165,c3346,c4303,c4294,c7189,c8339,c1198,c680,c9480,c0336,c228,c6393,c0290,c2373,c463,c369,c7268,c8100,c4278,c9202,c6448,c630,c9272,c8417,c1169,c2451,c3302,c9424,c3388,c541,c847,c4156,c565,c2365,c4350,c9339,c386,c646,c8249,c2350,c874,c8209,c3123,c6329,c19,c4274,c4188,c5267,c2191,c1409,c6471,c1354,c7199,c9312,c6405,c3309,c1278,c198,c5496,c4123,c9439,c0225,c6354,c0238,c958,c5253,c2232,c1434,c27,c1266,c355,c7312,c5440,c9420,c30,c5472,c919,c3430,c8380,c2480,c0166,c6358,c6193,c1288,c716,c1135,c3293,c6481,c5207,c3292,c6226,c5330,c7405,c7313,c5313,c5481,c0361,c1458,c2226,c5206,c123,c4310,c581,c8424,c311,c3161,c1331,c222,c2212,c4457,c058,c1297,c2171,c8461,c2388,c2231,c7212,c8137,c0380,c528,c4258 );

input x0;
input x1;
input x2;
input x3;
input x4;
input x5;
input x6;
input x7;
input x8;
input x9;
input x10;
input x11;
input x12;
input x13;
input x14;
input x15;
input x16;
input x17;
input x18;
input x19;
input x20;
input x21;
input x22;
input x23;
input x24;
input x25;
input x26;
input x27;
input x28;
input x29;
input x30;
input x31;
input x32;
input x33;
input x34;
input x35;
input x36;
input x37;
input x38;
input x39;
input x40;
input x41;
input x42;
input x43;
input x44;
input x45;
input x46;
input x47;
input x48;
input x49;
input x50;
input x51;
input x52;
input x53;
input x54;
input x55;
input x56;
input x57;
input x58;
input x59;
input x60;
input x61;
input x62;
input x63;
input x64;
input x65;
input x66;
input x67;
input x68;
input x69;
input x70;
input x71;
input x72;
input x73;
input x74;
input x75;
input x76;
input x77;
input x78;
input x79;
input x80;
input x81;
input x82;
input x83;
input x84;
input x85;
input x86;
input x87;
input x88;
input x89;
input x90;
input x91;
input x92;
input x93;
input x94;
input x95;
input x96;
input x97;
input x98;
input x99;
input x100;
input x101;
input x102;
input x103;
input x104;
input x105;
input x106;
input x107;
input x108;
input x109;
input x110;
input x111;
input x112;
input x113;
input x114;
input x115;
input x116;
input x117;
input x118;
input x119;
input x120;
input x121;
input x122;
input x123;
input x124;
input x125;
input x126;
input x127;
input x128;
input x129;
input x130;
input x131;
input x132;
input x133;
input x134;
input x135;
input x136;
input x137;
input x138;
input x139;
input x140;
input x141;
input x142;
input x143;
input x144;
input x145;
input x146;
input x147;
input x148;
input x149;
input x150;
input x151;
input x152;
input x153;
input x154;
input x155;
input x156;
input x157;
input x158;
input x159;
input x160;
input x161;
input x162;
input x163;
input x164;
input x165;
input x166;
input x167;
input x168;
input x169;
input x170;
input x171;
input x172;
input x173;
input x174;
input x175;
input x176;
input x177;
input x178;
input x179;
input x180;
input x181;
input x182;
input x183;
input x184;
input x185;
input x186;
input x187;
input x188;
input x189;
input x190;
input x191;
input x192;
input x193;
input x194;
input x195;
input x196;
input x197;
input x198;
input x199;
input x200;
input x201;
input x202;
input x203;
input x204;
input x205;
input x206;
input x207;
input x208;
input x209;
input x210;
input x211;
input x212;
input x213;
input x214;
input x215;
input x216;
input x217;
input x218;
input x219;
input x220;
input x221;
input x222;
input x223;
input x224;
input x225;
input x226;
input x227;
input x228;
input x229;
input x230;
input x231;
input x232;
input x233;
input x234;
input x235;
input x236;
input x237;
input x238;
input x239;
input x240;
input x241;
input x242;
input x243;
input x244;
input x245;
input x246;
input x247;
input x248;
input x249;
input x250;
input x251;
input x252;
input x253;
input x254;
input x255;
input x256;
input x257;
input x258;
input x259;
input x260;
input x261;
input x262;
input x263;
input x264;
input x265;
input x266;
input x267;
input x268;
input x269;
input x270;
input x271;
input x272;
input x273;
input x274;
input x275;
input x276;
input x277;
input x278;
input x279;
input x280;
input x281;
input x282;
input x283;
input x284;
input x285;
input x286;
input x287;
input x288;
input x289;
input x290;
input x291;
input x292;
input x293;
input x294;
input x295;
input x296;
input x297;
input x298;
input x299;
input x300;
input x301;
input x302;
input x303;
input x304;
input x305;
input x306;
input x307;
input x308;
input x309;
input x310;
input x311;
input x312;
input x313;
input x314;
input x315;
input x316;
input x317;
input x318;
input x319;
input x320;
input x321;
input x322;
input x323;
input x324;
input x325;
input x326;
input x327;
input x328;
input x329;
input x330;
input x331;
input x332;
input x333;
input x334;
input x335;
input x336;
input x337;
input x338;
input x339;
input x340;
input x341;
input x342;
input x343;
input x344;
input x345;
input x346;
input x347;
input x348;
input x349;
input x350;
input x351;
input x352;
input x353;
input x354;
input x355;
input x356;
input x357;
input x358;
input x359;
input x360;
input x361;
input x362;
input x363;
input x364;
input x365;
input x366;
input x367;
input x368;
input x369;
input x370;
input x371;
input x372;
input x373;
input x374;
input x375;
input x376;
input x377;
input x378;
input x379;
input x380;
input x381;
input x382;
input x383;
input x384;
input x385;
input x386;
input x387;
input x388;
input x389;
input x390;
input x391;
input x392;
input x393;
input x394;
input x395;
input x396;
input x397;
input x398;
input x399;
input x400;
input x401;
input x402;
input x403;
input x404;
input x405;
input x406;
input x407;
input x408;
input x409;
input x410;
input x411;
input x412;
input x413;
input x414;
input x415;
input x416;
input x417;
input x418;
input x419;
input x420;
input x421;
input x422;
input x423;
input x424;
input x425;
input x426;
input x427;
input x428;
input x429;
input x430;
input x431;
input x432;
input x433;
input x434;
input x435;
input x436;
input x437;
input x438;
input x439;
input x440;
input x441;
input x442;
input x443;
input x444;
input x445;
input x446;
input x447;
input x448;
input x449;
input x450;
input x451;
input x452;
input x453;
input x454;
input x455;
input x456;
input x457;
input x458;
input x459;
input x460;
input x461;
input x462;
input x463;
input x464;
input x465;
input x466;
input x467;
input x468;
input x469;
input x470;
input x471;
input x472;
input x473;
input x474;
input x475;
input x476;
input x477;
input x478;
input x479;
input x480;
input x481;
input x482;
input x483;
input x484;
input x485;
input x486;
input x487;
input x488;
input x489;
input x490;
input x491;
input x492;
input x493;
input x494;
input x495;
input x496;
input x497;
input x498;
input x499;
input x500;
input x501;
input x502;
input x503;
input x504;
input x505;
input x506;
input x507;
input x508;
input x509;
input x510;
input x511;
input x512;
input x513;
input x514;
input x515;
input x516;
input x517;
input x518;
input x519;
input x520;
input x521;
input x522;
input x523;
input x524;
input x525;
input x526;
input x527;
input x528;
input x529;
input x530;
input x531;
input x532;
input x533;
input x534;
input x535;
input x536;
input x537;
input x538;
input x539;
input x540;
input x541;
input x542;
input x543;
input x544;
input x545;
input x546;
input x547;
input x548;
input x549;
input x550;
input x551;
input x552;
input x553;
input x554;
input x555;
input x556;
input x557;
input x558;
input x559;
input x560;
input x561;
input x562;
input x563;
input x564;
input x565;
input x566;
input x567;
input x568;
input x569;
input x570;
input x571;
input x572;
input x573;
input x574;
input x575;
input x576;
input x577;
input x578;
input x579;
input x580;
input x581;
input x582;
input x583;
input x584;
input x585;
input x586;
input x587;
input x588;
input x589;
input x590;
input x591;
input x592;
input x593;
input x594;
input x595;
input x596;
input x597;
input x598;
input x599;
input x600;
input x601;
input x602;
input x603;
input x604;
input x605;
input x606;
input x607;
input x608;
input x609;
input x610;
input x611;
input x612;
input x613;
input x614;
input x615;
input x616;
input x617;
input x618;
input x619;
input x620;
input x621;
input x622;
input x623;
input x624;
input x625;
input x626;
input x627;
input x628;
input x629;
input x630;
input x631;
input x632;
input x633;
input x634;
input x635;
input x636;
input x637;
input x638;
input x639;
input x640;
input x641;
input x642;
input x643;
input x644;
input x645;
input x646;
input x647;
input x648;
input x649;
input x650;
input x651;
input x652;
input x653;
input x654;
input x655;
input x656;
input x657;
input x658;
input x659;
input x660;
input x661;
input x662;
input x663;
input x664;
input x665;
input x666;
input x667;
input x668;
input x669;
input x670;
input x671;
input x672;
input x673;
input x674;
input x675;
input x676;
input x677;
input x678;
input x679;
input x680;
input x681;
input x682;
input x683;
input x684;
input x685;
input x686;
input x687;
input x688;
input x689;
input x690;
input x691;
input x692;
input x693;
input x694;
input x695;
input x696;
input x697;
input x698;
input x699;
input x700;
input x701;
input x702;
input x703;
input x704;
input x705;
input x706;
input x707;
input x708;
input x709;
input x710;
input x711;
input x712;
input x713;
input x714;
input x715;
input x716;
input x717;
input x718;
input x719;
input x720;
input x721;
input x722;
input x723;
input x724;
input x725;
input x726;
input x727;
input x728;
input x729;
input x730;
input x731;
input x732;
input x733;
input x734;
input x735;
input x736;
input x737;
input x738;
input x739;
input x740;
input x741;
input x742;
input x743;
input x744;
input x745;
input x746;
input x747;
input x748;
input x749;
input x750;
input x751;
input x752;
input x753;
input x754;
input x755;
input x756;
input x757;
input x758;
input x759;
input x760;
input x761;
input x762;
input x763;
input x764;
input x765;
input x766;
input x767;
input x768;
input x769;
input x770;
input x771;
input x772;
input x773;
input x774;
input x775;
input x776;
input x777;
input x778;
input x779;
input x780;
input x781;
input x782;
input x783;
output c3401;
output c1490;
output c5398;
output c7286;
output c439;
output c8240;
output c947;
output c4206;
output c2455;
output c152;
output c9300;
output c1113;
output c079;
output c3229;
output c8483;
output c969;
output c0269;
output c0366;
output c3285;
output c2162;
output c196;
output c3187;
output c8271;
output c136;
output c8471;
output c3480;
output c0371;
output c8104;
output c8242;
output c4330;
output c679;
output c6498;
output c5202;
output c5341;
output c473;
output c7454;
output c950;
output c6430;
output c6416;
output c6252;
output c298;
output c2366;
output c6422;
output c7102;
output c6294;
output c613;
output c753;
output c866;
output c0120;
output c8491;
output c7231;
output c195;
output c0334;
output c215;
output c1200;
output c2224;
output c54;
output c6353;
output c736;
output c7330;
output c1346;
output c4456;
output c8252;
output c3264;
output c137;
output c5319;
output c9241;
output c5363;
output c134;
output c6370;
output c7457;
output c4226;
output c5272;
output c7333;
output c8453;
output c1318;
output c371;
output c4183;
output c2298;
output c9210;
output c3391;
output c9196;
output c5484;
output c5451;
output c6327;
output c1498;
output c0381;
output c0415;
output c5339;
output c8468;
output c4460;
output c1411;
output c4110;
output c6113;
output c2313;
output c0324;
output c4348;
output c7345;
output c9322;
output c2426;
output c673;
output c9408;
output c4319;
output c4358;
output c9244;
output c3235;
output c4401;
output c531;
output c9165;
output c2367;
output c1465;
output c3299;
output c31;
output c6130;
output c3462;
output c773;
output c034;
output c8345;
output c5335;
output c7250;
output c7147;
output c8322;
output c2260;
output c4259;
output c2241;
output c395;
output c644;
output c1342;
output c8108;
output c6271;
output c5478;
output c619;
output c7285;
output c3303;
output c5224;
output c6278;
output c1316;
output c990;
output c3288;
output c6232;
output c479;
output c2218;
output c0491;
output c725;
output c6166;
output c6427;
output c4293;
output c1388;
output c6381;
output c970;
output c1353;
output c4222;
output c8245;
output c9329;
output c2108;
output c4404;
output c7464;
output c9164;
output c7271;
output c713;
output c1299;
output c4162;
output c7200;
output c5216;
output c5197;
output c8297;
output c3322;
output c9104;
output c284;
output c7223;
output c6142;
output c8109;
output c5294;
output c15;
output c655;
output c6339;
output c1275;
output c241;
output c636;
output c6249;
output c1420;
output c5191;
output c855;
output c1432;
output c7221;
output c1234;
output c3387;
output c676;
output c8436;
output c3461;
output c7213;
output c563;
output c1327;
output c3298;
output c5220;
output c4363;
output c2429;
output c1231;
output c3376;
output c3177;
output c8118;
output c3381;
output c6291;
output c211;
output c8329;
output c3443;
output c1466;
output c3331;
output c6434;
output c7182;
output c589;
output c7280;
output c3478;
output c7365;
output c6272;
output c364;
output c4291;
output c2267;
output c3195;
output c1469;
output c3252;
output c7337;
output c818;
output c3199;
output c0463;
output c0455;
output c917;
output c2114;
output c0123;
output c6264;
output c3435;
output c7245;
output c75;
output c9381;
output c3441;
output c4158;
output c1373;
output c7311;
output c0449;
output c3188;
output c7485;
output c1291;
output c6101;
output c1247;
output c3368;
output c6388;
output c2436;
output c2169;
output c143;
output c5252;
output c0487;
output c0256;
output c6236;
output c0435;
output c1340;
output c3448;
output c4414;
output c865;
output c8192;
output c6103;
output c3231;
output c7488;
output c2486;
output c3428;
output c3207;
output c6305;
output c233;
output c487;
output c8190;
output c0157;
output c9222;
output c9268;
output c8200;
output c3330;
output c0335;
output c6350;
output c5177;
output c2179;
output c5218;
output c3297;
output c2184;
output c3383;
output c7355;
output c0175;
output c5413;
output c1328;
output c5338;
output c5133;
output c992;
output c728;
output c0474;
output c89;
output c0447;
output c653;
output c7346;
output c711;
output c263;
output c914;
output c166;
output c7321;
output c7323;
output c7297;
output c7387;
output c8390;
output c9110;
output c942;
output c8466;
output c1106;
output c9371;
output c4114;
output c4221;
output c2322;
output c7450;
output c794;
output c0212;
output c4224;
output c553;
output c2269;
output c341;
output c8400;
output c2402;
output c3247;
output c0244;
output c4235;
output c76;
output c4495;
output c7113;
output c4230;
output c06;
output c8432;
output c9434;
output c9145;
output c7414;
output c161;
output c8125;
output c0254;
output c6100;
output c420;
output c7371;
output c8480;
output c640;
output c1268;
output c4428;
output c576;
output c6359;
output c458;
output c2462;
output c090;
output c3116;
output c5105;
output c690;
output c9308;
output c5258;
output c545;
output c0227;
output c462;
output c9201;
output c3417;
output c710;
output c443;
output c6231;
output c7139;
output c5350;
output c261;
output c1225;
output c0482;
output c5163;
output c9203;
output c3390;
output c2473;
output c6431;
output c789;
output c5382;
output c1241;
output c3260;
output c391;
output c0468;
output c081;
output c9160;
output c0428;
output c0265;
output c712;
output c5183;
output c8404;
output c2188;
output c6445;
output c2432;
output c859;
output c5389;
output c6367;
output c6243;
output c0287;
output c7194;
output c7195;
output c0398;
output c8127;
output c4246;
output c3342;
output c8235;
output c7201;
output c8144;
output c471;
output c3216;
output c6451;
output c556;
output c3238;
output c33;
output c2453;
output c0427;
output c2122;
output c9292;
output c8310;
output c5136;
output c0483;
output c8318;
output c7209;
output c933;
output c839;
output c862;
output c3282;
output c8462;
output c8237;
output c8317;
output c1453;
output c8267;
output c5275;
output c3453;
output c7149;
output c1159;
output c951;
output c6380;
output c3174;
output c2444;
output c3254;
output c6450;
output c2472;
output c9162;
output c8444;
output c8472;
output c7219;
output c8306;
output c3436;
output c3464;
output c1240;
output c2150;
output c6493;
output c4487;
output c3361;
output c4269;
output c6241;
output c4125;
output c8319;
output c9426;
output c287;
output c5357;
output c0253;
output c5390;
output c8187;
output c9346;
output c7421;
output c6134;
output c1473;
output c2204;
output c8386;
output c8259;
output c1398;
output c9126;
output c0306;
output c863;
output c1155;
output c6334;
output c237;
output c071;
output c62;
output c749;
output c7172;
output c7352;
output c431;
output c7498;
output c5140;
output c5443;
output c1153;
output c083;
output c040;
output c218;
output c9141;
output c7494;
output c5376;
output c0350;
output c5381;
output c9149;
output c0125;
output c6242;
output c2126;
output c3477;
output c4225;
output c7409;
output c2239;
output c0281;
output c8223;
output c1127;
output c6171;
output c4204;
output c8403;
output c1248;
output c1441;
output c212;
output c8183;
output c9199;
output c7295;
output c6131;
output c8156;
output c0189;
output c1306;
output c2450;
output c0264;
output c7165;
output c5166;
output c3371;
output c258;
output c5142;
output c1363;
output c9475;
output c6330;
output c4313;
output c91;
output c987;
output c6382;
output c3408;
output c8478;
output c9343;
output c850;
output c4106;
output c7445;
output c5474;
output c4413;
output c498;
output c6110;
output c7410;
output c4470;
output c7325;
output c1492;
output c068;
output c9299;
output c188;
output c025;
output c6136;
output c551;
output c7395;
output c1108;
output c423;
output c788;
output c3313;
output c2198;
output c8191;
output c9198;
output c8464;
output c9236;
output c61;
output c0387;
output c4100;
output c4177;
output c4129;
output c5115;
output c3122;
output c8388;
output c5119;
output c699;
output c5269;
output c482;
output c3409;
output c812;
output c3220;
output c9447;
output c784;
output c7444;
output c5471;
output c9364;
output c8314;
output c2401;
output c5238;
output c340;
output c3319;
output c9115;
output c1220;
output c6296;
output c0144;
output c0198;
output c1481;
output c2306;
output c2483;
output c0365;
output c9266;
output c8338;
output c0156;
output c2297;
output c4433;
output c9209;
output c046;
output c5212;
output c6155;
output c2248;
output c6220;
output c6146;
output c6317;
output c3492;
output c493;
output c573;
output c717;
output c2255;
output c9250;
output c076;
output c0304;
output c5372;
output c1372;
output c2328;
output c7456;
output c766;
output c0229;
output c5486;
output c4190;
output c0394;
output c9390;
output c8307;
output c5404;
output c1415;
output c0258;
output c4327;
output c8331;
output c348;
output c7292;
output c5309;
output c8206;
output c3159;
output c6248;
output c9180;
output c250;
output c6208;
output c3402;
output c7356;
output c339;
output c2112;
output c6384;
output c4290;
output c0214;
output c3283;
output c7117;
output c3400;
output c8397;
output c9288;
output c5113;
output c4402;
output c7307;
output c3148;
output c777;
output c6428;
output c7400;
output c1167;
output c0297;
output c623;
output c012;
output c2499;
output c9175;
output c3339;
output c6436;
output c7234;
output c321;
output c6293;
output c4390;
output c5491;
output c0465;
output c7279;
output c3194;
output c2156;
output c2430;
output c5282;
output c5380;
output c6214;
output c0312;
output c543;
output c0112;
output c396;
output c894;
output c3175;
output c4335;
output c9430;
output c8167;
output c5375;
output c0280;
output c021;
output c483;
output c0457;
output c6304;
output c1228;
output c7112;
output c5316;
output c6153;
output c6132;
output c0382;
output c199;
output c0385;
output c7125;
output c1475;
output c9176;
output c4176;
output c7141;
output c7226;
output c9304;
output c4196;
output c5345;
output c8325;
output c518;
output c1180;
output c2181;
output c8333;
output c6139;
output c5203;
output c650;
output c4112;
output c4325;
output c3263;
output c8258;
output c8262;
output c964;
output c9453;
output c1381;
output c7393;
output c9135;
output c3259;
output c4217;
output c189;
output c7495;
output c2186;
output c4374;
output c5296;
output c0400;
output c4130;
output c7187;
output c3241;
output c6473;
output c8399;
output c5280;
output c110;
output c1209;
output c635;
output c519;
output c5233;
output c6412;
output c1134;
output c612;
output c9310;
output c4286;
output c3485;
output c7374;
output c828;
output c2484;
output c4160;
output c3350;
output c617;
output c3149;
output c3218;
output c4298;
output c7466;
output c8121;
output c0218;
output c117;
output c289;
output c6140;
output c0126;
output c056;
output c3192;
output c3294;
output c2403;
output c4408;
output c674;
output c2476;
output c6224;
output c5353;
output c989;
output c3336;
output c4480;
output c4145;
output c5435;
output c0476;
output c7242;
output c547;
output c5368;
output c4139;
output c2318;
output c8215;
output c1238;
output c9182;
output c844;
output c4107;
output c4279;
output c1164;
output c194;
output c746;
output c8286;
output c7217;
output c3173;
output c3483;
output c0338;
output c891;
output c0127;
output c5449;
output c2394;
output c4387;
output c583;
output c1128;
output c834;
output c172;
output c2138;
output c760;
output c4321;
output c2201;
output c669;
output c4435;
output c4189;
output c0456;
output c4416;
output c0442;
output c6477;
output c3333;
output c835;
output c6141;
output c5208;
output c359;
output c5124;
output c610;
output c6483;
output c6230;
output c1282;
output c71;
output c525;
output c2203;
output c0135;
output c7150;
output c82;
output c848;
output c0110;
output c169;
output c1197;
output c7294;
output c9465;
output c4429;
output c4334;
output c0376;
output c8236;
output c447;
output c5165;
output c3459;
output c6240;
output c452;
output c2101;
output c3106;
output c9163;
output c0215;
output c5242;
output c125;
output c63;
output c765;
output c0163;
output c4193;
output c414;
output c4243;
output c114;
output c974;
output c4205;
output c3234;
output c22;
output c7233;
output c0369;
output c3410;
output c9116;
output c2194;
output c0409;
output c3332;
output c3171;
output c4257;
output c7246;
output c2358;
output c6297;
output c979;
output c3165;
output c3343;
output c4339;
output c7127;
output c0174;
output c572;
output c2331;
output c3181;
output c790;
output c8363;
output c575;
output c593;
output c0329;
output c366;
output c570;
output c4281;
output c6426;
output c1468;
output c4137;
output c167;
output c0310;
output c4120;
output c9237;
output c822;
output c0496;
output c080;
output c6184;
output c181;
output c3245;
output c5193;
output c6341;
output c7434;
output c825;
output c5460;
output c7403;
output c9290;
output c316;
output c6108;
output c5226;
output c4273;
output c6250;
output c9332;
output c956;
output c1349;
output c450;
output c171;
output c779;
output c6210;
output c1196;
output c976;
output c28;
output c8327;
output c982;
output c840;
output c0300;
output c1311;
output c6383;
output c7303;
output c2123;
output c5109;
output c7220;
output c6443;
output c3164;
output c7426;
output c2339;
output c5239;
output c3112;
output c1345;
output c1283;
output c5446;
output c7310;
output c665;
output c4352;
output c9356;
output c795;
output c2332;
output c4449;
output c8248;
output c9138;
output c8184;
output c8112;
output c9464;
output c6326;
output c0141;
output c07;
output c3270;
output c4212;
output c5384;
output c6345;
output c7357;
output c9369;
output c8175;
output c5118;
output c4295;
output c0116;
output c3365;
output c4307;
output c48;
output c7439;
output c0425;
output c2315;
output c0454;
output c8202;
output c9151;
output c2151;
output c4288;
output c1190;
output c6259;
output c9183;
output c6127;
output c7190;
output c8168;
output c780;
output c2434;
output c9384;
output c434;
output c4373;
output c6183;
output c3138;
output c160;
output c8186;
output c8456;
output c9234;
output c6352;
output c7477;
output c3424;
output c8394;
output c5402;
output c2288;
output c0453;
output c030;
output c2414;
output c4102;
output c4333;
output c1269;
output c4474;
output c2102;
output c857;
output c7133;
output c2423;
output c3243;
output c4447;
output c2235;
output c1243;
output c5123;
output c9276;
output c1150;
output c2246;
output c356;
output c9321;
output c577;
output c0140;
output c0313;
output c2498;
output c1211;
output c684;
output c1455;
output c0302;
output c3135;
output c2487;
output c3121;
output c888;
output c2145;
output c1274;
output c9494;
output c7342;
output c5168;
output c1338;
output c2304;
output c819;
output c1111;
output c4410;
output c1360;
output c5255;
output c4135;
output c9136;
output c3414;
output c4317;
output c5304;
output c6470;
output c7120;
output c3244;
output c1221;
output c7389;
output c1380;
output c072;
output c6129;
output c2404;
output c7230;
output c0199;
output c873;
output c5434;
output c2243;
output c911;
output c7399;
output c1483;
output c7467;
output c0275;
output c0337;
output c9233;
output c9281;
output c8197;
output c5205;
output c675;
output c7416;
output c1391;
output c3153;
output c846;
output c5321;
output c1460;
output c7351;
output c836;
output c3266;
output c381;
output c4371;
output c9121;
output c9311;
output c2211;
output c5122;
output c5217;
output c9345;
output c8169;
output c6338;
output c4260;
output c530;
output c9286;
output c8123;
output c14;
output c0498;
output c8298;
output c4418;
output c745;
output c149;
output c3219;
output c8342;
output c4364;
output c843;
output c8376;
output c3226;
output c5361;
output c3119;
output c2433;
output c7132;
output c775;
output c3262;
output c213;
output c3422;
output c7316;
output c7288;
output c3305;
output c4232;
output c5222;
output c3446;
output c9320;
output c9347;
output c6356;
output c4493;
output c0240;
output c177;
output c0402;
output c0160;
output c6209;
output c4454;
output c7218;
output c031;
output c2466;
output c3113;
output c0448;
output c9229;
output c6363;
output c8194;
output c0315;
output c6168;
output c6206;
output c6314;
output c0416;
output c3484;
output c6397;
output c754;
output c2431;
output c5179;
output c9471;
output c5388;
output c8225;
output c8229;
output c392;
output c4452;
output c6195;
output c5236;
output c7274;
output c427;
output c275;
output c8295;
output c4385;
output c418;
output c5427;
output c896;
output c9350;
output c5150;
output c5495;
output c4486;
output c4461;
output c629;
output c9359;
output c435;
output c3460;
output c1419;
output c2361;
output c925;
output c4415;
output c3102;
output c7479;
output c7180;
output c639;
output c3248;
output c5303;
output c469;
output c324;
output c1129;
output c662;
output c6275;
output c0327;
output c7106;
output c6467;
output c0401;
output c1174;
output c226;
output c2311;
output c932;
output c5181;
output c5129;
output c7465;
output c4328;
output c668;
output c0161;
output c68;
output c842;
output c049;
output c2289;
output c78;
output c7227;
output c5470;
output c5442;
output c8341;
output c496;
output c1255;
output c9108;
output c4168;
output c0311;
output c5359;
output c0115;
output c093;
output c7487;
output c9275;
output c9267;
output c5180;
output c8401;
output c2352;
output c279;
output c9440;
output c5106;
output c9212;
output c353;
output c95;
output c772;
output c9194;
output c3169;
output c8357;
output c1203;
output c7244;
output c4430;
output c1204;
output c6105;
output c3139;
output c9386;
output c5270;
output c9122;
output c2441;
output c569;
output c9442;
output c7343;
output c637;
output c8135;
output c5171;
output c6219;
output c743;
output c1384;
output c759;
output c098;
output c2442;
output c4383;
output c590;
output c3431;
output c0231;
output c7304;
output c3337;
output c4157;
output c1448;
output c2369;
output c468;
output c2277;
output c1280;
output c6286;
output c7305;
output c1343;
output c8359;
output c43;
output c6449;
output c7455;
output c84;
output c6119;
output c8181;
output c730;
output c4265;
output c7211;
output c3327;
output c8230;
output c4375;
output c8385;
output c5128;
output c1326;
output c889;
output c6182;
output c3452;
output c7140;
output c3329;
output c7257;
output c72;
output c8281;
output c692;
output c515;
output c7151;
output c955;
output c4432;
output c2368;
output c2425;
output c1216;
output c2301;
output c9134;
output c8178;
output c810;
output c5286;
output c560;
output c128;
output c4367;
output c1229;
output c6281;
output c8162;
output c8154;
output c3198;
output c6411;
output c3438;
output c3257;
output c2355;
output c7459;
output c4141;
output c6178;
output c2412;
output c0462;
output c9353;
output c387;
output c881;
output c7348;
output c8113;
output c2270;
output c9481;
output c3114;
output c3205;
output c1301;
output c3221;
output c1145;
output c3103;
output c9366;
output c0344;
output c5188;
output c440;
output c1329;
output c8365;
output c7329;
output c1287;
output c2159;
output c2262;
output c1371;
output c2274;
output c8343;
output c8373;
output c426;
output c582;
output c6116;
output c4331;
output c0220;
output c6179;
output c075;
output c2475;
output c4147;
output c5134;
output c7196;
output c1207;
output c7255;
output c6161;
output c1487;
output c0285;
output c4151;
output c6435;
output c5433;
output c315;
output c1339;
output c0249;
output c1140;
output c6458;
output c086;
output c1452;
output c5201;
output c2494;
output c111;
output c9449;
output c8459;
output c6223;
output c2175;
output c1124;
output c8351;
output c7484;
output c3454;
output c8347;
output c5457;
output c4411;
output c6292;
output c6124;
output c4136;
output c8448;
output c0323;
output c2464;
output c323;
output c5211;
output c2386;
output c0478;
output c0388;
output c7388;
output c0467;
output c5137;
output c5172;
output c8222;
output c1489;
output c9216;
output c0352;
output c2215;
output c9252;
output c9223;
output c9277;
output c268;
output c3228;
output c7162;
output c312;
output c9263;
output c2392;
output c4292;
output c592;
output c2164;
output c895;
output c9396;
output c965;
output c5189;
output c9291;
output c6313;
output c1114;
output c916;
output c1296;
output c085;
output c1232;
output c9309;
output c9407;
output c3240;
output c7447;
output c5110;
output c8411;
output c9107;
output c2193;
output c3306;
output c7283;
output c2479;
output c4266;
output c5302;
output c5424;
output c4194;
output c7490;
output c0472;
output c478;
output c9477;
output c3384;
output c1142;
output c7349;
output c633;
output c1257;
output c7225;
output c0331;
output c6306;
output c786;
output c36;
output c8176;
output c6322;
output c647;
output c9363;
output c3489;
output c3184;
output c052;
output c6320;
output c2439;
output c1364;
output c7273;
output c8257;
output c5408;
output c7236;
output c2185;
output c0274;
output c4166;
output c8484;
output c722;
output c9181;
output c354;
output c1401;
output c0164;
output c063;
output c8330;
output c2252;
output c5223;
output c475;
output c7458;
output c4301;
output c2146;
output c7469;
output c4372;
output c8410;
output c7378;
output c6174;
output c796;
output c4312;
output c9358;
output c0404;
output c7142;
output c059;
output c6181;
output c0370;
output c9451;
output c3321;
output c033;
output c4250;
output c752;
output c3267;
output c7193;
output c8247;
output c9178;
output c0348;
output c3211;
output c1271;
output c4494;
output c88;
output c4475;
output c0403;
output c0250;
output c628;
output c77;
output c3287;
output c9344;
output c4285;
output c7110;
output c5441;
output c4153;
output c8114;
output c3307;
output c2183;
output c5334;
output c9326;
output c2343;
output c3268;
output c9285;
output c1400;
output c4437;
output c4329;
output c6328;
output c16;
output c757;
output c131;
output c1183;
output c37;
output c4308;
output c884;
output c7446;
output c9226;
output c9114;
output c4417;
output c967;
output c4439;
output c6246;
output c2163;
output c3364;
output c7436;
output c0145;
output c3251;
output c7402;
output c5245;
output c5156;
output c7478;
output c245;
output c4150;
output c7468;
output c069;
output c5412;
output c17;
output c521;
output c257;
output c6390;
output c876;
output c5263;
output c4473;
output c0206;
output c9456;
output c1244;
output c0173;
output c2353;
output c8469;
output c4490;
output c6438;
output c56;
output c4116;
output c5248;
output c1480;
output c3326;
output c295;
output c1403;
output c817;
output c2259;
output c798;
output c599;
output c5432;
output c0192;
output c5186;
output c1166;
output c1252;
output c2417;
output c094;
output c7105;
output c1446;
output c0188;
output c6461;
output c0246;
output c1224;
output c6469;
output c2121;
output c689;
output c0417;
output c532;
output c42;
output c2247;
output c8221;
output c8250;
output c6347;
output c959;
output c2329;
output c9130;
output c6391;
output c9305;
output c998;
output c7100;
output c8292;
output c03;
output c4377;
output c0484;
output c5439;
output c1462;
output c5146;
output c078;
output c9379;
output c555;
output c296;
output c0405;
output c349;
output c3455;
output c574;
output c0266;
output c764;
output c4341;
output c5494;
output c7264;
output c9255;
output c0396;
output c7361;
output c9102;
output c347;
output c1214;
output c099;
output c1186;
output c1428;
output c4245;
output c5190;
output c1276;
output c2275;
output c7425;
output c8352;
output c6442;
output c2174;
output c7418;
output c6159;
output c1467;
output c34;
output c0392;
output c4214;
output c0397;
output c883;
output c813;
output c2314;
output c9156;
output c0113;
output c8487;
output c724;
output c8278;
output c755;
output c620;
output c7224;
output c731;
output c9186;
output c1109;
output c9211;
output c8253;
output c520;
output c0317;
output c0407;
output c3128;
output c6107;
output c5378;
output c962;
output c5315;
output c467;
output c4272;
output c8446;
output c9422;
output c45;
output c0309;
output c73;
output c548;
output c0142;
output c1152;
output c165;
output c3463;
output c2317;
output c7462;
output c5130;
output c0185;
output c0495;
output c552;
output c983;
output c7126;
output c2397;
output c3110;
output c0356;
output c8362;
output c8449;
output c6495;
output c7143;
output c1394;
output c5469;
output c8203;
output c491;
output c4237;
output c3272;
output c9144;
output c5452;
output c0460;
output c5237;
output c557;
output c7430;
output c112;
output c9323;
output c6454;
output c768;
output c7198;
output c8294;
output c4209;
output c2490;
output c1178;
output c1457;
output c792;
output c0339;
output c3362;
output c4173;
output c8336;
output c864;
output c2338;
output c2491;
output c984;
output c2154;
output c1437;
output c6394;
output c4247;
output c6118;
output c6480;
output c3423;
output c1181;
output c3232;
output c9499;
output c6419;
output c7101;
output c9485;
output c769;
output c5284;
output c3276;
output c122;
output c3214;
output c4197;
output c8101;
output c6269;
output c6408;
output c8498;
output c0393;
output c3356;
output c1350;
output c8420;
output c9303;
output c1223;
output c4202;
output c6463;
output c8243;
output c9306;
output c3354;
output c9242;
output c9120;
output c350;
output c9374;
output c8497;
output c5371;
output c838;
output c2229;
output c7207;
output c8289;
output c9432;
output c2292;
output c8296;
output c6488;
output c288;
output c8396;
output c3210;
output c7344;
output c9331;
output c0114;
output c4419;
output c0391;
output c3490;
output c2225;
output c1463;
output c8355;
output c8110;
output c3236;
output c9261;
output c373;
output c7491;
output c0191;
output c4356;
output c2419;
output c8208;
output c2468;
output c036;
output c3407;
output c791;
output c6482;
output c622;
output c1431;
output c961;
output c2197;
output c4315;
output c5173;
output c4398;
output c8427;
output c2155;
output c9433;
output c9296;
output c3233;
output c7214;
output c7319;
output c367;
output c264;
output c376;
output c4431;
output c645;
output c912;
output c7270;
output c4231;
output c060;
output c3355;
output c1456;
output c0284;
output c0421;
output c3166;
output c5182;
output c6409;
output c494;
output c3405;
output c9132;
output c8337;
output c3465;
output c4425;
output c524;
output c5214;
output c2172;
output c248;
output c7258;
output c1300;
output c8475;
output c2348;
output c977;
output c2460;
output c317;
output c6299;
output c4389;
output c8490;
output c4393;
output c7375;
output c0136;
output c6258;
output c4179;
output c8264;
output c8130;
output c2467;
output c4282;
output c824;
output c2461;
output c8389;
output c2321;
output c5403;
output c6444;
output c9395;
output c2384;
output c2233;
output c9490;
output c5445;
output c3386;
output c538;
output c915;
output c4164;
output c841;
output c1396;
output c9335;
output c041;
output c9105;
output c8321;
output c444;
output c6163;
output c8305;
output c9330;
output c0195;
output c0466;
output c2308;
output c0479;
output c6268;
output c5141;
output c6489;
output c0236;
output c937;
output c5326;
output c6122;
output c614;
output c1406;
output c9417;
output c1270;
output c0245;
output c7197;
output c9497;
output c8251;
output c413;
output c2242;
output c6192;
output c024;
output c2190;
output c4219;
output c0440;
output c0325;
output c5400;
output c3141;
output c762;
output c18;
output c5417;
output c0223;
output c8470;
output c1389;
output c0257;
output c529;
output c9123;
output c1488;
output c3304;
output c2228;
output c1491;
output c2111;
output c0117;
output c7204;
output c9462;
output c0438;
output c280;
output c3470;
output c641;
output c7239;
output c9167;
output c591;
output c7124;
output c0293;
output c5370;
output c018;
output c130;
output c1348;
output c9319;
output c4300;
output c671;
output c9169;
output c9450;
output c9314;
output c7266;
output c9192;
output c9455;
output c4472;
output c871;
output c2299;
output c6154;
output c1334;
output c0133;
output c4340;
output c1459;
output c285;
output c4304;
output c94;
output c718;
output c6282;
output c446;
output c7131;
output c5488;
output c5260;
output c5268;
output c6369;
output c3353;
output c140;
output c2359;
output c7496;
output c2128;
output c734;
output c8116;
output c9142;
output c1385;
output c2223;
output c930;
output c453;
output c7134;
output c5342;
output c0276;
output c4346;
output c6361;
output c089;
output c2438;
output c0434;
output c0259;
output c6287;
output c1298;
output c7160;
output c744;
output c2381;
output c1416;
output c5401;
output c0303;
output c7169;
output c6349;
output c2396;
output c8211;
output c9402;
output c3380;
output c6218;
output c0151;
output c3156;
output c8353;
output c7269;
output c3345;
output c7453;
output c8146;
output c7340;
output c3488;
output c3144;
output c6207;
output c7298;
output c8435;
output c5436;
output c0103;
output c9298;
output c5347;
output c0122;
output c2263;
output c9405;
output c973;
output c6111;
output c6490;
output c6355;
output c4233;
output c7390;
output c7287;
output c6298;
output c0341;
output c0459;
output c9348;
output c7372;
output c6439;
output c9370;
output c1193;
output c2363;
output c2496;
output c1235;
output c0295;
output c1254;
output c7184;
output c1279;
output c5479;
output c7115;
output c8131;
output c13;
output c93;
output c658;
output c6187;
output c0235;
output c1454;
output c9342;
output c7347;
output c6368;
output c497;
output c8474;
output c6216;
output c2178;
output c9385;
output c6485;
output c2210;
output c492;
output c1263;
output c8422;
output c338;
output c1286;
output c2236;
output c6312;
output c2360;
output c6365;
output c7384;
output c47;
output c6151;
output c170;
output c429;
output c7253;
output c2495;
output c9179;
output c0182;
output c0201;
output c2261;
output c3392;
output c8273;
output c0143;
output c9474;
output c9247;
output c3104;
output c921;
output c9172;
output c1239;
output c2349;
output c9297;
output c422;
output c0277;
output c0408;
output c2115;
output c9441;
output c2251;
output c0176;
output c9109;
output c2199;
output c019;
output c7415;
output c913;
output c3444;
output c1330;
output c2240;
output c118;
output c8102;
output c4403;
output c9283;
output c5354;
output c2165;
output c9428;
output c4143;
output c9340;
output c240;
output c1118;
output c3152;
output c6186;
output c4484;
output c972;
output c121;
output c2459;
output c4208;
output c3209;
output c4499;
output c379;
output c5259;
output c2157;
output c0321;
output c5145;
output c5311;
output c3147;
output c2207;
output c9131;
output c8285;
output c278;
output c5101;
output c1205;
output c682;
output c6188;
output c0159;
output c3255;
output c020;
output c6255;
output c6348;
output c774;
output c8372;
output c488;
output c4239;
output c7176;
output c244;
output c4174;
output c251;
output c397;
output c449;
output c861;
output c6309;
output c83;
output c0252;
output c5153;
output c7483;
output c5476;
output c4111;
output c2100;
output c7481;
output c3286;
output c815;
output c1277;
output c892;
output c4399;
output c1116;
output c135;
output c156;
output c6440;
output c8421;
output c4170;
output c657;
output c5421;
output c1461;
output c3109;
output c4322;
output c4388;
output c4421;
output c49;
output c0412;
output c0128;
output c0316;
output c523;
output c9452;
output c7206;
output c1387;
output c1177;
output c416;
output c9153;
output c1414;
output c4353;
output c9271;
output c2176;
output c991;
output c92;
output c5423;
output c1479;
output c9476;
output c8103;
output c382;
output c5349;
output c3183;
output c29;
output c9206;
output c1378;
output c8288;
output c6373;
output c85;
output c0205;
output c8374;
output c6266;
output c6396;
output c362;
output c1451;
output c2375;
output c5228;
output c5149;
output c8228;
output c1195;
output c8276;
output c351;
output c115;
output c8270;
output c380;
output c8492;
output c174;
output c477;
output c7205;
output c7135;
output c0389;
output c46;
output c1313;
output c9282;
output c084;
output c7407;
output c3499;
output c0450;
output c3341;
output c7386;
output c4443;
output c0147;
output c4234;
output c0158;
output c6245;
output c2173;
output c5366;
output c9398;
output c247;
output c0384;
output c3469;
output c0121;
output c8485;
output c8360;
output c0461;
output c3447;
output c829;
output c9378;
output c3379;
output c2217;
output c554;
output c4210;
output c2379;
output c1261;
output c8379;
output c9302;
output c5336;
output c8160;
output c0139;
output c331;
output c5116;
output c470;
output c6261;
output c6475;
output c634;
output c4444;
output c1450;
output c4103;
output c5132;
output c1139;
output c8106;
output c2427;
output c7431;
output c51;
output c7277;
output c273;
output c5210;
output c8179;
output c6325;
output c522;
output c0282;
output c9101;
output c7480;
output c8166;
output c9376;
output c2457;
output c3242;
output c981;
output c7364;
output c1314;
output c8234;
output c782;
output c142;
output c1315;
output c3334;
output c8308;
output c4351;
output c116;
output c512;
output c3456;
output c926;
output c3155;
output c9438;
output c3497;
output c6180;
output c045;
output c8152;
output c1312;
output c1310;
output c4228;
output c98;
output c9318;
output c1133;
output c6228;
output c6117;
output c7440;
output c1320;
output c7366;
output c6137;
output c9380;
output c5293;
output c5152;
output c0263;
output c8148;
output c5241;
output c191;
output c4192;
output c526;
output c7369;
output c2333;
output c5393;
output c3450;
output c9333;
output c7203;
output c4394;
output c6189;
output c495;
output c7276;
output c3352;
output c1262;
output c0213;
output c1425;
output c8290;
output c4113;
output c9461;
output c4284;
output c0262;
output c5249;
output c180;
output c1438;
output c90;
output c5346;
output c0497;
output c7417;
output c0202;
output c096;
output c327;
output c1176;
output c1141;
output c0330;
output c0445;
output c8473;
output c6260;
output c1210;
output c4146;
output c3143;
output c5144;
output c797;
output c0219;
output c335;
output c0154;
output c0107;
output c0314;
output c7103;
output c7383;
output c291;
output c0399;
output c6280;
output c6386;
output c3160;
output c86;
output c770;
output c6316;
output c2391;
output c8133;
output c1433;
output c9403;
output c4241;
output c1383;
output c6239;
output c8430;
output c3136;
output c9357;
output c827;
output c4203;
output c3290;
output c182;
output c8437;
output c0167;
output c5264;
output c0118;
output c5178;
output c954;
output c3389;
output c3275;
output c8226;
output c9187;
output c0357;
output c3273;
output c8241;
output c2202;
output c3300;
output c7397;
output c7210;
output c8188;
output c1405;
output c246;
output c3193;
output c4380;
output c480;
output c8476;
output c516;
output c8212;
output c4483;
output c451;
output c1148;
output c0299;
output c1256;
output c5215;
output c6360;
output c4381;
output c1355;
output c1302;
output c4491;
output c6378;
output c3158;
output c6413;
output c0261;
output c6125;
output c4109;
output c8440;
output c2330;
output c5231;
output c1100;
output c459;
output c2393;
output c9489;
output c9100;
output c1202;
output c6215;
output c4326;
output c9473;
output c9488;
output c5337;
output c9444;
output c0251;
output c9301;
output c1304;
output c6247;
output c4395;
output c0255;
output c8328;
output c3310;
output c9365;
output c2409;
output c0172;
output c2398;
output c2182;
output c3434;
output c3473;
output c8486;
output c1402;
output c113;
output c3363;
output c5147;
output c763;
output c26;
output c7332;
output c7111;
output c3279;
output c2395;
output c7476;
output c6476;
output c9189;
output c7123;
output c0486;
output c814;
output c4478;
output c6229;
output c3374;
output c533;
output c936;
output c4488;
output c9325;
output c179;
output c943;
output c5377;
output c4442;
output c4122;
output c8282;
output c1464;
output c3367;
output c6357;
output c0481;
output c7259;
output c5461;
output c4365;
output c6374;
output c1294;
output c7301;
output c5199;
output c0494;
output c7289;
output c9315;
output c852;
output c3280;
output c9328;
output c4223;
output c3118;
output c6465;
output c0152;
output c2279;
output c8443;
output c254;
output c4361;
output c1217;
output c3101;
output c7291;
output c3439;
output c157;
output c7472;
output c6263;
output c23;
output c3324;
output c3132;
output c1429;
output c425;
output c6289;
output c7119;
output c8304;
output c6170;
output c2416;
output c2144;
output c7166;
output c2148;
output c2280;
output c0228;
output c1259;
output c3397;
output c5374;
output c5428;
output c4355;
output c457;
output c9401;
output c7118;
output c0105;
output c6221;
output c0132;
output c3351;
output c1281;
output c1482;
output c0439;
output c3476;
output c3125;
output c232;
output c0180;
output c536;
output c4117;
output c5406;
output c3382;
output c5314;
output c2195;
output c3360;
output c8477;
output c4152;
output c793;
output c5462;
output c2287;
output c1290;
output c9257;
output c5289;
output c5104;
output c559;
output c8155;
output c0101;
output c0475;
output c360;
output c9334;
output c7473;
output c5437;
output c5121;
output c6418;
output c6167;
output c448;
output c8316;
output c616;
output c9117;
output c6484;
output c1123;
output c5473;
output c4349;
output c039;
output c60;
output c544;
output c9147;
output c3357;
output c042;
output c9217;
output c8377;
output c0243;
output c923;
output c6202;
output c3396;
output c4323;
output c5379;
output c8120;
output c2307;
output c466;
output c0278;
output c7254;
output c1417;
output c0187;
output c082;
output c5139;
output c8153;
output c928;
output c6112;
output c5170;
output c1362;
output c5362;
output c5243;
output c5312;
output c2106;
output c69;
output c5301;
output c0137;
output c3317;
output c8418;
output c4338;
output c3117;
output c3457;
output c7406;
output c3375;
output c9278;
output c952;
output c9478;
output c5383;
output c0270;
output c6417;
output c0138;
output c1147;
output c2265;
output c0222;
output c9260;
output c953;
output c8441;
output c1143;
output c6121;
output c1182;
output c1418;
output c8277;
output c7350;
output c2124;
output c1305;
output c8254;
output c0413;
output c09;
output c2281;
output c3246;
output c6407;
output c2372;
output c823;
output c1317;
output c3178;
output c236;
output c869;
output c293;
output c0414;
output c3182;
output c6128;
output c8143;
output c837;
output c5453;
output c2340;
output c6497;
output c9204;
output c9454;
output c0296;
output c6285;
output c0234;
output c3127;
output c1168;
output c8216;
output c2327;
output c9214;
output c8177;
output c5425;
output c4213;
output c428;
output c173;
output c7275;
output c9251;
output c6277;
output c162;
output c3284;
output c6244;
output c993;
output c1390;
output c1212;
output c6265;
output c8413;
output c4104;
output c4140;
output c5143;
output c931;
output c0319;
output c9129;
output c3189;
output c6303;
output c8164;
output c562;
output c8275;
output c740;
output c150;
output c5477;
output c3130;
output c0130;
output c061;
output c6420;
output c9316;
output c139;
output c4476;
output c8423;
output c652;
output c6145;
output c3150;
output c155;
output c517;
output c9177;
output c2220;
output c698;
output c2147;
output c4354;
output c1367;
output c1344;
output c6172;
output c4276;
output c5256;
output c7104;
output c8412;
output c878;
output c05;
output c0184;
output c9227;
output c0429;
output c4159;
output c2300;
output c6169;
output c0383;
output c7368;
output c5240;
output c811;
output c6106;
output c266;
output c087;
output c141;
output c4412;
output c8284;
output c7267;
output c4128;
output c6375;
output c0345;
output c9409;
output c558;
output c2271;
output c4267;
output c597;
output c9185;
output c1173;
output c945;
output c4236;
output c193;
output c374;
output c3421;
output c252;
output c6491;
output c7412;
output c8238;
output c8416;
output c272;
output c163;
output c5409;
output c070;
output c70;
output c816;
output c7128;
output c3308;
output c2488;
output c5490;
output c8244;
output c2411;
output c6425;
output c9368;
output c9436;
output c8147;
output c8132;
output c1191;
output c2341;
output c4132;
output c9492;
output c2166;
output c9360;
output c2129;
output c1470;
output c1249;
output c1377;
output c2320;
output c853;
output c7320;
output c858;
output c0423;
output c9191;
output c1242;
output c748;
output c9419;
output c5117;
output c7441;
output c6197;
output c8457;
output c3466;
output c7334;
output c7174;
output c2127;
output c3359;
output c5467;
output c3180;
output c490;
output c4485;
output c0349;
output c6288;
output c1478;
output c3170;
output c7442;
output c3176;
output c3498;
output c1309;
output c5221;
output c9197;
output c2481;
output c417;
output c4366;
output c5415;
output c1375;
output c546;
output c0492;
output c5297;
output c0360;
output c8279;
output c1272;
output c023;
output c621;
output c877;
output c066;
output c975;
output c2238;
output c7492;
output c997;
output c6185;
output c8332;
output c9256;
output c8182;
output c3215;
output c0436;
output c1352;
output c7261;
output c1332;
output c0237;
output c1267;
output c6432;
output c6198;
output c7154;
output c9399;
output c2276;
output c3320;
output c59;
output c5318;
output c7427;
output c3486;
output c65;
output c7168;
output c0165;
output c4127;
output c146;
output c0342;
output c79;
output c8163;
output c8415;
output c678;
output c5174;
output c8493;
output c186;
output c6196;
output c346;
output c5247;
output c4498;
output c9243;
output c1436;
output c2216;
output c4434;
output c6233;
output c527;
output c7130;
output c1101;
output c3265;
output c1499;
output c3271;
output c0390;
output c7252;
output c9337;
output c8218;
output c2406;
output c1265;
output c778;
output c7216;
output c3403;
output c3494;
output c0471;
output c9249;
output c4318;
output c941;
output c7404;
output c8366;
output c9139;
output c3393;
output c262;
output c3433;
output c6227;
output c5364;
output c1423;
output c1237;
output c626;
output c375;
output c0209;
output c4186;
output c7422;
output c899;
output c5246;
output c0343;
output c0374;
output c2370;
output c7475;
output c2400;
output c0488;
output c9460;
output c8439;
output c4489;
output c015;
output c2465;
output c5131;
output c9119;
output c2135;
output c4118;
output c4218;
output c3269;
output c9193;
output c6331;
output c3415;
output c5277;
output c5391;
output c1131;
output c8407;
output c4344;
output c6311;
output c2192;
output c7358;
output c1121;
output c9412;
output c1236;
output c3369;
output c1335;
output c017;
output c9170;
output c4172;
output c7474;
output c1495;
output c9388;
output c1412;
output c64;
output c5344;
output c3212;
output c0373;
output c2326;
output c994;
output c4263;
output c8405;
output c223;
output c4441;
output c5444;
output c7153;
output c9459;
output c3111;
output c6441;
output c9354;
output c99;
output c4481;
output c9472;
output c6123;
output c5164;
output c0441;
output c6144;
output c7413;
output c0432;
output c4242;
output c2383;
output c0232;
output c5169;
output c6403;
output c8198;
output c971;
output c2448;
output c4154;
output c890;
output c4178;
output c7370;
output c0333;
output c6447;
output c299;
output c411;
output c2107;
output c3411;
output c585;
output c377;
output c8488;
output c5176;
output c8256;
output c4459;
output c6211;
output c534;
output c4101;
output c8151;
output c0437;
output c2474;
output c5112;
output c4216;
output c6395;
output c9415;
output c5455;
output c0242;
output c8392;
output c5483;
output c2214;
output c2482;
output c4368;
output c3261;
output c6423;
output c7247;
output c2254;
output c0217;
output c249;
output c0153;
output c037;
output c4240;
output c7326;
output c1376;
output c2376;
output c3200;
output c5410;
output c9313;
output c6310;
output c733;
output c9414;
output c0326;
output c7336;
output c0368;
output c1336;
output c2334;
output c6323;
output c2250;
output c1104;
output c8224;
output c154;
output c7420;
output c783;
output c265;
output c7159;
output c8479;
output c5126;
output c4360;
output c259;
output c394;
output c7155;
output c2424;
output c6201;
output c0149;
output c2161;
output c8161;
output c3253;
output c0367;
output c7433;
output c2208;
output c7392;
output c3404;
output c6452;
output c8455;
output c8301;
output c6387;
output c9220;
output c21;
output c2385;
output c4271;
output c9225;
output c1445;
output c057;
output c9213;
output c412;
output c3419;
output c1130;
output c9352;
output c7470;
output c187;
output c5194;
output c0490;
output c6459;
output c8105;
output c129;
output c286;
output c1246;
output c2132;
output c8463;
output c1162;
output c0451;
output c8107;
output c9391;
output c25;
output c2415;
output c9289;
output c8438;
output c5498;
output c0109;
output c6114;
output c663;
output c8451;
output c1219;
output c833;
output c1427;
output c175;
output c011;
output c2258;
output c9159;
output c3312;
output c9140;
output c0129;
output c4138;
output c74;
output c4426;
output c8141;
output c2362;
output c849;
output c4405;
output c0419;
output c7186;
output c2291;
output c4119;
output c697;
output c924;
output c3378;
output c7449;
output c1110;
output c4370;
output c5250;
output c0207;
output c0272;
output c9143;
output c0328;
output c9400;
output c3203;
output c6270;
output c7443;
output c5229;
output c8335;
output c7185;
output c2196;
output c4131;
output c7235;
output c9137;
output c6372;
output c1189;
output c9221;
output c8299;
output c4108;
output c1333;
output c4144;
output c8122;
output c5482;
output c738;
output c5333;
output c219;
output c5485;
output c7114;
output c693;
output c0196;
output c1136;
output c0241;
output c3185;
output c9274;
output c1119;
output c0170;
output c5185;
output c7178;
output c6156;
output c0354;
output c695;
output c0186;
output c132;
output c168;
output c539;
output c4262;
output c3347;
output c0124;
output c5307;
output c9207;
output c7290;
output c5369;
output c3140;
output c1201;
output c445;
output c9125;
output c5405;
output c2452;
output c615;
output c9238;
output c729;
output c1160;
output c9200;
output c0418;
output c5291;
output c6494;
output c6267;
output c7138;
output c3451;
output c8136;
output c4169;
output c221;
output c410;
output c946;
output c880;
output c5175;
output c0221;
output c8313;
output c6204;
output c5279;
output c9418;
output c5151;
output c8128;
output c2237;
output c9284;
output c7158;
output c7122;
output c5138;
output c9253;
output c1393;
output c9270;
output c1472;
output c8207;
output c938;
output c0430;
output c8312;
output c9446;
output c00;
output c0267;
output c0322;
output c887;
output c5305;
output c4391;
output c9495;
output c1192;
output c239;
output c826;
output c944;
output c7499;
output c7164;
output c8433;
output c0420;
output c1397;
output c8280;
output c9362;
output c9427;
output c7152;
output c0433;
output c8195;
output c342;
output c7108;
output c856;
output c8467;
output c2445;
output c5135;
output c656;
output c5120;
output c7148;
output c7367;
output c2346;
output c489;
output c6222;
output c1486;
output c5200;
output c2446;
output c7362;
output c7222;
output c0362;
output c2283;
output c2104;
output c2109;
output c3377;
output c8367;
output c2447;
output c643;
output c0100;
output c8268;
output c073;
output c255;
output c333;
output c4467;
output c4397;
output c1366;
output c2312;
output c751;
output c1213;
output c7489;
output c3213;
output c8274;
output c4124;
output c1284;
output c2110;
output c8115;
output c2485;
output c8445;
output c5328;
output c9279;
output c5367;
output c9443;
output c4283;
output c4496;
output c028;
output c5285;
output c7373;
output c885;
output c935;
output c1494;
output c097;
output c4466;
output c9128;
output c6371;
output c9262;
output c787;
output c2336;
output c5426;
output c8419;
output c510;
output c5127;
output c9184;
output c0308;
output c5351;
output c8465;
output c0452;
output c5499;
output c2152;
output c910;
output c2105;
output c4492;
output c8170;
output c8499;
output c5308;
output c4400;
output c9486;
output c8300;
output c1253;
output c5298;
output c720;
output c4378;
output c6389;
output c511;
output c1245;
output c571;
output c5299;
output c96;
output c6321;
output c980;
output c7471;
output c1175;
output c5323;
output c2180;
output c7493;
output c7248;
output c238;
output c8157;
output c4436;
output c8447;
output c1382;
output c1138;
output c948;
output c750;
output c5324;
output c185;
output c8382;
output c1341;
output c158;
output c6401;
output c9155;
output c8324;
output c3338;
output c3301;
output c1188;
output c055;
output c1222;
output c5261;
output c985;
output c322;
output c292;
output c1426;
output c384;
output c7318;
output c383;
output c8145;
output c5317;
output c6377;
output c9146;
output c6376;
output c026;
output c5184;
output c2458;
output c5465;
output c566;
output c966;
output c785;
output c6343;
output c9467;
output c6333;
output c5234;
output c5266;
output c7278;
output c2295;
output c3274;
output c0131;
output c3230;
output c8460;
output c1439;
output c1324;
output c9484;
output c9111;
output c5219;
output c7181;
output c0226;
output c120;
output c1407;
output c587;
output c5114;
output c398;
output c9248;
output c053;
output c2470;
output c934;
output c0294;
output c2302;
output c1120;
output c4468;
output c4270;
output c3204;
output c6276;
output c2408;
output c436;
output c1289;
output c9382;
output c074;
output c4287;
output c1442;
output c0181;
output c649;
output c9273;
output c6148;
output c696;
output c6295;
output c3120;
output c3340;
output c9265;
output c963;
output c821;
output c3395;
output c7324;
output c4280;
output c320;
output c4195;
output c022;
output c2310;
output c04;
output c2469;
output c691;
output c3190;
output c9173;
output c0340;
output c2206;
output c7353;
output c735;
output c3154;
output c5454;
output c567;
output c9171;
output c9317;
output c190;
output c3427;
output c1374;
output c077;
output c1154;
output c3133;
output c24;
output c2149;
output c6499;
output c2428;
output c7137;
output c588;
output c7363;
output c0119;
output c138;
output c8269;
output c9157;
output c1386;
output c430;
output c5198;
output c6262;
output c6399;
output c922;
output c3131;
output c742;
output c1156;
output c8320;
output c4424;
output c1392;
output c3385;
output c8371;
output c0148;
output c8431;
output c7411;
output c4211;
output c5430;
output c6496;
output c1171;
output c3491;
output c4220;
output c4343;
output c0260;
output c334;
output c8201;
output c4336;
output c719;
output c5161;
output c5157;
output c8140;
output c7228;
output c8450;
output c3151;
output c1443;
output c7381;
output c3314;
output c7328;
output c5419;
output c8309;
output c6217;
output c5288;
output c3429;
output c1474;
output c0364;
output c5373;
output c3258;
output c088;
output c9377;
output c8111;
output c5329;
output c4453;
output c8302;
output c50;
output c044;
output c456;
output c0208;
output c4450;
output c7376;
output c2227;
output c6308;
output c7327;
output c5450;
output c9231;
output c231;
output c2471;
output c8291;
output c7161;
output c9389;
output c2177;
output c1137;
output c4386;
output c561;
output c5411;
output c3142;
output c3425;
output c8426;
output c0248;
output c4438;
output c6424;
output c7146;
output c6486;
output c0386;
output c767;
output c0320;
output c2380;
output c0426;
output c4187;
output c9416;
output c6446;
output c2118;
output c184;
output c9295;
output c1322;
output c3468;
output c4185;
output c6414;
output c0271;
output c9367;
output c2410;
output c3481;
output c694;
output c9493;
output c2492;
output c9232;
output c1413;
output c0239;
output c7429;
output c8171;
output c8129;
output c2443;
output c3325;
output c2364;
output c095;
output c271;
output c6162;
output c2117;
output c3163;
output c8378;
output c294;
output c549;
output c6437;
output c8489;
output c9205;
output c9287;
output c7183;
output c0200;
output c365;
output c8261;
output c3146;
output c3277;
output c358;
output c8185;
output c9483;
output c6143;
output c8496;
output c8227;
output c8232;
output c1358;
output c5306;
output c6468;
output c2290;
output c927;
output c2187;
output c2244;
output c8344;
output c4215;
output c715;
output c4134;
output c737;
output c9393;
output c0286;
output c683;
output c2278;
output c9406;
output c40;
output c6364;
output c4337;
output c4420;
output c2390;
output c6126;
output c0230;
output c651;
output c0178;
output c6462;
output c886;
output c7116;
output c2160;
output c7109;
output c4409;
output c8174;
output c7215;
output c3196;
output c9392;
output c7408;
output c0406;
output c872;
output c4440;
output c4446;
output c642;
output c9264;
output c2354;
output c9372;
output c9373;
output c7359;
output c1208;
output c0183;
output c5418;
output c133;
output c659;
output c1185;
output c0162;
output c5107;
output c5100;
output c4445;
output c0446;
output c7145;
output c4256;
output c464;
output c8204;
output c0289;
output c8381;
output c8193;
output c9133;
output c5287;
output c6324;
output c3426;
output c9258;
output c5310;
output c537;
output c0268;
output c1125;
output c3344;
output c3227;
output c2371;
output c378;
output c1163;
output c2249;
output c176;
output c5422;
output c8495;
output c1144;
output c6290;
output c97;
output c8454;
output c2205;
output c2454;
output c685;
output c0477;
output c7202;
output c4406;
output c0470;
output c5448;
output c3137;
output c0353;
output c918;
output c7460;
output c960;
output c4306;
output c7308;
output c4255;
output c1132;
output c8354;
output c9158;
output c9411;
output c81;
output c4244;
output c875;
output c6302;
output c4277;
output c39;
output c1308;
output c7435;
output c5155;
output c5204;
output c8414;
output c87;
output c9148;
output c9466;
output c8406;
output c3256;
output c310;
output c476;
output c336;
output c5416;
output c1194;
output c8334;
output c345;
output c6301;
output c5340;
output c5162;
output c0458;
output c8239;
output c7341;
output c0351;
output c681;
output c4121;
output c5492;
output c065;
output c415;
output c2120;
output c2344;
output c568;
output c832;
output c2222;
output c7315;
output c7121;
output c9336;
output c6274;
output c145;
output c7360;
output c6200;
output c3186;
output c4268;
output c8395;
output c8387;
output c968;
output c739;
output c5396;
output c6366;
output c3482;
output c253;
output c5356;
output c5273;
output c7377;
output c0410;
output c2357;
output c1303;
output c2477;
output c3278;
output c1149;
output c2143;
output c5196;
output c5274;
output c666;
output c0108;
output c6429;
output c6332;
output c7398;
output c8356;
output c6133;
output c2142;
output c1151;
output c9269;
output c8402;
output c3348;
output c5209;
output c3168;
output c7432;
output c4227;
output c5187;
output c5365;
output c6346;
output c3281;
output c01;
output c677;
output c939;
output c598;
output c5322;
output c6238;
output c4455;
output c4175;
output c3370;
output c2230;
output c2103;
output c0279;
output c6205;
output c9404;
output c5167;
output c421;
output c1251;
output c867;
output c067;
output c1435;
output c2141;
output c4200;
output c1112;
output c995;
output c6158;
output c2440;
output c8231;
output c8134;
output c035;
output c6257;
output c3394;
output c648;
output c6235;
output c66;
output c9161;
output c6336;
output c243;
output c4142;
output c9410;
output c0292;
output c820;
output c4345;
output c6318;
output c0473;
output c0155;
output c3373;
output c5360;
output c625;
output c9375;
output c6402;
output c047;
output c461;
output c2282;
output c1161;
output c747;
output c050;
output c092;
output c0493;
output c329;
output c0318;
output c3318;
output c2294;
output c313;
output c3145;
output c514;
output c3335;
output c7299;
output c1493;
output c8429;
output c0358;
output c2437;
output c8199;
output c4149;
output c7256;
output c7331;
output c596;
output c1476;
output c4161;
output c9435;
output c3398;
output c9152;
output c4422;
output c7191;
output c1359;
output c3328;
output c2319;
output c8384;
output c2221;
output c67;
output c5327;
output c7335;
output c1199;
output c8265;
output c3172;
output c9254;
output c7177;
output c4379;
output c830;
output c6199;
output c4302;
output c3358;
output c7272;
output c6406;
output c8139;
output c3296;
output c5487;
output c164;
output c474;
output c2356;
output c7241;
output c3222;
output c957;
output c2136;
output c0424;
output c8233;
output c1356;
output c1369;
output c234;
output c4427;
output c3202;
output c3129;
output c016;
output c062;
output c9235;
output c7385;
output c4314;
output c687;
output c1187;
output c7380;
output c4382;
output c3366;
output c41;
output c6212;
output c2418;
output c627;
output c4148;
output c5394;
output c2345;
output c7452;
output c442;
output c3289;
output c8323;
output c2449;
output c8393;
output c2256;
output c2342;
output c5108;
output c064;
output c7229;
output c6138;
output c6478;
output c6307;
output c6421;
output c586;
output c1126;
output c721;
output c3197;
output c460;
output c8370;
output c126;
output c210;
output c5271;
output c9361;
output c6479;
output c1146;
output c3420;
output c0355;
output c4342;
output c8255;
output c276;
output c3126;
output c274;
output c9230;
output c868;
output c1122;
output c4392;
output c5158;
output c52;
output c2200;
output c1477;
output c02;
output c6319;
output c7296;
output c7306;
output c6273;
output c1496;
output c0298;
output c3474;
output c4369;
output c229;
output c8172;
output c091;
output c8173;
output c6492;
output c7208;
output c3416;
output c3449;
output c9224;
output c4126;
output c9245;
output c6237;
output c4297;
output c5392;
output c6213;
output c0177;
output c2303;
output c4362;
output c9341;
output c58;
output c0379;
output c1117;
output c3249;
output c3162;
output c2134;
output c1444;
output c6283;
output c5431;
output c1440;
output c594;
output c5276;
output c486;
output c595;
output c9195;
output c385;
output c38;
output c632;
output c5192;
output c6147;
output c4191;
output c6379;
output c1421;
output c3239;
output c5463;
output c756;
output c9324;
output c2133;
output c5230;
output c4249;
output c667;
output c6160;
output c2219;
output c0134;
output c0307;
output c6173;
output c2137;
output c4359;
output c8340;
output c5459;
output c1285;
output c9124;
output c8283;
output c5292;
output c831;
output c8434;
output c3479;
output c1105;
output c9463;
output c9218;
output c147;
output c9168;
output c455;
output c4482;
output c8138;
output c0210;
output c3225;
output c014;
output c3372;
output c399;
output c1447;
output c242;
output c9113;
output c5358;
output c5283;
output c0288;
output c3323;
output c197;
output c433;
output c5290;
output c20;
output c277;
output c2189;
output c2377;
output c8180;
output c9293;
output c8346;
output c1399;
output c4309;
output c1273;
output c1395;
output c7423;
output c2420;
output c5493;
output c5480;
output c714;
output c1258;
output c920;
output c9470;
output c5159;
output c2268;
output c5352;
output c5257;
output c8266;
output c8189;
output c153;
output c5102;
output c2139;
output c119;
output c578;
output c0283;
output c727;
output c4182;
output c9338;
output c513;
output c5497;
output c1485;
output c7314;
output c2234;
output c5348;
output c3471;
output c7157;
output c949;
output c9349;
output c1410;
output c2435;
output c6176;
output c432;
output c4396;
output c5262;
output c8481;
output c9166;
output c879;
output c8350;
output c53;
output c1321;
output c1103;
output c7136;
output c1165;
output c8159;
output c32;
output c986;
output c4407;
output c7282;
output c3349;
output c5385;
output c7300;
output c4316;
output c7338;
output c3458;
output c8442;
output c7171;
output c8428;
output c7424;
output c3124;
output c661;
output c2273;
output c8452;
output c5265;
output c6455;
output c0106;
output c361;
output c4105;
output c2119;
output c1230;
output c4320;
output c9219;
output c7175;
output c1347;
output c290;
output c5254;
output c5160;
output c882;
output c1497;
output c3108;
output c6190;
output c5468;
output c4357;
output c4229;
output c2493;
output c7265;
output c454;
output c7382;
output c776;
output c4289;
output c5281;
output c8217;
output c9112;
output c2389;
output c8246;
output c6456;
output c9190;
output c0378;
output c4163;
output c4198;
output c4275;
output c4253;
output c3467;
output c224;
output c5447;
output c1264;
output c1102;
output c6464;
output c8260;
output c7461;
output c732;
output c2351;
output c618;
output c5458;
output c1172;
output c9174;
output c3418;
output c3399;
output c0216;
output c013;
output c6340;
output c5332;
output c4423;
output c540;
output c7396;
output c5300;
output c9394;
output c1206;
output c9448;
output c2296;
output c6102;
output c1449;
output c319;
output c0480;
output c485;
output c8494;
output c5464;
output c8326;
output c3191;
output c438;
output c0489;
output c761;
output c0171;
output c929;
output c1370;
output c7240;
output c441;
output c9103;
output c1471;
output c6254;
output c4376;
output c893;
output c260;
output c726;
output c4238;
output c1404;
output c686;
output c144;
output c611;
output c0363;
output c0111;
output c7163;
output c9429;
output c8311;
output c4261;
output c0375;
output c5244;
output c357;
output c3157;
output c5125;
output c9307;
output c44;
output c2293;
output c7173;
output c8287;
output c3107;
output c3115;
output c660;
output c7428;
output c624;
output c0168;
output c6253;
output c0204;
output c283;
output c1368;
output c5420;
output c1484;
output c9327;
output c2422;
output c7448;
output c8124;
output c3445;
output c7419;
output c8165;
output c9491;
output c6460;
output c481;
output c9294;
output c7486;
output c051;
output c3315;
output c9387;
output c9469;
output c6466;
output c484;
output c389;
output c0444;
output c225;
output c5475;
output c5489;
output c0485;
output c9458;
output c151;
output c7179;
output c3432;
output c370;
output c6351;
output c897;
output c8263;
output c1379;
output c564;
output c5251;
output c5148;
output c6400;
output c4252;
output c0211;
output c3413;
output c214;
output c235;
output c0233;
output c8210;
output c1227;
output c4311;
output c7284;
output c1430;
output c5456;
output c741;
output c4251;
output c330;
output c2116;
output c860;
output c6362;
output c029;
output c352;
output c8398;
output c127;
output c363;
output c6115;
output c0102;
output c7339;
output c3201;
output c8315;
output c9498;
output c368;
output c1179;
output c4199;
output c344;
output c2309;
output c7451;
output c1351;
output c5407;
output c3472;
output c0224;
output c9188;
output c124;
output c1250;
output c393;
output c7317;
output c1260;
output c5399;
output c148;
output c2382;
output c7238;
output c8213;
output c2399;
output c7438;
output c3105;
output c9240;
output c5343;
output c9208;
output c6225;
output c6487;
output c6474;
output c7281;
output c0332;
output c2286;
output c220;
output c1357;
output c0194;
output c2305;
output c1422;
output c8391;
output c1323;
output c8205;
output c8361;
output c6433;
output c5325;
output c1319;
output c6177;
output c8158;
output c6157;
output c6109;
output c297;
output c5213;
output c771;
output c9487;
output c8219;
output c1408;
output c4184;
output c8214;
output c854;
output c281;
output c217;
output c670;
output c328;
output c043;
output c2168;
output c424;
output c2387;
output c1107;
output c4465;
output c5232;
output c5225;
output c178;
output c3493;
output c9423;
output c638;
output c9425;
output c0431;
output c183;
output c5154;
output c2113;
output c269;
output c8364;
output c6251;
output c437;
output c6152;
output c2324;
output c390;
output c4133;
output c7107;
output c9445;
output c3224;
output c9482;
output c0377;
output c9383;
output c6165;
output c3250;
output c2405;
output c4477;
output c5438;
output c4171;
output c55;
output c0422;
output c9479;
output c9413;
output c1424;
output c5320;
output c3167;
output c4264;
output c4471;
output c2456;
output c6344;
output c9246;
output c6256;
output c7251;
output c7391;
output c8142;
output c7232;
output c1170;
output c35;
output c8383;
output c230;
output c2125;
output c6472;
output c2335;
output c6385;
output c12;
output c7237;
output c325;
output c6135;
output c9228;
output c1361;
output c9457;
output c1218;
output c6457;
output c2266;
output c5466;
output c579;
output c8150;
output c4463;
output c1325;
output c0499;
output c799;
output c8458;
output c0347;
output c2213;
output c542;
output c999;
output c6279;
output c2489;
output c465;
output c372;
output c7192;
output c7263;
output c654;
output c3291;
output c535;
output c631;
output c2378;
output c3179;
output c282;
output c7249;
output c0169;
output c0372;
output c256;
output c8119;
output c5111;
output c6175;
output c2497;
output c1293;
output c4254;
output c6203;
output c2463;
output c2347;
output c4201;
output c8272;
output c9154;
output c3475;
output c8303;
output c80;
output c326;
output c3412;
output c9118;
output c0193;
output c4458;
output c1157;
output c940;
output c7302;
output c851;
output c318;
output c7309;
output c343;
output c7167;
output c4347;
output c1233;
output c1295;
output c4462;
output c8126;
output c8293;
output c1292;
output c5195;
output c584;
output c4296;
output c6234;
output c5386;
output c8149;
output c4324;
output c1215;
output c8425;
output c2413;
output c5103;
output c9355;
output c048;
output c337;
output c7188;
output c8220;
output c4167;
output c6392;
output c4155;
output c5397;
output c8409;
output c5235;
output c6150;
output c5395;
output c1337;
output c7156;
output c3495;
output c6410;
output c4384;
output c0104;
output c2421;
output c4479;
output c8349;
output c8196;
output c5278;
output c0469;
output c9397;
output c7322;
output c2478;
output c4469;
output c2170;
output c3437;
output c2153;
output c3496;
output c8375;
output c6335;
output c6315;
output c9127;
output c5414;
output c996;
output c781;
output c0190;
output c9106;
output c7401;
output c0359;
output c2245;
output c4248;
output c4299;
output c672;
output c6194;
output c6120;
output c227;
output c1307;
output c4451;
output c9280;
output c3442;
output c3217;
output c027;
output c2325;
output c723;
output c5227;
output c6337;
output c3223;
output c845;
output c4115;
output c2264;
output c4332;
output c3237;
output c0247;
output c1226;
output c6104;
output c9468;
output c550;
output c5429;
output c054;
output c7129;
output c4464;
output c6415;
output c192;
output c010;
output c388;
output c9215;
output c159;
output c7463;
output c5331;
output c2374;
output c9239;
output c419;
output c267;
output c032;
output c4448;
output c4497;
output c0146;
output c0291;
output c038;
output c0305;
output c9259;
output c9496;
output c3206;
output c664;
output c8368;
output c0395;
output c10;
output c3311;
output c7170;
output c3487;
output c688;
output c6284;
output c0346;
output c8369;
output c2131;
output c6191;
output c1365;
output c2285;
output c2316;
output c216;
output c6342;
output c9421;
output c2284;
output c7394;
output c499;
output c4180;
output c0464;
output c0273;
output c2337;
output c08;
output c270;
output c2253;
output c2158;
output c4207;
output c8348;
output c2209;
output c3208;
output c5295;
output c0150;
output c3316;
output c4181;
output c11;
output c7482;
output c988;
output c0179;
output c2407;
output c332;
output c6404;
output c4305;
output c8482;
output c6453;
output c7379;
output c898;
output c870;
output c5355;
output c1115;
output c5387;
output c0443;
output c3295;
output c0197;
output c7437;
output c2130;
output c3134;
output c0203;
output c6398;
output c6300;
output c9150;
output c0411;
output c2323;
output c2257;
output c1158;
output c2140;
output c7354;
output c472;
output c7262;
output c7260;
output c2272;
output c3100;
output c9351;
output c9431;
output c3406;
output c57;
output c7243;
output c0301;
output c8358;
output c6149;
output c8117;
output c6164;
output c1184;
output c3440;
output c7144;
output c758;
output c7497;
output c978;
output c580;
output c7293;
output c8408;
output c314;
output c2167;
output c9437;
output c4165;
output c3346;
output c4303;
output c4294;
output c7189;
output c8339;
output c1198;
output c680;
output c9480;
output c0336;
output c228;
output c6393;
output c0290;
output c2373;
output c463;
output c369;
output c7268;
output c8100;
output c4278;
output c9202;
output c6448;
output c630;
output c9272;
output c8417;
output c1169;
output c2451;
output c3302;
output c9424;
output c3388;
output c541;
output c847;
output c4156;
output c565;
output c2365;
output c4350;
output c9339;
output c386;
output c646;
output c8249;
output c2350;
output c874;
output c8209;
output c3123;
output c6329;
output c19;
output c4274;
output c4188;
output c5267;
output c2191;
output c1409;
output c6471;
output c1354;
output c7199;
output c9312;
output c6405;
output c3309;
output c1278;
output c198;
output c5496;
output c4123;
output c9439;
output c0225;
output c6354;
output c0238;
output c958;
output c5253;
output c2232;
output c1434;
output c27;
output c1266;
output c355;
output c7312;
output c5440;
output c9420;
output c30;
output c5472;
output c919;
output c3430;
output c8380;
output c2480;
output c0166;
output c6358;
output c6193;
output c1288;
output c716;
output c1135;
output c3293;
output c6481;
output c5207;
output c3292;
output c6226;
output c5330;
output c7405;
output c7313;
output c5313;
output c5481;
output c0361;
output c1458;
output c2226;
output c5206;
output c123;
output c4310;
output c581;
output c8424;
output c311;
output c3161;
output c1331;
output c222;
output c2212;
output c4457;
output c058;
output c1297;
output c2171;
output c8461;
output c2388;
output c2231;
output c7212;
output c8137;
output c0380;
output c528;
output c4258;

assign c00 =  x339 &  x367 &  x472 &  x480 & ~x14;
assign c02 =  x285 &  x313 &  x684 &  x739 &  x749 & ~x2 & ~x362;
assign c04 =  x215 & ~x50 & ~x273 & ~x278 & ~x356 & ~x592;
assign c06 = ~x494 & ~x510 & ~x525 & ~x581 & ~x750;
assign c08 =  x764 & ~x21 & ~x61 & ~x388 & ~x478 & ~x667;
assign c010 = ~x13 & ~x15 & ~x22 & ~x23 & ~x40 & ~x42 & ~x140 & ~x170 & ~x336 & ~x391 & ~x415 & ~x416 & ~x451 & ~x472 & ~x478 & ~x536 & ~x584 & ~x612 & ~x620 & ~x674 & ~x761 & ~x773;
assign c012 =  x343 &  x651 &  x679 &  x733 &  x735 & ~x13;
assign c014 =  x199 & ~x224 & ~x392;
assign c016 =  x271 &  x489 & ~x52 & ~x252 & ~x508 & ~x534 & ~x557 & ~x563 & ~x619 & ~x641 & ~x646 & ~x734 & ~x758 & ~x766 & ~x768;
assign c018 =  x143;
assign c020 =  x269 &  x317 &  x658 & ~x388 & ~x750;
assign c022 =  x454 &  x679 & ~x40 & ~x279 & ~x337;
assign c024 = ~x307 & ~x438 & ~x494 & ~x525 & ~x559 & ~x582 & ~x694 & ~x750 & ~x758 & ~x762;
assign c026 =  x303 &  x369 &  x721;
assign c028 =  x241 &  x317 &  x461 &  x517 &  x541 &  x546 &  x574 &  x600 &  x606 &  x630 & ~x7 & ~x53 & ~x54 & ~x392 & ~x555 & ~x582 & ~x588 & ~x725 & ~x774;
assign c030 = ~x525 & ~x538 & ~x550 & ~x555 & ~x576 & ~x580 & ~x581;
assign c032 =  x44 &  x162 &  x239 &  x737 & ~x1 & ~x5 & ~x22 & ~x23 & ~x54 & ~x109 & ~x167 & ~x196 & ~x225 & ~x253 & ~x278 & ~x279 & ~x365 & ~x474 & ~x507 & ~x557 & ~x562 & ~x581 & ~x587 & ~x593 & ~x609 & ~x613 & ~x618 & ~x642 & ~x670 & ~x673 & ~x694;
assign c034 =  x220 &  x248 & ~x308 & ~x392;
assign c036 =  x274 & ~x1 & ~x55 & ~x113 & ~x138 & ~x199 & ~x253 & ~x333 & ~x445 & ~x505 & ~x509 & ~x557 & ~x592 & ~x620 & ~x621 & ~x670 & ~x706 & ~x725 & ~x750;
assign c038 =  x624 &  x767 &  x769 &  x770 &  x772 & ~x145 & ~x200 & ~x370;
assign c040 = ~x409 & ~x438 & ~x477 & ~x523 & ~x649 & ~x668 & ~x750;
assign c042 =  x214 &  x624 & ~x4 & ~x276 & ~x304 & ~x413 & ~x496 & ~x592 & ~x612 & ~x613;
assign c044 =  x243 &  x518 &  x662 &  x693 &  x721 & ~x23 & ~x58 & ~x167 & ~x363 & ~x394 & ~x565 & ~x612;
assign c046 = ~x114 & ~x196 & ~x333 & ~x391 & ~x453 & ~x455 & ~x510 & ~x554 & ~x592 & ~x594 & ~x612 & ~x670 & ~x702 & ~x709 & ~x735;
assign c048 =  x48 & ~x54 & ~x335 & ~x592 & ~x670 & ~x721;
assign c050 = ~x353 & ~x438 & ~x495 & ~x555 & ~x750;
assign c052 =  x42 &  x218 &  x285 &  x286 & ~x6 & ~x22 & ~x23 & ~x78 & ~x107 & ~x109 & ~x363 & ~x419 & ~x562 & ~x638;
assign c054 = ~x94 & ~x128 & ~x160 & ~x188 & ~x219 & ~x477 & ~x497 & ~x535 & ~x750 & ~x754;
assign c056 =  x162 &  x382 &  x547 &  x632 & ~x1 & ~x19 & ~x22 & ~x23 & ~x54 & ~x81 & ~x113 & ~x115 & ~x140 & ~x170 & ~x196 & ~x362 & ~x364 & ~x393 & ~x446 & ~x447 & ~x454 & ~x510 & ~x534 & ~x538 & ~x584 & ~x613 & ~x614 & ~x617 & ~x621 & ~x622 & ~x639 & ~x649 & ~x672 & ~x698 & ~x731 & ~x761 & ~x762 & ~x781 & ~x783;
assign c058 = ~x23 & ~x85 & ~x326 & ~x392 & ~x409 & ~x438 & ~x532 & ~x592 & ~x648 & ~x750 & ~x762 & ~x781;
assign c060 =  x748 & ~x104;
assign c062 =  x227 & ~x23 & ~x54 & ~x167 & ~x364 & ~x756;
assign c064 =  x624 & ~x24 & ~x53 & ~x254 & ~x335 & ~x391 & ~x424 & ~x445 & ~x477 & ~x592 & ~x612 & ~x670 & ~x676 & ~x727 & ~x766 & ~x767 & ~x769 & ~x782;
assign c066 = ~x497 & ~x513 & ~x581 & ~x626;
assign c068 =  x326 &  x405 &  x625 &  x657 & ~x60 & ~x109 & ~x137 & ~x308 & ~x455 & ~x511;
assign c070 =  x764 & ~x10 & ~x167 & ~x528;
assign c072 =  x118 &  x173 &  x201 &  x229 &  x288 &  x630 &  x715 & ~x22 & ~x392 & ~x445 & ~x478 & ~x649;
assign c074 = ~x432 & ~x511 & ~x655;
assign c076 =  x289 &  x351 & ~x30 & ~x119 & ~x167 & ~x175 & ~x195 & ~x385 & ~x506 & ~x592 & ~x642 & ~x648 & ~x703 & ~x705 & ~x781;
assign c078 =  x651 &  x678 &  x679 &  x708 &  x735 & ~x2 & ~x15 & ~x645;
assign c080 =  x243 &  x317 &  x460 &  x577 &  x578 &  x713 & ~x142 & ~x356 & ~x394 & ~x694 & ~x727;
assign c082 = ~x129 & ~x413 & ~x441 & ~x471 & ~x594 & ~x772;
assign c084 =  x200 &  x229 &  x247 &  x256 &  x274 &  x276 & ~x4;
assign c086 = ~x371 & ~x454 & ~x459 & ~x497 & ~x554 & ~x734 & ~x759;
assign c088 =  x255 & ~x7 & ~x55 & ~x771;
assign c090 = ~x650 & ~x655 & ~x709 & ~x738 & ~x767 & ~x769;
assign c092 =  x191 &  x219 &  x302 & ~x28 & ~x278 & ~x309 & ~x365 & ~x392 & ~x422 & ~x479 & ~x533 & ~x644 & ~x755;
assign c094 =  x243 &  x263 &  x628 &  x631 &  x658 &  x685 &  x720 & ~x89 & ~x117 & ~x218 & ~x304 & ~x311 & ~x762;
assign c096 =  x607 & ~x188 & ~x412;
assign c098 =  x214 &  x233 &  x603 &  x625 &  x658 & ~x91 & ~x413;
assign c0100 =  x214 &  x266 &  x290 &  x401 &  x407 &  x489 &  x541 &  x545 &  x546 &  x597 &  x600 &  x684 &  x713 & ~x142 & ~x278 & ~x336 & ~x395 & ~x440 & ~x477 & ~x502 & ~x611 & ~x617 & ~x673;
assign c0102 =  x42 &  x288 &  x685 &  x765 &  x769 & ~x454 & ~x498;
assign c0104 = ~x5 & ~x19 & ~x180 & ~x361 & ~x413 & ~x455 & ~x581 & ~x592 & ~x610 & ~x638 & ~x704 & ~x750 & ~x754;
assign c0106 =  x339 &  x367 &  x369;
assign c0108 = ~x93 & ~x160 & ~x357 & ~x454 & ~x554 & ~x555 & ~x586 & ~x655;
assign c0110 =  x247 &  x598 & ~x283 & ~x394 & ~x650 & ~x668 & ~x697 & ~x754;
assign c0112 =  x40 &  x134 & ~x5 & ~x24 & ~x27 & ~x54 & ~x55 & ~x57 & ~x86 & ~x139 & ~x141 & ~x143 & ~x165 & ~x196 & ~x222 & ~x251 & ~x392 & ~x394 & ~x416 & ~x426 & ~x445 & ~x453 & ~x454 & ~x471 & ~x476 & ~x500 & ~x501 & ~x508 & ~x510 & ~x535 & ~x561 & ~x583 & ~x586 & ~x590 & ~x592 & ~x594 & ~x611 & ~x612 & ~x617 & ~x621 & ~x644 & ~x670 & ~x699 & ~x702 & ~x704 & ~x725 & ~x728 & ~x750 & ~x760;
assign c0114 =  x146 & ~x471 & ~x472 & ~x767;
assign c0116 =  x219 &  x228 &  x285 & ~x37 & ~x769;
assign c0118 = ~x223 & ~x464 & ~x494 & ~x549;
assign c0120 = ~x93 & ~x129 & ~x130 & ~x308 & ~x361 & ~x385 & ~x415 & ~x525 & ~x554 & ~x566;
assign c0122 = ~x377 & ~x606 & ~x676;
assign c0124 = ~x94 & ~x445 & ~x565 & ~x602 & ~x604 & ~x605 & ~x638;
assign c0126 =  x18 & ~x29 & ~x338 & ~x367 & ~x502 & ~x613 & ~x670 & ~x677 & ~x723 & ~x756 & ~x774;
assign c0128 = ~x130 & ~x510 & ~x603 & ~x604 & ~x605;
assign c0130 =  x229 &  x274 &  x605 & ~x390 & ~x508 & ~x510 & ~x724;
assign c0132 =  x339 &  x359 &  x367 & ~x28;
assign c0134 =  x260 &  x288 &  x434 &  x517 &  x595 &  x629 &  x651 & ~x13 & ~x52 & ~x118 & ~x392 & ~x781;
assign c0136 =  x158 &  x624 &  x628 &  x678 &  x679 & ~x11 & ~x169 & ~x555 & ~x730 & ~x756;
assign c0138 = ~x371 & ~x597;
assign c0140 =  x246 &  x340 & ~x336 & ~x640 & ~x750;
assign c0142 =  x17 &  x233 &  x624 &  x769 &  x772 & ~x731;
assign c0144 =  x108;
assign c0146 =  x215 &  x270 &  x692 & ~x161 & ~x173 & ~x230 & ~x537 & ~x559 & ~x761;
assign c0148 =  x108;
assign c0150 =  x200 &  x201 &  x246 &  x257 &  x285 & ~x612;
assign c0152 =  x289 &  x574 &  x597 &  x602 &  x624 &  x628 & ~x28 & ~x51 & ~x116 & ~x337 & ~x649 & ~x703;
assign c0154 = ~x413 & ~x711 & ~x714 & ~x768;
assign c0156 =  x625 &  x687 &  x716 &  x741 &  x767 &  x769 &  x770 &  x771 &  x772 & ~x6 & ~x25 & ~x61 & ~x141 & ~x199 & ~x308 & ~x334 & ~x335 & ~x337 & ~x338 & ~x360 & ~x361 & ~x391 & ~x394 & ~x413 & ~x424 & ~x472 & ~x499 & ~x500 & ~x508 & ~x556 & ~x558 & ~x584 & ~x590 & ~x594 & ~x617 & ~x644 & ~x678 & ~x781;
assign c0158 = ~x93 & ~x512 & ~x713 & ~x766;
assign c0160 =  x78 &  x107 &  x220 & ~x112 & ~x224 & ~x308 & ~x671 & ~x700 & ~x726;
assign c0162 = ~x456 & ~x485 & ~x627 & ~x750;
assign c0164 =  x164 & ~x364;
assign c0166 =  x121 &  x243 &  x261 &  x314 &  x413 &  x497 &  x568 &  x609 &  x623 &  x624 &  x708 &  x748 &  x749 & ~x24 & ~x57 & ~x391 & ~x587;
assign c0168 =  x242 &  x540 &  x658 &  x708 &  x735 &  x737 &  x763 & ~x392 & ~x448 & ~x759;
assign c0170 =  x289 &  x317 &  x319 &  x346 &  x373 &  x458 &  x488 &  x489 &  x517 &  x543 &  x598 &  x601 &  x603 &  x624 &  x629 &  x632 &  x652 &  x658 &  x715 &  x744 & ~x1 & ~x13 & ~x23 & ~x29 & ~x80 & ~x111 & ~x219 & ~x255 & ~x283 & ~x284 & ~x394 & ~x395 & ~x396 & ~x397 & ~x448 & ~x504 & ~x562 & ~x564 & ~x592 & ~x611 & ~x639 & ~x668;
assign c0172 = ~x119 & ~x211 & ~x426 & ~x454 & ~x472 & ~x511 & ~x555 & ~x705;
assign c0174 =  x368 &  x396 &  x452 &  x623 &  x624 & ~x13;
assign c0176 =  x220 &  x637 &  x665 & ~x337 & ~x392;
assign c0178 = ~x413 & ~x471 & ~x472 & ~x655;
assign c0180 = ~x23 & ~x51 & ~x53 & ~x80 & ~x81 & ~x88 & ~x136 & ~x180 & ~x226 & ~x282 & ~x335 & ~x388 & ~x392 & ~x413 & ~x441 & ~x442 & ~x453 & ~x454 & ~x471 & ~x477 & ~x482 & ~x507 & ~x510 & ~x538 & ~x554 & ~x561 & ~x581 & ~x582 & ~x617 & ~x642 & ~x670 & ~x676 & ~x698 & ~x701 & ~x704 & ~x729 & ~x750 & ~x754 & ~x759 & ~x762 & ~x777;
assign c0182 =  x274 & ~x19 & ~x23 & ~x221 & ~x445 & ~x469 & ~x508 & ~x525 & ~x566 & ~x609 & ~x749;
assign c0184 = ~x445 & ~x455 & ~x626 & ~x627 & ~x650 & ~x681;
assign c0186 =  x70 &  x77 & ~x29 & ~x61 & ~x142 & ~x284 & ~x308 & ~x421 & ~x508 & ~x592 & ~x676;
assign c0188 =  x371 &  x595 &  x651 &  x679 &  x708 & ~x40 & ~x223;
assign c0190 =  x143;
assign c0192 =  x44 &  x173 &  x201 &  x257 & ~x7 & ~x88 & ~x311 & ~x648 & ~x728 & ~x749;
assign c0194 =  x9 &  x215 &  x243 &  x289 &  x434 &  x518 &  x547 &  x598 &  x599 &  x601 &  x602 &  x624 &  x630 & ~x308 & ~x388 & ~x592;
assign c0196 = ~x93 & ~x102 & ~x104 & ~x413 & ~x455;
assign c0198 =  x652 &  x681 &  x769 &  x770 &  x771 & ~x191;
assign c0200 =  x243 &  x465 &  x489 &  x546 &  x574 &  x596 &  x597 &  x658 &  x686 &  x713 &  x745 & ~x171 & ~x173 & ~x611 & ~x695 & ~x762;
assign c0202 = ~x14 & ~x412 & ~x714 & ~x766 & ~x767;
assign c0204 = ~x67 & ~x129 & ~x371 & ~x455;
assign c0206 =  x241 &  x262 &  x268 &  x290 &  x317 &  x374 &  x431 &  x460 &  x486 &  x574 &  x597 &  x598 & ~x34 & ~x84 & ~x114 & ~x141 & ~x220 & ~x250 & ~x307 & ~x357 & ~x369 & ~x413 & ~x422 & ~x441 & ~x554 & ~x556 & ~x592 & ~x617 & ~x721 & ~x755 & ~x756;
assign c0208 =  x47 &  x651 &  x715 &  x746 & ~x13 & ~x303;
assign c0210 =  x215 &  x233 &  x461 &  x518 &  x603 &  x658 & ~x145 & ~x342 & ~x589 & ~x592;
assign c0212 =  x485 &  x574 &  x597 &  x628 &  x743 & ~x88 & ~x107 & ~x194 & ~x253 & ~x284 & ~x370 & ~x413 & ~x417 & ~x469 & ~x511 & ~x527 & ~x566 & ~x638 & ~x650 & ~x668 & ~x704 & ~x727 & ~x749 & ~x754;
assign c0214 =  x17 & ~x25 & ~x54 & ~x79 & ~x389 & ~x392 & ~x419 & ~x448 & ~x472 & ~x478 & ~x554 & ~x581 & ~x592 & ~x614 & ~x620 & ~x667 & ~x668 & ~x676 & ~x696 & ~x698 & ~x723 & ~x753;
assign c0216 =  x338 &  x339;
assign c0218 =  x117 &  x369 &  x735;
assign c0220 = ~x93 & ~x153 & ~x193 & ~x441 & ~x471 & ~x472 & ~x525 & ~x640 & ~x706;
assign c0222 = ~x130 & ~x156 & ~x370 & ~x413 & ~x440 & ~x441 & ~x468 & ~x510 & ~x563 & ~x565 & ~x649;
assign c0224 =  x105 &  x243 &  x708 &  x735 &  x769 &  x771;
assign c0226 = ~x354 & ~x371 & ~x379 & ~x494;
assign c0228 =  x77 & ~x7 & ~x22 & ~x87 & ~x445 & ~x448 & ~x473 & ~x534 & ~x584 & ~x592 & ~x594 & ~x615 & ~x754;
assign c0230 =  x369 &  x452 &  x735 &  x749;
assign c0232 =  x76 & ~x413 & ~x581 & ~x774;
assign c0234 =  x242 &  x266 &  x513 &  x570 &  x602 &  x603 &  x631 &  x635 &  x657 &  x770 & ~x22 & ~x23 & ~x91 & ~x167 & ~x304 & ~x449 & ~x455 & ~x476 & ~x595 & ~x670;
assign c0236 =  x212 &  x214 &  x233 &  x242 &  x264 &  x271 &  x434 &  x460 &  x461 &  x485 &  x488 &  x518 &  x547 &  x575 &  x603 &  x606 &  x635 & ~x22 & ~x56 & ~x114 & ~x167 & ~x192 & ~x248 & ~x254 & ~x309 & ~x419 & ~x448 & ~x455 & ~x613 & ~x615 & ~x701;
assign c0238 = ~x463 & ~x597 & ~x733;
assign c0240 =  x63 & ~x3 & ~x7 & ~x29 & ~x58 & ~x86 & ~x87 & ~x88 & ~x112 & ~x166 & ~x224 & ~x309 & ~x370 & ~x413 & ~x448 & ~x474 & ~x497 & ~x500 & ~x558 & ~x582 & ~x586 & ~x618 & ~x621 & ~x639 & ~x642 & ~x643 & ~x644 & ~x694 & ~x728 & ~x779;
assign c0242 =  x173 &  x201 &  x597 & ~x220 & ~x617 & ~x637 & ~x674 & ~x721 & ~x750 & ~x754;
assign c0244 =  x285 &  x312 &  x340 &  x415 & ~x16;
assign c0246 =  x430 & ~x5 & ~x23 & ~x55 & ~x87 & ~x107 & ~x113 & ~x165 & ~x193 & ~x222 & ~x249 & ~x250 & ~x306 & ~x311 & ~x313 & ~x340 & ~x358 & ~x370 & ~x388 & ~x398 & ~x420 & ~x503 & ~x525 & ~x531 & ~x532 & ~x537 & ~x561 & ~x581 & ~x584 & ~x591 & ~x592 & ~x594 & ~x609 & ~x611 & ~x615 & ~x617 & ~x668 & ~x675 & ~x676 & ~x698 & ~x700 & ~x704 & ~x705 & ~x733 & ~x750 & ~x761 & ~x774 & ~x779 & ~x783;
assign c0248 =  x457 &  x574 &  x603 &  x652 &  x658 & ~x119 & ~x167 & ~x667 & ~x726 & ~x733 & ~x749;
assign c0250 = ~x211 & ~x212 & ~x399 & ~x413 & ~x475 & ~x554;
assign c0252 =  x274 & ~x7 & ~x23 & ~x85 & ~x280 & ~x472 & ~x504 & ~x557 & ~x561 & ~x566 & ~x642 & ~x648 & ~x650 & ~x695 & ~x701 & ~x704 & ~x721 & ~x750 & ~x756 & ~x780;
assign c0254 =  x9 &  x215 &  x624 &  x625 &  x629;
assign c0256 = ~x54 & ~x74 & ~x81 & ~x93 & ~x104 & ~x114 & ~x125 & ~x128 & ~x162 & ~x170 & ~x307 & ~x335 & ~x503 & ~x507 & ~x535 & ~x563 & ~x583 & ~x584 & ~x589 & ~x617 & ~x620 & ~x641 & ~x642 & ~x754 & ~x757 & ~x781 & ~x782;
assign c0258 =  x118 & ~x23 & ~x28 & ~x59 & ~x79 & ~x81 & ~x88 & ~x109 & ~x166 & ~x167 & ~x168 & ~x195 & ~x225 & ~x251 & ~x282 & ~x305 & ~x309 & ~x336 & ~x361 & ~x415 & ~x426 & ~x501 & ~x510 & ~x559 & ~x561 & ~x564 & ~x584 & ~x592 & ~x593 & ~x618 & ~x622 & ~x649 & ~x668 & ~x670 & ~x693 & ~x727 & ~x750 & ~x777 & ~x778;
assign c0260 =  x204 &  x233 &  x624 &  x763 & ~x110 & ~x141 & ~x449 & ~x559 & ~x588 & ~x642;
assign c0262 = ~x412 & ~x413 & ~x426 & ~x554 & ~x705 & ~x766 & ~x767 & ~x771 & ~x772 & ~x777;
assign c0264 =  x567 &  x679 & ~x13 & ~x15 & ~x16 & ~x29 & ~x40 & ~x41 & ~x54 & ~x57 & ~x618 & ~x754;
assign c0266 =  x289 &  x380 & ~x13 & ~x42 & ~x146 & ~x194 & ~x197 & ~x256 & ~x308 & ~x450 & ~x505 & ~x561 & ~x617 & ~x759;
assign c0268 = ~x168 & ~x365 & ~x383 & ~x411 & ~x438 & ~x494 & ~x551;
assign c0270 =  x262 &  x351 &  x431 &  x602 &  x629 &  x657 & ~x252 & ~x312 & ~x338 & ~x412 & ~x468 & ~x586 & ~x592 & ~x594 & ~x615 & ~x646 & ~x750 & ~x762;
assign c0272 =  x76 &  x105 &  x133 &  x162 & ~x416 & ~x445 & ~x693 & ~x754;
assign c0274 =  x679 &  x734 &  x748 & ~x13 & ~x505;
assign c0276 =  x764 &  x765 &  x767 &  x769 & ~x167 & ~x397 & ~x611 & ~x703 & ~x754;
assign c0278 = ~x29 & ~x61 & ~x74 & ~x93 & ~x120 & ~x128 & ~x130 & ~x426 & ~x445 & ~x454 & ~x510;
assign c0280 =  x158 &  x212 &  x326 &  x433 &  x490 &  x578 &  x597 &  x658 & ~x55 & ~x562 & ~x609 & ~x723 & ~x733 & ~x774;
assign c0282 =  x214 &  x215 &  x353 &  x429 &  x485 &  x568 & ~x15 & ~x302 & ~x391 & ~x555 & ~x585;
assign c0284 =  x97 &  x126 &  x242 &  x243 &  x257 &  x285 &  x331 &  x369 &  x460 &  x601 & ~x779;
assign c0286 =  x349 &  x597 & ~x34 & ~x83 & ~x84 & ~x167 & ~x222 & ~x311 & ~x335 & ~x371 & ~x385 & ~x413 & ~x422 & ~x441 & ~x530 & ~x555 & ~x561 & ~x706 & ~x721 & ~x727 & ~x733 & ~x735;
assign c0288 =  x42 &  x70 &  x233 &  x603 &  x770 &  x771 &  x772 & ~x511 & ~x594;
assign c0290 =  x227 & ~x48 & ~x759;
assign c0292 =  x178 &  x597 &  x598 &  x601 & ~x112 & ~x114 & ~x195 & ~x361 & ~x371 & ~x413 & ~x477 & ~x532 & ~x590 & ~x641 & ~x707 & ~x735 & ~x750;
assign c0294 =  x233 &  x769 & ~x170 & ~x356 & ~x455;
assign c0296 =  x226;
assign c0298 =  x107 & ~x306 & ~x647 & ~x781;
assign c0300 =  x164;
assign c0302 =  x214 &  x297 &  x488 &  x602 &  x603 & ~x20 & ~x60 & ~x87 & ~x107 & ~x111 & ~x119 & ~x144 & ~x166 & ~x171 & ~x173 & ~x219 & ~x226 & ~x336 & ~x343 & ~x371 & ~x420 & ~x483 & ~x504 & ~x562 & ~x565 & ~x613 & ~x619 & ~x667 & ~x669 & ~x705 & ~x728 & ~x753 & ~x761;
assign c0304 = ~x320 & ~x455 & ~x513 & ~x597;
assign c0306 =  x288 &  x289 &  x658 & ~x280 & ~x284 & ~x310 & ~x455 & ~x726;
assign c0308 = ~x93 & ~x94 & ~x120 & ~x128 & ~x413 & ~x705;
assign c0310 =  x765 &  x769 &  x771 &  x775 & ~x37 & ~x336;
assign c0312 = ~x371 & ~x597 & ~x684;
assign c0314 =  x226;
assign c0316 =  x256 &  x258 & ~x5 & ~x24 & ~x61 & ~x112 & ~x642 & ~x761 & ~x781;
assign c0318 =  x76 &  x105 &  x375 &  x624 &  x685 &  x770 &  x771 & ~x392 & ~x705;
assign c0320 = ~x441 & ~x482 & ~x512 & ~x516 & ~x517;
assign c0322 =  x136;
assign c0324 = ~x212 & ~x238 & ~x413 & ~x566 & ~x592 & ~x721 & ~x749 & ~x759;
assign c0326 =  x651 &  x679 & ~x334 & ~x384 & ~x440 & ~x504;
assign c0328 =  x430 &  x568 &  x625 &  x678 &  x680 &  x706 &  x708 &  x735 & ~x13 & ~x170 & ~x224 & ~x589;
assign c0330 =  x78 & ~x23 & ~x57 & ~x170 & ~x251 & ~x255 & ~x391 & ~x417 & ~x423 & ~x450 & ~x451 & ~x473 & ~x475 & ~x505 & ~x561 & ~x700 & ~x724 & ~x752 & ~x759 & ~x782;
assign c0332 =  x162 &  x471 &  x749;
assign c0334 = ~x127 & ~x161 & ~x253 & ~x425 & ~x426 & ~x509 & ~x510 & ~x525 & ~x529 & ~x592 & ~x612 & ~x613 & ~x668 & ~x723;
assign c0336 =  x214 &  x321 &  x405 &  x462 &  x485 &  x541 &  x602 &  x624 & ~x1 & ~x22 & ~x79 & ~x112 & ~x531 & ~x731 & ~x749;
assign c0338 =  x200 &  x202 & ~x1 & ~x19 & ~x22 & ~x23 & ~x167 & ~x336 & ~x622;
assign c0340 = ~x114 & ~x492 & ~x495 & ~x510 & ~x694 & ~x750 & ~x762;
assign c0342 =  x184 &  x205 &  x233 &  x261 &  x263 &  x289 &  x317 &  x630 & ~x22 & ~x23 & ~x52 & ~x142 & ~x283 & ~x311 & ~x455 & ~x539 & ~x695 & ~x734;
assign c0344 =  x105 &  x129 &  x133 &  x160 & ~x5 & ~x304 & ~x391 & ~x619 & ~x637 & ~x667 & ~x694 & ~x700 & ~x701 & ~x722 & ~x750;
assign c0346 =  x268 &  x326 &  x461 &  x487 &  x573 &  x629 & ~x4 & ~x55 & ~x56 & ~x60 & ~x284 & ~x455 & ~x511 & ~x555 & ~x558 & ~x721 & ~x750;
assign c0348 = ~x463 & ~x604 & ~x657 & ~x658 & ~x686;
assign c0350 =  x248 & ~x0 & ~x1 & ~x2 & ~x61 & ~x280 & ~x531 & ~x673 & ~x783;
assign c0352 = ~x150 & ~x440 & ~x510 & ~x750;
assign c0354 =  x77 &  x78 & ~x254 & ~x391 & ~x448 & ~x479 & ~x759;
assign c0356 =  x255 & ~x772;
assign c0358 =  x69 &  x233 &  x271 &  x327 &  x489 &  x547 &  x574 &  x575 & ~x441;
assign c0360 = ~x354 & ~x355 & ~x384 & ~x412 & ~x494;
assign c0362 =  x15 &  x134 &  x219 &  x229;
assign c0364 = ~x74 & ~x92 & ~x102 & ~x129 & ~x357 & ~x413;
assign c0366 =  x215 &  x316 &  x624 &  x683 &  x735 &  x765 &  x769;
assign c0368 =  x132 & ~x377;
assign c0370 = ~x178 & ~x413 & ~x472 & ~x497 & ~x525 & ~x637 & ~x750;
assign c0372 =  x310;
assign c0374 = ~x102 & ~x111 & ~x120 & ~x139 & ~x142 & ~x156 & ~x158 & ~x165 & ~x193 & ~x388 & ~x503 & ~x581 & ~x592 & ~x621 & ~x749 & ~x782;
assign c0376 = ~x224 & ~x238 & ~x371 & ~x597 & ~x622;
assign c0378 = ~x566 & ~x574 & ~x713;
assign c0380 = ~x29 & ~x388 & ~x400 & ~x446 & ~x455 & ~x538 & ~x557 & ~x766;
assign c0382 =  x317 &  x345 &  x597 &  x656 & ~x54 & ~x356 & ~x750;
assign c0384 =  x198;
assign c0386 = ~x74 & ~x94 & ~x602 & ~x612;
assign c0388 =  x285 & ~x2 & ~x22 & ~x55 & ~x58 & ~x140 & ~x142 & ~x224 & ~x277 & ~x391 & ~x395 & ~x445 & ~x472 & ~x565 & ~x612 & ~x617 & ~x641 & ~x644 & ~x645 & ~x647 & ~x695 & ~x702 & ~x704 & ~x705 & ~x727;
assign c0390 = ~x492 & ~x494 & ~x603 & ~x604 & ~x605;
assign c0392 =  x143;
assign c0394 =  x650 &  x706 & ~x13 & ~x15 & ~x41 & ~x54 & ~x419 & ~x728;
assign c0396 =  x369 &  x678 & ~x15;
assign c0398 =  x19 & ~x13 & ~x476;
assign c0400 =  x208 &  x426 &  x454 &  x601 &  x679 &  x681 & ~x10 & ~x57 & ~x334;
assign c0402 =  x20;
assign c0404 =  x214 &  x515 &  x546 &  x550 &  x578 &  x597 &  x607 & ~x29 & ~x137 & ~x558 & ~x591 & ~x704 & ~x735 & ~x766;
assign c0406 = ~x440 & ~x603 & ~x605;
assign c0408 = ~x93 & ~x277 & ~x438 & ~x482 & ~x508 & ~x524 & ~x554 & ~x582 & ~x617 & ~x639 & ~x759;
assign c0410 = ~x313 & ~x370 & ~x427 & ~x639 & ~x705 & ~x714 & ~x750 & ~x767 & ~x768;
assign c0412 =  x214 &  x261 &  x317 & ~x13 & ~x147 & ~x282 & ~x337 & ~x472 & ~x753;
assign c0414 =  x71 & ~x0 & ~x8 & ~x21 & ~x25 & ~x27 & ~x50 & ~x55 & ~x59 & ~x82 & ~x87 & ~x109 & ~x141 & ~x169 & ~x170 & ~x193 & ~x195 & ~x196 & ~x253 & ~x282 & ~x308 & ~x334 & ~x341 & ~x342 & ~x360 & ~x361 & ~x368 & ~x394 & ~x396 & ~x398 & ~x413 & ~x414 & ~x421 & ~x425 & ~x426 & ~x441 & ~x442 & ~x445 & ~x448 & ~x449 & ~x454 & ~x455 & ~x481 & ~x500 & ~x509 & ~x510 & ~x511 & ~x525 & ~x527 & ~x533 & ~x555 & ~x565 & ~x566 & ~x593 & ~x594 & ~x609 & ~x614 & ~x637 & ~x645 & ~x646 & ~x648 & ~x649 & ~x695 & ~x696 & ~x706 & ~x721 & ~x724 & ~x727 & ~x728 & ~x729 & ~x733 & ~x750 & ~x751 & ~x758 & ~x761 & ~x762 & ~x777 & ~x781;
assign c0416 =  x229 &  x257 &  x274 &  x285 &  x303 &  x330 &  x358 &  x656 &  x658;
assign c0418 =  x285 &  x313 &  x624 &  x685 &  x735 &  x749 & ~x23;
assign c0420 = ~x379 & ~x525 & ~x578 & ~x583 & ~x750;
assign c0422 =  x70 &  x289 &  x743 &  x771 &  x772 & ~x3 & ~x55 & ~x165 & ~x343 & ~x371 & ~x399 & ~x474 & ~x638 & ~x645 & ~x754;
assign c0424 = ~x343 & ~x511 & ~x637 & ~x766;
assign c0426 =  x191 & ~x7 & ~x29 & ~x54 & ~x280 & ~x306 & ~x308 & ~x336 & ~x397 & ~x426 & ~x474 & ~x557 & ~x561 & ~x562 & ~x563 & ~x592 & ~x612 & ~x622 & ~x649 & ~x667 & ~x706;
assign c0428 =  x243 &  x411 &  x747 &  x769 &  x770 &  x771 & ~x28 & ~x57 & ~x58 & ~x60 & ~x371 & ~x426 & ~x454 & ~x566 & ~x610;
assign c0430 =  x243 &  x658 &  x748 & ~x22 & ~x104 & ~x479;
assign c0432 = ~x455 & ~x625 & ~x627 & ~x681 & ~x738 & ~x750 & ~x771;
assign c0434 = ~x355 & ~x603 & ~x606 & ~x632 & ~x633 & ~x658 & ~x750;
assign c0436 =  x97 &  x241 &  x298 &  x405 &  x493 &  x517 &  x575 &  x601 &  x603 &  x658 & ~x392 & ~x455 & ~x511 & ~x531 & ~x592 & ~x623 & ~x640 & ~x706 & ~x726;
assign c0438 = ~x409 & ~x410 & ~x492 & ~x494 & ~x495;
assign c0440 =  x288 &  x596 &  x597 &  x657 &  x658 &  x714 & ~x57 & ~x108 & ~x277 & ~x391 & ~x581 & ~x614 & ~x618 & ~x731;
assign c0442 = ~x195 & ~x220 & ~x251 & ~x255 & ~x283 & ~x335 & ~x337 & ~x343 & ~x370 & ~x391 & ~x426 & ~x446 & ~x455 & ~x469 & ~x472 & ~x538 & ~x592 & ~x595 & ~x650 & ~x675 & ~x732 & ~x734 & ~x750 & ~x752 & ~x766 & ~x767 & ~x768 & ~x772;
assign c0444 =  x116 &  x144 & ~x23 & ~x645;
assign c0446 =  x317 &  x351 &  x487 &  x708 &  x714 &  x770 &  x771 &  x772 & ~x62 & ~x339;
assign c0448 =  x662 & ~x3 & ~x307 & ~x336 & ~x361 & ~x375 & ~x413 & ~x415 & ~x478 & ~x555 & ~x581 & ~x584 & ~x618 & ~x700 & ~x733;
assign c0450 =  x173 &  x174 &  x201 &  x598 &  x737 & ~x199 & ~x253 & ~x538 & ~x554 & ~x648 & ~x670;
assign c0452 =  x164 & ~x335;
assign c0454 =  x284 & ~x0 & ~x57 & ~x167 & ~x280 & ~x336 & ~x363 & ~x391 & ~x482 & ~x510 & ~x534 & ~x584 & ~x645 & ~x670 & ~x701 & ~x783;
assign c0456 =  x77 & ~x22 & ~x58 & ~x60 & ~x391 & ~x472 & ~x534 & ~x564 & ~x585 & ~x590 & ~x613 & ~x671 & ~x678 & ~x763 & ~x781;
assign c0458 =  x542 &  x595 &  x651 &  x652 &  x679 & ~x13 & ~x40 & ~x41 & ~x671;
assign c0460 =  x199 & ~x167;
assign c0462 =  x98 &  x298 &  x317 &  x430 &  x431 &  x520 &  x545 &  x571 &  x572 &  x573 &  x574 &  x597 &  x598 &  x600 &  x605 &  x632 &  x654 &  x680 &  x681 &  x686 &  x708 &  x711 &  x767 &  x771 &  x772 &  x773 & ~x20 & ~x55 & ~x56 & ~x81 & ~x140 & ~x167 & ~x195 & ~x196 & ~x280 & ~x336 & ~x361 & ~x392 & ~x394 & ~x423 & ~x450 & ~x480 & ~x501 & ~x502 & ~x529 & ~x558 & ~x561 & ~x584 & ~x587 & ~x592 & ~x642 & ~x671 & ~x702 & ~x705 & ~x706 & ~x723 & ~x724 & ~x730 & ~x783;
assign c0464 =  x162 &  x330 &  x665 &  x735 &  x748;
assign c0466 =  x288 &  x764 & ~x21 & ~x58 & ~x85 & ~x170 & ~x223 & ~x337 & ~x500 & ~x555 & ~x621 & ~x696 & ~x724 & ~x731 & ~x780;
assign c0468 =  x679 & ~x5 & ~x22 & ~x25 & ~x31 & ~x193 & ~x280 & ~x384 & ~x412 & ~x420 & ~x505 & ~x532 & ~x586 & ~x702 & ~x723 & ~x759;
assign c0470 =  x274 &  x285 &  x286 &  x314 &  x331 &  x341 &  x359 &  x369 &  x376 &  x415 &  x452 &  x679 &  x685 & ~x559;
assign c0472 =  x304 & ~x20 & ~x29 & ~x87 & ~x88 & ~x166 & ~x196 & ~x564 & ~x617 & ~x677 & ~x702 & ~x727 & ~x779 & ~x780;
assign c0474 =  x136;
assign c0476 = ~x158 & ~x178 & ~x455 & ~x497;
assign c0478 =  x218 & ~x588 & ~x670 & ~x728 & ~x734 & ~x751;
assign c0480 =  x46 &  x47 &  x77 & ~x22 & ~x58 & ~x167 & ~x360 & ~x415 & ~x448 & ~x532 & ~x561 & ~x562 & ~x706;
assign c0482 = ~x19 & ~x53 & ~x92 & ~x160 & ~x283 & ~x413 & ~x455 & ~x468 & ~x499 & ~x526 & ~x529 & ~x585 & ~x695 & ~x760;
assign c0484 = ~x93 & ~x426 & ~x478 & ~x508 & ~x657 & ~x766;
assign c0486 = ~x347 & ~x510 & ~x517 & ~x567 & ~x750;
assign c0488 =  x233 &  x271 &  x289 &  x375 &  x488 &  x596 &  x602 &  x744 & ~x134 & ~x167 & ~x444 & ~x701 & ~x752;
assign c0490 =  x215 & ~x15 & ~x41 & ~x80 & ~x138 & ~x172 & ~x224 & ~x249 & ~x283 & ~x451 & ~x472 & ~x502 & ~x562 & ~x563 & ~x612 & ~x617 & ~x642 & ~x674 & ~x725 & ~x755;
assign c0492 =  x171;
assign c0494 =  x595 &  x651 & ~x15 & ~x40 & ~x41 & ~x505 & ~x617;
assign c0496 =  x430 & ~x21 & ~x28 & ~x160 & ~x284 & ~x416 & ~x422 & ~x425 & ~x426 & ~x427 & ~x447 & ~x511 & ~x584 & ~x614 & ~x621 & ~x695 & ~x750 & ~x764;
assign c0498 =  x454 &  x575 &  x679 &  x706 &  x708 & ~x13 & ~x307;
assign c01 =  x10 &  x38 &  x40 &  x66 &  x67 &  x102 &  x124 &  x184 &  x324 &  x353 &  x432 &  x458 &  x738 & ~x5 & ~x254 & ~x449;
assign c03 =  x404 &  x655 & ~x230 & ~x567 & ~x664 & ~x679 & ~x692;
assign c05 =  x325 & ~x201 & ~x247 & ~x275 & ~x289;
assign c07 =  x195;
assign c09 =  x113;
assign c011 =  x210 &  x217 &  x492 &  x538 &  x566 &  x638 & ~x250;
assign c013 =  x66 &  x67 &  x237 &  x542 &  x739 & ~x312 & ~x623 & ~x677;
assign c015 =  x168;
assign c017 =  x337 &  x470;
assign c019 =  x364;
assign c021 =  x67 &  x72 &  x92 &  x128 & ~x77 & ~x163 & ~x443 & ~x698;
assign c023 = ~x47 & ~x65 & ~x75 & ~x314 & ~x323 & ~x411;
assign c025 =  x307;
assign c027 =  x390;
assign c029 =  x324 &  x711 &  x717 & ~x161 & ~x692;
assign c033 =  x56;
assign c035 =  x503;
assign c037 =  x190 &  x324 &  x356 &  x416 &  x442 &  x470 &  x528;
assign c039 = ~x246 & ~x692 & ~x720 & ~x748;
assign c041 =  x179 &  x267 &  x711 & ~x48 & ~x202 & ~x472 & ~x775;
assign c043 =  x128 &  x156 & ~x203 & ~x244 & ~x300 & ~x444;
assign c045 =  x750 & ~x406;
assign c047 =  x35 &  x49 &  x62 &  x493;
assign c049 =  x564 & ~x95;
assign c051 = ~x48 & ~x232 & ~x243 & ~x244 & ~x288 & ~x415;
assign c053 =  x24;
assign c055 =  x84;
assign c057 =  x29;
assign c059 =  x167;
assign c061 = ~x47 & ~x50 & ~x77 & ~x229 & ~x256 & ~x664 & ~x748;
assign c063 =  x476;
assign c065 =  x364;
assign c067 = ~x16 & ~x65 & ~x240 & ~x273 & ~x716;
assign c069 =  x781;
assign c071 =  x112;
assign c073 =  x299 &  x384 & ~x32 & ~x48 & ~x143 & ~x200 & ~x282 & ~x341 & ~x388 & ~x703;
assign c075 =  x334 & ~x289;
assign c077 =  x563 &  x594;
assign c079 = ~x381;
assign c081 =  x525 & ~x46 & ~x48 & ~x77 & ~x136;
assign c083 =  x391;
assign c085 = ~x46 & ~x234 & ~x380 & ~x683;
assign c087 =  x363;
assign c089 =  x757;
assign c091 =  x344 &  x408 &  x638 & ~x108;
assign c093 =  x757;
assign c095 =  x780;
assign c097 =  x674;
assign c099 =  x335 &  x559;
assign c0101 =  x159 &  x203 &  x216 &  x245 &  x259 &  x266 &  x301 &  x325 &  x353 &  x356 &  x371 &  x381 &  x384 &  x412 &  x426 &  x432 &  x437 &  x510 &  x512 &  x539;
assign c0103 = ~x204 & ~x232 & ~x272 & ~x369;
assign c0105 = ~x215 & ~x352 & ~x743;
assign c0107 = ~x240 & ~x380 & ~x543;
assign c0109 = ~x39 & ~x204 & ~x429;
assign c0111 =  x189 &  x324 &  x328 &  x329 &  x356 &  x442 &  x443 &  x528;
assign c0113 =  x475;
assign c0115 =  x615;
assign c0117 =  x128 &  x264 &  x295 &  x432 &  x711 & ~x118 & ~x190 & ~x218 & ~x386 & ~x608 & ~x623;
assign c0119 =  x384 &  x525 & ~x742;
assign c0121 =  x156 & ~x229 & ~x568;
assign c0123 =  x28;
assign c0125 = ~x73 & ~x407 & ~x571;
assign c0127 =  x294 &  x385 &  x526 &  x593 &  x610;
assign c0129 =  x101 &  x153 &  x175 &  x179 &  x208 &  x209 &  x210 &  x291 &  x321 &  x379 &  x381 &  x402 &  x405 &  x436 &  x717 & ~x77 & ~x113 & ~x115 & ~x135 & ~x137 & ~x140 & ~x144 & ~x162 & ~x222 & ~x331 & ~x780;
assign c0131 =  x251;
assign c0133 =  x67 &  x68 &  x150 &  x184 &  x210 &  x211 &  x239 &  x291 &  x325 &  x381 &  x408 &  x463 &  x486 &  x492 &  x494 & ~x5 & ~x27 & ~x48 & ~x78 & ~x171 & ~x200 & ~x218 & ~x228 & ~x366 & ~x447 & ~x480 & ~x763;
assign c0135 =  x695;
assign c0137 =  x390 & ~x691;
assign c0139 = ~x100 & ~x202 & ~x246 & ~x568;
assign c0141 =  x649 &  x666 & ~x220;
assign c0143 =  x704;
assign c0145 =  x40 &  x74 &  x92 &  x179 &  x207 &  x267 &  x324 &  x436 &  x464 &  x579 & ~x8 & ~x33 & ~x478;
assign c0147 =  x279;
assign c0149 =  x412 & ~x10 & ~x17 & ~x32 & ~x77 & ~x105 & ~x224 & ~x248 & ~x366 & ~x367 & ~x390 & ~x422 & ~x452 & ~x759;
assign c0151 =  x22;
assign c0153 =  x783;
assign c0155 =  x643;
assign c0157 =  x505;
assign c0159 = ~x96 & ~x380 & ~x661;
assign c0161 =  x71 &  x344 &  x412 & ~x11 & ~x77 & ~x220 & ~x276 & ~x366 & ~x447 & ~x500;
assign c0163 =  x418;
assign c0165 =  x73 &  x104 &  x124 &  x128 &  x160 &  x188 &  x203 &  x211 &  x273 &  x466 & ~x77 & ~x362 & ~x734 & ~x761;
assign c0167 =  x273 &  x370 &  x510 &  x593 &  x610;
assign c0169 =  x616;
assign c0171 = ~x75 & ~x187 & ~x203 & ~x259 & ~x260 & ~x330;
assign c0173 =  x195;
assign c0175 =  x67 &  x188 &  x203 &  x204 &  x244 &  x245 &  x319 &  x348 &  x717 & ~x530 & ~x588 & ~x592 & ~x672 & ~x677 & ~x762;
assign c0179 = ~x64 & ~x69 & ~x259 & ~x290 & ~x485;
assign c0181 =  x85;
assign c0183 =  x629 &  x746 & ~x247 & ~x289;
assign c0185 = ~x207 & ~x208 & ~x380 & ~x515 & ~x683;
assign c0187 =  x14 &  x717 & ~x64 & ~x765;
assign c0189 = ~x73 & ~x430 & ~x745;
assign c0191 =  x446;
assign c0193 =  x756;
assign c0195 =  x167;
assign c0197 =  x14 & ~x23 & ~x134 & ~x138 & ~x144 & ~x163 & ~x173 & ~x189 & ~x228 & ~x247 & ~x248 & ~x251 & ~x420 & ~x422 & ~x446 & ~x451 & ~x561;
assign c0199 = ~x236 & ~x494 & ~x736;
assign c0201 =  x563;
assign c0203 =  x252;
assign c0205 =  x123 & ~x174 & ~x203 & ~x244 & ~x272 & ~x386;
assign c0207 = ~x319 & ~x348 & ~x437 & ~x707;
assign c0209 =  x141;
assign c0211 =  x448;
assign c0213 =  x464 &  x627 & ~x148 & ~x176 & ~x231 & ~x246 & ~x258;
assign c0215 =  x68 &  x120 &  x211 &  x661 &  x737 & ~x77 & ~x134 & ~x534 & ~x665;
assign c0217 =  x756;
assign c0219 = ~x64 & ~x256 & ~x434 & ~x545 & ~x601;
assign c0221 =  x14 & ~x20 & ~x77 & ~x135 & ~x224 & ~x310 & ~x367 & ~x474 & ~x506 & ~x765 & ~x782;
assign c0223 =  x168;
assign c0225 =  x668 & ~x314;
assign c0227 =  x84;
assign c0229 =  x279;
assign c0231 =  x615;
assign c0233 =  x296 &  x328 &  x528;
assign c0235 = ~x401 & ~x690 & ~x748;
assign c0237 =  x57;
assign c0239 =  x23;
assign c0241 =  x85;
assign c0243 =  x783;
assign c0245 =  x101 &  x123 &  x188 &  x210 &  x237 &  x409 &  x494 &  x607 &  x717 &  x718 & ~x34 & ~x55 & ~x228 & ~x278 & ~x308 & ~x313 & ~x340 & ~x366 & ~x387 & ~x475 & ~x555 & ~x560 & ~x610 & ~x695 & ~x697 & ~x754;
assign c0247 =  x167;
assign c0249 =  x10 &  x96 &  x176 &  x211 &  x322 &  x468 &  x493 & ~x86 & ~x389;
assign c0251 = ~x73 & ~x98 & ~x204;
assign c0253 =  x669;
assign c0257 =  x704;
assign c0259 = ~x46 & ~x47 & ~x437 & ~x689;
assign c0261 =  x68 &  x71 &  x96 &  x99 &  x127 &  x153 &  x210 &  x267 &  x291 &  x324 &  x346 &  x348 &  x380 &  x400 &  x456 &  x466 &  x493 &  x495 &  x577 & ~x48 & ~x51 & ~x62 & ~x89 & ~x307 & ~x388 & ~x393 & ~x424 & ~x589 & ~x703 & ~x753 & ~x781;
assign c0263 =  x510 &  x527;
assign c0265 =  x74 &  x96 &  x124 &  x125 &  x128 &  x182 &  x207 &  x237 &  x292 &  x403 &  x492 &  x494 &  x549 &  x717 &  x736 & ~x173 & ~x230 & ~x310 & ~x330 & ~x646 & ~x730;
assign c0267 =  x67 &  x102 &  x158 &  x325 &  x466 &  x495 & ~x117 & ~x191 & ~x526;
assign c0269 = ~x45 & ~x203 & ~x262;
assign c0271 =  x758;
assign c0273 =  x14 & ~x64 & ~x736;
assign c0275 =  x67 &  x154 &  x209 &  x319 &  x380 & ~x62 & ~x77 & ~x80 & ~x115 & ~x171 & ~x247 & ~x307 & ~x331 & ~x775 & ~x780;
assign c0277 =  x781;
assign c0279 =  x280;
assign c0281 =  x36 &  x37 &  x102 &  x103 &  x104 &  x128 &  x149 &  x158 &  x161 &  x175 &  x176 &  x182 &  x188 &  x210 &  x217 &  x244 &  x245 &  x272 &  x300 &  x301 &  x324 &  x328 &  x350 &  x400 &  x403 &  x404 &  x412 &  x428 &  x492 &  x495 &  x552 &  x571 &  x635 &  x661 & ~x0 & ~x85 & ~x87 & ~x114;
assign c0285 =  x156 &  x181 &  x211 &  x711 & ~x173 & ~x244 & ~x259 & ~x330 & ~x504 & ~x638;
assign c0287 =  x751;
assign c0289 =  x756;
assign c0291 = ~x46 & ~x231 & ~x545 & ~x568;
assign c0293 =  x167;
assign c0295 = ~x11 & ~x38 & ~x683;
assign c0297 =  x616;
assign c0299 =  x72 &  x524 & ~x47 & ~x77 & ~x557;
assign c0303 =  x93 &  x240 & ~x77 & ~x229;
assign c0305 =  x307;
assign c0307 =  x74 &  x125 &  x352 &  x717 & ~x692;
assign c0309 =  x203 &  x230 &  x273 &  x323 &  x325 &  x328 &  x538 &  x566 & ~x753 & ~x760 & ~x778;
assign c0311 = ~x72 & ~x186 & ~x736;
assign c0313 =  x14 & ~x77 & ~x134 & ~x161 & ~x249 & ~x256 & ~x259 & ~x272 & ~x301 & ~x302;
assign c0315 =  x66 &  x73 &  x74 &  x96 &  x103 &  x104 &  x131 &  x158 &  x176 &  x209 &  x238 &  x239 &  x319 &  x324 &  x325 &  x381 &  x403 &  x459 &  x548 &  x655 &  x660 &  x714 &  x774 & ~x83 & ~x110 & ~x165 & ~x254 & ~x334 & ~x341 & ~x424 & ~x675 & ~x723;
assign c0317 = ~x97 & ~x185 & ~x233;
assign c0319 =  x566;
assign c0321 =  x448;
assign c0323 = ~x47 & ~x262 & ~x368 & ~x691 & ~x736;
assign c0325 =  x418 & ~x234;
assign c0327 = ~x16 & ~x46 & ~x215 & ~x329;
assign c0329 =  x615;
assign c0331 =  x139;
assign c0333 =  x723;
assign c0335 =  x196;
assign c0337 =  x511 &  x525 &  x539 &  x555;
assign c0339 =  x161 &  x273 &  x291 &  x325 &  x356 &  x435 &  x552 &  x593;
assign c0341 = ~x46 & ~x47 & ~x64 & ~x231 & ~x257 & ~x286 & ~x287 & ~x312 & ~x315;
assign c0343 =  x67 &  x68 &  x153 &  x211 &  x348 &  x493 &  x633 & ~x19 & ~x22 & ~x33 & ~x35 & ~x105 & ~x168 & ~x285 & ~x528 & ~x561 & ~x613 & ~x701 & ~x775;
assign c0345 =  x37 &  x67 &  x74 &  x101 &  x104 &  x120 &  x122 &  x123 &  x124 &  x127 &  x128 &  x148 &  x150 &  x211 &  x235 &  x240 &  x293 &  x294 &  x324 &  x348 &  x377 &  x409 &  x464 &  x516 &  x520 &  x658 &  x718 &  x719 &  x736 & ~x20 & ~x80 & ~x338 & ~x448 & ~x449 & ~x589 & ~x705 & ~x761;
assign c0347 =  x37 &  x92 &  x101 &  x175 &  x187 &  x188 &  x209 &  x211 &  x231 &  x237 &  x273 &  x292 &  x325 &  x348 &  x350 &  x434 &  x457 &  x520 &  x548 &  x603 &  x709 &  x718 & ~x82 & ~x86 & ~x113 & ~x171 & ~x280 & ~x445 & ~x447 & ~x472 & ~x528 & ~x584 & ~x701 & ~x761;
assign c0349 =  x211 &  x655 & ~x230 & ~x244 & ~x316;
assign c0351 =  x4;
assign c0353 =  x532;
assign c0355 =  x728;
assign c0357 =  x683 & ~x48 & ~x77 & ~x105 & ~x204 & ~x229 & ~x231 & ~x232 & ~x286 & ~x330 & ~x342;
assign c0359 =  x96 &  x128 &  x438 &  x690 & ~x201 & ~x453 & ~x623;
assign c0361 =  x502;
assign c0363 =  x559;
assign c0365 =  x124 &  x182 &  x235 &  x291 &  x292 & ~x30 & ~x202 & ~x244 & ~x273 & ~x301 & ~x475 & ~x565;
assign c0367 =  x223 & ~x215;
assign c0369 =  x57;
assign c0371 =  x6 &  x588;
assign c0373 = ~x45 & ~x124 & ~x233 & ~x683;
assign c0375 =  x676;
assign c0377 =  x324 &  x648;
assign c0379 =  x620;
assign c0381 = ~x162 & ~x204 & ~x216 & ~x244 & ~x257 & ~x259 & ~x288 & ~x341 & ~x396;
assign c0383 =  x445;
assign c0385 =  x26;
assign c0389 =  x189 &  x230 &  x273 &  x324 &  x442 &  x566 &  x593;
assign c0391 =  x690 & ~x330 & ~x692 & ~x748;
assign c0393 =  x758;
assign c0395 =  x121 & ~x75 & ~x747;
assign c0399 =  x555 & ~x108 & ~x117;
assign c0401 =  x559;
assign c0403 =  x371 &  x416 &  x440 &  x526;
assign c0405 =  x527 &  x695;
assign c0407 =  x139;
assign c0409 =  x179 &  x272 &  x324 &  x328 &  x342 &  x426 &  x440 &  x442 & ~x777;
assign c0411 =  x67 &  x124 &  x127 &  x151 &  x156 &  x188 &  x296 &  x322 &  x325 &  x495 &  x627 &  x710 &  x739 & ~x77 & ~x90 & ~x694 & ~x695;
assign c0413 = ~x64 & ~x259 & ~x568 & ~x636 & ~x664;
assign c0415 =  x478;
assign c0417 = ~x47 & ~x231 & ~x269 & ~x301 & ~x342 & ~x720;
assign c0419 =  x124 &  x128 &  x324 &  x711 & ~x65;
assign c0421 =  x356 &  x511 &  x554 & ~x35 & ~x48 & ~x49;
assign c0423 =  x446;
assign c0425 =  x469 & ~x64 & ~x117 & ~x136 & ~x222;
assign c0427 =  x699;
assign c0429 =  x616;
assign c0431 = ~x286 & ~x434 & ~x571;
assign c0433 =  x492 & ~x75 & ~x204 & ~x217 & ~x243 & ~x273 & ~x301 & ~x386 & ~x613;
assign c0435 =  x14 &  x66 &  x324 &  x352;
assign c0437 = ~x214 & ~x233 & ~x541 & ~x661;
assign c0439 = ~x17 & ~x45 & ~x95 & ~x177 & ~x232;
assign c0441 =  x123 &  x466 & ~x173 & ~x664;
assign c0443 =  x123 &  x211 & ~x316;
assign c0445 = ~x176 & ~x204 & ~x215 & ~x259 & ~x288 & ~x314;
assign c0447 =  x363;
assign c0449 =  x82 &  x476;
assign c0451 =  x307;
assign c0453 =  x307;
assign c0455 =  x44 &  x72 &  x95 &  x126 &  x183 & ~x146 & ~x692;
assign c0457 = ~x65 & ~x116 & ~x215 & ~x246 & ~x288;
assign c0459 = ~x75 & ~x185 & ~x231 & ~x236 & ~x314;
assign c0461 =  x505;
assign c0463 =  x307;
assign c0465 =  x728;
assign c0467 =  x501;
assign c0469 =  x620;
assign c0471 =  x300 &  x400 & ~x229;
assign c0473 =  x447;
assign c0475 = ~x286 & ~x289 & ~x316;
assign c0477 =  x55;
assign c0479 = ~x17 & ~x232 & ~x245 & ~x288 & ~x664;
assign c0481 =  x723 & ~x32;
assign c0483 =  x671;
assign c0485 =  x476;
assign c0487 = ~x64 & ~x98 & ~x127 & ~x181 & ~x237 & ~x258 & ~x265;
assign c0489 =  x643;
assign c0491 =  x470 &  x510 & ~x745;
assign c0493 =  x704;
assign c0495 =  x189 &  x424 &  x554;
assign c0497 =  x421;
assign c0499 =  x648;
assign c10 =  x111;
assign c12 =  x25;
assign c14 = ~x69 & ~x86 & ~x97 & ~x187 & ~x355 & ~x389;
assign c16 =  x45 &  x157 &  x180 &  x712 & ~x90 & ~x107 & ~x169 & ~x308 & ~x386 & ~x536 & ~x566 & ~x594 & ~x646 & ~x648 & ~x674 & ~x695 & ~x697 & ~x722 & ~x742;
assign c18 =  x7;
assign c110 = ~x461 & ~x511 & ~x629;
assign c112 = ~x25 & ~x163 & ~x233 & ~x288 & ~x305 & ~x307 & ~x315 & ~x316 & ~x411 & ~x417 & ~x469 & ~x513 & ~x568 & ~x569 & ~x597 & ~x602 & ~x680;
assign c114 =  x747 & ~x434 & ~x629 & ~x685;
assign c116 =  x30;
assign c118 =  x721;
assign c120 =  x45 &  x495 &  x551 &  x687 & ~x692 & ~x776;
assign c122 = ~x32 & ~x85 & ~x257 & ~x334 & ~x378 & ~x434 & ~x537 & ~x611 & ~x645 & ~x742;
assign c124 =  x348 &  x488 &  x685 & ~x103 & ~x108 & ~x134 & ~x163 & ~x191 & ~x203 & ~x307 & ~x397 & ~x482 & ~x513 & ~x673;
assign c126 =  x579 &  x594 &  x624;
assign c128 =  x408 & ~x317 & ~x513 & ~x681;
assign c130 = ~x44 & ~x345 & ~x465 & ~x737;
assign c132 =  x644;
assign c134 =  x49 &  x482 &  x708 &  x736;
assign c136 =  x20 &  x203 &  x580;
assign c138 =  x759;
assign c140 = ~x205 & ~x439 & ~x513 & ~x708;
assign c142 =  x103 & ~x119 & ~x231 & ~x276 & ~x305 & ~x385 & ~x440 & ~x602 & ~x693;
assign c144 =  x45 &  x126 &  x268 &  x466 &  x521 & ~x546 & ~x617;
assign c146 =  x315 &  x679;
assign c148 =  x291 &  x460 & ~x0 & ~x6 & ~x31 & ~x54 & ~x60 & ~x92 & ~x136 & ~x144 & ~x175 & ~x176 & ~x188 & ~x199 & ~x202 & ~x216 & ~x231 & ~x255 & ~x258 & ~x276 & ~x288 & ~x301 & ~x303 & ~x307 & ~x317 & ~x336 & ~x373 & ~x416 & ~x426 & ~x428 & ~x439 & ~x441 & ~x448 & ~x477 & ~x485 & ~x497 & ~x506 & ~x513 & ~x529 & ~x530 & ~x538 & ~x566 & ~x567 & ~x585 & ~x620 & ~x639 & ~x648 & ~x669 & ~x677 & ~x706 & ~x707 & ~x761 & ~x763;
assign c150 =  x45 &  x315 &  x373 &  x607 &  x681 &  x765 & ~x730;
assign c152 =  x95 &  x345 &  x428 &  x456 &  x540 &  x765 & ~x80 & ~x284 & ~x534;
assign c154 =  x112;
assign c156 =  x317 &  x345 &  x401 & ~x12 & ~x328 & ~x568;
assign c158 =  x691 &  x734;
assign c160 =  x342;
assign c162 =  x436 & ~x215 & ~x345 & ~x513 & ~x738;
assign c164 =  x547 & ~x60 & ~x288 & ~x327 & ~x365 & ~x411 & ~x466 & ~x495 & ~x552 & ~x738;
assign c166 =  x512 &  x607 &  x717 & ~x601;
assign c168 =  x73 &  x181 &  x241 &  x270 &  x289 &  x317 &  x373 &  x376 &  x432 &  x551 & ~x30 & ~x77 & ~x139 & ~x286 & ~x677 & ~x699 & ~x732;
assign c170 =  x121 &  x262 &  x289 &  x710 & ~x188 & ~x216;
assign c172 =  x130 &  x207 &  x211 &  x520 & ~x14 & ~x315 & ~x316 & ~x502 & ~x552 & ~x569 & ~x597 & ~x635 & ~x652;
assign c174 = ~x0 & ~x43 & ~x140 & ~x316 & ~x427 & ~x485 & ~x513 & ~x527 & ~x654;
assign c176 =  x39 &  x68 &  x210 &  x319 &  x381 &  x436 &  x599 & ~x64 & ~x230 & ~x246 & ~x288 & ~x366 & ~x385 & ~x411 & ~x467 & ~x479 & ~x513 & ~x753;
assign c178 =  x9 &  x14;
assign c180 =  x241 &  x321 &  x376 &  x492 & ~x65 & ~x104 & ~x176 & ~x177 & ~x247 & ~x345 & ~x401 & ~x421 & ~x496 & ~x523 & ~x702 & ~x738 & ~x783;
assign c182 =  x435 & ~x371 & ~x373 & ~x449 & ~x495 & ~x542 & ~x610 & ~x652;
assign c184 =  x373 &  x399;
assign c186 = ~x232 & ~x382 & ~x513 & ~x709 & ~x737;
assign c188 =  x45 &  x124 &  x270 &  x321 &  x689 & ~x495;
assign c190 =  x157 &  x354 & ~x65 & ~x467 & ~x513 & ~x636 & ~x652 & ~x737;
assign c192 =  x392;
assign c194 =  x72 &  x240 &  x373 &  x400 &  x401 &  x428 &  x466 &  x484 &  x495 &  x540 &  x607 &  x624 &  x680 &  x736 & ~x55 & ~x286 & ~x453 & ~x502 & ~x585 & ~x615 & ~x778;
assign c196 =  x20 &  x175 &  x595;
assign c198 = ~x44 & ~x465 & ~x549;
assign c1100 =  x16 &  x328 &  x345 &  x495 &  x551;
assign c1102 =  x102 &  x289 &  x291 &  x323 &  x345 &  x352 &  x355 &  x401 &  x437 &  x439 &  x463 &  x491 &  x523 &  x551 &  x575 &  x598 & ~x35 & ~x90 & ~x144 & ~x161 & ~x170 & ~x224 & ~x252 & ~x286 & ~x306 & ~x309 & ~x396 & ~x511 & ~x584 & ~x611 & ~x669 & ~x672 & ~x705 & ~x782;
assign c1104 =  x10 &  x14 & ~x470 & ~x676;
assign c1106 =  x19 & ~x602;
assign c1108 =  x512 &  x652 & ~x685;
assign c1110 = ~x44 & ~x71 & ~x145 & ~x365 & ~x496;
assign c1112 = ~x70 & ~x150;
assign c1114 =  x14 &  x17 &  x19 &  x72 &  x262 &  x271 & ~x6 & ~x257 & ~x448 & ~x563 & ~x722 & ~x723 & ~x732;
assign c1116 =  x8;
assign c1118 = ~x352 & ~x380 & ~x741;
assign c1120 =  x226;
assign c1122 =  x293 &  x459 & ~x176 & ~x466;
assign c1124 =  x765 & ~x655;
assign c1126 =  x118 &  x607 &  x666;
assign c1128 =  x13 &  x16 &  x355 &  x541 & ~x229 & ~x453 & ~x482;
assign c1130 =  x270 & ~x575;
assign c1132 =  x644 &  x669;
assign c1134 = ~x263 & ~x439;
assign c1136 =  x44 &  x45 &  x151 &  x372 &  x373 &  x376 &  x400 &  x430 &  x551 &  x579 &  x659 &  x765 &  x766 & ~x1 & ~x5 & ~x472 & ~x500;
assign c1138 =  x45 &  x775 & ~x742;
assign c1140 =  x72 &  x156 &  x233 &  x326 &  x580 &  x607 &  x680 &  x765;
assign c1142 =  x19 & ~x247;
assign c1144 =  x408 & ~x317 & ~x335 & ~x382 & ~x401 & ~x410 & ~x485 & ~x513 & ~x595 & ~x623 & ~x738;
assign c1146 =  x644;
assign c1148 =  x43 &  x47 &  x74 &  x97 &  x125 &  x130 &  x212 &  x266 &  x270 &  x355 &  x429 &  x521 &  x606 &  x634 &  x662 &  x681 & ~x5 & ~x28 & ~x30 & ~x51 & ~x110 & ~x136 & ~x248 & ~x275 & ~x363 & ~x364 & ~x421 & ~x501 & ~x536 & ~x587 & ~x643 & ~x725 & ~x754;
assign c1150 =  x83;
assign c1152 = ~x147 & ~x226 & ~x233 & ~x345 & ~x355 & ~x401 & ~x485 & ~x513 & ~x523 & ~x578 & ~x581 & ~x607 & ~x619 & ~x625 & ~x636 & ~x667;
assign c1154 =  x45 &  x131 &  x158 &  x210 &  x262 &  x270 &  x289 &  x298 &  x326 &  x354 &  x383 & ~x26 & ~x27 & ~x50 & ~x202 & ~x285 & ~x310 & ~x367 & ~x448 & ~x454 & ~x470 & ~x481 & ~x511 & ~x567 & ~x595 & ~x620 & ~x637 & ~x696 & ~x753;
assign c1156 =  x624 &  x708 & ~x629 & ~x713;
assign c1158 = ~x3 & ~x135 & ~x221 & ~x378 & ~x399 & ~x434 & ~x483 & ~x553 & ~x567 & ~x673;
assign c1160 =  x30;
assign c1162 =  x54;
assign c1164 =  x45 &  x773 & ~x77 & ~x399 & ~x426 & ~x664 & ~x692 & ~x776;
assign c1166 =  x153 &  x402 &  x599 & ~x336 & ~x461 & ~x586;
assign c1168 =  x289 &  x290 &  x492 & ~x62 & ~x115 & ~x147 & ~x313 & ~x356 & ~x528 & ~x652;
assign c1170 =  x131 &  x176 &  x428 &  x765;
assign c1172 =  x312;
assign c1174 =  x20 &  x342;
assign c1176 =  x226 &  x283;
assign c1178 =  x20 &  x343;
assign c1180 =  x105 & ~x685;
assign c1182 =  x10 &  x15 &  x155 &  x205 &  x463 & ~x118 & ~x197 & ~x275 & ~x338 & ~x749;
assign c1184 =  x345 & ~x72 & ~x221 & ~x574 & ~x741;
assign c1186 =  x212 &  x233 &  x289 &  x488 & ~x2 & ~x313 & ~x315 & ~x330 & ~x336 & ~x343 & ~x412 & ~x423 & ~x510 & ~x617 & ~x663 & ~x675 & ~x702 & ~x735;
assign c1188 =  x45 &  x67 & ~x57 & ~x82 & ~x258 & ~x306 & ~x392 & ~x477 & ~x490 & ~x503 & ~x756 & ~x782;
assign c1190 =  x615;
assign c1192 =  x45 &  x400 &  x410 &  x512 &  x540 &  x551 &  x607 &  x624 &  x652 &  x736 & ~x118;
assign c1194 =  x16 &  x17 &  x261 & ~x188 & ~x247;
assign c1196 = ~x73 & ~x439 & ~x523 & ~x652;
assign c1198 = ~x130 & ~x158 & ~x159 & ~x382 & ~x513;
assign c1200 =  x45 &  x93 &  x100 &  x435 &  x439 &  x523 &  x548 &  x551 &  x743 &  x773 & ~x35 & ~x90 & ~x309 & ~x588;
assign c1202 =  x317 & ~x81 & ~x107 & ~x273 & ~x299 & ~x304 & ~x423 & ~x652;
assign c1204 =  x2;
assign c1206 =  x407 & ~x382 & ~x401 & ~x523 & ~x578 & ~x689;
assign c1208 =  x35 &  x621 & ~x573;
assign c1210 =  x297 &  x346 &  x378 &  x437 &  x684 & ~x15 & ~x301 & ~x513 & ~x737;
assign c1212 =  x373 & ~x0 & ~x518 & ~x742;
assign c1214 = ~x40 & ~x263 & ~x353 & ~x466;
assign c1216 =  x68 &  x94 &  x773 & ~x51 & ~x54 & ~x171 & ~x216 & ~x244 & ~x363 & ~x367 & ~x368 & ~x387 & ~x393 & ~x400 & ~x415 & ~x496 & ~x596 & ~x652 & ~x749;
assign c1218 =  x289 & ~x106 & ~x467 & ~x495 & ~x503 & ~x523 & ~x736;
assign c1220 =  x105 &  x175 &  x274 &  x454 &  x511 &  x595 &  x736;
assign c1222 =  x44 &  x235 &  x345 &  x401 &  x458 &  x712 & ~x88 & ~x413 & ~x427 & ~x428 & ~x455 & ~x523 & ~x596 & ~x622 & ~x652 & ~x693 & ~x694 & ~x708 & ~x727 & ~x760;
assign c1224 = ~x159 & ~x467 & ~x513 & ~x541 & ~x550 & ~x710;
assign c1226 =  x289 & ~x0 & ~x142 & ~x365 & ~x602;
assign c1228 =  x105 &  x734;
assign c1230 =  x624 & ~x546 & ~x742;
assign c1232 =  x10 &  x11 &  x14 &  x205 &  x289 &  x485 &  x548 &  x576 &  x658 & ~x419;
assign c1234 =  x671;
assign c1236 =  x10 &  x11 &  x13 & ~x133 & ~x198 & ~x412;
assign c1238 = ~x12 & ~x434 & ~x602;
assign c1240 = ~x629;
assign c1242 =  x20 &  x286 &  x343;
assign c1244 = ~x42 & ~x43 & ~x70 & ~x158 & ~x358 & ~x646;
assign c1246 =  x208 &  x321 &  x322 &  x375 & ~x191 & ~x382 & ~x505 & ~x662;
assign c1248 =  x105 &  x624 &  x734;
assign c1250 =  x532;
assign c1252 =  x28;
assign c1254 =  x39 &  x45 &  x122 &  x319 &  x324 &  x325 &  x488 &  x492 &  x516 &  x687 & ~x62 & ~x84 & ~x216 & ~x395 & ~x512 & ~x556 & ~x647 & ~x652 & ~x722;
assign c1256 =  x45 & ~x135 & ~x434 & ~x602;
assign c1258 =  x72 &  x93 &  x263 &  x288 &  x316 &  x353 &  x400 &  x428 &  x439 &  x512 &  x540 &  x652 &  x716 &  x736 & ~x60 & ~x253;
assign c1260 =  x126 &  x465 & ~x136 & ~x400 & ~x485;
assign c1262 =  x560;
assign c1264 =  x429 & ~x553 & ~x748;
assign c1266 =  x68 &  x399 &  x551 &  x681 &  x688 & ~x252;
assign c1268 =  x20 &  x356 &  x580;
assign c1270 =  x550 & ~x575;
assign c1272 =  x20 &  x147;
assign c1274 =  x76 &  x764 & ~x655;
assign c1278 = ~x139 & ~x224 & ~x246 & ~x275 & ~x288 & ~x303 & ~x333 & ~x366 & ~x389 & ~x412 & ~x425 & ~x496 & ~x558 & ~x574 & ~x595 & ~x602 & ~x619 & ~x622 & ~x636 & ~x669;
assign c1280 =  x645;
assign c1282 = ~x220 & ~x284 & ~x382 & ~x401 & ~x438 & ~x450 & ~x485 & ~x494 & ~x513 & ~x559 & ~x585 & ~x676 & ~x708;
assign c1284 =  x764;
assign c1286 =  x608 &  x652 & ~x630;
assign c1288 =  x10 & ~x349;
assign c1290 =  x294 & ~x64 & ~x466 & ~x606 & ~x633 & ~x680;
assign c1292 =  x588;
assign c1294 =  x463 & ~x53 & ~x103 & ~x187 & ~x192 & ~x201 & ~x215 & ~x217 & ~x260 & ~x271 & ~x298 & ~x305 & ~x382 & ~x466 & ~x485 & ~x501 & ~x523 & ~x537 & ~x591 & ~x607 & ~x614 & ~x730 & ~x753;
assign c1296 =  x125 & ~x36 & ~x356 & ~x602;
assign c1298 =  x756;
assign c1300 =  x45 &  x345 &  x654 & ~x686;
assign c1302 =  x289 &  x317 &  x345 & ~x87 & ~x161 & ~x300 & ~x427 & ~x495 & ~x509 & ~x607;
assign c1304 =  x45 &  x95 &  x100 &  x298 &  x463 &  x570 & ~x36 & ~x143 & ~x161 & ~x229 & ~x427 & ~x441 & ~x525 & ~x553 & ~x623 & ~x624 & ~x754 & ~x763;
assign c1306 =  x36 & ~x490 & ~x742;
assign c1308 =  x374 & ~x232 & ~x287 & ~x485 & ~x513;
assign c1310 = ~x23 & ~x188 & ~x228 & ~x602 & ~x636 & ~x676 & ~x721 & ~x736;
assign c1312 =  x10 &  x13 &  x317 & ~x192;
assign c1314 =  x235 &  x289 &  x292 &  x345 &  x407 &  x541 &  x542 &  x773 & ~x86 & ~x200 & ~x201 & ~x244 & ~x398 & ~x412 & ~x539;
assign c1316 =  x14 &  x20 &  x231;
assign c1318 =  x39 &  x68 &  x72 &  x349 &  x520 & ~x144 & ~x146 & ~x175 & ~x188 & ~x316 & ~x400 & ~x444 & ~x496 & ~x512 & ~x552 & ~x635 & ~x677 & ~x700 & ~x706;
assign c1320 =  x49 &  x162;
assign c1322 =  x588;
assign c1324 =  x421;
assign c1326 =  x68 &  x100 &  x289 &  x344 &  x659 & ~x33 & ~x495;
assign c1328 =  x344 &  x345 &  x484 &  x765 & ~x169 & ~x478 & ~x769;
assign c1330 =  x736 & ~x712;
assign c1332 =  x456 &  x484 &  x634 &  x653 &  x765 & ~x62 & ~x594 & ~x638;
assign c1334 =  x2;
assign c1336 =  x14 &  x16 &  x157 &  x242 &  x270 &  x458 &  x488 & ~x52 & ~x334 & ~x507;
assign c1338 =  x73 &  x317 &  x318 &  x322 &  x347 &  x400 &  x579 &  x607 &  x635 &  x765 & ~x50 & ~x77 & ~x202 & ~x218 & ~x641 & ~x778;
assign c1340 =  x30;
assign c1342 =  x403 & ~x490 & ~x629;
assign c1344 =  x743 & ~x329 & ~x410 & ~x537 & ~x550 & ~x569 & ~x681;
assign c1346 =  x439 &  x551 &  x765 & ~x0 & ~x424 & ~x693;
assign c1348 =  x21 &  x343;
assign c1350 =  x207 & ~x316 & ~x382 & ~x439 & ~x450 & ~x483 & ~x485 & ~x511 & ~x610 & ~x652;
assign c1352 =  x160 &  x373 &  x568 & ~x193;
assign c1354 =  x11 &  x487 & ~x287 & ~x400 & ~x508;
assign c1356 =  x435 & ~x205 & ~x345 & ~x373 & ~x466 & ~x560 & ~x626 & ~x654;
assign c1358 =  x454 &  x764;
assign c1360 =  x218 &  x342 &  x369 &  x397;
assign c1362 =  x429 & ~x136 & ~x166 & ~x277 & ~x336 & ~x503 & ~x518 & ~x615 & ~x685 & ~x740 & ~x743 & ~x768 & ~x769;
assign c1364 = ~x71 & ~x99;
assign c1366 =  x10 &  x14 & ~x0;
assign c1368 =  x20 &  x342;
assign c1370 =  x616;
assign c1372 =  x54 & ~x546;
assign c1374 =  x41 &  x44 &  x45 &  x74 &  x154 &  x289 &  x326 & ~x412;
assign c1376 =  x476;
assign c1378 =  x42 &  x45 &  x100 &  x151 &  x157 &  x183 &  x319 &  x376 &  x404 &  x576 & ~x3 & ~x4 & ~x24 & ~x26 & ~x140 & ~x172 & ~x188 & ~x192 & ~x252 & ~x302 & ~x307 & ~x315 & ~x332 & ~x335 & ~x363 & ~x364 & ~x368 & ~x385 & ~x394 & ~x428 & ~x440 & ~x478 & ~x479 & ~x495 & ~x540 & ~x551 & ~x568 & ~x579 & ~x583 & ~x612 & ~x615 & ~x636 & ~x647 & ~x671 & ~x702 & ~x723 & ~x726 & ~x779;
assign c1380 =  x40 &  x70 &  x157 & ~x24 & ~x91 & ~x216 & ~x244 & ~x274 & ~x412 & ~x455 & ~x484 & ~x495 & ~x523 & ~x636 & ~x640 & ~x707;
assign c1382 =  x308;
assign c1384 =  x14 & ~x75 & ~x467;
assign c1386 =  x45 &  x93 &  x634 & ~x308 & ~x671 & ~x714;
assign c1388 =  x10 &  x11 &  x13 & ~x2 & ~x5 & ~x202 & ~x419 & ~x441 & ~x646;
assign c1390 =  x323 &  x435 & ~x35 & ~x131 & ~x132 & ~x601 & ~x713;
assign c1392 =  x235 & ~x167 & ~x391 & ~x503 & ~x517 & ~x585 & ~x602 & ~x742 & ~x783;
assign c1394 = ~x99 & ~x327 & ~x512 & ~x689;
assign c1396 = ~x44 & ~x214 & ~x355;
assign c1398 = ~x119 & ~x172 & ~x258 & ~x396 & ~x434 & ~x448 & ~x581 & ~x624 & ~x641 & ~x652 & ~x669 & ~x771 & ~x778;
assign c1400 =  x1;
assign c1402 =  x19 & ~x479;
assign c1404 =  x20 & ~x658 & ~x742;
assign c1406 =  x45 &  x327 &  x344 &  x411 &  x523 & ~x330 & ~x497 & ~x595 & ~x675;
assign c1408 =  x48;
assign c1410 = ~x378 & ~x420 & ~x434 & ~x496 & ~x546 & ~x602 & ~x636;
assign c1412 =  x671;
assign c1414 =  x20 &  x373;
assign c1416 =  x484 &  x680 & ~x43 & ~x725;
assign c1418 =  x40 &  x131 &  x270 &  x514 & ~x194 & ~x602;
assign c1420 =  x622 &  x748 & ~x629;
assign c1422 =  x11 &  x72 &  x157 & ~x111 & ~x160 & ~x400 & ~x452 & ~x511 & ~x704;
assign c1424 = ~x72 & ~x434 & ~x518 & ~x602 & ~x742;
assign c1426 =  x627 & ~x43 & ~x69 & ~x70 & ~x131 & ~x367;
assign c1428 =  x36 &  x624 & ~x629 & ~x713;
assign c1430 =  x48 &  x371 &  x512;
assign c1432 = ~x71 & ~x100 & ~x652;
assign c1434 =  x484 & ~x685;
assign c1436 =  x123 &  x127 &  x402 & ~x333 & ~x391 & ~x490;
assign c1438 =  x123 &  x153 &  x178 &  x293 &  x402 &  x577 &  x633 & ~x317 & ~x345 & ~x535;
assign c1440 =  x547 & ~x13 & ~x43 & ~x158 & ~x286 & ~x287 & ~x299 & ~x418 & ~x483 & ~x694 & ~x697 & ~x776;
assign c1442 =  x20 & ~x712;
assign c1444 =  x42 & ~x350 & ~x454 & ~x575 & ~x652 & ~x771;
assign c1446 = ~x214 & ~x268 & ~x316 & ~x480;
assign c1448 =  x121 &  x242 &  x289 &  x401 &  x411 &  x429 &  x439 &  x579 &  x635 & ~x553;
assign c1450 =  x261 &  x401 &  x435 & ~x220 & ~x573 & ~x629;
assign c1452 =  x644;
assign c1454 =  x19 &  x262 & ~x136 & ~x192 & ~x278 & ~x338;
assign c1456 =  x291 &  x488 & ~x56 & ~x65 & ~x85 & ~x141 & ~x221 & ~x248 & ~x438 & ~x448 & ~x466 & ~x467 & ~x470 & ~x474 & ~x553 & ~x606 & ~x668 & ~x754 & ~x761 & ~x778;
assign c1458 =  x631 & ~x401 & ~x549 & ~x746;
assign c1460 =  x45 &  x131 &  x210 &  x242 &  x400 &  x428 &  x429 &  x512 &  x540 &  x652 &  x680 & ~x305 & ~x557;
assign c1462 = ~x69 & ~x97 & ~x218 & ~x316 & ~x411 & ~x447 & ~x694 & ~x707;
assign c1464 =  x14 & ~x316 & ~x513 & ~x555;
assign c1466 =  x547 & ~x131 & ~x187 & ~x382 & ~x655;
assign c1468 =  x402 &  x409 &  x655 & ~x2 & ~x7 & ~x24 & ~x34 & ~x50 & ~x53 & ~x62 & ~x79 & ~x114 & ~x134 & ~x198 & ~x218 & ~x228 & ~x230 & ~x246 & ~x303 & ~x311 & ~x314 & ~x358 & ~x363 & ~x387 & ~x396 & ~x413 & ~x426 & ~x444 & ~x452 & ~x453 & ~x478 & ~x499 & ~x500 & ~x502 & ~x509 & ~x536 & ~x553 & ~x583 & ~x587 & ~x609 & ~x637 & ~x742 & ~x752 & ~x754 & ~x756 & ~x783;
assign c1470 =  x206 &  x236 &  x322 &  x381 &  x405 &  x632 & ~x35 & ~x164 & ~x173 & ~x259 & ~x280 & ~x287 & ~x355 & ~x400 & ~x452 & ~x495 & ~x523 & ~x554 & ~x607 & ~x624 & ~x625 & ~x703 & ~x732 & ~x736 & ~x751;
assign c1472 =  x345 & ~x147 & ~x259 & ~x286 & ~x467 & ~x469 & ~x495 & ~x496 & ~x643;
assign c1474 =  x84;
assign c1476 =  x147 & ~x518 & ~x629 & ~x685 & ~x714;
assign c1478 =  x21 &  x454 &  x580;
assign c1480 =  x381 & ~x205 & ~x466 & ~x568;
assign c1482 =  x660 & ~x314 & ~x513 & ~x569 & ~x652;
assign c1484 =  x34 & ~x629;
assign c1486 =  x13 &  x16 &  x213 & ~x21 & ~x65 & ~x252 & ~x618;
assign c1488 =  x242 &  x431 &  x465 &  x483 &  x484 &  x595 &  x624 &  x651 & ~x30 & ~x77 & ~x282 & ~x646 & ~x673 & ~x779;
assign c1490 =  x184 & ~x259 & ~x410 & ~x452 & ~x513 & ~x605;
assign c1492 =  x55;
assign c1494 =  x45 & ~x283 & ~x434 & ~x462 & ~x568 & ~x575;
assign c1496 =  x755;
assign c1498 =  x83;
assign c11 =  x770;
assign c13 = ~x403 & ~x406 & ~x407;
assign c15 = ~x74 & ~x295 & ~x407;
assign c17 = ~x74 & ~x96 & ~x126;
assign c19 =  x770;
assign c111 =  x745 &  x769 &  x770 &  x771;
assign c113 =  x215 &  x299 &  x352 &  x627 &  x740 & ~x37 & ~x332 & ~x395;
assign c115 =  x152 &  x658 &  x683 &  x744 & ~x3 & ~x21 & ~x91 & ~x108 & ~x169 & ~x191 & ~x194 & ~x252 & ~x285 & ~x343 & ~x391 & ~x425 & ~x456 & ~x509 & ~x636 & ~x646 & ~x665 & ~x669 & ~x677;
assign c117 =  x272 & ~x607 & ~x718;
assign c119 =  x598 &  x740 &  x770 & ~x10 & ~x368 & ~x396 & ~x420 & ~x616;
assign c121 =  x296 &  x549 &  x745 &  x769 &  x770;
assign c123 =  x737 &  x770;
assign c125 =  x186 &  x269 &  x320 &  x405 &  x520 &  x597 &  x653 &  x681 &  x737 & ~x28 & ~x111 & ~x357 & ~x387 & ~x721 & ~x765;
assign c127 = ~x435 & ~x437 & ~x543 & ~x663;
assign c129 =  x351 &  x376 &  x487 &  x488 &  x494 &  x514 &  x516 &  x544 &  x548 &  x573 &  x600 & ~x31 & ~x33 & ~x79 & ~x113 & ~x142 & ~x166 & ~x193 & ~x196 & ~x306 & ~x311 & ~x338 & ~x340 & ~x392 & ~x420 & ~x422 & ~x701 & ~x754 & ~x770 & ~x772;
assign c131 =  x720 & ~x161 & ~x733;
assign c133 =  x427 &  x574 & ~x6 & ~x10 & ~x51 & ~x63 & ~x64 & ~x76 & ~x135 & ~x144 & ~x225 & ~x284 & ~x335;
assign c135 =  x78;
assign c137 = ~x3 & ~x74 & ~x94 & ~x124 & ~x125;
assign c139 =  x64 &  x65 &  x574 & ~x454;
assign c141 =  x189 &  x515 &  x656 & ~x27 & ~x167 & ~x336 & ~x337;
assign c143 =  x180 &  x264 &  x543 &  x709 & ~x14 & ~x678;
assign c145 = ~x86 & ~x113 & ~x194 & ~x375 & ~x403 & ~x431 & ~x487 & ~x532 & ~x544 & ~x587 & ~x607 & ~x615;
assign c147 =  x658 & ~x66 & ~x74 & ~x78 & ~x94 & ~x112 & ~x113;
assign c149 = ~x181 & ~x182 & ~x754;
assign c151 =  x92 &  x629 &  x630;
assign c153 = ~x600 & ~x604 & ~x635 & ~x708;
assign c155 =  x154 &  x655 & ~x262 & ~x290 & ~x298 & ~x317 & ~x734;
assign c157 =  x720 & ~x14 & ~x693;
assign c159 =  x359;
assign c161 =  x441 & ~x396 & ~x748 & ~x772;
assign c163 =  x473;
assign c165 = ~x74 & ~x105 & ~x133 & ~x153 & ~x154;
assign c167 =  x714 &  x742 & ~x25 & ~x175 & ~x213 & ~x279 & ~x336;
assign c169 =  x265 & ~x20 & ~x62;
assign c171 =  x163;
assign c173 =  x658 &  x746 &  x769 & ~x537;
assign c175 =  x390;
assign c177 =  x94 &  x155 &  x522 &  x571 &  x602 &  x627 &  x658 & ~x62 & ~x82 & ~x140 & ~x197 & ~x249 & ~x281 & ~x310 & ~x311 & ~x766;
assign c179 =  x546 & ~x85 & ~x213 & ~x467 & ~x551 & ~x566 & ~x679;
assign c181 =  x43 &  x351 &  x602 &  x740 &  x743 &  x769;
assign c183 =  x155 &  x490 &  x519 &  x571 &  x575 &  x627 &  x742 & ~x3 & ~x10 & ~x34 & ~x35 & ~x141 & ~x165 & ~x249 & ~x341 & ~x360 & ~x361 & ~x425 & ~x449 & ~x504 & ~x508 & ~x529 & ~x537 & ~x592 & ~x617 & ~x733;
assign c185 =  x212 &  x548 &  x658 &  x689 & ~x83 & ~x167 & ~x509 & ~x703 & ~x772;
assign c187 =  x176 &  x539 & ~x190 & ~x563;
assign c189 =  x64 &  x92 &  x742;
assign c191 = ~x209 & ~x210 & ~x322;
assign c193 = ~x103 & ~x124 & ~x125 & ~x126 & ~x195 & ~x773;
assign c195 =  x92 &  x155 & ~x18 & ~x414 & ~x642 & ~x700 & ~x722;
assign c197 = ~x125 & ~x149 & ~x185 & ~x773;
assign c199 = ~x379 & ~x403 & ~x408 & ~x751;
assign c1101 =  x520 &  x543 &  x658 &  x685 & ~x39 & ~x51 & ~x139 & ~x498 & ~x561 & ~x614 & ~x775;
assign c1103 =  x41 &  x180 &  x602 &  x658 &  x683 &  x715 &  x742 &  x744 & ~x27 & ~x29 & ~x270 & ~x301 & ~x414 & ~x456 & ~x644;
assign c1105 = ~x10 & ~x180 & ~x209 & ~x773;
assign c1107 =  x244 &  x658 &  x745 & ~x614 & ~x782;
assign c1109 = ~x108 & ~x238 & ~x265;
assign c1111 =  x178 &  x203 &  x259 &  x273 &  x330;
assign c1113 =  x686 & ~x297;
assign c1115 =  x273 &  x385 &  x413 &  x544;
assign c1117 =  x92 &  x575 &  x745 & ~x732;
assign c1119 =  x64 &  x76;
assign c1121 =  x761;
assign c1123 =  x331;
assign c1125 =  x658 &  x711 &  x744 &  x769 & ~x17 & ~x30 & ~x413 & ~x692 & ~x703;
assign c1127 = ~x209 & ~x224 & ~x656;
assign c1129 =  x78;
assign c1131 =  x549 &  x714 & ~x22 & ~x66 & ~x74 & ~x364 & ~x760;
assign c1133 =  x639;
assign c1135 =  x64 & ~x464;
assign c1137 =  x443;
assign c1139 =  x658 &  x740 &  x745 &  x770;
assign c1141 =  x732;
assign c1143 =  x441 & ~x36 & ~x52 & ~x89;
assign c1145 =  x548 &  x577 &  x625 &  x746 & ~x14 & ~x230;
assign c1147 =  x120 &  x718 & ~x79 & ~x339 & ~x564 & ~x750;
assign c1149 = ~x279 & ~x294 & ~x295 & ~x661;
assign c1151 =  x325 & ~x154;
assign c1153 =  x92 &  x742 &  x745;
assign c1155 = ~x140 & ~x291 & ~x294 & ~x661 & ~x667;
assign c1157 = ~x88 & ~x111 & ~x139 & ~x420 & ~x435 & ~x437 & ~x504 & ~x509 & ~x530 & ~x587 & ~x644 & ~x647 & ~x725 & ~x758 & ~x783;
assign c1159 =  x66 &  x489 & ~x716;
assign c1161 =  x69 &  x97 & ~x51 & ~x109 & ~x112 & ~x250 & ~x257 & ~x269 & ~x278 & ~x284 & ~x297 & ~x308 & ~x474 & ~x532 & ~x579 & ~x696 & ~x700 & ~x702 & ~x725;
assign c1163 =  x542 &  x548 &  x599 &  x658 &  x659 &  x739 & ~x62 & ~x82 & ~x104 & ~x116 & ~x121 & ~x133 & ~x142 & ~x192 & ~x203 & ~x224 & ~x225 & ~x228 & ~x247 & ~x343 & ~x364 & ~x369 & ~x388 & ~x449 & ~x535 & ~x556 & ~x583 & ~x615 & ~x644 & ~x648 & ~x674 & ~x724 & ~x725 & ~x750;
assign c1165 =  x98 &  x630 &  x692;
assign c1167 =  x97 &  x215 &  x630 & ~x45;
assign c1169 = ~x209 & ~x239;
assign c1171 =  x690 & ~x14 & ~x455 & ~x772;
assign c1173 =  x155 &  x157 &  x236 &  x742 & ~x3 & ~x326;
assign c1175 = ~x556 & ~x656 & ~x713 & ~x716;
assign c1177 =  x12 &  x378 &  x399 & ~x772;
assign c1179 = ~x154;
assign c1181 =  x740 &  x769 &  x770 & ~x14 & ~x779;
assign c1183 = ~x14 & ~x56 & ~x291;
assign c1185 =  x548 &  x654 &  x658 &  x716 &  x742 & ~x13 & ~x14 & ~x51 & ~x108 & ~x369 & ~x775;
assign c1187 =  x655 &  x770 & ~x14;
assign c1189 =  x66 &  x92 &  x713 &  x745 & ~x359 & ~x725;
assign c1191 = ~x103 & ~x184 & ~x185 & ~x262;
assign c1193 = ~x124 & ~x660;
assign c1195 = ~x10 & ~x37 & ~x108 & ~x152 & ~x310 & ~x755 & ~x780;
assign c1197 =  x120 &  x244 &  x517 & ~x223 & ~x612;
assign c1199 =  x493 &  x548 &  x571 &  x625 &  x653 &  x742 &  x746 & ~x7 & ~x9 & ~x109 & ~x221 & ~x359 & ~x414 & ~x423 & ~x593 & ~x699 & ~x725 & ~x733 & ~x751 & ~x782;
assign c1201 =  x207 &  x720 &  x742 & ~x447;
assign c1203 = ~x262 & ~x269 & ~x290;
assign c1205 =  x70 &  x238 &  x317 &  x402 &  x462 &  x517 &  x571 &  x625 & ~x60 & ~x109 & ~x333 & ~x340 & ~x419 & ~x526 & ~x644;
assign c1207 = ~x432 & ~x632 & ~x644;
assign c1209 = ~x403 & ~x406 & ~x408;
assign c1211 =  x384 & ~x20 & ~x46 & ~x757 & ~x775;
assign c1213 = ~x78 & ~x125 & ~x622 & ~x716;
assign c1215 = ~x14 & ~x86 & ~x121 & ~x460 & ~x477 & ~x564;
assign c1217 =  x155 &  x744 & ~x47 & ~x62 & ~x92 & ~x446 & ~x583 & ~x702 & ~x772;
assign c1219 =  x189 &  x323 &  x631 & ~x56 & ~x110 & ~x139 & ~x338;
assign c1221 =  x404 &  x636 &  x658 & ~x771 & ~x772;
assign c1223 =  x64;
assign c1225 =  x581 & ~x18 & ~x21 & ~x422 & ~x450 & ~x752 & ~x779;
assign c1227 = ~x211 & ~x435;
assign c1229 =  x97 &  x351 &  x438 &  x548 &  x769 &  x770 &  x771 & ~x197 & ~x250 & ~x451 & ~x530 & ~x588 & ~x783;
assign c1231 =  x742 & ~x6 & ~x346 & ~x526 & ~x533 & ~x613 & ~x751;
assign c1233 =  x352 & ~x194 & ~x707 & ~x717 & ~x738 & ~x764 & ~x781;
assign c1235 =  x549 &  x770;
assign c1237 =  x133 &  x658 & ~x252 & ~x504 & ~x671 & ~x782;
assign c1239 =  x745 &  x746 &  x769 &  x770;
assign c1241 = ~x576 & ~x627 & ~x777;
assign c1243 =  x64 &  x75 & ~x395 & ~x615;
assign c1245 = ~x526 & ~x576 & ~x600 & ~x638 & ~x663;
assign c1247 =  x64 &  x179 &  x210 &  x494 & ~x108 & ~x368 & ~x416 & ~x564;
assign c1249 =  x210 &  x629 &  x654 &  x710 &  x742 & ~x300 & ~x373 & ~x423 & ~x732;
assign c1251 = ~x75 & ~x164 & ~x224 & ~x435 & ~x775;
assign c1253 =  x415;
assign c1255 =  x70 &  x230 & ~x111 & ~x170 & ~x332 & ~x364 & ~x474 & ~x755;
assign c1257 = ~x32 & ~x82 & ~x632 & ~x644 & ~x653 & ~x660 & ~x696 & ~x752 & ~x773;
assign c1259 =  x742 & ~x232;
assign c1261 =  x745 & ~x10 & ~x56 & ~x262 & ~x364 & ~x447 & ~x473;
assign c1263 =  x676;
assign c1265 =  x658 &  x667;
assign c1267 =  x471 &  x499;
assign c1269 = ~x66 & ~x94 & ~x184;
assign c1271 =  x150 &  x236 &  x266 &  x434 &  x738 &  x742 &  x745 & ~x21 & ~x82 & ~x416 & ~x650;
assign c1273 =  x119 &  x549 &  x658;
assign c1275 =  x347 &  x655 &  x687 &  x742 & ~x6 & ~x20 & ~x262 & ~x306 & ~x317 & ~x450 & ~x534 & ~x562 & ~x614 & ~x666;
assign c1277 =  x70 &  x296 &  x406 &  x488 &  x602 &  x658 &  x740 &  x769 &  x770 &  x771 & ~x416 & ~x473;
assign c1279 =  x96 &  x155 &  x295 &  x325 &  x408 &  x513 &  x514 &  x549 & ~x252 & ~x713 & ~x772 & ~x773;
assign c1281 =  x261 &  x547 &  x575 &  x609 & ~x781;
assign c1283 =  x69 & ~x436 & ~x460;
assign c1285 =  x92 &  x120 & ~x621;
assign c1287 =  x770 & ~x14;
assign c1289 = ~x138 & ~x450 & ~x460 & ~x576 & ~x641 & ~x747 & ~x775;
assign c1291 =  x303;
assign c1293 =  x69 &  x629 &  x658 &  x742 & ~x242;
assign c1295 =  x70 &  x128 &  x517 &  x543 &  x544 &  x742 & ~x552 & ~x560 & ~x612 & ~x775;
assign c1297 =  x769 &  x770 &  x771 & ~x32;
assign c1299 =  x517 &  x658 &  x740 & ~x197 & ~x772;
assign c1301 =  x230 &  x273 & ~x527 & ~x679;
assign c1303 =  x268 & ~x154 & ~x444 & ~x732;
assign c1305 =  x770 & ~x92 & ~x298 & ~x559 & ~x644;
assign c1307 =  x245 &  x273 & ~x224 & ~x477 & ~x772 & ~x776;
assign c1309 = ~x435 & ~x498 & ~x632;
assign c1311 = ~x544 & ~x608 & ~x632 & ~x661;
assign c1313 =  x63 &  x75;
assign c1315 =  x148 &  x413 &  x441 & ~x702;
assign c1317 =  x258 &  x272 & ~x1 & ~x31 & ~x198 & ~x476 & ~x587 & ~x616 & ~x699 & ~x774 & ~x775;
assign c1319 =  x120 & ~x168 & ~x197 & ~x224 & ~x250 & ~x610 & ~x708 & ~x758 & ~x776;
assign c1321 =  x264 &  x600 &  x770 & ~x92 & ~x194 & ~x250 & ~x281 & ~x283 & ~x311 & ~x360 & ~x386 & ~x525 & ~x554 & ~x556 & ~x587 & ~x731 & ~x775;
assign c1323 =  x769 &  x770 & ~x121;
assign c1325 =  x378 &  x546 &  x742 &  x746 & ~x10 & ~x137 & ~x335;
assign c1327 = ~x1 & ~x10 & ~x103 & ~x114 & ~x133 & ~x325 & ~x779;
assign c1329 =  x598 &  x769 &  x770;
assign c1331 =  x360;
assign c1333 = ~x14 & ~x375 & ~x403;
assign c1335 =  x266 &  x320 &  x376 &  x434 &  x491 &  x548 &  x599 & ~x51 & ~x81 & ~x113 & ~x262 & ~x473 & ~x584 & ~x594 & ~x703;
assign c1337 =  x63 & ~x594;
assign c1339 =  x630 & ~x297;
assign c1341 =  x153 &  x746 &  x769 &  x770 &  x771;
assign c1343 = ~x14 & ~x57 & ~x126 & ~x772;
assign c1345 =  x329 &  x330 &  x358 &  x488 & ~x26 & ~x30;
assign c1347 =  x499;
assign c1349 =  x43 &  x548 &  x658 & ~x108 & ~x526;
assign c1351 =  x658 &  x742 &  x745 & ~x364 & ~x386 & ~x504 & ~x773;
assign c1353 =  x179 &  x180 &  x465 & ~x14 & ~x32 & ~x420 & ~x509 & ~x717;
assign c1355 =  x267 &  x548 &  x602 & ~x10 & ~x92 & ~x168 & ~x202 & ~x229 & ~x230 & ~x250 & ~x306 & ~x389 & ~x453 & ~x559 & ~x613 & ~x620 & ~x700 & ~x724 & ~x772;
assign c1357 = ~x14 & ~x52 & ~x60 & ~x137 & ~x197 & ~x211 & ~x250 & ~x252 & ~x351 & ~x463 & ~x721 & ~x725 & ~x731 & ~x751 & ~x775 & ~x783;
assign c1359 =  x658 &  x687 & ~x4 & ~x5 & ~x57 & ~x79 & ~x80 & ~x89 & ~x135 & ~x174 & ~x195 & ~x223 & ~x262 & ~x280 & ~x312 & ~x390 & ~x533 & ~x534 & ~x538 & ~x563 & ~x566 & ~x581 & ~x613 & ~x615 & ~x617 & ~x666 & ~x672 & ~x754 & ~x758 & ~x761 & ~x780 & ~x781;
assign c1361 = ~x14 & ~x51 & ~x88 & ~x142 & ~x202 & ~x715 & ~x716 & ~x718 & ~x758 & ~x759;
assign c1363 =  x705 & ~x197 & ~x776;
assign c1365 =  x546 &  x769 &  x770 & ~x113 & ~x369;
assign c1367 =  x602 &  x658 &  x714 &  x739 &  x740 &  x742 & ~x25 & ~x80 & ~x89 & ~x201 & ~x228 & ~x302 & ~x325 & ~x416 & ~x470 & ~x509 & ~x705 & ~x725;
assign c1369 = ~x14 & ~x51 & ~x238;
assign c1371 = ~x14 & ~x168 & ~x280 & ~x295;
assign c1373 =  x125 &  x465 &  x600 &  x630 & ~x5 & ~x51 & ~x78 & ~x89 & ~x165 & ~x168 & ~x171 & ~x249 & ~x303 & ~x341 & ~x396 & ~x418 & ~x425 & ~x473 & ~x475 & ~x501 & ~x536 & ~x559 & ~x645 & ~x723 & ~x728 & ~x730 & ~x772 & ~x782;
assign c1375 =  x329 & ~x5 & ~x7 & ~x20 & ~x34 & ~x56 & ~x57 & ~x84 & ~x752;
assign c1377 =  x44 & ~x492;
assign c1379 =  x518 &  x548 &  x742 &  x746 & ~x671 & ~x727;
assign c1381 =  x249;
assign c1383 =  x387 & ~x748;
assign c1385 =  x219;
assign c1387 = ~x161 & ~x200 & ~x238 & ~x275 & ~x448 & ~x473 & ~x508 & ~x619 & ~x642 & ~x645 & ~x646 & ~x695 & ~x704 & ~x779;
assign c1389 =  x77 & ~x414;
assign c1391 =  x215 &  x348 &  x524 &  x539 & ~x23;
assign c1393 = ~x54 & ~x92 & ~x169 & ~x336 & ~x586 & ~x626 & ~x628 & ~x655 & ~x713 & ~x716 & ~x773;
assign c1395 =  x273 & ~x60 & ~x141 & ~x197 & ~x366 & ~x389 & ~x772;
assign c1397 =  x244 &  x413 &  x441 & ~x197;
assign c1399 =  x96 &  x123 &  x127 &  x153 &  x209 &  x295 &  x433 &  x548 &  x577 &  x598 &  x628 &  x658 & ~x81 & ~x84 & ~x168 & ~x196 & ~x247 & ~x252 & ~x336 & ~x340 & ~x391 & ~x395 & ~x397 & ~x445 & ~x447 & ~x479 & ~x501 & ~x528 & ~x530 & ~x585 & ~x617 & ~x696 & ~x725 & ~x759 & ~x770 & ~x772;
assign c1401 = ~x223 & ~x224 & ~x237 & ~x308 & ~x754 & ~x755 & ~x777 & ~x782;
assign c1403 =  x720 &  x770;
assign c1405 =  x770 & ~x206;
assign c1407 =  x188 &  x204 &  x658;
assign c1409 = ~x210 & ~x239;
assign c1411 =  x70 &  x235 &  x268 &  x405 &  x516 &  x548 &  x602 &  x630 &  x658 & ~x17 & ~x245 & ~x420 & ~x475 & ~x509 & ~x722 & ~x749 & ~x768;
assign c1413 =  x273 &  x351 & ~x86 & ~x249 & ~x250 & ~x367 & ~x421 & ~x559 & ~x756;
assign c1415 =  x43 & ~x408;
assign c1417 =  x125 &  x566;
assign c1419 = ~x493 & ~x548 & ~x570;
assign c1421 = ~x11 & ~x75 & ~x230 & ~x764 & ~x772 & ~x775;
assign c1423 =  x69 &  x270 &  x510 & ~x48 & ~x169;
assign c1425 =  x164;
assign c1427 =  x155 &  x187 &  x625 &  x745 &  x746 & ~x751;
assign c1429 =  x510 &  x630 & ~x256;
assign c1431 =  x546 &  x571 &  x603 & ~x51 & ~x75 & ~x718 & ~x773;
assign c1433 = ~x5 & ~x6 & ~x7 & ~x8 & ~x54 & ~x81 & ~x107 & ~x113 & ~x166 & ~x169 & ~x195 & ~x196 & ~x224 & ~x226 & ~x249 & ~x252 & ~x334 & ~x362 & ~x472 & ~x475 & ~x478 & ~x702 & ~x715 & ~x716 & ~x717 & ~x776 & ~x783;
assign c1435 =  x163;
assign c1437 =  x603 &  x769 &  x770 &  x772 & ~x420 & ~x509 & ~x582;
assign c1439 =  x43 &  x492 &  x571 &  x601 &  x658 &  x745 & ~x10 & ~x11;
assign c1441 =  x68 &  x92 & ~x476 & ~x702;
assign c1443 =  x465 &  x491 &  x599 & ~x14 & ~x92 & ~x103 & ~x399 & ~x695 & ~x772;
assign c1445 = ~x1 & ~x59 & ~x74 & ~x124 & ~x125 & ~x126 & ~x716 & ~x718 & ~x738 & ~x773;
assign c1447 = ~x154 & ~x663 & ~x688;
assign c1449 =  x120 &  x176 &  x188 &  x546;
assign c1451 =  x244 &  x603 &  x737;
assign c1453 =  x742 &  x745 &  x769 &  x770;
assign c1455 = ~x298 & ~x348 & ~x408;
assign c1457 = ~x10 & ~x21 & ~x59 & ~x91 & ~x105 & ~x148 & ~x164 & ~x184 & ~x185 & ~x190 & ~x197 & ~x222 & ~x249 & ~x280 & ~x421 & ~x676 & ~x698 & ~x758 & ~x775;
assign c1459 =  x720;
assign c1461 = ~x267 & ~x351 & ~x521;
assign c1463 =  x200;
assign c1465 = ~x42 & ~x83 & ~x209 & ~x781;
assign c1467 =  x96 &  x97 &  x406 &  x408 &  x577 &  x602 &  x630 & ~x63 & ~x113 & ~x170 & ~x225 & ~x509 & ~x772;
assign c1469 = ~x0 & ~x251 & ~x509 & ~x556 & ~x561 & ~x592 & ~x632 & ~x638;
assign c1471 =  x43 &  x92 &  x517 &  x661;
assign c1473 =  x639;
assign c1475 =  x302 & ~x730;
assign c1477 =  x376 &  x683 &  x686 &  x687 & ~x45 & ~x368 & ~x450 & ~x764;
assign c1479 = ~x265 & ~x266 & ~x775;
assign c1481 = ~x14 & ~x94 & ~x128 & ~x208;
assign c1483 =  x64;
assign c1485 =  x517 &  x544 &  x684 &  x743 &  x745 &  x769 &  x770 &  x771 & ~x81 & ~x161 & ~x174;
assign c1487 = ~x14 & ~x24 & ~x83 & ~x112 & ~x169 & ~x170 & ~x238 & ~x253 & ~x365 & ~x476 & ~x588 & ~x642 & ~x759;
assign c1489 = ~x38 & ~x111 & ~x126 & ~x154 & ~x235 & ~x283 & ~x364;
assign c1491 =  x720 &  x742 & ~x113;
assign c1493 =  x629 &  x720 &  x742 &  x743 &  x745 &  x769 & ~x113 & ~x724;
assign c1495 =  x557;
assign c1497 =  x630 &  x658 &  x770 & ~x149;
assign c1499 = ~x619 & ~x634 & ~x663 & ~x683 & ~x735 & ~x754 & ~x772;
assign c20 =  x90 &  x175 &  x489 & ~x87 & ~x198 & ~x283 & ~x395 & ~x504 & ~x591;
assign c22 =  x68 &  x244 &  x273 &  x330 &  x433 &  x442 &  x464 &  x493 &  x525 &  x542 &  x547 &  x550 &  x582 &  x599 &  x622 &  x628 &  x632 &  x657 &  x660 &  x663 &  x678 &  x750 & ~x5 & ~x6 & ~x19 & ~x60 & ~x61 & ~x75 & ~x77 & ~x163 & ~x172 & ~x195 & ~x197 & ~x199 & ~x200 & ~x223 & ~x252 & ~x256 & ~x275 & ~x276 & ~x311 & ~x360 & ~x393 & ~x394 & ~x416 & ~x447 & ~x448 & ~x502 & ~x507 & ~x560 & ~x590 & ~x616 & ~x618 & ~x700 & ~x726 & ~x754;
assign c24 =  x512 &  x514 &  x610 &  x655 &  x709 &  x710 &  x711 &  x715 &  x778 & ~x19 & ~x56 & ~x88 & ~x111 & ~x140 & ~x227 & ~x254 & ~x278 & ~x365 & ~x474 & ~x477 & ~x478 & ~x504 & ~x590 & ~x703;
assign c26 = ~x31 & ~x32 & ~x50 & ~x115 & ~x166 & ~x277 & ~x310 & ~x364 & ~x384 & ~x440 & ~x506 & ~x671 & ~x740 & ~x741 & ~x742 & ~x745 & ~x771 & ~x773;
assign c28 =  x91 &  x204 &  x212 &  x319 &  x349 &  x481 &  x550 &  x604 & ~x27 & ~x282 & ~x304 & ~x770 & ~x774;
assign c210 =  x721 & ~x628 & ~x631 & ~x657;
assign c212 =  x331 &  x370 &  x387 & ~x278 & ~x665 & ~x672;
assign c214 =  x44 & ~x25 & ~x26 & ~x58 & ~x88 & ~x107 & ~x136 & ~x144 & ~x164 & ~x170 & ~x200 & ~x220 & ~x227 & ~x249 & ~x250 & ~x282 & ~x306 & ~x309 & ~x336 & ~x364 & ~x389 & ~x391 & ~x419 & ~x424 & ~x438 & ~x446 & ~x476 & ~x616 & ~x668 & ~x697 & ~x699 & ~x726 & ~x727 & ~x729 & ~x757 & ~x759;
assign c216 =  x192;
assign c218 =  x42 & ~x98 & ~x390 & ~x402;
assign c220 = ~x54 & ~x71 & ~x223 & ~x227 & ~x729 & ~x738 & ~x741 & ~x745 & ~x763 & ~x783;
assign c222 = ~x58 & ~x206 & ~x222 & ~x280 & ~x295 & ~x335 & ~x365 & ~x378 & ~x472 & ~x503 & ~x504 & ~x530 & ~x670 & ~x697;
assign c224 =  x750 & ~x249 & ~x275 & ~x682 & ~x683 & ~x686 & ~x689 & ~x714 & ~x717 & ~x719 & ~x745;
assign c226 =  x777 & ~x116 & ~x194 & ~x196 & ~x275 & ~x443 & ~x556 & ~x618 & ~x639 & ~x770 & ~x773;
assign c228 =  x247 &  x779;
assign c230 =  x125 &  x159 &  x160 &  x179 &  x206 &  x217 &  x231 &  x232 &  x244 &  x245 &  x298 &  x302 &  x345 &  x349 &  x354 &  x358 &  x370 &  x381 &  x402 &  x411 &  x434 &  x454 &  x458 &  x520 &  x538 &  x549 &  x570 &  x573 &  x594 &  x600 &  x602 &  x603 &  x604 &  x653 &  x722 & ~x33 & ~x110 & ~x113 & ~x138 & ~x167 & ~x193 & ~x225 & ~x228 & ~x252 & ~x254 & ~x282 & ~x308 & ~x336 & ~x337 & ~x339 & ~x362 & ~x390 & ~x473 & ~x476 & ~x501 & ~x502 & ~x535 & ~x560 & ~x587 & ~x642 & ~x670 & ~x697 & ~x700 & ~x725 & ~x727;
assign c232 = ~x330 & ~x382 & ~x388 & ~x410 & ~x423 & ~x424 & ~x531;
assign c234 =  x68 &  x175 &  x232 &  x599 &  x609 &  x627 &  x679 &  x681 &  x685 & ~x7 & ~x48 & ~x52 & ~x88 & ~x107 & ~x139 & ~x219 & ~x226 & ~x248 & ~x250 & ~x275 & ~x283 & ~x304 & ~x305 & ~x333 & ~x360 & ~x388 & ~x395 & ~x591 & ~x644 & ~x724 & ~x779;
assign c236 =  x398 & ~x1 & ~x4 & ~x24 & ~x25 & ~x26 & ~x27 & ~x29 & ~x30 & ~x52 & ~x55 & ~x56 & ~x58 & ~x85 & ~x86 & ~x109 & ~x110 & ~x112 & ~x138 & ~x142 & ~x143 & ~x165 & ~x168 & ~x169 & ~x194 & ~x222 & ~x254 & ~x281 & ~x305 & ~x307 & ~x308 & ~x334 & ~x362 & ~x363 & ~x392 & ~x418 & ~x420 & ~x446 & ~x448 & ~x473 & ~x476 & ~x501 & ~x503 & ~x588 & ~x616 & ~x642 & ~x644 & ~x671 & ~x699 & ~x700 & ~x701 & ~x726 & ~x729 & ~x738 & ~x741 & ~x742 & ~x744 & ~x754 & ~x761 & ~x762 & ~x766 & ~x767 & ~x771 & ~x775 & ~x782 & ~x783;
assign c238 =  x46 &  x162 &  x259 &  x303 &  x387 &  x434 &  x549 &  x633 &  x708 & ~x60 & ~x222;
assign c240 = ~x10 & ~x26 & ~x103 & ~x104 & ~x132 & ~x421 & ~x523;
assign c242 = ~x4 & ~x8 & ~x21 & ~x22 & ~x23 & ~x26 & ~x34 & ~x61 & ~x81 & ~x87 & ~x88 & ~x113 & ~x137 & ~x140 & ~x164 & ~x169 & ~x172 & ~x192 & ~x195 & ~x199 & ~x226 & ~x228 & ~x250 & ~x281 & ~x283 & ~x304 & ~x309 & ~x332 & ~x335 & ~x365 & ~x367 & ~x390 & ~x417 & ~x420 & ~x445 & ~x448 & ~x475 & ~x501 & ~x529 & ~x535 & ~x540 & ~x558 & ~x614 & ~x615 & ~x616 & ~x617 & ~x644 & ~x701 & ~x703 & ~x731 & ~x740 & ~x741 & ~x742 & ~x743 & ~x745 & ~x746 & ~x759 & ~x770 & ~x775;
assign c244 =  x104 &  x161 &  x434 & ~x15 & ~x78 & ~x221 & ~x283 & ~x422;
assign c246 =  x752 & ~x4 & ~x665;
assign c248 = ~x245 & ~x570;
assign c250 = ~x76 & ~x164 & ~x179 & ~x332 & ~x333 & ~x334 & ~x338 & ~x395 & ~x424 & ~x445 & ~x450 & ~x451 & ~x478 & ~x502 & ~x528 & ~x529 & ~x531 & ~x556 & ~x586 & ~x642 & ~x725 & ~x741 & ~x769 & ~x770 & ~x771 & ~x772;
assign c252 =  x511 &  x749 & ~x0 & ~x30 & ~x56 & ~x86 & ~x105 & ~x116 & ~x138 & ~x141 & ~x142 & ~x144 & ~x145 & ~x191 & ~x200 & ~x226 & ~x249 & ~x253 & ~x255 & ~x275 & ~x303 & ~x309 & ~x311 & ~x312 & ~x340 & ~x362 & ~x367 & ~x368 & ~x423 & ~x443 & ~x448 & ~x476 & ~x532 & ~x585 & ~x612 & ~x615 & ~x616 & ~x618 & ~x729 & ~x764 & ~x765 & ~x767 & ~x771 & ~x774;
assign c254 = ~x303 & ~x545 & ~x571;
assign c256 = ~x281 & ~x354 & ~x390 & ~x438 & ~x473 & ~x474 & ~x586 & ~x767 & ~x770 & ~x771 & ~x775;
assign c258 =  x41 & ~x21 & ~x73 & ~x79 & ~x98 & ~x227 & ~x282 & ~x445 & ~x502 & ~x503;
assign c260 =  x312 &  x396 &  x424 & ~x34;
assign c262 = ~x271 & ~x436 & ~x439 & ~x492;
assign c264 =  x173 &  x201 &  x257 &  x330 &  x375 &  x441 &  x544 &  x601 &  x733 & ~x34 & ~x49 & ~x115 & ~x530 & ~x557 & ~x672;
assign c266 =  x315 &  x518 & ~x27 & ~x79 & ~x85 & ~x227 & ~x249 & ~x255 & ~x360 & ~x474 & ~x682 & ~x683 & ~x686 & ~x689 & ~x690 & ~x698 & ~x714 & ~x719 & ~x745 & ~x769;
assign c268 =  x160 &  x190 &  x387 & ~x562;
assign c270 = ~x172 & ~x283 & ~x446 & ~x478 & ~x540 & ~x712 & ~x713 & ~x717 & ~x740 & ~x741 & ~x746;
assign c272 = ~x41 & ~x770;
assign c274 =  x102 &  x189 &  x414 &  x489 & ~x192 & ~x646 & ~x710 & ~x712 & ~x714 & ~x717 & ~x719 & ~x726;
assign c276 =  x62 &  x228;
assign c278 =  x317 &  x401 & ~x10 & ~x12 & ~x15 & ~x114 & ~x172 & ~x253 & ~x614 & ~x678;
assign c280 =  x772 &  x774;
assign c282 =  x256 &  x648;
assign c284 =  x273 &  x329 &  x351 &  x438 &  x514 &  x516 &  x554 & ~x7 & ~x23 & ~x83 & ~x163 & ~x171 & ~x192 & ~x227 & ~x332 & ~x420 & ~x477 & ~x500 & ~x645 & ~x719 & ~x730 & ~x780;
assign c286 =  x175 &  x301 &  x414 &  x576 &  x628 & ~x8 & ~x15 & ~x33 & ~x49 & ~x228 & ~x760;
assign c288 =  x778 & ~x228 & ~x275 & ~x303 & ~x748 & ~x755 & ~x757 & ~x782;
assign c290 =  x749 & ~x6 & ~x35 & ~x52 & ~x64 & ~x133 & ~x190 & ~x221 & ~x360 & ~x387 & ~x419 & ~x770 & ~x772;
assign c292 =  x411 & ~x20 & ~x34 & ~x109 & ~x172 & ~x364 & ~x391 & ~x416 & ~x424 & ~x450 & ~x501 & ~x586 & ~x680 & ~x700 & ~x731;
assign c294 = ~x377 & ~x379 & ~x406 & ~x434 & ~x436 & ~x490 & ~x491 & ~x546;
assign c296 =  x191 &  x247 &  x331 &  x359 & ~x164;
assign c298 = ~x28 & ~x56 & ~x58 & ~x59 & ~x83 & ~x107 & ~x112 & ~x113 & ~x137 & ~x138 & ~x141 & ~x168 & ~x194 & ~x220 & ~x221 & ~x225 & ~x226 & ~x227 & ~x254 & ~x280 & ~x304 & ~x305 & ~x310 & ~x334 & ~x337 & ~x360 & ~x363 & ~x364 & ~x389 & ~x392 & ~x444 & ~x445 & ~x446 & ~x447 & ~x449 & ~x473 & ~x501 & ~x506 & ~x531 & ~x552 & ~x585 & ~x613 & ~x615 & ~x636 & ~x645 & ~x697 & ~x701 & ~x728 & ~x738 & ~x740 & ~x741 & ~x744 & ~x745 & ~x746 & ~x755 & ~x770 & ~x773 & ~x775 & ~x776;
assign c2100 = ~x107 & ~x170 & ~x276 & ~x279 & ~x304 & ~x332 & ~x360 & ~x402 & ~x446 & ~x450 & ~x618;
assign c2102 =  x132 & ~x172 & ~x219 & ~x283 & ~x303 & ~x310 & ~x331 & ~x710 & ~x712 & ~x714 & ~x717 & ~x769 & ~x773;
assign c2104 =  x734 & ~x219 & ~x332 & ~x620 & ~x683 & ~x710;
assign c2106 = ~x68 & ~x72 & ~x169 & ~x193 & ~x199 & ~x226 & ~x276 & ~x333 & ~x336 & ~x390 & ~x533 & ~x558 & ~x559 & ~x740 & ~x746 & ~x767 & ~x773 & ~x775;
assign c2108 =  x454 &  x498 &  x717 &  x778 & ~x91 & ~x195 & ~x279 & ~x310 & ~x393 & ~x533 & ~x697;
assign c2110 =  x518 & ~x0 & ~x167 & ~x227 & ~x474 & ~x539 & ~x561 & ~x595 & ~x766 & ~x770;
assign c2112 = ~x153 & ~x154 & ~x277 & ~x367 & ~x439 & ~x495 & ~x769;
assign c2114 =  x371 &  x457 &  x492 &  x576 &  x750 & ~x23 & ~x27 & ~x28 & ~x49 & ~x62 & ~x136 & ~x137 & ~x163 & ~x200 & ~x227 & ~x249 & ~x304 & ~x333 & ~x388 & ~x395 & ~x417 & ~x473 & ~x535 & ~x696 & ~x699 & ~x729 & ~x738 & ~x741 & ~x742 & ~x747 & ~x756 & ~x757;
assign c2116 =  x132 &  x148 &  x322 &  x358 &  x407 &  x432 &  x520 &  x653 & ~x85 & ~x88 & ~x110 & ~x311 & ~x473 & ~x475 & ~x735 & ~x741;
assign c2118 =  x276 &  x528;
assign c2120 =  x70 &  x159 &  x160 &  x175 &  x288 &  x430 &  x431 &  x432 &  x486 &  x517 &  x654 &  x707 & ~x56 & ~x219 & ~x283 & ~x390 & ~x726 & ~x729;
assign c2122 =  x175 &  x190 &  x273 &  x298 &  x300 &  x430 &  x491 &  x706 & ~x59 & ~x78 & ~x83 & ~x195 & ~x221 & ~x255 & ~x360 & ~x388 & ~x420 & ~x504 & ~x532 & ~x619 & ~x755;
assign c2124 =  x45 &  x187 &  x385 &  x426 & ~x2 & ~x12 & ~x15 & ~x27 & ~x49 & ~x56 & ~x135 & ~x138 & ~x172 & ~x226 & ~x421 & ~x504;
assign c2126 = ~x98 & ~x103 & ~x439;
assign c2128 =  x767 &  x774 & ~x256 & ~x333;
assign c2130 = ~x75 & ~x132 & ~x410 & ~x521;
assign c2132 =  x534;
assign c2134 =  x204 &  x469 &  x542 &  x711 &  x714 &  x778 & ~x116 & ~x171 & ~x196 & ~x281 & ~x445 & ~x449 & ~x450 & ~x753 & ~x754 & ~x769 & ~x780;
assign c2136 = ~x73 & ~x75 & ~x128 & ~x274 & ~x302 & ~x415 & ~x449 & ~x473 & ~x762;
assign c2138 = ~x2 & ~x29 & ~x30 & ~x50 & ~x56 & ~x58 & ~x87 & ~x138 & ~x192 & ~x196 & ~x198 & ~x226 & ~x275 & ~x279 & ~x306 & ~x335 & ~x367 & ~x389 & ~x395 & ~x418 & ~x419 & ~x422 & ~x467 & ~x523 & ~x534 & ~x563 & ~x585 & ~x587 & ~x615 & ~x672 & ~x740 & ~x745 & ~x757 & ~x767;
assign c2140 =  x456 &  x511 &  x737 &  x778;
assign c2142 =  x556 &  x724 & ~x15;
assign c2144 =  x715 &  x724;
assign c2146 =  x76 &  x190 &  x425 &  x621 & ~x391 & ~x451 & ~x586 & ~x675 & ~x763 & ~x781;
assign c2148 =  x44 &  x68 &  x322 &  x432 &  x435 &  x521 &  x547 &  x549 &  x653 &  x738 & ~x1 & ~x2 & ~x11 & ~x256 & ~x283;
assign c2150 =  x105 &  x161 & ~x15;
assign c2152 =  x407 &  x408 &  x454 &  x522 &  x711 &  x750 & ~x82 & ~x91 & ~x105 & ~x226 & ~x228 & ~x283 & ~x530 & ~x558 & ~x757;
assign c2154 =  x502;
assign c2156 =  x451 &  x507;
assign c2158 = ~x97 & ~x401 & ~x571;
assign c2160 = ~x104 & ~x138 & ~x226 & ~x332 & ~x361 & ~x362 & ~x451 & ~x501 & ~x521 & ~x550;
assign c2162 = ~x75 & ~x104 & ~x302 & ~x439 & ~x495 & ~x669;
assign c2164 =  x43 &  x72 &  x245 &  x287 &  x385 &  x386 &  x410 &  x442 &  x461 &  x490 &  x518 &  x520 &  x545 &  x549 &  x573 &  x633 &  x653 &  x662 &  x683 &  x688 &  x778 & ~x5 & ~x31 & ~x33 & ~x85 & ~x86 & ~x87 & ~x142 & ~x164 & ~x166 & ~x195 & ~x222 & ~x283 & ~x419 & ~x475 & ~x477 & ~x587 & ~x590 & ~x642 & ~x726 & ~x731 & ~x754;
assign c2166 =  x46 &  x247 &  x331 & ~x8 & ~x170 & ~x730;
assign c2168 =  x433 &  x773 &  x774 & ~x312;
assign c2170 = ~x0 & ~x18 & ~x20 & ~x23 & ~x52 & ~x60 & ~x81 & ~x114 & ~x116 & ~x141 & ~x165 & ~x169 & ~x227 & ~x256 & ~x283 & ~x355 & ~x361 & ~x390 & ~x418 & ~x419 & ~x422 & ~x472 & ~x507 & ~x619 & ~x673 & ~x675 & ~x745 & ~x763 & ~x768 & ~x770;
assign c2172 =  x619;
assign c2174 =  x395 & ~x649;
assign c2176 =  x37 &  x47 &  x387 & ~x304;
assign c2178 =  x135 &  x556;
assign c2180 =  x105 &  x230 &  x460 &  x544 & ~x14 & ~x23 & ~x618;
assign c2182 = ~x34 & ~x106 & ~x153 & ~x275 & ~x305 & ~x334 & ~x391 & ~x421 & ~x423 & ~x445 & ~x472 & ~x501 & ~x502 & ~x505 & ~x507 & ~x528 & ~x533 & ~x562 & ~x614 & ~x618 & ~x641 & ~x644 & ~x746 & ~x770 & ~x771;
assign c2184 =  x413 & ~x5 & ~x52 & ~x56 & ~x85 & ~x114 & ~x410 & ~x417 & ~x450 & ~x670 & ~x755;
assign c2186 =  x37 &  x591 &  x619;
assign c2188 = ~x496;
assign c2190 =  x135;
assign c2192 =  x675 & ~x678;
assign c2194 = ~x271 & ~x330 & ~x409;
assign c2196 =  x129 &  x147 &  x204 &  x288 &  x296 &  x297 &  x300 &  x301 &  x322 &  x382 &  x404 &  x434 &  x494 &  x519 &  x547 &  x581 &  x750 & ~x22 & ~x110 & ~x138 & ~x200 & ~x360 & ~x365 & ~x504 & ~x775 & ~x779;
assign c2198 =  x290 & ~x111 & ~x523;
assign c2200 =  x11 &  x37 &  x189 &  x461 & ~x53 & ~x89 & ~x194 & ~x197 & ~x226 & ~x500 & ~x701;
assign c2202 =  x626 &  x710 &  x711 &  x715 & ~x54 & ~x104 & ~x219 & ~x255 & ~x275 & ~x303 & ~x335;
assign c2204 =  x76 &  x133 & ~x15 & ~x163;
assign c2206 =  x394;
assign c2208 =  x128 &  x316 &  x623 & ~x27 & ~x29 & ~x109 & ~x198 & ~x201 & ~x229 & ~x255 & ~x283 & ~x334 & ~x613 & ~x674 & ~x779;
assign c2210 = ~x8 & ~x35 & ~x78 & ~x110 & ~x185 & ~x186 & ~x254 & ~x309 & ~x333 & ~x339 & ~x360 & ~x388 & ~x396 & ~x416 & ~x417 & ~x444 & ~x473 & ~x480 & ~x507 & ~x534 & ~x587 & ~x760 & ~x770 & ~x782;
assign c2212 =  x423 & ~x677;
assign c2214 = ~x10 & ~x18 & ~x74 & ~x81 & ~x171 & ~x219 & ~x275 & ~x284 & ~x331 & ~x334 & ~x340 & ~x362 & ~x365 & ~x472 & ~x480 & ~x501 & ~x504 & ~x506 & ~x589 & ~x615 & ~x640 & ~x670 & ~x695 & ~x726;
assign c2216 =  x366;
assign c2218 = ~x20 & ~x25 & ~x30 & ~x56 & ~x140 & ~x172 & ~x185 & ~x193 & ~x197 & ~x200 & ~x215 & ~x251 & ~x419 & ~x445 & ~x502 & ~x507 & ~x615 & ~x644 & ~x645 & ~x725 & ~x758 & ~x765;
assign c2220 =  x765 &  x768 &  x772 &  x773 &  x774 & ~x6 & ~x78;
assign c2222 =  x131 &  x149 &  x522 &  x654 &  x656 & ~x58 & ~x78 & ~x249 & ~x278 & ~x388 & ~x391 & ~x416 & ~x559 & ~x726 & ~x742 & ~x743 & ~x745 & ~x758;
assign c2224 =  x173 &  x387 &  x668;
assign c2226 = ~x217 & ~x272 & ~x521;
assign c2228 =  x581 &  x749 & ~x118 & ~x162 & ~x172 & ~x227 & ~x247 & ~x275 & ~x283 & ~x303 & ~x396 & ~x443 & ~x723 & ~x770;
assign c2230 =  x454 & ~x483;
assign c2232 =  x246 & ~x15 & ~x58 & ~x200;
assign c2234 =  x190 &  x218 &  x245 &  x246 &  x413 &  x460 &  x489 &  x622 &  x750 & ~x170 & ~x192 & ~x222 & ~x668;
assign c2236 =  x40 & ~x30 & ~x56 & ~x68 & ~x170 & ~x227 & ~x390 & ~x474 & ~x698 & ~x728 & ~x770 & ~x773;
assign c2238 =  x614;
assign c2240 =  x134 &  x163 &  x556;
assign c2242 =  x133 &  x414 &  x470 & ~x15 & ~x83 & ~x165 & ~x276 & ~x280 & ~x417 & ~x505 & ~x531 & ~x613 & ~x757;
assign c2244 =  x367;
assign c2246 = ~x23 & ~x109 & ~x250 & ~x483 & ~x539 & ~x738 & ~x739 & ~x781;
assign c2248 =  x204 &  x693 & ~x60 & ~x118 & ~x275 & ~x283 & ~x309 & ~x396 & ~x480 & ~x773;
assign c2250 =  x72 &  x173 &  x398 &  x599 &  x686 & ~x200 & ~x364 & ~x423 & ~x619;
assign c2252 =  x16 &  x95 &  x486 &  x487 &  x519 &  x573 &  x622 &  x628 &  x658 &  x666 &  x711 &  x714 & ~x23 & ~x53 & ~x56 & ~x112 & ~x225 & ~x255 & ~x309 & ~x334 & ~x366 & ~x614 & ~x616 & ~x697 & ~x753;
assign c2254 =  x354 & ~x2 & ~x60 & ~x225 & ~x283 & ~x307 & ~x309 & ~x337 & ~x503 & ~x504 & ~x682 & ~x685 & ~x686 & ~x688 & ~x689 & ~x691 & ~x710 & ~x715 & ~x767;
assign c2256 =  x315 & ~x265 & ~x266 & ~x765;
assign c2258 = ~x244 & ~x446 & ~x464 & ~x547;
assign c2260 = ~x125 & ~x378 & ~x501 & ~x504 & ~x532;
assign c2262 = ~x418 & ~x503 & ~x570 & ~x571 & ~x574 & ~x578 & ~x644;
assign c2264 = ~x2 & ~x23 & ~x26 & ~x164 & ~x194 & ~x199 & ~x255 & ~x277 & ~x310 & ~x333 & ~x364 & ~x372 & ~x390 & ~x456 & ~x507 & ~x559 & ~x560 & ~x619 & ~x645 & ~x670 & ~x744 & ~x754 & ~x768 & ~x772;
assign c2266 =  x71 &  x100 &  x125 &  x204 &  x266 &  x314 &  x315 &  x317 &  x351 &  x398 &  x414 &  x433 &  x442 &  x462 &  x522 &  x538 &  x655 &  x657 &  x681 &  x750 & ~x20 & ~x22 & ~x31 & ~x33 & ~x51 & ~x58 & ~x59 & ~x79 & ~x80 & ~x88 & ~x105 & ~x171 & ~x249 & ~x255 & ~x282 & ~x306 & ~x310 & ~x332 & ~x360 & ~x391 & ~x418 & ~x445 & ~x477 & ~x532 & ~x617 & ~x643 & ~x645 & ~x698 & ~x729 & ~x730 & ~x766 & ~x771;
assign c2268 =  x92 &  x94 &  x133 &  x202 &  x215 &  x258 &  x264 &  x287 &  x322 &  x385 &  x403 &  x633 &  x681 &  x685 & ~x166 & ~x168 & ~x195 & ~x224 & ~x227 & ~x304 & ~x311 & ~x393 & ~x504 & ~x585 & ~x591 & ~x700 & ~x726 & ~x754;
assign c2270 = ~x1 & ~x5 & ~x25 & ~x30 & ~x32 & ~x33 & ~x36 & ~x47 & ~x48 & ~x54 & ~x56 & ~x57 & ~x74 & ~x77 & ~x80 & ~x86 & ~x87 & ~x88 & ~x102 & ~x103 & ~x104 & ~x110 & ~x112 & ~x113 & ~x116 & ~x133 & ~x140 & ~x144 & ~x164 & ~x169 & ~x172 & ~x192 & ~x220 & ~x222 & ~x250 & ~x276 & ~x279 & ~x282 & ~x304 & ~x305 & ~x307 & ~x337 & ~x360 & ~x361 & ~x365 & ~x417 & ~x421 & ~x422 & ~x446 & ~x479 & ~x502 & ~x534 & ~x556 & ~x557 & ~x559 & ~x586 & ~x587 & ~x588 & ~x590 & ~x614 & ~x615 & ~x642 & ~x644 & ~x671 & ~x673 & ~x700 & ~x725 & ~x726 & ~x729 & ~x753 & ~x759 & ~x760 & ~x771 & ~x782;
assign c2272 =  x173 &  x722 &  x778 & ~x227 & ~x283 & ~x312;
assign c2274 = ~x60 & ~x75 & ~x79 & ~x84 & ~x104 & ~x165 & ~x302 & ~x495 & ~x507;
assign c2276 =  x201 &  x328 &  x695 & ~x89 & ~x196 & ~x451 & ~x504 & ~x672 & ~x707 & ~x770;
assign c2278 = ~x103 & ~x151 & ~x186 & ~x361 & ~x417 & ~x477 & ~x500 & ~x530 & ~x762;
assign c2280 =  x175 & ~x84 & ~x109 & ~x193 & ~x200 & ~x221 & ~x304 & ~x616 & ~x661 & ~x759;
assign c2282 =  x158 &  x204 &  x402 &  x434 &  x491 &  x492 &  x514 &  x569 &  x605 &  x625 &  x632 &  x651 & ~x6 & ~x54 & ~x59 & ~x111 & ~x115 & ~x141 & ~x144 & ~x227 & ~x229 & ~x303 & ~x360 & ~x362 & ~x387 & ~x396 & ~x421 & ~x473 & ~x476 & ~x558 & ~x584 & ~x591 & ~x644;
assign c2284 =  x706 & ~x191 & ~x229 & ~x275 & ~x535 & ~x613 & ~x710 & ~x714 & ~x717;
assign c2286 =  x731 & ~x566 & ~x678 & ~x758;
assign c2288 =  x711 &  x745 &  x746 & ~x27 & ~x103 & ~x107 & ~x136 & ~x558 & ~x673;
assign c2290 = ~x2 & ~x21 & ~x22 & ~x25 & ~x49 & ~x57 & ~x141 & ~x192 & ~x224 & ~x225 & ~x249 & ~x250 & ~x277 & ~x279 & ~x281 & ~x364 & ~x448 & ~x528 & ~x552 & ~x729 & ~x740 & ~x742 & ~x767 & ~x773;
assign c2292 =  x44 & ~x294 & ~x464 & ~x492;
assign c2294 =  x314 & ~x3 & ~x32 & ~x53 & ~x85 & ~x166 & ~x168 & ~x210 & ~x222 & ~x226 & ~x250 & ~x252 & ~x306 & ~x309 & ~x391 & ~x392 & ~x449 & ~x478 & ~x533 & ~x558 & ~x674 & ~x726;
assign c2296 = ~x78 & ~x112 & ~x178 & ~x184 & ~x185 & ~x186 & ~x195 & ~x199 & ~x222 & ~x249 & ~x252 & ~x255 & ~x276 & ~x278 & ~x304 & ~x307 & ~x333 & ~x362 & ~x367 & ~x390 & ~x395 & ~x416 & ~x450 & ~x479 & ~x501 & ~x505 & ~x530 & ~x532 & ~x643 & ~x697 & ~x770 & ~x772;
assign c2298 =  x581 & ~x0 & ~x9 & ~x279 & ~x361 & ~x392 & ~x495 & ~x523;
assign c2300 =  x583 &  x772 &  x775;
assign c2302 = ~x29 & ~x78 & ~x110 & ~x138 & ~x143 & ~x163 & ~x167 & ~x171 & ~x248 & ~x249 & ~x275 & ~x279 & ~x283 & ~x303 & ~x310 & ~x313 & ~x333 & ~x367 & ~x389 & ~x393 & ~x444 & ~x449 & ~x477 & ~x501 & ~x502 & ~x507 & ~x563 & ~x619 & ~x646 & ~x673 & ~x697 & ~x710 & ~x712 & ~x714 & ~x716 & ~x717 & ~x740 & ~x741 & ~x746 & ~x754 & ~x767 & ~x768;
assign c2304 =  x37 & ~x15 & ~x84 & ~x136 & ~x169 & ~x191 & ~x283 & ~x673 & ~x702 & ~x724 & ~x726 & ~x759 & ~x773;
assign c2306 =  x75 &  x244 &  x414 &  x463 &  x509 &  x516 &  x521 &  x543 & ~x14 & ~x15 & ~x22 & ~x83 & ~x109 & ~x168 & ~x200 & ~x227 & ~x445 & ~x476 & ~x529 & ~x646 & ~x699;
assign c2308 = ~x56 & ~x103 & ~x104 & ~x105 & ~x116 & ~x133 & ~x140 & ~x145 & ~x162 & ~x275 & ~x284 & ~x446 & ~x473 & ~x474 & ~x477 & ~x507 & ~x533 & ~x592 & ~x667 & ~x732 & ~x779 & ~x783;
assign c2310 = ~x7 & ~x78 & ~x84 & ~x88 & ~x107 & ~x111 & ~x137 & ~x138 & ~x163 & ~x178 & ~x179 & ~x185 & ~x191 & ~x220 & ~x227 & ~x228 & ~x255 & ~x276 & ~x281 & ~x309 & ~x332 & ~x334 & ~x360 & ~x363 & ~x389 & ~x391 & ~x422 & ~x423 & ~x446 & ~x502 & ~x505 & ~x528 & ~x646 & ~x673 & ~x726 & ~x758 & ~x765;
assign c2312 =  x42 & ~x25 & ~x26 & ~x31 & ~x66 & ~x100 & ~x103 & ~x104 & ~x227 & ~x250 & ~x283 & ~x390 & ~x393 & ~x423 & ~x446 & ~x450 & ~x476 & ~x501 & ~x674 & ~x701;
assign c2314 =  x749 &  x777 & ~x199 & ~x275 & ~x367 & ~x444 & ~x480 & ~x648 & ~x770 & ~x772;
assign c2316 =  x76 & ~x169 & ~x283 & ~x390 & ~x745;
assign c2318 = ~x0 & ~x2 & ~x144 & ~x195 & ~x198 & ~x226 & ~x254 & ~x255 & ~x276 & ~x279 & ~x283 & ~x335 & ~x389 & ~x395 & ~x445 & ~x449 & ~x474 & ~x505 & ~x507 & ~x529 & ~x530 & ~x557 & ~x567 & ~x595 & ~x670 & ~x675 & ~x698 & ~x703 & ~x740 & ~x745 & ~x747 & ~x769;
assign c2320 =  x144 &  x675;
assign c2322 = ~x266 & ~x322 & ~x334 & ~x350 & ~x351 & ~x474 & ~x504;
assign c2324 =  x173 &  x244 &  x407 &  x426 &  x549 &  x576 &  x648 & ~x6 & ~x24 & ~x34 & ~x58 & ~x227 & ~x333 & ~x531;
assign c2326 =  x76 &  x161 &  x458 &  x463 &  x487 &  x594 & ~x4 & ~x198 & ~x255 & ~x283 & ~x304;
assign c2328 =  x175 &  x341 &  x375 &  x526 &  x549 &  x751 &  x779 & ~x80 & ~x109 & ~x226 & ~x283;
assign c2330 =  x124 &  x330 &  x385 &  x434 &  x463 &  x549 &  x577 &  x654 &  x687 &  x710 &  x778 & ~x27 & ~x33 & ~x53 & ~x110 & ~x194 & ~x200 & ~x276 & ~x278 & ~x335 & ~x363 & ~x388 & ~x446 & ~x449 & ~x618;
assign c2332 =  x68 &  x349 &  x352 &  x684 & ~x0 & ~x191 & ~x277 & ~x283 & ~x480 & ~x588 & ~x726 & ~x756 & ~x777;
assign c2334 = ~x245 & ~x515 & ~x545;
assign c2336 =  x563 &  x647 & ~x14;
assign c2338 =  x641;
assign c2340 =  x62 & ~x504 & ~x559 & ~x770;
assign c2342 = ~x78 & ~x103 & ~x302 & ~x428;
assign c2344 =  x200;
assign c2346 = ~x4 & ~x32 & ~x52 & ~x56 & ~x81 & ~x87 & ~x138 & ~x221 & ~x252 & ~x253 & ~x277 & ~x279 & ~x305 & ~x333 & ~x335 & ~x337 & ~x399 & ~x427 & ~x502 & ~x530 & ~x531 & ~x588 & ~x644 & ~x738 & ~x767;
assign c2348 =  x37 &  x46 &  x260 &  x356 &  x404 &  x582 & ~x416;
assign c2350 =  x11 &  x62 &  x398;
assign c2352 = ~x1 & ~x20 & ~x22 & ~x25 & ~x30 & ~x54 & ~x58 & ~x79 & ~x81 & ~x82 & ~x86 & ~x87 & ~x104 & ~x107 & ~x113 & ~x115 & ~x137 & ~x169 & ~x199 & ~x213 & ~x334 & ~x390 & ~x421 & ~x422 & ~x447 & ~x474 & ~x518 & ~x521 & ~x534 & ~x589 & ~x614 & ~x644 & ~x646 & ~x671 & ~x673 & ~x726 & ~x727 & ~x756 & ~x757;
assign c2354 =  x161 &  x244 &  x407 &  x462 &  x778 & ~x5 & ~x86 & ~x111 & ~x275 & ~x360 & ~x503 & ~x506 & ~x534 & ~x700 & ~x729;
assign c2356 =  x228 &  x368;
assign c2358 =  x367;
assign c2360 =  x76 &  x133 &  x160 &  x189 &  x301 &  x399 &  x434 & ~x34 & ~x227 & ~x311 & ~x394 & ~x479 & ~x561 & ~x589;
assign c2362 = ~x30 & ~x61 & ~x66 & ~x78 & ~x79 & ~x91 & ~x111 & ~x119 & ~x163 & ~x220 & ~x251 & ~x283 & ~x333 & ~x337 & ~x361 & ~x390 & ~x392 & ~x419 & ~x445 & ~x500 & ~x559 & ~x726 & ~x727 & ~x740 & ~x741 & ~x744 & ~x745 & ~x766 & ~x769 & ~x775;
assign c2364 = ~x191 & ~x220 & ~x275 & ~x654 & ~x656 & ~x660 & ~x661 & ~x662 & ~x683 & ~x686 & ~x689 & ~x745 & ~x770 & ~x775;
assign c2366 =  x200 &  x396;
assign c2368 = ~x22 & ~x31 & ~x32 & ~x55 & ~x80 & ~x85 & ~x104 & ~x167 & ~x281 & ~x333 & ~x347 & ~x350 & ~x446 & ~x529 & ~x533 & ~x561 & ~x729 & ~x757;
assign c2370 = ~x0 & ~x8 & ~x9 & ~x21 & ~x25 & ~x28 & ~x33 & ~x35 & ~x48 & ~x50 & ~x55 & ~x57 & ~x61 & ~x81 & ~x82 & ~x83 & ~x85 & ~x110 & ~x115 & ~x136 & ~x138 & ~x139 & ~x140 & ~x142 & ~x163 & ~x185 & ~x195 & ~x198 & ~x200 & ~x227 & ~x228 & ~x248 & ~x255 & ~x278 & ~x279 & ~x284 & ~x304 & ~x311 & ~x334 & ~x336 & ~x360 & ~x365 & ~x388 & ~x390 & ~x391 & ~x395 & ~x416 & ~x422 & ~x423 & ~x444 & ~x446 & ~x451 & ~x472 & ~x473 & ~x501 & ~x503 & ~x506 & ~x530 & ~x533 & ~x561 & ~x563 & ~x589 & ~x612 & ~x613 & ~x643 & ~x644 & ~x646 & ~x669 & ~x675 & ~x699 & ~x701 & ~x731 & ~x753 & ~x755 & ~x759 & ~x760 & ~x771 & ~x775 & ~x780 & ~x783;
assign c2372 =  x189 &  x288 &  x463 & ~x192 & ~x219 & ~x276 & ~x285 & ~x312;
assign c2374 =  x444 & ~x15 & ~x31;
assign c2376 =  x37 &  x648 &  x716;
assign c2378 =  x520 &  x663 &  x779 & ~x54 & ~x170 & ~x227 & ~x735;
assign c2380 = ~x59 & ~x226 & ~x306 & ~x316 & ~x333 & ~x344 & ~x419 & ~x450 & ~x559 & ~x642 & ~x767 & ~x781;
assign c2382 = ~x7 & ~x9 & ~x19 & ~x23 & ~x32 & ~x36 & ~x103 & ~x104 & ~x107 & ~x135 & ~x162 & ~x164 & ~x169 & ~x173 & ~x190 & ~x192 & ~x196 & ~x201 & ~x225 & ~x246 & ~x275 & ~x284 & ~x302 & ~x303 & ~x332 & ~x338 & ~x395 & ~x396 & ~x415 & ~x477 & ~x502 & ~x506 & ~x508 & ~x557 & ~x558 & ~x562 & ~x585 & ~x591 & ~x612 & ~x639 & ~x642 & ~x673 & ~x726 & ~x779;
assign c2384 =  x618;
assign c2386 =  x189 &  x257 &  x322 &  x683 &  x695 &  x710 &  x714 & ~x82 & ~x85 & ~x107 & ~x250 & ~x361 & ~x448;
assign c2388 =  x173 &  x425 & ~x395 & ~x618 & ~x619 & ~x641;
assign c2390 = ~x271 & ~x434 & ~x464 & ~x492 & ~x521 & ~x549;
assign c2392 =  x462 & ~x21 & ~x61 & ~x116 & ~x192 & ~x226 & ~x312 & ~x423 & ~x679 & ~x707 & ~x745 & ~x774;
assign c2394 =  x427 & ~x27 & ~x193 & ~x200 & ~x392 & ~x416 & ~x513 & ~x530 & ~x535 & ~x556 & ~x557 & ~x647 & ~x758 & ~x782;
assign c2396 =  x187 &  x218 &  x627 &  x715 & ~x54 & ~x107 & ~x192 & ~x252 & ~x752 & ~x759 & ~x769;
assign c2398 =  x37 &  x132 &  x458 &  x554 &  x571 & ~x57 & ~x60 & ~x88 & ~x109 & ~x140 & ~x196 & ~x390 & ~x392 & ~x393 & ~x504 & ~x588 & ~x671 & ~x701 & ~x763;
assign c2400 =  x244 &  x458 &  x517 &  x573 &  x633 &  x651 & ~x54 & ~x145 & ~x164 & ~x166 & ~x171 & ~x227 & ~x419 & ~x583;
assign c2402 =  x327 &  x350 &  x377 &  x577 & ~x8 & ~x163 & ~x164 & ~x172 & ~x224 & ~x275 & ~x276 & ~x303 & ~x334 & ~x340 & ~x360 & ~x364 & ~x366 & ~x391 & ~x396 & ~x422 & ~x449 & ~x480 & ~x536 & ~x555 & ~x611 & ~x667 & ~x676 & ~x696 & ~x700;
assign c2404 =  x69 &  x161 &  x291 &  x427 &  x463 &  x484 &  x681 &  x711 &  x745 & ~x88 & ~x166 & ~x171 & ~x227 & ~x367 & ~x395 & ~x445 & ~x473 & ~x613 & ~x617 & ~x641 & ~x670 & ~x729;
assign c2406 = ~x128 & ~x530 & ~x572 & ~x574;
assign c2408 = ~x25 & ~x73 & ~x82 & ~x98 & ~x140 & ~x143 & ~x196 & ~x199 & ~x226 & ~x248 & ~x281 & ~x283 & ~x335 & ~x417 & ~x418 & ~x422 & ~x448 & ~x474 & ~x501 & ~x503 & ~x504 & ~x534 & ~x765 & ~x766 & ~x767;
assign c2410 =  x129 & ~x139 & ~x162 & ~x171 & ~x173 & ~x218 & ~x246 & ~x250 & ~x312 & ~x340 & ~x502 & ~x535 & ~x589 & ~x730 & ~x732;
assign c2412 =  x273 &  x300 &  x649 &  x687 &  x711 &  x750 & ~x88 & ~x199 & ~x256 & ~x275 & ~x283;
assign c2414 =  x201 &  x441 &  x733 & ~x3 & ~x21 & ~x27 & ~x32 & ~x110 & ~x172 & ~x192 & ~x305 & ~x393 & ~x645 & ~x679 & ~x700 & ~x703 & ~x754 & ~x767;
assign c2416 =  x76 &  x256 &  x368;
assign c2418 =  x128 &  x259 &  x347 &  x410 &  x458 &  x511 &  x600 &  x632 &  x686 &  x716 & ~x4 & ~x52 & ~x78 & ~x90 & ~x104 & ~x200 & ~x311 & ~x448 & ~x531 & ~x586 & ~x780;
assign c2420 =  x380 & ~x66 & ~x107 & ~x256 & ~x275 & ~x564;
assign c2422 =  x641;
assign c2424 = ~x3 & ~x97 & ~x141 & ~x248 & ~x250 & ~x305 & ~x334 & ~x422 & ~x474 & ~x505 & ~x506 & ~x571 & ~x616 & ~x726;
assign c2426 =  x147 &  x230 &  x762 & ~x48 & ~x110 & ~x275 & ~x312 & ~x445 & ~x507 & ~x588 & ~x612 & ~x615 & ~x640 & ~x675 & ~x702;
assign c2428 =  x247 &  x640 &  x742;
assign c2430 =  x72 &  x155 &  x158 &  x232 &  x483 &  x762 & ~x0 & ~x1 & ~x24 & ~x27 & ~x34 & ~x51 & ~x57 & ~x168 & ~x200 & ~x284 & ~x387 & ~x506 & ~x584 & ~x612;
assign c2432 =  x104 &  x439 & ~x284 & ~x390 & ~x710 & ~x717 & ~x719 & ~x743;
assign c2434 =  x10 &  x16 &  x37 &  x330 &  x683;
assign c2436 =  x300 &  x357 &  x386 &  x398 &  x410 &  x434 &  x458 &  x510 &  x571 &  x683 &  x711 &  x750 & ~x0 & ~x26 & ~x27 & ~x113 & ~x172 & ~x252 & ~x275 & ~x276 & ~x283 & ~x304 & ~x305;
assign c2438 =  x91 &  x98 &  x243 &  x264 &  x299 &  x345 &  x439 &  x493 &  x519 & ~x78 & ~x200 & ~x332 & ~x335 & ~x395 & ~x444 & ~x507 & ~x668 & ~x726 & ~x753 & ~x781;
assign c2440 =  x117 &  x368 & ~x535;
assign c2442 = ~x135 & ~x223 & ~x248 & ~x388 & ~x446 & ~x477 & ~x479 & ~x504 & ~x531 & ~x535 & ~x558 & ~x561 & ~x595 & ~x615 & ~x651 & ~x737 & ~x742 & ~x744 & ~x746 & ~x756 & ~x763 & ~x764 & ~x768 & ~x772 & ~x773;
assign c2444 =  x245 &  x370 &  x375 &  x462 &  x655 & ~x276 & ~x278 & ~x281 & ~x559 & ~x595 & ~x770;
assign c2446 =  x175 &  x177 &  x189 &  x216 &  x298 &  x372 &  x380 &  x405 &  x414 &  x442 &  x483 &  x498 &  x511 &  x542 &  x547 &  x567 &  x604 &  x655 &  x682 &  x722 & ~x221 & ~x283 & ~x307 & ~x309 & ~x312 & ~x368 & ~x447 & ~x449 & ~x451 & ~x612 & ~x616 & ~x670 & ~x672 & ~x703 & ~x730 & ~x754 & ~x757 & ~x760;
assign c2448 = ~x0 & ~x22 & ~x33 & ~x52 & ~x82 & ~x87 & ~x110 & ~x116 & ~x138 & ~x213 & ~x215 & ~x243 & ~x255 & ~x282 & ~x309 & ~x337 & ~x339 & ~x360 & ~x391 & ~x445 & ~x449 & ~x452 & ~x505 & ~x531 & ~x700 & ~x702 & ~x730 & ~x758 & ~x767 & ~x768;
assign c2450 =  x69 &  x295 &  x296 &  x297 &  x301 &  x378 &  x406 &  x441 &  x454 &  x489 &  x511 &  x515 &  x526 &  x545 &  x549 &  x554 &  x566 &  x570 &  x595 &  x679 &  x706 & ~x2 & ~x5 & ~x8 & ~x80 & ~x108 & ~x139 & ~x166 & ~x197 & ~x220 & ~x222 & ~x229 & ~x277 & ~x312 & ~x338 & ~x392 & ~x417 & ~x446 & ~x448 & ~x559 & ~x586 & ~x726;
assign c2452 =  x37 &  x472 &  x500 &  x528 & ~x58;
assign c2454 =  x297 &  x409 &  x543 & ~x171 & ~x200 & ~x528 & ~x614 & ~x645 & ~x710 & ~x712 & ~x719 & ~x730 & ~x731 & ~x741 & ~x745;
assign c2456 = ~x433 & ~x434 & ~x439 & ~x493 & ~x767 & ~x770;
assign c2458 = ~x272 & ~x455;
assign c2460 =  x106 & ~x33 & ~x59 & ~x391 & ~x757;
assign c2462 =  x144;
assign c2464 =  x648 &  x767;
assign c2466 =  x200 &  x228 &  x340 &  x396;
assign c2468 =  x121 &  x542 &  x722 & ~x107 & ~x228 & ~x229 & ~x275 & ~x303 & ~x702;
assign c2470 =  x534;
assign c2472 =  x395;
assign c2474 =  x173 &  x577 &  x599 &  x621 &  x648 & ~x591;
assign c2476 =  x458 & ~x53 & ~x282 & ~x444 & ~x533 & ~x561 & ~x707 & ~x724 & ~x738 & ~x741 & ~x747;
assign c2478 =  x776;
assign c2480 =  x15 &  x189 &  x438 &  x470 &  x554 &  x576 &  x630 &  x658 &  x750 &  x778 & ~x34 & ~x51 & ~x87 & ~x116 & ~x194 & ~x249 & ~x311 & ~x333 & ~x367 & ~x697 & ~x699 & ~x701 & ~x728 & ~x780 & ~x782;
assign c2482 = ~x35 & ~x56 & ~x83 & ~x170 & ~x199 & ~x200 & ~x218 & ~x227 & ~x254 & ~x277 & ~x282 & ~x302 & ~x330 & ~x331 & ~x361 & ~x362 & ~x368 & ~x505 & ~x529 & ~x592 & ~x738 & ~x740 & ~x742 & ~x745 & ~x757 & ~x782;
assign c2484 =  x121 &  x152 &  x160 &  x300 &  x549 &  x573 &  x693 & ~x162 & ~x172 & ~x219 & ~x227 & ~x256 & ~x275 & ~x283 & ~x303 & ~x387 & ~x500 & ~x591 & ~x671 & ~x753 & ~x775;
assign c2486 =  x367;
assign c2488 = ~x151 & ~x153 & ~x154 & ~x275 & ~x303 & ~x331 & ~x333 & ~x423 & ~x534 & ~x585 & ~x645 & ~x646 & ~x742 & ~x770;
assign c2490 =  x90 & ~x227 & ~x742 & ~x770;
assign c2492 =  x69 &  x175 &  x413 &  x442 &  x463 &  x492 &  x762 & ~x23 & ~x28 & ~x83 & ~x105 & ~x108 & ~x199 & ~x253 & ~x284 & ~x335 & ~x337 & ~x417 & ~x530 & ~x559 & ~x591 & ~x614 & ~x780;
assign c2494 =  x200 &  x642;
assign c2496 =  x204 &  x270 &  x288 &  x385 &  x400 &  x434 &  x493 &  x516 &  x656 &  x711 &  x714 &  x715 & ~x56 & ~x104 & ~x171 & ~x253 & ~x311 & ~x334 & ~x587 & ~x730;
assign c2498 =  x70 &  x302 &  x432 &  x463 &  x571 &  x655 &  x779 & ~x83 & ~x283 & ~x335 & ~x590 & ~x755;
assign c21 = ~x11 & ~x39 & ~x47;
assign c23 =  x109;
assign c25 =  x182 &  x267 &  x329 &  x342 &  x353 &  x372 &  x407 &  x409 &  x427 &  x437 &  x483 &  x495 &  x499 &  x521 &  x552 &  x580 &  x594 &  x624 &  x651 &  x663 &  x677 &  x679 &  x692 &  x720 & ~x3 & ~x110 & ~x116 & ~x390 & ~x391 & ~x417 & ~x420 & ~x587;
assign c27 =  x39 &  x45 &  x67 &  x213 &  x216 &  x232 &  x237 &  x273 &  x342 &  x374 &  x406 &  x413 &  x440 &  x467 &  x483 &  x487 &  x496 &  x525 &  x537 &  x552 &  x611 &  x637 &  x652 &  x679 &  x707 & ~x137 & ~x500 & ~x534 & ~x561 & ~x563 & ~x586 & ~x755;
assign c29 =  x39 & ~x452 & ~x453 & ~x565 & ~x592 & ~x610 & ~x733;
assign c211 =  x93 &  x99 &  x147 &  x149 &  x155 &  x158 &  x180 &  x203 &  x236 &  x262 &  x324 &  x326 &  x350 &  x380 &  x386 &  x398 &  x399 &  x403 &  x429 &  x430 &  x431 &  x441 &  x454 &  x462 &  x466 &  x515 &  x537 &  x578 &  x583 &  x600 &  x637 &  x665 &  x676 & ~x10 & ~x18 & ~x36 & ~x46 & ~x47 & ~x51 & ~x54 & ~x89 & ~x106 & ~x167 & ~x278 & ~x365 & ~x392 & ~x501 & ~x503 & ~x530 & ~x587 & ~x669 & ~x699 & ~x700 & ~x702 & ~x754 & ~x783;
assign c213 =  x166;
assign c215 =  x156 &  x186 &  x210 &  x327 &  x354 &  x376 &  x465 &  x580 &  x693 &  x734 &  x761 & ~x736;
assign c217 =  x44 &  x190 & ~x442 & ~x453 & ~x498 & ~x611 & ~x733;
assign c219 = ~x39;
assign c221 = ~x385 & ~x553;
assign c225 =  x502;
assign c227 =  x278;
assign c229 =  x32;
assign c231 =  x362;
assign c233 =  x57;
assign c235 =  x447;
assign c237 =  x2;
assign c239 =  x194;
assign c241 = ~x44;
assign c243 = ~x442 & ~x470 & ~x526 & ~x553 & ~x583 & ~x694 & ~x732;
assign c245 =  x92 &  x97 &  x157 &  x177 &  x208 &  x213 &  x272 &  x292 &  x318 &  x325 &  x345 &  x355 &  x356 &  x379 &  x409 &  x410 &  x464 &  x482 &  x565 & ~x36 & ~x46 & ~x47 & ~x77 & ~x113 & ~x141 & ~x168 & ~x278 & ~x391 & ~x475 & ~x476 & ~x562 & ~x614 & ~x615 & ~x674 & ~x766;
assign c247 = ~x17 & ~x36 & ~x45;
assign c249 =  x55;
assign c251 = ~x45 & ~x47 & ~x121;
assign c253 = ~x414 & ~x593 & ~x608;
assign c255 = ~x636 & ~x637 & ~x751;
assign c257 =  x335;
assign c259 =  x391;
assign c261 =  x12 &  x39 &  x189 &  x213 &  x271 &  x294 &  x371 &  x377 &  x412 &  x443 &  x569 &  x620 & ~x47 & ~x63 & ~x142 & ~x529 & ~x587 & ~x700;
assign c263 =  x285 &  x319 &  x325 &  x327 &  x347 &  x356 &  x373 &  x376 &  x379 &  x383 &  x384 &  x414 &  x433 &  x436 &  x470 &  x485 &  x508 &  x509 &  x526 &  x527 &  x545 &  x565 &  x577 &  x606 &  x610 &  x635 & ~x17 & ~x36 & ~x46 & ~x57 & ~x111 & ~x168 & ~x224 & ~x365 & ~x392 & ~x502 & ~x503 & ~x531 & ~x532 & ~x644 & ~x776;
assign c265 = ~x342 & ~x371;
assign c267 =  x12 &  x205 &  x208 &  x234 &  x400 &  x495 &  x516 &  x541 &  x599 &  x611 &  x636 &  x652 &  x659 &  x734 & ~x47 & ~x59 & ~x77 & ~x113 & ~x362 & ~x559 & ~x698;
assign c269 =  x153 &  x188 &  x285 &  x350 &  x354 &  x676 & ~x31 & ~x47 & ~x766;
assign c271 =  x140;
assign c273 =  x447;
assign c275 =  x83;
assign c277 =  x447;
assign c279 =  x466 &  x524 &  x761 & ~x36 & ~x47 & ~x736;
assign c281 =  x644;
assign c283 = ~x42 & ~x96;
assign c285 =  x587;
assign c287 = ~x17 & ~x36 & ~x45 & ~x46 & ~x48 & ~x251 & ~x636;
assign c289 =  x477;
assign c291 =  x399 &  x429 &  x468 &  x496 &  x513 &  x524 &  x538 &  x594 &  x601 &  x637 & ~x7 & ~x17 & ~x19 & ~x35 & ~x45 & ~x46 & ~x47 & ~x55;
assign c293 =  x361;
assign c295 = ~x14 & ~x39;
assign c297 = ~x234 & ~x329 & ~x385;
assign c299 =  x52;
assign c2101 =  x169;
assign c2103 =  x55;
assign c2105 =  x93 &  x179 &  x744 & ~x82 & ~x251 & ~x390 & ~x478 & ~x620 & ~x649 & ~x668 & ~x675 & ~x695 & ~x696 & ~x702 & ~x704 & ~x728 & ~x732 & ~x733 & ~x755;
assign c2107 =  x86;
assign c2109 =  x6;
assign c2111 =  x82;
assign c2113 =  x41 & ~x453 & ~x481 & ~x498 & ~x565 & ~x733;
assign c2117 =  x166;
assign c2119 = ~x120 & ~x175 & ~x202;
assign c2121 =  x194;
assign c2123 =  x83;
assign c2125 = ~x42;
assign c2127 = ~x413 & ~x426;
assign c2129 =  x66 &  x184 &  x210 &  x215 &  x327 &  x354 &  x405 &  x508 &  x537 &  x553 & ~x3 & ~x7 & ~x36 & ~x46 & ~x116 & ~x333 & ~x474 & ~x501 & ~x589;
assign c2131 = ~x291 & ~x684;
assign c2133 =  x448;
assign c2135 =  x13 &  x92 &  x154 &  x180 &  x262 &  x269 &  x314 &  x322 &  x324 &  x328 &  x347 &  x522 &  x537 & ~x1 & ~x4 & ~x18 & ~x46 & ~x47 & ~x58 & ~x77 & ~x87 & ~x112 & ~x279 & ~x473 & ~x617 & ~x776;
assign c2137 = ~x37 & ~x45 & ~x47 & ~x148;
assign c2139 =  x114;
assign c2141 =  x137;
assign c2143 =  x99 &  x126 &  x181 &  x207 &  x466 &  x492 & ~x587 & ~x610 & ~x649 & ~x705;
assign c2145 =  x336;
assign c2147 =  x392;
assign c2149 = ~x233 & ~x262;
assign c2151 =  x34 &  x35 &  x48 &  x127 &  x623;
assign c2153 =  x181 &  x386 &  x536 &  x552 &  x554 &  x676 & ~x36 & ~x58 & ~x673 & ~x720;
assign c2155 =  x169;
assign c2157 = ~x526 & ~x555 & ~x580 & ~x607;
assign c2159 =  x307;
assign c2161 =  x52;
assign c2163 =  x66 &  x102 &  x124 &  x154 &  x157 &  x179 &  x185 &  x209 &  x233 &  x235 &  x265 &  x270 &  x271 &  x287 &  x315 &  x318 &  x321 &  x345 &  x353 &  x354 &  x372 &  x375 &  x382 &  x433 &  x461 &  x463 &  x466 &  x483 &  x488 &  x511 &  x517 &  x523 &  x568 &  x572 &  x580 &  x626 &  x634 &  x636 &  x652 &  x657 &  x683 &  x684 &  x687 &  x690 &  x692 &  x709 &  x710 &  x717 &  x720 &  x738 &  x741 &  x742 & ~x23 & ~x30 & ~x86 & ~x108 & ~x136 & ~x194 & ~x226 & ~x308 & ~x392 & ~x504 & ~x531 & ~x557 & ~x643 & ~x674 & ~x729 & ~x756 & ~x781;
assign c2165 =  x32;
assign c2167 =  x447;
assign c2169 =  x59;
assign c2171 = ~x463 & ~x684;
assign c2173 = ~x413;
assign c2175 =  x250;
assign c2177 =  x363;
assign c2179 =  x109;
assign c2181 =  x551 &  x552 &  x691 & ~x453 & ~x668 & ~x676;
assign c2183 = ~x315 & ~x485;
assign c2185 = ~x553 & ~x554 & ~x611 & ~x636;
assign c2187 = ~x17;
assign c2189 = ~x607 & ~x636;
assign c2191 =  x195;
assign c2193 =  x308;
assign c2195 =  x59;
assign c2197 =  x96 &  x150 &  x234 &  x273 &  x348 &  x374 &  x429 &  x469 &  x522 &  x524 &  x568 &  x570 &  x637 &  x652 &  x658 &  x665 &  x692 &  x717 &  x736 & ~x2 & ~x4 & ~x31 & ~x167 & ~x198 & ~x472;
assign c2199 =  x41 &  x151 &  x154 &  x210 &  x213 &  x406 &  x457 &  x496 &  x539 &  x552 &  x580 &  x636 & ~x18 & ~x559 & ~x733;
assign c2201 =  x152 &  x374 &  x436 &  x468 &  x579 &  x664 & ~x139 & ~x341;
assign c2203 =  x12 &  x42 &  x66 &  x125 &  x241 &  x242 &  x246 &  x293 &  x299 &  x301 &  x353 &  x401 &  x415 &  x431 &  x457 &  x465 &  x482 &  x498 &  x517 &  x633 &  x682 & ~x47 & ~x48 & ~x85 & ~x112 & ~x170 & ~x221 & ~x339 & ~x529 & ~x615;
assign c2205 = ~x37 & ~x38 & ~x289;
assign c2207 = ~x47 & ~x262;
assign c2209 = ~x596 & ~x636 & ~x637;
assign c2211 =  x411 & ~x175 & ~x230;
assign c2213 = ~x371 & ~x453 & ~x565;
assign c2215 =  x700;
assign c2217 =  x4;
assign c2219 =  x134 & ~x397 & ~x453 & ~x481 & ~x509 & ~x704;
assign c2221 =  x55;
assign c2225 =  x221;
assign c2227 =  x365;
assign c2229 =  x316 & ~x2 & ~x6 & ~x10 & ~x11 & ~x17 & ~x36 & ~x45 & ~x46 & ~x47 & ~x113 & ~x141 & ~x450 & ~x615 & ~x617 & ~x618 & ~x647 & ~x697 & ~x726 & ~x727 & ~x765;
assign c2231 =  x109;
assign c2233 =  x38 & ~x470;
assign c2235 =  x353 &  x372 &  x432 &  x459 &  x471 &  x496 &  x511 &  x537 &  x580 &  x607 &  x626 &  x627 &  x634 &  x636 &  x639 &  x653 &  x655 &  x659 & ~x11 & ~x17 & ~x18 & ~x22 & ~x56 & ~x84 & ~x116 & ~x165 & ~x225 & ~x700;
assign c2237 = ~x517;
assign c2239 =  x502;
assign c2241 =  x13 &  x238 &  x269 &  x271 &  x292 &  x319 &  x373 &  x523 &  x552 &  x574 &  x630 &  x656 & ~x17 & ~x19 & ~x36 & ~x47 & ~x115 & ~x192 & ~x251 & ~x279;
assign c2243 =  x440 & ~x39;
assign c2245 =  x12 &  x14 &  x93 &  x94 &  x97 &  x130 &  x146 &  x153 &  x156 &  x179 &  x180 &  x185 &  x190 &  x209 &  x212 &  x260 &  x343 &  x353 &  x356 &  x371 &  x378 &  x401 &  x410 &  x413 &  x429 &  x457 &  x491 &  x510 &  x523 &  x632 &  x637 & ~x47 & ~x114 & ~x249 & ~x252 & ~x279 & ~x305 & ~x393 & ~x473 & ~x505 & ~x561 & ~x616 & ~x617;
assign c2247 =  x456 &  x466 &  x538 &  x610 &  x621 &  x652 & ~x9 & ~x27 & ~x118 & ~x174;
assign c2249 = ~x17 & ~x45;
assign c2251 =  x92 &  x152 &  x156 &  x209 &  x264 &  x329 &  x408 &  x427 &  x513 &  x551 &  x607 &  x636 &  x652 &  x679 &  x684 &  x738 &  x747 & ~x143 & ~x561 & ~x672 & ~x733 & ~x761;
assign c2253 = ~x733;
assign c2255 =  x376 &  x387 &  x457 &  x466 &  x523 &  x552 &  x624 &  x626 &  x761 & ~x739;
assign c2257 =  x32;
assign c2259 =  x448;
assign c2261 =  x17 &  x738;
assign c2263 =  x137;
assign c2265 = ~x45;
assign c2267 =  x81;
assign c2269 =  x39 & ~x498 & ~x527 & ~x566 & ~x611 & ~x704;
assign c2271 =  x65 &  x154 &  x259 &  x299 &  x372 &  x466 &  x467 &  x652 &  x691 &  x707 &  x720 &  x769;
assign c2273 =  x39 &  x213 &  x239 &  x245 &  x429 &  x466 &  x551 &  x683 & ~x313;
assign c2275 =  x40 &  x130 &  x154 &  x210 &  x214 &  x236 &  x237 &  x407 &  x408 &  x457 &  x466 &  x467 &  x512 &  x603 &  x655 &  x680 & ~x31 & ~x59 & ~x341 & ~x367 & ~x422 & ~x560 & ~x648 & ~x699;
assign c2277 =  x448;
assign c2279 =  x186 &  x209 &  x210 &  x214 &  x238 &  x321 &  x352 &  x413 &  x427 &  x438 &  x457 &  x466 &  x545 &  x549 &  x551 &  x570 &  x578 &  x711 &  x738 &  x741 & ~x18 & ~x27 & ~x55 & ~x168 & ~x195 & ~x732;
assign c2281 = ~x39 & ~x45 & ~x121;
assign c2283 =  x7;
assign c2285 =  x475;
assign c2287 =  x94 &  x99 &  x146 &  x154 &  x184 &  x208 &  x236 &  x237 &  x265 &  x288 &  x326 &  x353 &  x354 &  x376 &  x406 &  x414 &  x425 &  x431 &  x485 &  x498 &  x519 &  x525 &  x537 &  x566 &  x597 &  x620 &  x650 & ~x17 & ~x26 & ~x35 & ~x36 & ~x46 & ~x47 & ~x109 & ~x138 & ~x163 & ~x170 & ~x306 & ~x334 & ~x393 & ~x394 & ~x419 & ~x450 & ~x506 & ~x561 & ~x646 & ~x783;
assign c2289 =  x192;
assign c2291 =  x57;
assign c2293 =  x114;
assign c2295 =  x14 &  x72 &  x95 &  x181 &  x265 &  x289 &  x300 &  x346 &  x348 &  x490 &  x523 &  x597 & ~x10 & ~x17 & ~x46 & ~x47 & ~x391;
assign c2297 = ~x518 & ~x685;
assign c2299 = ~x580 & ~x610;
assign c2303 =  x51;
assign c2305 =  x55;
assign c2307 = ~x298;
assign c2309 = ~x385 & ~x607;
assign c2311 =  x361;
assign c2313 = ~x39;
assign c2315 = ~x652 & ~x666;
assign c2317 = ~x469 & ~x470 & ~x554 & ~x649;
assign c2319 = ~x317;
assign c2321 =  x468 &  x510 & ~x17 & ~x46 & ~x47 & ~x211;
assign c2323 =  x280;
assign c2325 = ~x204;
assign c2327 = ~x46 & ~x289;
assign c2329 =  x162 &  x324 &  x521 &  x572 &  x612 &  x624 & ~x17 & ~x736;
assign c2331 =  x466 & ~x42;
assign c2333 =  x93 &  x176 &  x205 &  x212 &  x216 &  x238 &  x291 &  x293 &  x315 &  x326 &  x327 &  x350 &  x355 &  x356 &  x378 &  x425 &  x426 &  x455 &  x457 &  x458 &  x463 &  x466 &  x510 &  x525 &  x547 &  x554 &  x575 &  x598 &  x600 &  x603 &  x604 &  x610 &  x626 &  x637 & ~x17 & ~x36 & ~x46 & ~x47 & ~x59 & ~x80 & ~x89 & ~x113 & ~x194 & ~x226 & ~x254 & ~x279 & ~x310 & ~x419 & ~x447 & ~x532 & ~x587 & ~x588 & ~x699 & ~x702 & ~x726 & ~x774 & ~x775;
assign c2335 = ~x342;
assign c2337 =  x363;
assign c2339 = ~x175;
assign c2341 =  x10 & ~x553;
assign c2343 =  x194;
assign c2345 =  x23;
assign c2347 = ~x198 & ~x454 & ~x498 & ~x722;
assign c2349 =  x169;
assign c2351 =  x278;
assign c2353 =  x42 &  x260 &  x347 &  x485 &  x516 &  x570 &  x578 &  x609 & ~x17 & ~x45 & ~x46 & ~x47 & ~x53 & ~x142 & ~x166 & ~x280 & ~x333 & ~x335 & ~x669;
assign c2355 =  x24;
assign c2357 =  x55;
assign c2359 =  x238 &  x266 &  x294 &  x355 &  x440 &  x455 &  x566 &  x598 & ~x36 & ~x37 & ~x45 & ~x46 & ~x775;
assign c2363 =  x169;
assign c2365 =  x48;
assign c2367 =  x12 &  x14 &  x39 &  x208 &  x238 &  x245 &  x269 &  x297 &  x397 &  x401 &  x457 &  x466 &  x468 &  x496 &  x523 &  x552 &  x581 &  x634 & ~x18 & ~x47 & ~x48 & ~x51 & ~x335 & ~x502 & ~x645 & ~x758;
assign c2369 =  x47 & ~x593 & ~x610;
assign c2371 = ~x599;
assign c2373 =  x363;
assign c2375 =  x13 &  x67 &  x93 &  x120 &  x159 &  x175 &  x213 &  x233 &  x235 &  x238 &  x287 &  x292 &  x301 &  x318 &  x320 &  x325 &  x345 &  x353 &  x379 &  x426 &  x454 &  x455 &  x457 &  x466 &  x497 &  x498 &  x515 &  x520 &  x523 &  x541 &  x574 &  x578 &  x582 &  x601 &  x626 &  x660 & ~x9 & ~x17 & ~x20 & ~x21 & ~x36 & ~x47 & ~x59 & ~x63 & ~x77 & ~x81 & ~x107 & ~x117 & ~x164 & ~x194 & ~x196 & ~x252 & ~x254 & ~x276 & ~x305 & ~x307 & ~x363 & ~x616 & ~x643 & ~x644 & ~x700;
assign c2377 = ~x343;
assign c2379 =  x363;
assign c2381 =  x36 & ~x470;
assign c2383 = ~x121 & ~x180;
assign c2385 = ~x120 & ~x317;
assign c2387 =  x127 &  x154 &  x205 &  x207 &  x211 &  x240 &  x272 &  x287 &  x342 &  x382 &  x402 &  x462 &  x492 &  x513 &  x521 &  x523 &  x546 &  x548 &  x549 &  x572 &  x576 &  x624 &  x638 &  x652 &  x667 &  x694 & ~x5 & ~x11 & ~x18 & ~x139 & ~x277 & ~x534 & ~x586 & ~x589 & ~x614 & ~x756 & ~x767;
assign c2389 = ~x202 & ~x721;
assign c2391 = ~x147;
assign c2395 =  x249;
assign c2397 = ~x45 & ~x263 & ~x711 & ~x749;
assign c2399 = ~x175 & ~x204;
assign c2401 =  x169;
assign c2403 =  x179 & ~x453 & ~x498 & ~x538;
assign c2405 = ~x17 & ~x204;
assign c2407 =  x249;
assign c2409 =  x180 &  x212 &  x235 &  x242 &  x376 &  x377 &  x523 &  x596 &  x609 &  x761 & ~x24 & ~x36 & ~x613 & ~x745;
assign c2411 = ~x17 & ~x36 & ~x46 & ~x47 & ~x76 & ~x211;
assign c2413 =  x587;
assign c2415 =  x102 &  x206 &  x291 &  x324 &  x325 &  x328 &  x354 &  x384 &  x408 &  x437 &  x459 &  x468 &  x550 &  x551 &  x552 &  x636 &  x679 &  x682 &  x692 &  x720 & ~x26 & ~x28 & ~x169 & ~x226 & ~x253 & ~x310 & ~x390 & ~x445 & ~x446 & ~x561 & ~x618 & ~x778;
assign c2417 =  x151 &  x156 &  x158 &  x179 &  x186 &  x213 &  x241 &  x267 &  x269 &  x294 &  x315 &  x316 &  x344 &  x385 &  x429 &  x441 &  x456 &  x481 &  x485 &  x495 &  x498 &  x543 &  x552 &  x578 &  x580 &  x595 &  x627 &  x629 &  x651 &  x652 &  x655 &  x661 &  x662 &  x667 & ~x167 & ~x221 & ~x308 & ~x447 & ~x770 & ~x774 & ~x775;
assign c2419 =  x71 &  x188 &  x289 &  x322 &  x329 &  x374 &  x439 &  x465 &  x483 &  x522 &  x523 &  x570 &  x580 &  x626 &  x635 &  x714 &  x717 & ~x4 & ~x390 & ~x419 & ~x446 & ~x618 & ~x670 & ~x695 & ~x731 & ~x732 & ~x778;
assign c2421 = ~x17 & ~x37 & ~x47 & ~x96;
assign c2423 = ~x637 & ~x664;
assign c2425 =  x362;
assign c2427 =  x84;
assign c2429 =  x211 &  x238 &  x239 &  x244 &  x265 &  x289 &  x317 &  x405 &  x426 &  x429 &  x455 &  x457 &  x466 &  x483 &  x496 &  x525 &  x539 &  x552 &  x568 &  x574 &  x580 &  x595 &  x609 &  x624 &  x636 &  x650 &  x692 & ~x22 & ~x31 & ~x86 & ~x140 & ~x141 & ~x275 & ~x281 & ~x308 & ~x333 & ~x337 & ~x364 & ~x447 & ~x504 & ~x505 & ~x534 & ~x557 & ~x591 & ~x617 & ~x672 & ~x697 & ~x757;
assign c2431 = ~x45 & ~x46 & ~x47 & ~x184;
assign c2433 =  x141;
assign c2435 =  x7;
assign c2437 =  x59;
assign c2439 =  x57;
assign c2441 = ~x36 & ~x184;
assign c2443 =  x26;
assign c2445 = ~x569 & ~x580;
assign c2447 = ~x554 & ~x636;
assign c2449 =  x128 &  x205 &  x210 &  x242 &  x319 &  x320 &  x326 &  x400 &  x403 &  x441 &  x456 &  x457 &  x468 &  x481 &  x483 &  x490 &  x497 &  x517 &  x525 &  x537 &  x542 &  x580 &  x593 &  x625 &  x638 &  x662 & ~x24 & ~x27 & ~x29 & ~x51 & ~x110 & ~x112 & ~x118 & ~x194 & ~x222 & ~x338 & ~x451 & ~x535 & ~x731 & ~x755;
assign c2451 =  x71 &  x152 &  x157 &  x180 &  x205 &  x209 &  x323 &  x379 &  x399 &  x439 &  x469 &  x482 &  x483 &  x524 &  x537 &  x571 &  x580 &  x594 &  x597 &  x607 &  x609 &  x611 &  x630 &  x652 &  x653 &  x676 &  x678 &  x732 &  x761 & ~x21 & ~x142 & ~x171 & ~x504 & ~x586 & ~x587 & ~x614;
assign c2453 =  x644;
assign c2455 = ~x412 & ~x413 & ~x470;
assign c2457 =  x448;
assign c2459 = ~x38 & ~x45 & ~x263;
assign c2461 = ~x208;
assign c2463 = ~x11 & ~x17 & ~x47 & ~x96 & ~x158;
assign c2465 =  x447;
assign c2467 =  x588;
assign c2469 = ~x189;
assign c2471 =  x59;
assign c2473 =  x782;
assign c2475 = ~x39 & ~x204;
assign c2477 =  x50;
assign c2479 =  x559;
assign c2481 =  x7;
assign c2483 =  x42 &  x316 &  x344 & ~x0 & ~x18 & ~x21 & ~x36 & ~x37 & ~x45 & ~x46 & ~x47 & ~x76 & ~x77 & ~x80 & ~x107 & ~x112 & ~x220 & ~x306 & ~x334 & ~x391 & ~x417 & ~x418 & ~x422 & ~x447 & ~x474 & ~x698 & ~x702 & ~x736 & ~x748 & ~x753;
assign c2485 = ~x69 & ~x121;
assign c2487 =  x27;
assign c2489 =  x756;
assign c2493 =  x334;
assign c2495 =  x1;
assign c2497 =  x71 &  x176 &  x178 &  x179 &  x181 &  x210 &  x212 &  x240 &  x267 &  x272 &  x288 &  x324 &  x341 &  x353 &  x358 &  x380 &  x402 &  x441 &  x466 &  x468 &  x488 &  x496 &  x515 &  x548 &  x554 &  x555 &  x569 &  x571 &  x579 &  x621 &  x622 &  x658 & ~x0 & ~x4 & ~x8 & ~x27 & ~x32 & ~x47 & ~x49 & ~x108 & ~x141 & ~x226 & ~x251 & ~x253 & ~x307 & ~x334 & ~x361 & ~x393 & ~x449 & ~x473 & ~x561 & ~x764;
assign c2499 = ~x17 & ~x45 & ~x47 & ~x152;
assign c30 =  x37 &  x132 &  x148 &  x245 &  x546 & ~x0 & ~x62 & ~x90 & ~x113 & ~x449 & ~x506 & ~x642 & ~x649 & ~x779;
assign c32 =  x74 &  x132 &  x329 & ~x191 & ~x217 & ~x219 & ~x255 & ~x313 & ~x396 & ~x612 & ~x678 & ~x735;
assign c34 =  x102 &  x741 &  x750;
assign c36 =  x439 & ~x204 & ~x272 & ~x334 & ~x558 & ~x560 & ~x700;
assign c38 =  x429 & ~x107 & ~x275 & ~x493 & ~x503 & ~x534;
assign c310 =  x271 & ~x6 & ~x28 & ~x52 & ~x60 & ~x85 & ~x112 & ~x114 & ~x117 & ~x136 & ~x191 & ~x200 & ~x228 & ~x306 & ~x326 & ~x416 & ~x472 & ~x618 & ~x636 & ~x648 & ~x667 & ~x669 & ~x678 & ~x679 & ~x693 & ~x704 & ~x705 & ~x751 & ~x760 & ~x761 & ~x764 & ~x776 & ~x777;
assign c312 = ~x231 & ~x329 & ~x381 & ~x522 & ~x550;
assign c314 =  x37 &  x371 &  x455 &  x499;
assign c316 = ~x128 & ~x499 & ~x735 & ~x750;
assign c318 =  x37 &  x76 &  x537 &  x738 & ~x391 & ~x395 & ~x562;
assign c320 =  x677;
assign c322 = ~x67 & ~x81 & ~x227 & ~x282 & ~x332 & ~x334 & ~x361 & ~x388 & ~x417 & ~x471 & ~x506 & ~x584 & ~x596 & ~x652 & ~x669 & ~x698 & ~x750;
assign c324 =  x37 &  x47 &  x174 &  x217 &  x684 & ~x4 & ~x29 & ~x200 & ~x222 & ~x251 & ~x280 & ~x367 & ~x390 & ~x447 & ~x533 & ~x558 & ~x617;
assign c326 =  x15 &  x44 &  x47 &  x148 &  x517 & ~x29 & ~x54 & ~x113 & ~x165 & ~x249 & ~x254 & ~x394;
assign c328 =  x66 &  x125 &  x148 &  x178 &  x267 &  x434 &  x490 &  x713 & ~x5 & ~x52 & ~x62 & ~x77 & ~x90 & ~x220 & ~x339 & ~x420 & ~x446 & ~x527 & ~x566 & ~x590 & ~x609 & ~x642 & ~x679 & ~x733;
assign c330 =  x99 &  x124 &  x129 &  x151 &  x154 &  x182 &  x212 &  x267 &  x293 &  x350 &  x408 &  x522 &  x574 &  x577 &  x690 & ~x9 & ~x22 & ~x23 & ~x25 & ~x28 & ~x57 & ~x61 & ~x81 & ~x111 & ~x140 & ~x192 & ~x226 & ~x258 & ~x281 & ~x315 & ~x339 & ~x394 & ~x453 & ~x614 & ~x643 & ~x669;
assign c332 = ~x242 & ~x342 & ~x771;
assign c334 =  x348 & ~x195 & ~x345;
assign c336 =  x422;
assign c338 =  x319 & ~x1 & ~x29 & ~x78 & ~x80 & ~x106 & ~x228 & ~x381 & ~x472 & ~x531 & ~x580 & ~x724 & ~x757;
assign c340 = ~x273 & ~x333 & ~x548;
assign c342 = ~x285 & ~x471 & ~x604;
assign c344 =  x132 &  x148 & ~x0 & ~x19 & ~x20 & ~x59 & ~x79 & ~x91 & ~x107 & ~x247 & ~x255 & ~x282 & ~x474 & ~x506 & ~x679 & ~x751;
assign c346 =  x36 &  x37 &  x47 &  x64 &  x91 &  x119 &  x738 & ~x250 & ~x303 & ~x311;
assign c348 = ~x8 & ~x23 & ~x24 & ~x69 & ~x90 & ~x143 & ~x336 & ~x476 & ~x619 & ~x700 & ~x708;
assign c350 =  x6;
assign c352 =  x366;
assign c354 = ~x79 & ~x199 & ~x234 & ~x248 & ~x326 & ~x389 & ~x473 & ~x558 & ~x774;
assign c356 =  x630 & ~x1 & ~x34 & ~x89 & ~x115 & ~x139 & ~x141 & ~x169 & ~x247 & ~x274 & ~x275 & ~x282 & ~x285 & ~x337 & ~x340 & ~x447 & ~x452 & ~x512 & ~x531 & ~x552 & ~x554 & ~x567 & ~x580 & ~x581 & ~x608 & ~x615 & ~x647 & ~x651 & ~x667 & ~x669 & ~x671 & ~x679 & ~x704 & ~x753;
assign c358 = ~x436;
assign c360 = ~x24 & ~x133 & ~x231 & ~x253 & ~x282 & ~x296 & ~x593;
assign c362 =  x63 &  x509;
assign c364 =  x690 & ~x270;
assign c366 =  x37 &  x91 &  x234 & ~x23 & ~x59 & ~x194 & ~x248 & ~x282 & ~x334 & ~x336 & ~x367 & ~x475 & ~x500 & ~x674 & ~x779;
assign c368 =  x65 &  x189 &  x735 &  x739 &  x741 &  x743 &  x748 & ~x250 & ~x255 & ~x448 & ~x619 & ~x760;
assign c370 =  x38 &  x722 &  x741;
assign c372 = ~x25 & ~x31 & ~x43 & ~x61 & ~x62 & ~x63 & ~x77 & ~x78 & ~x107 & ~x137 & ~x196 & ~x308 & ~x335 & ~x618 & ~x641 & ~x701;
assign c374 =  x38 &  x74 &  x75 &  x91 &  x119 &  x210 &  x370 & ~x192 & ~x728 & ~x730;
assign c376 = ~x128 & ~x709;
assign c378 =  x263 &  x624 &  x625 & ~x217 & ~x220 & ~x232 & ~x336 & ~x472 & ~x701 & ~x754;
assign c380 =  x405 &  x658 & ~x9 & ~x200 & ~x401 & ~x705;
assign c382 =  x123 &  x151 &  x236 &  x264 &  x267 &  x373 &  x433 &  x456 &  x521 &  x543 &  x575 &  x659 &  x680 &  x739 & ~x3 & ~x57 & ~x114 & ~x249 & ~x259 & ~x308 & ~x358 & ~x393 & ~x612 & ~x671;
assign c384 =  x65 &  x287 &  x686 & ~x104 & ~x679;
assign c386 = ~x66 & ~x466;
assign c388 = ~x0 & ~x8 & ~x29 & ~x32 & ~x80 & ~x141 & ~x203 & ~x225 & ~x247 & ~x259 & ~x306 & ~x310 & ~x313 & ~x336 & ~x359 & ~x361 & ~x363 & ~x388 & ~x396 & ~x416 & ~x424 & ~x445 & ~x447 & ~x474 & ~x475 & ~x476 & ~x477 & ~x557 & ~x588 & ~x616 & ~x709 & ~x721 & ~x728 & ~x732 & ~x750 & ~x751 & ~x754 & ~x757;
assign c390 = ~x354;
assign c392 =  x65 &  x91 &  x119 &  x133 &  x154 &  x511 &  x512 &  x635 & ~x534 & ~x779;
assign c394 = ~x134 & ~x259 & ~x273 & ~x329 & ~x357 & ~x438 & ~x449 & ~x453 & ~x482 & ~x509;
assign c396 =  x371 & ~x8 & ~x15 & ~x119 & ~x248 & ~x275 & ~x477 & ~x735;
assign c398 =  x75 & ~x62 & ~x146 & ~x387 & ~x581 & ~x596 & ~x650 & ~x651 & ~x693 & ~x782;
assign c3100 =  x37 &  x46 &  x91 &  x456 &  x457 &  x513 &  x546 &  x604 &  x663 &  x737 & ~x139 & ~x220 & ~x224 & ~x281 & ~x361 & ~x389 & ~x444 & ~x531 & ~x672 & ~x673;
assign c3102 =  x339;
assign c3104 =  x450;
assign c3106 =  x64 &  x92 &  x133 &  x161 &  x688 &  x709 &  x744 &  x748 & ~x3 & ~x220 & ~x589 & ~x778;
assign c3108 = ~x296 & ~x301 & ~x423 & ~x623;
assign c3110 = ~x241 & ~x274 & ~x330 & ~x453 & ~x552 & ~x731 & ~x776 & ~x779;
assign c3112 = ~x27 & ~x78 & ~x90 & ~x113 & ~x163 & ~x170 & ~x173 & ~x196 & ~x465 & ~x476;
assign c3114 =  x37 &  x412 &  x537 & ~x138;
assign c3116 =  x37 &  x122 &  x405 & ~x5 & ~x29 & ~x62 & ~x143 & ~x247 & ~x388 & ~x590 & ~x608 & ~x675 & ~x760 & ~x782;
assign c3118 =  x153 &  x322 & ~x93 & ~x134 & ~x172 & ~x259 & ~x538;
assign c3120 =  x37 &  x553 &  x737 &  x748 & ~x89 & ~x110 & ~x140 & ~x165 & ~x227 & ~x338 & ~x754 & ~x761;
assign c3122 =  x607 & ~x86 & ~x165 & ~x197 & ~x204 & ~x216 & ~x231 & ~x246 & ~x287 & ~x358 & ~x398 & ~x643;
assign c3124 =  x75 &  x412 &  x509;
assign c3126 = ~x173 & ~x552 & ~x777;
assign c3128 = ~x70 & ~x78 & ~x219 & ~x251 & ~x470 & ~x499 & ~x612 & ~x723 & ~x775;
assign c3130 =  x41 &  x545 &  x573 &  x602 &  x710 & ~x0 & ~x10 & ~x23 & ~x56 & ~x104 & ~x107 & ~x134 & ~x162 & ~x171 & ~x172 & ~x189 & ~x200 & ~x224 & ~x225 & ~x228 & ~x230 & ~x255 & ~x278 & ~x282 & ~x286 & ~x336 & ~x367 & ~x390 & ~x393 & ~x426 & ~x532 & ~x584 & ~x591 & ~x701 & ~x731 & ~x735 & ~x754;
assign c3132 = ~x73 & ~x134 & ~x373 & ~x693;
assign c3134 =  x101 &  x181 &  x240 &  x325 &  x327 &  x351 &  x408 &  x518 &  x546 &  x628 &  x629 &  x659 &  x686 &  x743 & ~x1 & ~x2 & ~x6 & ~x8 & ~x29 & ~x35 & ~x61 & ~x62 & ~x81 & ~x161 & ~x195 & ~x197 & ~x248 & ~x275 & ~x306 & ~x340 & ~x396 & ~x415 & ~x416 & ~x454 & ~x478 & ~x482 & ~x510 & ~x588 & ~x589 & ~x590 & ~x613 & ~x646 & ~x671 & ~x701 & ~x706 & ~x730 & ~x749 & ~x776 & ~x779;
assign c3136 =  x123 &  x125 &  x129 &  x154 &  x182 &  x213 &  x291 &  x298 &  x354 &  x377 &  x383 &  x409 &  x410 &  x513 &  x517 &  x568 &  x575 &  x577 &  x578 &  x596 &  x659 &  x662 &  x690 &  x692 &  x746 & ~x26 & ~x30 & ~x57 & ~x58 & ~x87 & ~x110 & ~x114 & ~x137 & ~x170 & ~x220 & ~x309 & ~x333 & ~x391 & ~x443 & ~x446 & ~x475 & ~x499 & ~x503 & ~x529 & ~x558 & ~x587 & ~x613 & ~x614 & ~x726 & ~x728 & ~x760 & ~x783;
assign c3138 =  x271 & ~x55 & ~x283 & ~x326 & ~x330 & ~x639 & ~x704 & ~x722 & ~x751 & ~x781;
assign c3140 =  x74 &  x91 &  x119 &  x243 &  x384 &  x398 &  x491 &  x683 & ~x81 & ~x169 & ~x250 & ~x534 & ~x560 & ~x590 & ~x670 & ~x730 & ~x781;
assign c3142 = ~x652;
assign c3144 = ~x5 & ~x35 & ~x39 & ~x44 & ~x61 & ~x62 & ~x76 & ~x104 & ~x133 & ~x140 & ~x188 & ~x309 & ~x337 & ~x361 & ~x506;
assign c3146 = ~x239 & ~x414;
assign c3148 = ~x156 & ~x595 & ~x764;
assign c3150 =  x132 & ~x327;
assign c3152 =  x188 & ~x345;
assign c3154 =  x769 & ~x10 & ~x62 & ~x82 & ~x85 & ~x133 & ~x203 & ~x579 & ~x779;
assign c3156 =  x151 & ~x200 & ~x469;
assign c3158 = ~x190 & ~x222 & ~x247 & ~x415 & ~x454 & ~x487;
assign c3160 =  x322 &  x377 &  x513 &  x541 & ~x1 & ~x61 & ~x83 & ~x327 & ~x554 & ~x639 & ~x674 & ~x702 & ~x755;
assign c3162 =  x396;
assign c3164 =  x101 &  x290 &  x439 & ~x25 & ~x176 & ~x307 & ~x336;
assign c3166 =  x132 &  x160 & ~x134 & ~x372 & ~x400 & ~x583;
assign c3168 =  x148 & ~x317;
assign c3170 = ~x67 & ~x69 & ~x72 & ~x223 & ~x531 & ~x703;
assign c3172 =  x634 & ~x28 & ~x29 & ~x53 & ~x134 & ~x138 & ~x145 & ~x170 & ~x196 & ~x199 & ~x200 & ~x251 & ~x274 & ~x281 & ~x289 & ~x336 & ~x444 & ~x554 & ~x611 & ~x667 & ~x725 & ~x776;
assign c3174 = ~x463;
assign c3176 =  x129 &  x241 &  x243 &  x545 &  x742 & ~x5 & ~x62 & ~x78 & ~x113 & ~x138 & ~x140 & ~x142 & ~x161 & ~x162 & ~x449 & ~x534 & ~x623 & ~x776;
assign c3178 =  x545 & ~x29 & ~x78 & ~x114 & ~x134 & ~x225 & ~x275 & ~x281 & ~x304 & ~x426 & ~x472 & ~x476 & ~x499 & ~x532 & ~x596 & ~x652 & ~x679 & ~x707 & ~x754;
assign c3180 =  x65 &  x344 &  x384 &  x385 & ~x53 & ~x275 & ~x622 & ~x668;
assign c3182 =  x38 &  x65 &  x94 &  x385 &  x398 &  x456 &  x468 &  x484 &  x566 &  x630 & ~x587;
assign c3184 =  x6;
assign c3186 = ~x203 & ~x231 & ~x426 & ~x548 & ~x589;
assign c3188 =  x129 &  x157 &  x208 &  x236 &  x267 &  x373 &  x734 &  x735 & ~x53 & ~x54 & ~x59 & ~x85 & ~x111 & ~x166 & ~x284 & ~x392 & ~x448 & ~x562 & ~x589 & ~x643 & ~x760;
assign c3190 =  x181 &  x371 & ~x203;
assign c3192 =  x456 &  x499;
assign c3194 =  x208 &  x296 &  x680 & ~x301 & ~x509 & ~x651;
assign c3196 =  x133 & ~x58 & ~x220 & ~x287 & ~x300 & ~x343 & ~x531 & ~x587 & ~x731;
assign c3198 =  x157 &  x435 &  x455 &  x659 &  x766 & ~x0 & ~x451 & ~x611 & ~x679;
assign c3200 = ~x390 & ~x407;
assign c3202 =  x63 &  x65 &  x370;
assign c3204 =  x124 &  x242 &  x377 &  x428 &  x518 &  x635 &  x657 & ~x59 & ~x114 & ~x315 & ~x359 & ~x667;
assign c3206 = ~x7 & ~x23 & ~x112 & ~x163 & ~x190 & ~x191 & ~x203 & ~x258 & ~x286 & ~x301 & ~x313 & ~x317 & ~x343 & ~x356 & ~x358 & ~x359 & ~x428 & ~x447 & ~x484 & ~x501 & ~x538 & ~x641 & ~x651 & ~x668 & ~x678;
assign c3208 =  x101 &  x160 &  x189 &  x739 &  x747 & ~x62 & ~x107 & ~x669;
assign c3210 =  x36 &  x37 &  x91 &  x486 &  x597 &  x744 & ~x3 & ~x32 & ~x113 & ~x170 & ~x219 & ~x220 & ~x248 & ~x310 & ~x331 & ~x359 & ~x393 & ~x449 & ~x476 & ~x478 & ~x503 & ~x530 & ~x647 & ~x730 & ~x758 & ~x762 & ~x779;
assign c3212 = ~x73 & ~x249;
assign c3214 =  x127 &  x487 &  x692 &  x719 &  x741 &  x748 &  x749 & ~x20 & ~x35 & ~x52 & ~x56 & ~x107 & ~x251 & ~x308 & ~x476 & ~x589 & ~x644 & ~x758;
assign c3216 =  x215 & ~x11 & ~x382 & ~x454;
assign c3218 =  x37 &  x370 &  x439 &  x626 & ~x562;
assign c3220 =  x379 &  x490 &  x577 & ~x29 & ~x52 & ~x173 & ~x309 & ~x362 & ~x427 & ~x568 & ~x672 & ~x676 & ~x750 & ~x755;
assign c3222 = ~x436 & ~x453;
assign c3224 =  x38 &  x748 &  x749 & ~x306 & ~x534;
assign c3226 =  x748 &  x749 &  x750;
assign c3228 =  x311;
assign c3230 =  x290 &  x292 &  x541 &  x636 &  x710 &  x739 &  x748 &  x749 &  x769 & ~x757;
assign c3232 =  x64 &  x124 &  x125 &  x184 &  x294 &  x433 &  x546 &  x573 &  x741 &  x743 & ~x22 & ~x62 & ~x134 & ~x219 & ~x282 & ~x309 & ~x310 & ~x336 & ~x476 & ~x479 & ~x563 & ~x703 & ~x781;
assign c3234 = ~x86 & ~x289 & ~x298;
assign c3236 = ~x103 & ~x365 & ~x432;
assign c3238 =  x659 &  x745 & ~x3 & ~x86 & ~x169 & ~x256 & ~x333 & ~x709;
assign c3240 = ~x1 & ~x6 & ~x8 & ~x70 & ~x88 & ~x141 & ~x142 & ~x170 & ~x201 & ~x218 & ~x222 & ~x275 & ~x277 & ~x278 & ~x282 & ~x333 & ~x368 & ~x449 & ~x450 & ~x451 & ~x471 & ~x475 & ~x499 & ~x559 & ~x612 & ~x618 & ~x641 & ~x642 & ~x665 & ~x725 & ~x730 & ~x732 & ~x749 & ~x754 & ~x760 & ~x779;
assign c3242 =  x101 &  x125 &  x210 &  x271 &  x405 &  x517 &  x545 &  x548 &  x600 & ~x1 & ~x113 & ~x133 & ~x202 & ~x229 & ~x310 & ~x362 & ~x393 & ~x478 & ~x580 & ~x594 & ~x610 & ~x612 & ~x618 & ~x665 & ~x782;
assign c3244 =  x65 &  x148 &  x315 & ~x524;
assign c3246 =  x41 & ~x258 & ~x297 & ~x314 & ~x330 & ~x467 & ~x580 & ~x641 & ~x748;
assign c3248 =  x105 &  x735 & ~x85 & ~x590;
assign c3250 =  x328 &  x738 & ~x161 & ~x249 & ~x534 & ~x567 & ~x609;
assign c3252 =  x517 &  x545 &  x573 & ~x230 & ~x273 & ~x312 & ~x495 & ~x510 & ~x757;
assign c3254 =  x105 &  x122 &  x468 &  x511 & ~x3 & ~x54 & ~x86 & ~x220;
assign c3256 =  x37 &  x749 &  x750;
assign c3258 = ~x200 & ~x407;
assign c3260 = ~x241 & ~x301 & ~x382 & ~x466;
assign c3262 = ~x133 & ~x231 & ~x232 & ~x259 & ~x270 & ~x299 & ~x355 & ~x454;
assign c3264 = ~x134 & ~x270;
assign c3266 =  x573 & ~x93 & ~x133 & ~x230 & ~x274 & ~x313 & ~x569 & ~x678 & ~x751;
assign c3268 =  x417;
assign c3270 =  x64 &  x384 &  x398 &  x537;
assign c3272 =  x124 &  x125 &  x126 &  x236 &  x349 &  x354 &  x377 &  x383 &  x434 &  x462 &  x571 &  x575 &  x598 &  x625 &  x654 & ~x0 & ~x27 & ~x30 & ~x55 & ~x231 & ~x311;
assign c3274 =  x216 &  x634 & ~x248 & ~x763;
assign c3276 =  x64 &  x189 &  x217 & ~x90 & ~x224;
assign c3278 =  x71 &  x292 &  x433 &  x491 &  x545 &  x742 & ~x31 & ~x52 & ~x53 & ~x113 & ~x249 & ~x287 & ~x303 & ~x389 & ~x423 & ~x471 & ~x756 & ~x782;
assign c3280 =  x65 &  x97 &  x766 & ~x9 & ~x22 & ~x48 & ~x85 & ~x679;
assign c3282 =  x21;
assign c3284 =  x43 & ~x655;
assign c3286 = ~x68;
assign c3288 =  x461 &  x513 &  x597 &  x690 & ~x5 & ~x27 & ~x54 & ~x88 & ~x114 & ~x327 & ~x562 & ~x564 & ~x723;
assign c3290 =  x240 & ~x0 & ~x1 & ~x14 & ~x16 & ~x23 & ~x29 & ~x30 & ~x34 & ~x43 & ~x58 & ~x108 & ~x170 & ~x195 & ~x222 & ~x282 & ~x393 & ~x475 & ~x669 & ~x706 & ~x724;
assign c3292 = ~x29 & ~x436 & ~x454;
assign c3294 = ~x29 & ~x100 & ~x110 & ~x165 & ~x392 & ~x497 & ~x728 & ~x764;
assign c3296 = ~x219 & ~x463;
assign c3298 =  x65 &  x370 &  x398 & ~x251 & ~x334 & ~x621;
assign c3300 =  x294 &  x513 & ~x58 & ~x299 & ~x762;
assign c3302 = ~x259 & ~x261 & ~x271 & ~x300 & ~x427 & ~x454 & ~x725;
assign c3304 =  x322 &  x430 & ~x135 & ~x277 & ~x317 & ~x446 & ~x534;
assign c3306 =  x11 &  x45 &  x66 &  x132 &  x160 &  x241 &  x377 &  x654 &  x663 &  x711 &  x712 &  x717 & ~x27 & ~x54 & ~x112 & ~x135 & ~x140 & ~x165 & ~x169 & ~x191 & ~x251 & ~x283 & ~x336 & ~x389 & ~x393 & ~x475 & ~x476 & ~x532 & ~x533 & ~x586 & ~x590 & ~x641 & ~x750 & ~x781;
assign c3308 =  x377 &  x748 & ~x59 & ~x107 & ~x272 & ~x274 & ~x306 & ~x387 & ~x392 & ~x783;
assign c3310 = ~x68 & ~x298;
assign c3312 = ~x271 & ~x275 & ~x427 & ~x482 & ~x499;
assign c3314 =  x16 &  x36 &  x65 &  x745;
assign c3316 =  x128 &  x153 &  x211 &  x322 &  x373 &  x378 &  x464 &  x546 &  x575 &  x680 &  x692 &  x739 & ~x2 & ~x22 & ~x51 & ~x53 & ~x142 & ~x166 & ~x252 & ~x443 & ~x476 & ~x504 & ~x703;
assign c3318 =  x46 &  x47 &  x64 &  x74 &  x147 &  x513 &  x713 & ~x4 & ~x28 & ~x87 & ~x108 & ~x110 & ~x136 & ~x138 & ~x191 & ~x198 & ~x222 & ~x252 & ~x336 & ~x392 & ~x417 & ~x590 & ~x622 & ~x638 & ~x649 & ~x701 & ~x723 & ~x728 & ~x730 & ~x779;
assign c3320 =  x376 &  x466 & ~x81 & ~x138 & ~x145 & ~x221 & ~x255 & ~x256 & ~x309 & ~x327 & ~x336 & ~x362 & ~x421 & ~x447 & ~x476 & ~x479 & ~x501 & ~x558 & ~x565 & ~x619 & ~x639 & ~x669 & ~x671 & ~x677 & ~x728 & ~x730 & ~x751 & ~x752;
assign c3322 = ~x0 & ~x29 & ~x53 & ~x60 & ~x167 & ~x196 & ~x247 & ~x254 & ~x282 & ~x341 & ~x358 & ~x454 & ~x484 & ~x504 & ~x531 & ~x563 & ~x620 & ~x642 & ~x669 & ~x722 & ~x771 & ~x778 & ~x783;
assign c3324 =  x127 &  x129 &  x148 &  x350 &  x432 &  x465 &  x547 & ~x10 & ~x54 & ~x137 & ~x164 & ~x200 & ~x219 & ~x276 & ~x332 & ~x335 & ~x584 & ~x595 & ~x731;
assign c3326 = ~x85 & ~x96 & ~x377;
assign c3328 = ~x66 & ~x165 & ~x301 & ~x332 & ~x466 & ~x704 & ~x731;
assign c3330 = ~x8 & ~x171 & ~x268 & ~x305 & ~x332 & ~x427 & ~x506 & ~x536 & ~x557 & ~x592 & ~x615 & ~x645 & ~x649 & ~x696;
assign c3332 =  x349 &  x545 &  x633 & ~x221 & ~x271 & ~x356 & ~x730;
assign c3334 =  x36 &  x91 &  x105;
assign c3336 = ~x221 & ~x242 & ~x244 & ~x254 & ~x273 & ~x441 & ~x568 & ~x580 & ~x773;
assign c3338 =  x317 & ~x29 & ~x274 & ~x427 & ~x454 & ~x524;
assign c3340 =  x64 &  x122 &  x370 &  x663 &  x741 & ~x27 & ~x331;
assign c3342 = ~x69 & ~x118 & ~x133 & ~x134 & ~x190 & ~x422 & ~x534 & ~x561 & ~x679 & ~x705;
assign c3344 =  x400 & ~x159 & ~x220 & ~x282;
assign c3346 =  x311 &  x478;
assign c3348 =  x157 &  x741 & ~x113 & ~x138 & ~x250 & ~x274 & ~x418 & ~x496 & ~x589 & ~x721;
assign c3350 = ~x182 & ~x367 & ~x505 & ~x665 & ~x679 & ~x703 & ~x752 & ~x753;
assign c3352 =  x41 &  x45 &  x64 &  x489 & ~x0 & ~x2 & ~x4 & ~x22 & ~x24 & ~x27 & ~x29 & ~x61 & ~x107 & ~x113 & ~x134 & ~x171 & ~x221 & ~x229 & ~x360 & ~x363 & ~x453 & ~x474 & ~x501 & ~x535 & ~x589 & ~x615 & ~x701 & ~x724 & ~x728 & ~x761 & ~x779;
assign c3354 = ~x466 & ~x485 & ~x541 & ~x569;
assign c3356 =  x45 &  x72 &  x74 &  x91 &  x119 &  x147 &  x174 &  x568 & ~x1 & ~x24 & ~x61 & ~x112 & ~x113 & ~x200 & ~x222 & ~x366 & ~x449 & ~x474 & ~x502 & ~x592 & ~x727;
assign c3358 =  x422;
assign c3360 =  x37 &  x677;
assign c3362 =  x95 &  x211 &  x212 &  x463 &  x540 &  x659 &  x682 &  x743 & ~x0 & ~x2 & ~x28 & ~x52 & ~x87 & ~x114 & ~x140 & ~x143 & ~x256 & ~x272 & ~x309 & ~x330 & ~x336 & ~x362 & ~x365 & ~x394 & ~x418 & ~x449 & ~x470 & ~x475 & ~x589 & ~x613 & ~x699 & ~x701 & ~x724 & ~x728;
assign c3364 =  x261 & ~x78 & ~x514 & ~x534;
assign c3366 = ~x170 & ~x203 & ~x229 & ~x485 & ~x523 & ~x679;
assign c3368 =  x124 &  x129 &  x213 &  x405 &  x462 &  x518 &  x570 &  x577 &  x713 & ~x29 & ~x215 & ~x416 & ~x503 & ~x761;
assign c3370 = ~x301 & ~x408 & ~x603;
assign c3372 = ~x73 & ~x569;
assign c3374 =  x121 &  x177 &  x236 &  x322 &  x352 &  x376 &  x378 &  x407 &  x462 &  x491 &  x546 &  x606 &  x628 &  x629 &  x631 &  x713 & ~x20 & ~x25 & ~x27 & ~x58 & ~x82 & ~x107 & ~x114 & ~x116 & ~x144 & ~x162 & ~x170 & ~x221 & ~x226 & ~x230 & ~x283 & ~x387 & ~x390 & ~x449 & ~x497 & ~x502 & ~x503 & ~x582 & ~x637 & ~x665 & ~x666 & ~x674 & ~x725 & ~x733;
assign c3376 =  x433 & ~x297 & ~x470 & ~x693;
assign c3378 =  x746 & ~x4 & ~x12 & ~x24 & ~x28 & ~x30 & ~x59 & ~x143 & ~x221 & ~x277 & ~x327 & ~x424 & ~x472 & ~x476 & ~x583 & ~x588 & ~x639 & ~x695 & ~x762;
assign c3380 =  x374 &  x405 &  x546 &  x577 &  x599 &  x657 &  x658 &  x741 & ~x26 & ~x27 & ~x32 & ~x50 & ~x78 & ~x90 & ~x138 & ~x169 & ~x173 & ~x191 & ~x196 & ~x222 & ~x277 & ~x307 & ~x311 & ~x312 & ~x337 & ~x415 & ~x425 & ~x440 & ~x479 & ~x504 & ~x533 & ~x553 & ~x584 & ~x594 & ~x622 & ~x677 & ~x695 & ~x705 & ~x750 & ~x754 & ~x777;
assign c3382 =  x292 &  x770 & ~x53 & ~x84 & ~x145 & ~x165 & ~x275 & ~x327 & ~x389 & ~x450 & ~x590 & ~x641 & ~x723;
assign c3384 =  x636 & ~x231 & ~x244;
assign c3386 =  x124 &  x129 &  x462 &  x690 &  x742 & ~x90 & ~x105 & ~x171 & ~x217 & ~x230 & ~x274 & ~x330 & ~x332 & ~x471 & ~x473 & ~x533 & ~x590 & ~x609 & ~x679 & ~x701 & ~x735 & ~x778;
assign c3388 =  x294 &  x517 &  x577 & ~x1 & ~x26 & ~x82 & ~x108 & ~x195 & ~x218 & ~x250 & ~x388 & ~x411 & ~x502 & ~x592 & ~x779;
assign c3390 =  x37 &  x65 &  x636 &  x677 &  x735 & ~x195 & ~x281 & ~x306 & ~x391 & ~x534 & ~x782;
assign c3392 =  x127 &  x129 &  x157 &  x545 &  x605 & ~x105 & ~x139 & ~x160 & ~x223 & ~x309 & ~x332 & ~x338 & ~x396 & ~x454 & ~x534 & ~x585 & ~x637 & ~x664 & ~x726;
assign c3394 =  x546 & ~x174 & ~x219 & ~x224 & ~x373 & ~x388 & ~x443 & ~x701;
assign c3396 = ~x93 & ~x411 & ~x467;
assign c3398 = ~x44 & ~x67 & ~x68 & ~x336;
assign c3400 =  x65 &  x70 &  x101 &  x153 &  x379 &  x430 &  x487 &  x489 &  x494 &  x513 &  x545 &  x599 &  x629 &  x685 &  x745 & ~x24 & ~x29 & ~x78 & ~x107 & ~x113 & ~x133 & ~x134 & ~x163 & ~x198 & ~x250 & ~x251 & ~x364 & ~x478 & ~x534 & ~x583 & ~x589 & ~x609 & ~x611 & ~x638 & ~x639 & ~x648 & ~x701;
assign c3402 =  x65 &  x462 &  x766 & ~x76 & ~x105 & ~x425 & ~x589 & ~x651 & ~x679 & ~x748 & ~x779;
assign c3404 = ~x5 & ~x28 & ~x29 & ~x44 & ~x69 & ~x80 & ~x764;
assign c3406 = ~x96 & ~x542;
assign c3408 =  x517 &  x545 &  x630 &  x631 & ~x2 & ~x8 & ~x19 & ~x27 & ~x51 & ~x57 & ~x77 & ~x85 & ~x103 & ~x114 & ~x115 & ~x144 & ~x147 & ~x160 & ~x161 & ~x172 & ~x194 & ~x203 & ~x216 & ~x219 & ~x220 & ~x221 & ~x222 & ~x227 & ~x231 & ~x244 & ~x248 & ~x257 & ~x286 & ~x339 & ~x342 & ~x358 & ~x359 & ~x364 & ~x384 & ~x414 & ~x421 & ~x423 & ~x425 & ~x426 & ~x443 & ~x445 & ~x446 & ~x453 & ~x534 & ~x536 & ~x561 & ~x562 & ~x564 & ~x590 & ~x669 & ~x694 & ~x704 & ~x726 & ~x732 & ~x750 & ~x751 & ~x759 & ~x761;
assign c3410 =  x354 & ~x381 & ~x583;
assign c3412 =  x103 &  x122 &  x371 &  x384 &  x412 &  x464 & ~x48 & ~x107 & ~x217 & ~x219 & ~x534 & ~x611;
assign c3414 = ~x266 & ~x522;
assign c3416 =  x101 &  x213 &  x231 &  x405 &  x408 &  x491 &  x493 &  x598 &  x605 &  x686 &  x710 &  x713 &  x743 & ~x111 & ~x133 & ~x219 & ~x281 & ~x336 & ~x442 & ~x470 & ~x639 & ~x649 & ~x749 & ~x758 & ~x761 & ~x776;
assign c3418 =  x366;
assign c3420 =  x734 & ~x231 & ~x309;
assign c3422 =  x37 &  x119 &  x481;
assign c3424 = ~x234 & ~x289;
assign c3426 =  x245 &  x545 &  x766 & ~x35 & ~x671;
assign c3428 =  x65 &  x132 &  x189 &  x629 & ~x5 & ~x335 & ~x427 & ~x727 & ~x751 & ~x783;
assign c3430 = ~x175 & ~x379;
assign c3432 =  x36 & ~x27 & ~x190 & ~x282 & ~x287 & ~x331 & ~x701;
assign c3434 =  x65 &  x122 &  x177 &  x357 &  x463 &  x542 &  x632 &  x658 &  x741 &  x742 &  x747 & ~x52 & ~x194 & ~x197 & ~x226 & ~x363 & ~x615 & ~x649 & ~x676 & ~x723;
assign c3436 = ~x28 & ~x51 & ~x58 & ~x108 & ~x222 & ~x255 & ~x258 & ~x273 & ~x277 & ~x331 & ~x548 & ~x671 & ~x728;
assign c3438 =  x517 & ~x8 & ~x21 & ~x190 & ~x193 & ~x251 & ~x326 & ~x420 & ~x479 & ~x672;
assign c3440 =  x311;
assign c3442 =  x101 &  x124 &  x127 &  x152 &  x179 &  x320 &  x516 &  x545 &  x546 &  x573 &  x742 & ~x5 & ~x29 & ~x55 & ~x60 & ~x133 & ~x138 & ~x141 & ~x203 & ~x229 & ~x245 & ~x280 & ~x359 & ~x368 & ~x423 & ~x426 & ~x451 & ~x471 & ~x534 & ~x594 & ~x612 & ~x619 & ~x641 & ~x674 & ~x699 & ~x754;
assign c3444 =  x11 &  x65 &  x70 &  x103 &  x237 &  x294 &  x384 &  x487 &  x517 &  x545 &  x738 & ~x2 & ~x24 & ~x29 & ~x222 & ~x473 & ~x534;
assign c3446 = ~x4 & ~x57 & ~x116 & ~x223 & ~x230 & ~x308 & ~x313 & ~x369 & ~x449 & ~x641 & ~x642 & ~x655 & ~x672 & ~x729;
assign c3448 =  x324 &  x457 &  x748 &  x749 &  x766 & ~x25 & ~x170 & ~x196 & ~x591 & ~x673;
assign c3450 =  x132 & ~x2 & ~x29 & ~x49 & ~x106 & ~x111 & ~x112 & ~x114 & ~x139 & ~x163 & ~x198 & ~x225 & ~x275 & ~x336 & ~x364 & ~x367 & ~x419 & ~x421 & ~x447 & ~x472 & ~x483 & ~x503 & ~x590 & ~x622 & ~x693 & ~x706 & ~x730 & ~x759 & ~x779;
assign c3452 = ~x88 & ~x497 & ~x513;
assign c3454 =  x356 &  x385 & ~x13 & ~x30 & ~x80 & ~x138 & ~x306 & ~x366 & ~x642 & ~x678 & ~x729;
assign c3456 = ~x104 & ~x134 & ~x289 & ~x356 & ~x372 & ~x539 & ~x552;
assign c3458 = ~x231 & ~x271 & ~x289 & ~x327 & ~x367 & ~x701;
assign c3460 = ~x484 & ~x572;
assign c3462 = ~x134 & ~x192 & ~x332 & ~x380 & ~x388 & ~x448 & ~x498 & ~x665 & ~x705;
assign c3464 = ~x73 & ~x266 & ~x453;
assign c3466 =  x315 & ~x345;
assign c3468 =  x159 & ~x33 & ~x60 & ~x83 & ~x145 & ~x173 & ~x192 & ~x220 & ~x298 & ~x333 & ~x508 & ~x612 & ~x615 & ~x618 & ~x707 & ~x734 & ~x764 & ~x778 & ~x782;
assign c3470 =  x65 &  x66 &  x122 &  x155 &  x315 &  x384 &  x404 &  x681 &  x713 &  x738 & ~x22 & ~x87 & ~x144 & ~x559 & ~x611 & ~x647 & ~x694;
assign c3472 =  x65 &  x385 & ~x89 & ~x112 & ~x397 & ~x594 & ~x610;
assign c3474 =  x36 &  x565;
assign c3476 =  x332;
assign c3478 =  x375 &  x546 &  x686 &  x747 & ~x61 & ~x78 & ~x367 & ~x454 & ~x484 & ~x679 & ~x703 & ~x756;
assign c3480 =  x275 &  x366;
assign c3482 = ~x356 & ~x464 & ~x776;
assign c3484 = ~x29 & ~x103 & ~x121 & ~x231 & ~x272 & ~x274 & ~x299 & ~x300 & ~x427 & ~x483 & ~x509 & ~x531;
assign c3486 = ~x18 & ~x28 & ~x43 & ~x62 & ~x78 & ~x107 & ~x196 & ~x197 & ~x200 & ~x504 & ~x531 & ~x760 & ~x779;
assign c3488 =  x47 &  x91 &  x370 & ~x733;
assign c3490 =  x329 & ~x133 & ~x667 & ~x755;
assign c3492 =  x128 &  x152 &  x185 &  x188 &  x241 &  x319 &  x349 &  x378 &  x517 &  x541 &  x548 &  x577 &  x658 &  x686 &  x687 &  x689 &  x691 &  x713 &  x717 &  x739 &  x740 &  x742 & ~x26 & ~x29 & ~x51 & ~x77 & ~x107 & ~x112 & ~x138 & ~x169 & ~x170 & ~x193 & ~x195 & ~x198 & ~x199 & ~x224 & ~x226 & ~x249 & ~x275 & ~x280 & ~x282 & ~x336 & ~x416 & ~x419 & ~x442 & ~x535 & ~x645 & ~x670 & ~x672 & ~x674 & ~x678 & ~x698 & ~x700 & ~x703 & ~x724 & ~x725 & ~x730;
assign c3494 =  x262 &  x540 & ~x142 & ~x229 & ~x260 & ~x388 & ~x426 & ~x507 & ~x582 & ~x669 & ~x727 & ~x754;
assign c3496 = ~x4 & ~x11 & ~x541 & ~x709;
assign c3498 = ~x71 & ~x493;
assign c31 =  x70 &  x97 & ~x406 & ~x490;
assign c33 =  x145 &  x201 &  x259;
assign c35 = ~x40 & ~x46 & ~x122;
assign c37 =  x13 &  x521 & ~x574;
assign c39 =  x173 &  x231;
assign c311 =  x611;
assign c313 =  x98 & ~x434;
assign c315 =  x134 &  x275;
assign c317 =  x131 &  x234 &  x269 &  x288 &  x321 &  x323 &  x373 &  x495 &  x608 &  x655 & ~x417 & ~x445 & ~x479 & ~x506 & ~x565 & ~x722 & ~x759;
assign c319 =  x498 &  x610 & ~x474;
assign c321 =  x362;
assign c323 =  x14 &  x151 &  x263 & ~x120 & ~x476 & ~x645;
assign c325 =  x170;
assign c327 =  x146 &  x173 &  x231 &  x258 & ~x763;
assign c329 =  x258 &  x286 &  x290 &  x301 &  x326 &  x344 &  x411 &  x433 &  x681 &  x687 & ~x308 & ~x555 & ~x646 & ~x780;
assign c331 =  x491 & ~x211;
assign c333 = ~x290 & ~x740;
assign c335 =  x69 &  x153 &  x159 &  x214 &  x289 &  x317 &  x326 &  x355 &  x375 &  x376 &  x486 &  x521 &  x655 & ~x27 & ~x46 & ~x248 & ~x310 & ~x587;
assign c337 = ~x7 & ~x537;
assign c339 = ~x663 & ~x718 & ~x742;
assign c343 =  x219;
assign c345 =  x219 & ~x666;
assign c347 = ~x46 & ~x186 & ~x243;
assign c349 =  x733 & ~x770;
assign c351 =  x106 &  x157 &  x259 &  x737 & ~x8 & ~x394 & ~x475 & ~x526 & ~x537 & ~x583 & ~x723 & ~x751;
assign c353 =  x583 &  x723;
assign c355 = ~x186 & ~x236;
assign c357 = ~x691 & ~x744 & ~x746 & ~x769 & ~x772;
assign c359 =  x14 &  x593;
assign c361 =  x326 &  x454 &  x516 &  x594 &  x631 & ~x387 & ~x614;
assign c363 =  x390;
assign c365 =  x301 &  x454 &  x460 &  x594 & ~x80 & ~x192 & ~x388;
assign c367 =  x180 &  x213 &  x543 &  x712 & ~x251 & ~x332 & ~x523 & ~x582 & ~x663 & ~x736;
assign c369 = ~x290 & ~x291 & ~x347;
assign c371 = ~x737 & ~x739 & ~x745;
assign c373 =  x655 & ~x350 & ~x378;
assign c375 =  x427 &  x454 &  x482 &  x638;
assign c377 = ~x130 & ~x263 & ~x626 & ~x712;
assign c379 =  x212 & ~x658 & ~x714;
assign c381 =  x39 &  x180 &  x269 &  x319 &  x323 &  x492 & ~x612 & ~x624 & ~x691 & ~x720 & ~x736 & ~x737;
assign c383 = ~x291 & ~x348 & ~x656;
assign c385 =  x555 &  x695;
assign c387 =  x19;
assign c389 =  x377 &  x426 &  x454 &  x482 &  x510 &  x581 & ~x35 & ~x79 & ~x140 & ~x388 & ~x528;
assign c391 = ~x235 & ~x543;
assign c393 = ~x75 & ~x291 & ~x516 & ~x631 & ~x687;
assign c395 = ~x75 & ~x291;
assign c397 =  x695;
assign c399 = ~x37 & ~x45 & ~x149 & ~x178 & ~x205;
assign c3101 =  x150 &  x267 &  x323 & ~x201 & ~x218 & ~x252 & ~x304 & ~x397 & ~x443 & ~x591 & ~x648 & ~x725 & ~x742;
assign c3103 =  x231 &  x650 & ~x201;
assign c3105 =  x235 &  x326 &  x465 &  x572 &  x605 &  x626 &  x680 &  x714 &  x739 &  x767 & ~x7 & ~x21 & ~x116 & ~x189 & ~x218 & ~x285 & ~x305 & ~x445 & ~x481 & ~x503 & ~x530 & ~x538 & ~x650 & ~x694 & ~x695 & ~x725 & ~x727 & ~x761;
assign c3107 =  x191;
assign c3109 = ~x476 & ~x615 & ~x701 & ~x718 & ~x738 & ~x745 & ~x769;
assign c3111 =  x67 &  x258 &  x301 &  x317 &  x459 &  x621 & ~x79;
assign c3113 =  x709 & ~x46 & ~x47 & ~x64 & ~x209;
assign c3115 = ~x75 & ~x120 & ~x350;
assign c3117 =  x173 &  x231;
assign c3119 =  x314 &  x622;
assign c3121 =  x15 &  x96 &  x683 & ~x120 & ~x496;
assign c3123 =  x62;
assign c3125 =  x219;
assign c3127 =  x210 &  x238 &  x351 &  x684 & ~x64 & ~x115 & ~x364 & ~x445 & ~x506 & ~x731 & ~x770;
assign c3129 =  x182 &  x683 & ~x490 & ~x518;
assign c3131 = ~x544;
assign c3133 =  x121 &  x231 &  x288 &  x289 &  x399 &  x427 &  x429 &  x464 &  x539 &  x567 &  x581 &  x609 &  x656 &  x718 & ~x0 & ~x418 & ~x444 & ~x479 & ~x529 & ~x673 & ~x699 & ~x782;
assign c3135 =  x205 &  x289 &  x317 &  x318 &  x323 &  x404 &  x411 &  x518 &  x521 &  x549 &  x550 &  x604 &  x679 &  x718 & ~x14 & ~x199 & ~x284 & ~x304 & ~x313 & ~x330 & ~x364 & ~x425 & ~x469 & ~x611 & ~x754;
assign c3137 =  x15 &  x150 &  x262 &  x291 & ~x342 & ~x736;
assign c3139 = ~x75 & ~x186 & ~x544 & ~x626;
assign c3143 =  x761;
assign c3145 =  x454 & ~x770;
assign c3147 = ~x75 & ~x127 & ~x159 & ~x177 & ~x690;
assign c3149 = ~x291 & ~x634 & ~x744;
assign c3151 =  x493 & ~x378 & ~x518;
assign c3153 =  x386 &  x414 &  x594 & ~x500;
assign c3155 =  x90;
assign c3157 =  x176 &  x241 &  x404 &  x432 &  x434 &  x693 &  x744 &  x745 & ~x613 & ~x621;
assign c3159 =  x69 & ~x517 & ~x741 & ~x769;
assign c3161 = ~x45 & ~x131 & ~x209;
assign c3163 =  x607 &  x764 &  x765 &  x767 &  x774 &  x775 & ~x7 & ~x472 & ~x780;
assign c3165 =  x153 &  x177 &  x181 &  x242 &  x266 &  x289 &  x290 &  x458 &  x550 &  x569 &  x571 & ~x58 & ~x109 & ~x144 & ~x191 & ~x280 & ~x287 & ~x302 & ~x360 & ~x391 & ~x476 & ~x479 & ~x526 & ~x566 & ~x592 & ~x610 & ~x616 & ~x645 & ~x698 & ~x704 & ~x705;
assign c3167 =  x14 &  x411 &  x427 &  x465 &  x548 &  x549 &  x581 & ~x52 & ~x115 & ~x145 & ~x170 & ~x306 & ~x337 & ~x451 & ~x479;
assign c3169 =  x464 &  x572 &  x767 & ~x686;
assign c3171 =  x610 & ~x117 & ~x145;
assign c3173 =  x303;
assign c3175 =  x333;
assign c3177 = ~x75 & ~x206 & ~x265 & ~x322;
assign c3179 =  x18 &  x289 &  x298 &  x432 &  x572 & ~x174 & ~x247 & ~x419 & ~x470;
assign c3181 = ~x717 & ~x744 & ~x745;
assign c3183 =  x118 &  x231;
assign c3185 =  x118 &  x231 &  x259 & ~x50;
assign c3187 =  x182 & ~x630 & ~x714;
assign c3189 =  x453 &  x665;
assign c3191 =  x173 & ~x539;
assign c3193 =  x639;
assign c3195 =  x118 &  x190 & ~x441 & ~x530;
assign c3197 = ~x319 & ~x716 & ~x772;
assign c3199 = ~x319 & ~x404;
assign c3201 =  x248;
assign c3203 =  x173 & ~x537;
assign c3205 =  x140;
assign c3207 =  x173 &  x202 &  x231 &  x259;
assign c3209 =  x182 &  x184 &  x627 & ~x316 & ~x663;
assign c3211 = ~x383 & ~x718 & ~x737 & ~x769;
assign c3213 = ~x12 & ~x177 & ~x206 & ~x209;
assign c3215 =  x359;
assign c3217 =  x314 &  x621;
assign c3219 = ~x46 & ~x126 & ~x154 & ~x210 & ~x237;
assign c3221 =  x390;
assign c3223 =  x289 &  x298 &  x521 &  x540 &  x543 &  x679 & ~x29 & ~x366 & ~x370 & ~x395 & ~x553 & ~x566 & ~x646;
assign c3225 = ~x717 & ~x739 & ~x740;
assign c3227 = ~x16 & ~x65 & ~x127 & ~x158;
assign c3229 =  x732;
assign c3231 =  x465 &  x632 &  x662 &  x679 &  x683 &  x719 &  x768 & ~x57 & ~x117 & ~x174 & ~x393 & ~x475 & ~x751;
assign c3233 =  x620;
assign c3235 =  x15 & ~x372;
assign c3237 =  x239 &  x487 &  x520 &  x767 & ~x0;
assign c3239 =  x733 & ~x770;
assign c3241 =  x162 & ~x33 & ~x554;
assign c3243 =  x303;
assign c3245 =  x678 &  x706 &  x777;
assign c3247 = ~x11 & ~x158 & ~x205 & ~x210 & ~x236;
assign c3249 = ~x206 & ~x207 & ~x212;
assign c3251 =  x40 &  x118 &  x229;
assign c3253 =  x128 & ~x120 & ~x518 & ~x748;
assign c3255 =  x62 &  x259;
assign c3257 =  x15 &  x123 &  x159 &  x210 &  x290 &  x297 &  x403 &  x515 &  x655 &  x689 & ~x64 & ~x313 & ~x749;
assign c3259 =  x76 &  x289 & ~x189;
assign c3261 =  x441;
assign c3263 = ~x149 & ~x207 & ~x663;
assign c3265 =  x762;
assign c3267 =  x454 &  x650;
assign c3269 =  x162 &  x231 & ~x553;
assign c3271 = ~x177 & ~x186 & ~x291;
assign c3273 =  x534;
assign c3275 =  x173 & ~x636;
assign c3277 =  x11 & ~x188 & ~x383 & ~x540;
assign c3279 = ~x40 & ~x123;
assign c3281 = ~x179 & ~x578;
assign c3283 = ~x11 & ~x46 & ~x210;
assign c3285 =  x90 &  x219;
assign c3287 = ~x75 & ~x383 & ~x597 & ~x606 & ~x634 & ~x774;
assign c3289 = ~x120 & ~x691 & ~x737 & ~x741 & ~x769;
assign c3291 = ~x94 & ~x124 & ~x689;
assign c3293 = ~x539 & ~x545 & ~x574 & ~x601 & ~x630;
assign c3295 =  x454 &  x482 & ~x77 & ~x275 & ~x641;
assign c3297 =  x257;
assign c3299 =  x555;
assign c3301 =  x627 &  x712 & ~x742;
assign c3303 =  x14 &  x510 & ~x77;
assign c3305 = ~x265 & ~x323 & ~x352;
assign c3307 =  x257 &  x462;
assign c3309 = ~x178 & ~x208 & ~x236;
assign c3311 = ~x65 & ~x207 & ~x212;
assign c3313 =  x498;
assign c3315 =  x130 &  x262 &  x270 &  x289 &  x318 &  x373 &  x516 &  x521 &  x679 & ~x198 & ~x304 & ~x308 & ~x525 & ~x583;
assign c3317 =  x159 &  x182 &  x289 &  x427 &  x521 &  x569 &  x581 &  x609 &  x681 & ~x35 & ~x167;
assign c3319 =  x90;
assign c3321 =  x14 &  x295 &  x627 & ~x770 & ~x776;
assign c3323 =  x557 &  x703;
assign c3325 =  x18 &  x205 &  x767 & ~x200 & ~x253 & ~x471 & ~x529 & ~x536 & ~x611 & ~x670 & ~x762;
assign c3327 =  x121 &  x131 &  x150 &  x205 &  x233 &  x261 &  x289 &  x352 &  x576 &  x681 &  x687 &  x716 &  x767 & ~x26 & ~x145 & ~x539;
assign c3329 = ~x46 & ~x47 & ~x293 & ~x295;
assign c3331 =  x652 & ~x210;
assign c3333 =  x242 &  x608 &  x655 &  x707 &  x768 & ~x110 & ~x147 & ~x446;
assign c3335 =  x150 &  x204 &  x233 &  x240 &  x270 &  x289 &  x293 &  x321 &  x457 &  x459 &  x462 &  x521 &  x579 &  x595 &  x600 &  x652 &  x683 &  x713 &  x767 &  x768 & ~x4 & ~x26 & ~x250 & ~x279 & ~x306 & ~x338 & ~x389 & ~x395 & ~x446 & ~x475 & ~x478 & ~x530 & ~x536 & ~x642 & ~x645 & ~x697 & ~x758;
assign c3337 = ~x263 & ~x543 & ~x544;
assign c3339 =  x14 & ~x518;
assign c3341 =  x74 &  x159 &  x215 &  x262 &  x289 &  x299 &  x350 &  x406 &  x409 &  x513 &  x628 &  x636 &  x651 &  x679 &  x683 &  x720 &  x740 & ~x7 & ~x34 & ~x110 & ~x136 & ~x286 & ~x334 & ~x370 & ~x443 & ~x610 & ~x619 & ~x701 & ~x781;
assign c3343 =  x148 &  x260 &  x262 &  x269 &  x271 &  x318 &  x323 &  x345 &  x404 &  x406 &  x429 &  x461 &  x521 &  x569 &  x570 &  x571 &  x635 &  x659 &  x681 &  x711 &  x715 &  x737 &  x740 &  x768 & ~x56 & ~x113 & ~x116 & ~x168 & ~x173 & ~x253 & ~x277 & ~x281 & ~x304 & ~x366 & ~x474 & ~x529 & ~x560 & ~x563 & ~x584 & ~x672 & ~x675 & ~x697 & ~x723;
assign c3345 = ~x122 & ~x159 & ~x215 & ~x295;
assign c3347 =  x515 &  x571 &  x628 & ~x340 & ~x362 & ~x378 & ~x481;
assign c3349 =  x45 & ~x518 & ~x742;
assign c3351 = ~x47 & ~x158 & ~x179 & ~x319;
assign c3353 =  x257 &  x639;
assign c3355 =  x11 & ~x148 & ~x216 & ~x383 & ~x579 & ~x663;
assign c3357 = ~x639 & ~x663 & ~x737 & ~x745;
assign c3359 =  x761;
assign c3361 = ~x684 & ~x716;
assign c3363 =  x15 &  x150 &  x768 & ~x35 & ~x422 & ~x540 & ~x696;
assign c3365 =  x92 &  x151 &  x187 &  x289 &  x400 &  x467 &  x738 & ~x13 & ~x310 & ~x667;
assign c3367 =  x19 &  x260 & ~x145;
assign c3369 =  x158 &  x576 & ~x344 & ~x551;
assign c3371 =  x508;
assign c3373 =  x558 &  x729;
assign c3375 =  x628 & ~x191 & ~x630 & ~x770;
assign c3377 =  x231;
assign c3379 =  x248;
assign c3381 =  x234 &  x260 &  x270 &  x289 &  x316 &  x372 &  x379 &  x383 &  x404 &  x405 &  x428 &  x433 &  x436 &  x462 &  x488 &  x524 &  x549 &  x567 &  x569 &  x608 &  x609 &  x634 &  x689 &  x717 & ~x0 & ~x2 & ~x50 & ~x52 & ~x196 & ~x225 & ~x359 & ~x363 & ~x500 & ~x506 & ~x559 & ~x643 & ~x646 & ~x669 & ~x702 & ~x755 & ~x758;
assign c3383 = ~x322 & ~x574 & ~x630 & ~x737;
assign c3385 = ~x47 & ~x291 & ~x516;
assign c3387 = ~x157 & ~x177 & ~x404;
assign c3389 = ~x625;
assign c3391 = ~x11 & ~x12 & ~x75 & ~x94 & ~x122;
assign c3393 =  x73 &  x214 &  x262 &  x330 &  x344 &  x408 &  x427 &  x428 &  x603 &  x626 &  x627 & ~x21 & ~x50 & ~x312 & ~x418 & ~x584 & ~x697;
assign c3395 = ~x290 & ~x743 & ~x744 & ~x772;
assign c3397 = ~x206;
assign c3399 = ~x717 & ~x738;
assign c3401 = ~x95 & ~x157 & ~x178 & ~x233;
assign c3403 =  x258 &  x639;
assign c3405 =  x186 & ~x91 & ~x597;
assign c3407 =  x40 &  x71 &  x178 &  x212 & ~x77 & ~x105 & ~x140 & ~x148 & ~x300 & ~x309 & ~x316 & ~x414 & ~x427 & ~x501 & ~x568 & ~x624 & ~x672 & ~x702 & ~x735 & ~x765;
assign c3409 =  x655 & ~x518 & ~x693;
assign c3411 = ~x627 & ~x661;
assign c3413 =  x222;
assign c3415 = ~x40 & ~x126;
assign c3417 =  x171;
assign c3419 = ~x737 & ~x745 & ~x769;
assign c3421 = ~x626 & ~x663 & ~x711;
assign c3423 =  x453 &  x497 & ~x8 & ~x247 & ~x448;
assign c3425 = ~x132 & ~x383 & ~x597 & ~x691 & ~x770;
assign c3427 =  x372 & ~x45;
assign c3429 = ~x605;
assign c3431 =  x231 &  x344 &  x375 & ~x284 & ~x766;
assign c3433 =  x248;
assign c3435 =  x14 &  x38 & ~x540;
assign c3437 =  x14 &  x67 &  x125 &  x178 &  x432 &  x768 & ~x34 & ~x88 & ~x338 & ~x559 & ~x650 & ~x702 & ~x763;
assign c3439 = ~x130 & ~x627 & ~x656;
assign c3441 =  x331;
assign c3443 =  x219;
assign c3445 = ~x372 & ~x653 & ~x690;
assign c3447 =  x158 &  x159 &  x242 &  x262 &  x269 &  x271 &  x383 &  x438 &  x492 &  x547 &  x712 &  x716 &  x740 & ~x0 & ~x24 & ~x283 & ~x338 & ~x370 & ~x441 & ~x442 & ~x452 & ~x526 & ~x565 & ~x647 & ~x674 & ~x783;
assign c3449 =  x184 &  x239 & ~x518;
assign c3451 =  x248;
assign c3453 =  x262 &  x431 & ~x553 & ~x658;
assign c3455 = ~x149 & ~x627 & ~x656;
assign c3457 =  x93 &  x130 &  x177 &  x182 &  x261 &  x263 &  x265 &  x270 &  x289 &  x347 &  x406 &  x460 &  x519 &  x571 &  x740 &  x743 &  x767 & ~x4 & ~x6 & ~x108 & ~x140 & ~x144 & ~x162 & ~x218 & ~x226 & ~x230 & ~x245 & ~x247 & ~x274 & ~x282 & ~x285 & ~x305 & ~x342 & ~x397 & ~x420 & ~x506 & ~x536 & ~x563 & ~x674 & ~x701 & ~x755;
assign c3459 =  x498 &  x526 &  x638;
assign c3461 = ~x120 & ~x130 & ~x157 & ~x158 & ~x178;
assign c3463 =  x78 &  x767;
assign c3465 =  x44 &  x582 &  x638;
assign c3467 = ~x120 & ~x630 & ~x663 & ~x742;
assign c3469 =  x242 &  x260 &  x353 &  x374 &  x461 &  x486 &  x491 &  x523 &  x548 &  x651 &  x767 & ~x22 & ~x161 & ~x252 & ~x340 & ~x480 & ~x530 & ~x564 & ~x723;
assign c3471 =  x131 &  x158 &  x159 &  x178 &  x262 &  x265 &  x289 &  x326 &  x354 &  x355 &  x401 &  x404 &  x430 &  x460 &  x461 &  x490 &  x516 &  x544 &  x545 &  x547 &  x552 &  x604 &  x718 &  x738 &  x740 & ~x2 & ~x54 & ~x80 & ~x82 & ~x83 & ~x110 & ~x113 & ~x116 & ~x145 & ~x162 & ~x163 & ~x164 & ~x170 & ~x171 & ~x192 & ~x246 & ~x253 & ~x254 & ~x256 & ~x276 & ~x307 & ~x310 & ~x330 & ~x340 & ~x366 & ~x389 & ~x442 & ~x451 & ~x499 & ~x500 & ~x529 & ~x533 & ~x557 & ~x564 & ~x585 & ~x617 & ~x618 & ~x672 & ~x674 & ~x702 & ~x731 & ~x753 & ~x759 & ~x760 & ~x762;
assign c3473 =  x270 &  x289 &  x382 &  x491 &  x521 &  x522 &  x570 &  x604 &  x718 &  x767 & ~x11 & ~x26 & ~x27 & ~x145 & ~x363 & ~x385 & ~x414 & ~x417 & ~x425 & ~x533 & ~x537 & ~x591 & ~x646 & ~x648;
assign c3475 = ~x46 & ~x214 & ~x349;
assign c3477 = ~x47 & ~x153 & ~x178 & ~x204;
assign c3479 =  x15 &  x745 & ~x742;
assign c3481 = ~x122 & ~x214 & ~x265;
assign c3483 = ~x132 & ~x358 & ~x489 & ~x517;
assign c3485 =  x78;
assign c3489 =  x341;
assign c3491 =  x611;
assign c3493 = ~x95 & ~x716 & ~x717 & ~x772;
assign c3495 =  x256;
assign c3497 = ~x290 & ~x319 & ~x346 & ~x430;
assign c3499 =  x248;
assign c40 =  x134 &  x219 &  x331 &  x752 & ~x28 & ~x168;
assign c42 =  x231 &  x568 & ~x197 & ~x224 & ~x250 & ~x615 & ~x708 & ~x738 & ~x745 & ~x746 & ~x747 & ~x756 & ~x771;
assign c44 =  x43 &  x462 & ~x54 & ~x653 & ~x711 & ~x772 & ~x773;
assign c46 = ~x680 & ~x719 & ~x739 & ~x749 & ~x757 & ~x771;
assign c48 = ~x5 & ~x37 & ~x53 & ~x57 & ~x61 & ~x79 & ~x82 & ~x85 & ~x90 & ~x107 & ~x116 & ~x140 & ~x143 & ~x171 & ~x248 & ~x305 & ~x365 & ~x393 & ~x420 & ~x586 & ~x691 & ~x708 & ~x709 & ~x717 & ~x718 & ~x719 & ~x720 & ~x727 & ~x736 & ~x737 & ~x738 & ~x739 & ~x740 & ~x741 & ~x742 & ~x744 & ~x745 & ~x746 & ~x754 & ~x758 & ~x765;
assign c410 = ~x3 & ~x20 & ~x114 & ~x521;
assign c412 =  x299 &  x662 & ~x3 & ~x145 & ~x219 & ~x247 & ~x309 & ~x364 & ~x651 & ~x693;
assign c414 = ~x26 & ~x35 & ~x96 & ~x472 & ~x475 & ~x528 & ~x534 & ~x757 & ~x769;
assign c416 =  x355 & ~x1 & ~x47 & ~x62 & ~x162 & ~x172 & ~x190 & ~x218 & ~x229 & ~x247 & ~x257 & ~x359 & ~x473 & ~x500 & ~x536 & ~x650 & ~x692 & ~x697 & ~x727;
assign c418 =  x285 &  x341 &  x555 & ~x3 & ~x18 & ~x19 & ~x24 & ~x112 & ~x169 & ~x171 & ~x198 & ~x255 & ~x388 & ~x419 & ~x477 & ~x479 & ~x507 & ~x531 & ~x535 & ~x559 & ~x562 & ~x698 & ~x708 & ~x728 & ~x729 & ~x737 & ~x738 & ~x739 & ~x740 & ~x741 & ~x742 & ~x744 & ~x745 & ~x747 & ~x765 & ~x766 & ~x769;
assign c420 =  x231 &  x412 &  x454 &  x456 &  x468 &  x568 &  x595 &  x596 &  x690 & ~x29 & ~x87 & ~x145 & ~x444 & ~x472 & ~x476 & ~x780;
assign c422 =  x259 &  x316 &  x320 &  x357 &  x457 &  x546 &  x638 &  x679 &  x692 & ~x111 & ~x171 & ~x219 & ~x255 & ~x416 & ~x444 & ~x447 & ~x562 & ~x703 & ~x727 & ~x754 & ~x781;
assign c424 =  x14 &  x175 &  x238 &  x357 &  x494 &  x612 & ~x51 & ~x108 & ~x224 & ~x364 & ~x781;
assign c426 = ~x17 & ~x78 & ~x135 & ~x272 & ~x381 & ~x474 & ~x587 & ~x617;
assign c428 =  x42 & ~x249 & ~x473 & ~x653 & ~x690 & ~x711 & ~x713 & ~x718 & ~x719 & ~x739;
assign c430 = ~x3 & ~x9 & ~x33 & ~x36 & ~x60 & ~x62 & ~x63 & ~x89 & ~x113 & ~x116 & ~x135 & ~x163 & ~x248 & ~x295 & ~x311 & ~x421 & ~x445 & ~x531 & ~x532 & ~x534 & ~x560 & ~x587 & ~x615 & ~x730 & ~x753 & ~x757 & ~x770 & ~x776;
assign c432 = ~x79 & ~x118 & ~x219 & ~x247 & ~x301 & ~x615 & ~x625 & ~x678;
assign c434 =  x228 &  x696 &  x750;
assign c436 =  x97 & ~x16 & ~x76 & ~x708 & ~x709 & ~x710 & ~x711 & ~x737 & ~x739 & ~x740 & ~x745 & ~x747;
assign c438 =  x284 &  x341 &  x703 & ~x222;
assign c440 =  x244 &  x318 &  x577 &  x685 &  x690 & ~x16 & ~x87 & ~x92 & ~x307;
assign c442 =  x267 &  x483 &  x512 &  x652 &  x718 & ~x134 & ~x135 & ~x420 & ~x700 & ~x776;
assign c444 =  x201 &  x229 &  x268 &  x314 &  x368 &  x412 &  x439 &  x456 &  x512 &  x568 &  x605 &  x662 & ~x35 & ~x77 & ~x87;
assign c446 = ~x3 & ~x37 & ~x64 & ~x134 & ~x146 & ~x162 & ~x174 & ~x190 & ~x201 & ~x276 & ~x396 & ~x499 & ~x612 & ~x665 & ~x668 & ~x678 & ~x754;
assign c448 =  x259 &  x356 &  x400 &  x568 &  x637 &  x665 &  x714 & ~x28 & ~x87 & ~x472;
assign c450 = ~x290 & ~x292 & ~x769;
assign c452 =  x13 &  x349 &  x631 & ~x27 & ~x219 & ~x247 & ~x284 & ~x447 & ~x749 & ~x762 & ~x779;
assign c454 =  x182 &  x564 &  x707 &  x735 & ~x2 & ~x27 & ~x194 & ~x224 & ~x615 & ~x671 & ~x726;
assign c456 =  x725;
assign c458 =  x183 &  x208 &  x238 &  x243 &  x289 &  x314 &  x344 &  x521 &  x596 &  x684 & ~x18 & ~x24 & ~x133 & ~x134 & ~x282 & ~x673;
assign c460 = ~x3 & ~x29 & ~x48 & ~x82 & ~x85 & ~x112 & ~x192 & ~x224 & ~x249 & ~x262 & ~x333 & ~x336 & ~x337 & ~x389 & ~x393 & ~x418 & ~x419 & ~x448 & ~x474 & ~x479 & ~x493 & ~x558 & ~x615 & ~x619 & ~x643 & ~x673 & ~x697 & ~x753 & ~x757 & ~x758 & ~x780;
assign c462 =  x13 &  x214 &  x714 & ~x166 & ~x172 & ~x248 & ~x419 & ~x444 & ~x445 & ~x528 & ~x530 & ~x668 & ~x724 & ~x734;
assign c464 =  x330 &  x639 &  x651 &  x683 &  x687 &  x692 &  x720 & ~x50 & ~x57 & ~x310;
assign c466 = ~x26 & ~x37 & ~x51 & ~x62 & ~x163 & ~x315 & ~x415 & ~x421 & ~x530 & ~x612 & ~x668;
assign c468 =  x316 & ~x3 & ~x37 & ~x46 & ~x58 & ~x62 & ~x77 & ~x110 & ~x197 & ~x250 & ~x254 & ~x280 & ~x282 & ~x367 & ~x472 & ~x503 & ~x504 & ~x533 & ~x615 & ~x618 & ~x737 & ~x738 & ~x739 & ~x741 & ~x744 & ~x745 & ~x746 & ~x747 & ~x773;
assign c470 =  x179 &  x314 &  x441 &  x708 &  x714 & ~x91;
assign c472 =  x184 &  x231 &  x235 &  x291 &  x357 &  x551 &  x573 &  x596 &  x623 &  x628 &  x651 &  x692 &  x720 & ~x25 & ~x78 & ~x86 & ~x141 & ~x171 & ~x280 & ~x421 & ~x669 & ~x782;
assign c474 =  x245 &  x717 & ~x2 & ~x3 & ~x106 & ~x111 & ~x119 & ~x134 & ~x146 & ~x162 & ~x255 & ~x282 & ~x393 & ~x758;
assign c476 =  x237 &  x484 &  x552 &  x568 &  x608 &  x624 &  x692 & ~x3 & ~x247 & ~x504 & ~x612 & ~x618 & ~x640 & ~x668 & ~x780;
assign c478 = ~x107 & ~x127 & ~x234 & ~x269 & ~x363;
assign c480 =  x178 &  x271 &  x346 &  x372 &  x443 &  x467 &  x573 &  x715 &  x719 & ~x22 & ~x106 & ~x134 & ~x504 & ~x645 & ~x728;
assign c482 =  x372 & ~x22 & ~x91 & ~x118 & ~x119 & ~x133 & ~x162 & ~x190 & ~x218 & ~x247 & ~x591 & ~x706 & ~x725 & ~x765;
assign c484 =  x356 &  x750 & ~x6 & ~x58 & ~x76 & ~x86 & ~x107 & ~x142 & ~x224 & ~x252 & ~x311 & ~x389 & ~x503 & ~x531 & ~x618 & ~x673 & ~x700 & ~x728 & ~x737 & ~x738 & ~x739 & ~x740 & ~x743 & ~x745 & ~x746 & ~x747 & ~x757 & ~x759 & ~x765 & ~x769 & ~x773;
assign c486 = ~x1 & ~x21 & ~x35 & ~x48 & ~x50 & ~x62 & ~x106 & ~x134 & ~x219 & ~x222 & ~x304 & ~x311 & ~x368 & ~x423 & ~x486 & ~x534 & ~x588 & ~x671 & ~x754 & ~x783;
assign c488 =  x719 &  x768 & ~x2 & ~x26 & ~x51 & ~x163 & ~x201 & ~x219 & ~x615 & ~x640 & ~x645 & ~x780 & ~x783;
assign c490 =  x659 & ~x0 & ~x5 & ~x6 & ~x7 & ~x8 & ~x10 & ~x11 & ~x17 & ~x19 & ~x24 & ~x25 & ~x26 & ~x27 & ~x28 & ~x29 & ~x30 & ~x31 & ~x32 & ~x33 & ~x34 & ~x48 & ~x49 & ~x50 & ~x51 & ~x53 & ~x57 & ~x78 & ~x79 & ~x85 & ~x86 & ~x107 & ~x110 & ~x111 & ~x112 & ~x135 & ~x137 & ~x140 & ~x142 & ~x143 & ~x145 & ~x167 & ~x172 & ~x173 & ~x191 & ~x194 & ~x198 & ~x199 & ~x201 & ~x219 & ~x224 & ~x225 & ~x247 & ~x249 & ~x254 & ~x255 & ~x278 & ~x280 & ~x285 & ~x305 & ~x306 & ~x307 & ~x310 & ~x311 & ~x334 & ~x335 & ~x336 & ~x337 & ~x360 & ~x364 & ~x389 & ~x391 & ~x392 & ~x395 & ~x421 & ~x422 & ~x423 & ~x447 & ~x476 & ~x501 & ~x503 & ~x504 & ~x529 & ~x530 & ~x532 & ~x534 & ~x535 & ~x558 & ~x559 & ~x586 & ~x587 & ~x589 & ~x590 & ~x616 & ~x617 & ~x642 & ~x645 & ~x670 & ~x672 & ~x698 & ~x699 & ~x702 & ~x706 & ~x726 & ~x727 & ~x749 & ~x754 & ~x755 & ~x759 & ~x762 & ~x780 & ~x783;
assign c492 =  x355 & ~x162 & ~x678 & ~x692 & ~x706 & ~x780;
assign c494 =  x400 &  x526 &  x552 &  x568 &  x611 & ~x27 & ~x108 & ~x361 & ~x416 & ~x646 & ~x727;
assign c496 = ~x244 & ~x278 & ~x305 & ~x348 & ~x534 & ~x754;
assign c498 = ~x34 & ~x59 & ~x107 & ~x278 & ~x393 & ~x407 & ~x435 & ~x450 & ~x505 & ~x530 & ~x644;
assign c4100 = ~x272 & ~x515;
assign c4102 =  x623 & ~x28 & ~x49 & ~x504 & ~x615 & ~x684 & ~x758;
assign c4104 =  x42 &  x229 &  x235 &  x340 &  x396 &  x496 &  x521 &  x554 &  x598 &  x608 & ~x7 & ~x25 & ~x55 & ~x109 & ~x167 & ~x251 & ~x504;
assign c4106 =  x356 &  x662 & ~x20 & ~x133 & ~x134 & ~x504 & ~x558 & ~x615 & ~x762 & ~x775 & ~x777 & ~x783;
assign c4108 =  x181 &  x235 &  x546 &  x554 &  x687 &  x715 &  x720 & ~x83 & ~x145 & ~x336 & ~x673 & ~x758;
assign c4110 =  x200;
assign c4112 =  x752 & ~x720 & ~x745 & ~x771;
assign c4114 =  x201 & ~x46 & ~x737 & ~x743;
assign c4116 =  x14 & ~x2 & ~x24 & ~x391 & ~x396 & ~x650 & ~x705 & ~x721 & ~x727;
assign c4118 =  x289 &  x355 &  x543 &  x546 & ~x62 & ~x247 & ~x364 & ~x392 & ~x419 & ~x472 & ~x668 & ~x706 & ~x721 & ~x723 & ~x778 & ~x780;
assign c4120 =  x45 &  x235 &  x314 &  x443 &  x484 &  x567 &  x568 &  x580 &  x651 &  x665 &  x721 & ~x109 & ~x782;
assign c4122 =  x355 & ~x30 & ~x82 & ~x110 & ~x169 & ~x194 & ~x201 & ~x280 & ~x284 & ~x304 & ~x312 & ~x332 & ~x333 & ~x339 & ~x359 & ~x364 & ~x416 & ~x528 & ~x668 & ~x678 & ~x692 & ~x753 & ~x765 & ~x774 & ~x775;
assign c4124 = ~x0 & ~x4 & ~x5 & ~x7 & ~x8 & ~x11 & ~x18 & ~x19 & ~x20 & ~x21 & ~x24 & ~x25 & ~x27 & ~x29 & ~x30 & ~x31 & ~x33 & ~x34 & ~x37 & ~x50 & ~x51 & ~x52 & ~x53 & ~x54 & ~x55 & ~x56 & ~x58 & ~x59 & ~x61 & ~x78 & ~x79 & ~x80 & ~x83 & ~x84 & ~x86 & ~x87 & ~x107 & ~x108 & ~x115 & ~x116 & ~x136 & ~x137 & ~x141 & ~x142 & ~x165 & ~x168 & ~x169 & ~x170 & ~x171 & ~x191 & ~x192 & ~x193 & ~x194 & ~x196 & ~x197 & ~x198 & ~x199 & ~x200 & ~x201 & ~x220 & ~x221 & ~x222 & ~x223 & ~x224 & ~x226 & ~x229 & ~x249 & ~x251 & ~x253 & ~x254 & ~x255 & ~x256 & ~x276 & ~x278 & ~x280 & ~x281 & ~x283 & ~x284 & ~x303 & ~x305 & ~x306 & ~x307 & ~x309 & ~x310 & ~x311 & ~x312 & ~x333 & ~x336 & ~x340 & ~x361 & ~x362 & ~x363 & ~x365 & ~x368 & ~x388 & ~x391 & ~x392 & ~x393 & ~x416 & ~x418 & ~x419 & ~x421 & ~x423 & ~x444 & ~x449 & ~x472 & ~x474 & ~x476 & ~x479 & ~x502 & ~x505 & ~x506 & ~x529 & ~x530 & ~x531 & ~x534 & ~x535 & ~x558 & ~x563 & ~x586 & ~x587 & ~x589 & ~x613 & ~x614 & ~x615 & ~x616 & ~x617 & ~x641 & ~x642 & ~x643 & ~x672 & ~x698 & ~x700 & ~x703 & ~x706 & ~x726 & ~x730 & ~x731 & ~x755 & ~x756 & ~x758 & ~x764 & ~x781 & ~x783;
assign c4126 = ~x81 & ~x559 & ~x615 & ~x627 & ~x634 & ~x685 & ~x712;
assign c4128 =  x14 &  x45 &  x205 &  x568 &  x572 &  x596 &  x609 &  x637 &  x639 &  x690 & ~x728;
assign c4130 =  x44 &  x400 &  x581 &  x596 &  x637 &  x691 & ~x27 & ~x60 & ~x82 & ~x112 & ~x169 & ~x222 & ~x248 & ~x278 & ~x311 & ~x390 & ~x452 & ~x536 & ~x591 & ~x612 & ~x640 & ~x697 & ~x756;
assign c4132 =  x13 &  x42 &  x184 &  x216 &  x218 &  x329 &  x349 &  x372 &  x551 &  x596 & ~x77 & ~x111 & ~x167 & ~x278 & ~x393 & ~x419 & ~x474 & ~x502 & ~x560 & ~x644 & ~x726 & ~x771;
assign c4134 =  x272 &  x383 &  x483 &  x484 &  x524 &  x608 &  x747 & ~x27 & ~x140 & ~x195 & ~x417 & ~x530 & ~x642 & ~x758 & ~x777 & ~x780;
assign c4136 = ~x208 & ~x644 & ~x737 & ~x738 & ~x739 & ~x740;
assign c4138 =  x316 & ~x24 & ~x51 & ~x60 & ~x77 & ~x82 & ~x194 & ~x222 & ~x339 & ~x363 & ~x394 & ~x472 & ~x503 & ~x507 & ~x532 & ~x558 & ~x668 & ~x673 & ~x720 & ~x727 & ~x737 & ~x738 & ~x739 & ~x740 & ~x742 & ~x744 & ~x746 & ~x758 & ~x767 & ~x769 & ~x773;
assign c4140 = ~x1 & ~x2 & ~x3 & ~x6 & ~x17 & ~x27 & ~x28 & ~x33 & ~x47 & ~x48 & ~x49 & ~x62 & ~x63 & ~x77 & ~x107 & ~x173 & ~x219 & ~x226 & ~x284 & ~x304 & ~x339 & ~x419 & ~x436 & ~x475 & ~x590 & ~x615 & ~x670 & ~x671 & ~x698 & ~x726 & ~x763 & ~x775;
assign c4142 =  x270 &  x345 & ~x10 & ~x26 & ~x145 & ~x190 & ~x201 & ~x218 & ~x222 & ~x247 & ~x275 & ~x359 & ~x364 & ~x474 & ~x476 & ~x591 & ~x617 & ~x646 & ~x648 & ~x668 & ~x692 & ~x694 & ~x696 & ~x698 & ~x727 & ~x781;
assign c4144 = ~x18 & ~x21 & ~x25 & ~x90 & ~x169 & ~x197 & ~x251 & ~x276 & ~x305 & ~x306 & ~x615 & ~x617 & ~x681 & ~x708 & ~x711 & ~x718 & ~x719 & ~x736 & ~x739 & ~x742 & ~x744 & ~x745;
assign c4146 =  x182 &  x731 &  x752 & ~x27 & ~x60 & ~x78 & ~x84 & ~x195;
assign c4148 = ~x48 & ~x60 & ~x351 & ~x407 & ~x419 & ~x758;
assign c4150 =  x382 & ~x16 & ~x36 & ~x54 & ~x110 & ~x161 & ~x173 & ~x190 & ~x191 & ~x196 & ~x201 & ~x281 & ~x362 & ~x389 & ~x502 & ~x747 & ~x774;
assign c4152 =  x38 &  x179 &  x233 &  x568 &  x747 & ~x780;
assign c4154 = ~x2 & ~x59 & ~x79 & ~x107 & ~x165 & ~x318 & ~x376;
assign c4156 = ~x269 & ~x318 & ~x765;
assign c4158 =  x235 &  x265 &  x266 &  x295 &  x518 &  x551 &  x568 &  x579 &  x623 &  x651 &  x686 &  x687 &  x744 & ~x29 & ~x113 & ~x311 & ~x613 & ~x645 & ~x674;
assign c4160 = ~x4 & ~x5 & ~x8 & ~x17 & ~x19 & ~x21 & ~x24 & ~x32 & ~x34 & ~x35 & ~x37 & ~x48 & ~x62 & ~x76 & ~x82 & ~x86 & ~x87 & ~x90 & ~x110 & ~x111 & ~x164 & ~x168 & ~x197 & ~x198 & ~x223 & ~x224 & ~x248 & ~x250 & ~x305 & ~x306 & ~x334 & ~x338 & ~x339 & ~x417 & ~x419 & ~x473 & ~x530 & ~x532 & ~x534 & ~x535 & ~x557 & ~x563 & ~x586 & ~x587 & ~x614 & ~x616 & ~x645 & ~x669 & ~x708 & ~x727 & ~x736 & ~x737 & ~x738 & ~x739 & ~x740 & ~x741 & ~x744 & ~x746 & ~x747 & ~x757 & ~x758 & ~x759 & ~x766 & ~x769 & ~x770 & ~x771 & ~x774;
assign c4162 =  x71 &  x327 &  x461 &  x514 &  x518 & ~x2 & ~x22 & ~x25 & ~x30 & ~x336 & ~x389 & ~x447 & ~x502 & ~x588 & ~x653 & ~x726 & ~x754;
assign c4164 = ~x0 & ~x2 & ~x6 & ~x7 & ~x8 & ~x22 & ~x23 & ~x32 & ~x52 & ~x79 & ~x106 & ~x135 & ~x170 & ~x171 & ~x172 & ~x249 & ~x267 & ~x281 & ~x306 & ~x333 & ~x337 & ~x363 & ~x389 & ~x421 & ~x446 & ~x476 & ~x500 & ~x507 & ~x530 & ~x562 & ~x613 & ~x615 & ~x619 & ~x645 & ~x672 & ~x673 & ~x726 & ~x728 & ~x759 & ~x765 & ~x767;
assign c4166 =  x456 &  x484 &  x524 &  x565 &  x609 &  x637 &  x713 & ~x219;
assign c4168 = ~x208 & ~x262 & ~x304 & ~x307;
assign c4170 = ~x11 & ~x36 & ~x44 & ~x84 & ~x172 & ~x308 & ~x390 & ~x613;
assign c4172 = ~x18 & ~x46 & ~x224 & ~x229 & ~x340 & ~x499 & ~x507 & ~x535 & ~x721;
assign c4174 = ~x5 & ~x28 & ~x119 & ~x146 & ~x172 & ~x174 & ~x362 & ~x408 & ~x421 & ~x730;
assign c4176 =  x400 &  x467 & ~x201 & ~x219 & ~x480 & ~x639 & ~x679 & ~x707 & ~x749;
assign c4178 = ~x208 & ~x301;
assign c4180 =  x456 &  x634 &  x746 & ~x28 & ~x133 & ~x218 & ~x219 & ~x762;
assign c4182 = ~x232 & ~x712;
assign c4184 =  x261 &  x290 &  x293 &  x350 &  x578 &  x604 &  x690 & ~x18 & ~x20 & ~x164 & ~x190 & ~x588 & ~x619 & ~x668 & ~x671 & ~x679 & ~x706 & ~x757;
assign c4186 =  x468 &  x484 &  x552 &  x595 &  x608 &  x683 &  x768 & ~x167 & ~x762;
assign c4188 =  x329 &  x372 &  x440 &  x484 &  x568 &  x608 & ~x118 & ~x674;
assign c4190 = ~x262 & ~x381 & ~x769;
assign c4192 =  x206 &  x456 &  x568 &  x652 &  x662 &  x690 &  x714 & ~x198 & ~x247 & ~x252 & ~x777;
assign c4194 =  x219 &  x461 &  x511 &  x528 &  x568;
assign c4196 =  x322 &  x580 &  x692 & ~x62 & ~x118 & ~x146 & ~x168 & ~x219 & ~x221 & ~x335 & ~x338 & ~x339 & ~x393 & ~x757 & ~x781;
assign c4198 = ~x201 & ~x219 & ~x247 & ~x257 & ~x498 & ~x556 & ~x623 & ~x693;
assign c4200 =  x13 & ~x18 & ~x27 & ~x53 & ~x201 & ~x226 & ~x247 & ~x248 & ~x281 & ~x284 & ~x419 & ~x679 & ~x700 & ~x701;
assign c4202 =  x42 &  x331 & ~x4 & ~x23 & ~x51 & ~x53 & ~x87 & ~x112 & ~x137 & ~x165 & ~x170 & ~x336 & ~x362 & ~x560 & ~x643 & ~x711 & ~x728 & ~x739 & ~x740 & ~x745 & ~x771 & ~x783;
assign c4204 =  x235 &  x444 & ~x253;
assign c4206 =  x42 &  x233 &  x257 &  x275 &  x324 &  x331 &  x368 &  x377 &  x433 &  x528 &  x579 & ~x2 & ~x141 & ~x560;
assign c4208 =  x354 &  x662 & ~x18 & ~x26 & ~x62 & ~x88 & ~x90 & ~x104 & ~x172 & ~x197 & ~x693;
assign c4210 = ~x263 & ~x277 & ~x333 & ~x706;
assign c4212 =  x201 &  x399 &  x408 &  x637 & ~x3 & ~x109 & ~x746;
assign c4214 =  x270 &  x298 & ~x64 & ~x133 & ~x134 & ~x146 & ~x308 & ~x365 & ~x534 & ~x651 & ~x721;
assign c4216 =  x13 &  x647;
assign c4218 =  x400 &  x411 &  x546 & ~x62 & ~x90 & ~x201 & ~x247 & ~x472 & ~x507 & ~x640 & ~x693 & ~x749;
assign c4220 =  x271 &  x675 &  x696 & ~x27 & ~x59 & ~x62 & ~x193 & ~x252 & ~x617 & ~x727;
assign c4222 =  x596 & ~x133 & ~x162 & ~x762;
assign c4224 = ~x51 & ~x109 & ~x253 & ~x403 & ~x419 & ~x474 & ~x475 & ~x534 & ~x554;
assign c4226 =  x175 &  x230 &  x275 &  x331 &  x443 &  x552 &  x556 &  x638 & ~x249 & ~x618;
assign c4228 =  x13 &  x14 &  x154 &  x552 &  x608 &  x620 & ~x88;
assign c4230 =  x409 &  x750 & ~x5 & ~x8 & ~x35 & ~x46 & ~x48 & ~x54 & ~x84 & ~x107 & ~x192 & ~x227 & ~x615 & ~x737 & ~x738 & ~x739 & ~x740 & ~x741 & ~x742 & ~x744 & ~x745 & ~x746 & ~x758 & ~x769 & ~x771;
assign c4232 =  x13 &  x16 &  x400 &  x552 & ~x51 & ~x284 & ~x362 & ~x532 & ~x727 & ~x762;
assign c4234 =  x71 &  x266 &  x354 &  x356 & ~x28 & ~x48 & ~x62 & ~x164 & ~x173 & ~x201 & ~x305 & ~x391 & ~x532 & ~x643 & ~x706 & ~x779;
assign c4236 =  x275 &  x314 &  x331 &  x554 &  x584 &  x612 &  x668 &  x696 &  x732 &  x751 & ~x615 & ~x769;
assign c4238 =  x12 &  x14 &  x314 &  x443 &  x470 &  x552 & ~x52 & ~x106 & ~x305 & ~x505 & ~x531;
assign c4240 = ~x262 & ~x740;
assign c4242 =  x266 &  x317 &  x379 &  x405 &  x441 &  x469 & ~x25 & ~x26 & ~x30 & ~x55 & ~x82 & ~x112 & ~x172 & ~x192 & ~x201 & ~x224 & ~x335 & ~x340 & ~x390 & ~x417 & ~x528 & ~x558 & ~x613 & ~x668 & ~x702 & ~x724 & ~x728 & ~x759 & ~x762;
assign c4244 =  x154 &  x205 &  x352 &  x433 &  x526 & ~x2 & ~x3 & ~x17 & ~x29 & ~x48 & ~x63 & ~x142 & ~x171 & ~x221 & ~x280 & ~x615 & ~x643 & ~x673 & ~x698 & ~x726 & ~x737 & ~x738 & ~x739 & ~x745 & ~x765 & ~x768 & ~x774;
assign c4246 = ~x145 & ~x284 & ~x528 & ~x584 & ~x617 & ~x668 & ~x696 & ~x700 & ~x717 & ~x718 & ~x719 & ~x738 & ~x739 & ~x740 & ~x744 & ~x745 & ~x746 & ~x769;
assign c4248 =  x288 &  x289 &  x290 &  x550 &  x658 &  x660 &  x714 &  x716 & ~x28 & ~x30 & ~x55 & ~x78 & ~x90 & ~x105 & ~x119 & ~x172 & ~x173 & ~x194 & ~x219 & ~x255 & ~x280 & ~x310 & ~x339 & ~x368 & ~x388 & ~x390 & ~x393 & ~x445 & ~x533 & ~x534 & ~x585 & ~x591 & ~x615 & ~x641 & ~x642 & ~x645 & ~x671 & ~x697 & ~x726 & ~x727 & ~x782;
assign c4250 =  x38 &  x331 &  x484 &  x522 &  x552 &  x638 &  x665 &  x721 & ~x141 & ~x419 & ~x532;
assign c4252 = ~x24 & ~x62 & ~x119 & ~x146 & ~x408;
assign c4254 =  x631 & ~x51 & ~x76 & ~x106 & ~x112 & ~x133 & ~x134 & ~x145 & ~x229 & ~x312 & ~x361 & ~x450 & ~x530 & ~x589 & ~x703 & ~x759 & ~x765 & ~x777;
assign c4256 =  x175 &  x235 &  x312 &  x647 & ~x364;
assign c4258 =  x271 &  x378 &  x718 & ~x162 & ~x190 & ~x391 & ~x623 & ~x651 & ~x721 & ~x778;
assign c4260 =  x155 &  x230 &  x697 & ~x278 & ~x721;
assign c4262 =  x11 &  x13 &  x14 &  x265 &  x747;
assign c4264 = ~x9 & ~x111 & ~x163 & ~x256 & ~x339 & ~x362 & ~x364 & ~x431 & ~x445 & ~x503 & ~x505 & ~x671 & ~x673;
assign c4266 =  x201 &  x528 &  x552 &  x554;
assign c4268 =  x215 &  x662 & ~x17 & ~x170 & ~x201 & ~x219 & ~x247 & ~x650;
assign c4270 =  x182 &  x184 &  x202 &  x300 &  x341 &  x359 &  x426 &  x443 &  x514 &  x571 &  x601 &  x603 &  x610 & ~x22 & ~x24 & ~x30 & ~x50 & ~x51 & ~x78 & ~x80 & ~x113 & ~x221 & ~x222 & ~x223 & ~x255 & ~x280 & ~x305 & ~x307 & ~x338 & ~x449 & ~x614 & ~x615 & ~x671 & ~x672 & ~x726 & ~x754 & ~x767 & ~x770 & ~x773;
assign c4272 = ~x26 & ~x127 & ~x241 & ~x324 & ~x354 & ~x382;
assign c4274 =  x231 &  x442 &  x467 &  x554 &  x582 &  x608 &  x651 &  x687 &  x693 &  x707 & ~x112 & ~x618;
assign c4276 = ~x24 & ~x25 & ~x161 & ~x253 & ~x390 & ~x521 & ~x584;
assign c4278 =  x70 &  x552 & ~x183;
assign c4280 =  x750 & ~x29 & ~x37 & ~x48 & ~x62 & ~x63 & ~x85 & ~x87 & ~x115 & ~x172 & ~x194 & ~x221 & ~x282 & ~x362 & ~x364 & ~x366 & ~x473 & ~x502 & ~x531 & ~x559 & ~x673 & ~x699 & ~x726 & ~x737 & ~x738 & ~x743 & ~x744 & ~x745 & ~x746 & ~x768 & ~x769 & ~x780;
assign c4282 = ~x7 & ~x21 & ~x29 & ~x30 & ~x49 & ~x50 & ~x56 & ~x85 & ~x201 & ~x247 & ~x253 & ~x256 & ~x363 & ~x472 & ~x552 & ~x558 & ~x580 & ~x669 & ~x678 & ~x727;
assign c4284 = ~x3 & ~x24 & ~x30 & ~x197 & ~x298 & ~x533 & ~x617 & ~x741 & ~x766 & ~x768;
assign c4286 =  x467 &  x526 &  x608 &  x610 &  x637 &  x651 &  x720 & ~x0 & ~x50 & ~x619;
assign c4288 =  x288 &  x779 & ~x0 & ~x35 & ~x36 & ~x49 & ~x50 & ~x54 & ~x57 & ~x59 & ~x62 & ~x82 & ~x135 & ~x249 & ~x252 & ~x276 & ~x419 & ~x475 & ~x613 & ~x758 & ~x765 & ~x767 & ~x770 & ~x773;
assign c4290 = ~x431;
assign c4292 = ~x23 & ~x250 & ~x280 & ~x320 & ~x348 & ~x613 & ~x644 & ~x765;
assign c4294 =  x13 &  x14 &  x152 &  x288 &  x295 &  x299 &  x400 &  x467 &  x486 &  x494 &  x517 &  x550 &  x551 &  x603 &  x648 & ~x25 & ~x33 & ~x49 & ~x62 & ~x78 & ~x113 & ~x192 & ~x419 & ~x587 & ~x615 & ~x616 & ~x618 & ~x700;
assign c4296 = ~x2 & ~x3 & ~x10 & ~x16 & ~x56 & ~x111 & ~x145 & ~x173 & ~x252 & ~x275 & ~x312 & ~x331 & ~x340 & ~x474 & ~x498 & ~x500 & ~x559 & ~x678 & ~x679 & ~x694 & ~x749 & ~x774;
assign c4298 =  x231 &  x331 &  x512 &  x552 &  x568 &  x610 &  x639 &  x655 & ~x5 & ~x53 & ~x62 & ~x304 & ~x506 & ~x531 & ~x673 & ~x700;
assign c4300 =  x239 &  x314 &  x321 &  x349 &  x682 & ~x20 & ~x48 & ~x133 & ~x134 & ~x162 & ~x163 & ~x247 & ~x248 & ~x256 & ~x475 & ~x671 & ~x754 & ~x757;
assign c4302 =  x45 &  x69 &  x218 &  x331 &  x427 &  x668 & ~x3 & ~x26 & ~x50 & ~x62 & ~x168 & ~x194 & ~x281 & ~x617;
assign c4304 =  x345 & ~x11 & ~x218 & ~x274 & ~x332 & ~x680;
assign c4306 =  x316 &  x751 & ~x4 & ~x19 & ~x29 & ~x30 & ~x47 & ~x60 & ~x61 & ~x62 & ~x82 & ~x83 & ~x85 & ~x107 & ~x113 & ~x143 & ~x168 & ~x225 & ~x251 & ~x253 & ~x311 & ~x333 & ~x337 & ~x360 & ~x361 & ~x364 & ~x417 & ~x422 & ~x502 & ~x504 & ~x532 & ~x559 & ~x590 & ~x613 & ~x643 & ~x670 & ~x698 & ~x727 & ~x742 & ~x755 & ~x767 & ~x768 & ~x774;
assign c4308 = ~x222 & ~x264 & ~x470 & ~x543;
assign c4310 =  x13 &  x14 &  x16 &  x233 &  x234 &  x326 &  x329 &  x369 &  x470 &  x484 & ~x7 & ~x196 & ~x278 & ~x282 & ~x419 & ~x698 & ~x756;
assign c4312 =  x13 &  x14 &  x16 &  x44 &  x205 &  x318 &  x384 &  x400 &  x430 &  x438 &  x492 &  x655 & ~x4 & ~x29 & ~x48 & ~x50 & ~x57 & ~x62 & ~x78 & ~x79 & ~x81 & ~x87 & ~x113 & ~x141 & ~x198 & ~x221 & ~x226 & ~x253 & ~x278 & ~x305 & ~x393 & ~x643 & ~x698 & ~x700 & ~x782;
assign c4314 =  x638 &  x731 &  x752 & ~x62 & ~x306;
assign c4316 =  x148 &  x229 &  x297 &  x396 &  x526 &  x536 &  x567 &  x648 & ~x2 & ~x87 & ~x113;
assign c4318 =  x569 &  x609 &  x734 &  x779 & ~x199 & ~x251 & ~x476 & ~x558 & ~x773;
assign c4320 = ~x10 & ~x21 & ~x23 & ~x28 & ~x29 & ~x48 & ~x54 & ~x60 & ~x62 & ~x88 & ~x108 & ~x112 & ~x117 & ~x119 & ~x145 & ~x163 & ~x174 & ~x191 & ~x201 & ~x219 & ~x247 & ~x275 & ~x280 & ~x282 & ~x306 & ~x312 & ~x388 & ~x393 & ~x451 & ~x453 & ~x472 & ~x529 & ~x561 & ~x668 & ~x669 & ~x671 & ~x698 & ~x728 & ~x730 & ~x759 & ~x765 & ~x767 & ~x773 & ~x780;
assign c4322 =  x42 &  x98 &  x288 & ~x2 & ~x8 & ~x20 & ~x25 & ~x33 & ~x55 & ~x57 & ~x60 & ~x82 & ~x86 & ~x111 & ~x167 & ~x196 & ~x199 & ~x222 & ~x227 & ~x249 & ~x251 & ~x282 & ~x390 & ~x392 & ~x418 & ~x532 & ~x559 & ~x560 & ~x645 & ~x681 & ~x756;
assign c4324 =  x687 & ~x133 & ~x174 & ~x190 & ~x218 & ~x678;
assign c4326 = ~x174 & ~x264;
assign c4328 =  x298 &  x300 &  x321 &  x372 &  x580 &  x630 &  x692 &  x714 &  x720 & ~x31 & ~x162 & ~x227 & ~x256 & ~x282 & ~x644 & ~x698;
assign c4330 =  x585;
assign c4332 = ~x17 & ~x191 & ~x231 & ~x263 & ~x348 & ~x617;
assign c4334 =  x14 &  x181 & ~x19 & ~x77 & ~x87 & ~x226 & ~x616 & ~x617 & ~x698 & ~x737 & ~x738 & ~x739 & ~x745 & ~x757 & ~x766 & ~x768 & ~x773;
assign c4336 =  x331 &  x344 &  x359 &  x387 & ~x110 & ~x113 & ~x141 & ~x197 & ~x337 & ~x737 & ~x739 & ~x740 & ~x741 & ~x744 & ~x745 & ~x746 & ~x782;
assign c4338 =  x229 &  x443 &  x484 &  x552 &  x595 &  x665;
assign c4340 =  x356 &  x400 &  x567 &  x573 &  x609 &  x636 & ~x18 & ~x24 & ~x134 & ~x190 & ~x247 & ~x416 & ~x419 & ~x474 & ~x668 & ~x779;
assign c4342 =  x158 &  x205 &  x230 &  x257 &  x265 &  x272 &  x275 &  x300 &  x303 &  x415 &  x439 &  x453 &  x467 &  x554 &  x648 &  x696 & ~x1 & ~x4 & ~x8 & ~x30 & ~x58 & ~x59 & ~x78 & ~x136 & ~x198 & ~x249 & ~x253 & ~x279 & ~x280 & ~x310 & ~x364 & ~x418 & ~x530 & ~x532 & ~x757;
assign c4344 = ~x22 & ~x90 & ~x183 & ~x336 & ~x364 & ~x368 & ~x615 & ~x669 & ~x672 & ~x730 & ~x769 & ~x770;
assign c4346 =  x289 &  x687 &  x690 &  x718 & ~x14 & ~x48 & ~x118 & ~x133 & ~x142 & ~x247 & ~x253 & ~x474 & ~x531 & ~x645;
assign c4348 =  x41 &  x247 &  x331 &  x406 &  x492 &  x514 &  x552 &  x580 &  x595 &  x638 & ~x55 & ~x86 & ~x108 & ~x112 & ~x225 & ~x448 & ~x587;
assign c4350 = ~x598 & ~x613 & ~x711 & ~x739;
assign c4352 =  x13 & ~x37 & ~x48 & ~x59 & ~x393 & ~x698 & ~x738 & ~x739 & ~x740;
assign c4354 =  x231 &  x708 & ~x119 & ~x276 & ~x338 & ~x776;
assign c4356 =  x11 &  x12 &  x14 &  x15 & ~x87 & ~x145 & ~x196 & ~x248 & ~x337 & ~x446;
assign c4358 =  x201 &  x228 &  x256 &  x350 &  x648 & ~x504 & ~x615;
assign c4360 =  x99 &  x175 &  x231 &  x271 &  x288 &  x290 &  x317 &  x322 &  x327 &  x341 &  x427 &  x443 &  x456 &  x462 &  x525 &  x554 &  x567 &  x609 &  x652 &  x665 & ~x58 & ~x112 & ~x113 & ~x135 & ~x534 & ~x674 & ~x783;
assign c4362 =  x567 & ~x27 & ~x29 & ~x114 & ~x308 & ~x449 & ~x615 & ~x645 & ~x681 & ~x684 & ~x708 & ~x710;
assign c4364 =  x648 & ~x26 & ~x30 & ~x32 & ~x34 & ~x51 & ~x56 & ~x59 & ~x85 & ~x115 & ~x142 & ~x166 & ~x168 & ~x170 & ~x253 & ~x282 & ~x390 & ~x419 & ~x476 & ~x559 & ~x589 & ~x680 & ~x782;
assign c4366 = ~x21 & ~x36 & ~x48 & ~x87 & ~x135 & ~x163 & ~x310 & ~x339 & ~x419 & ~x445 & ~x515 & ~x559 & ~x586 & ~x730 & ~x758;
assign c4368 =  x13 &  x462 & ~x5 & ~x54 & ~x62 & ~x83 & ~x110 & ~x145 & ~x196 & ~x201 & ~x224 & ~x279 & ~x419 & ~x721 & ~x756 & ~x761 & ~x780;
assign c4370 = ~x291 & ~x324;
assign c4372 =  x266 &  x269 &  x368 &  x552 & ~x26 & ~x55 & ~x109 & ~x112 & ~x113 & ~x167 & ~x221 & ~x250 & ~x587 & ~x671;
assign c4374 =  x151 &  x175 &  x552 &  x609 &  x623 &  x637 &  x648 &  x651 &  x679;
assign c4376 = ~x262 & ~x272;
assign c4378 =  x409 &  x461 &  x464 &  x492 &  x605 & ~x8 & ~x20 & ~x30 & ~x163 & ~x219 & ~x223 & ~x247 & ~x312 & ~x445 & ~x615 & ~x617 & ~x706 & ~x750 & ~x757 & ~x758 & ~x779;
assign c4380 =  x201 &  x368 &  x424 &  x564 &  x631 &  x751 & ~x0 & ~x47 & ~x48;
assign c4382 =  x175 &  x215 &  x229 &  x640 & ~x3 & ~x87 & ~x364;
assign c4384 =  x298 &  x411 &  x412 &  x517 &  x687 & ~x8 & ~x27 & ~x49 & ~x62 & ~x110 & ~x190 & ~x194 & ~x249 & ~x303 & ~x310 & ~x443 & ~x472 & ~x503 & ~x615 & ~x668 & ~x698 & ~x726 & ~x749;
assign c4386 = ~x190 & ~x219 & ~x284 & ~x477 & ~x556 & ~x577;
assign c4388 =  x42 &  x300 &  x303 &  x415 &  x427 &  x438 &  x568 &  x638 & ~x5 & ~x62 & ~x78 & ~x364 & ~x419 & ~x535 & ~x671 & ~x726 & ~x757;
assign c4390 =  x69 & ~x21 & ~x23 & ~x24 & ~x54 & ~x87 & ~x107 & ~x110 & ~x138 & ~x163 & ~x168 & ~x169 & ~x183 & ~x223 & ~x249 & ~x280 & ~x281 & ~x282 & ~x305 & ~x306 & ~x393 & ~x417 & ~x450 & ~x472 & ~x474 & ~x586 & ~x591 & ~x643 & ~x670 & ~x729 & ~x757 & ~x776;
assign c4392 = ~x51 & ~x55 & ~x83 & ~x85 & ~x142 & ~x196 & ~x250 & ~x252 & ~x307 & ~x336 & ~x366 & ~x375 & ~x474 & ~x475 & ~x532 & ~x618 & ~x727;
assign c4394 =  x733 & ~x16 & ~x37 & ~x59 & ~x90 & ~x141 & ~x449 & ~x534 & ~x702 & ~x737 & ~x738 & ~x740 & ~x742 & ~x744 & ~x745;
assign c4396 =  x124 &  x459 & ~x90 & ~x110 & ~x193 & ~x507 & ~x591 & ~x711 & ~x738 & ~x739;
assign c4398 =  x275 &  x331 &  x406 &  x528 &  x567 &  x570 &  x596 & ~x20 & ~x27 & ~x31 & ~x85 & ~x113 & ~x699 & ~x782;
assign c4400 =  x400 &  x412 &  x568 &  x684 & ~x27 & ~x60 & ~x80 & ~x616 & ~x617 & ~x745 & ~x772 & ~x783;
assign c4402 =  x69 & ~x1 & ~x199 & ~x615 & ~x633 & ~x641 & ~x737 & ~x739 & ~x741 & ~x745 & ~x747 & ~x766;
assign c4404 =  x289 &  x345 & ~x46 & ~x47 & ~x62 & ~x76 & ~x85 & ~x118 & ~x146 & ~x172 & ~x174 & ~x201 & ~x218 & ~x247 & ~x312 & ~x359 & ~x416 & ~x480 & ~x535 & ~x693 & ~x780;
assign c4406 =  x14 &  x275 &  x396 &  x415;
assign c4408 = ~x2 & ~x5 & ~x21 & ~x27 & ~x30 & ~x32 & ~x34 & ~x48 & ~x59 & ~x171 & ~x201 & ~x209 & ~x248 & ~x252 & ~x278 & ~x422 & ~x451 & ~x478 & ~x503 & ~x586 & ~x700 & ~x702 & ~x755 & ~x764;
assign c4410 =  x262 &  x345 &  x631 & ~x36 & ~x76 & ~x79 & ~x145 & ~x162 & ~x163 & ~x173 & ~x190 & ~x218 & ~x219 & ~x228 & ~x275 & ~x276 & ~x419 & ~x445 & ~x508 & ~x588 & ~x698 & ~x721;
assign c4412 =  x313 & ~x46 & ~x50 & ~x165 & ~x532 & ~x720 & ~x737 & ~x738 & ~x742 & ~x743 & ~x744 & ~x745 & ~x746 & ~x747 & ~x768 & ~x770 & ~x772;
assign c4414 =  x234 &  x261 &  x602 &  x630 & ~x28 & ~x48 & ~x76 & ~x87 & ~x118 & ~x145 & ~x146 & ~x173 & ~x419 & ~x451 & ~x528 & ~x765;
assign c4416 =  x265 &  x272 &  x327 &  x383 &  x470 &  x603 &  x655 &  x662 &  x719 & ~x4 & ~x21 & ~x22 & ~x25 & ~x29 & ~x35 & ~x85 & ~x111 & ~x137 & ~x140 & ~x164 & ~x171 & ~x219 & ~x248 & ~x447 & ~x502 & ~x503 & ~x674 & ~x728 & ~x757 & ~x779;
assign c4418 =  x13 &  x14 &  x349 &  x356 &  x429 & ~x25 & ~x27 & ~x50 & ~x87 & ~x115 & ~x143 & ~x219 & ~x226 & ~x279 & ~x389 & ~x472 & ~x563 & ~x586 & ~x589 & ~x734 & ~x749;
assign c4420 = ~x17 & ~x190 & ~x201 & ~x247 & ~x248 & ~x359 & ~x648 & ~x665 & ~x678 & ~x708 & ~x774;
assign c4422 =  x261 &  x517 & ~x48 & ~x360 & ~x396 & ~x472 & ~x623 & ~x680 & ~x749;
assign c4424 =  x12 & ~x36 & ~x54 & ~x671 & ~x708 & ~x709 & ~x718 & ~x736 & ~x739 & ~x743 & ~x746 & ~x768;
assign c4426 = ~x8 & ~x48 & ~x49 & ~x76 & ~x135 & ~x252 & ~x282 & ~x361 & ~x388 & ~x389 & ~x478 & ~x507 & ~x532 & ~x535 & ~x615 & ~x690 & ~x691 & ~x708 & ~x710 & ~x711 & ~x712 & ~x713 & ~x716 & ~x718 & ~x719 & ~x737 & ~x739 & ~x740 & ~x741 & ~x742 & ~x744 & ~x746 & ~x758 & ~x764 & ~x768 & ~x769;
assign c4428 = ~x249 & ~x652 & ~x653 & ~x740;
assign c4430 =  x238 &  x298 &  x299 &  x467 &  x688 & ~x18 & ~x28 & ~x59 & ~x78 & ~x118 & ~x119 & ~x133 & ~x135 & ~x137 & ~x219 & ~x225 & ~x251 & ~x671 & ~x702 & ~x783;
assign c4432 =  x327 & ~x18 & ~x78 & ~x166 & ~x308 & ~x568 & ~x706 & ~x722 & ~x749;
assign c4434 = ~x232 & ~x348 & ~x768;
assign c4436 =  x585;
assign c4438 =  x427 &  x443 &  x494 &  x575 & ~x6 & ~x48 & ~x110 & ~x115 & ~x134 & ~x219 & ~x224 & ~x252 & ~x421 & ~x504 & ~x535 & ~x559 & ~x586 & ~x757;
assign c4440 = ~x198 & ~x244 & ~x472 & ~x505 & ~x768 & ~x769 & ~x773;
assign c4442 =  x14 &  x456 &  x484 &  x567 & ~x252 & ~x645 & ~x749;
assign c4444 =  x229 &  x257 &  x316 &  x325 &  x347 &  x377 &  x405 &  x412 &  x482 &  x514 &  x564 &  x638 &  x648 &  x732 &  x751 & ~x0 & ~x5 & ~x21 & ~x32 & ~x62 & ~x112 & ~x113 & ~x197 & ~x418 & ~x615 & ~x617 & ~x672 & ~x700 & ~x754 & ~x769 & ~x781;
assign c4446 =  x15 &  x484 & ~x364 & ~x710;
assign c4448 =  x235 &  x386 &  x554 &  x564 &  x581 &  x621 &  x624 &  x652 & ~x21 & ~x22 & ~x63 & ~x137 & ~x196 & ~x222 & ~x336 & ~x364 & ~x419 & ~x773 & ~x782;
assign c4450 = ~x272 & ~x348;
assign c4452 =  x43 &  x242 &  x271 &  x349 &  x372 &  x408 &  x492 &  x546 &  x602 &  x712 & ~x4 & ~x25 & ~x26 & ~x201 & ~x219 & ~x223 & ~x275 & ~x305 & ~x312 & ~x340 & ~x361 & ~x390 & ~x472 & ~x535 & ~x559 & ~x668 & ~x749 & ~x755 & ~x761 & ~x778;
assign c4454 =  x355 & ~x17 & ~x119 & ~x190 & ~x202 & ~x218 & ~x338 & ~x389 & ~x498 & ~x693;
assign c4456 = ~x208 & ~x421 & ~x737;
assign c4458 = ~x8 & ~x76 & ~x90 & ~x114 & ~x172 & ~x668 & ~x708 & ~x717 & ~x718 & ~x719 & ~x720 & ~x737 & ~x738 & ~x739 & ~x740 & ~x741 & ~x742 & ~x744 & ~x746 & ~x747;
assign c4460 =  x231 &  x294 &  x596 &  x623 &  x635 &  x651 &  x665 &  x742 &  x747 & ~x28 & ~x55 & ~x57 & ~x504;
assign c4462 =  x751 & ~x27 & ~x33 & ~x103;
assign c4464 =  x436 & ~x19 & ~x683 & ~x687 & ~x711 & ~x738;
assign c4466 = ~x172 & ~x477 & ~x502 & ~x580 & ~x708 & ~x709 & ~x710 & ~x711 & ~x718 & ~x719 & ~x727 & ~x737 & ~x738 & ~x739 & ~x740 & ~x741 & ~x742 & ~x745 & ~x747;
assign c4468 =  x238 &  x297 &  x344 &  x427 &  x604 &  x636 &  x692 & ~x27 & ~x32 & ~x58 & ~x118 & ~x134 & ~x171 & ~x172 & ~x194 & ~x219 & ~x251 & ~x394 & ~x504 & ~x726 & ~x758;
assign c4470 =  x243 &  x262 &  x326 &  x349 &  x440 &  x462 &  x577 & ~x35 & ~x36 & ~x54 & ~x113 & ~x219 & ~x247 & ~x256 & ~x280 & ~x445 & ~x530 & ~x615 & ~x644 & ~x645 & ~x668 & ~x679 & ~x696 & ~x763;
assign c4472 =  x692 &  x712 &  x720 & ~x19 & ~x91 & ~x586;
assign c4474 =  x289 &  x354 & ~x54 & ~x117 & ~x134 & ~x196 & ~x201 & ~x228 & ~x282 & ~x533 & ~x693 & ~x706 & ~x721;
assign c4476 =  x244 &  x267 &  x272 &  x295 &  x351 &  x357 &  x435 &  x484 &  x540 &  x608 &  x623 &  x637 &  x665 &  x679 &  x693 & ~x112 & ~x276 & ~x284 & ~x305 & ~x312 & ~x339 & ~x447 & ~x559 & ~x586 & ~x591 & ~x726 & ~x780;
assign c4478 = ~x18 & ~x21 & ~x31 & ~x35 & ~x36 & ~x49 & ~x63 & ~x226 & ~x284 & ~x472 & ~x499 & ~x530 & ~x534 & ~x558 & ~x640 & ~x701 & ~x720 & ~x737 & ~x738 & ~x739 & ~x740 & ~x745 & ~x746 & ~x747 & ~x768 & ~x773 & ~x780;
assign c4480 =  x331 &  x752 & ~x252 & ~x362 & ~x419 & ~x420 & ~x736 & ~x737 & ~x738;
assign c4482 =  x157 &  x325 &  x368 &  x396 &  x472 &  x492 &  x577 &  x584 & ~x7 & ~x22 & ~x56 & ~x61 & ~x112 & ~x115 & ~x249 & ~x306 & ~x419 & ~x559 & ~x589 & ~x615;
assign c4484 =  x350 & ~x25 & ~x28 & ~x61 & ~x64 & ~x119 & ~x133 & ~x134 & ~x219 & ~x247 & ~x279 & ~x363 & ~x503 & ~x735;
assign c4486 = ~x231 & ~x438 & ~x768;
assign c4488 = ~x16 & ~x90 & ~x172 & ~x301 & ~x359 & ~x391 & ~x393 & ~x534 & ~x719;
assign c4490 =  x259 &  x315 &  x400 &  x540 &  x568 &  x637 &  x638 &  x692 &  x693 &  x721 & ~x618;
assign c4492 =  x241 &  x322 & ~x10 & ~x46 & ~x64 & ~x133 & ~x162 & ~x172 & ~x190 & ~x246 & ~x285 & ~x303 & ~x340 & ~x615 & ~x757;
assign c4494 =  x12 &  x14 &  x15 &  x234 &  x238 &  x290 &  x322 &  x344 &  x481 &  x543 &  x648 & ~x8 & ~x19 & ~x26 & ~x57 & ~x78 & ~x88 & ~x142 & ~x277 & ~x362 & ~x420 & ~x531 & ~x699 & ~x771;
assign c4496 =  x154 &  x179 &  x184 &  x235 &  x265 &  x288 &  x313 &  x346 &  x408 &  x409 &  x493 &  x568 &  x594 &  x610 &  x631 &  x638 &  x653 & ~x2 & ~x3 & ~x26 & ~x30 & ~x33 & ~x36 & ~x57 & ~x61 & ~x87 & ~x137 & ~x163 & ~x165 & ~x192 & ~x226 & ~x227 & ~x249 & ~x477 & ~x559 & ~x613 & ~x616 & ~x641 & ~x674 & ~x697 & ~x727 & ~x758 & ~x768 & ~x771 & ~x781;
assign c4498 =  x751 & ~x30 & ~x34 & ~x56 & ~x57 & ~x76 & ~x78 & ~x79 & ~x254 & ~x276 & ~x304 & ~x333 & ~x394 & ~x419 & ~x449 & ~x531 & ~x559 & ~x614 & ~x643 & ~x669 & ~x699 & ~x720 & ~x736 & ~x737 & ~x738 & ~x740 & ~x741 & ~x745 & ~x746 & ~x747 & ~x767 & ~x768 & ~x780;
assign c41 = ~x72 & ~x97;
assign c43 =  x24 &  x419;
assign c45 =  x278;
assign c47 =  x193;
assign c49 = ~x384 & ~x496 & ~x566;
assign c411 = ~x182;
assign c413 =  x107;
assign c415 = ~x97 & ~x99;
assign c417 =  x766 & ~x425 & ~x565;
assign c419 = ~x545;
assign c421 =  x73 &  x91 &  x93 &  x96 &  x98 &  x102 &  x104 &  x157 &  x184 &  x260 &  x296 &  x358 &  x378 &  x466 &  x488 &  x520 &  x663 &  x666 &  x722 & ~x33 & ~x45 & ~x167 & ~x365 & ~x391 & ~x422 & ~x503 & ~x535 & ~x728 & ~x763;
assign c423 =  x19;
assign c425 =  x157 &  x264 &  x292 &  x660 & ~x314 & ~x398 & ~x666;
assign c427 =  x104 &  x706 & ~x39 & ~x760;
assign c429 = ~x126 & ~x155 & ~x236;
assign c431 =  x306;
assign c433 = ~x411 & ~x565 & ~x581 & ~x621;
assign c435 =  x615;
assign c437 = ~x455 & ~x524 & ~x567;
assign c439 =  x237 &  x291 & ~x425 & ~x426 & ~x525 & ~x609;
assign c441 =  x77 &  x135;
assign c443 =  x36 &  x62;
assign c445 =  x165;
assign c447 =  x7;
assign c449 =  x17;
assign c451 =  x17 &  x89;
assign c453 = ~x385 & ~x398;
assign c455 = ~x604;
assign c457 = ~x182 & ~x188;
assign c459 =  x137;
assign c461 = ~x258 & ~x413 & ~x483;
assign c463 =  x135;
assign c465 =  x2;
assign c467 =  x157 &  x184 &  x460 &  x463 &  x549 &  x660 &  x739 &  x740 & ~x7 & ~x107 & ~x109 & ~x254 & ~x336 & ~x364 & ~x443 & ~x448 & ~x509 & ~x537 & ~x560 & ~x565 & ~x566 & ~x587 & ~x610;
assign c469 =  x363;
assign c471 = ~x121 & ~x261 & ~x608 & ~x636 & ~x664;
assign c473 =  x76 &  x96 &  x133 &  x183 &  x509 &  x621 & ~x14;
assign c475 =  x72 &  x94 &  x96 &  x99 &  x104 &  x119 &  x125 &  x128 &  x161 &  x177 &  x185 &  x208 &  x258 &  x262 &  x273 &  x302 &  x414 &  x430 &  x432 &  x437 &  x459 &  x460 &  x471 &  x490 &  x491 &  x525 &  x526 &  x649 &  x661 &  x678 &  x705 &  x706 &  x722 &  x734 & ~x9 & ~x17 & ~x254 & ~x338 & ~x765 & ~x782;
assign c477 = ~x238;
assign c479 = ~x120 & ~x126;
assign c481 =  x67 &  x119 &  x463 &  x508 &  x677 & ~x13 & ~x389;
assign c483 = ~x122 & ~x374;
assign c485 =  x769 & ~x509 & ~x581;
assign c487 =  x107;
assign c489 =  x104 &  x189 &  x706 &  x770;
assign c491 = ~x313 & ~x373 & ~x398 & ~x565;
assign c493 =  x137;
assign c495 = ~x405 & ~x579 & ~x602;
assign c497 = ~x176;
assign c499 =  x755;
assign c4101 =  x94 &  x295 &  x543 &  x773 & ~x51 & ~x306 & ~x509 & ~x537 & ~x647 & ~x666;
assign c4103 = ~x157 & ~x491;
assign c4105 = ~x188 & ~x384;
assign c4107 = ~x125 & ~x182;
assign c4109 =  x40 &  x73 &  x74 &  x91 &  x93 &  x96 &  x105 &  x119 &  x125 &  x185 &  x296 &  x330 &  x350 &  x382 &  x397 &  x453 &  x462 &  x485 &  x494 &  x513 &  x523 &  x653 &  x659 &  x677 & ~x110 & ~x171 & ~x395 & ~x445 & ~x476 & ~x586 & ~x672 & ~x698;
assign c4111 =  x49;
assign c4113 =  x113 &  x225;
assign c4115 =  x18;
assign c4117 =  x18;
assign c4119 =  x280;
assign c4121 =  x17 &  x74 & ~x286 & ~x511;
assign c4123 =  x19;
assign c4125 =  x135 & ~x637;
assign c4127 =  x208 &  x237 & ~x341 & ~x398 & ~x470 & ~x510 & ~x610;
assign c4129 =  x106 & ~x511;
assign c4131 =  x78;
assign c4133 =  x63 &  x64 &  x90 &  x189 &  x480 & ~x13 & ~x389;
assign c4135 =  x135 & ~x314;
assign c4137 = ~x65 & ~x125;
assign c4139 = ~x495 & ~x602;
assign c4141 =  x362;
assign c4143 = ~x126;
assign c4145 = ~x125 & ~x235 & ~x236 & ~x237;
assign c4147 =  x773 & ~x386;
assign c4149 = ~x261;
assign c4151 =  x17 & ~x372 & ~x455;
assign c4153 = ~x547;
assign c4155 =  x88;
assign c4157 =  x78;
assign c4159 =  x503;
assign c4161 =  x26;
assign c4163 = ~x355 & ~x371;
assign c4165 =  x46 & ~x286;
assign c4167 = ~x97 & ~x98 & ~x266;
assign c4169 = ~x98;
assign c4171 =  x141;
assign c4173 = ~x120 & ~x126 & ~x155;
assign c4175 =  x711 & ~x356;
assign c4177 =  x476;
assign c4179 =  x418;
assign c4181 = ~x399 & ~x411;
assign c4183 =  x617;
assign c4185 =  x90 & ~x14;
assign c4187 =  x138 &  x643;
assign c4189 = ~x70 & ~x98 & ~x182;
assign c4191 =  x587;
assign c4193 = ~x327 & ~x483;
assign c4195 =  x96 &  x104 &  x376 &  x382 &  x566 &  x663 &  x745 & ~x38 & ~x277;
assign c4197 = ~x461 & ~x658 & ~x660 & ~x661;
assign c4199 =  x727;
assign c4201 =  x52;
assign c4203 =  x25;
assign c4205 =  x91 &  x96 &  x104 &  x161 &  x185 &  x206 &  x211 &  x217 &  x231 &  x246 &  x273 &  x285 &  x373 &  x399 &  x427 &  x460 &  x493 &  x522 &  x525 &  x526 &  x630 &  x677 &  x689 &  x722 & ~x164 & ~x170 & ~x194 & ~x276 & ~x309 & ~x417 & ~x418 & ~x420 & ~x757 & ~x775 & ~x777;
assign c4207 = ~x98;
assign c4209 = ~x430 & ~x573 & ~x621;
assign c4211 =  x309;
assign c4213 = ~x97 & ~x716;
assign c4215 =  x224;
assign c4217 = ~x122 & ~x126;
assign c4219 = ~x126;
assign c4221 =  x137;
assign c4223 = ~x16 & ~x125 & ~x182;
assign c4225 =  x93 &  x119 & ~x39 & ~x54 & ~x65;
assign c4227 =  x47 & ~x595;
assign c4229 =  x137;
assign c4231 =  x531 &  x561;
assign c4233 = ~x72 & ~x97 & ~x714;
assign c4235 = ~x147 & ~x373;
assign c4237 =  x560;
assign c4239 =  x532;
assign c4241 =  x645;
assign c4243 = ~x157;
assign c4245 =  x37 &  x64 &  x75 &  x76 &  x185 & ~x12 & ~x13;
assign c4247 = ~x69 & ~x125 & ~x153;
assign c4249 =  x292 &  x488 & ~x245 & ~x364 & ~x386 & ~x398 & ~x426 & ~x454 & ~x470 & ~x510 & ~x537 & ~x554 & ~x565 & ~x566 & ~x621 & ~x643;
assign c4251 =  x63 &  x76 &  x90 &  x104 &  x105 &  x118 &  x132 &  x183 & ~x770;
assign c4253 =  x643;
assign c4255 =  x51 &  x391;
assign c4257 =  x8;
assign c4259 = ~x126;
assign c4261 =  x112;
assign c4263 =  x68 &  x75 &  x96 &  x157 &  x520 & ~x12 & ~x15 & ~x61 & ~x196 & ~x643 & ~x727;
assign c4265 = ~x153 & ~x182;
assign c4267 = ~x330 & ~x345 & ~x425 & ~x527 & ~x611 & ~x621;
assign c4269 =  x115;
assign c4271 = ~x434;
assign c4273 =  x167;
assign c4275 =  x91 &  x94 &  x661 &  x722 & ~x38;
assign c4277 =  x68 &  x73 &  x91 &  x93 &  x96 &  x104 &  x159 &  x161 &  x203 &  x212 &  x294 &  x347 &  x358 &  x458 &  x513 &  x525 &  x565 &  x659 &  x663 &  x677 &  x722 & ~x504 & ~x506 & ~x559 & ~x562 & ~x588;
assign c4279 =  x212 &  x459 &  x488 &  x575 & ~x217 & ~x257 & ~x258 & ~x286 & ~x313;
assign c4281 =  x36 &  x64 &  x94 &  x272 &  x295 &  x326 &  x376 &  x680 &  x681 & ~x24 & ~x109 & ~x361 & ~x388 & ~x394;
assign c4283 =  x37 &  x117 &  x298 &  x685 & ~x389;
assign c4285 =  x197;
assign c4287 =  x774;
assign c4289 = ~x70 & ~x99;
assign c4291 =  x100 &  x488 &  x773 & ~x397 & ~x610;
assign c4293 = ~x125 & ~x236;
assign c4295 = ~x72;
assign c4297 =  x112;
assign c4299 = ~x372;
assign c4301 =  x76 &  x104 &  x258 &  x321 & ~x12 & ~x14 & ~x81 & ~x394 & ~x478;
assign c4303 =  x62;
assign c4305 =  x306;
assign c4307 = ~x42 & ~x71;
assign c4309 = ~x65;
assign c4311 =  x251;
assign c4313 = ~x370 & ~x440 & ~x608 & ~x609;
assign c4315 = ~x126;
assign c4317 = ~x122 & ~x573;
assign c4319 = ~x573;
assign c4321 =  x8;
assign c4323 = ~x237;
assign c4325 = ~x42 & ~x98;
assign c4327 =  x44 &  x68 &  x70 &  x73 &  x91 &  x94 &  x96 &  x104 &  x129 &  x132 &  x146 &  x157 &  x159 &  x161 &  x179 &  x185 &  x234 &  x271 &  x321 &  x325 &  x352 &  x403 &  x453 &  x458 &  x467 &  x481 &  x491 &  x497 &  x520 &  x526 &  x601 &  x602 &  x657 &  x677 &  x706 &  x722 & ~x84 & ~x110 & ~x193 & ~x250 & ~x305 & ~x530 & ~x585 & ~x670 & ~x675 & ~x753 & ~x759;
assign c4329 =  x37 &  x76 &  x90 &  x190 &  x382 &  x583 & ~x333 & ~x361;
assign c4331 =  x68 &  x96 &  x209 &  x492 &  x520 &  x660 & ~x337 & ~x483 & ~x511 & ~x776;
assign c4333 =  x64 &  x75 &  x94 &  x522 &  x600 & ~x12 & ~x15 & ~x89 & ~x107 & ~x193 & ~x362 & ~x366 & ~x417 & ~x423 & ~x473 & ~x504;
assign c4335 =  x390;
assign c4337 =  x40 &  x67 &  x73 &  x96 &  x104 &  x132 &  x160 &  x161 &  x203 &  x274 &  x329 &  x499 &  x520 &  x522 &  x573 &  x626 &  x687 &  x695 & ~x36 & ~x38 & ~x367;
assign c4339 =  x237 &  x683 &  x744 & ~x217 & ~x230 & ~x302 & ~x369 & ~x414 & ~x426 & ~x566 & ~x610 & ~x751;
assign c4341 =  x474;
assign c4343 = ~x148 & ~x239;
assign c4345 =  x128 &  x154 &  x321 & ~x161 & ~x338 & ~x358 & ~x387 & ~x414 & ~x425 & ~x565 & ~x704 & ~x762 & ~x779;
assign c4347 =  x6;
assign c4349 =  x76 &  x119 &  x132 &  x147 &  x161 &  x174 &  x183 &  x208 &  x214 &  x593 &  x649 & ~x14 & ~x311 & ~x558;
assign c4351 =  x197;
assign c4353 =  x77 &  x97 & ~x282;
assign c4355 = ~x635 & ~x658;
assign c4357 =  x418;
assign c4359 =  x194;
assign c4361 =  x560;
assign c4363 =  x278;
assign c4365 =  x78;
assign c4367 = ~x412 & ~x413 & ~x441 & ~x510 & ~x566 & ~x581;
assign c4369 = ~x153;
assign c4371 = ~x573;
assign c4373 =  x57;
assign c4375 =  x165;
assign c4377 =  x561;
assign c4379 =  x363;
assign c4381 =  x253;
assign c4383 = ~x373 & ~x621 & ~x778;
assign c4385 =  x101 &  x182 & ~x358 & ~x426 & ~x469 & ~x537 & ~x565 & ~x611;
assign c4387 =  x55 &  x112;
assign c4389 = ~x350 & ~x551;
assign c4391 =  x64 &  x76 &  x94 &  x97 &  x177 &  x185 &  x187 &  x565 &  x598 & ~x14 & ~x60 & ~x143 & ~x164 & ~x585 & ~x641 & ~x754;
assign c4393 =  x477;
assign c4395 =  x419;
assign c4397 = ~x65 & ~x242;
assign c4399 =  x10 &  x69 &  x70 &  x466 &  x600 & ~x558;
assign c4401 = ~x413 & ~x426 & ~x609 & ~x637;
assign c4403 = ~x154;
assign c4405 =  x75 &  x76 &  x90 &  x98 &  x105 &  x217 &  x245 &  x302 &  x346 &  x471 &  x481 &  x519 &  x527 &  x565 &  x625 & ~x394 & ~x534;
assign c4407 =  x142;
assign c4409 =  x86;
assign c4411 = ~x405 & ~x686;
assign c4413 =  x117 &  x688;
assign c4415 =  x166;
assign c4417 = ~x413 & ~x427;
assign c4419 =  x418;
assign c4421 =  x25;
assign c4423 = ~x242 & ~x630;
assign c4425 =  x458 &  x520 &  x599 & ~x342 & ~x358 & ~x470 & ~x566 & ~x621;
assign c4427 =  x28;
assign c4429 =  x71 &  x95 &  x129 &  x153 &  x264 &  x323 &  x432 &  x739 &  x740 &  x742 & ~x170 & ~x369 & ~x560 & ~x562 & ~x565 & ~x591 & ~x610 & ~x621 & ~x676;
assign c4431 = ~x72 & ~x126;
assign c4433 =  x335;
assign c4435 =  x81;
assign c4439 =  x392;
assign c4441 =  x363;
assign c4443 =  x278 &  x478;
assign c4445 = ~x126 & ~x153 & ~x182;
assign c4447 =  x21;
assign c4449 =  x363;
assign c4451 =  x210 &  x708 & ~x581;
assign c4453 =  x278;
assign c4457 = ~x42 & ~x97;
assign c4459 =  x51;
assign c4461 = ~x567 & ~x686;
assign c4463 =  x419;
assign c4465 =  x165;
assign c4467 = ~x120 & ~x125 & ~x182;
assign c4469 =  x10 &  x296 &  x660 & ~x7 & ~x58 & ~x279 & ~x472 & ~x505;
assign c4471 =  x46 & ~x442 & ~x482;
assign c4473 =  x56 & ~x371;
assign c4475 = ~x358 & ~x412 & ~x553 & ~x565;
assign c4477 =  x195;
assign c4479 =  x78;
assign c4481 = ~x372 & ~x427;
assign c4483 =  x107;
assign c4485 =  x109;
assign c4487 = ~x72;
assign c4489 = ~x270 & ~x286 & ~x621;
assign c4491 =  x222;
assign c4493 =  x196;
assign c4495 = ~x205 & ~x317 & ~x350;
assign c4497 =  x197;
assign c4499 =  x153 &  x287 &  x457 &  x655 &  x738 & ~x582 & ~x610 & ~x611 & ~x761;
assign c50 =  x220 &  x428 &  x567;
assign c52 =  x369 &  x436 & ~x1 & ~x43 & ~x46 & ~x47 & ~x102 & ~x119 & ~x148 & ~x156 & ~x336 & ~x622 & ~x634 & ~x636 & ~x681 & ~x686 & ~x697 & ~x708 & ~x716 & ~x720 & ~x733 & ~x751 & ~x767 & ~x777;
assign c54 =  x454 &  x513 & ~x403;
assign c56 =  x135;
assign c58 =  x651 &  x652 & ~x288 & ~x395 & ~x450;
assign c510 =  x481 & ~x240 & ~x548 & ~x569;
assign c512 =  x481 & ~x36 & ~x44 & ~x78 & ~x86 & ~x103 & ~x190 & ~x192 & ~x234 & ~x241 & ~x283 & ~x285 & ~x447 & ~x574 & ~x649 & ~x728;
assign c514 =  x436 &  x454 &  x483 & ~x45 & ~x111 & ~x118 & ~x159 & ~x186 & ~x270 & ~x692 & ~x699 & ~x709 & ~x722 & ~x748;
assign c516 =  x265 & ~x8 & ~x89 & ~x152 & ~x185 & ~x202 & ~x204 & ~x213 & ~x243 & ~x259 & ~x282 & ~x311 & ~x312 & ~x676 & ~x697 & ~x703 & ~x711 & ~x712;
assign c518 =  x512 &  x514 & ~x569 & ~x689;
assign c520 =  x398 &  x505 &  x569;
assign c522 =  x426 &  x451 &  x454 & ~x16 & ~x269 & ~x270 & ~x306 & ~x313 & ~x604 & ~x694;
assign c524 =  x342;
assign c526 =  x218 & ~x354 & ~x535;
assign c528 =  x613 & ~x607 & ~x722;
assign c530 =  x538 &  x567 & ~x347;
assign c532 =  x538 &  x539 & ~x186 & ~x258 & ~x288 & ~x423 & ~x477 & ~x740 & ~x743;
assign c534 = ~x326 & ~x518 & ~x540 & ~x541 & ~x542 & ~x546 & ~x569;
assign c536 =  x427 &  x537 &  x569 &  x571 & ~x53 & ~x664;
assign c538 =  x454 &  x482 &  x534 &  x540 &  x568 & ~x46 & ~x114 & ~x145 & ~x180 & ~x636 & ~x692 & ~x716;
assign c540 =  x325 &  x355 & ~x76 & ~x373 & ~x435 & ~x450;
assign c542 = ~x13 & ~x42 & ~x129 & ~x166 & ~x180 & ~x257 & ~x284 & ~x293 & ~x391 & ~x450 & ~x459 & ~x589 & ~x645 & ~x698 & ~x705 & ~x776;
assign c544 =  x481 &  x509 & ~x315 & ~x460;
assign c546 =  x158 & ~x450 & ~x477 & ~x478 & ~x506;
assign c548 =  x399 &  x480 &  x481 & ~x107 & ~x346 & ~x447 & ~x579 & ~x630 & ~x650 & ~x663 & ~x740 & ~x742 & ~x744;
assign c550 =  x454 & ~x269 & ~x270 & ~x570;
assign c552 =  x266 &  x398 &  x509 & ~x391 & ~x736;
assign c554 =  x453 & ~x269 & ~x539 & ~x543 & ~x548 & ~x552 & ~x578;
assign c556 =  x386 &  x413 & ~x24 & ~x88 & ~x285 & ~x313 & ~x405 & ~x433 & ~x434 & ~x478;
assign c558 =  x539 &  x567 &  x572 & ~x73 & ~x128 & ~x532 & ~x722;
assign c560 = ~x40 & ~x77 & ~x102 & ~x137 & ~x295 & ~x325 & ~x326 & ~x447 & ~x531 & ~x588 & ~x633 & ~x666 & ~x692 & ~x700 & ~x706 & ~x711 & ~x777;
assign c562 =  x398 &  x536 &  x539 &  x569 & ~x281;
assign c564 =  x103 &  x713;
assign c566 =  x595 &  x613 & ~x154 & ~x450 & ~x451 & ~x616;
assign c568 =  x521 & ~x377 & ~x378;
assign c570 =  x76;
assign c572 =  x667 & ~x477 & ~x480;
assign c574 =  x736 & ~x456;
assign c576 =  x679 & ~x509;
assign c578 =  x604 & ~x508 & ~x514 & ~x559;
assign c580 =  x162;
assign c582 = ~x184 & ~x386 & ~x389 & ~x594 & ~x596 & ~x715;
assign c584 =  x397 &  x481 &  x541 & ~x185 & ~x578;
assign c586 =  x266 &  x481 & ~x596;
assign c588 =  x428 & ~x143 & ~x241 & ~x269 & ~x575 & ~x621 & ~x638 & ~x643 & ~x675 & ~x686 & ~x698;
assign c590 =  x426 & ~x16 & ~x96 & ~x116 & ~x269 & ~x447 & ~x562 & ~x565 & ~x574 & ~x575 & ~x580 & ~x588 & ~x700 & ~x708 & ~x711 & ~x728 & ~x748 & ~x769 & ~x770 & ~x777;
assign c592 =  x266 &  x481 & ~x102 & ~x103 & ~x241 & ~x242 & ~x281 & ~x691 & ~x703;
assign c594 =  x524 & ~x406 & ~x407;
assign c596 = ~x85 & ~x98 & ~x149 & ~x174 & ~x215 & ~x287 & ~x291 & ~x413 & ~x477 & ~x478 & ~x480 & ~x739;
assign c598 =  x531;
assign c5100 =  x623 &  x641 & ~x71 & ~x340 & ~x477;
assign c5102 =  x537 & ~x14 & ~x138 & ~x154 & ~x391 & ~x478 & ~x506;
assign c5104 =  x425 &  x537 &  x540 &  x567 & ~x650;
assign c5106 =  x426 &  x481 & ~x177 & ~x269 & ~x270 & ~x656 & ~x657 & ~x686 & ~x743;
assign c5108 =  x219 &  x538;
assign c5110 =  x159 & ~x450 & ~x477 & ~x646;
assign c5112 =  x565 & ~x295 & ~x326;
assign c5114 =  x239 & ~x33 & ~x258;
assign c5116 =  x509 &  x537 &  x539 & ~x399 & ~x477 & ~x531 & ~x749;
assign c5118 = ~x65 & ~x181 & ~x186 & ~x202 & ~x221 & ~x241 & ~x388 & ~x504 & ~x561 & ~x569 & ~x572 & ~x574 & ~x578 & ~x582 & ~x627 & ~x650 & ~x663 & ~x665 & ~x675 & ~x724 & ~x738;
assign c5120 =  x565 &  x581 & ~x506;
assign c5122 =  x299 & ~x124 & ~x323 & ~x531 & ~x761;
assign c5124 =  x713 & ~x540;
assign c5126 = ~x8 & ~x16 & ~x26 & ~x70 & ~x74 & ~x89 & ~x106 & ~x149 & ~x159 & ~x162 & ~x180 & ~x255 & ~x282 & ~x356 & ~x363 & ~x477 & ~x504 & ~x559 & ~x688 & ~x692 & ~x698 & ~x717 & ~x746;
assign c5128 =  x595 &  x596 &  x611 & ~x739 & ~x740;
assign c5130 =  x641 & ~x579;
assign c5132 = ~x18 & ~x81 & ~x149 & ~x166 & ~x206 & ~x360 & ~x362 & ~x477 & ~x506 & ~x579 & ~x588 & ~x720 & ~x729 & ~x753;
assign c5134 = ~x69 & ~x124 & ~x163 & ~x176 & ~x181 & ~x193 & ~x349 & ~x377 & ~x661 & ~x664;
assign c5136 =  x481 & ~x197 & ~x242 & ~x364 & ~x561 & ~x565 & ~x568 & ~x569 & ~x573 & ~x575 & ~x634 & ~x685 & ~x686 & ~x721 & ~x742;
assign c5138 = ~x12 & ~x36 & ~x38 & ~x40 & ~x150 & ~x204 & ~x253 & ~x256 & ~x286 & ~x309 & ~x378 & ~x406 & ~x407 & ~x435;
assign c5140 = ~x44 & ~x55 & ~x69 & ~x70 & ~x98 & ~x150 & ~x232 & ~x258 & ~x356 & ~x373 & ~x478 & ~x688 & ~x767 & ~x774;
assign c5142 =  x613 &  x641 & ~x154 & ~x506;
assign c5144 =  x165 & ~x19;
assign c5146 = ~x11 & ~x40 & ~x69 & ~x74 & ~x77 & ~x97 & ~x113 & ~x118 & ~x122 & ~x151 & ~x162 & ~x166 & ~x236 & ~x241 & ~x285 & ~x291 & ~x310 & ~x445 & ~x563 & ~x575 & ~x609 & ~x611 & ~x655 & ~x675 & ~x699 & ~x715 & ~x745 & ~x754 & ~x779;
assign c5148 =  x730;
assign c5150 =  x357 & ~x128 & ~x349 & ~x434 & ~x435;
assign c5152 = ~x25 & ~x67 & ~x114 & ~x121 & ~x151 & ~x174 & ~x325 & ~x508 & ~x543 & ~x688 & ~x722 & ~x733;
assign c5154 =  x538 &  x566 & ~x70 & ~x231 & ~x235 & ~x343 & ~x366 & ~x478 & ~x671 & ~x674 & ~x739;
assign c5156 =  x566 & ~x99 & ~x166 & ~x202 & ~x321 & ~x478;
assign c5158 =  x534 &  x539 & ~x233 & ~x341 & ~x639;
assign c5160 = ~x14 & ~x37 & ~x38 & ~x48 & ~x77 & ~x102 & ~x111 & ~x124 & ~x125 & ~x129 & ~x132 & ~x150 & ~x172 & ~x208 & ~x221 & ~x241 & ~x417 & ~x447 & ~x563 & ~x565 & ~x567 & ~x577 & ~x579 & ~x599 & ~x647 & ~x652 & ~x666 & ~x720 & ~x740;
assign c5162 =  x299 &  x300 & ~x14 & ~x18 & ~x45 & ~x79 & ~x115 & ~x144 & ~x149 & ~x152 & ~x154 & ~x179 & ~x197 & ~x199 & ~x204 & ~x232 & ~x280 & ~x281 & ~x286 & ~x313 & ~x316 & ~x357 & ~x364 & ~x711 & ~x719 & ~x721 & ~x723 & ~x739 & ~x750 & ~x758 & ~x771 & ~x779;
assign c5164 = ~x15 & ~x19 & ~x70 & ~x72 & ~x75 & ~x82 & ~x86 & ~x113 & ~x125 & ~x147 & ~x149 & ~x153 & ~x392 & ~x405 & ~x406 & ~x433 & ~x434 & ~x717;
assign c5166 = ~x208 & ~x268 & ~x270 & ~x508 & ~x518 & ~x539 & ~x550 & ~x571 & ~x581 & ~x672;
assign c5168 =  x537 &  x539 &  x540 & ~x351;
assign c5170 =  x567 & ~x407;
assign c5172 =  x481 &  x567 &  x568 &  x569 & ~x120 & ~x166 & ~x187 & ~x261 & ~x637;
assign c5174 = ~x121 & ~x149 & ~x227 & ~x344 & ~x391 & ~x392 & ~x403 & ~x447 & ~x509 & ~x525 & ~x552 & ~x671 & ~x759;
assign c5176 =  x533 & ~x447;
assign c5178 =  x533 &  x539;
assign c5180 = ~x362 & ~x507 & ~x541 & ~x546 & ~x547 & ~x552 & ~x570 & ~x574 & ~x578 & ~x579 & ~x580 & ~x655 & ~x685 & ~x762 & ~x777;
assign c5182 =  x76 &  x681 & ~x563;
assign c5184 =  x306;
assign c5186 =  x431 &  x482 & ~x70 & ~x71 & ~x213 & ~x447 & ~x579;
assign c5188 =  x134 &  x684;
assign c5190 = ~x150 & ~x162 & ~x182 & ~x234 & ~x269 & ~x567 & ~x604 & ~x606 & ~x646;
assign c5192 =  x603 & ~x323;
assign c5194 = ~x60 & ~x104 & ~x105 & ~x241 & ~x416 & ~x567 & ~x578 & ~x579 & ~x582 & ~x609 & ~x666 & ~x674 & ~x676 & ~x685 & ~x688 & ~x703 & ~x741 & ~x745;
assign c5196 =  x468 &  x482 & ~x4 & ~x65 & ~x70 & ~x151 & ~x159 & ~x171 & ~x350 & ~x364 & ~x394 & ~x676 & ~x686 & ~x693;
assign c5198 =  x767 & ~x458 & ~x479;
assign c5200 =  x218 &  x594 & ~x751;
assign c5202 =  x595 & ~x152 & ~x157 & ~x303;
assign c5204 =  x238;
assign c5206 =  x369 & ~x185;
assign c5208 = ~x68 & ~x187 & ~x284 & ~x314 & ~x349 & ~x378 & ~x407 & ~x656 & ~x707 & ~x747;
assign c5210 =  x509 &  x551 & ~x186 & ~x240 & ~x681 & ~x770;
assign c5212 = ~x341 & ~x395 & ~x509 & ~x552;
assign c5214 =  x524 & ~x4 & ~x45 & ~x166 & ~x176 & ~x281 & ~x291 & ~x407 & ~x745;
assign c5216 =  x162;
assign c5218 =  x359 &  x448 &  x539 &  x543 & ~x111;
assign c5220 =  x430 &  x454 & ~x30 & ~x73 & ~x116 & ~x269 & ~x310 & ~x362 & ~x419 & ~x657 & ~x712;
assign c5222 =  x267 &  x540 & ~x345 & ~x368;
assign c5224 =  x735;
assign c5226 =  x239 & ~x379;
assign c5228 =  x484 & ~x318 & ~x418 & ~x575;
assign c5230 =  x399 & ~x98 & ~x107 & ~x154 & ~x187 & ~x349 & ~x715;
assign c5232 =  x481 &  x539 &  x569 & ~x91 & ~x242;
assign c5234 =  x425 & ~x100 & ~x159 & ~x269 & ~x270 & ~x507 & ~x539 & ~x540 & ~x543 & ~x546 & ~x547 & ~x548 & ~x550 & ~x552 & ~x554 & ~x556 & ~x565 & ~x609 & ~x650 & ~x658 & ~x704 & ~x771;
assign c5236 = ~x523 & ~x537 & ~x539 & ~x542 & ~x546 & ~x550 & ~x572 & ~x582 & ~x728;
assign c5238 =  x481 & ~x112 & ~x128 & ~x135 & ~x269 & ~x270 & ~x562 & ~x565 & ~x581 & ~x630 & ~x668 & ~x705 & ~x719 & ~x762;
assign c5240 =  x434 & ~x62 & ~x119 & ~x174 & ~x175 & ~x289 & ~x363 & ~x386 & ~x389 & ~x532 & ~x622 & ~x756;
assign c5242 = ~x14 & ~x18 & ~x39 & ~x70 & ~x71 & ~x85 & ~x149 & ~x198 & ~x255 & ~x258 & ~x280 & ~x281 & ~x312 & ~x313 & ~x422 & ~x506 & ~x523 & ~x537 & ~x538 & ~x551 & ~x552 & ~x714 & ~x717;
assign c5244 = ~x23 & ~x24 & ~x129 & ~x325 & ~x388 & ~x520 & ~x577 & ~x650 & ~x694 & ~x706 & ~x711 & ~x729 & ~x733;
assign c5246 =  x425 & ~x359 & ~x540 & ~x546;
assign c5248 =  x451 & ~x508 & ~x579;
assign c5250 =  x134;
assign c5252 = ~x40 & ~x269 & ~x390 & ~x505 & ~x508 & ~x539 & ~x711 & ~x733;
assign c5254 =  x510 & ~x13 & ~x22 & ~x39 & ~x45 & ~x62 & ~x73 & ~x84 & ~x147 & ~x156 & ~x170 & ~x177 & ~x204 & ~x205 & ~x208 & ~x240 & ~x285 & ~x345 & ~x447 & ~x587 & ~x617 & ~x653 & ~x688 & ~x742 & ~x750;
assign c5256 =  x681 & ~x509 & ~x619;
assign c5258 =  x732;
assign c5260 =  x48;
assign c5262 =  x238 &  x239 &  x508 &  x512 & ~x214;
assign c5264 =  x557 & ~x356 & ~x424;
assign c5266 =  x427 &  x481 & ~x43 & ~x63 & ~x349 & ~x606 & ~x631 & ~x671 & ~x703;
assign c5268 =  x371 &  x481 & ~x149 & ~x337;
assign c5270 =  x425 &  x453 & ~x10 & ~x111 & ~x164 & ~x182 & ~x185 & ~x186 & ~x212 & ~x240 & ~x254 & ~x270 & ~x570 & ~x575 & ~x638;
assign c5272 =  x239 &  x538 & ~x158 & ~x405;
assign c5274 =  x701;
assign c5276 =  x397 &  x502 & ~x309 & ~x578 & ~x675 & ~x759;
assign c5278 = ~x298 & ~x518 & ~x523 & ~x537 & ~x539 & ~x542 & ~x565;
assign c5280 =  x477 &  x537 &  x541 & ~x215;
assign c5282 =  x565 & ~x232 & ~x517 & ~x709;
assign c5284 = ~x42 & ~x54 & ~x325 & ~x475 & ~x537 & ~x540 & ~x546 & ~x616 & ~x638;
assign c5286 =  x359 & ~x4 & ~x69 & ~x321 & ~x433 & ~x434;
assign c5288 =  x373 &  x477 &  x480 &  x507 &  x538 &  x541 & ~x223 & ~x607 & ~x717 & ~x722;
assign c5290 =  x76 & ~x454;
assign c5292 =  x453 & ~x46 & ~x403;
assign c5294 =  x218 & ~x1 & ~x8 & ~x14 & ~x15 & ~x16 & ~x19 & ~x24 & ~x41 & ~x47 & ~x60 & ~x63 & ~x65 & ~x66 & ~x76 & ~x78 & ~x97 & ~x105 & ~x142 & ~x144 & ~x154 & ~x159 & ~x168 & ~x174 & ~x176 & ~x177 & ~x179 & ~x181 & ~x186 & ~x204 & ~x222 & ~x235 & ~x263 & ~x287 & ~x309 & ~x341 & ~x364 & ~x532 & ~x615 & ~x634 & ~x643 & ~x661 & ~x672 & ~x680 & ~x682 & ~x683 & ~x687 & ~x691 & ~x704 & ~x706 & ~x720 & ~x722 & ~x725 & ~x728 & ~x738 & ~x741 & ~x742 & ~x743 & ~x745 & ~x748 & ~x774 & ~x782;
assign c5296 =  x481 & ~x128 & ~x447 & ~x554 & ~x582;
assign c5298 =  x398 &  x509 &  x538 & ~x339;
assign c5300 =  x539 & ~x350 & ~x689;
assign c5302 =  x220 & ~x326;
assign c5304 =  x264 &  x428;
assign c5306 =  x415 & ~x65 & ~x123 & ~x406 & ~x435;
assign c5308 =  x539 & ~x129 & ~x283;
assign c5310 =  x537 &  x540 & ~x177 & ~x232 & ~x269 & ~x337 & ~x587 & ~x697 & ~x765;
assign c5312 =  x454 & ~x520 & ~x539 & ~x542;
assign c5314 = ~x5 & ~x184 & ~x233 & ~x240 & ~x548 & ~x550 & ~x580 & ~x616 & ~x631;
assign c5316 =  x278 & ~x379;
assign c5318 =  x276 &  x509 &  x514 &  x515 & ~x230 & ~x234 & ~x318 & ~x345 & ~x469 & ~x705;
assign c5320 =  x484 & ~x154 & ~x240 & ~x447 & ~x564 & ~x582 & ~x587;
assign c5322 =  x106;
assign c5324 =  x454 & ~x112 & ~x152 & ~x166 & ~x180 & ~x215 & ~x241 & ~x263 & ~x447 & ~x548 & ~x569 & ~x572 & ~x636 & ~x638 & ~x646 & ~x708 & ~x714 & ~x720 & ~x748 & ~x766 & ~x771;
assign c5326 =  x536 &  x537 &  x539 & ~x138 & ~x366 & ~x565 & ~x611 & ~x666 & ~x712 & ~x722 & ~x735 & ~x771 & ~x780;
assign c5328 =  x537;
assign c5330 =  x480 &  x527 &  x538 &  x540 & ~x42 & ~x99 & ~x125 & ~x180 & ~x199 & ~x254 & ~x289 & ~x559 & ~x616 & ~x741;
assign c5332 =  x266 & ~x13 & ~x14 & ~x61 & ~x82 & ~x96 & ~x108 & ~x204 & ~x254 & ~x312 & ~x315 & ~x336 & ~x339 & ~x378 & ~x393 & ~x587 & ~x699 & ~x758;
assign c5334 =  x264 & ~x70 & ~x202 & ~x283 & ~x309 & ~x629 & ~x646 & ~x673 & ~x719;
assign c5336 =  x468 &  x533 &  x534 & ~x422;
assign c5338 =  x510 &  x539 & ~x447 & ~x548;
assign c5340 =  x369 & ~x4 & ~x74 & ~x145 & ~x556 & ~x646 & ~x674 & ~x678 & ~x704 & ~x715 & ~x766 & ~x770;
assign c5342 =  x451 & ~x74 & ~x270 & ~x507 & ~x541 & ~x546 & ~x552 & ~x554 & ~x570 & ~x579;
assign c5344 =  x679 & ~x511;
assign c5346 =  x334 &  x624 & ~x258;
assign c5348 =  x537 &  x541 &  x567 &  x568 & ~x608 & ~x767 & ~x771;
assign c5350 = ~x24 & ~x33 & ~x79 & ~x134 & ~x136 & ~x145 & ~x200 & ~x263 & ~x395 & ~x477 & ~x478 & ~x531 & ~x560 & ~x575 & ~x578 & ~x579 & ~x627 & ~x643 & ~x655 & ~x658 & ~x680 & ~x685 & ~x720 & ~x742 & ~x747 & ~x752;
assign c5352 =  x731;
assign c5354 = ~x233 & ~x323 & ~x480 & ~x506 & ~x509 & ~x511 & ~x527 & ~x537;
assign c5356 =  x482 & ~x121 & ~x243 & ~x269 & ~x534 & ~x570 & ~x574;
assign c5358 = ~x356 & ~x403 & ~x538 & ~x540 & ~x542;
assign c5360 =  x569 & ~x55 & ~x62 & ~x69 & ~x102 & ~x115 & ~x179 & ~x197 & ~x237 & ~x575 & ~x622 & ~x626 & ~x627 & ~x712 & ~x727 & ~x734 & ~x751 & ~x756;
assign c5362 =  x733;
assign c5364 =  x398 &  x477 &  x507;
assign c5366 = ~x102 & ~x269 & ~x368 & ~x476 & ~x531 & ~x569 & ~x654 & ~x716;
assign c5368 =  x509 &  x592 & ~x47 & ~x127 & ~x376 & ~x658;
assign c5370 =  x264 & ~x36 & ~x65 & ~x83 & ~x98 & ~x180 & ~x283 & ~x340 & ~x766;
assign c5372 =  x622 & ~x315 & ~x345 & ~x400 & ~x563 & ~x615;
assign c5374 =  x537 &  x538 & ~x179 & ~x459 & ~x715;
assign c5376 =  x565 & ~x477 & ~x507;
assign c5378 = ~x3 & ~x4 & ~x14 & ~x18 & ~x49 & ~x55 & ~x68 & ~x81 & ~x90 & ~x262 & ~x312 & ~x409 & ~x422 & ~x447 & ~x450 & ~x478 & ~x503 & ~x590 & ~x691 & ~x700 & ~x742 & ~x745 & ~x755;
assign c5380 =  x106;
assign c5382 =  x507 & ~x269 & ~x418;
assign c5384 =  x669 & ~x722;
assign c5386 =  x595 &  x613 & ~x181 & ~x450 & ~x478 & ~x533;
assign c5388 =  x370 &  x454 & ~x179 & ~x291 & ~x318 & ~x666 & ~x703 & ~x741;
assign c5390 = ~x321 & ~x433 & ~x435 & ~x480;
assign c5392 =  x621;
assign c5394 =  x540 & ~x3 & ~x117 & ~x262 & ~x422 & ~x424 & ~x480;
assign c5396 = ~x39 & ~x355 & ~x356 & ~x477 & ~x542;
assign c5398 = ~x14 & ~x18 & ~x64 & ~x118 & ~x179 & ~x198 & ~x322 & ~x478 & ~x506 & ~x536 & ~x539 & ~x540 & ~x541 & ~x542 & ~x636 & ~x703 & ~x705;
assign c5400 =  x264;
assign c5402 = ~x236 & ~x269 & ~x287 & ~x417 & ~x575 & ~x577 & ~x620 & ~x649 & ~x652 & ~x660;
assign c5404 =  x78;
assign c5406 =  x549 & ~x185 & ~x317 & ~x613 & ~x734;
assign c5408 = ~x240 & ~x241 & ~x388 & ~x551 & ~x596 & ~x657;
assign c5410 =  x406 & ~x65 & ~x71 & ~x111 & ~x176 & ~x204 & ~x228 & ~x441 & ~x506 & ~x508 & ~x533;
assign c5412 =  x164;
assign c5414 =  x384 & ~x379 & ~x447 & ~x661 & ~x691 & ~x764 & ~x768;
assign c5416 =  x631 & ~x371 & ~x406 & ~x435;
assign c5420 =  x539 & ~x97 & ~x514;
assign c5422 = ~x96 & ~x113 & ~x259 & ~x260 & ~x368 & ~x378 & ~x406 & ~x407;
assign c5424 = ~x67 & ~x89 & ~x129 & ~x130 & ~x149 & ~x313 & ~x368 & ~x478 & ~x507 & ~x508 & ~x525 & ~x531 & ~x533 & ~x552 & ~x562 & ~x580 & ~x590 & ~x617 & ~x720;
assign c5426 =  x582 & ~x257 & ~x347 & ~x374 & ~x506;
assign c5428 =  x239 &  x481 &  x539;
assign c5430 =  x539 & ~x98 & ~x433;
assign c5432 =  x476 &  x536 &  x568;
assign c5434 =  x189 &  x621 &  x622;
assign c5436 =  x454 & ~x18 & ~x78 & ~x179 & ~x185 & ~x240 & ~x241 & ~x242 & ~x270 & ~x565 & ~x571 & ~x572 & ~x574 & ~x577 & ~x578 & ~x582 & ~x596 & ~x606 & ~x652 & ~x691 & ~x731;
assign c5438 =  x264 &  x266 & ~x288;
assign c5440 =  x503;
assign c5442 =  x237 & ~x126 & ~x532 & ~x676;
assign c5444 =  x483 &  x537 &  x538 & ~x69 & ~x128 & ~x285 & ~x343 & ~x422 & ~x506;
assign c5446 =  x509 & ~x101 & ~x119 & ~x534 & ~x568 & ~x569 & ~x577 & ~x649 & ~x740 & ~x746;
assign c5448 = ~x2 & ~x4 & ~x5 & ~x14 & ~x55 & ~x66 & ~x74 & ~x88 & ~x95 & ~x122 & ~x128 & ~x156 & ~x166 & ~x168 & ~x180 & ~x185 & ~x187 & ~x191 & ~x208 & ~x213 & ~x236 & ~x282 & ~x308 & ~x318 & ~x363 & ~x364 & ~x395 & ~x396 & ~x418 & ~x578 & ~x617 & ~x623 & ~x639 & ~x659 & ~x662 & ~x667 & ~x689 & ~x714 & ~x722 & ~x733 & ~x738 & ~x740 & ~x768;
assign c5450 =  x681 & ~x513;
assign c5452 =  x679 & ~x174 & ~x287 & ~x552 & ~x694;
assign c5454 =  x450 & ~x268 & ~x548;
assign c5456 =  x603 & ~x459 & ~x508 & ~x530 & ~x590;
assign c5458 =  x265 &  x512 & ~x319 & ~x716;
assign c5460 =  x162 &  x677;
assign c5462 =  x211 & ~x350;
assign c5464 =  x451 & ~x270 & ~x534 & ~x539 & ~x540 & ~x542 & ~x550;
assign c5466 =  x509 & ~x127 & ~x259 & ~x416 & ~x607 & ~x741 & ~x745;
assign c5468 =  x105;
assign c5470 = ~x14 & ~x45 & ~x118 & ~x128 & ~x152 & ~x305 & ~x309 & ~x323 & ~x706 & ~x722 & ~x736 & ~x738 & ~x740 & ~x745;
assign c5472 =  x102 &  x712;
assign c5474 =  x393 &  x397 & ~x577;
assign c5476 =  x739;
assign c5478 =  x237 & ~x97 & ~x149 & ~x725;
assign c5480 = ~x10 & ~x108 & ~x115 & ~x116 & ~x224 & ~x234 & ~x412 & ~x422 & ~x423 & ~x504 & ~x506 & ~x508 & ~x729 & ~x761 & ~x780;
assign c5482 =  x567 & ~x64 & ~x78 & ~x94 & ~x114 & ~x127 & ~x128 & ~x144 & ~x178 & ~x223 & ~x372 & ~x477 & ~x480 & ~x506 & ~x507 & ~x716 & ~x719 & ~x742 & ~x764 & ~x766;
assign c5484 =  x509 &  x512 &  x566 &  x567 & ~x61 & ~x177 & ~x233 & ~x263 & ~x290 & ~x314 & ~x337 & ~x708 & ~x712 & ~x736;
assign c5486 =  x358 &  x454 & ~x7 & ~x118 & ~x123 & ~x125 & ~x137 & ~x221 & ~x241 & ~x570 & ~x573 & ~x575 & ~x577 & ~x654 & ~x715 & ~x733 & ~x747;
assign c5488 =  x239 & ~x540 & ~x711;
assign c5490 =  x407 & ~x8 & ~x14 & ~x32 & ~x45 & ~x59 & ~x63 & ~x70 & ~x100 & ~x103 & ~x106 & ~x116 & ~x117 & ~x145 & ~x149 & ~x173 & ~x195 & ~x197 & ~x200 & ~x204 & ~x205 & ~x229 & ~x230 & ~x257 & ~x261 & ~x283 & ~x313 & ~x335 & ~x357 & ~x391 & ~x450 & ~x588 & ~x617 & ~x643 & ~x664 & ~x676 & ~x686 & ~x689 & ~x692 & ~x706 & ~x744 & ~x769;
assign c5492 =  x505 &  x506 &  x507;
assign c5494 = ~x28 & ~x40 & ~x87 & ~x97 & ~x111 & ~x229 & ~x233 & ~x288 & ~x378 & ~x407 & ~x480 & ~x716 & ~x745;
assign c5496 =  x162 &  x603;
assign c5498 =  x631 &  x708 & ~x372 & ~x538;
assign c51 =  x295 &  x349 &  x351 &  x354 &  x382 &  x387 &  x418 &  x443 &  x474 &  x491 &  x509 & ~x29 & ~x51 & ~x77 & ~x111 & ~x136 & ~x158 & ~x165 & ~x246 & ~x641 & ~x662 & ~x733;
assign c53 =  x353 &  x361 &  x439 &  x443 &  x445 &  x473 &  x474 & ~x35 & ~x53 & ~x77 & ~x104 & ~x109 & ~x110 & ~x130 & ~x132 & ~x145 & ~x148 & ~x162 & ~x163 & ~x165 & ~x166 & ~x170 & ~x189 & ~x191 & ~x192 & ~x207 & ~x213 & ~x218 & ~x220 & ~x222 & ~x265 & ~x592 & ~x599 & ~x612 & ~x645 & ~x650 & ~x695 & ~x708 & ~x723 & ~x763;
assign c55 = ~x18 & ~x51 & ~x104 & ~x191 & ~x217 & ~x274 & ~x314 & ~x329 & ~x450 & ~x478 & ~x482 & ~x498 & ~x499 & ~x500 & ~x501 & ~x529 & ~x565 & ~x585 & ~x647 & ~x675 & ~x697 & ~x755 & ~x766 & ~x777;
assign c57 =  x193 &  x521 &  x590;
assign c59 = ~x26 & ~x59 & ~x83 & ~x84 & ~x175 & ~x207 & ~x272 & ~x273 & ~x301 & ~x494 & ~x495 & ~x498 & ~x501 & ~x557 & ~x675 & ~x679;
assign c511 =  x68 & ~x501;
assign c513 =  x214 &  x245 &  x275 &  x384 &  x474 & ~x397 & ~x398;
assign c515 =  x258;
assign c517 =  x646;
assign c519 = ~x247 & ~x382 & ~x472 & ~x501 & ~x528 & ~x696;
assign c521 =  x244 &  x277 &  x351 &  x411 & ~x397;
assign c523 =  x91;
assign c525 =  x15;
assign c527 =  x387 &  x413 &  x443 & ~x112 & ~x148 & ~x159 & ~x170 & ~x199 & ~x217 & ~x226 & ~x236 & ~x247 & ~x262 & ~x273 & ~x299 & ~x301 & ~x328 & ~x617 & ~x636 & ~x755 & ~x757;
assign c529 =  x204;
assign c531 =  x742;
assign c533 =  x349 &  x351 &  x377 &  x379 &  x385 &  x390 &  x417 &  x441 &  x443 &  x469 &  x497 & ~x0 & ~x67 & ~x76 & ~x77 & ~x86 & ~x109 & ~x110 & ~x117 & ~x123 & ~x125 & ~x145 & ~x154 & ~x155 & ~x226 & ~x227 & ~x234 & ~x243 & ~x245 & ~x262 & ~x342 & ~x589 & ~x605 & ~x686 & ~x688 & ~x694 & ~x718 & ~x720 & ~x727 & ~x736 & ~x743 & ~x761 & ~x779;
assign c535 =  x717;
assign c537 =  x323 &  x347 &  x349 &  x375 &  x401 & ~x527 & ~x585 & ~x668 & ~x711;
assign c539 =  x305 &  x323 &  x326 &  x359 &  x361 &  x387 &  x413 &  x414 &  x464 &  x474 & ~x13 & ~x31 & ~x33 & ~x40 & ~x61 & ~x69 & ~x118 & ~x125 & ~x136 & ~x171 & ~x198 & ~x219 & ~x232 & ~x287 & ~x307 & ~x316 & ~x342 & ~x620 & ~x626 & ~x661 & ~x697 & ~x733 & ~x737;
assign c541 =  x97 & ~x529;
assign c543 =  x231;
assign c545 =  x325 &  x382 &  x403 &  x417 &  x418 &  x432 &  x443 &  x464 &  x465 &  x469 &  x472 & ~x3 & ~x6 & ~x9 & ~x20 & ~x35 & ~x37 & ~x39 & ~x47 & ~x50 & ~x80 & ~x109 & ~x126 & ~x217 & ~x223 & ~x246 & ~x312 & ~x313 & ~x363 & ~x619 & ~x627 & ~x648 & ~x694 & ~x699 & ~x713 & ~x720 & ~x739 & ~x746 & ~x771;
assign c547 =  x634 & ~x108 & ~x418 & ~x644;
assign c549 =  x242 &  x277 &  x351 &  x382 &  x411 &  x490 & ~x395;
assign c551 =  x272 &  x325 &  x361 &  x384 &  x600;
assign c553 =  x294 &  x375 &  x382 &  x405 &  x472 &  x474 &  x542 &  x556 & ~x35 & ~x664;
assign c555 =  x213 &  x270 &  x489 &  x524 & ~x427;
assign c557 =  x39;
assign c559 = ~x271 & ~x438 & ~x439 & ~x495 & ~x501 & ~x502;
assign c561 =  x42 & ~x529;
assign c563 = ~x276 & ~x304 & ~x415 & ~x430 & ~x500 & ~x501 & ~x528 & ~x563 & ~x585 & ~x759;
assign c565 =  x270 &  x275 &  x298 &  x302 &  x304 &  x405 &  x406 &  x417 &  x489 &  x491;
assign c567 =  x93;
assign c569 =  x467 &  x472 & ~x219 & ~x236 & ~x239 & ~x288 & ~x301 & ~x329 & ~x368 & ~x567 & ~x590;
assign c571 =  x69;
assign c573 =  x41;
assign c575 = ~x141 & ~x466 & ~x486 & ~x495 & ~x502 & ~x579 & ~x765;
assign c577 =  x771;
assign c579 =  x380 &  x385 &  x388 &  x404 &  x405 &  x417 &  x433 &  x437 &  x440 &  x445 &  x471 &  x474 & ~x31 & ~x34 & ~x110 & ~x173 & ~x191 & ~x218 & ~x221 & ~x288 & ~x560 & ~x626 & ~x639 & ~x644 & ~x648 & ~x654 & ~x658 & ~x663 & ~x665 & ~x686 & ~x687;
assign c581 =  x256;
assign c583 =  x14;
assign c585 =  x347 &  x372 &  x398 & ~x191 & ~x209 & ~x218 & ~x244 & ~x245 & ~x250 & ~x260 & ~x274 & ~x301 & ~x307 & ~x528 & ~x562 & ~x585 & ~x593 & ~x594 & ~x632 & ~x670 & ~x723 & ~x738;
assign c587 =  x325 & ~x162 & ~x301 & ~x498 & ~x500 & ~x501 & ~x678;
assign c589 =  x39;
assign c591 =  x242 &  x303 &  x325 &  x433 &  x467 &  x489 & ~x426;
assign c593 =  x499 &  x517 &  x520 &  x579 & ~x402;
assign c595 =  x275 &  x606 & ~x457;
assign c597 =  x361 &  x389 &  x390 & ~x5 & ~x50 & ~x140 & ~x189 & ~x261 & ~x262 & ~x501 & ~x599 & ~x612 & ~x745 & ~x775 & ~x782;
assign c599 =  x411 &  x474 & ~x256 & ~x265 & ~x294 & ~x295 & ~x348 & ~x660;
assign c5101 =  x202;
assign c5103 =  x41;
assign c5105 =  x287;
assign c5107 =  x326 &  x352 &  x380 &  x411 &  x443 & ~x122 & ~x207 & ~x374 & ~x402 & ~x426;
assign c5109 =  x258;
assign c5111 =  x214 &  x241 &  x270 &  x272 &  x275 &  x276 &  x300 &  x304 &  x325 &  x326 &  x327 &  x359 &  x382 &  x386 & ~x0 & ~x54;
assign c5113 =  x636 & ~x162;
assign c5115 = ~x408 & ~x438 & ~x465 & ~x502;
assign c5117 =  x688;
assign c5119 =  x743 & ~x500;
assign c5121 =  x243 &  x275 &  x359 &  x460 &  x520 &  x548 &  x573;
assign c5123 =  x41;
assign c5125 = ~x353 & ~x415 & ~x472 & ~x499 & ~x500 & ~x501;
assign c5127 = ~x382 & ~x460 & ~x515 & ~x529;
assign c5129 =  x41 & ~x549;
assign c5131 =  x324 &  x355 &  x360 &  x377 &  x403 &  x411 &  x415 &  x443 &  x472 & ~x42 & ~x83 & ~x99 & ~x165 & ~x221 & ~x255 & ~x264 & ~x335 & ~x394 & ~x652 & ~x705 & ~x762 & ~x764;
assign c5133 =  x259;
assign c5135 =  x302 &  x499 &  x606 & ~x457;
assign c5137 =  x273 &  x275 &  x302 &  x382 &  x489 &  x491 &  x548 & ~x370;
assign c5139 = ~x211 & ~x380 & ~x437 & ~x495 & ~x501 & ~x502 & ~x529 & ~x570 & ~x698;
assign c5141 =  x408 &  x411 &  x415 &  x442 &  x470 &  x494 &  x550 &  x553 &  x578 &  x579 & ~x36 & ~x85 & ~x168 & ~x170 & ~x198 & ~x207 & ~x285 & ~x365 & ~x718;
assign c5143 =  x349 &  x390 &  x445 &  x474 & ~x239 & ~x301;
assign c5145 =  x43;
assign c5147 =  x322 &  x390 & ~x30 & ~x84 & ~x100 & ~x110 & ~x127 & ~x211 & ~x245 & ~x262 & ~x271 & ~x299 & ~x611 & ~x612 & ~x647 & ~x689 & ~x692;
assign c5149 =  x688 & ~x307;
assign c5151 =  x232;
assign c5153 = ~x246 & ~x299 & ~x303 & ~x472 & ~x500 & ~x557;
assign c5155 = ~x219;
assign c5157 =  x202;
assign c5159 =  x349 &  x354 &  x355 &  x382 &  x384 &  x437 &  x441 &  x443 &  x444 & ~x8 & ~x16 & ~x68 & ~x86 & ~x124 & ~x134 & ~x160 & ~x203 & ~x219 & ~x243 & ~x252 & ~x301 & ~x503 & ~x646 & ~x674 & ~x741;
assign c5161 =  x68 & ~x473 & ~x501;
assign c5163 =  x89;
assign c5165 =  x325 &  x380 &  x417 &  x443 &  x457 &  x465 &  x471 &  x474 &  x491 &  x513 & ~x7 & ~x18 & ~x66 & ~x68 & ~x94 & ~x97 & ~x112 & ~x136 & ~x165 & ~x191 & ~x219 & ~x221 & ~x223 & ~x232 & ~x233 & ~x251 & ~x255 & ~x262 & ~x560 & ~x616 & ~x622 & ~x662 & ~x671 & ~x683 & ~x684 & ~x697 & ~x728 & ~x751 & ~x755 & ~x758 & ~x760;
assign c5167 =  x349 &  x382 &  x471 & ~x53 & ~x98 & ~x106 & ~x222 & ~x247 & ~x301 & ~x329 & ~x532 & ~x585 & ~x599 & ~x612 & ~x618 & ~x678 & ~x728 & ~x741 & ~x766;
assign c5169 =  x69 & ~x446;
assign c5171 =  x375 &  x404 &  x405 &  x409 &  x415 &  x417 &  x431 &  x432 &  x459 & ~x33 & ~x53 & ~x58 & ~x60 & ~x62 & ~x80 & ~x160 & ~x210 & ~x264 & ~x279 & ~x280 & ~x366 & ~x593 & ~x616 & ~x645 & ~x679 & ~x717 & ~x755 & ~x781;
assign c5173 =  x320 &  x322 &  x347 &  x372 &  x412 &  x417 &  x418 &  x443 & ~x41 & ~x96 & ~x114 & ~x119 & ~x156 & ~x214 & ~x617 & ~x631 & ~x756;
assign c5175 =  x270 &  x382 &  x387 &  x405 &  x409 &  x417 &  x431 &  x445 &  x464 &  x466 &  x491 & ~x39 & ~x74 & ~x313 & ~x342 & ~x392 & ~x664 & ~x673 & ~x741 & ~x752 & ~x757 & ~x758;
assign c5177 =  x185 &  x191 &  x213 &  x243 &  x304;
assign c5179 =  x213 &  x300 &  x381 &  x383 &  x387 &  x572 &  x584;
assign c5181 = ~x355;
assign c5183 =  x324 &  x417 &  x443 &  x468 &  x470 &  x472 &  x473 &  x474 & ~x0 & ~x20 & ~x21 & ~x103 & ~x107 & ~x143 & ~x166 & ~x186 & ~x273 & ~x274 & ~x300 & ~x301 & ~x313 & ~x366 & ~x393 & ~x561 & ~x591 & ~x595 & ~x602 & ~x630 & ~x666 & ~x687 & ~x697 & ~x698 & ~x708 & ~x717 & ~x747 & ~x773;
assign c5185 =  x242 &  x247 &  x277 &  x300 &  x301 &  x405;
assign c5187 =  x321 &  x349 &  x375 &  x382 &  x383 &  x385 &  x401 &  x417 &  x444 & ~x35 & ~x182 & ~x257 & ~x274 & ~x591 & ~x601 & ~x647 & ~x649 & ~x653 & ~x698 & ~x700 & ~x703 & ~x777;
assign c5189 =  x206;
assign c5191 =  x635 &  x663 & ~x278;
assign c5193 =  x380 &  x386 &  x387 &  x388 &  x435 &  x443 &  x472 &  x558 &  x574 &  x578;
assign c5195 =  x470 &  x474 & ~x34 & ~x46 & ~x57 & ~x90 & ~x138 & ~x145 & ~x163 & ~x188 & ~x198 & ~x207 & ~x246 & ~x259 & ~x266 & ~x275 & ~x307 & ~x329 & ~x605 & ~x698 & ~x732 & ~x773;
assign c5197 =  x128 &  x411 &  x619;
assign c5199 =  x310;
assign c5201 =  x256;
assign c5203 =  x38;
assign c5205 =  x322 &  x418 &  x474 & ~x188 & ~x216 & ~x301 & ~x328 & ~x503;
assign c5207 = ~x191 & ~x426 & ~x500 & ~x501 & ~x502 & ~x527 & ~x757;
assign c5209 =  x362 &  x410 &  x418 &  x474 & ~x239 & ~x300 & ~x301 & ~x394 & ~x591 & ~x600 & ~x612 & ~x637;
assign c5213 =  x382 &  x590;
assign c5215 =  x297 &  x322 &  x375 &  x377 &  x383 &  x402 &  x404 &  x417 &  x434 &  x435 &  x460 &  x472 &  x489 &  x490 &  x494 &  x517 & ~x149;
assign c5217 =  x230;
assign c5219 =  x744;
assign c5221 =  x191 &  x382 &  x491;
assign c5223 =  x345 &  x346 &  x356 & ~x4 & ~x29 & ~x164 & ~x207 & ~x217 & ~x218 & ~x219 & ~x245 & ~x308 & ~x560 & ~x690 & ~x697;
assign c5225 =  x716;
assign c5227 =  x178;
assign c5229 =  x635 & ~x191;
assign c5231 =  x11;
assign c5233 =  x191 &  x272 &  x275 &  x325;
assign c5235 =  x275 &  x590;
assign c5237 =  x41;
assign c5239 =  x214 &  x275 &  x304 &  x324 &  x443 &  x501;
assign c5241 =  x241 &  x324 &  x326 &  x381 &  x441 &  x442 &  x443 &  x491 &  x584;
assign c5243 =  x146;
assign c5245 =  x286;
assign c5247 =  x256;
assign c5249 =  x325 &  x327 &  x355 &  x359 &  x382 &  x386 &  x411 &  x466 &  x488 &  x612 & ~x54 & ~x251;
assign c5251 =  x202;
assign c5253 =  x213 &  x241 &  x275 &  x297 &  x331 &  x517;
assign c5255 =  x42;
assign c5257 =  x304 &  x323 &  x325 &  x382 &  x383 &  x385 &  x388 &  x404 &  x416 &  x417 &  x446 &  x462 &  x489 &  x496 & ~x94 & ~x116 & ~x147;
assign c5261 =  x323 &  x383 &  x415 &  x444 &  x468 & ~x3 & ~x22 & ~x36 & ~x51 & ~x54 & ~x61 & ~x75 & ~x79 & ~x84 & ~x100 & ~x104 & ~x106 & ~x110 & ~x111 & ~x128 & ~x160 & ~x173 & ~x183 & ~x210 & ~x221 & ~x231 & ~x236 & ~x239 & ~x264 & ~x301 & ~x394 & ~x602 & ~x604 & ~x614 & ~x643 & ~x686 & ~x700 & ~x707 & ~x754 & ~x757 & ~x776 & ~x783;
assign c5263 =  x260 &  x316;
assign c5265 =  x322 &  x325 &  x375 &  x380 &  x382 &  x404 &  x417 &  x465 & ~x54 & ~x119 & ~x134 & ~x137 & ~x219 & ~x245 & ~x599 & ~x689;
assign c5267 =  x746;
assign c5269 =  x122;
assign c5271 =  x359 &  x377 &  x382 &  x404 &  x443 &  x463 &  x469 &  x489 &  x491 &  x493 &  x524 & ~x236 & ~x393 & ~x761;
assign c5273 =  x241 &  x268 &  x273 &  x303 &  x324 &  x351 &  x520 &  x612;
assign c5275 =  x606 &  x665;
assign c5277 =  x202;
assign c5279 =  x360 &  x379 &  x382 &  x383 &  x384 &  x390 &  x474 &  x490 &  x513 & ~x65 & ~x115 & ~x162 & ~x184 & ~x197 & ~x253 & ~x314 & ~x599 & ~x609 & ~x630 & ~x721;
assign c5281 =  x203;
assign c5283 =  x214 &  x275 &  x301 &  x325 &  x388 &  x472;
assign c5285 =  x717;
assign c5287 =  x42 & ~x473;
assign c5289 =  x747;
assign c5291 =  x260;
assign c5293 =  x746;
assign c5295 =  x717;
assign c5297 =  x310;
assign c5299 =  x590 &  x618;
assign c5301 =  x13;
assign c5303 =  x321 &  x324 &  x354 &  x385 &  x388 &  x405 &  x407 &  x418 &  x465 &  x491 & ~x3 & ~x9 & ~x17 & ~x22 & ~x32 & ~x60 & ~x69 & ~x76 & ~x80 & ~x105 & ~x110 & ~x132 & ~x154 & ~x156 & ~x179 & ~x288 & ~x715 & ~x735 & ~x760 & ~x769 & ~x781;
assign c5305 =  x242 &  x275 &  x323 &  x325 &  x331 &  x359 &  x360 &  x382 &  x405 &  x529 & ~x206 & ~x691;
assign c5307 =  x355 &  x377 &  x380 &  x413 &  x433 &  x443 &  x465 &  x467 &  x470 &  x489 &  x491 &  x496 &  x499 &  x518 & ~x24 & ~x31 & ~x33 & ~x48 & ~x51 & ~x58 & ~x59 & ~x63 & ~x70 & ~x81 & ~x83 & ~x87 & ~x89 & ~x90 & ~x92 & ~x103 & ~x108 & ~x115 & ~x120 & ~x157 & ~x165 & ~x174 & ~x176 & ~x177 & ~x191 & ~x195 & ~x197 & ~x200 & ~x201 & ~x219 & ~x225 & ~x226 & ~x230 & ~x246 & ~x257 & ~x280 & ~x334 & ~x337 & ~x364 & ~x365 & ~x420 & ~x700 & ~x782;
assign c5309 =  x231;
assign c5311 =  x241 &  x244 &  x275 &  x304 &  x381 &  x388 &  x490 &  x529 & ~x426;
assign c5313 =  x313;
assign c5315 =  x118;
assign c5317 =  x405 &  x411 &  x489 & ~x95 & ~x284 & ~x316 & ~x402 & ~x773;
assign c5319 =  x295 &  x320 &  x322 &  x347 &  x360 &  x375 &  x382 &  x401 &  x404 &  x429 & ~x98 & ~x104 & ~x224 & ~x244 & ~x245 & ~x273 & ~x627 & ~x642 & ~x678 & ~x695;
assign c5321 = ~x51 & ~x299 & ~x301 & ~x471 & ~x500 & ~x501 & ~x557;
assign c5323 =  x602 &  x607 &  x614 & ~x363;
assign c5325 =  x268 &  x320 &  x449 & ~x299;
assign c5327 =  x606 & ~x29 & ~x107 & ~x191 & ~x588 & ~x728 & ~x776;
assign c5329 = ~x54 & ~x430 & ~x495 & ~x515;
assign c5331 =  x286;
assign c5333 =  x349 &  x357 &  x361 &  x375 &  x380 &  x382 &  x384 &  x388 &  x403 &  x405 &  x417 &  x442 &  x459 &  x463 &  x465 &  x467 &  x490 &  x493 & ~x16 & ~x18 & ~x54 & ~x111 & ~x143 & ~x164 & ~x624 & ~x683 & ~x727;
assign c5335 =  x297 &  x361 &  x362 &  x382 &  x384 &  x417 &  x442 &  x446 &  x463 &  x470 &  x473 &  x474 & ~x8 & ~x12 & ~x23 & ~x30 & ~x42 & ~x44 & ~x69 & ~x87 & ~x103 & ~x112 & ~x114 & ~x118 & ~x126 & ~x159 & ~x179 & ~x181 & ~x208 & ~x211 & ~x219 & ~x233 & ~x620 & ~x642 & ~x653 & ~x670 & ~x697 & ~x716 & ~x744 & ~x746 & ~x762 & ~x765;
assign c5337 =  x283;
assign c5339 =  x43;
assign c5341 =  x324 &  x351 &  x358 &  x380 &  x382 &  x385 &  x473 &  x491 &  x524 &  x554 &  x573 &  x574 &  x577 &  x578 &  x579 & ~x285 & ~x755;
assign c5343 =  x270 &  x301 &  x303 &  x323 &  x380 &  x382 &  x467 &  x489;
assign c5345 =  x382 &  x606 & ~x402 & ~x457;
assign c5347 =  x273 &  x381 &  x382 &  x404 &  x405 &  x411 &  x413 &  x437 &  x473 &  x492 &  x542 & ~x224 & ~x229 & ~x309 & ~x689 & ~x699 & ~x757;
assign c5349 =  x259;
assign c5351 =  x242 &  x275 &  x298 &  x381 &  x471 &  x489 &  x490 & ~x426;
assign c5353 =  x213 &  x326 &  x331 &  x351 &  x380 &  x382 &  x405 & ~x150;
assign c5355 =  x96 & ~x501;
assign c5357 =  x362 & ~x273 & ~x299 & ~x304 & ~x327;
assign c5359 =  x233 & ~x136;
assign c5361 =  x275 &  x304 &  x326 &  x489 & ~x402;
assign c5363 =  x309;
assign c5365 =  x380 &  x382 &  x470 &  x472 &  x494 &  x548 &  x573 & ~x427;
assign c5367 =  x14;
assign c5369 =  x382 &  x418 & ~x24 & ~x184 & ~x244 & ~x525 & ~x526 & ~x591;
assign c5371 =  x320 &  x372 &  x374 &  x401 &  x415 &  x417 & ~x211 & ~x585 & ~x775;
assign c5373 =  x213 &  x241 &  x272 &  x301 &  x302 &  x323 &  x387 &  x405 &  x491 &  x499;
assign c5375 =  x320 &  x349 &  x372 &  x375 &  x403 & ~x529 & ~x630;
assign c5377 = ~x348 & ~x430 & ~x486 & ~x494 & ~x495 & ~x499;
assign c5379 =  x255;
assign c5381 =  x259;
assign c5383 =  x633;
assign c5385 =  x43;
assign c5387 = ~x297 & ~x439 & ~x515 & ~x549 & ~x557;
assign c5389 =  x354 &  x377 & ~x6 & ~x246 & ~x291 & ~x299 & ~x328 & ~x329 & ~x619;
assign c5391 =  x270 &  x274 &  x275 &  x304 &  x355 &  x358 &  x411 &  x417 &  x493 & ~x60 & ~x396 & ~x399 & ~x401 & ~x452;
assign c5393 =  x322 &  x325 &  x389 &  x417 &  x471 & ~x197 & ~x219 & ~x525 & ~x564 & ~x598 & ~x627 & ~x659;
assign c5395 = ~x217 & ~x275 & ~x500 & ~x501 & ~x502 & ~x530;
assign c5397 =  x214 &  x221 &  x272 &  x304 &  x411;
assign c5399 =  x320 &  x322 &  x323 &  x349 &  x375 &  x377 &  x382 &  x383 &  x386 &  x404 &  x431 &  x432 &  x465 & ~x82 & ~x341 & ~x736 & ~x746 & ~x756;
assign c5401 =  x242 &  x270 &  x330 &  x354 &  x382 &  x383 &  x460 &  x489 & ~x341 & ~x398;
assign c5403 =  x447 & ~x137 & ~x219 & ~x250 & ~x392 & ~x666;
assign c5405 =  x68;
assign c5407 =  x662 &  x688;
assign c5409 =  x248 &  x276 &  x590 & ~x428;
assign c5411 =  x40;
assign c5413 =  x355 &  x417 &  x474 & ~x172 & ~x220 & ~x244 & ~x258 & ~x301 & ~x329 & ~x647;
assign c5415 =  x463 &  x572 &  x628 &  x630 &  x633;
assign c5417 =  x213 &  x304 &  x381 &  x612;
assign c5419 =  x331 &  x358 &  x377 &  x403 &  x411 &  x416 &  x432 &  x491 & ~x504;
assign c5421 =  x322 &  x418 & ~x238 & ~x276 & ~x301 & ~x599;
assign c5423 =  x93;
assign c5425 = ~x410 & ~x414 & ~x488 & ~x501 & ~x502 & ~x528;
assign c5427 =  x320 &  x325 &  x372 & ~x19 & ~x174 & ~x182 & ~x192 & ~x217 & ~x219 & ~x237 & ~x243 & ~x245 & ~x246 & ~x301 & ~x302 & ~x503 & ~x623 & ~x632 & ~x649 & ~x680 & ~x767;
assign c5429 =  x242 &  x293 &  x320 &  x330 &  x375 &  x431;
assign c5431 =  x247 &  x274 &  x275 &  x301 &  x304 &  x325 &  x383 &  x387 &  x411 &  x517 &  x518 & ~x426;
assign c5433 =  x295 &  x320 &  x347 &  x349 &  x361 &  x375 &  x405 &  x418 &  x435 &  x472 &  x474;
assign c5435 =  x123;
assign c5437 =  x318 &  x395;
assign c5439 =  x204;
assign c5441 =  x361 &  x382 &  x413 &  x436 &  x441 &  x467 &  x489 &  x491 &  x558 & ~x336 & ~x397;
assign c5443 =  x269 &  x275 &  x325 &  x351 &  x381 &  x443 &  x460 &  x471 &  x524 &  x548 & ~x3 & ~x121 & ~x260 & ~x369 & ~x756;
assign c5445 =  x320 &  x346 &  x347 &  x362 &  x400 &  x429 &  x442 &  x443 & ~x7 & ~x28 & ~x117 & ~x247 & ~x503 & ~x576 & ~x583 & ~x619 & ~x660 & ~x685 & ~x690 & ~x708 & ~x748 & ~x776;
assign c5447 =  x656 &  x661 &  x688 &  x717;
assign c5449 =  x311;
assign c5451 =  x274 &  x302 &  x381 &  x385 &  x467 &  x521 &  x600;
assign c5453 =  x234;
assign c5455 =  x241 &  x244 &  x268 &  x275 &  x301 &  x304 &  x325;
assign c5459 = ~x196 & ~x217 & ~x492 & ~x501 & ~x502 & ~x638 & ~x652 & ~x717 & ~x769;
assign c5461 =  x380 &  x383 &  x385 &  x417 &  x439 &  x441 &  x446 &  x465 &  x467 &  x471 &  x474 &  x496 & ~x1 & ~x81 & ~x92 & ~x266 & ~x675 & ~x730 & ~x750 & ~x765;
assign c5463 =  x353 &  x375 &  x377 &  x432 & ~x369 & ~x524 & ~x613 & ~x760;
assign c5465 =  x122;
assign c5467 =  x176;
assign c5469 =  x275 &  x304 &  x384 &  x467 &  x493 &  x548;
assign c5471 =  x284;
assign c5473 =  x310;
assign c5475 =  x212 &  x215 &  x221 &  x327;
assign c5477 = ~x382 & ~x493 & ~x495 & ~x501 & ~x502;
assign c5479 = ~x439 & ~x449 & ~x502 & ~x529 & ~x530;
assign c5481 =  x354 &  x382 &  x606 &  x626 &  x628;
assign c5483 =  x202;
assign c5485 = ~x4 & ~x34 & ~x116 & ~x430 & ~x466 & ~x494 & ~x499 & ~x501;
assign c5487 =  x215 &  x297 &  x304 &  x383 &  x491 &  x548 &  x573 &  x600;
assign c5489 =  x322 &  x323 &  x349 &  x351 &  x375 &  x382 &  x404 &  x405 &  x406 &  x443 &  x444 &  x462 &  x463 &  x488 &  x490 & ~x7 & ~x26 & ~x27 & ~x71 & ~x85 & ~x93 & ~x119 & ~x122 & ~x126 & ~x141 & ~x149 & ~x150 & ~x154 & ~x161 & ~x197 & ~x285 & ~x289 & ~x312 & ~x634 & ~x639 & ~x647 & ~x668 & ~x681 & ~x692 & ~x703 & ~x729 & ~x766 & ~x768;
assign c5491 = ~x426 & ~x470 & ~x498 & ~x499 & ~x500 & ~x501 & ~x528;
assign c5493 =  x318 &  x345 &  x396 &  x417;
assign c5495 =  x243 &  x272 &  x275 &  x325 &  x411;
assign c5497 =  x320 &  x347 &  x372 &  x375 & ~x218 & ~x525 & ~x528;
assign c5499 =  x320 &  x346 &  x347 &  x375 &  x376 &  x380 &  x382 &  x402 &  x403 &  x415 & ~x180 & ~x214 & ~x225 & ~x245 & ~x591 & ~x647 & ~x679;
assign c60 =  x130 &  x183 &  x271 &  x405 &  x489 &  x608 &  x636 & ~x362 & ~x454 & ~x615 & ~x644 & ~x650 & ~x669;
assign c62 =  x75 &  x123 &  x452 &  x620 &  x624 &  x636;
assign c64 =  x344 &  x404 &  x406 &  x428 &  x546 &  x679 &  x769 & ~x143 & ~x195 & ~x416 & ~x475 & ~x560 & ~x639 & ~x696 & ~x729;
assign c66 =  x73 &  x103 &  x119 &  x213 &  x435 &  x601 &  x653 & ~x46 & ~x416;
assign c68 = ~x61 & ~x202 & ~x304 & ~x362 & ~x416 & ~x477 & ~x656 & ~x684;
assign c610 = ~x656;
assign c612 =  x230 &  x377 &  x401 &  x604 & ~x12 & ~x13 & ~x15 & ~x58 & ~x166 & ~x555 & ~x669 & ~x697 & ~x732;
assign c614 = ~x274 & ~x627;
assign c616 =  x98 &  x133 &  x739 & ~x38;
assign c618 = ~x11 & ~x492;
assign c620 =  x322 &  x636 &  x652 & ~x107 & ~x469 & ~x642 & ~x728;
assign c622 =  x66 &  x471 &  x510 &  x636 &  x752;
assign c624 = ~x16 & ~x182 & ~x626;
assign c626 =  x72 &  x205 &  x214 &  x266 &  x269 &  x429 &  x490 &  x513 & ~x4 & ~x32 & ~x137 & ~x198 & ~x282 & ~x284 & ~x385 & ~x424 & ~x555 & ~x640 & ~x644 & ~x699 & ~x751;
assign c628 =  x47 &  x121 &  x245 &  x286 &  x636 & ~x16;
assign c630 =  x358 &  x541 &  x653 &  x686 & ~x19 & ~x45 & ~x109 & ~x138 & ~x254 & ~x763;
assign c632 =  x237 &  x266 &  x347 &  x350 &  x378 &  x407 &  x459 &  x495 &  x517 &  x547 &  x598 & ~x26 & ~x57 & ~x78 & ~x88 & ~x109 & ~x166 & ~x281 & ~x284 & ~x340 & ~x363 & ~x365 & ~x449 & ~x452 & ~x473 & ~x475 & ~x478 & ~x505 & ~x527 & ~x558 & ~x559 & ~x586 & ~x588 & ~x644 & ~x646 & ~x667 & ~x674 & ~x676 & ~x697 & ~x705 & ~x727 & ~x762 & ~x779 & ~x781;
assign c634 =  x39 &  x155 &  x210 &  x234 &  x295 &  x378 & ~x5 & ~x79 & ~x228 & ~x285 & ~x333 & ~x591 & ~x621;
assign c636 =  x15 &  x40 &  x742 & ~x46 & ~x50 & ~x478 & ~x562 & ~x645 & ~x763 & ~x783;
assign c638 = ~x297 & ~x380;
assign c640 =  x35 &  x48 &  x188 &  x203 &  x496 &  x521 &  x580 &  x651 &  x659 &  x664 & ~x27 & ~x28 & ~x82 & ~x137 & ~x140 & ~x141 & ~x252 & ~x448 & ~x701 & ~x755;
assign c642 =  x75 &  x155 &  x186 &  x262 &  x343 &  x347 &  x359 &  x377 &  x516 &  x601 &  x623 &  x636 & ~x83 & ~x109 & ~x167 & ~x249 & ~x421 & ~x449 & ~x700;
assign c644 =  x242 &  x258 &  x260 &  x287 &  x315 &  x343 &  x374 &  x376 &  x380 &  x436 &  x459 &  x492 &  x553 & ~x0 & ~x1 & ~x14 & ~x15 & ~x16 & ~x41 & ~x82 & ~x84 & ~x139 & ~x166 & ~x279 & ~x531;
assign c646 =  x75 &  x133 &  x331 &  x592 & ~x163;
assign c648 =  x118 &  x146 &  x483 &  x497 &  x687 &  x743 & ~x2 & ~x26 & ~x363 & ~x419 & ~x671 & ~x752 & ~x778;
assign c650 =  x105 &  x207 &  x230 &  x286 &  x344 &  x629 &  x652 &  x769 & ~x141 & ~x310 & ~x364 & ~x365 & ~x476 & ~x532 & ~x615 & ~x699 & ~x757;
assign c652 =  x210 &  x258 &  x297 &  x322 &  x377 &  x487 & ~x10 & ~x331 & ~x416 & ~x473 & ~x699;
assign c654 =  x75 &  x76 &  x103 &  x207 &  x266 &  x268 &  x298 &  x467 &  x495 &  x548 &  x568 &  x595 &  x627 &  x655 &  x679 & ~x31 & ~x58 & ~x107 & ~x420 & ~x588 & ~x672;
assign c656 =  x231 &  x441 &  x480 &  x507 & ~x142 & ~x168 & ~x194 & ~x365 & ~x422 & ~x446 & ~x616 & ~x781;
assign c658 =  x231 &  x312 &  x314 &  x357 &  x387 & ~x15 & ~x281 & ~x779;
assign c660 =  x120 &  x125 &  x186 &  x260 &  x330 &  x356 &  x433 &  x685 & ~x10 & ~x172 & ~x312 & ~x419 & ~x590 & ~x675;
assign c662 =  x49 &  x344 &  x455 & ~x112 & ~x251;
assign c664 = ~x186 & ~x319 & ~x416;
assign c666 = ~x130 & ~x185 & ~x448;
assign c668 =  x293 &  x343 &  x432 &  x440 &  x456 &  x496 &  x520 &  x721 &  x749 & ~x13 & ~x80 & ~x725;
assign c670 =  x315 &  x414 & ~x25 & ~x38 & ~x222 & ~x765;
assign c672 = ~x11 & ~x379;
assign c674 =  x92 &  x94 &  x103 &  x126 &  x323 &  x546 & ~x38 & ~x46 & ~x448 & ~x697;
assign c676 =  x243 &  x350 &  x462 &  x463 &  x546 &  x575 &  x578 &  x602 & ~x192 & ~x193 & ~x199 & ~x247 & ~x254 & ~x275 & ~x282 & ~x313 & ~x505 & ~x531 & ~x564 & ~x582 & ~x762;
assign c678 =  x40 &  x95 &  x121 &  x179 &  x202 &  x234 &  x238 &  x266 &  x295 &  x320 &  x330 &  x343 &  x350 &  x490 &  x527 &  x578 &  x634 &  x648 &  x750 & ~x89 & ~x107;
assign c680 = ~x297 & ~x682;
assign c682 =  x384 &  x439 &  x464 &  x518 &  x575 &  x652 &  x680 & ~x4 & ~x78 & ~x396 & ~x445 & ~x696;
assign c684 =  x210 &  x330 &  x518 &  x769 & ~x46;
assign c686 = ~x217 & ~x315 & ~x468;
assign c688 =  x325 &  x357 &  x387 &  x518 &  x536 &  x637 & ~x5 & ~x28 & ~x50 & ~x60 & ~x87 & ~x141 & ~x164 & ~x168 & ~x193 & ~x198 & ~x306 & ~x309 & ~x418 & ~x421;
assign c690 = ~x184 & ~x512;
assign c692 =  x105 &  x609 &  x752 & ~x192 & ~x250 & ~x766;
assign c694 = ~x514;
assign c696 = ~x158;
assign c698 =  x66 &  x73 &  x271 &  x551 &  x627 &  x658 & ~x17 & ~x18 & ~x52 & ~x54 & ~x111 & ~x136 & ~x137 & ~x169 & ~x170 & ~x200 & ~x221 & ~x228 & ~x253 & ~x254 & ~x281 & ~x311 & ~x335 & ~x367 & ~x394 & ~x449 & ~x560 & ~x561 & ~x562 & ~x641 & ~x670 & ~x764 & ~x774 & ~x780;
assign c6100 =  x133 &  x330 &  x687 & ~x38 & ~x46 & ~x194 & ~x250;
assign c6102 =  x92 & ~x38 & ~x48 & ~x197 & ~x276 & ~x307 & ~x729;
assign c6104 =  x61 &  x440 &  x608 & ~x30 & ~x140 & ~x252 & ~x532 & ~x700 & ~x757;
assign c6106 =  x161 &  x358 &  x414 &  x498 & ~x5 & ~x17 & ~x25 & ~x34 & ~x753;
assign c6108 =  x258 &  x303 &  x679 &  x693 & ~x252 & ~x392 & ~x505 & ~x640;
assign c6110 =  x414 &  x686 & ~x38 & ~x46 & ~x505;
assign c6112 =  x314 &  x343 &  x454 &  x741 & ~x11 & ~x200;
assign c6114 =  x265 &  x314 &  x345 &  x665 & ~x13 & ~x15 & ~x16 & ~x49 & ~x421 & ~x757;
assign c6116 =  x339 & ~x24 & ~x53 & ~x724;
assign c6118 =  x91 &  x209 &  x210 &  x232 &  x319 &  x328 &  x329 &  x381 &  x465 &  x550 &  x628 &  x686 & ~x9 & ~x47 & ~x53 & ~x78 & ~x80 & ~x82 & ~x107 & ~x110 & ~x168 & ~x171 & ~x280 & ~x365 & ~x447 & ~x450 & ~x506 & ~x644 & ~x756;
assign c6120 = ~x411 & ~x430;
assign c6122 = ~x74 & ~x520;
assign c6124 =  x60;
assign c6126 =  x59;
assign c6128 =  x636 & ~x141 & ~x146 & ~x226 & ~x441 & ~x593 & ~x611 & ~x674;
assign c6130 =  x269 &  x322 &  x345 &  x401 & ~x144 & ~x280 & ~x360 & ~x362 & ~x363 & ~x368 & ~x445 & ~x449 & ~x450 & ~x502 & ~x507 & ~x560 & ~x645 & ~x647 & ~x696 & ~x766;
assign c6132 =  x75 &  x637 &  x752;
assign c6134 =  x76 &  x536 & ~x163;
assign c6136 =  x217 &  x245 &  x597 &  x625 & ~x11 & ~x45 & ~x61 & ~x165 & ~x363 & ~x618 & ~x696;
assign c6138 =  x370 & ~x28 & ~x34 & ~x38 & ~x57 & ~x333 & ~x392 & ~x618 & ~x728;
assign c6140 =  x238 &  x328 &  x604 &  x679 &  x680 &  x689 &  x720 &  x742 & ~x224 & ~x392 & ~x476 & ~x588 & ~x611 & ~x639 & ~x676 & ~x724 & ~x732 & ~x781;
assign c6142 =  x595 &  x601 &  x636 & ~x20 & ~x23 & ~x31 & ~x55 & ~x280 & ~x364 & ~x447 & ~x565 & ~x593 & ~x640 & ~x644 & ~x672 & ~x696 & ~x699 & ~x700 & ~x751;
assign c6144 =  x461 &  x555 & ~x10 & ~x137 & ~x334 & ~x396;
assign c6146 =  x45 &  x233 &  x519 & ~x84 & ~x168 & ~x279 & ~x342 & ~x358 & ~x366 & ~x398 & ~x498 & ~x585 & ~x647 & ~x757 & ~x761;
assign c6148 =  x15 & ~x46 & ~x445 & ~x539;
assign c6150 =  x41 &  x44 &  x63 &  x75 &  x98 &  x156 &  x176 &  x268 &  x323 &  x349 &  x409 &  x459 &  x484 &  x487 &  x493 &  x521 &  x574 &  x575 &  x604 & ~x25 & ~x30 & ~x49 & ~x79 & ~x88 & ~x196 & ~x277 & ~x365 & ~x445 & ~x673 & ~x763;
assign c6152 =  x344 &  x427 &  x580 &  x652 & ~x4 & ~x14 & ~x195 & ~x620 & ~x639 & ~x668 & ~x695;
assign c6154 =  x266 &  x292 &  x322 &  x377 &  x513 & ~x20 & ~x25 & ~x58 & ~x250 & ~x252 & ~x448 & ~x682;
assign c6156 =  x63 &  x64 &  x75 &  x181 &  x602 &  x636 &  x724 & ~x88;
assign c6158 = ~x122 & ~x331 & ~x416;
assign c6160 =  x119 &  x328 & ~x17 & ~x45 & ~x106 & ~x361 & ~x699;
assign c6162 = ~x46 & ~x375 & ~x766;
assign c6164 = ~x46 & ~x186 & ~x381;
assign c6166 =  x35 & ~x0 & ~x12 & ~x20 & ~x53 & ~x55 & ~x60 & ~x79 & ~x137 & ~x169 & ~x195 & ~x196 & ~x560 & ~x587 & ~x672 & ~x759 & ~x783;
assign c6168 =  x61 &  x300 &  x412 & ~x29 & ~x754;
assign c6170 = ~x129 & ~x319;
assign c6172 =  x63 &  x75 &  x148 &  x230 &  x244 &  x518 &  x536 &  x565 &  x612 & ~x166 & ~x167 & ~x448 & ~x561;
assign c6174 =  x128 &  x373 &  x509 &  x585 & ~x362;
assign c6176 =  x118 &  x322 &  x564 &  x665 & ~x59 & ~x163 & ~x199 & ~x765;
assign c6178 =  x435 &  x557 & ~x6 & ~x142 & ~x221 & ~x278 & ~x306 & ~x336 & ~x779;
assign c6180 =  x267 &  x269 &  x323 &  x324 &  x349 &  x485 &  x568 &  x652 & ~x7 & ~x16 & ~x23 & ~x27 & ~x53 & ~x135 & ~x144 & ~x169 & ~x337 & ~x416 & ~x443 & ~x447 & ~x448 & ~x450 & ~x451 & ~x471 & ~x560 & ~x563 & ~x584 & ~x588 & ~x614 & ~x761;
assign c6182 =  x452 &  x585 & ~x3 & ~x14;
assign c6184 = ~x46 & ~x464;
assign c6186 =  x63 &  x752 & ~x474;
assign c6188 = ~x17 & ~x122 & ~x140 & ~x388 & ~x390 & ~x535 & ~x585 & ~x586 & ~x587;
assign c6190 =  x401 & ~x13 & ~x14 & ~x24 & ~x28 & ~x81 & ~x84 & ~x143 & ~x198 & ~x310 & ~x365 & ~x420 & ~x718 & ~x728;
assign c6192 = ~x17 & ~x46 & ~x136 & ~x479 & ~x527 & ~x530 & ~x536 & ~x583 & ~x759 & ~x762;
assign c6194 =  x273 &  x369 &  x536 & ~x13 & ~x16 & ~x29 & ~x35 & ~x140 & ~x142 & ~x225 & ~x783;
assign c6196 = ~x158 & ~x467;
assign c6198 =  x479 &  x585;
assign c6200 =  x65 &  x103 &  x232 &  x322 &  x327 &  x544 &  x575 &  x579 &  x602 &  x608 &  x631 &  x636 &  x652 &  x686 &  x707 & ~x249 & ~x251 & ~x278 & ~x308 & ~x395 & ~x444 & ~x448 & ~x479 & ~x504 & ~x671 & ~x728 & ~x779;
assign c6202 =  x103 &  x214 &  x264 &  x289 &  x350 &  x405 &  x495 &  x520 &  x657 & ~x55 & ~x80 & ~x143 & ~x256 & ~x312 & ~x334 & ~x396 & ~x420 & ~x421 & ~x502 & ~x582 & ~x612 & ~x617 & ~x640 & ~x673 & ~x674 & ~x731 & ~x732 & ~x755 & ~x780;
assign c6204 =  x119 & ~x106 & ~x451 & ~x735 & ~x760 & ~x766 & ~x783;
assign c6206 =  x62 & ~x6 & ~x13 & ~x16 & ~x34 & ~x141 & ~x365 & ~x421 & ~x423 & ~x783;
assign c6208 =  x143;
assign c6210 = ~x464;
assign c6212 =  x400 &  x577 &  x623 &  x652 & ~x57 & ~x393 & ~x471 & ~x537 & ~x555 & ~x563;
assign c6214 =  x67 &  x234 &  x267 &  x296 &  x378 &  x383 &  x597 &  x603 & ~x82 & ~x85 & ~x165 & ~x247 & ~x252 & ~x503 & ~x536 & ~x556 & ~x621 & ~x668 & ~x759;
assign c6216 =  x161 &  x230 &  x408 &  x544 &  x599 &  x654 &  x689 &  x715 & ~x46 & ~x47 & ~x764;
assign c6218 =  x64 &  x65 &  x75 &  x92 &  x120 &  x214 &  x293 &  x294 &  x460 &  x464 &  x467 & ~x7 & ~x35 & ~x60 & ~x111 & ~x113 & ~x143 & ~x168 & ~x191 & ~x194 & ~x199 & ~x200 & ~x220 & ~x306 & ~x332 & ~x450 & ~x531 & ~x590 & ~x646;
assign c6220 =  x36 &  x187 &  x411 &  x412 & ~x2 & ~x16 & ~x51 & ~x138 & ~x196 & ~x223 & ~x306 & ~x620;
assign c6222 =  x262 &  x298 & ~x217 & ~x426;
assign c6224 = ~x269 & ~x542;
assign c6226 = ~x45 & ~x319;
assign c6228 =  x60;
assign c6230 =  x103 & ~x45 & ~x64 & ~x669 & ~x748;
assign c6232 = ~x38 & ~x428;
assign c6234 =  x232 &  x387 &  x455 &  x491 & ~x620 & ~x673 & ~x696;
assign c6236 =  x203 &  x266 &  x330 &  x457 &  x563 & ~x3 & ~x25 & ~x110 & ~x192 & ~x305 & ~x775;
assign c6238 =  x35 &  x455 &  x651 & ~x5 & ~x58 & ~x84 & ~x137 & ~x337 & ~x392 & ~x393 & ~x700 & ~x755;
assign c6240 =  x36 &  x235 &  x261 & ~x476 & ~x640 & ~x677 & ~x732;
assign c6242 =  x95 &  x495 &  x519 & ~x315 & ~x398 & ~x497 & ~x528 & ~x555 & ~x610;
assign c6244 = ~x46 & ~x655;
assign c6246 = ~x458;
assign c6248 = ~x376;
assign c6250 = ~x238 & ~x297 & ~x466;
assign c6252 = ~x11 & ~x239 & ~x467;
assign c6254 =  x67 &  x75 &  x105 &  x203 &  x260 &  x620 &  x640 &  x668 & ~x54 & ~x226;
assign c6256 = ~x45 & ~x365 & ~x389 & ~x468 & ~x476 & ~x496 & ~x762;
assign c6258 = ~x269 & ~x319;
assign c6260 =  x291 &  x319 &  x345 &  x602 &  x680 & ~x86 & ~x134 & ~x135 & ~x192 & ~x342 & ~x398 & ~x445 & ~x560 & ~x586 & ~x590 & ~x778;
assign c6262 =  x546 &  x569 & ~x56 & ~x80 & ~x144 & ~x228 & ~x274 & ~x285 & ~x315 & ~x357 & ~x498 & ~x531 & ~x593 & ~x753 & ~x759;
assign c6264 = ~x411 & ~x514;
assign c6266 = ~x359 & ~x594 & ~x682 & ~x752;
assign c6268 =  x63 &  x752 & ~x310;
assign c6270 =  x118 &  x331 & ~x615 & ~x639 & ~x728 & ~x751 & ~x781;
assign c6272 =  x104 &  x378 &  x595 & ~x10 & ~x34 & ~x60 & ~x112 & ~x169 & ~x193 & ~x256 & ~x647;
assign c6274 = ~x45 & ~x383;
assign c6276 =  x373 &  x710 & ~x38 & ~x46 & ~x757 & ~x765;
assign c6278 =  x119 &  x741 & ~x46 & ~x529;
assign c6280 = ~x38 & ~x358 & ~x457;
assign c6282 =  x101 &  x149 &  x213 &  x769 & ~x17 & ~x37 & ~x50 & ~x364;
assign c6284 =  x262 &  x266 &  x268 &  x291 &  x321 &  x324 &  x327 &  x346 &  x354 &  x381 &  x406 &  x408 &  x439 &  x460 &  x466 &  x494 &  x495 & ~x26 & ~x162 & ~x223 & ~x278 & ~x446 & ~x477 & ~x500 & ~x671 & ~x761 & ~x766;
assign c6286 =  x63 &  x245 &  x322 &  x387 &  x415 &  x425 &  x438 &  x536 &  x580 &  x608 &  x636 & ~x30 & ~x672 & ~x764 & ~x775;
assign c6288 =  x260 &  x286 & ~x11 & ~x39 & ~x446 & ~x504 & ~x505 & ~x561;
assign c6290 = ~x202 & ~x484 & ~x624;
assign c6292 =  x42 & ~x376 & ~x766;
assign c6294 = ~x498 & ~x507 & ~x682;
assign c6296 =  x668 & ~x30 & ~x137 & ~x200 & ~x615 & ~x765;
assign c6298 = ~x11 & ~x467;
assign c6300 =  x59;
assign c6302 =  x36 &  x47 &  x273 &  x368 &  x412 &  x437 &  x455 & ~x762;
assign c6304 =  x581 &  x752 & ~x140 & ~x737;
assign c6306 =  x43 &  x267 &  x327 &  x489 &  x492 &  x571 &  x680 & ~x79 & ~x305 & ~x342 & ~x426 & ~x471 & ~x481 & ~x610;
assign c6308 =  x416 &  x452 & ~x249 & ~x310 & ~x762 & ~x764;
assign c6310 =  x282;
assign c6312 = ~x17 & ~x158 & ~x337 & ~x453;
assign c6314 =  x205 &  x511 &  x549 &  x623 & ~x13 & ~x14 & ~x15 & ~x165 & ~x280 & ~x309 & ~x333 & ~x533 & ~x761 & ~x778;
assign c6316 =  x73 &  x132 &  x344 &  x425 &  x429 &  x689 & ~x46 & ~x114 & ~x277 & ~x305;
assign c6318 =  x92 &  x322 &  x350 & ~x47 & ~x168 & ~x249 & ~x501 & ~x618 & ~x765 & ~x766;
assign c6320 =  x326 &  x328 &  x686 &  x749 & ~x527;
assign c6322 =  x284 &  x343 & ~x583 & ~x702 & ~x730;
assign c6324 =  x579 & ~x135 & ~x198 & ~x315 & ~x341 & ~x413 & ~x416 & ~x426;
assign c6326 =  x283 & ~x646 & ~x780;
assign c6328 =  x146 &  x625 &  x744 & ~x8 & ~x18 & ~x46 & ~x534 & ~x748 & ~x754 & ~x775;
assign c6330 =  x311 & ~x16 & ~x22;
assign c6332 = ~x235 & ~x309 & ~x530 & ~x641 & ~x766;
assign c6334 =  x92 &  x97 &  x104 &  x162 &  x177 &  x179 &  x190 &  x231 &  x234 &  x238 &  x243 &  x261 &  x323 &  x387 &  x406 &  x452 &  x495 &  x579 &  x595 & ~x673 & ~x761;
assign c6336 =  x284 &  x330 &  x369 & ~x15 & ~x751 & ~x755 & ~x761 & ~x779;
assign c6338 =  x43 &  x330 &  x384 &  x657 & ~x74 & ~x419 & ~x619 & ~x673;
assign c6340 = ~x10 & ~x45 & ~x107 & ~x351;
assign c6342 =  x440 &  x460 &  x636 &  x679 & ~x136 & ~x426 & ~x696 & ~x752;
assign c6344 =  x66 &  x74 &  x91 &  x131 &  x182 &  x573 &  x716 & ~x10 & ~x25 & ~x78 & ~x253 & ~x364 & ~x474 & ~x776;
assign c6346 =  x38 &  x75 &  x91 &  x104 &  x118 &  x182 &  x273 &  x330 &  x343 &  x344 &  x345 &  x353 &  x406 &  x410 &  x427 &  x430 &  x463 &  x490 &  x545 &  x576 &  x627 &  x630 & ~x54 & ~x111 & ~x196 & ~x754 & ~x762;
assign c6348 =  x210 &  x395 & ~x752;
assign c6350 = ~x6 & ~x13 & ~x31 & ~x110 & ~x166 & ~x225 & ~x362 & ~x681 & ~x699;
assign c6352 =  x230 & ~x15 & ~x39 & ~x164;
assign c6354 =  x203 & ~x38 & ~x45 & ~x46 & ~x64 & ~x646 & ~x748;
assign c6356 =  x73 &  x91 &  x133 &  x244 &  x321 &  x359 &  x384 &  x399 &  x491 &  x525 &  x556 &  x612 & ~x8 & ~x79 & ~x83 & ~x221 & ~x362;
assign c6358 =  x284 &  x357 & ~x222 & ~x365 & ~x618 & ~x674 & ~x751;
assign c6360 =  x35 &  x286 &  x328 &  x399 & ~x15 & ~x250 & ~x282 & ~x307 & ~x308 & ~x364 & ~x448;
assign c6362 =  x319 &  x484 &  x573 & ~x2 & ~x35 & ~x79 & ~x247 & ~x392 & ~x640 & ~x647 & ~x754;
assign c6364 =  x132 &  x202 &  x315 &  x683 & ~x2 & ~x9 & ~x45 & ~x85 & ~x110 & ~x141 & ~x220 & ~x335 & ~x703 & ~x731 & ~x758;
assign c6366 = ~x208 & ~x241 & ~x439;
assign c6368 = ~x17 & ~x74 & ~x430;
assign c6370 =  x330 &  x685 &  x691 & ~x45;
assign c6372 =  x118 &  x323 &  x630 &  x683 &  x711 & ~x28 & ~x88 & ~x227 & ~x725 & ~x731 & ~x732 & ~x733 & ~x753 & ~x761 & ~x778;
assign c6374 =  x274 &  x603 & ~x46 & ~x478 & ~x533 & ~x675 & ~x728;
assign c6376 =  x65 &  x75 &  x121 &  x261 &  x326 &  x382 &  x401 &  x408 & ~x135 & ~x174;
assign c6378 =  x270 &  x458 &  x468 &  x574 &  x636 &  x707 & ~x593 & ~x780;
assign c6380 =  x75 &  x343 & ~x3 & ~x47 & ~x644;
assign c6382 = ~x376;
assign c6384 =  x264 &  x536 &  x668 & ~x172 & ~x220;
assign c6386 = ~x101 & ~x269;
assign c6388 = ~x404 & ~x466 & ~x549;
assign c6390 =  x103 &  x537 &  x718 & ~x38;
assign c6392 = ~x184 & ~x492 & ~x652;
assign c6394 =  x12 &  x91 &  x92 &  x231 &  x414 &  x691 & ~x107 & ~x138 & ~x192 & ~x222 & ~x227 & ~x338 & ~x782;
assign c6396 =  x97 &  x100 &  x132 &  x161 &  x184 &  x186 &  x206 &  x214 &  x231 &  x237 &  x266 &  x290 &  x321 &  x349 &  x350 &  x380 &  x457 &  x514 &  x516 &  x575 &  x597 &  x631 &  x652 &  x683 &  x686 & ~x29 & ~x61 & ~x83 & ~x87 & ~x111 & ~x163 & ~x250 & ~x308 & ~x393 & ~x447 & ~x507 & ~x562 & ~x702 & ~x776;
assign c6398 = ~x383 & ~x571;
assign c6400 =  x60;
assign c6402 =  x452 &  x630 &  x636 & ~x56 & ~x338 & ~x763 & ~x766;
assign c6404 = ~x494;
assign c6406 =  x93 &  x102 &  x231 &  x317 & ~x1 & ~x37 & ~x45 & ~x227;
assign c6408 =  x266 &  x439 &  x456 &  x486 &  x623 &  x633 &  x679 &  x692 & ~x25 & ~x112 & ~x198 & ~x477 & ~x557 & ~x582 & ~x592 & ~x647 & ~x700 & ~x779;
assign c6410 =  x468 &  x492 &  x636 & ~x12 & ~x16 & ~x506 & ~x555 & ~x582 & ~x615 & ~x645;
assign c6412 =  x570 &  x686 & ~x2 & ~x29 & ~x34 & ~x35 & ~x194 & ~x249 & ~x421 & ~x454 & ~x469 & ~x471 & ~x505 & ~x507 & ~x535 & ~x581 & ~x778;
assign c6414 =  x75 &  x244 &  x271 &  x301 &  x387 &  x405 &  x536 &  x624 &  x627 & ~x255 & ~x588 & ~x765;
assign c6416 = ~x11 & ~x347 & ~x684 & ~x766;
assign c6418 =  x12 &  x302 &  x652 &  x685 & ~x46 & ~x62 & ~x109 & ~x114 & ~x166 & ~x591;
assign c6420 =  x178 &  x236 &  x608 &  x652 & ~x1 & ~x86 & ~x107 & ~x425 & ~x442 & ~x454 & ~x696;
assign c6422 =  x36 &  x229 &  x317 &  x320 &  x328 &  x345 &  x408 & ~x2 & ~x11 & ~x16 & ~x142;
assign c6424 =  x231 &  x242 & ~x39 & ~x308 & ~x418;
assign c6426 =  x219 &  x231 &  x245 &  x272 &  x315 &  x371 &  x552 &  x623 &  x624 &  x684 &  x686 & ~x223 & ~x252 & ~x758 & ~x779;
assign c6428 =  x12 &  x69 &  x73 &  x92 &  x266 &  x290 &  x294 &  x354 &  x522 & ~x27 & ~x47 & ~x50 & ~x57 & ~x136 & ~x223 & ~x278 & ~x476 & ~x505 & ~x532 & ~x560 & ~x563 & ~x669 & ~x699;
assign c6430 =  x653 &  x709 & ~x45 & ~x226 & ~x449 & ~x702;
assign c6432 =  x343 & ~x205;
assign c6434 =  x60;
assign c6436 =  x348 &  x400 &  x404 &  x429 &  x493 &  x545 &  x546 &  x575 &  x680 &  x714 & ~x275 & ~x285 & ~x358 & ~x362 & ~x479 & ~x584 & ~x779;
assign c6438 =  x323 &  x485 &  x490 &  x608 &  x680 & ~x424 & ~x475 & ~x482 & ~x526 & ~x611 & ~x762;
assign c6440 =  x10 &  x294 &  x350 &  x547 & ~x193 & ~x531 & ~x555 & ~x557 & ~x640 & ~x675 & ~x724;
assign c6442 = ~x376 & ~x686;
assign c6444 =  x121 &  x320 &  x349 &  x433 &  x434 &  x578 &  x686 & ~x83 & ~x370 & ~x498 & ~x582 & ~x702;
assign c6446 =  x339 & ~x675;
assign c6448 =  x238 &  x327 &  x495 & ~x145 & ~x275 & ~x419 & ~x471 & ~x502 & ~x558 & ~x704 & ~x779;
assign c6450 = ~x235 & ~x541;
assign c6452 = ~x237 & ~x347;
assign c6454 =  x34 &  x61;
assign c6456 =  x597 & ~x45 & ~x135 & ~x227 & ~x423 & ~x675 & ~x781;
assign c6458 =  x210 &  x231 &  x355 &  x385 &  x602 &  x657 & ~x57 & ~x640 & ~x751;
assign c6460 =  x119 &  x161 &  x214 &  x343 & ~x46 & ~x117;
assign c6462 =  x372 &  x380 &  x408 &  x462 &  x464 &  x468 &  x599 &  x602 &  x689 &  x693 &  x707 & ~x55 & ~x363 & ~x532 & ~x620 & ~x752 & ~x779;
assign c6464 =  x326 &  x330 &  x376 &  x493 &  x684 &  x688 &  x718 &  x750 & ~x54 & ~x79 & ~x163 & ~x167 & ~x169;
assign c6466 =  x75 &  x180 &  x314 &  x321 &  x406 &  x452 & ~x227 & ~x311 & ~x394;
assign c6468 =  x367 & ~x308;
assign c6470 =  x104 &  x182 &  x211 &  x271 &  x372 &  x383 &  x406 &  x486 &  x493 &  x546 &  x570 &  x575 &  x655 &  x686 &  x769 & ~x25 & ~x57 & ~x110 & ~x138 & ~x251 & ~x254 & ~x281 & ~x392 & ~x423 & ~x446 & ~x534 & ~x535 & ~x555 & ~x565 & ~x613 & ~x670 & ~x761;
assign c6472 =  x401 & ~x627;
assign c6474 =  x119 &  x288 &  x318 &  x600 &  x601 &  x655 &  x658 & ~x5 & ~x6 & ~x20 & ~x46 & ~x53 & ~x116 & ~x135 & ~x140 & ~x193 & ~x308 & ~x309 & ~x310 & ~x333 & ~x367 & ~x473 & ~x501 & ~x502 & ~x616 & ~x775;
assign c6476 =  x35 &  x36 &  x48 &  x384 &  x455 &  x520 &  x688 & ~x420 & ~x727;
assign c6478 =  x182 &  x209 &  x322 &  x405 &  x489 &  x601 & ~x4 & ~x12 & ~x60 & ~x85 & ~x310 & ~x363 & ~x422 & ~x442 & ~x450 & ~x471 & ~x481 & ~x506 & ~x647 & ~x697 & ~x731 & ~x753 & ~x781;
assign c6480 = ~x39 & ~x410;
assign c6482 =  x75 &  x581 &  x752 & ~x169;
assign c6484 =  x327 &  x462 &  x484 &  x496 &  x549 &  x573 &  x636 &  x654 &  x692 & ~x421 & ~x453 & ~x477 & ~x591;
assign c6486 =  x327 &  x405 &  x458 &  x487 &  x495 &  x547 &  x596 &  x686 &  x720 & ~x28 & ~x164 & ~x169 & ~x223 & ~x342 & ~x506 & ~x700 & ~x725 & ~x757;
assign c6488 =  x302 & ~x38 & ~x113 & ~x339 & ~x764;
assign c6490 = ~x184;
assign c6492 =  x259 &  x322 &  x384 &  x387 &  x432 &  x526 &  x536 &  x554 & ~x34 & ~x86 & ~x142 & ~x310 & ~x393 & ~x394 & ~x585;
assign c6494 =  x50;
assign c6496 =  x731 & ~x748 & ~x771;
assign c6498 = ~x180 & ~x439;
assign c61 = ~x299 & ~x300 & ~x534 & ~x666;
assign c63 =  x739 & ~x3 & ~x21 & ~x26 & ~x81 & ~x190 & ~x528 & ~x622 & ~x665 & ~x672 & ~x693 & ~x706 & ~x728;
assign c65 = ~x434 & ~x489;
assign c67 =  x736 &  x764 &  x765;
assign c69 =  x392;
assign c611 = ~x406 & ~x409 & ~x633 & ~x746;
assign c613 =  x613;
assign c615 =  x503;
assign c617 =  x566 &  x568 & ~x91 & ~x92;
assign c619 =  x466 & ~x69 & ~x70 & ~x204;
assign c621 =  x223;
assign c623 =  x0;
assign c625 = ~x226 & ~x340 & ~x363 & ~x415 & ~x445 & ~x532 & ~x608 & ~x623 & ~x664 & ~x719 & ~x720;
assign c627 =  x11 &  x16 &  x273 &  x691 &  x736;
assign c629 =  x222;
assign c631 =  x70 &  x175 &  x237 & ~x24 & ~x113 & ~x360 & ~x384 & ~x440;
assign c635 = ~x24 & ~x27 & ~x80 & ~x141 & ~x226 & ~x278 & ~x308 & ~x333 & ~x392 & ~x413 & ~x420 & ~x423 & ~x427 & ~x444 & ~x453 & ~x455 & ~x471 & ~x506 & ~x511 & ~x528 & ~x595 & ~x613 & ~x616 & ~x622 & ~x623 & ~x639 & ~x646 & ~x665 & ~x693 & ~x694 & ~x734 & ~x756 & ~x759;
assign c637 = ~x68 & ~x289 & ~x662;
assign c639 =  x40 &  x181 &  x457 &  x516 &  x626 &  x662 &  x682 & ~x19 & ~x91 & ~x92 & ~x111 & ~x333 & ~x366 & ~x783;
assign c641 =  x392;
assign c643 =  x43 &  x97 &  x435 &  x543 &  x547 &  x606 &  x709 &  x765 &  x766 &  x768 &  x773 &  x774 &  x775 & ~x59 & ~x529;
assign c645 = ~x119 & ~x288;
assign c647 = ~x124 & ~x286 & ~x287;
assign c649 =  x175 &  x181 &  x212 &  x375 &  x424 &  x508 &  x510 &  x550 &  x633 & ~x753 & ~x769 & ~x770;
assign c653 = ~x92 & ~x118 & ~x127 & ~x741 & ~x742;
assign c655 = ~x98 & ~x181 & ~x236;
assign c657 =  x40 &  x42 &  x122 &  x130 &  x215 &  x316 &  x319 &  x409 &  x435 &  x438 &  x441 &  x485 &  x662 & ~x63 & ~x76 & ~x79 & ~x85 & ~x116 & ~x134 & ~x277 & ~x534;
assign c659 = ~x67 & ~x148 & ~x258;
assign c661 =  x606 &  x660 & ~x47 & ~x91 & ~x104 & ~x118;
assign c663 =  x0;
assign c665 = ~x70 & ~x286;
assign c667 =  x261 &  x466 &  x628 &  x634 &  x748 & ~x7 & ~x113 & ~x197 & ~x306 & ~x397 & ~x447 & ~x472 & ~x481 & ~x530 & ~x622 & ~x640 & ~x671 & ~x705;
assign c669 =  x16 & ~x111 & ~x452 & ~x622 & ~x665 & ~x706;
assign c671 =  x130 &  x131 &  x181 &  x204 &  x236 &  x245 &  x262 &  x264 &  x294 &  x296 &  x300 &  x373 &  x375 &  x437 &  x457 &  x465 &  x509 &  x516 &  x546 &  x573 &  x694 &  x705 &  x722 & ~x33 & ~x86 & ~x169 & ~x225 & ~x311 & ~x503 & ~x741 & ~x742 & ~x743 & ~x744 & ~x745 & ~x747 & ~x769;
assign c673 =  x160 &  x175 &  x259 & ~x387 & ~x499 & ~x637 & ~x693 & ~x702 & ~x706;
assign c675 = ~x231 & ~x288;
assign c677 = ~x155 & ~x216;
assign c679 =  x605 &  x634 &  x692 &  x765 &  x766 &  x774 &  x775;
assign c681 =  x739 & ~x356 & ~x384 & ~x412 & ~x645;
assign c683 = ~x266 & ~x578 & ~x716;
assign c685 =  x77 &  x219 &  x230 &  x275 &  x550 &  x662 & ~x367;
assign c687 =  x739 & ~x26 & ~x88 & ~x134 & ~x146 & ~x195 & ~x201 & ~x227 & ~x446 & ~x474 & ~x561 & ~x563 & ~x668 & ~x693 & ~x701 & ~x727 & ~x753;
assign c689 =  x403 &  x413 &  x482 &  x523 &  x596 &  x599 & ~x25 & ~x105 & ~x781;
assign c691 =  x70 &  x182 &  x605 & ~x110 & ~x311 & ~x497 & ~x511 & ~x525 & ~x591 & ~x666 & ~x673;
assign c693 =  x26;
assign c695 =  x212 &  x272 &  x402 &  x544 & ~x108 & ~x415 & ~x622 & ~x665;
assign c697 =  x762 &  x777;
assign c699 = ~x71 & ~x634;
assign c6101 =  x654 &  x660 &  x746 & ~x104 & ~x118 & ~x134 & ~x474;
assign c6103 =  x435 &  x736 & ~x368 & ~x619 & ~x637 & ~x665 & ~x678 & ~x693 & ~x706;
assign c6105 = ~x43 & ~x66 & ~x258 & ~x313;
assign c6107 =  x11 &  x14;
assign c6109 =  x30;
assign c6111 =  x336;
assign c6113 = ~x68 & ~x70 & ~x230;
assign c6115 =  x96 & ~x104 & ~x109 & ~x118 & ~x134 & ~x173 & ~x218 & ~x219 & ~x246 & ~x335 & ~x449 & ~x585 & ~x645 & ~x674 & ~x698 & ~x726;
assign c6117 =  x40 &  x130 &  x625 &  x744 &  x747 & ~x7 & ~x23 & ~x387 & ~x388 & ~x693 & ~x694 & ~x703 & ~x734;
assign c6119 =  x89 &  x106 &  x633 &  x736 &  x737 & ~x56;
assign c6121 =  x89 &  x654 &  x711;
assign c6125 = ~x65 & ~x93 & ~x118 & ~x148 & ~x176 & ~x181 & ~x210;
assign c6127 =  x148 &  x183 &  x232 &  x240 &  x403 &  x404 &  x433 & ~x87 & ~x308 & ~x504 & ~x562 & ~x741 & ~x742 & ~x745 & ~x746 & ~x753 & ~x770;
assign c6129 =  x56;
assign c6131 =  x149 &  x229 &  x237 &  x426 &  x430 &  x516 &  x621 &  x625 &  x705 & ~x164 & ~x477 & ~x697 & ~x741 & ~x742 & ~x744 & ~x756 & ~x769;
assign c6133 = ~x67 & ~x71 & ~x160;
assign c6135 =  x145 &  x191 &  x219 &  x256 &  x379 &  x625 & ~x281;
assign c6137 =  x69 &  x236 &  x272 &  x341 &  x509 &  x513 &  x527 &  x542 &  x543 &  x544 &  x649 & ~x8 & ~x30 & ~x31 & ~x701 & ~x741 & ~x742 & ~x743 & ~x745 & ~x769;
assign c6139 =  x420;
assign c6141 =  x41 &  x155 &  x201 &  x330 &  x517 &  x547 &  x705 &  x732 & ~x725;
assign c6143 = ~x40 & ~x98;
assign c6145 = ~x69 & ~x232;
assign c6147 =  x11 & ~x8;
assign c6149 =  x498 & ~x685 & ~x687 & ~x690 & ~x714 & ~x716;
assign c6151 =  x54;
assign c6153 =  x362;
assign c6155 =  x44 &  x125 &  x131 &  x341 &  x373 &  x435 &  x514 &  x599 &  x629 &  x649 &  x705 &  x761 & ~x59 & ~x88;
assign c6157 = ~x285 & ~x300 & ~x356 & ~x396 & ~x399 & ~x412 & ~x424 & ~x427 & ~x537 & ~x640 & ~x759;
assign c6159 =  x121 &  x375 &  x632 & ~x310 & ~x552 & ~x608;
assign c6161 =  x124 &  x125 &  x376 &  x654 & ~x609 & ~x637 & ~x648 & ~x665 & ~x706;
assign c6163 =  x85;
assign c6165 =  x120 &  x191 &  x748 & ~x141 & ~x361 & ~x538 & ~x558;
assign c6167 = ~x2 & ~x4 & ~x10 & ~x25 & ~x32 & ~x33 & ~x36 & ~x47 & ~x48 & ~x56 & ~x60 & ~x75 & ~x81 & ~x91 & ~x92 & ~x104 & ~x118 & ~x119 & ~x133 & ~x134 & ~x140 & ~x142 & ~x146 & ~x166 & ~x223 & ~x307 & ~x336 & ~x615 & ~x725 & ~x759;
assign c6169 =  x504;
assign c6171 =  x17 &  x635 &  x774 & ~x142;
assign c6173 =  x43 &  x125 &  x543 &  x662 & ~x7 & ~x50 & ~x91 & ~x134 & ~x146 & ~x252 & ~x364 & ~x419 & ~x420 & ~x642 & ~x756;
assign c6175 =  x500 &  x528 &  x541 &  x684 &  x709;
assign c6177 =  x195;
assign c6179 =  x44 &  x130 &  x380 &  x403 &  x435 &  x497 & ~x91 & ~x105 & ~x134;
assign c6181 =  x392;
assign c6183 =  x748;
assign c6185 =  x138;
assign c6187 = ~x0 & ~x6 & ~x21 & ~x135 & ~x164 & ~x166 & ~x254 & ~x449 & ~x475 & ~x561 & ~x563 & ~x608 & ~x613 & ~x642 & ~x664 & ~x708 & ~x719 & ~x720 & ~x730 & ~x736;
assign c6189 =  x44 &  x70 &  x409 &  x461 &  x515 &  x661 &  x689 &  x739 & ~x171 & ~x397 & ~x445 & ~x508 & ~x564 & ~x665 & ~x666 & ~x678 & ~x695 & ~x705 & ~x706;
assign c6191 = ~x9 & ~x463 & ~x713 & ~x741 & ~x742 & ~x769;
assign c6193 = ~x69 & ~x97 & ~x125 & ~x148;
assign c6195 = ~x489 & ~x517 & ~x742 & ~x744;
assign c6197 =  x22;
assign c6201 = ~x70 & ~x97 & ~x124 & ~x181;
assign c6203 =  x147 &  x435 &  x436 &  x626 &  x736 & ~x86 & ~x509 & ~x622 & ~x694 & ~x729;
assign c6205 =  x122 &  x131 &  x217 &  x238 &  x240 &  x351 &  x397 &  x606 &  x723 &  x733 &  x751 & ~x310 & ~x392 & ~x502 & ~x561 & ~x644 & ~x700 & ~x744 & ~x745;
assign c6207 =  x251;
assign c6209 = ~x288;
assign c6211 =  x55;
assign c6213 =  x14 &  x566 & ~x5 & ~x105 & ~x134;
assign c6215 =  x403 &  x519 &  x735 & ~x316;
assign c6217 =  x600 &  x739 &  x768 & ~x287;
assign c6219 =  x192 & ~x510;
assign c6221 =  x501;
assign c6223 =  x28;
assign c6225 =  x766 &  x767 &  x771 &  x774 &  x775;
assign c6227 =  x42 &  x706 & ~x419 & ~x701 & ~x709 & ~x713 & ~x714 & ~x715 & ~x719 & ~x740 & ~x741 & ~x742 & ~x745 & ~x746 & ~x764 & ~x769;
assign c6229 =  x11 &  x70 &  x736;
assign c6231 =  x448;
assign c6233 =  x698;
assign c6235 =  x446;
assign c6237 = ~x70 & ~x93 & ~x202;
assign c6239 =  x24;
assign c6241 =  x307;
assign c6243 = ~x201 & ~x596 & ~x636 & ~x637 & ~x708;
assign c6245 =  x172 &  x173 &  x191 &  x219 &  x464 &  x551 &  x568 & ~x165 & ~x198 & ~x502;
assign c6247 =  x96 &  x102 &  x124 &  x130 &  x147 &  x180 &  x212 &  x246 &  x269 &  x302 &  x341 &  x373 &  x439 &  x442 &  x514 &  x517 &  x538 &  x582 &  x599 &  x611 &  x621 &  x625 &  x660 &  x666 & ~x8 & ~x116 & ~x141 & ~x164 & ~x249 & ~x254 & ~x364 & ~x448 & ~x561 & ~x585 & ~x641 & ~x701 & ~x769 & ~x770;
assign c6249 =  x43 &  x130 &  x175 &  x181 &  x229 &  x438 &  x467 &  x513 &  x538 &  x554 &  x621 &  x705 & ~x730 & ~x741 & ~x742 & ~x745;
assign c6253 =  x337;
assign c6255 =  x40 &  x229 &  x269 &  x328 &  x341 &  x424 &  x514 &  x606 &  x611 &  x621 &  x649 &  x662 &  x663 &  x723 & ~x769;
assign c6257 =  x219 &  x293 &  x410 &  x583 & ~x769;
assign c6259 =  x532;
assign c6261 = ~x66 & ~x67 & ~x103 & ~x127 & ~x132 & ~x154;
assign c6263 =  x364;
assign c6265 = ~x489 & ~x657 & ~x658 & ~x685;
assign c6267 =  x97 &  x218 &  x313 & ~x107 & ~x115 & ~x279 & ~x738 & ~x741 & ~x742 & ~x745 & ~x766 & ~x770;
assign c6269 = ~x5 & ~x29 & ~x65 & ~x91 & ~x92 & ~x103 & ~x104 & ~x114 & ~x118 & ~x120 & ~x132 & ~x134 & ~x146 & ~x147 & ~x160 & ~x171 & ~x190 & ~x201;
assign c6271 =  x130 &  x155 &  x211 &  x216 &  x232 &  x236 &  x240 &  x292 &  x293 &  x320 &  x326 &  x330 &  x341 &  x385 &  x414 &  x432 &  x433 &  x461 &  x492 &  x518 &  x519 &  x547 &  x573 &  x610 &  x611 &  x723 & ~x30 & ~x54 & ~x78 & ~x109 & ~x226 & ~x253 & ~x502 & ~x534 & ~x669 & ~x674 & ~x728 & ~x741 & ~x742 & ~x744 & ~x745 & ~x746 & ~x767 & ~x769 & ~x776;
assign c6273 =  x446;
assign c6275 =  x248 &  x611;
assign c6277 =  x14 &  x328 &  x344 &  x567 & ~x20 & ~x24 & ~x30 & ~x63 & ~x107 & ~x134 & ~x283 & ~x417 & ~x476 & ~x727;
assign c6279 = ~x91 & ~x118 & ~x166 & ~x201 & ~x339 & ~x368 & ~x618 & ~x623 & ~x680;
assign c6281 =  x139;
assign c6283 =  x153 &  x231 &  x236 &  x268 &  x324 &  x341 &  x397 &  x457 &  x460 &  x463 &  x541 &  x565 &  x621 &  x705 & ~x85 & ~x86 & ~x223 & ~x226 & ~x304 & ~x339 & ~x738 & ~x740 & ~x741 & ~x770;
assign c6285 = ~x65 & ~x229 & ~x258 & ~x287;
assign c6287 =  x457 &  x683 & ~x91 & ~x104 & ~x105;
assign c6289 =  x448;
assign c6291 = ~x271 & ~x299 & ~x300 & ~x609;
assign c6293 = ~x161 & ~x246 & ~x326 & ~x619;
assign c6295 = ~x400 & ~x401 & ~x452 & ~x664;
assign c6299 =  x211 &  x486 &  x544 &  x660 &  x779;
assign c6301 =  x444 &  x584 &  x639 &  x710;
assign c6303 =  x477;
assign c6305 =  x196;
assign c6307 =  x39 &  x399 &  x552 &  x566 & ~x105 & ~x249 & ~x311;
assign c6309 =  x70 &  x129 &  x210 &  x237 &  x243 &  x328 &  x381 &  x438 &  x441 &  x465 &  x546 &  x548 &  x605 &  x630 &  x634 &  x682 &  x711 &  x746 & ~x1 & ~x8 & ~x52 & ~x54 & ~x57 & ~x58 & ~x195 & ~x255 & ~x449 & ~x504 & ~x586 & ~x590 & ~x641 & ~x645 & ~x667 & ~x675 & ~x700;
assign c6311 = ~x52 & ~x109 & ~x171 & ~x335 & ~x401 & ~x423 & ~x452 & ~x479 & ~x537 & ~x733 & ~x754 & ~x755;
assign c6315 =  x139;
assign c6317 =  x172 &  x191 &  x219 & ~x566;
assign c6319 = ~x7 & ~x30 & ~x64 & ~x65 & ~x91 & ~x92 & ~x103 & ~x104 & ~x107 & ~x118 & ~x132 & ~x134 & ~x146 & ~x161 & ~x171 & ~x201 & ~x225 & ~x227 & ~x228 & ~x365 & ~x394 & ~x533 & ~x675 & ~x732;
assign c6321 =  x477;
assign c6323 =  x25 &  x756;
assign c6325 =  x599 &  x627 &  x633 &  x688 & ~x61 & ~x79 & ~x104 & ~x146 & ~x228 & ~x275 & ~x452 & ~x562 & ~x612 & ~x754;
assign c6327 =  x38 &  x155 &  x493 &  x597 & ~x623;
assign c6329 = ~x258 & ~x579 & ~x635 & ~x664 & ~x708 & ~x720;
assign c6331 =  x276 &  x304 &  x676;
assign c6335 =  x130 &  x357 &  x678 &  x706 & ~x115 & ~x503 & ~x585 & ~x714 & ~x715 & ~x716 & ~x742 & ~x747;
assign c6337 =  x497 &  x513 &  x553 & ~x5 & ~x53 & ~x91 & ~x92 & ~x104 & ~x105;
assign c6339 =  x1;
assign c6341 =  x70 &  x599 &  x737 &  x765 &  x766 &  x774 & ~x51 & ~x733;
assign c6343 =  x455 &  x526 & ~x92;
assign c6345 =  x475;
assign c6347 =  x44 &  x131 &  x190 &  x436 &  x457 &  x733 & ~x7 & ~x738 & ~x741 & ~x742 & ~x745 & ~x746;
assign c6349 =  x417;
assign c6351 =  x588;
assign c6353 =  x121 &  x145 &  x155 &  x218 &  x514 &  x550 &  x582 &  x621 &  x666 &  x694 & ~x613 & ~x769;
assign c6355 =  x128 &  x179 &  x209 & ~x117 & ~x146 & ~x246 & ~x330;
assign c6357 =  x781;
assign c6359 = ~x96 & ~x206 & ~x243 & ~x261;
assign c6361 =  x145 &  x211 &  x219 & ~x310 & ~x769;
assign c6363 =  x43 &  x119 &  x175 &  x183 &  x229 &  x313 &  x378 &  x433 &  x516 &  x694 &  x722 & ~x198 & ~x365 & ~x742 & ~x745 & ~x746 & ~x769 & ~x770;
assign c6365 =  x136;
assign c6367 =  x344 & ~x517;
assign c6369 =  x55;
assign c6373 = ~x120 & ~x177 & ~x216 & ~x316;
assign c6375 = ~x19 & ~x90 & ~x91 & ~x146 & ~x201 & ~x401;
assign c6377 =  x588;
assign c6379 =  x566 & ~x644 & ~x708 & ~x710 & ~x713 & ~x716 & ~x719 & ~x741 & ~x744 & ~x746 & ~x752 & ~x769;
assign c6381 = ~x261 & ~x288 & ~x693;
assign c6383 =  x38 &  x97 &  x121 &  x147 &  x291 &  x436 &  x578 &  x599 & ~x196 & ~x252 & ~x361 & ~x623 & ~x651 & ~x727;
assign c6385 =  x392;
assign c6387 =  x99 &  x122 &  x654 & ~x118 & ~x201 & ~x452 & ~x694;
assign c6389 = ~x69 & ~x119 & ~x210;
assign c6391 =  x764 &  x765 & ~x31 & ~x114;
assign c6393 =  x166;
assign c6395 = ~x201 & ~x260 & ~x271 & ~x272;
assign c6397 =  x464 & ~x65 & ~x91 & ~x92 & ~x103 & ~x104 & ~x120 & ~x146;
assign c6399 = ~x147 & ~x312 & ~x372 & ~x608 & ~x664;
assign c6401 =  x250;
assign c6403 =  x41 &  x70 &  x153 &  x175 &  x186 &  x205 &  x216 &  x231 &  x268 &  x358 &  x397 &  x425 &  x438 &  x439 &  x542 &  x565 &  x566 &  x583 &  x610 &  x611 &  x627 &  x632 &  x639 &  x649 &  x678 & ~x9 & ~x28 & ~x33 & ~x79 & ~x84 & ~x142 & ~x198 & ~x506 & ~x615 & ~x670;
assign c6405 =  x410 &  x494 &  x545 &  x547 &  x566 &  x581 & ~x52 & ~x91 & ~x105 & ~x671;
assign c6407 = ~x99 & ~x120 & ~x125 & ~x127 & ~x153 & ~x154 & ~x159 & ~x181;
assign c6409 =  x403 &  x766 & ~x693 & ~x694 & ~x706;
assign c6413 =  x11 &  x17 &  x130 &  x571 & ~x727;
assign c6415 =  x244 & ~x32 & ~x77 & ~x107 & ~x146 & ~x201 & ~x246 & ~x508 & ~x537 & ~x693;
assign c6417 =  x763;
assign c6419 =  x195;
assign c6421 =  x544 &  x600 & ~x19 & ~x33 & ~x64 & ~x75 & ~x79 & ~x91 & ~x104 & ~x117 & ~x142 & ~x146 & ~x164 & ~x783;
assign c6425 =  x756;
assign c6427 =  x757;
assign c6429 =  x229 &  x466 &  x662 &  x751 & ~x613 & ~x769 & ~x770;
assign c6431 =  x123 &  x151 &  x158 &  x205 &  x206 &  x241 &  x245 &  x261 &  x269 &  x375 &  x400 &  x405 &  x410 &  x522 &  x546 &  x547 &  x638 &  x649 &  x666 &  x705 & ~x220 & ~x337 & ~x363 & ~x388 & ~x586 & ~x725 & ~x769 & ~x770;
assign c6433 = ~x204 & ~x232 & ~x341 & ~x343 & ~x720 & ~x775;
assign c6435 =  x399 &  x522 &  x538 &  x606 & ~x47 & ~x105 & ~x146 & ~x586;
assign c6437 =  x54;
assign c6439 =  x14 &  x436 &  x550 &  x610 &  x678 & ~x50 & ~x77 & ~x134;
assign c6441 =  x479 &  x507 &  x675;
assign c6443 = ~x120 & ~x202 & ~x204 & ~x231;
assign c6445 =  x148 &  x175 &  x774 & ~x564 & ~x706;
assign c6447 =  x516 &  x553 & ~x0 & ~x76 & ~x91 & ~x104 & ~x107 & ~x118 & ~x138;
assign c6449 =  x477;
assign c6451 =  x252;
assign c6453 =  x77 &  x122 &  x191 &  x736 & ~x510 & ~x783;
assign c6455 =  x44 &  x379 &  x488 &  x525 &  x566 &  x654 & ~x18 & ~x91;
assign c6457 =  x728;
assign c6459 = ~x92 & ~x231 & ~x261;
assign c6461 =  x124 &  x145 &  x147 &  x236 &  x458 &  x509 &  x639 &  x663 &  x677 &  x723 &  x751;
assign c6463 =  x191 & ~x665 & ~x753;
assign c6465 =  x42 &  x106 & ~x566;
assign c6467 =  x44 &  x122 &  x187 &  x207 &  x322 &  x376 &  x379 &  x403 &  x433 &  x492 &  x516 &  x542 &  x602 & ~x9 & ~x56 & ~x138 & ~x168 & ~x305 & ~x340 & ~x365 & ~x415 & ~x589 & ~x693 & ~x724 & ~x780;
assign c6469 = ~x118 & ~x285 & ~x371 & ~x406;
assign c6471 = ~x127 & ~x409 & ~x435;
assign c6473 = ~x93 & ~x97 & ~x154 & ~x156 & ~x160;
assign c6475 =  x644;
assign c6477 =  x70 &  x94 &  x121 &  x124 &  x127 &  x129 &  x130 &  x131 &  x148 &  x159 &  x175 &  x179 &  x183 &  x203 &  x211 &  x212 &  x296 &  x353 &  x376 &  x379 &  x404 &  x460 &  x467 &  x493 &  x541 &  x606 &  x633 &  x681 &  x712 &  x740 &  x742 &  x747 &  x748 & ~x32 & ~x52 & ~x56 & ~x80 & ~x86 & ~x166 & ~x250 & ~x361 & ~x367 & ~x645 & ~x725;
assign c6479 =  x698;
assign c6481 =  x167;
assign c6483 = ~x65 & ~x67 & ~x92 & ~x97 & ~x98 & ~x120;
assign c6487 = ~x67 & ~x119 & ~x148 & ~x174 & ~x232;
assign c6489 =  x3;
assign c6491 =  x629 &  x654 &  x739 & ~x301 & ~x369 & ~x452 & ~x592;
assign c6493 =  x107 &  x192 & ~x370;
assign c6495 =  x778 & ~x745 & ~x752 & ~x769;
assign c6497 =  x251;
assign c6499 =  x72 &  x121 &  x130 &  x145 &  x173 &  x191 &  x201 &  x212 &  x219 &  x326 &  x352 &  x402 &  x626 &  x632 &  x748 & ~x502 & ~x642 & ~x698 & ~x759;
assign c70 = ~x301 & ~x440 & ~x655;
assign c74 =  x292 &  x318 & ~x88 & ~x648 & ~x708;
assign c76 =  x646;
assign c78 =  x214 & ~x47 & ~x50 & ~x54 & ~x78 & ~x89 & ~x119 & ~x134 & ~x255 & ~x280 & ~x290 & ~x335 & ~x369 & ~x598 & ~x600 & ~x703 & ~x704 & ~x707 & ~x712 & ~x717 & ~x732 & ~x739 & ~x760 & ~x763 & ~x773;
assign c710 =  x185 &  x296 &  x380 &  x415 &  x445 &  x486 &  x513 &  x521 &  x524 & ~x42 & ~x138 & ~x230 & ~x313 & ~x450 & ~x503 & ~x770;
assign c712 =  x614 &  x635 & ~x42 & ~x179 & ~x452 & ~x477;
assign c714 = ~x30 & ~x134 & ~x163 & ~x198 & ~x260 & ~x480 & ~x540 & ~x619 & ~x628 & ~x708 & ~x771;
assign c716 =  x482 &  x590 &  x632;
assign c718 =  x495 &  x559 &  x577 & ~x17 & ~x71 & ~x179 & ~x181 & ~x231 & ~x237 & ~x257 & ~x260 & ~x280 & ~x287 & ~x367 & ~x420 & ~x690 & ~x698;
assign c720 = ~x38 & ~x42 & ~x66 & ~x113 & ~x116 & ~x133 & ~x152 & ~x177 & ~x211 & ~x217 & ~x220 & ~x223 & ~x234 & ~x238 & ~x246 & ~x250 & ~x265 & ~x272 & ~x300 & ~x301 & ~x311 & ~x328 & ~x329 & ~x330 & ~x618 & ~x652 & ~x670 & ~x707;
assign c722 =  x386 &  x417 & ~x30 & ~x92 & ~x133 & ~x184 & ~x209 & ~x211 & ~x255 & ~x260 & ~x540 & ~x589 & ~x640 & ~x671 & ~x674 & ~x680 & ~x701 & ~x757;
assign c724 =  x403 &  x430 &  x516 &  x606 & ~x42 & ~x102 & ~x163 & ~x372 & ~x399;
assign c726 = ~x156 & ~x211 & ~x250 & ~x318 & ~x453 & ~x480 & ~x481 & ~x482 & ~x681 & ~x778;
assign c728 =  x215 &  x633 & ~x82 & ~x147 & ~x179 & ~x342 & ~x420 & ~x453;
assign c730 =  x587 & ~x45 & ~x193 & ~x680;
assign c732 = ~x44 & ~x78 & ~x133 & ~x164 & ~x185 & ~x454 & ~x586 & ~x707 & ~x729 & ~x769;
assign c734 =  x320 &  x321 &  x346 &  x372 & ~x30 & ~x31 & ~x33 & ~x47 & ~x82 & ~x86 & ~x134 & ~x139 & ~x144 & ~x163 & ~x164 & ~x198 & ~x231 & ~x252 & ~x253 & ~x309 & ~x503 & ~x619 & ~x622 & ~x637 & ~x648 & ~x664 & ~x726 & ~x757 & ~x758;
assign c736 = ~x30 & ~x133 & ~x209 & ~x260 & ~x293 & ~x347 & ~x399 & ~x453 & ~x596 & ~x605;
assign c738 =  x242 & ~x19 & ~x28 & ~x37 & ~x45 & ~x60 & ~x108 & ~x119 & ~x126 & ~x127 & ~x153 & ~x163 & ~x182 & ~x195 & ~x205 & ~x223 & ~x280 & ~x568 & ~x625 & ~x628 & ~x664 & ~x672 & ~x675 & ~x680 & ~x708 & ~x726 & ~x745 & ~x757 & ~x773 & ~x776;
assign c740 =  x325 &  x329 &  x331 &  x360 &  x403 &  x456 &  x457 &  x515 &  x520 & ~x8 & ~x23 & ~x31 & ~x34 & ~x71 & ~x89 & ~x179 & ~x229 & ~x252 & ~x259 & ~x280 & ~x284 & ~x309 & ~x315 & ~x318 & ~x339 & ~x343 & ~x397 & ~x398 & ~x424 & ~x588 & ~x615 & ~x646 & ~x664 & ~x698 & ~x704 & ~x759 & ~x782;
assign c742 =  x434 &  x578 & ~x42 & ~x54 & ~x57 & ~x59 & ~x70 & ~x119 & ~x124 & ~x144 & ~x173 & ~x175 & ~x179 & ~x235 & ~x619 & ~x626 & ~x636 & ~x749;
assign c744 =  x380 &  x458 &  x522 & ~x42 & ~x102 & ~x166 & ~x177 & ~x192 & ~x220 & ~x266 & ~x598 & ~x700 & ~x753;
assign c746 =  x293 &  x319 &  x372 & ~x221 & ~x246 & ~x619 & ~x625 & ~x655;
assign c748 =  x156 &  x332 & ~x643;
assign c750 =  x130 &  x243;
assign c752 =  x382 &  x436 &  x464 &  x471 &  x487 &  x496 &  x520 &  x521 & ~x31 & ~x49 & ~x68 & ~x97 & ~x107 & ~x116 & ~x125 & ~x135 & ~x203 & ~x211 & ~x223 & ~x267 & ~x316 & ~x363 & ~x641 & ~x656 & ~x671 & ~x708 & ~x719 & ~x727 & ~x739 & ~x749 & ~x763 & ~x766 & ~x768 & ~x779 & ~x781;
assign c754 =  x187 &  x301 &  x357 &  x418 &  x517 & ~x48 & ~x206 & ~x225 & ~x231 & ~x233 & ~x503 & ~x727 & ~x734;
assign c756 =  x349 &  x373 &  x403 &  x428 &  x456 &  x491 & ~x11 & ~x19 & ~x38 & ~x62 & ~x588 & ~x623 & ~x648 & ~x656 & ~x687 & ~x706 & ~x722 & ~x730 & ~x732 & ~x772;
assign c758 = ~x246 & ~x482 & ~x485;
assign c760 =  x382 &  x456 &  x484 &  x604 & ~x17 & ~x19 & ~x48 & ~x75 & ~x83 & ~x85 & ~x117 & ~x120 & ~x133 & ~x156 & ~x191 & ~x195 & ~x198 & ~x223 & ~x254 & ~x317 & ~x339 & ~x647 & ~x650 & ~x677 & ~x707 & ~x737 & ~x758;
assign c762 =  x186 &  x187 &  x358 &  x361 &  x606 & ~x47 & ~x290 & ~x338 & ~x345 & ~x643 & ~x766;
assign c764 =  x362 &  x379 &  x382 &  x439 &  x446 &  x462 &  x463 & ~x4 & ~x25 & ~x30 & ~x36 & ~x37 & ~x43 & ~x45 & ~x53 & ~x54 & ~x60 & ~x63 & ~x78 & ~x83 & ~x93 & ~x107 & ~x111 & ~x113 & ~x117 & ~x120 & ~x123 & ~x142 & ~x149 & ~x166 & ~x174 & ~x177 & ~x181 & ~x199 & ~x203 & ~x205 & ~x227 & ~x230 & ~x238 & ~x254 & ~x258 & ~x280 & ~x282 & ~x286 & ~x288 & ~x291 & ~x343 & ~x397 & ~x588 & ~x589 & ~x616 & ~x641 & ~x653 & ~x654 & ~x662 & ~x664 & ~x666 & ~x667 & ~x670 & ~x678 & ~x688 & ~x697 & ~x706 & ~x721 & ~x726 & ~x737 & ~x743 & ~x769;
assign c766 =  x402 &  x606 & ~x152 & ~x163 & ~x200 & ~x661;
assign c768 =  x211 &  x326 &  x474 &  x486 &  x541 &  x551 & ~x14 & ~x32 & ~x50 & ~x97 & ~x138 & ~x147 & ~x176 & ~x289 & ~x343 & ~x424 & ~x425 & ~x451 & ~x477 & ~x756;
assign c770 =  x242 &  x326 &  x332 &  x353 &  x382 &  x387 &  x388 &  x413 &  x483 &  x487 &  x551 & ~x41 & ~x43 & ~x44 & ~x45 & ~x50 & ~x78 & ~x86 & ~x129 & ~x133 & ~x134 & ~x135 & ~x152 & ~x160 & ~x220 & ~x221 & ~x255 & ~x317 & ~x367 & ~x370 & ~x448 & ~x698 & ~x704 & ~x705 & ~x708 & ~x714 & ~x750 & ~x756 & ~x758 & ~x761 & ~x766 & ~x769 & ~x775;
assign c772 = ~x163 & ~x164 & ~x480 & ~x481 & ~x511 & ~x625;
assign c774 =  x378 &  x379 &  x402 &  x406 &  x483 &  x578 & ~x6 & ~x31 & ~x42 & ~x45 & ~x52 & ~x75 & ~x76 & ~x80 & ~x83 & ~x108 & ~x157 & ~x190 & ~x335 & ~x616 & ~x652 & ~x655 & ~x698 & ~x727 & ~x771;
assign c776 = ~x23 & ~x29 & ~x33 & ~x38 & ~x42 & ~x44 & ~x47 & ~x53 & ~x62 & ~x67 & ~x68 & ~x85 & ~x96 & ~x99 & ~x104 & ~x105 & ~x106 & ~x113 & ~x125 & ~x126 & ~x130 & ~x134 & ~x142 & ~x144 & ~x162 & ~x182 & ~x196 & ~x198 & ~x223 & ~x260 & ~x290 & ~x317 & ~x337 & ~x372 & ~x392 & ~x426 & ~x454 & ~x563 & ~x599 & ~x644 & ~x669 & ~x678 & ~x695 & ~x708 & ~x711 & ~x721 & ~x741 & ~x748 & ~x758 & ~x760 & ~x781;
assign c778 =  x298 &  x380 &  x404 & ~x10 & ~x17 & ~x29 & ~x68 & ~x70 & ~x105 & ~x144 & ~x223 & ~x290 & ~x569 & ~x580 & ~x589 & ~x647 & ~x683 & ~x695 & ~x702 & ~x727 & ~x767 & ~x777;
assign c780 =  x605 &  x606 &  x609 & ~x2 & ~x14 & ~x18 & ~x32 & ~x42 & ~x53 & ~x57 & ~x58 & ~x102 & ~x104 & ~x158 & ~x160 & ~x168 & ~x174 & ~x222 & ~x228 & ~x230 & ~x233 & ~x287 & ~x288 & ~x308 & ~x363 & ~x681 & ~x691 & ~x704 & ~x708 & ~x731 & ~x746 & ~x779;
assign c782 =  x351 &  x384 &  x405 &  x408 & ~x23 & ~x28 & ~x41 & ~x43 & ~x69 & ~x83 & ~x88 & ~x114 & ~x119 & ~x129 & ~x142 & ~x154 & ~x165 & ~x198 & ~x201 & ~x227 & ~x316 & ~x448 & ~x598 & ~x664 & ~x671 & ~x757 & ~x769;
assign c784 =  x242 &  x430 &  x577 &  x578 & ~x193 & ~x628 & ~x688;
assign c786 =  x328 &  x362 &  x410 &  x413 &  x418 & ~x17 & ~x66 & ~x67 & ~x68 & ~x70 & ~x80 & ~x88 & ~x89 & ~x97 & ~x223 & ~x227 & ~x480 & ~x704 & ~x707;
assign c788 =  x244 &  x303 &  x353 &  x486 &  x497 & ~x2 & ~x12 & ~x20 & ~x44 & ~x47 & ~x58 & ~x67 & ~x69 & ~x97 & ~x114 & ~x125 & ~x135 & ~x193 & ~x226 & ~x289 & ~x293 & ~x313 & ~x370 & ~x396 & ~x420 & ~x451 & ~x677 & ~x687 & ~x696 & ~x704 & ~x707 & ~x731 & ~x773;
assign c790 =  x634 & ~x13 & ~x33 & ~x40 & ~x41 & ~x44 & ~x79 & ~x89 & ~x93 & ~x100 & ~x115 & ~x135 & ~x149 & ~x152 & ~x165 & ~x191 & ~x195 & ~x224 & ~x252 & ~x254 & ~x314 & ~x342 & ~x370 & ~x397 & ~x422 & ~x424 & ~x425 & ~x451 & ~x673 & ~x678 & ~x680 & ~x705 & ~x707 & ~x710 & ~x724 & ~x760 & ~x765 & ~x778;
assign c792 =  x532 &  x561 & ~x66 & ~x531;
assign c794 =  x375 &  x383 &  x384 & ~x30 & ~x47 & ~x86 & ~x116 & ~x528 & ~x600;
assign c796 =  x158 &  x474 & ~x44 & ~x230;
assign c798 =  x387 & ~x37 & ~x79 & ~x88 & ~x108 & ~x163 & ~x260 & ~x261 & ~x314 & ~x528 & ~x529 & ~x640 & ~x655 & ~x674 & ~x677 & ~x725 & ~x770 & ~x778;
assign c7100 =  x185 &  x239 &  x521 & ~x42 & ~x50 & ~x133 & ~x222 & ~x475 & ~x670 & ~x695 & ~x698 & ~x738 & ~x755;
assign c7102 =  x477 & ~x502;
assign c7104 =  x445 & ~x6 & ~x125 & ~x300;
assign c7106 =  x389 &  x494 & ~x7 & ~x14 & ~x23 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x47 & ~x52 & ~x71 & ~x72 & ~x83 & ~x117 & ~x227 & ~x251 & ~x283 & ~x287 & ~x316 & ~x345 & ~x363 & ~x451 & ~x480 & ~x481 & ~x701 & ~x730 & ~x757 & ~x758 & ~x764 & ~x768 & ~x769 & ~x780;
assign c7108 = ~x43 & ~x50 & ~x68 & ~x108 & ~x113 & ~x137 & ~x153 & ~x173 & ~x210 & ~x214 & ~x216 & ~x228 & ~x243 & ~x245 & ~x272 & ~x274 & ~x300 & ~x301 & ~x302 & ~x317 & ~x593 & ~x621 & ~x700 & ~x726 & ~x731 & ~x738 & ~x747;
assign c7110 =  x79;
assign c7112 =  x443 &  x456 &  x551 & ~x41 & ~x116 & ~x126 & ~x253 & ~x566 & ~x708;
assign c7114 =  x244 &  x246 &  x300 &  x355 &  x378 &  x382 &  x418 &  x463 &  x491 &  x492 &  x518 &  x563 &  x604 & ~x77 & ~x115 & ~x169 & ~x179 & ~x262 & ~x290 & ~x315 & ~x339 & ~x343 & ~x424 & ~x503 & ~x644 & ~x737 & ~x757;
assign c7116 =  x407 &  x463 & ~x42 & ~x66 & ~x126 & ~x133 & ~x210 & ~x250 & ~x501 & ~x625 & ~x695 & ~x711 & ~x753 & ~x758;
assign c7118 =  x368;
assign c7120 =  x633 &  x634 &  x637 & ~x73 & ~x264 & ~x344 & ~x374 & ~x739;
assign c7122 =  x550 & ~x246 & ~x300;
assign c7124 =  x434 &  x470 &  x487 &  x540 &  x541 & ~x41 & ~x53 & ~x147 & ~x206 & ~x226 & ~x307 & ~x315 & ~x370 & ~x480 & ~x677 & ~x765 & ~x778 & ~x779;
assign c7126 =  x159 &  x274 &  x471;
assign c7128 =  x326 &  x360 &  x434 &  x631 &  x632 &  x634 &  x635 & ~x54 & ~x95 & ~x174 & ~x176 & ~x230 & ~x288 & ~x290 & ~x339 & ~x343 & ~x344 & ~x373 & ~x392 & ~x399 & ~x426 & ~x450 & ~x452;
assign c7130 = ~x301 & ~x456 & ~x628;
assign c7132 =  x321 &  x375 &  x428 &  x456 &  x550 & ~x68 & ~x125 & ~x156 & ~x316 & ~x339 & ~x503;
assign c7134 =  x215 &  x389 &  x458 &  x516 & ~x36 & ~x41 & ~x51 & ~x70 & ~x97 & ~x101 & ~x108 & ~x226 & ~x267 & ~x286 & ~x316 & ~x338 & ~x369 & ~x448 & ~x695 & ~x700 & ~x707 & ~x714 & ~x722 & ~x745 & ~x748 & ~x783;
assign c7136 =  x292 &  x372;
assign c7138 = ~x337 & ~x511 & ~x512 & ~x636 & ~x757 & ~x774;
assign c7140 = ~x17 & ~x30 & ~x47 & ~x68 & ~x73 & ~x120 & ~x125 & ~x133 & ~x135 & ~x154 & ~x175 & ~x210 & ~x234 & ~x282 & ~x363 & ~x539 & ~x587 & ~x596 & ~x598 & ~x600 & ~x654 & ~x670 & ~x674 & ~x679 & ~x681 & ~x707 & ~x735 & ~x741 & ~x743 & ~x748 & ~x751;
assign c7142 =  x362 &  x469 &  x632 & ~x55 & ~x89 & ~x206 & ~x341 & ~x365 & ~x772 & ~x782;
assign c7144 = ~x189 & ~x226 & ~x451 & ~x482 & ~x596 & ~x628;
assign c7146 =  x321 &  x449 & ~x36 & ~x81 & ~x133 & ~x301 & ~x626;
assign c7148 =  x293 &  x320 &  x345 & ~x246 & ~x753;
assign c7150 =  x321 &  x347 &  x349 &  x373 &  x374 &  x429 &  x450 &  x456 & ~x13 & ~x41 & ~x42 & ~x45 & ~x126 & ~x144 & ~x205 & ~x589 & ~x642 & ~x700;
assign c7152 =  x422 &  x449 &  x451 &  x452 &  x483 & ~x54 & ~x244;
assign c7154 =  x349 &  x403 &  x429 &  x430 &  x445 & ~x36 & ~x42 & ~x51 & ~x54 & ~x163 & ~x195 & ~x628 & ~x666 & ~x675 & ~x682 & ~x695;
assign c7156 =  x423 & ~x66 & ~x245;
assign c7158 =  x297 &  x378 &  x414 &  x458 &  x462 &  x522 &  x555 &  x604 &  x606 & ~x0 & ~x5 & ~x8 & ~x69 & ~x93 & ~x163 & ~x191 & ~x201 & ~x226 & ~x237 & ~x255 & ~x369 & ~x373 & ~x732 & ~x749 & ~x750 & ~x765;
assign c7160 =  x577 &  x578 & ~x41 & ~x66 & ~x209 & ~x265 & ~x593 & ~x625 & ~x701 & ~x749;
assign c7162 =  x498 & ~x266 & ~x301 & ~x330;
assign c7164 =  x293 &  x319 &  x352 &  x375 &  x386 & ~x34 & ~x44 & ~x50 & ~x87 & ~x195 & ~x610 & ~x613 & ~x638 & ~x655 & ~x669 & ~x724 & ~x744 & ~x746 & ~x760;
assign c7166 =  x186 &  x418 &  x526 &  x577 &  x579 & ~x137 & ~x206 & ~x318;
assign c7168 =  x418 &  x491 & ~x272 & ~x301;
assign c7170 =  x379 & ~x503 & ~x543 & ~x544 & ~x545 & ~x625;
assign c7172 = ~x272 & ~x455;
assign c7174 =  x660;
assign c7176 =  x297 &  x323 &  x403 &  x484 &  x606 & ~x2 & ~x40 & ~x50 & ~x67 & ~x70 & ~x125 & ~x135 & ~x161 & ~x172 & ~x179 & ~x226 & ~x261 & ~x265 & ~x287 & ~x364 & ~x373 & ~x392 & ~x694 & ~x707 & ~x768 & ~x776;
assign c7178 =  x299 &  x327 &  x390 &  x483 &  x496 & ~x63 & ~x110 & ~x114 & ~x135 & ~x227 & ~x261 & ~x314 & ~x566 & ~x642 & ~x689 & ~x701 & ~x704 & ~x716 & ~x748 & ~x752 & ~x781;
assign c7180 =  x352 &  x362 &  x632 & ~x206 & ~x451 & ~x452;
assign c7182 = ~x510;
assign c7184 =  x349 &  x378 &  x403 &  x456 &  x491 & ~x15 & ~x42 & ~x45 & ~x54 & ~x64 & ~x69 & ~x76 & ~x107 & ~x116 & ~x121 & ~x134 & ~x136 & ~x149 & ~x171 & ~x178 & ~x217 & ~x265 & ~x396 & ~x503 & ~x738 & ~x750;
assign c7186 =  x379 &  x462 &  x575 &  x576 &  x577 &  x578 &  x579 & ~x4 & ~x7 & ~x16 & ~x17 & ~x19 & ~x28 & ~x30 & ~x31 & ~x33 & ~x38 & ~x40 & ~x43 & ~x46 & ~x69 & ~x73 & ~x95 & ~x96 & ~x119 & ~x123 & ~x131 & ~x132 & ~x133 & ~x135 & ~x154 & ~x160 & ~x164 & ~x168 & ~x177 & ~x207 & ~x209 & ~x222 & ~x223 & ~x228 & ~x258 & ~x282 & ~x284 & ~x291 & ~x392 & ~x448 & ~x588 & ~x589 & ~x616 & ~x619 & ~x633 & ~x637 & ~x643 & ~x647 & ~x660 & ~x677 & ~x680 & ~x682 & ~x695 & ~x697 & ~x707 & ~x711 & ~x722 & ~x743 & ~x745 & ~x748 & ~x753 & ~x756 & ~x770 & ~x775 & ~x779;
assign c7188 = ~x15 & ~x38 & ~x42 & ~x78 & ~x89 & ~x97 & ~x182 & ~x236 & ~x426 & ~x452 & ~x482 & ~x629 & ~x669 & ~x695 & ~x759;
assign c7190 =  x402 & ~x300 & ~x628;
assign c7192 =  x298 &  x411 &  x434 &  x444 & ~x12 & ~x14 & ~x15 & ~x17 & ~x31 & ~x37 & ~x38 & ~x47 & ~x49 & ~x63 & ~x77 & ~x99 & ~x116 & ~x125 & ~x154 & ~x156 & ~x161 & ~x163 & ~x174 & ~x189 & ~x208 & ~x209 & ~x224 & ~x251 & ~x259 & ~x261 & ~x279 & ~x286 & ~x313 & ~x578 & ~x587 & ~x619 & ~x634 & ~x638 & ~x683 & ~x698 & ~x700 & ~x708 & ~x711 & ~x768 & ~x776 & ~x780;
assign c7194 =  x349 &  x378 &  x403 &  x456 & ~x10 & ~x14 & ~x31 & ~x67 & ~x82 & ~x93 & ~x182 & ~x265 & ~x266 & ~x640 & ~x655 & ~x669 & ~x683 & ~x781;
assign c7196 =  x349 &  x403 &  x428 &  x429 & ~x125 & ~x153 & ~x205 & ~x259 & ~x282 & ~x335 & ~x556 & ~x636 & ~x643 & ~x651 & ~x671 & ~x724;
assign c7198 =  x158 &  x159 &  x186 &  x187;
assign c7200 =  x471 &  x483 &  x576 &  x578 & ~x60 & ~x67 & ~x68 & ~x135 & ~x164 & ~x166 & ~x179 & ~x198 & ~x211 & ~x220 & ~x225 & ~x284 & ~x641 & ~x698 & ~x761;
assign c7202 =  x470 & ~x134 & ~x142 & ~x177 & ~x190 & ~x191 & ~x219 & ~x272 & ~x328 & ~x619 & ~x654 & ~x680;
assign c7204 =  x403 &  x428 &  x578 & ~x265;
assign c7206 =  x158 &  x389 &  x471 &  x551 & ~x42 & ~x44 & ~x70 & ~x114 & ~x234 & ~x258 & ~x728 & ~x781;
assign c7208 =  x474 & ~x266 & ~x300 & ~x301;
assign c7210 =  x213 &  x380 & ~x42 & ~x73 & ~x77 & ~x116 & ~x217 & ~x451;
assign c7212 =  x215 &  x332 &  x352 &  x388 &  x517 & ~x12 & ~x23 & ~x24 & ~x96 & ~x116 & ~x139 & ~x154 & ~x157 & ~x178 & ~x182 & ~x183 & ~x225 & ~x315 & ~x318 & ~x370 & ~x393 & ~x423 & ~x451 & ~x693 & ~x707 & ~x712 & ~x728 & ~x731 & ~x732 & ~x750 & ~x759;
assign c7214 =  x491 &  x517 & ~x100 & ~x182 & ~x272 & ~x284 & ~x300 & ~x301 & ~x655 & ~x671 & ~x675 & ~x680 & ~x739 & ~x755;
assign c7216 =  x298 &  x332 &  x417 &  x550 & ~x75 & ~x126 & ~x178 & ~x266 & ~x267 & ~x373 & ~x680 & ~x695 & ~x724 & ~x749;
assign c7218 = ~x49 & ~x145 & ~x208 & ~x211 & ~x220 & ~x453 & ~x455 & ~x627 & ~x655 & ~x712;
assign c7220 =  x352 &  x402 &  x413 &  x428 &  x429 &  x456 &  x505 &  x524 & ~x27 & ~x44 & ~x64 & ~x78 & ~x125 & ~x126 & ~x139 & ~x152 & ~x153 & ~x154 & ~x161 & ~x217 & ~x340 & ~x448 & ~x617 & ~x643 & ~x671 & ~x680 & ~x709 & ~x716 & ~x722 & ~x733 & ~x741 & ~x764 & ~x773 & ~x779 & ~x781;
assign c7222 =  x455 &  x604 &  x606 & ~x119 & ~x182 & ~x424 & ~x647 & ~x698 & ~x749 & ~x768;
assign c7224 =  x301 &  x381 &  x384 &  x406 &  x418 & ~x14 & ~x15 & ~x35 & ~x60 & ~x128 & ~x147 & ~x195 & ~x229 & ~x364 & ~x596 & ~x607 & ~x636 & ~x696 & ~x758 & ~x772;
assign c7226 =  x664 & ~x374;
assign c7228 =  x293 &  x345 & ~x77 & ~x272 & ~x273;
assign c7230 =  x334 &  x362 &  x633 & ~x47 & ~x223 & ~x344;
assign c7232 = ~x344 & ~x511 & ~x512 & ~x598;
assign c7234 =  x242 &  x325 &  x326 &  x351 &  x361 &  x380 &  x384 &  x411 &  x418 &  x444 &  x461 &  x464 &  x519 &  x563 &  x604 &  x606 & ~x38 & ~x45 & ~x58 & ~x113 & ~x117 & ~x230 & ~x253 & ~x287 & ~x289 & ~x365 & ~x367 & ~x683 & ~x712 & ~x727 & ~x732 & ~x765;
assign c7236 =  x187 &  x472 &  x541 &  x579 &  x591 & ~x374 & ~x671;
assign c7238 =  x293 &  x319 &  x372 & ~x246 & ~x652 & ~x701 & ~x708 & ~x770;
assign c7240 = ~x300;
assign c7242 =  x357 &  x387 &  x500 &  x604 &  x605 &  x606 & ~x1 & ~x5 & ~x12 & ~x49 & ~x96 & ~x100 & ~x128 & ~x184 & ~x196 & ~x200 & ~x209 & ~x225 & ~x226 & ~x258 & ~x283 & ~x367 & ~x673;
assign c7244 = ~x474 & ~x495 & ~x616;
assign c7246 =  x663;
assign c7248 = ~x211 & ~x236 & ~x300 & ~x320 & ~x481;
assign c7250 =  x464 &  x577 &  x578 & ~x15 & ~x35 & ~x53 & ~x100 & ~x127 & ~x179 & ~x195 & ~x199 & ~x335 & ~x371 & ~x610 & ~x611 & ~x613 & ~x635 & ~x662 & ~x669 & ~x763 & ~x773 & ~x774;
assign c7252 =  x362 &  x384 & ~x105 & ~x156 & ~x266 & ~x504 & ~x597 & ~x628 & ~x728;
assign c7254 =  x444 & ~x46 & ~x73 & ~x86 & ~x92 & ~x129 & ~x153 & ~x182 & ~x185 & ~x186 & ~x191 & ~x211 & ~x212 & ~x219 & ~x230 & ~x244 & ~x245 & ~x259 & ~x272 & ~x284 & ~x300 & ~x301 & ~x307 & ~x593 & ~x595 & ~x598 & ~x611 & ~x616 & ~x618 & ~x729 & ~x735 & ~x749 & ~x757 & ~x769;
assign c7256 = ~x78 & ~x127 & ~x134 & ~x397 & ~x485 & ~x540 & ~x735 & ~x769;
assign c7258 =  x661;
assign c7260 =  x293 &  x319 &  x349 &  x372;
assign c7262 =  x418 & ~x275 & ~x301 & ~x596 & ~x598 & ~x617 & ~x619;
assign c7264 =  x349 &  x375 &  x402 &  x428 &  x460 &  x478 &  x483 & ~x8 & ~x42 & ~x45 & ~x46 & ~x55 & ~x59 & ~x66 & ~x87 & ~x89 & ~x116 & ~x133 & ~x135 & ~x136 & ~x142 & ~x152 & ~x154 & ~x161 & ~x165 & ~x190 & ~x226 & ~x309 & ~x310 & ~x336 & ~x339 & ~x589 & ~x619 & ~x631 & ~x641 & ~x655 & ~x670 & ~x677 & ~x695 & ~x708 & ~x719 & ~x723 & ~x726 & ~x737 & ~x743 & ~x763 & ~x768 & ~x770;
assign c7266 =  x186 &  x242 &  x298 &  x306 & ~x41 & ~x69 & ~x98 & ~x225 & ~x365 & ~x398 & ~x588;
assign c7268 = ~x328 & ~x544 & ~x545;
assign c7270 =  x559 & ~x15 & ~x163 & ~x679 & ~x708 & ~x735;
assign c7272 =  x382 &  x384 &  x411 &  x491 & ~x15 & ~x42 & ~x50 & ~x77 & ~x83 & ~x116 & ~x129 & ~x131 & ~x158 & ~x169 & ~x174 & ~x265 & ~x266 & ~x372 & ~x419 & ~x589 & ~x659 & ~x702;
assign c7274 =  x418 &  x470 &  x491 & ~x39 & ~x50 & ~x89 & ~x95 & ~x104 & ~x160 & ~x193 & ~x235 & ~x260 & ~x337 & ~x363 & ~x567 & ~x580 & ~x708 & ~x719 & ~x772;
assign c7276 =  x321 &  x345 &  x450;
assign c7278 = ~x50 & ~x96 & ~x153 & ~x482 & ~x483 & ~x628 & ~x681;
assign c7280 =  x386 &  x438 &  x491 & ~x79 & ~x134 & ~x139 & ~x164 & ~x195 & ~x217 & ~x253 & ~x314 & ~x397 & ~x596 & ~x616 & ~x693 & ~x749 & ~x761;
assign c7282 =  x270 &  x298 &  x349 &  x380 &  x403 &  x404 &  x410 &  x467 & ~x5 & ~x12 & ~x36 & ~x46 & ~x47 & ~x61 & ~x64 & ~x66 & ~x67 & ~x81 & ~x88 & ~x94 & ~x114 & ~x121 & ~x125 & ~x129 & ~x142 & ~x151 & ~x153 & ~x157 & ~x167 & ~x198 & ~x201 & ~x233 & ~x234 & ~x236 & ~x251 & ~x281 & ~x284 & ~x335 & ~x475 & ~x503 & ~x617 & ~x644 & ~x649 & ~x656 & ~x682 & ~x696 & ~x704 & ~x707 & ~x708 & ~x726 & ~x738 & ~x762 & ~x763;
assign c7284 =  x417 &  x461 & ~x75 & ~x86 & ~x152 & ~x217 & ~x226 & ~x256 & ~x370 & ~x423 & ~x566 & ~x641 & ~x680 & ~x687 & ~x695 & ~x708;
assign c7286 =  x319 &  x451 & ~x22 & ~x27 & ~x246 & ~x250 & ~x589 & ~x686;
assign c7288 =  x270 &  x355 &  x379 &  x380 &  x389 &  x404 &  x410 &  x445 &  x495 & ~x2 & ~x7 & ~x20 & ~x23 & ~x31 & ~x40 & ~x42 & ~x50 & ~x107 & ~x134 & ~x155 & ~x169 & ~x182 & ~x193 & ~x195 & ~x196 & ~x231 & ~x308 & ~x313 & ~x336 & ~x603 & ~x636 & ~x640 & ~x675 & ~x695 & ~x703 & ~x776;
assign c7290 =  x387 &  x440 &  x442 &  x477 &  x491 &  x521 & ~x15 & ~x42 & ~x54 & ~x58 & ~x66 & ~x78 & ~x105 & ~x108 & ~x114 & ~x126 & ~x130 & ~x133 & ~x134 & ~x136 & ~x159 & ~x211 & ~x225 & ~x226 & ~x229 & ~x235 & ~x252 & ~x337 & ~x366 & ~x397 & ~x619 & ~x634 & ~x638 & ~x695 & ~x708 & ~x753;
assign c7292 =  x186 &  x187 &  x354 &  x408 &  x442 &  x460 &  x468 & ~x26 & ~x51 & ~x230 & ~x279 & ~x311 & ~x337 & ~x339 & ~x392 & ~x559;
assign c7294 =  x418 & ~x220 & ~x250 & ~x272 & ~x300 & ~x301;
assign c7296 =  x461 &  x661 & ~x76 & ~x397 & ~x426;
assign c7298 = ~x220 & ~x250 & ~x290 & ~x440;
assign c7300 =  x403 &  x604 &  x606 & ~x453 & ~x503;
assign c7302 =  x130;
assign c7304 =  x293 &  x319 &  x320 &  x372 & ~x23 & ~x42 & ~x47 & ~x50 & ~x89 & ~x177 & ~x208 & ~x697;
assign c7306 =  x243 &  x483 &  x500 & ~x50 & ~x567 & ~x643;
assign c7308 = ~x473 & ~x497 & ~x521;
assign c7310 =  x332 &  x634 & ~x2 & ~x39 & ~x74 & ~x96 & ~x142 & ~x150 & ~x424 & ~x451 & ~x731 & ~x744 & ~x748 & ~x759 & ~x770;
assign c7312 = ~x300 & ~x511 & ~x512;
assign c7314 =  x422 &  x449 &  x451 &  x452 & ~x108 & ~x222 & ~x503;
assign c7316 = ~x17 & ~x501 & ~x521 & ~x599;
assign c7318 =  x349 &  x375 &  x402 &  x427 & ~x266 & ~x619 & ~x628;
assign c7320 =  x186 &  x243 & ~x23 & ~x41 & ~x47 & ~x57 & ~x96 & ~x227 & ~x641 & ~x678 & ~x695 & ~x697 & ~x700 & ~x732 & ~x768;
assign c7322 =  x325 &  x604 &  x605 &  x606 &  x607 & ~x2 & ~x13 & ~x15 & ~x24 & ~x31 & ~x36 & ~x40 & ~x68 & ~x76 & ~x84 & ~x86 & ~x92 & ~x117 & ~x137 & ~x147 & ~x149 & ~x162 & ~x166 & ~x190 & ~x195 & ~x200 & ~x201 & ~x227 & ~x229 & ~x230 & ~x337 & ~x372 & ~x448 & ~x642 & ~x643 & ~x654 & ~x656 & ~x658 & ~x674 & ~x675 & ~x682 & ~x701 & ~x731 & ~x742 & ~x751 & ~x758 & ~x766;
assign c7324 =  x449 & ~x160 & ~x217 & ~x220 & ~x272 & ~x330 & ~x628 & ~x723;
assign c7326 =  x380 &  x382 &  x417 &  x442 &  x460 & ~x1 & ~x4 & ~x7 & ~x14 & ~x17 & ~x21 & ~x33 & ~x43 & ~x48 & ~x53 & ~x74 & ~x82 & ~x83 & ~x86 & ~x89 & ~x102 & ~x111 & ~x115 & ~x123 & ~x127 & ~x139 & ~x149 & ~x150 & ~x165 & ~x178 & ~x194 & ~x196 & ~x230 & ~x231 & ~x232 & ~x258 & ~x311 & ~x314 & ~x337 & ~x343 & ~x372 & ~x397 & ~x425 & ~x532 & ~x587 & ~x644 & ~x649 & ~x669 & ~x686 & ~x703 & ~x716 & ~x721 & ~x749 & ~x753 & ~x762 & ~x763 & ~x764 & ~x770 & ~x777;
assign c7328 =  x243 &  x357 &  x379 &  x607 & ~x119 & ~x133 & ~x265 & ~x451 & ~x680 & ~x763;
assign c7330 =  x660 & ~x373 & ~x401 & ~x452;
assign c7332 =  x362 &  x475 & ~x12 & ~x17 & ~x43 & ~x167 & ~x279 & ~x366 & ~x586 & ~x747;
assign c7334 =  x327 &  x460 &  x487 & ~x35 & ~x266 & ~x398 & ~x566 & ~x651 & ~x697 & ~x773;
assign c7336 = ~x373 & ~x423 & ~x425 & ~x542 & ~x619;
assign c7338 = ~x96 & ~x134 & ~x156 & ~x198 & ~x206 & ~x230 & ~x261 & ~x342 & ~x453 & ~x480 & ~x481 & ~x664 & ~x671 & ~x738;
assign c7340 =  x532 &  x592;
assign c7342 =  x333;
assign c7344 =  x349 &  x362 &  x606 & ~x47 & ~x101 & ~x167 & ~x281 & ~x315 & ~x699 & ~x777;
assign c7346 = ~x81 & ~x133 & ~x163 & ~x250 & ~x481 & ~x482 & ~x485;
assign c7348 =  x266 &  x319 &  x345 & ~x665;
assign c7350 =  x213 &  x429 &  x456 &  x521 & ~x108 & ~x209 & ~x222 & ~x223 & ~x283 & ~x312 & ~x339 & ~x369 & ~x370 & ~x531 & ~x707 & ~x745 & ~x777;
assign c7352 =  x349 &  x578 & ~x42 & ~x66 & ~x184 & ~x191 & ~x230 & ~x642 & ~x684 & ~x691 & ~x777;
assign c7354 =  x470 & ~x37 & ~x133 & ~x156 & ~x157 & ~x208 & ~x211 & ~x221 & ~x224 & ~x248 & ~x250 & ~x265 & ~x272 & ~x300 & ~x301 & ~x589 & ~x593 & ~x598 & ~x616 & ~x626 & ~x628 & ~x637 & ~x707 & ~x741 & ~x757 & ~x770;
assign c7356 =  x423 &  x449 & ~x14 & ~x36 & ~x160 & ~x238 & ~x611 & ~x719 & ~x775;
assign c7358 = ~x49 & ~x96 & ~x164 & ~x251 & ~x495 & ~x500 & ~x501 & ~x596 & ~x707;
assign c7360 =  x321 &  x374 & ~x77 & ~x152 & ~x300 & ~x301 & ~x599 & ~x617 & ~x714 & ~x763;
assign c7362 = ~x17 & ~x47 & ~x89 & ~x146 & ~x217 & ~x301 & ~x482 & ~x561 & ~x615 & ~x635 & ~x695;
assign c7364 =  x269 &  x378 &  x380 &  x388 &  x404 &  x405 &  x408 &  x429 &  x430 &  x440 &  x456 &  x460 &  x483 &  x550 & ~x30 & ~x68 & ~x70 & ~x71 & ~x73 & ~x80 & ~x95 & ~x97 & ~x119 & ~x135 & ~x151 & ~x161 & ~x163 & ~x167 & ~x168 & ~x174 & ~x191 & ~x195 & ~x264 & ~x265 & ~x365 & ~x398 & ~x424 & ~x688 & ~x715 & ~x731 & ~x732 & ~x754 & ~x757 & ~x759 & ~x763;
assign c7366 =  x215 &  x418 &  x458 &  x562 &  x604 &  x606 & ~x12 & ~x112 & ~x260 & ~x364 & ~x367 & ~x450;
assign c7368 = ~x15 & ~x16 & ~x21 & ~x42 & ~x73 & ~x91 & ~x97 & ~x142 & ~x165 & ~x198 & ~x209 & ~x211 & ~x223 & ~x226 & ~x282 & ~x308 & ~x309 & ~x314 & ~x454 & ~x599 & ~x605 & ~x613 & ~x616 & ~x687 & ~x701 & ~x707 & ~x743;
assign c7370 =  x349 &  x418 &  x438 & ~x4 & ~x7 & ~x125 & ~x126 & ~x150 & ~x163 & ~x554 & ~x671 & ~x684 & ~x763;
assign c7372 =  x187 &  x242 &  x243 &  x331 &  x403 &  x429 &  x488 & ~x7 & ~x96 & ~x114 & ~x179 & ~x198 & ~x225 & ~x341 & ~x365 & ~x707 & ~x711 & ~x718 & ~x740 & ~x754 & ~x775;
assign c7374 =  x332 &  x474 &  x633 & ~x42 & ~x168 & ~x370 & ~x373 & ~x451 & ~x777;
assign c7376 = ~x163 & ~x452 & ~x501;
assign c7378 =  x186 &  x187 &  x302 &  x360 &  x418 & ~x8 & ~x12 & ~x50 & ~x421;
assign c7380 =  x326 &  x604 &  x606 & ~x220 & ~x619;
assign c7382 = ~x66 & ~x133 & ~x157 & ~x430 & ~x453 & ~x456 & ~x771;
assign c7384 = ~x440;
assign c7386 = ~x37 & ~x60 & ~x113 & ~x125 & ~x175 & ~x208 & ~x282 & ~x372 & ~x397 & ~x540 & ~x627 & ~x628 & ~x671 & ~x708 & ~x757;
assign c7388 =  x241 &  x242 &  x306 &  x357 & ~x38 & ~x66 & ~x152 & ~x208 & ~x223 & ~x341 & ~x370 & ~x426 & ~x448 & ~x451 & ~x756 & ~x776;
assign c7390 =  x471 &  x577 &  x578 & ~x0 & ~x3 & ~x29 & ~x30 & ~x36 & ~x42 & ~x143 & ~x150 & ~x156 & ~x164 & ~x182 & ~x190 & ~x193 & ~x195 & ~x260 & ~x307 & ~x308 & ~x561 & ~x624 & ~x660 & ~x671 & ~x680 & ~x688 & ~x736 & ~x739 & ~x762 & ~x770 & ~x780 & ~x782;
assign c7392 =  x215 & ~x12 & ~x47 & ~x57 & ~x148 & ~x163 & ~x169 & ~x205 & ~x209 & ~x222 & ~x229 & ~x284 & ~x289 & ~x321 & ~x347 & ~x368 & ~x616 & ~x710 & ~x772;
assign c7394 =  x362 &  x410 & ~x21 & ~x23 & ~x47 & ~x48 & ~x53 & ~x67 & ~x74 & ~x96 & ~x104 & ~x116 & ~x128 & ~x226 & ~x229 & ~x256 & ~x258 & ~x287 & ~x556 & ~x589 & ~x619 & ~x687 & ~x703 & ~x705 & ~x765 & ~x769;
assign c7396 =  x578 & ~x73 & ~x75 & ~x140 & ~x160 & ~x163 & ~x198 & ~x598;
assign c7398 =  x187 &  x326 &  x353 &  x354 &  x378 &  x379 &  x429 & ~x23 & ~x63 & ~x152 & ~x226 & ~x317 & ~x701 & ~x720 & ~x776;
assign c7400 =  x333 &  x362 &  x633 & ~x44 & ~x66 & ~x235 & ~x451;
assign c7402 =  x634 &  x635 &  x638 & ~x15 & ~x18 & ~x24 & ~x31 & ~x35 & ~x152 & ~x169 & ~x287 & ~x372 & ~x374 & ~x399;
assign c7404 =  x213 &  x277 &  x305 &  x333 &  x564 &  x623;
assign c7406 =  x384 & ~x37 & ~x217 & ~x523 & ~x529;
assign c7408 = ~x193 & ~x385 & ~x439;
assign c7410 =  x374 & ~x133 & ~x524;
assign c7412 =  x349 &  x374 &  x400 &  x441 &  x445 &  x455 & ~x9 & ~x125 & ~x313;
assign c7414 =  x349 &  x375 &  x383 &  x445 & ~x117 & ~x118 & ~x175 & ~x220 & ~x244 & ~x319 & ~x710;
assign c7416 =  x242 &  x387 &  x491 & ~x2 & ~x57 & ~x76 & ~x93 & ~x154 & ~x193 & ~x200 & ~x211 & ~x217 & ~x220 & ~x235 & ~x282 & ~x335 & ~x336 & ~x675 & ~x679 & ~x719 & ~x759 & ~x763;
assign c7418 = ~x42 & ~x272 & ~x454;
assign c7420 =  x379 &  x402 &  x491 &  x578 & ~x20 & ~x37 & ~x48 & ~x68 & ~x139 & ~x165 & ~x211 & ~x315 & ~x643 & ~x683 & ~x701 & ~x760 & ~x768;
assign c7422 =  x333 &  x384 &  x484 &  x549 &  x550 & ~x31 & ~x42 & ~x45 & ~x50 & ~x52 & ~x68 & ~x95 & ~x96 & ~x116 & ~x147 & ~x163 & ~x164 & ~x182 & ~x195 & ~x198 & ~x209 & ~x284 & ~x308 & ~x392 & ~x609 & ~x637 & ~x681 & ~x694 & ~x770;
assign c7424 = ~x220 & ~x222 & ~x272 & ~x300 & ~x301 & ~x328 & ~x356 & ~x711;
assign c7426 =  x440 &  x605 &  x606 & ~x74 & ~x109 & ~x116 & ~x150 & ~x158 & ~x176 & ~x193 & ~x260 & ~x373 & ~x392 & ~x616 & ~x641 & ~x679 & ~x721 & ~x769;
assign c7428 =  x158 &  x186 &  x189 &  x446 & ~x44 & ~x50 & ~x206 & ~x232 & ~x759;
assign c7430 =  x390 &  x474 & ~x89 & ~x134 & ~x266 & ~x321 & ~x451 & ~x614 & ~x778;
assign c7432 =  x186 &  x243 &  x514 & ~x13 & ~x220 & ~x222 & ~x695 & ~x760 & ~x782;
assign c7434 =  x293 &  x319 & ~x189 & ~x613 & ~x628 & ~x646 & ~x665 & ~x741 & ~x770 & ~x772;
assign c7436 = ~x35 & ~x113 & ~x116 & ~x133 & ~x246 & ~x265 & ~x342 & ~x424 & ~x453 & ~x589 & ~x671 & ~x770;
assign c7438 =  x158 &  x213 &  x242;
assign c7440 =  x242 &  x354 &  x388 &  x471 &  x508 & ~x29 & ~x42 & ~x50 & ~x152 & ~x162 & ~x163 & ~x182 & ~x222 & ~x262 & ~x337 & ~x448 & ~x616 & ~x695 & ~x712 & ~x736 & ~x738;
assign c7442 =  x321 &  x379 &  x400 &  x429 &  x451 &  x452 &  x477 & ~x14 & ~x40 & ~x45 & ~x60 & ~x79 & ~x103 & ~x108 & ~x144 & ~x160 & ~x619 & ~x746;
assign c7444 =  x215 &  x242 &  x244 &  x269 &  x417 &  x496 &  x538 &  x604 &  x605 &  x606 & ~x100 & ~x284 & ~x287 & ~x288 & ~x647 & ~x707;
assign c7446 = ~x42 & ~x209 & ~x223 & ~x453 & ~x510 & ~x651 & ~x695 & ~x708;
assign c7448 =  x144 &  x213;
assign c7450 = ~x32 & ~x423 & ~x426 & ~x453 & ~x481 & ~x485 & ~x773;
assign c7452 =  x634 & ~x132 & ~x135 & ~x345 & ~x618 & ~x649;
assign c7454 =  x518 &  x634 &  x637 & ~x182 & ~x222 & ~x397 & ~x707 & ~x739;
assign c7456 =  x471 & ~x47 & ~x113 & ~x133 & ~x163 & ~x190 & ~x228 & ~x236 & ~x282 & ~x539 & ~x540 & ~x561 & ~x595 & ~x619 & ~x626 & ~x640 & ~x708 & ~x712 & ~x725 & ~x726 & ~x758;
assign c7458 = ~x272 & ~x387 & ~x455;
assign c7460 =  x349 &  x428 &  x429 &  x456 &  x477 &  x490 & ~x11 & ~x70 & ~x77 & ~x102 & ~x116 & ~x126 & ~x147 & ~x156 & ~x170 & ~x194 & ~x223 & ~x265 & ~x287 & ~x632 & ~x655 & ~x681 & ~x707 & ~x708 & ~x713 & ~x728 & ~x769;
assign c7462 =  x332 &  x349 &  x380 &  x402 &  x404 &  x471 &  x483 &  x484 &  x491 &  x514 & ~x21 & ~x100 & ~x114 & ~x336 & ~x369 & ~x475 & ~x589 & ~x656 & ~x670 & ~x719 & ~x758;
assign c7464 =  x185 &  x522 & ~x45 & ~x119 & ~x137 & ~x144 & ~x152 & ~x182 & ~x209 & ~x261 & ~x503 & ~x531 & ~x723 & ~x737;
assign c7466 =  x380 &  x404 &  x429 &  x444 &  x456 &  x495 & ~x15 & ~x41 & ~x47 & ~x67 & ~x118 & ~x146 & ~x230 & ~x231 & ~x234 & ~x264 & ~x265 & ~x282 & ~x308 & ~x318 & ~x346 & ~x392 & ~x423 & ~x531 & ~x646 & ~x689 & ~x690 & ~x697 & ~x701 & ~x710 & ~x714 & ~x736 & ~x772;
assign c7468 =  x321 &  x373 &  x423 &  x426 & ~x58 & ~x88 & ~x100 & ~x137 & ~x153 & ~x200 & ~x207 & ~x227 & ~x315 & ~x699 & ~x704 & ~x712;
assign c7470 = ~x17 & ~x42 & ~x47 & ~x69 & ~x73 & ~x91 & ~x117 & ~x148 & ~x160 & ~x173 & ~x182 & ~x191 & ~x198 & ~x209 & ~x217 & ~x220 & ~x222 & ~x226 & ~x308 & ~x337 & ~x348 & ~x585 & ~x599 & ~x600 & ~x628 & ~x632 & ~x638 & ~x641 & ~x680 & ~x719;
assign c7472 =  x242 & ~x41 & ~x42 & ~x44 & ~x57 & ~x115 & ~x140 & ~x145 & ~x167 & ~x223 & ~x226 & ~x251 & ~x307 & ~x308 & ~x392 & ~x584 & ~x624 & ~x631 & ~x653 & ~x656 & ~x681 & ~x697 & ~x731 & ~x735 & ~x761;
assign c7474 =  x415 & ~x42 & ~x68 & ~x80 & ~x116 & ~x133 & ~x136 & ~x142 & ~x211 & ~x337 & ~x364 & ~x529 & ~x598 & ~x611 & ~x618 & ~x619 & ~x681 & ~x707 & ~x726 & ~x744 & ~x763 & ~x766;
assign c7476 =  x354 & ~x19 & ~x20 & ~x42 & ~x92 & ~x97 & ~x113 & ~x126 & ~x130 & ~x150 & ~x152 & ~x164 & ~x169 & ~x210 & ~x267 & ~x339 & ~x363 & ~x365 & ~x426 & ~x664 & ~x674 & ~x697 & ~x698 & ~x706;
assign c7478 = ~x31 & ~x80 & ~x95 & ~x116 & ~x134 & ~x163 & ~x182 & ~x203 & ~x211 & ~x265 & ~x282 & ~x294 & ~x392 & ~x399 & ~x447 & ~x453 & ~x454 & ~x705 & ~x707 & ~x721 & ~x758 & ~x762;
assign c7480 =  x293 &  x319 &  x372 &  x450 & ~x200 & ~x222 & ~x252 & ~x711 & ~x717;
assign c7482 =  x277 &  x293 &  x320 & ~x6 & ~x18 & ~x21 & ~x38 & ~x51 & ~x55 & ~x66 & ~x70 & ~x114 & ~x116 & ~x118 & ~x128 & ~x134 & ~x196 & ~x257 & ~x516 & ~x680 & ~x708 & ~x715 & ~x718 & ~x747 & ~x764 & ~x766 & ~x780 & ~x782;
assign c7484 =  x354 &  x419 & ~x364;
assign c7486 =  x375 & ~x32 & ~x156 & ~x163 & ~x191 & ~x226 & ~x282 & ~x543 & ~x544 & ~x708;
assign c7488 = ~x230 & ~x234 & ~x250 & ~x451 & ~x482 & ~x483 & ~x561 & ~x712;
assign c7490 =  x474 &  x518 &  x550 & ~x23 & ~x33 & ~x36 & ~x49 & ~x73 & ~x96 & ~x106 & ~x136 & ~x137 & ~x140 & ~x192 & ~x193 & ~x222 & ~x266 & ~x292 & ~x367 & ~x642 & ~x644 & ~x684 & ~x690 & ~x697 & ~x703 & ~x734 & ~x754 & ~x770 & ~x772 & ~x773 & ~x783;
assign c7492 =  x403 &  x428 &  x578 & ~x236 & ~x338 & ~x589;
assign c7494 =  x269 &  x405 &  x418 & ~x54 & ~x56 & ~x120 & ~x203 & ~x307 & ~x335 & ~x582 & ~x616 & ~x619 & ~x636 & ~x640 & ~x668 & ~x724;
assign c7496 =  x382 &  x386 & ~x21 & ~x24 & ~x56 & ~x57 & ~x79 & ~x92 & ~x106 & ~x114 & ~x127 & ~x133 & ~x135 & ~x157 & ~x165 & ~x178 & ~x195 & ~x207 & ~x209 & ~x223 & ~x227 & ~x233 & ~x371 & ~x397 & ~x420 & ~x531 & ~x557 & ~x615 & ~x616 & ~x617 & ~x643 & ~x680 & ~x692 & ~x695 & ~x708 & ~x712 & ~x730 & ~x757 & ~x759 & ~x767;
assign c7498 =  x402 &  x403 &  x456 &  x477 & ~x49 & ~x86 & ~x120 & ~x126 & ~x134 & ~x182 & ~x210 & ~x251 & ~x264 & ~x317 & ~x503 & ~x589 & ~x645 & ~x653 & ~x655 & ~x671 & ~x674 & ~x687 & ~x724;
assign c71 =  x282;
assign c73 =  x220 &  x537 &  x569 &  x584 & ~x659;
assign c75 =  x235;
assign c77 = ~x248 & ~x276 & ~x305 & ~x395 & ~x418 & ~x443 & ~x445 & ~x446 & ~x564 & ~x586 & ~x610 & ~x641;
assign c79 =  x105;
assign c711 =  x330 & ~x349 & ~x406 & ~x408;
assign c713 =  x425 & ~x389;
assign c715 =  x42;
assign c717 =  x295 &  x473 &  x584 &  x585 &  x612 &  x613 & ~x280 & ~x659;
assign c719 =  x207;
assign c721 = ~x404 & ~x405 & ~x432 & ~x433 & ~x461;
assign c723 =  x151;
assign c725 =  x233;
assign c727 =  x584 &  x611 & ~x634;
assign c729 =  x643;
assign c731 =  x369;
assign c733 = ~x5 & ~x7 & ~x24 & ~x28 & ~x53 & ~x150 & ~x286 & ~x390 & ~x394 & ~x396 & ~x417 & ~x418 & ~x559 & ~x562 & ~x586 & ~x599 & ~x611 & ~x630 & ~x640 & ~x681 & ~x743 & ~x758;
assign c735 =  x697;
assign c737 =  x221 &  x584 & ~x186;
assign c739 =  x453 & ~x417 & ~x418 & ~x576;
assign c741 =  x124;
assign c743 = ~x31 & ~x102 & ~x406 & ~x407 & ~x463 & ~x633 & ~x688 & ~x711;
assign c745 =  x191;
assign c747 =  x756;
assign c749 =  x696;
assign c751 =  x135;
assign c753 =  x612;
assign c755 = ~x145 & ~x251 & ~x268 & ~x270 & ~x274 & ~x276 & ~x305 & ~x334 & ~x395 & ~x506 & ~x535 & ~x548 & ~x551 & ~x556 & ~x579 & ~x582 & ~x661;
assign c757 =  x312;
assign c759 = ~x35 & ~x123 & ~x241 & ~x268 & ~x269 & ~x270 & ~x271 & ~x390 & ~x535 & ~x546 & ~x550 & ~x575 & ~x578 & ~x586;
assign c761 = ~x241 & ~x268 & ~x269 & ~x270 & ~x305 & ~x333 & ~x390 & ~x541 & ~x547 & ~x564 & ~x581;
assign c763 = ~x85 & ~x305 & ~x333 & ~x334 & ~x361 & ~x362 & ~x389 & ~x390 & ~x506 & ~x507 & ~x532 & ~x538 & ~x558 & ~x563 & ~x586 & ~x610;
assign c765 =  x220 &  x501 &  x537 &  x584 &  x594 &  x596 &  x611 & ~x159 & ~x717 & ~x724;
assign c767 =  x408 & ~x390 & ~x418 & ~x445;
assign c769 =  x533 &  x545 & ~x334;
assign c771 =  x176;
assign c773 =  x397 &  x425 & ~x390;
assign c775 =  x249 &  x546 &  x613 & ~x655;
assign c777 =  x50;
assign c781 =  x231;
assign c783 =  x248 &  x479 &  x506 &  x572;
assign c785 =  x537 & ~x407 & ~x449;
assign c787 = ~x350 & ~x352 & ~x380 & ~x463 & ~x464;
assign c791 =  x249 &  x501 &  x506 &  x534 &  x571 &  x572 & ~x347 & ~x659;
assign c793 =  x221 &  x247 &  x248 &  x249 &  x295 &  x466 &  x545 &  x569 &  x571 &  x585;
assign c795 =  x310;
assign c797 =  x425 &  x454 & ~x133 & ~x269 & ~x270 & ~x271 & ~x338 & ~x665;
assign c799 =  x466 & ~x390 & ~x415 & ~x417 & ~x418;
assign c7101 = ~x305 & ~x333 & ~x361 & ~x386 & ~x388 & ~x389 & ~x582;
assign c7105 = ~x293 & ~x405 & ~x406 & ~x407 & ~x435 & ~x463 & ~x606;
assign c7109 =  x137;
assign c7111 =  x603 &  x656;
assign c7113 =  x69;
assign c7115 =  x315;
assign c7117 =  x533 &  x584 & ~x401;
assign c7119 =  x335;
assign c7121 =  x651;
assign c7123 =  x506 &  x584 &  x593 &  x596 & ~x634;
assign c7125 =  x42;
assign c7127 =  x219 &  x612 & ~x159;
assign c7129 =  x39;
assign c7131 =  x145;
assign c7133 = ~x333 & ~x334 & ~x390 & ~x395 & ~x413 & ~x579 & ~x645;
assign c7135 =  x92;
assign c7137 =  x667;
assign c7139 =  x221 &  x641;
assign c7141 =  x682;
assign c7143 =  x137;
assign c7145 =  x248 &  x271 &  x540 &  x548 &  x584 &  x585;
assign c7147 =  x647;
assign c7149 =  x233;
assign c7151 =  x42;
assign c7153 =  x651;
assign c7155 =  x247 &  x248 &  x533 &  x556 &  x571 &  x585;
assign c7157 =  x13;
assign c7159 =  x183 &  x585;
assign c7161 =  x277 &  x356 &  x359 &  x479 &  x480 &  x489 &  x506 &  x511 &  x512 &  x528 &  x545 &  x571 &  x583 &  x584 &  x585 & ~x746;
assign c7163 =  x240 &  x268 &  x272 &  x533 &  x567 &  x582 &  x584 &  x595 &  x611 & ~x449;
assign c7165 =  x282;
assign c7167 =  x163;
assign c7169 =  x246 &  x586 & ~x306 & ~x428;
assign c7171 =  x233;
assign c7173 =  x783;
assign c7175 =  x46;
assign c7177 =  x596 &  x613 &  x641 & ~x663;
assign c7179 =  x557 & ~x269 & ~x690;
assign c7181 =  x219 &  x582 &  x611;
assign c7183 =  x360 & ~x249 & ~x390 & ~x417 & ~x418 & ~x443 & ~x444 & ~x445 & ~x446 & ~x752;
assign c7185 =  x205;
assign c7187 =  x69;
assign c7189 =  x44;
assign c7191 =  x122;
assign c7193 =  x260;
assign c7195 =  x248 &  x479 &  x480 &  x506 & ~x399;
assign c7197 = ~x297 & ~x305 & ~x339 & ~x361 & ~x548 & ~x549 & ~x563;
assign c7199 =  x235;
assign c7201 =  x425 & ~x3 & ~x130 & ~x154 & ~x270 & ~x535 & ~x552 & ~x574 & ~x597 & ~x609 & ~x667 & ~x674 & ~x733;
assign c7203 =  x466 & ~x390 & ~x415 & ~x417 & ~x418;
assign c7205 =  x275 &  x276 &  x277 &  x509 &  x537 &  x544 &  x554 &  x570 &  x571 & ~x98 & ~x117 & ~x592 & ~x603 & ~x622 & ~x623 & ~x628 & ~x631 & ~x673 & ~x776;
assign c7207 =  x622 &  x640 &  x651;
assign c7209 =  x537 &  x543 &  x556 &  x557 &  x567 &  x568 &  x570 &  x585 & ~x219 & ~x606 & ~x702;
assign c7211 =  x233;
assign c7213 =  x312;
assign c7215 =  x231;
assign c7217 =  x739;
assign c7219 =  x126;
assign c7221 =  x219 &  x569 &  x611;
assign c7223 =  x95;
assign c7225 =  x235;
assign c7227 =  x710;
assign c7229 =  x315;
assign c7231 =  x327 &  x433 &  x506 &  x507 &  x525 &  x538 &  x543 &  x545 &  x585 & ~x606;
assign c7233 =  x283;
assign c7235 =  x235;
assign c7237 =  x397 & ~x152 & ~x241 & ~x278 & ~x334 & ~x559;
assign c7239 = ~x305 & ~x389 & ~x492;
assign c7241 =  x312;
assign c7243 = ~x284 & ~x387 & ~x389 & ~x390;
assign c7245 = ~x59 & ~x81 & ~x406 & ~x407 & ~x434 & ~x435 & ~x462;
assign c7247 = ~x406 & ~x435 & ~x463;
assign c7249 =  x275 &  x322 &  x356 &  x416 &  x466 &  x479 &  x480 &  x506 &  x533 &  x536 &  x557 &  x568 & ~x74 & ~x623;
assign c7251 =  x736;
assign c7253 =  x248 &  x493 &  x556 &  x611;
assign c7255 =  x466 & ~x99 & ~x269 & ~x270 & ~x290 & ~x389 & ~x390 & ~x652;
assign c7257 =  x249 &  x506 &  x511 &  x546 & ~x214;
assign c7259 = ~x316 & ~x406 & ~x407 & ~x463 & ~x464 & ~x690;
assign c7261 =  x684;
assign c7263 =  x206;
assign c7265 =  x221 &  x602 &  x641;
assign c7267 =  x247 &  x612;
assign c7269 =  x247 & ~x333 & ~x402;
assign c7271 =  x310;
assign c7273 =  x193 &  x585;
assign c7275 =  x289;
assign c7277 =  x207;
assign c7279 =  x398 & ~x241 & ~x269 & ~x390;
assign c7281 =  x98;
assign c7283 =  x489 & ~x418 & ~x445 & ~x446;
assign c7285 =  x221 &  x247 &  x248 &  x585;
assign c7287 =  x585 &  x649 &  x651;
assign c7289 =  x235;
assign c7291 =  x397 & ~x222 & ~x240 & ~x241 & ~x262 & ~x269 & ~x311 & ~x313 & ~x700 & ~x771;
assign c7293 = ~x90 & ~x333 & ~x354 & ~x361 & ~x552 & ~x577;
assign c7295 =  x44;
assign c7297 =  x626 &  x653;
assign c7299 = ~x305 & ~x306 & ~x334 & ~x417 & ~x418 & ~x422 & ~x423 & ~x442 & ~x443 & ~x444 & ~x446 & ~x564 & ~x586 & ~x640 & ~x775;
assign c7301 = ~x406 & ~x407 & ~x435 & ~x436 & ~x463;
assign c7303 =  x279;
assign c7307 =  x683;
assign c7309 =  x260;
assign c7311 =  x695;
assign c7313 =  x335 & ~x382;
assign c7315 =  x220 &  x593 &  x612;
assign c7317 = ~x305 & ~x332 & ~x333 & ~x361 & ~x507;
assign c7319 =  x315;
assign c7321 =  x772;
assign c7323 =  x248 &  x506 & ~x187 & ~x660 & ~x690;
assign c7325 =  x600 &  x628 &  x655;
assign c7327 =  x194;
assign c7329 =  x204;
assign c7331 =  x370 & ~x394 & ~x396 & ~x417;
assign c7333 =  x116;
assign c7337 =  x611 &  x624;
assign c7339 =  x248 &  x501 &  x533 &  x557 &  x568 &  x585 &  x613;
assign c7341 = ~x417 & ~x444 & ~x445 & ~x576;
assign c7343 =  x248 &  x546 &  x557 & ~x18 & ~x371 & ~x606;
assign c7345 = ~x354 & ~x519;
assign c7347 = ~x83 & ~x406 & ~x407 & ~x435 & ~x436 & ~x463 & ~x464 & ~x689;
assign c7349 = ~x277 & ~x305 & ~x306 & ~x313 & ~x332 & ~x333 & ~x359 & ~x366 & ~x478;
assign c7351 =  x256;
assign c7353 = ~x26 & ~x147 & ~x172 & ~x309 & ~x332 & ~x333 & ~x338 & ~x360 & ~x361 & ~x386 & ~x394 & ~x504 & ~x564 & ~x614 & ~x701 & ~x715 & ~x780;
assign c7355 =  x179;
assign c7357 =  x669;
assign c7359 =  x258;
assign c7361 =  x453 & ~x268 & ~x269 & ~x270 & ~x390 & ~x551 & ~x552;
assign c7363 = ~x28 & ~x86 & ~x143 & ~x191 & ~x271 & ~x276 & ~x418 & ~x443 & ~x444 & ~x445 & ~x446 & ~x535 & ~x559 & ~x563 & ~x577 & ~x580 & ~x637 & ~x642 & ~x751;
assign c7365 =  x770;
assign c7367 =  x258;
assign c7369 =  x600 &  x624 &  x628 &  x655;
assign c7371 = ~x240 & ~x269 & ~x270 & ~x284 & ~x305 & ~x362 & ~x389 & ~x390 & ~x549 & ~x558;
assign c7373 = ~x193 & ~x240 & ~x248 & ~x389 & ~x390 & ~x541 & ~x551 & ~x558 & ~x564 & ~x581 & ~x663 & ~x693 & ~x720 & ~x779;
assign c7375 =  x163;
assign c7377 =  x257;
assign c7379 =  x234;
assign c7381 =  x457 & ~x32 & ~x61 & ~x240 & ~x270 & ~x306 & ~x394 & ~x417 & ~x418 & ~x576 & ~x656;
assign c7383 =  x336;
assign c7385 =  x249 &  x611 & ~x455;
assign c7387 = ~x406 & ~x407 & ~x421 & ~x422 & ~x433 & ~x435 & ~x449 & ~x751;
assign c7391 =  x289;
assign c7393 =  x313;
assign c7395 = ~x248 & ~x390 & ~x417 & ~x418 & ~x420 & ~x423 & ~x433 & ~x639 & ~x751;
assign c7397 =  x260;
assign c7399 =  x668;
assign c7401 = ~x305 & ~x330 & ~x333 & ~x358 & ~x361 & ~x362 & ~x385 & ~x386 & ~x388 & ~x389 & ~x390 & ~x505 & ~x559;
assign c7403 =  x683;
assign c7405 =  x506 &  x527 &  x583 &  x596 &  x611 & ~x532;
assign c7407 =  x57;
assign c7409 = ~x29 & ~x107 & ~x117 & ~x122 & ~x128 & ~x212 & ~x215 & ~x234 & ~x258 & ~x307 & ~x337 & ~x389 & ~x390 & ~x417 & ~x418 & ~x563 & ~x577 & ~x583 & ~x611 & ~x618 & ~x624 & ~x632 & ~x657 & ~x682 & ~x749 & ~x763;
assign c7411 =  x165;
assign c7413 = ~x205 & ~x251 & ~x389 & ~x390 & ~x416 & ~x417 & ~x418 & ~x577 & ~x581 & ~x616 & ~x730 & ~x774;
assign c7415 =  x583 &  x594 &  x626;
assign c7417 =  x126;
assign c7419 = ~x352 & ~x353 & ~x422 & ~x423 & ~x451;
assign c7421 =  x763;
assign c7423 =  x466 & ~x417 & ~x443 & ~x446;
assign c7425 =  x42;
assign c7427 =  x119;
assign c7429 =  x45;
assign c7431 =  x221 &  x585;
assign c7433 =  x234;
assign c7435 =  x669;
assign c7437 =  x359 &  x511 & ~x241 & ~x271 & ~x445 & ~x576;
assign c7439 = ~x3 & ~x30 & ~x62 & ~x196 & ~x252 & ~x282 & ~x324 & ~x325 & ~x352 & ~x353 & ~x354 & ~x381 & ~x382 & ~x691 & ~x708 & ~x780;
assign c7441 = ~x34 & ~x50 & ~x56 & ~x64 & ~x91 & ~x173 & ~x253 & ~x263 & ~x305 & ~x333 & ~x361 & ~x386 & ~x389 & ~x390 & ~x558 & ~x560 & ~x564 & ~x586 & ~x733 & ~x759;
assign c7443 = ~x350 & ~x352;
assign c7445 =  x217 &  x218 &  x570 & ~x375 & ~x740;
assign c7447 =  x247 &  x248 &  x506 &  x553 &  x584 & ~x400;
assign c7449 =  x309;
assign c7451 = ~x361;
assign c7453 =  x602 &  x611 &  x627 &  x651;
assign c7455 =  x398 & ~x269 & ~x270;
assign c7457 =  x285;
assign c7459 =  x285;
assign c7461 =  x585;
assign c7463 =  x133;
assign c7465 = ~x131 & ~x241 & ~x257 & ~x258 & ~x269 & ~x270 & ~x339 & ~x390 & ~x538 & ~x549 & ~x552 & ~x553 & ~x560 & ~x571 & ~x573 & ~x587 & ~x601 & ~x604;
assign c7467 =  x567 &  x613;
assign c7469 = ~x296 & ~x325 & ~x326 & ~x333 & ~x353 & ~x476;
assign c7471 =  x648;
assign c7473 =  x710;
assign c7475 =  x154;
assign c7477 =  x397 &  x425 & ~x268;
assign c7479 =  x249 &  x533 &  x556 &  x585;
assign c7481 =  x39;
assign c7483 =  x247 &  x248 &  x506 &  x546 & ~x428;
assign c7485 =  x725;
assign c7487 =  x315;
assign c7489 =  x260;
assign c7491 =  x267 &  x479 &  x506 &  x537 &  x566 &  x567 &  x584 &  x585;
assign c7493 = ~x215 & ~x241 & ~x242 & ~x270 & ~x390 & ~x417 & ~x418 & ~x574 & ~x751 & ~x771;
assign c7495 =  x479 &  x506 &  x556 &  x567 &  x568 &  x583 &  x584 &  x585 & ~x601;
assign c7497 =  x258;
assign c7499 =  x191 &  x585;
assign c80 = ~x100 & ~x456 & ~x485;
assign c82 = ~x45 & ~x187 & ~x217 & ~x271 & ~x273 & ~x345 & ~x349;
assign c84 =  x321 &  x323 &  x382 &  x384 & ~x651 & ~x666;
assign c86 = ~x157 & ~x272 & ~x299 & ~x301 & ~x302 & ~x323 & ~x328 & ~x441;
assign c88 =  x572 & ~x37 & ~x299 & ~x403 & ~x413;
assign c810 =  x448;
assign c812 =  x315 &  x533 & ~x218;
assign c814 = ~x45 & ~x76 & ~x126 & ~x266 & ~x267 & ~x440;
assign c816 = ~x45 & ~x239 & ~x265 & ~x267 & ~x293 & ~x294 & ~x296 & ~x316 & ~x320 & ~x321 & ~x324;
assign c818 =  x421 &  x562;
assign c820 =  x301 &  x354 & ~x510 & ~x540 & ~x624;
assign c822 =  x308;
assign c824 =  x437 &  x524 & ~x159 & ~x190;
assign c826 =  x500 & ~x101 & ~x127 & ~x682 & ~x684 & ~x685 & ~x692 & ~x714;
assign c828 =  x766 & ~x355;
assign c830 =  x5;
assign c832 = ~x455 & ~x486 & ~x540 & ~x541 & ~x570 & ~x623 & ~x651 & ~x679;
assign c834 = ~x467 & ~x468 & ~x470 & ~x485 & ~x486 & ~x487 & ~x496 & ~x522;
assign c836 = ~x98 & ~x155 & ~x305;
assign c838 =  x546 &  x635 &  x714 &  x716 &  x720 &  x734 &  x736 &  x742 & ~x228;
assign c840 =  x289 &  x293 &  x300 &  x384 & ~x657 & ~x665;
assign c842 =  x691 &  x766 & ~x62 & ~x105;
assign c844 =  x234 & ~x513 & ~x653 & ~x680;
assign c846 =  x502 &  x524 & ~x738;
assign c848 =  x152 & ~x684;
assign c850 =  x635 & ~x75 & ~x134 & ~x238;
assign c852 =  x659 &  x717 & ~x16 & ~x29 & ~x37 & ~x65 & ~x74 & ~x88 & ~x93 & ~x103 & ~x120 & ~x121 & ~x127 & ~x144 & ~x146 & ~x157 & ~x160 & ~x173 & ~x178 & ~x190 & ~x219 & ~x222 & ~x757;
assign c854 =  x392;
assign c856 = ~x426 & ~x428 & ~x442 & ~x519 & ~x526;
assign c858 =  x400 &  x523 &  x545 & ~x132 & ~x175 & ~x723 & ~x750;
assign c860 =  x356 &  x384 &  x501 & ~x39;
assign c862 =  x365;
assign c864 =  x336;
assign c866 =  x112;
assign c868 =  x447;
assign c870 =  x343 &  x400 &  x401 &  x523 &  x524 &  x545 &  x609 & ~x76 & ~x753;
assign c872 =  x290 &  x318 &  x345 &  x353 &  x427 &  x467 &  x519 &  x523 &  x524 &  x525 &  x552 &  x608 &  x636 &  x637 &  x651 &  x677 &  x685 &  x691 &  x692 &  x693 &  x714;
assign c874 =  x383 & ~x127 & ~x240 & ~x266 & ~x267;
assign c876 =  x51;
assign c878 = ~x347 & ~x463 & ~x486 & ~x494 & ~x498 & ~x513;
assign c880 = ~x10 & ~x38 & ~x217 & ~x238 & ~x243 & ~x272;
assign c882 =  x49 &  x50 &  x161;
assign c884 =  x326 &  x539 &  x608 &  x712 &  x714 &  x715 &  x716 &  x717 &  x718 &  x719 &  x740 &  x741 &  x743 &  x744 &  x745;
assign c886 =  x287 &  x348 &  x400 &  x427 &  x428 &  x456 &  x510 &  x511 &  x668 &  x677 &  x688 &  x693 &  x706;
assign c888 =  x51;
assign c890 =  x365;
assign c892 = ~x24 & ~x78 & ~x98 & ~x131 & ~x133 & ~x204 & ~x266 & ~x267 & ~x273 & ~x728;
assign c894 =  x634 &  x717 &  x741 &  x743 & ~x190 & ~x442 & ~x470 & ~x615;
assign c896 = ~x466 & ~x468 & ~x485 & ~x487 & ~x498 & ~x515;
assign c898 =  x552 &  x689 &  x690 &  x695 &  x706;
assign c8100 = ~x101;
assign c8102 =  x335;
assign c8104 =  x419;
assign c8106 =  x561;
assign c8108 =  x717 &  x734;
assign c8110 =  x334 & ~x627 & ~x679 & ~x685;
assign c8112 =  x55;
assign c8114 = ~x98 & ~x455 & ~x463 & ~x466 & ~x484;
assign c8116 =  x290 & ~x132 & ~x177 & ~x190 & ~x218;
assign c8118 = ~x39 & ~x45 & ~x154 & ~x233 & ~x246 & ~x265 & ~x293 & ~x329;
assign c8120 =  x325 &  x345 &  x348 &  x350 &  x351 &  x354 &  x372 &  x382 &  x436 &  x437 & ~x91 & ~x750 & ~x752 & ~x782;
assign c8122 =  x596 & ~x36 & ~x148 & ~x202 & ~x219 & ~x239 & ~x262 & ~x363;
assign c8124 =  x51 &  x315;
assign c8126 =  x263 &  x328 &  x361 &  x472 & ~x76;
assign c8128 =  x281 & ~x693;
assign c8130 =  x756;
assign c8132 =  x300 &  x318 &  x333 &  x356 &  x501;
assign c8134 =  x137;
assign c8136 =  x263 & ~x542 & ~x569 & ~x710;
assign c8138 =  x221 &  x290 &  x361 &  x622;
assign c8140 =  x764 & ~x70;
assign c8142 =  x561 & ~x246;
assign c8144 =  x521 &  x744 & ~x75;
assign c8146 =  x211 &  x236 &  x247 &  x329 &  x379 &  x524 &  x525 &  x637 &  x684 & ~x251 & ~x338 & ~x647;
assign c8148 =  x384 &  x401 &  x428 &  x539 &  x636 & ~x64 & ~x130 & ~x775;
assign c8150 =  x3;
assign c8152 = ~x10 & ~x50 & ~x103 & ~x118 & ~x188 & ~x204 & ~x219 & ~x246 & ~x260 & ~x267 & ~x272 & ~x274 & ~x293 & ~x295 & ~x301 & ~x729;
assign c8154 = ~x37 & ~x62 & ~x107 & ~x135 & ~x164 & ~x375 & ~x383 & ~x410 & ~x486 & ~x585;
assign c8156 =  x372 &  x719 & ~x145 & ~x388;
assign c8158 =  x371 &  x501;
assign c8160 =  x634 &  x660 &  x661 &  x685 &  x691 & ~x17 & ~x19 & ~x37 & ~x219 & ~x246 & ~x274 & ~x393 & ~x588;
assign c8162 =  x504;
assign c8164 =  x137 &  x639;
assign c8166 =  x227 &  x620;
assign c8168 = ~x98 & ~x314 & ~x409 & ~x426 & ~x435;
assign c8170 =  x511 &  x512 &  x522 & ~x266;
assign c8172 =  x49 &  x95 &  x213 &  x318 &  x688 & ~x643 & ~x673;
assign c8174 =  x280;
assign c8176 =  x783;
assign c8178 =  x560;
assign c8182 =  x432 &  x523 &  x545 &  x546 &  x549 & ~x66 & ~x77 & ~x133 & ~x154 & ~x155 & ~x190 & ~x777;
assign c8184 =  x282 & ~x103 & ~x656 & ~x686 & ~x735;
assign c8186 = ~x16 & ~x23 & ~x30 & ~x36 & ~x47 & ~x55 & ~x62 & ~x63 & ~x64 & ~x75 & ~x76 & ~x78 & ~x90 & ~x98 & ~x104 & ~x105 & ~x114 & ~x118 & ~x121 & ~x126 & ~x133 & ~x141 & ~x162 & ~x196 & ~x197 & ~x200 & ~x223 & ~x227 & ~x394 & ~x502 & ~x615;
assign c8188 =  x478 & ~x63;
assign c8190 =  x309 & ~x190;
assign c8192 =  x716 &  x717 &  x740 &  x741 &  x743 &  x744 & ~x17 & ~x64 & ~x120 & ~x133 & ~x146 & ~x174 & ~x190 & ~x196;
assign c8194 =  x691 & ~x238 & ~x266;
assign c8196 = ~x39 & ~x45 & ~x98 & ~x126 & ~x153 & ~x268 & ~x652 & ~x657 & ~x709 & ~x710;
assign c8198 =  x365;
assign c8200 =  x299 &  x321 &  x496 &  x524 & ~x102;
assign c8202 =  x447;
assign c8204 =  x159 & ~x597;
assign c8206 =  x281 & ~x132;
assign c8208 = ~x428 & ~x442 & ~x455 & ~x456 & ~x463 & ~x466 & ~x469;
assign c8210 = ~x106 & ~x343 & ~x375 & ~x383 & ~x440 & ~x457;
assign c8212 =  x165 &  x261;
assign c8214 =  x220 &  x398 &  x499 &  x637 &  x639 & ~x199;
assign c8216 =  x337;
assign c8218 =  x315 &  x399 &  x400 &  x459 & ~x692 & ~x699 & ~x710 & ~x720 & ~x729 & ~x749 & ~x750;
assign c8220 =  x429 &  x467 &  x514 &  x524 & ~x10 & ~x154 & ~x217;
assign c8222 = ~x121 & ~x243 & ~x271 & ~x273 & ~x293 & ~x300 & ~x301 & ~x469 & ~x498;
assign c8224 =  x429 &  x679 &  x732;
assign c8226 =  x281;
assign c8228 = ~x719;
assign c8230 =  x691 &  x718 & ~x98;
assign c8232 =  x364;
assign c8234 =  x344 &  x399 &  x428 &  x524 &  x596 &  x636 &  x692 &  x719 & ~x76 & ~x445 & ~x472;
assign c8236 = ~x36 & ~x46 & ~x92 & ~x98 & ~x155 & ~x240 & ~x273 & ~x275 & ~x293 & ~x294 & ~x295 & ~x296;
assign c8238 =  x298 &  x676 &  x694;
assign c8240 =  x196;
assign c8242 =  x427 &  x678 &  x705 &  x716;
assign c8244 = ~x441 & ~x457 & ~x485 & ~x486 & ~x510 & ~x515 & ~x522;
assign c8246 =  x263 &  x427 &  x501 &  x609;
assign c8248 =  x54;
assign c8250 =  x576 & ~x93 & ~x98 & ~x270 & ~x273;
assign c8252 =  x742 &  x766 & ~x87 & ~x134 & ~x218 & ~x470;
assign c8254 = ~x594 & ~x595;
assign c8256 =  x766 & ~x266 & ~x274;
assign c8258 =  x548 & ~x36 & ~x76 & ~x104 & ~x120 & ~x122 & ~x137 & ~x159 & ~x190 & ~x229 & ~x237 & ~x244;
assign c8260 =  x657 & ~x210 & ~x265 & ~x273;
assign c8262 =  x345 &  x390 &  x500 & ~x107;
assign c8264 =  x5;
assign c8266 =  x300 &  x384 & ~x654 & ~x683 & ~x684 & ~x711 & ~x722;
assign c8268 = ~x133 & ~x162 & ~x218 & ~x302 & ~x330 & ~x333 & ~x656 & ~x681;
assign c8270 =  x152 &  x399 &  x427 &  x428 &  x525 & ~x38 & ~x44 & ~x46 & ~x64 & ~x66 & ~x74;
assign c8272 = ~x39 & ~x107 & ~x133 & ~x134 & ~x187 & ~x210 & ~x217 & ~x331;
assign c8274 =  x766 & ~x76 & ~x77 & ~x119 & ~x133 & ~x176 & ~x215 & ~x243 & ~x265;
assign c8276 =  x113;
assign c8278 = ~x126 & ~x265 & ~x273 & ~x300 & ~x357 & ~x442;
assign c8280 =  x278 & ~x680 & ~x734 & ~x737;
assign c8282 =  x644;
assign c8284 =  x363;
assign c8286 =  x3;
assign c8288 =  x523 & ~x176 & ~x217 & ~x267;
assign c8290 =  x714 & ~x265 & ~x287 & ~x293;
assign c8292 =  x109 &  x611;
assign c8294 =  x398 &  x521 &  x663 & ~x212 & ~x266;
assign c8296 = ~x298 & ~x349 & ~x351 & ~x358;
assign c8298 =  x474 & ~x98 & ~x709;
assign c8300 =  x734 & ~x126 & ~x133;
assign c8302 =  x138;
assign c8304 =  x260 &  x276 &  x427 &  x677 & ~x37;
assign c8306 =  x393 &  x611;
assign c8308 =  x290 &  x433 & ~x712 & ~x733;
assign c8310 =  x1;
assign c8312 =  x196;
assign c8316 =  x364;
assign c8318 =  x137;
assign c8320 =  x605 &  x687 &  x718 & ~x244 & ~x273;
assign c8322 =  x273 &  x399 &  x499 &  x609 &  x637 &  x691 &  x692 &  x693 &  x695 &  x720;
assign c8324 =  x270 & ~x541 & ~x691;
assign c8326 = ~x154 & ~x182 & ~x189 & ~x265 & ~x274 & ~x302 & ~x331 & ~x441;
assign c8328 =  x290 &  x345 &  x411 & ~x3 & ~x7 & ~x651 & ~x655 & ~x656 & ~x666 & ~x680 & ~x684 & ~x694 & ~x702 & ~x705 & ~x721 & ~x768;
assign c8330 =  x177 &  x220 &  x354 &  x528 &  x581;
assign c8332 =  x14 &  x400 &  x624 & ~x71;
assign c8334 =  x224;
assign c8336 =  x282 & ~x679;
assign c8340 = ~x45 & ~x118 & ~x132 & ~x133 & ~x266 & ~x273;
assign c8342 = ~x99 & ~x133 & ~x399 & ~x628 & ~x679 & ~x685;
assign c8344 = ~x331;
assign c8346 =  x24;
assign c8348 = ~x539 & ~x540 & ~x626 & ~x627 & ~x677 & ~x681 & ~x706 & ~x710 & ~x779;
assign c8350 = ~x11 & ~x294 & ~x378 & ~x380;
assign c8354 =  x332 &  x398 & ~x93;
assign c8356 =  x14 &  x775 & ~x91;
assign c8358 = ~x78 & ~x242 & ~x265 & ~x269 & ~x272 & ~x274 & ~x299 & ~x300 & ~x329 & ~x441 & ~x444;
assign c8360 = ~x37 & ~x244 & ~x294 & ~x299 & ~x318;
assign c8362 =  x263 &  x264 &  x293 & ~x624 & ~x645 & ~x655 & ~x728;
assign c8364 =  x334 &  x351 &  x501 & ~x42 & ~x736;
assign c8366 =  x428 &  x717 & ~x132 & ~x203;
assign c8368 =  x461 &  x467 &  x579 & ~x76 & ~x155 & ~x182 & ~x752;
assign c8370 =  x336;
assign c8372 =  x263 &  x299 &  x356 & ~x569;
assign c8374 =  x384 &  x524 &  x691 &  x716 & ~x134 & ~x173;
assign c8376 =  x428 &  x474 &  x581 & ~x39;
assign c8378 =  x309 & ~x99;
assign c8380 =  x433 &  x436 &  x495 &  x523 &  x578 & ~x45 & ~x130;
assign c8382 =  x559;
assign c8384 =  x398 &  x429 &  x648 &  x687 &  x707;
assign c8386 =  x690 & ~x17 & ~x39 & ~x76 & ~x98 & ~x157 & ~x185 & ~x239;
assign c8388 =  x476;
assign c8390 = ~x65 & ~x71 & ~x245 & ~x471 & ~x482 & ~x510 & ~x526;
assign c8392 =  x338 & ~x146;
assign c8394 =  x427 &  x717 & ~x17 & ~x76 & ~x121;
assign c8396 =  x411 &  x461 &  x523 &  x551 & ~x10 & ~x29 & ~x34 & ~x36 & ~x45 & ~x92 & ~x120 & ~x133 & ~x279 & ~x304 & ~x756;
assign c8398 =  x336;
assign c8400 =  x532;
assign c8402 =  x315 &  x390;
assign c8404 =  x524 &  x569 & ~x10 & ~x99 & ~x182 & ~x267 & ~x269 & ~x448 & ~x477;
assign c8406 =  x432 &  x433 & ~x512 & ~x541 & ~x627 & ~x739;
assign c8408 =  x260 &  x298 &  x676 &  x691 &  x705;
assign c8410 =  x756;
assign c8412 = ~x69 & ~x99 & ~x115 & ~x119 & ~x132 & ~x189 & ~x190 & ~x200 & ~x204 & ~x210 & ~x226 & ~x246 & ~x267 & ~x294 & ~x331;
assign c8414 =  x308;
assign c8416 = ~x265 & ~x300 & ~x302 & ~x349 & ~x441 & ~x468 & ~x498;
assign c8418 =  x197;
assign c8420 = ~x99 & ~x110 & ~x127 & ~x455 & ~x588 & ~x609 & ~x654 & ~x663 & ~x680;
assign c8422 = ~x271;
assign c8424 =  x315 &  x334;
assign c8426 =  x263 &  x277 &  x385 &  x611 & ~x226;
assign c8428 =  x52;
assign c8430 =  x511 &  x690 & ~x76 & ~x98 & ~x133;
assign c8432 =  x759;
assign c8434 =  x714 & ~x103 & ~x358 & ~x414;
assign c8436 =  x718 & ~x10 & ~x210 & ~x754;
assign c8438 =  x168;
assign c8440 =  x3;
assign c8442 =  x79 &  x400 &  x678;
assign c8444 =  x356 & ~x569 & ~x628 & ~x667;
assign c8446 =  x694 &  x734 &  x766;
assign c8448 =  x223;
assign c8450 = ~x103 & ~x133 & ~x265 & ~x442 & ~x498;
assign c8452 =  x574 &  x577 &  x604 &  x687 &  x689 & ~x92 & ~x104 & ~x313;
assign c8454 =  x112;
assign c8456 =  x51 &  x66;
assign c8458 =  x438 & ~x76 & ~x99 & ~x103 & ~x161 & ~x164 & ~x240;
assign c8460 =  x308;
assign c8462 =  x14 &  x734 &  x743 &  x766;
assign c8464 = ~x218 & ~x271 & ~x272 & ~x345 & ~x441 & ~x442 & ~x469;
assign c8466 =  x677 &  x764;
assign c8468 =  x112;
assign c8470 =  x347 &  x411 & ~x49 & ~x99 & ~x133 & ~x197 & ~x421 & ~x588;
assign c8472 =  x427 &  x705 &  x722 &  x736 &  x738;
assign c8474 =  x79 &  x528;
assign c8476 =  x337;
assign c8478 = ~x513 & ~x569 & ~x710;
assign c8480 =  x400 &  x494 &  x519 &  x541 & ~x215 & ~x752;
assign c8482 =  x300 & ~x25 & ~x706 & ~x710 & ~x719 & ~x738;
assign c8484 =  x718 &  x735 & ~x92;
assign c8486 =  x514 &  x550 &  x601 & ~x240 & ~x301;
assign c8488 =  x137;
assign c8490 = ~x154 & ~x265 & ~x294 & ~x407 & ~x441;
assign c8492 =  x560;
assign c8494 =  x223;
assign c8496 =  x625 & ~x27 & ~x38 & ~x46 & ~x93 & ~x105 & ~x132 & ~x148 & ~x155 & ~x175 & ~x204 & ~x210 & ~x212 & ~x218 & ~x241;
assign c8498 =  x276 &  x401 &  x524 &  x691 &  x706 & ~x698;
assign c81 =  x748 & ~x307 & ~x453 & ~x482 & ~x509 & ~x528 & ~x620 & ~x675;
assign c83 =  x64 &  x652 & ~x80 & ~x588 & ~x620 & ~x667 & ~x675 & ~x700 & ~x703 & ~x729;
assign c85 =  x238 &  x266 &  x463 & ~x3 & ~x113 & ~x198 & ~x282 & ~x366 & ~x398;
assign c87 = ~x292 & ~x340 & ~x423 & ~x747;
assign c89 = ~x42 & ~x137 & ~x152 & ~x180 & ~x186 & ~x234 & ~x235 & ~x258 & ~x262 & ~x365 & ~x633 & ~x636 & ~x648 & ~x659 & ~x717 & ~x732 & ~x745;
assign c811 = ~x23 & ~x49 & ~x53 & ~x170 & ~x198 & ~x199 & ~x222 & ~x225 & ~x227 & ~x283 & ~x360 & ~x393 & ~x423 & ~x446 & ~x451 & ~x475 & ~x501 & ~x530 & ~x534 & ~x535 & ~x559 & ~x585 & ~x644 & ~x647 & ~x675 & ~x699 & ~x703 & ~x725 & ~x729 & ~x748 & ~x765;
assign c813 =  x40 &  x41 &  x42 &  x43 & ~x90 & ~x556;
assign c815 =  x64 &  x485 & ~x111 & ~x113 & ~x196 & ~x564 & ~x588 & ~x620;
assign c817 =  x69 &  x70 &  x594 & ~x23 & ~x49 & ~x366 & ~x474;
assign c819 =  x172 &  x228 & ~x29 & ~x505 & ~x761;
assign c821 = ~x33 & ~x234 & ~x262 & ~x337 & ~x339 & ~x562 & ~x591 & ~x606 & ~x633 & ~x661 & ~x662 & ~x689 & ~x748;
assign c823 = ~x166 & ~x213 & ~x235 & ~x236 & ~x544;
assign c825 =  x444 & ~x234 & ~x337 & ~x340;
assign c827 =  x444 & ~x635 & ~x636 & ~x663;
assign c829 = ~x14 & ~x283 & ~x304 & ~x311 & ~x359 & ~x368 & ~x400 & ~x508 & ~x530 & ~x620;
assign c831 =  x187 &  x215 &  x243 &  x485 &  x486 &  x492 &  x606 &  x623 &  x655 &  x656 &  x658 & ~x13 & ~x26 & ~x528 & ~x585 & ~x647 & ~x668 & ~x697 & ~x703;
assign c833 =  x101 &  x156 &  x157 &  x158 &  x182 &  x187 &  x217 &  x339 &  x396 &  x486 &  x656 &  x662 & ~x762;
assign c835 = ~x205 & ~x227 & ~x235 & ~x236 & ~x291 & ~x368 & ~x420 & ~x689 & ~x727 & ~x777;
assign c837 =  x698;
assign c839 =  x103 &  x118 &  x163 &  x199 &  x229 &  x303 & ~x53 & ~x224;
assign c841 =  x463 &  x736 & ~x5 & ~x31 & ~x52 & ~x366 & ~x368 & ~x370 & ~x388 & ~x396 & ~x418 & ~x474 & ~x500 & ~x509 & ~x583 & ~x585 & ~x588 & ~x590 & ~x620 & ~x675;
assign c843 =  x40 &  x69 & ~x23 & ~x112 & ~x139 & ~x166 & ~x193 & ~x199 & ~x220 & ~x280 & ~x308 & ~x310 & ~x361 & ~x478 & ~x502;
assign c845 =  x45 & ~x194 & ~x393 & ~x450 & ~x508 & ~x509 & ~x583 & ~x592 & ~x614;
assign c847 =  x397 &  x564 &  x751 & ~x112 & ~x419;
assign c849 =  x346 & ~x0 & ~x109 & ~x255 & ~x338 & ~x411 & ~x474 & ~x505 & ~x533 & ~x559 & ~x562;
assign c851 = ~x234 & ~x254 & ~x311 & ~x366 & ~x393 & ~x493 & ~x501;
assign c853 =  x453 & ~x180 & ~x575;
assign c855 =  x126 &  x127 &  x131 &  x150 &  x156 &  x187 &  x201 &  x202 &  x203 &  x204 &  x206 &  x210 &  x215 &  x230 &  x240 &  x241 &  x242 &  x258 &  x296 &  x313 &  x358 &  x368 &  x378 &  x397 &  x571 & ~x334;
assign c857 =  x65 &  x103 &  x158 &  x210 &  x257 &  x396 &  x598 & ~x80 & ~x588;
assign c859 =  x15 &  x68 &  x71 &  x98 & ~x49 & ~x80 & ~x168 & ~x251 & ~x279;
assign c861 = ~x163 & ~x186 & ~x207 & ~x234 & ~x543 & ~x562;
assign c863 =  x296 &  x324 &  x409 &  x437 &  x749 & ~x28 & ~x280 & ~x451 & ~x499 & ~x500 & ~x504 & ~x505 & ~x535 & ~x559 & ~x585 & ~x613 & ~x675;
assign c865 =  x445 &  x454 & ~x82 & ~x110 & ~x142 & ~x235 & ~x282 & ~x289 & ~x336 & ~x690 & ~x757 & ~x783;
assign c867 = ~x43 & ~x199 & ~x200 & ~x234 & ~x262 & ~x285 & ~x288 & ~x336 & ~x338 & ~x341 & ~x688 & ~x703 & ~x717 & ~x767;
assign c869 = ~x326 & ~x505 & ~x507 & ~x509 & ~x535 & ~x563 & ~x583;
assign c871 = ~x398 & ~x501 & ~x502 & ~x525;
assign c873 =  x295 &  x486 &  x598 & ~x14 & ~x86 & ~x501 & ~x530 & ~x534 & ~x535 & ~x560 & ~x611 & ~x612 & ~x616 & ~x781;
assign c875 = ~x326 & ~x353 & ~x523;
assign c877 =  x530 & ~x290 & ~x340;
assign c879 =  x349 & ~x143 & ~x368 & ~x508 & ~x525 & ~x554;
assign c881 = ~x227 & ~x232 & ~x284 & ~x311 & ~x562 & ~x603 & ~x631 & ~x703;
assign c883 =  x452 &  x453 &  x482 & ~x14 & ~x24 & ~x221 & ~x562 & ~x647;
assign c885 =  x268 &  x746 & ~x14 & ~x42 & ~x54 & ~x168 & ~x613;
assign c887 = ~x14 & ~x28 & ~x197 & ~x201 & ~x252 & ~x261 & ~x316 & ~x339 & ~x340 & ~x396 & ~x425 & ~x449 & ~x783;
assign c889 =  x296 &  x515 & ~x113 & ~x536 & ~x583 & ~x729;
assign c891 =  x171 &  x248 &  x305 &  x691;
assign c893 = ~x14 & ~x199 & ~x205 & ~x208 & ~x234 & ~x286 & ~x290 & ~x311 & ~x366 & ~x765;
assign c895 =  x453 & ~x14 & ~x21 & ~x50 & ~x590 & ~x633 & ~x735;
assign c897 =  x242 &  x598 &  x627 & ~x22 & ~x113 & ~x224 & ~x474 & ~x583 & ~x668 & ~x675 & ~x676;
assign c899 =  x157 &  x210 &  x303 &  x585 &  x619 &  x640 &  x641 & ~x84 & ~x109 & ~x420;
assign c8101 = ~x280 & ~x311 & ~x339 & ~x340 & ~x384 & ~x397 & ~x562;
assign c8103 =  x410 & ~x152 & ~x262 & ~x281 & ~x311 & ~x317 & ~x765;
assign c8105 =  x41 &  x42 &  x43 &  x44 & ~x87 & ~x225 & ~x279 & ~x335 & ~x367 & ~x388 & ~x530 & ~x535 & ~x585 & ~x619 & ~x647;
assign c8107 = ~x234 & ~x532 & ~x566 & ~x591 & ~x600 & ~x605 & ~x613 & ~x689;
assign c8109 =  x612 & ~x203 & ~x368 & ~x424;
assign c8111 =  x201 &  x231 &  x284 &  x313 &  x360 &  x396 &  x545 & ~x81 & ~x137 & ~x278 & ~x363;
assign c8113 =  x16 &  x42 & ~x253;
assign c8115 =  x506 &  x507 & ~x227 & ~x286 & ~x366 & ~x395;
assign c8117 =  x184 &  x360 &  x591 &  x619 &  x640 &  x641 & ~x280;
assign c8119 =  x653 & ~x335 & ~x340 & ~x368 & ~x454 & ~x508 & ~x563;
assign c8121 = ~x109 & ~x137 & ~x395 & ~x472 & ~x480 & ~x551 & ~x583 & ~x592 & ~x620 & ~x675 & ~x703 & ~x725;
assign c8123 = ~x19 & ~x152 & ~x180 & ~x199 & ~x286 & ~x312 & ~x340 & ~x342 & ~x368 & ~x395 & ~x716 & ~x747 & ~x755 & ~x761;
assign c8125 =  x463 &  x497 &  x750 & ~x23 & ~x308 & ~x334 & ~x416 & ~x478 & ~x559 & ~x590 & ~x613 & ~x753;
assign c8127 =  x103 & ~x41 & ~x474 & ~x480 & ~x501 & ~x505 & ~x508 & ~x584 & ~x613 & ~x618 & ~x701;
assign c8129 =  x296 &  x453 & ~x647 & ~x667 & ~x695;
assign c8131 = ~x366 & ~x393 & ~x411 & ~x474 & ~x564 & ~x583 & ~x585;
assign c8133 =  x410 &  x445 &  x473 &  x491 &  x543 & ~x261 & ~x316;
assign c8135 =  x73 &  x99 &  x100 &  x465 &  x487 &  x655 & ~x32 & ~x53 & ~x82 & ~x109 & ~x138 & ~x141 & ~x142 & ~x194 & ~x197 & ~x225 & ~x279 & ~x336 & ~x449 & ~x474 & ~x559 & ~x643 & ~x672 & ~x760;
assign c8137 = ~x227 & ~x234 & ~x340 & ~x374 & ~x402;
assign c8139 =  x135 & ~x252 & ~x454;
assign c8141 =  x625 & ~x3 & ~x41 & ~x114 & ~x199 & ~x339 & ~x340 & ~x360 & ~x368 & ~x480 & ~x535 & ~x647 & ~x675;
assign c8143 =  x206 &  x408 &  x718 & ~x534 & ~x589 & ~x620 & ~x621;
assign c8145 =  x463 & ~x58 & ~x340 & ~x500 & ~x613 & ~x636 & ~x675;
assign c8147 =  x530 & ~x236 & ~x262 & ~x312 & ~x634 & ~x649 & ~x659;
assign c8149 = ~x366 & ~x416 & ~x546 & ~x547 & ~x591 & ~x675 & ~x696;
assign c8151 =  x192 & ~x425;
assign c8153 =  x75 &  x212 &  x286 &  x597 &  x747 & ~x81 & ~x195 & ~x196 & ~x280 & ~x532;
assign c8155 =  x453 & ~x179 & ~x283 & ~x636 & ~x670;
assign c8157 =  x332 & ~x15 & ~x66 & ~x201 & ~x262;
assign c8159 =  x43 &  x44 &  x68 &  x69 &  x70 &  x71 & ~x532 & ~x588;
assign c8161 =  x408 &  x486 &  x516 &  x540 &  x598 &  x601 & ~x16 & ~x45 & ~x87 & ~x195 & ~x367 & ~x675 & ~x703;
assign c8163 = ~x15 & ~x284 & ~x319 & ~x451 & ~x616 & ~x744;
assign c8165 =  x410 &  x416 &  x423 &  x429 & ~x84 & ~x169 & ~x194 & ~x593 & ~x649;
assign c8167 =  x68 &  x397 &  x508 & ~x56 & ~x109 & ~x366 & ~x390 & ~x559 & ~x783;
assign c8169 =  x529 & ~x13 & ~x179 & ~x288 & ~x314 & ~x337 & ~x661 & ~x689;
assign c8171 = ~x319 & ~x402 & ~x559;
assign c8173 = ~x14 & ~x208 & ~x227 & ~x292 & ~x340 & ~x365 & ~x395 & ~x744;
assign c8175 = ~x254 & ~x257 & ~x552 & ~x585 & ~x636 & ~x675 & ~x770;
assign c8177 =  x43 &  x69 &  x71 &  x593 & ~x34;
assign c8179 =  x204 &  x232 &  x341 &  x359 &  x388 &  x423 & ~x80 & ~x137 & ~x559;
assign c8181 = ~x411 & ~x474 & ~x492;
assign c8183 =  x779;
assign c8185 =  x209 &  x650 &  x695 & ~x22 & ~x30 & ~x109 & ~x143 & ~x340 & ~x360 & ~x366 & ~x395 & ~x421 & ~x502 & ~x529 & ~x588 & ~x647;
assign c8187 =  x375 &  x739 & ~x199 & ~x279 & ~x283 & ~x368 & ~x472 & ~x480 & ~x585 & ~x639 & ~x647 & ~x777;
assign c8189 = ~x174 & ~x234 & ~x285 & ~x337 & ~x340 & ~x368 & ~x423 & ~x743 & ~x748;
assign c8191 =  x41 &  x42 &  x43 &  x44 & ~x3 & ~x8 & ~x19 & ~x27 & ~x34 & ~x50 & ~x55 & ~x60 & ~x80 & ~x81 & ~x113 & ~x137 & ~x141 & ~x165 & ~x168 & ~x171 & ~x193 & ~x199 & ~x226 & ~x252 & ~x254 & ~x280 & ~x282 & ~x307 & ~x310 & ~x335 & ~x336 & ~x361 & ~x362 & ~x366 & ~x391 & ~x420 & ~x446 & ~x478 & ~x561 & ~x589 & ~x617 & ~x698 & ~x729;
assign c8193 =  x440 & ~x279 & ~x286 & ~x312 & ~x340 & ~x636;
assign c8195 =  x15 &  x41 &  x42 &  x43 & ~x5 & ~x9 & ~x34 & ~x59 & ~x113 & ~x115 & ~x143 & ~x168 & ~x195 & ~x225 & ~x254 & ~x334 & ~x337 & ~x338 & ~x360 & ~x363 & ~x393 & ~x420 & ~x421 & ~x446 & ~x447 & ~x448 & ~x450 & ~x559 & ~x561 & ~x588 & ~x616 & ~x617 & ~x642 & ~x702 & ~x781;
assign c8197 =  x463 & ~x2 & ~x22 & ~x33 & ~x34 & ~x109 & ~x141 & ~x280 & ~x532 & ~x535 & ~x536 & ~x557 & ~x560 & ~x562 & ~x583 & ~x584 & ~x592 & ~x610 & ~x617 & ~x620 & ~x621 & ~x639 & ~x644 & ~x669 & ~x676 & ~x698 & ~x703 & ~x704 & ~x727 & ~x751 & ~x780 & ~x781;
assign c8199 =  x275 &  x303 &  x331 &  x359 &  x360 &  x472 &  x585 &  x641 & ~x23 & ~x26 & ~x137 & ~x251;
assign c8201 =  x408 &  x463 &  x465 & ~x2 & ~x13 & ~x44 & ~x53 & ~x480 & ~x505 & ~x509 & ~x556 & ~x620 & ~x727;
assign c8203 =  x536 &  x566 & ~x168 & ~x337 & ~x340 & ~x766;
assign c8205 =  x535 &  x536 & ~x227 & ~x311 & ~x366;
assign c8207 =  x132 &  x184 &  x564 & ~x280 & ~x389 & ~x474;
assign c8209 = ~x8 & ~x137 & ~x138 & ~x208 & ~x213 & ~x234 & ~x277 & ~x534 & ~x536 & ~x605;
assign c8211 =  x410 & ~x14 & ~x26 & ~x208 & ~x227 & ~x234 & ~x262 & ~x286 & ~x310 & ~x312 & ~x661 & ~x746 & ~x748 & ~x765 & ~x766;
assign c8213 =  x65 &  x103 &  x154 &  x204 &  x360 &  x368 & ~x25;
assign c8215 =  x44 &  x69 &  x71 & ~x2 & ~x90 & ~x559;
assign c8217 =  x342 &  x485 &  x733 & ~x169 & ~x253 & ~x255 & ~x311 & ~x393 & ~x417 & ~x671;
assign c8219 =  x573 & ~x23 & ~x151 & ~x176 & ~x206 & ~x227 & ~x229 & ~x231 & ~x255 & ~x282 & ~x286 & ~x310 & ~x340 & ~x366 & ~x368 & ~x395 & ~x643 & ~x689 & ~x701 & ~x741 & ~x748 & ~x775;
assign c8221 = ~x13 & ~x14 & ~x41 & ~x59 & ~x116 & ~x206 & ~x227 & ~x262 & ~x263 & ~x280 & ~x311 & ~x319 & ~x422 & ~x761;
assign c8223 =  x175 &  x243 &  x272 &  x314 &  x358 &  x386 &  x414 & ~x22 & ~x53 & ~x113 & ~x171 & ~x196 & ~x251 & ~x276 & ~x361 & ~x366 & ~x390 & ~x417 & ~x448 & ~x504 & ~x531 & ~x587;
assign c8225 = ~x0 & ~x27 & ~x196 & ~x411 & ~x417 & ~x451 & ~x478 & ~x502 & ~x527 & ~x560 & ~x563 & ~x613 & ~x618 & ~x781;
assign c8227 =  x750 & ~x32 & ~x54 & ~x80 & ~x114 & ~x225 & ~x227 & ~x249 & ~x252 & ~x282 & ~x390 & ~x391 & ~x417 & ~x421 & ~x446 & ~x476 & ~x561 & ~x757 & ~x774;
assign c8229 =  x510 & ~x141 & ~x251 & ~x340 & ~x365 & ~x366 & ~x633 & ~x661 & ~x715 & ~x718 & ~x722 & ~x767;
assign c8231 = ~x184 & ~x236 & ~x532 & ~x546 & ~x578 & ~x602 & ~x621;
assign c8233 =  x41 &  x43 &  x70 & ~x80 & ~x113 & ~x116 & ~x199 & ~x336 & ~x337 & ~x530 & ~x562 & ~x590 & ~x701;
assign c8235 =  x473 & ~x30 & ~x174 & ~x196 & ~x285 & ~x286 & ~x312;
assign c8237 =  x43 &  x70 & ~x50 & ~x337 & ~x505 & ~x703;
assign c8239 =  x750 & ~x5 & ~x57 & ~x170 & ~x195 & ~x227 & ~x252 & ~x282 & ~x283 & ~x338 & ~x363 & ~x389 & ~x420 & ~x590 & ~x645 & ~x765 & ~x781;
assign c8241 =  x47 & ~x6 & ~x25 & ~x56 & ~x113 & ~x114 & ~x390 & ~x393 & ~x449 & ~x450 & ~x473 & ~x507 & ~x529 & ~x588 & ~x701;
assign c8243 =  x119 &  x148 &  x541 &  x656 &  x746 &  x769 &  x770 & ~x616;
assign c8245 =  x444 & ~x14 & ~x227 & ~x233 & ~x262 & ~x636;
assign c8247 =  x185 &  x626 & ~x13 & ~x41 & ~x339 & ~x340 & ~x342 & ~x368 & ~x397 & ~x421;
assign c8249 =  x45 & ~x391 & ~x528 & ~x536 & ~x562 & ~x591 & ~x644 & ~x647 & ~x667 & ~x668 & ~x675 & ~x698 & ~x703;
assign c8251 = ~x227 & ~x258 & ~x280 & ~x339 & ~x340 & ~x342 & ~x366 & ~x368 & ~x395 & ~x688 & ~x744 & ~x766 & ~x767;
assign c8253 =  x42 &  x43 &  x329 &  x508 & ~x199;
assign c8255 =  x613 & ~x398;
assign c8257 =  x173 & ~x450 & ~x480 & ~x529 & ~x642;
assign c8259 = ~x225 & ~x292 & ~x544 & ~x689;
assign c8261 =  x121 &  x185 &  x187 &  x205 &  x232 &  x259 &  x266 &  x270 &  x292 &  x331 &  x368 &  x396 &  x444 &  x461 &  x486 &  x662 & ~x53 & ~x112 & ~x334 & ~x336;
assign c8263 =  x243 & ~x28 & ~x50 & ~x110 & ~x113 & ~x138 & ~x169 & ~x227 & ~x292 & ~x340 & ~x368 & ~x450 & ~x451 & ~x478 & ~x480 & ~x534;
assign c8265 =  x121 &  x175 &  x231 &  x426 & ~x80 & ~x227 & ~x283 & ~x308 & ~x418 & ~x449 & ~x589 & ~x765;
assign c8267 =  x64 &  x92 &  x204 &  x598 &  x680 & ~x23 & ~x28 & ~x647 & ~x667 & ~x675 & ~x729;
assign c8269 = ~x14 & ~x113 & ~x199 & ~x249 & ~x278 & ~x283 & ~x387 & ~x451 & ~x454 & ~x508 & ~x528 & ~x554 & ~x583 & ~x592 & ~x621 & ~x638 & ~x649 & ~x675 & ~x703;
assign c8271 =  x507 & ~x228 & ~x255 & ~x256 & ~x366 & ~x711;
assign c8273 =  x41 &  x43 &  x69 &  x70 &  x538 &  x654 & ~x54 & ~x109 & ~x168 & ~x198 & ~x222 & ~x225 & ~x227 & ~x278 & ~x279 & ~x281 & ~x307 & ~x363 & ~x418 & ~x474;
assign c8275 =  x243 &  x598 &  x625 & ~x27 & ~x340 & ~x368 & ~x748;
assign c8277 =  x40 &  x41 &  x69 & ~x49 & ~x473 & ~x475;
assign c8279 =  x296 &  x462 & ~x13 & ~x41 & ~x224 & ~x533 & ~x639 & ~x640;
assign c8281 = ~x8 & ~x13 & ~x26 & ~x148 & ~x152 & ~x200 & ~x206 & ~x227 & ~x236 & ~x256 & ~x283 & ~x286 & ~x311 & ~x337 & ~x339 & ~x340 & ~x616 & ~x690 & ~x742 & ~x744 & ~x770 & ~x783;
assign c8283 =  x65 &  x189 &  x621 & ~x80 & ~x109 & ~x113 & ~x140 & ~x420 & ~x450 & ~x531;
assign c8285 = ~x2 & ~x128 & ~x139 & ~x158 & ~x172 & ~x192 & ~x285 & ~x309 & ~x338 & ~x339 & ~x605 & ~x635 & ~x669 & ~x726 & ~x749 & ~x770;
assign c8287 =  x42 &  x43 &  x44 & ~x109 & ~x473 & ~x591 & ~x675 & ~x696 & ~x703;
assign c8289 = ~x295 & ~x319 & ~x474 & ~x600;
assign c8291 =  x78 &  x134 & ~x2 & ~x14 & ~x15 & ~x480;
assign c8293 =  x296 &  x352 &  x571 &  x598 & ~x194 & ~x196 & ~x284 & ~x304 & ~x308 & ~x448 & ~x472 & ~x479 & ~x501 & ~x531 & ~x647 & ~x675 & ~x703 & ~x780;
assign c8295 =  x18 & ~x3 & ~x57 & ~x112 & ~x195 & ~x308 & ~x363 & ~x365 & ~x366 & ~x420 & ~x421 & ~x473 & ~x505;
assign c8297 =  x39 & ~x0 & ~x54 & ~x225 & ~x283 & ~x360 & ~x366 & ~x423 & ~x472 & ~x473 & ~x502 & ~x507 & ~x676 & ~x701 & ~x703;
assign c8299 =  x424 & ~x60 & ~x250 & ~x335 & ~x560 & ~x602 & ~x636;
assign c8301 =  x71 &  x414 &  x751;
assign c8303 =  x410 & ~x14 & ~x96 & ~x199 & ~x286 & ~x340 & ~x342 & ~x425;
assign c8305 =  x41 &  x42 &  x43 & ~x52 & ~x82 & ~x165 & ~x193 & ~x340 & ~x361 & ~x390 & ~x417 & ~x446 & ~x558 & ~x589 & ~x701;
assign c8307 =  x553 &  x750 & ~x224 & ~x393 & ~x501 & ~x591 & ~x619 & ~x647 & ~x675 & ~x701;
assign c8309 =  x444 &  x585 & ~x226 & ~x260 & ~x421 & ~x531;
assign c8311 =  x154 &  x444 &  x585 &  x613 &  x614;
assign c8313 =  x453 & ~x130 & ~x149 & ~x180 & ~x207 & ~x253 & ~x255 & ~x309 & ~x630 & ~x632;
assign c8315 =  x471 & ~x1 & ~x15 & ~x54 & ~x59 & ~x72 & ~x122 & ~x234 & ~x255 & ~x260 & ~x261 & ~x262 & ~x282 & ~x290 & ~x340;
assign c8317 =  x518 &  x570 & ~x6 & ~x13 & ~x14 & ~x24 & ~x61 & ~x69 & ~x90 & ~x142 & ~x173 & ~x196 & ~x199 & ~x223 & ~x227 & ~x230 & ~x364 & ~x368 & ~x393 & ~x399 & ~x450;
assign c8319 =  x453 & ~x5 & ~x13 & ~x15 & ~x23 & ~x49 & ~x61 & ~x222 & ~x280 & ~x337 & ~x338 & ~x339 & ~x340 & ~x616 & ~x618 & ~x647 & ~x703 & ~x781;
assign c8321 = ~x319 & ~x340 & ~x433 & ~x480;
assign c8323 = ~x82 & ~x141 & ~x279 & ~x337 & ~x354 & ~x361 & ~x504 & ~x505 & ~x590 & ~x703 & ~x773;
assign c8325 =  x221;
assign c8327 =  x93 &  x133 &  x147 &  x189 &  x202 &  x230 &  x598 & ~x335 & ~x393 & ~x450;
assign c8329 =  x482 & ~x261 & ~x661 & ~x767;
assign c8331 = ~x14 & ~x125 & ~x184 & ~x390 & ~x554 & ~x556 & ~x621 & ~x639 & ~x648 & ~x777;
assign c8333 =  x346 &  x394 &  x396 &  x423 & ~x533;
assign c8335 =  x144 &  x145 & ~x109 & ~x166 & ~x449 & ~x474 & ~x559;
assign c8337 =  x147 &  x554 &  x564 &  x723 & ~x165 & ~x277 & ~x393 & ~x421 & ~x446 & ~x783;
assign c8339 = ~x33 & ~x137 & ~x147 & ~x207 & ~x228 & ~x234 & ~x254 & ~x257 & ~x282 & ~x284 & ~x285 & ~x310 & ~x311 & ~x337 & ~x504 & ~x607 & ~x633 & ~x635 & ~x661 & ~x689 & ~x747 & ~x762;
assign c8341 =  x175 &  x508 &  x509 &  x513 &  x723 & ~x165 & ~x169 & ~x279 & ~x362;
assign c8343 =  x295 &  x296 &  x598 & ~x15 & ~x41 & ~x227 & ~x279 & ~x339 & ~x340 & ~x368;
assign c8345 =  x305 & ~x7 & ~x13 & ~x231 & ~x255 & ~x287 & ~x307 & ~x310 & ~x338 & ~x587 & ~x741 & ~x762 & ~x763 & ~x766;
assign c8347 = ~x543 & ~x573 & ~x584;
assign c8349 =  x585 &  x590 &  x612 &  x641 & ~x279;
assign c8351 = ~x382 & ~x474 & ~x766;
assign c8353 =  x99 &  x584 &  x696 & ~x23 & ~x279 & ~x475;
assign c8355 = ~x171 & ~x179 & ~x180 & ~x181 & ~x200 & ~x206 & ~x222 & ~x229 & ~x232 & ~x233 & ~x253 & ~x254 & ~x258 & ~x261 & ~x262 & ~x284 & ~x315 & ~x340 & ~x366 & ~x661 & ~x663 & ~x675 & ~x687 & ~x688 & ~x716 & ~x743 & ~x744 & ~x745;
assign c8357 =  x68 &  x126 &  x465 &  x654 & ~x0 & ~x32 & ~x80 & ~x84 & ~x109 & ~x112 & ~x113 & ~x139 & ~x227 & ~x361 & ~x613 & ~x617;
assign c8359 =  x187 &  x621 & ~x80 & ~x90 & ~x417 & ~x473 & ~x474 & ~x559;
assign c8361 = ~x326 & ~x338 & ~x366 & ~x516 & ~x536;
assign c8363 =  x739 & ~x385 & ~x397 & ~x425 & ~x473 & ~x480 & ~x502 & ~x558 & ~x583 & ~x610 & ~x620 & ~x621 & ~x639 & ~x649 & ~x675 & ~x703;
assign c8365 = ~x138 & ~x141 & ~x198 & ~x225 & ~x366 & ~x368 & ~x385 & ~x387 & ~x396 & ~x454 & ~x472 & ~x483 & ~x497 & ~x505 & ~x533 & ~x675;
assign c8367 =  x42 &  x43 &  x44 &  x99 & ~x19 & ~x80 & ~x109 & ~x137 & ~x699;
assign c8369 = ~x15 & ~x26 & ~x41 & ~x60 & ~x113 & ~x227 & ~x255 & ~x286 & ~x311 & ~x338 & ~x339 & ~x340 & ~x368 & ~x397 & ~x425 & ~x450 & ~x451 & ~x453 & ~x454 & ~x480 & ~x505 & ~x532 & ~x534;
assign c8371 =  x192 & ~x480;
assign c8373 =  x135 & ~x425 & ~x480;
assign c8375 =  x101 &  x128 &  x129 &  x150 &  x284 &  x313 &  x320 &  x331 &  x376 &  x434 &  x486 &  x606 &  x661 & ~x6 & ~x137 & ~x168 & ~x279 & ~x672 & ~x728;
assign c8377 =  x158 &  x184 &  x214 &  x444 &  x584 &  x591 &  x619 &  x641 & ~x57 & ~x251 & ~x335 & ~x447;
assign c8379 =  x422 &  x449 & ~x610;
assign c8381 =  x105 &  x144 &  x256 &  x275 &  x283 & ~x196;
assign c8383 =  x383 &  x442 & ~x143 & ~x177 & ~x204 & ~x234 & ~x255 & ~x260 & ~x283 & ~x286 & ~x311 & ~x340 & ~x661 & ~x662 & ~x688 & ~x727 & ~x745;
assign c8385 =  x15 &  x41 &  x42 &  x43 & ~x83;
assign c8387 =  x201 & ~x24 & ~x27 & ~x508 & ~x527 & ~x528 & ~x532 & ~x558 & ~x562 & ~x563 & ~x588 & ~x589 & ~x591 & ~x593 & ~x616 & ~x668 & ~x675 & ~x702;
assign c8389 =  x481 & ~x186 & ~x285 & ~x311 & ~x648 & ~x675;
assign c8391 =  x70 &  x71 &  x397 &  x487 &  x564 & ~x6 & ~x23 & ~x137 & ~x141 & ~x168 & ~x196 & ~x225 & ~x393 & ~x560;
assign c8393 =  x175 &  x538 & ~x90 & ~x109 & ~x220 & ~x226 & ~x284 & ~x361 & ~x449 & ~x451 & ~x479 & ~x501 & ~x505 & ~x533 & ~x617 & ~x646 & ~x675;
assign c8395 =  x410 &  x453 & ~x575;
assign c8397 =  x98 &  x102 &  x134 &  x228 &  x568 & ~x139 & ~x504;
assign c8399 =  x64 &  x134 &  x145 &  x148 &  x256 &  x488 & ~x80 & ~x195 & ~x476 & ~x700;
assign c8401 =  x40 &  x41 &  x42 & ~x2 & ~x5 & ~x8 & ~x49 & ~x56 & ~x59 & ~x60 & ~x83 & ~x113 & ~x141 & ~x168 & ~x198 & ~x221 & ~x222 & ~x253 & ~x277 & ~x279 & ~x280 & ~x308 & ~x361 & ~x363 & ~x418 & ~x420 & ~x446 & ~x447 & ~x448 & ~x450 & ~x474 & ~x475 & ~x478 & ~x505 & ~x530 & ~x533 & ~x559 & ~x562 & ~x588 & ~x590 & ~x614 & ~x616 & ~x642 & ~x729 & ~x781;
assign c8403 =  x410 & ~x14 & ~x39 & ~x72 & ~x113 & ~x172 & ~x199 & ~x227 & ~x261 & ~x338 & ~x340 & ~x661;
assign c8405 = ~x23 & ~x168 & ~x311 & ~x338 & ~x339 & ~x366 & ~x393 & ~x395 & ~x396 & ~x411 & ~x473 & ~x474 & ~x500 & ~x559 & ~x562 & ~x588 & ~x669 & ~x725;
assign c8407 = ~x141 & ~x225 & ~x234 & ~x381 & ~x488;
assign c8409 =  x443 &  x444 & ~x84 & ~x252 & ~x262 & ~x264 & ~x311;
assign c8411 = ~x199 & ~x200 & ~x227 & ~x254 & ~x283 & ~x310 & ~x474 & ~x483 & ~x534 & ~x765;
assign c8413 =  x203 &  x750 & ~x584 & ~x675 & ~x703;
assign c8415 =  x331 & ~x290 & ~x721 & ~x765;
assign c8417 =  x178 &  x210 &  x238 &  x314 &  x324 &  x349 &  x375 &  x406 &  x518 &  x546 &  x604 & ~x2 & ~x30 & ~x88 & ~x138 & ~x141 & ~x198 & ~x227 & ~x249 & ~x309 & ~x418 & ~x698;
assign c8419 =  x266 &  x268 &  x324 &  x463 &  x606 &  x629 &  x653 & ~x146 & ~x199 & ~x227 & ~x360;
assign c8421 =  x266 &  x296 &  x352 &  x376 &  x381 &  x404 &  x486 &  x491 &  x492 &  x629 & ~x3 & ~x16 & ~x24 & ~x142 & ~x165 & ~x169 & ~x196 & ~x197 & ~x505 & ~x508 & ~x534 & ~x559 & ~x562 & ~x583 & ~x588 & ~x616 & ~x619 & ~x620 & ~x647 & ~x648 & ~x698 & ~x757;
assign c8423 =  x751 & ~x2;
assign c8425 =  x656 & ~x53 & ~x113 & ~x338 & ~x473 & ~x474 & ~x478 & ~x497 & ~x505 & ~x643 & ~x675 & ~x705;
assign c8427 =  x332 & ~x54 & ~x368 & ~x395;
assign c8429 = ~x234 & ~x284 & ~x340 & ~x583;
assign c8431 =  x68 &  x98 & ~x49 & ~x220 & ~x283 & ~x473 & ~x505;
assign c8433 =  x68 &  x69 &  x70 &  x554 &  x593 & ~x113 & ~x366;
assign c8435 =  x40 &  x68 &  x97 &  x127 &  x515 &  x607 &  x653 & ~x34 & ~x250;
assign c8437 =  x151 &  x209 &  x210 &  x243 &  x314 &  x537 &  x625 & ~x49 & ~x281;
assign c8439 = ~x186 & ~x227 & ~x263 & ~x561 & ~x603 & ~x636 & ~x688;
assign c8441 =  x43 &  x70 & ~x90 & ~x502;
assign c8443 = ~x198 & ~x199 & ~x234 & ~x286 & ~x340 & ~x402 & ~x429 & ~x480;
assign c8445 = ~x113 & ~x227 & ~x261 & ~x340 & ~x366 & ~x368 & ~x393 & ~x402;
assign c8447 = ~x156 & ~x186 & ~x263 & ~x282 & ~x284 & ~x312 & ~x338 & ~x339 & ~x602 & ~x620 & ~x658;
assign c8449 =  x68 &  x96 &  x97 &  x508 &  x564;
assign c8451 =  x750 & ~x6 & ~x26 & ~x50 & ~x78 & ~x109 & ~x113 & ~x164 & ~x251 & ~x334 & ~x472 & ~x473 & ~x533 & ~x590 & ~x613 & ~x669;
assign c8453 =  x585 & ~x338 & ~x422;
assign c8455 = ~x141 & ~x199 & ~x284 & ~x319 & ~x366 & ~x718 & ~x744 & ~x748;
assign c8457 = ~x23 & ~x80 & ~x109 & ~x165 & ~x340 & ~x368 & ~x390 & ~x415 & ~x523 & ~x584 & ~x585 & ~x696 & ~x703 & ~x704;
assign c8459 =  x214 &  x235 &  x240 &  x241 &  x262 &  x293 &  x381 &  x405 &  x457 &  x492 &  x540 &  x542 &  x652 & ~x13 & ~x620 & ~x703 & ~x730;
assign c8461 =  x210 &  x598 & ~x3 & ~x166 & ~x449 & ~x610;
assign c8463 =  x410 &  x470 &  x473 & ~x308 & ~x340 & ~x703;
assign c8465 =  x381 &  x403 &  x486 &  x487 &  x514 &  x576 &  x626 &  x629 &  x631 & ~x13 & ~x14 & ~x15 & ~x44 & ~x81 & ~x196 & ~x503 & ~x505 & ~x507 & ~x508 & ~x534 & ~x559 & ~x639 & ~x647 & ~x675 & ~x701 & ~x703;
assign c8467 =  x360 &  x585 &  x618 &  x641 & ~x141 & ~x448;
assign c8469 =  x158 &  x754;
assign c8471 =  x13 &  x41 & ~x2 & ~x7 & ~x8 & ~x53 & ~x59 & ~x60 & ~x109 & ~x114 & ~x137 & ~x141 & ~x143 & ~x166 & ~x168 & ~x222 & ~x226 & ~x279 & ~x280 & ~x282 & ~x337 & ~x389 & ~x393 & ~x450 & ~x478 & ~x505 & ~x533 & ~x560 & ~x729 & ~x757;
assign c8473 =  x64 &  x145 &  x286 &  x479 &  x529 & ~x23 & ~x54;
assign c8475 = ~x59 & ~x186 & ~x208 & ~x227 & ~x252 & ~x253 & ~x280 & ~x309 & ~x578 & ~x661;
assign c8477 =  x296 & ~x7 & ~x171 & ~x234 & ~x251 & ~x282 & ~x288 & ~x340;
assign c8479 =  x458 &  x486 & ~x33 & ~x137 & ~x141 & ~x168 & ~x195 & ~x227 & ~x252 & ~x254 & ~x280 & ~x309 & ~x311 & ~x359 & ~x360 & ~x366 & ~x367 & ~x388 & ~x390 & ~x393 & ~x395 & ~x415 & ~x423 & ~x448 & ~x478 & ~x507 & ~x586 & ~x644 & ~x669 & ~x675 & ~x781;
assign c8481 = ~x207 & ~x292 & ~x340 & ~x366 & ~x689;
assign c8483 =  x15 &  x42 &  x43 & ~x279 & ~x473;
assign c8485 = ~x23 & ~x234 & ~x280 & ~x325 & ~x366 & ~x465;
assign c8487 =  x69 &  x70 & ~x19 & ~x49 & ~x169 & ~x447 & ~x451 & ~x590 & ~x646;
assign c8489 =  x653 & ~x399 & ~x616 & ~x675;
assign c8491 = ~x179 & ~x199 & ~x234 & ~x285 & ~x290 & ~x311 & ~x340 & ~x688 & ~x689;
assign c8493 = ~x14 & ~x227 & ~x236 & ~x261 & ~x263 & ~x290 & ~x337 & ~x338 & ~x744 & ~x761 & ~x770;
assign c8495 =  x100 &  x127 &  x130 &  x184 &  x210 &  x296 &  x330 &  x564 &  x565 &  x652 & ~x111 & ~x280 & ~x338 & ~x393;
assign c8497 = ~x2 & ~x311 & ~x402 & ~x451 & ~x748 & ~x767;
assign c8499 =  x100 &  x130 &  x507 &  x508 &  x557 &  x585 &  x598 &  x613;
assign c90 =  x327 &  x387 &  x415 &  x470 &  x493 &  x501 &  x521 &  x530 &  x554 &  x555 &  x574 & ~x0 & ~x43 & ~x57 & ~x58 & ~x103 & ~x104 & ~x207 & ~x228 & ~x236 & ~x373 & ~x397 & ~x420 & ~x427 & ~x429 & ~x662 & ~x713 & ~x732 & ~x742 & ~x746 & ~x754 & ~x765;
assign c92 =  x496 &  x534 &  x535 &  x584 & ~x35 & ~x96 & ~x100 & ~x112 & ~x168 & ~x202 & ~x233 & ~x256 & ~x661;
assign c94 =  x274 &  x294 &  x358 & ~x252 & ~x594;
assign c96 =  x293 &  x303 &  x376 &  x543 &  x547 & ~x143 & ~x198 & ~x202 & ~x226 & ~x763 & ~x772;
assign c98 = ~x25 & ~x58 & ~x108 & ~x174 & ~x179 & ~x195 & ~x227 & ~x281 & ~x335 & ~x397 & ~x419 & ~x422 & ~x429 & ~x451 & ~x455 & ~x457 & ~x476 & ~x480 & ~x482 & ~x483 & ~x485 & ~x510 & ~x511 & ~x512;
assign c910 =  x387 &  x573 &  x583 &  x611 & ~x29 & ~x78 & ~x135 & ~x682 & ~x702 & ~x743 & ~x752 & ~x757;
assign c912 =  x212 &  x246 &  x247 &  x248 &  x273 &  x296 &  x304 &  x382 &  x517 &  x543 &  x624 &  x626 & ~x27 & ~x92 & ~x120 & ~x142 & ~x168 & ~x198 & ~x309 & ~x311 & ~x315 & ~x367 & ~x729;
assign c914 =  x619 &  x651 &  x656 & ~x400 & ~x455;
assign c916 =  x212 &  x354 &  x452 & ~x229 & ~x233 & ~x770;
assign c918 =  x467 &  x499 &  x520 &  x562 &  x598 & ~x29 & ~x107 & ~x113 & ~x123 & ~x161 & ~x174 & ~x206 & ~x230 & ~x254 & ~x345 & ~x425 & ~x504 & ~x698 & ~x705 & ~x750 & ~x755;
assign c920 =  x638 & ~x455 & ~x479 & ~x513;
assign c922 =  x321 &  x459 &  x488 & ~x10 & ~x157 & ~x206 & ~x567 & ~x605 & ~x680;
assign c924 =  x576 & ~x57 & ~x93 & ~x187 & ~x259 & ~x400 & ~x401 & ~x588 & ~x743;
assign c926 =  x467 &  x495 &  x584 & ~x8 & ~x22 & ~x42 & ~x56 & ~x58 & ~x59 & ~x134 & ~x152 & ~x157 & ~x162 & ~x171 & ~x206 & ~x401 & ~x633 & ~x703 & ~x765;
assign c928 =  x273 &  x326 &  x354 &  x406 &  x459 &  x462 &  x463 &  x488 &  x521 &  x541 &  x542 &  x546 & ~x13 & ~x18 & ~x30 & ~x42 & ~x72 & ~x76 & ~x77 & ~x81 & ~x103 & ~x104 & ~x108 & ~x111 & ~x120 & ~x121 & ~x122 & ~x126 & ~x129 & ~x131 & ~x133 & ~x134 & ~x143 & ~x151 & ~x158 & ~x168 & ~x173 & ~x174 & ~x178 & ~x180 & ~x197 & ~x198 & ~x199 & ~x206 & ~x223 & ~x231 & ~x262 & ~x287 & ~x290 & ~x291 & ~x308 & ~x335 & ~x345 & ~x366 & ~x427 & ~x476 & ~x504 & ~x675 & ~x689 & ~x698 & ~x706 & ~x713 & ~x718 & ~x726 & ~x734 & ~x735 & ~x736 & ~x737 & ~x738 & ~x739 & ~x752 & ~x761 & ~x765 & ~x769 & ~x783;
assign c930 =  x249 &  x452 & ~x226 & ~x596 & ~x680 & ~x769;
assign c932 = ~x68 & ~x84 & ~x144 & ~x157 & ~x480 & ~x481 & ~x511 & ~x707;
assign c934 =  x158 &  x187 &  x188 &  x410 &  x462 & ~x59 & ~x87 & ~x90 & ~x121 & ~x197 & ~x198 & ~x253 & ~x254 & ~x366 & ~x419 & ~x775;
assign c936 =  x522 &  x648 &  x683 & ~x36;
assign c938 = ~x24 & ~x39 & ~x131 & ~x206 & ~x419 & ~x429 & ~x455 & ~x483 & ~x484 & ~x765;
assign c940 =  x350 &  x387 &  x389 &  x478 &  x534 & ~x59 & ~x87 & ~x95 & ~x136 & ~x229 & ~x419 & ~x605 & ~x645 & ~x703 & ~x765;
assign c942 =  x293 &  x294 &  x320 &  x348 &  x446 & ~x126 & ~x149 & ~x185 & ~x723 & ~x763;
assign c944 =  x212 &  x267 &  x328 &  x331 &  x349 &  x383 &  x415 &  x493 &  x499 &  x502 &  x507 &  x526 &  x546 & ~x93 & ~x112 & ~x227 & ~x231 & ~x338 & ~x674 & ~x680 & ~x716 & ~x720 & ~x735 & ~x776;
assign c946 = ~x29 & ~x33 & ~x59 & ~x62 & ~x64 & ~x84 & ~x92 & ~x94 & ~x118 & ~x121 & ~x136 & ~x143 & ~x146 & ~x172 & ~x196 & ~x204 & ~x223 & ~x233 & ~x281 & ~x392 & ~x396 & ~x429 & ~x454 & ~x455 & ~x457 & ~x475 & ~x479 & ~x482 & ~x483 & ~x541 & ~x689;
assign c948 =  x348 &  x409 &  x410 &  x506 &  x541 &  x613 & ~x18 & ~x56 & ~x58 & ~x84 & ~x94 & ~x120 & ~x177 & ~x226 & ~x229 & ~x254 & ~x727 & ~x758 & ~x777;
assign c950 =  x506 &  x542 &  x543 &  x558 & ~x21 & ~x152 & ~x223 & ~x374 & ~x400 & ~x628 & ~x686;
assign c952 =  x609 & ~x9 & ~x12 & ~x31 & ~x35 & ~x44 & ~x59 & ~x66 & ~x67 & ~x92 & ~x95 & ~x112 & ~x122 & ~x140 & ~x149 & ~x169 & ~x179 & ~x201 & ~x204 & ~x205 & ~x226 & ~x229 & ~x252 & ~x281 & ~x289 & ~x337 & ~x362 & ~x396 & ~x400 & ~x401 & ~x453 & ~x532 & ~x728 & ~x744 & ~x758 & ~x761;
assign c954 =  x300 &  x303 &  x388 &  x486 & ~x43 & ~x113 & ~x136 & ~x137 & ~x214 & ~x291 & ~x577 & ~x596 & ~x613;
assign c956 = ~x60 & ~x80 & ~x112 & ~x170 & ~x281 & ~x315 & ~x397 & ~x401 & ~x429 & ~x448 & ~x455 & ~x482 & ~x483 & ~x485 & ~x509 & ~x511 & ~x513 & ~x538 & ~x567;
assign c958 =  x296 &  x359 &  x380 &  x383 &  x545 &  x572 &  x655 & ~x65 & ~x144 & ~x149 & ~x168 & ~x205 & ~x314 & ~x315 & ~x342;
assign c960 = ~x27 & ~x40 & ~x42 & ~x43 & ~x66 & ~x89 & ~x122 & ~x135 & ~x137 & ~x140 & ~x141 & ~x146 & ~x150 & ~x174 & ~x180 & ~x199 & ~x204 & ~x205 & ~x228 & ~x252 & ~x282 & ~x334 & ~x362 & ~x368 & ~x372 & ~x390 & ~x395 & ~x400 & ~x427 & ~x446 & ~x451 & ~x730 & ~x757 & ~x758 & ~x765 & ~x770 & ~x771 & ~x775;
assign c962 =  x296 &  x474 &  x507 & ~x35 & ~x79 & ~x84 & ~x93 & ~x105 & ~x113 & ~x149 & ~x170 & ~x185 & ~x209 & ~x229 & ~x367 & ~x396 & ~x400 & ~x559 & ~x643 & ~x654 & ~x664 & ~x695 & ~x710 & ~x734 & ~x759;
assign c964 =  x218 &  x246 &  x247 &  x330 &  x354 &  x380 &  x386 &  x546 & ~x31 & ~x57 & ~x68 & ~x84 & ~x94 & ~x117 & ~x120 & ~x223 & ~x225 & ~x258 & ~x393 & ~x447 & ~x771;
assign c966 =  x349 &  x376 &  x412 &  x562 &  x598 & ~x50 & ~x59 & ~x106 & ~x140 & ~x144 & ~x197 & ~x225 & ~x311 & ~x341 & ~x645 & ~x678 & ~x683 & ~x686 & ~x688 & ~x743;
assign c968 =  x626 & ~x3 & ~x480 & ~x483 & ~x509 & ~x747;
assign c970 =  x581 &  x584 & ~x115 & ~x126 & ~x129 & ~x155 & ~x176 & ~x177 & ~x192 & ~x362 & ~x400 & ~x617 & ~x720;
assign c972 =  x590;
assign c974 =  x544 &  x586 &  x610 &  x614 & ~x71 & ~x95 & ~x229 & ~x632 & ~x646 & ~x680 & ~x720 & ~x740;
assign c976 = ~x32 & ~x66 & ~x92 & ~x126 & ~x136 & ~x140 & ~x200 & ~x232 & ~x238 & ~x255 & ~x372 & ~x455 & ~x460 & ~x511;
assign c978 =  x350 &  x452 &  x519 &  x543 & ~x29 & ~x84 & ~x347;
assign c980 =  x239 &  x301 &  x304 &  x405 &  x450 &  x451 &  x453 & ~x13 & ~x42 & ~x56 & ~x59 & ~x126 & ~x134 & ~x149 & ~x617 & ~x720;
assign c982 =  x329 &  x438 &  x473 &  x478 &  x488 &  x494 &  x516 &  x540 &  x541 &  x608 & ~x10 & ~x40 & ~x61 & ~x62 & ~x79 & ~x92 & ~x232 & ~x255 & ~x288 & ~x316 & ~x687 & ~x724 & ~x739 & ~x750 & ~x755 & ~x762;
assign c984 =  x235;
assign c986 =  x105 &  x158 &  x496 & ~x27 & ~x64 & ~x396;
assign c988 =  x250 &  x348 &  x350 &  x376;
assign c990 =  x239 &  x240 &  x322 &  x350 &  x377 &  x404 &  x405 &  x484 & ~x45 & ~x57 & ~x59 & ~x153 & ~x587;
assign c992 =  x184 &  x212 &  x218 &  x246 &  x267 &  x328 & ~x12 & ~x121 & ~x197 & ~x335 & ~x396 & ~x763;
assign c994 =  x266 &  x267 &  x330 &  x383 &  x407 &  x417 &  x431 &  x471 &  x484 &  x522 & ~x11 & ~x28 & ~x59 & ~x84 & ~x93 & ~x97 & ~x101 & ~x108 & ~x201 & ~x285 & ~x288 & ~x615 & ~x646 & ~x660 & ~x679 & ~x689 & ~x711 & ~x736 & ~x746 & ~x750 & ~x776 & ~x780;
assign c996 = ~x16 & ~x126 & ~x148 & ~x168 & ~x264 & ~x343 & ~x400 & ~x431 & ~x475 & ~x482 & ~x483 & ~x484 & ~x538;
assign c998 = ~x183 & ~x460 & ~x479 & ~x680;
assign c9100 =  x266 &  x375 & ~x550;
assign c9102 =  x656 & ~x427 & ~x540 & ~x559 & ~x773;
assign c9104 =  x304 &  x305 &  x350 &  x358 &  x443 &  x493 &  x519 &  x546 & ~x12 & ~x129 & ~x135 & ~x136 & ~x153 & ~x185 & ~x209 & ~x235 & ~x282 & ~x291 & ~x364 & ~x401 & ~x646 & ~x654 & ~x657 & ~x744;
assign c9106 =  x160 &  x161 &  x184 &  x187 &  x217 & ~x88 & ~x392;
assign c9108 =  x351 &  x462 &  x494 &  x523 &  x573 & ~x32 & ~x42 & ~x206 & ~x226 & ~x279 & ~x339 & ~x370 & ~x429 & ~x455 & ~x671 & ~x702 & ~x749;
assign c9110 = ~x135 & ~x187 & ~x206 & ~x254 & ~x255 & ~x429 & ~x455;
assign c9112 =  x590 &  x668;
assign c9114 =  x266 &  x348 &  x414 &  x464 &  x599 & ~x11 & ~x24 & ~x34 & ~x59 & ~x312 & ~x315 & ~x662;
assign c9116 =  x293 &  x294 &  x325 &  x333 &  x348 &  x385 & ~x185 & ~x550 & ~x643;
assign c9118 =  x276 &  x301 &  x329 &  x380 &  x467 &  x468 & ~x111 & ~x177 & ~x214 & ~x596 & ~x677 & ~x737 & ~x773;
assign c9120 =  x610 & ~x9 & ~x35 & ~x58 & ~x69 & ~x92 & ~x123 & ~x137 & ~x140 & ~x168 & ~x172 & ~x177 & ~x254 & ~x259 & ~x319 & ~x347 & ~x372 & ~x400 & ~x401 & ~x480 & ~x511 & ~x761 & ~x775;
assign c9122 =  x411 &  x462 &  x496 &  x497 &  x534 &  x573 &  x581 & ~x2 & ~x120 & ~x126 & ~x153 & ~x255 & ~x283 & ~x284 & ~x285 & ~x288 & ~x425 & ~x589 & ~x631 & ~x666 & ~x728 & ~x755;
assign c9124 =  x246 &  x294 &  x322 &  x376 &  x613 & ~x719;
assign c9126 =  x295 &  x303 &  x304 &  x328 &  x383 &  x520 &  x543 & ~x102 & ~x134 & ~x180 & ~x186 & ~x198 & ~x202 & ~x233 & ~x255 & ~x374 & ~x400 & ~x732 & ~x773;
assign c9128 =  x424 &  x450 & ~x179 & ~x577;
assign c9130 = ~x47 & ~x72 & ~x235 & ~x456 & ~x458 & ~x617 & ~x648 & ~x649 & ~x718;
assign c9132 = ~x126 & ~x207 & ~x254 & ~x291 & ~x453 & ~x455 & ~x460 & ~x482 & ~x486 & ~x513 & ~x538;
assign c9134 =  x324 &  x489 &  x562 &  x576 & ~x5 & ~x9 & ~x16 & ~x18 & ~x26 & ~x51 & ~x69 & ~x72 & ~x94 & ~x121 & ~x123 & ~x127 & ~x180 & ~x337 & ~x455 & ~x675 & ~x703 & ~x712 & ~x721 & ~x735 & ~x772;
assign c9136 =  x581 & ~x65 & ~x145 & ~x172 & ~x173 & ~x313 & ~x337 & ~x345 & ~x401 & ~x455 & ~x458 & ~x587;
assign c9138 =  x648;
assign c9140 = ~x55 & ~x70 & ~x214 & ~x233 & ~x282 & ~x566 & ~x568 & ~x596 & ~x617 & ~x736 & ~x746;
assign c9142 =  x304 &  x330 &  x379 & ~x13 & ~x49 & ~x122 & ~x126 & ~x185 & ~x187 & ~x202 & ~x214 & ~x233 & ~x254 & ~x345 & ~x578 & ~x739;
assign c9144 =  x352 &  x414 &  x417 &  x450 &  x453 &  x457 &  x467 &  x468 &  x497 &  x525 &  x543 &  x553 & ~x27 & ~x31 & ~x35 & ~x66 & ~x68 & ~x112 & ~x140 & ~x155 & ~x169 & ~x223 & ~x253 & ~x265 & ~x342 & ~x617 & ~x645 & ~x655 & ~x688 & ~x707 & ~x726 & ~x727;
assign c9146 =  x494 &  x499 &  x500 &  x546 &  x549 &  x573 &  x584 & ~x18 & ~x24 & ~x51 & ~x56 & ~x58 & ~x68 & ~x78 & ~x126 & ~x264 & ~x338 & ~x347 & ~x401 & ~x423 & ~x429 & ~x702 & ~x776;
assign c9148 =  x304 &  x327 &  x480 &  x484 &  x496 &  x541 & ~x153 & ~x172 & ~x179 & ~x257 & ~x259 & ~x281 & ~x504 & ~x596 & ~x599 & ~x602 & ~x655 & ~x689;
assign c9150 =  x387 &  x508 &  x584 & ~x61 & ~x68 & ~x72 & ~x97 & ~x106 & ~x206 & ~x207 & ~x229 & ~x423 & ~x617 & ~x622 & ~x628 & ~x646;
assign c9152 =  x246 &  x249 &  x294 &  x303 &  x330 & ~x98 & ~x118 & ~x120 & ~x140 & ~x161 & ~x204 & ~x234 & ~x341 & ~x649 & ~x771;
assign c9154 = ~x13 & ~x18 & ~x26 & ~x27 & ~x28 & ~x41 & ~x56 & ~x58 & ~x97 & ~x98 & ~x99 & ~x101 & ~x108 & ~x113 & ~x114 & ~x115 & ~x133 & ~x137 & ~x140 & ~x143 & ~x151 & ~x202 & ~x224 & ~x226 & ~x231 & ~x237 & ~x279 & ~x290 & ~x309 & ~x397 & ~x400 & ~x425 & ~x429 & ~x450 & ~x455 & ~x457 & ~x483 & ~x701 & ~x734 & ~x747 & ~x756 & ~x765 & ~x783;
assign c9156 =  x249 &  x441 &  x488 & ~x175 & ~x262 & ~x596 & ~x599 & ~x743;
assign c9158 = ~x33 & ~x81 & ~x87 & ~x117 & ~x118 & ~x140 & ~x143 & ~x179 & ~x195 & ~x200 & ~x205 & ~x288 & ~x311 & ~x344 & ~x401 & ~x429 & ~x453 & ~x454 & ~x455 & ~x480 & ~x481 & ~x484 & ~x485 & ~x567 & ~x746;
assign c9160 =  x348 &  x543 &  x613 & ~x1 & ~x46 & ~x94 & ~x97 & ~x112 & ~x126 & ~x233 & ~x260 & ~x703 & ~x750 & ~x756 & ~x762;
assign c9162 =  x376 &  x429 &  x456 & ~x84 & ~x90 & ~x113 & ~x185 & ~x563 & ~x568 & ~x583 & ~x597 & ~x683 & ~x705;
assign c9164 =  x383 &  x387 &  x496 &  x530 &  x543 &  x546 &  x553 &  x556 &  x584 &  x585 & ~x27 & ~x58 & ~x90 & ~x95 & ~x106 & ~x125 & ~x145 & ~x150 & ~x230 & ~x338 & ~x342 & ~x364 & ~x393 & ~x400 & ~x633 & ~x688 & ~x704 & ~x713 & ~x720;
assign c9166 =  x526 &  x542 &  x558 &  x585 &  x586 & ~x6 & ~x31 & ~x56 & ~x126 & ~x146 & ~x150 & ~x223 & ~x233 & ~x396 & ~x590 & ~x623 & ~x633 & ~x648 & ~x651 & ~x655 & ~x683 & ~x743;
assign c9168 =  x163 &  x219 &  x246 &  x247;
assign c9170 =  x247 &  x383 &  x411 &  x441 &  x521 &  x522 &  x552 &  x573 & ~x76 & ~x87 & ~x88 & ~x93 & ~x97 & ~x112 & ~x229 & ~x260 & ~x311 & ~x372 & ~x429 & ~x448 & ~x755;
assign c9172 =  x47;
assign c9174 = ~x445 & ~x498 & ~x746;
assign c9176 =  x296 &  x304 &  x328 &  x333 &  x355 &  x385 &  x387 &  x388 &  x443 &  x446 &  x507 &  x520 &  x558 & ~x6 & ~x61 & ~x62 & ~x81 & ~x112 & ~x126 & ~x136 & ~x153 & ~x160 & ~x206 & ~x374 & ~x401 & ~x717 & ~x723;
assign c9178 =  x246 &  x247 &  x298 &  x384 &  x489 &  x536 &  x552 &  x567 &  x585 &  x611 & ~x58 & ~x78 & ~x89 & ~x122 & ~x170 & ~x171 & ~x204 & ~x233 & ~x289 & ~x363 & ~x365 & ~x367 & ~x709 & ~x719 & ~x730 & ~x747 & ~x748 & ~x777;
assign c9180 =  x267 &  x326 &  x354 &  x415 &  x438 &  x517 &  x518 & ~x6 & ~x24 & ~x28 & ~x31 & ~x36 & ~x37 & ~x59 & ~x113 & ~x148 & ~x199 & ~x223 & ~x258 & ~x281 & ~x288 & ~x314 & ~x362 & ~x372 & ~x419 & ~x475 & ~x717 & ~x758 & ~x783;
assign c9182 =  x452 &  x521 &  x523 &  x526 &  x556 & ~x13 & ~x47 & ~x56 & ~x74 & ~x87 & ~x96 & ~x142 & ~x167 & ~x176 & ~x202 & ~x210 & ~x257 & ~x291 & ~x311 & ~x319 & ~x373 & ~x655 & ~x672 & ~x771;
assign c9184 =  x19;
assign c9186 = ~x170 & ~x343 & ~x445 & ~x455 & ~x507 & ~x539 & ~x540;
assign c9188 =  x239 &  x267 &  x350 &  x450 &  x451 &  x452 & ~x56 & ~x72 & ~x127 & ~x144 & ~x775;
assign c9190 = ~x9 & ~x62 & ~x291 & ~x334 & ~x432 & ~x454 & ~x484 & ~x511 & ~x729;
assign c9192 =  x212 &  x706;
assign c9194 =  x299 &  x354 &  x575 & ~x56 & ~x92 & ~x115 & ~x138 & ~x150 & ~x204 & ~x373 & ~x427 & ~x452 & ~x455 & ~x479 & ~x482 & ~x483 & ~x615 & ~x727 & ~x746 & ~x775;
assign c9196 =  x424 & ~x578;
assign c9198 =  x558 & ~x174 & ~x185 & ~x578 & ~x611 & ~x613 & ~x721;
assign c9200 =  x452 &  x467 &  x518 & ~x44 & ~x92 & ~x136 & ~x187 & ~x201 & ~x214 & ~x215 & ~x248 & ~x319 & ~x337 & ~x344 & ~x345 & ~x587 & ~x596 & ~x602 & ~x649 & ~x719;
assign c9202 =  x304 &  x375 &  x387 &  x401 &  x546 &  x572 & ~x7 & ~x32 & ~x74 & ~x121 & ~x206 & ~x724 & ~x750 & ~x771 & ~x776;
assign c9204 =  x216 &  x436 &  x598 &  x611 &  x629;
assign c9206 =  x295 &  x350 &  x411 &  x513 &  x522 &  x527 &  x541 &  x561 &  x585 & ~x51 & ~x97 & ~x108 & ~x110 & ~x256 & ~x732 & ~x755 & ~x759 & ~x776;
assign c9208 =  x351 &  x517 &  x545 &  x583 &  x584 & ~x56 & ~x84 & ~x98 & ~x346 & ~x366 & ~x400 & ~x634 & ~x643 & ~x675 & ~x695;
assign c9210 = ~x433 & ~x453 & ~x457 & ~x482 & ~x483 & ~x679;
assign c9212 =  x239 &  x450 &  x542 & ~x56 & ~x188 & ~x713;
assign c9214 = ~x31 & ~x57 & ~x68 & ~x119 & ~x125 & ~x170 & ~x177 & ~x198 & ~x201 & ~x236 & ~x258 & ~x263 & ~x396 & ~x427 & ~x509 & ~x510 & ~x511 & ~x559 & ~x746 & ~x762 & ~x773 & ~x780;
assign c9216 = ~x21 & ~x58 & ~x85 & ~x118 & ~x126 & ~x136 & ~x206 & ~x262 & ~x288 & ~x319 & ~x334 & ~x340 & ~x362 & ~x371 & ~x511 & ~x772;
assign c9218 =  x266 &  x484 &  x543 &  x547 & ~x59 & ~x65 & ~x112 & ~x169 & ~x284;
assign c9220 =  x384 &  x545 &  x571 &  x653 & ~x337 & ~x482 & ~x643;
assign c9222 = ~x30 & ~x34 & ~x62 & ~x84 & ~x94 & ~x123 & ~x167 & ~x190 & ~x225 & ~x287 & ~x317 & ~x394 & ~x417 & ~x426 & ~x427 & ~x448 & ~x513 & ~x745;
assign c9224 =  x219 &  x245 &  x246 &  x247 &  x324 &  x376 &  x539 & ~x36 & ~x56 & ~x70 & ~x167 & ~x204 & ~x205 & ~x313 & ~x729 & ~x755 & ~x761;
assign c9226 =  x222 &  x353 &  x383 &  x467 & ~x12 & ~x27 & ~x44 & ~x45 & ~x56 & ~x61 & ~x127 & ~x151 & ~x225 & ~x235 & ~x365 & ~x710 & ~x718 & ~x741 & ~x772;
assign c9228 = ~x8 & ~x38 & ~x53 & ~x90 & ~x91 & ~x93 & ~x170 & ~x180 & ~x203 & ~x226 & ~x311 & ~x316 & ~x319 & ~x336 & ~x338 & ~x362 & ~x395 & ~x453 & ~x455 & ~x456 & ~x480 & ~x481 & ~x540 & ~x776 & ~x777;
assign c9230 = ~x140 & ~x177 & ~x182 & ~x202 & ~x311 & ~x393 & ~x514 & ~x515 & ~x538 & ~x569;
assign c9232 =  x348 &  x349 &  x520 &  x546 &  x598 &  x613 & ~x0 & ~x58 & ~x112 & ~x144 & ~x147 & ~x170 & ~x195 & ~x202 & ~x233 & ~x338 & ~x364 & ~x397 & ~x448 & ~x643 & ~x688 & ~x720 & ~x740 & ~x744 & ~x746 & ~x766 & ~x767 & ~x772;
assign c9234 =  x249 &  x272 &  x328 &  x411 &  x500 &  x501 &  x520 &  x540 &  x543 &  x573 & ~x7 & ~x40 & ~x45 & ~x64 & ~x75 & ~x92 & ~x106 & ~x128 & ~x146 & ~x159 & ~x168 & ~x173 & ~x177 & ~x182 & ~x206 & ~x291 & ~x343 & ~x713 & ~x719 & ~x723 & ~x730;
assign c9236 =  x410 &  x517 & ~x58 & ~x61 & ~x150 & ~x184 & ~x185 & ~x229 & ~x234 & ~x315 & ~x400 & ~x401 & ~x628 & ~x766;
assign c9238 =  x354 &  x435 &  x507 &  x585 & ~x56 & ~x136 & ~x143 & ~x169 & ~x373 & ~x396 & ~x617;
assign c9240 = ~x58 & ~x374 & ~x427 & ~x431 & ~x483 & ~x484 & ~x567;
assign c9242 =  x184 &  x212 &  x239 &  x614;
assign c9244 =  x329 &  x452 & ~x191 & ~x566 & ~x567 & ~x596 & ~x597 & ~x599 & ~x611 & ~x622;
assign c9246 =  x295 &  x414 &  x544 &  x545 &  x546 &  x597 &  x655 & ~x115 & ~x223 & ~x744;
assign c9248 =  x607 & ~x429 & ~x457 & ~x480;
assign c9250 =  x414 &  x473 &  x517 &  x530 & ~x54 & ~x56 & ~x58 & ~x71 & ~x121 & ~x134 & ~x158 & ~x185 & ~x193 & ~x209 & ~x214 & ~x215 & ~x218 & ~x316 & ~x623 & ~x654 & ~x676 & ~x677 & ~x682 & ~x721 & ~x753 & ~x762;
assign c9252 =  x158 &  x186 &  x187 &  x188 &  x218 &  x246 &  x355 & ~x1 & ~x3 & ~x4 & ~x34 & ~x56 & ~x60 & ~x90 & ~x142 & ~x231 & ~x256 & ~x284;
assign c9254 =  x184 &  x187 &  x218 &  x247 &  x299 & ~x10 & ~x29 & ~x45 & ~x59 & ~x99 & ~x339;
assign c9256 =  x219 &  x241 &  x246 &  x247 &  x304 &  x383 &  x405 &  x444 &  x488 &  x516 &  x522 & ~x43 & ~x68 & ~x79 & ~x88 & ~x118 & ~x144 & ~x171 & ~x229 & ~x233 & ~x342 & ~x363 & ~x702 & ~x741;
assign c9258 =  x239 &  x350 &  x450 &  x452 &  x538 & ~x56 & ~x136 & ~x765;
assign c9260 =  x350 &  x405 &  x493 &  x497 &  x545 &  x584 & ~x3 & ~x49 & ~x102 & ~x125 & ~x136 & ~x167 & ~x197 & ~x201 & ~x254 & ~x363 & ~x631 & ~x643 & ~x646 & ~x655 & ~x677 & ~x707 & ~x737;
assign c9262 =  x248 &  x415 &  x467 &  x543 &  x545 &  x590 &  x613 & ~x27 & ~x31 & ~x33 & ~x35 & ~x36 & ~x89 & ~x120 & ~x143 & ~x256 & ~x310 & ~x367 & ~x727;
assign c9264 =  x450 &  x452 &  x453 & ~x9 & ~x185 & ~x188 & ~x566 & ~x596;
assign c9266 =  x274 &  x450 &  x452 & ~x161;
assign c9268 =  x322 & ~x122 & ~x262 & ~x319 & ~x400 & ~x427 & ~x481 & ~x482;
assign c9270 =  x698;
assign c9272 = ~x35 & ~x53 & ~x90 & ~x198 & ~x229 & ~x268 & ~x307 & ~x391 & ~x400 & ~x514 & ~x689 & ~x741 & ~x742 & ~x761 & ~x766 & ~x770;
assign c9274 =  x293 &  x348 & ~x84 & ~x549 & ~x755;
assign c9276 =  x218 &  x219 &  x358 &  x548 &  x562 &  x573 & ~x3 & ~x12 & ~x17 & ~x33 & ~x56 & ~x83 & ~x87 & ~x112 & ~x114 & ~x118 & ~x143 & ~x144 & ~x171 & ~x202 & ~x338 & ~x364 & ~x365 & ~x419 & ~x767;
assign c9278 =  x266 &  x267 &  x449 &  x450 &  x451 & ~x112 & ~x173;
assign c9280 =  x300 &  x462 &  x467 &  x493 &  x519 &  x536 &  x608 &  x611 &  x612 &  x613 &  x614 & ~x0 & ~x1 & ~x5 & ~x11 & ~x24 & ~x27 & ~x29 & ~x36 & ~x42 & ~x51 & ~x53 & ~x56 & ~x67 & ~x70 & ~x81 & ~x93 & ~x94 & ~x99 & ~x101 & ~x105 & ~x108 & ~x114 & ~x120 & ~x196 & ~x198 & ~x202 & ~x226 & ~x234 & ~x253 & ~x280 & ~x338 & ~x369 & ~x633 & ~x649 & ~x658 & ~x660 & ~x688 & ~x724 & ~x728 & ~x750 & ~x763;
assign c9282 = ~x13 & ~x38 & ~x41 & ~x135 & ~x157 & ~x210 & ~x368 & ~x427 & ~x433 & ~x482 & ~x765;
assign c9284 =  x620 &  x657;
assign c9286 =  x352 &  x383 &  x496 &  x507 & ~x29 & ~x122 & ~x169 & ~x206 & ~x207 & ~x226 & ~x284 & ~x455 & ~x632 & ~x660 & ~x759;
assign c9288 =  x302 &  x304 &  x333 &  x389 &  x444 &  x493 &  x496 &  x499 &  x541 &  x544 &  x545 &  x557 & ~x8 & ~x52 & ~x57 & ~x59 & ~x64 & ~x112 & ~x149 & ~x162 & ~x182 & ~x205 & ~x223 & ~x233 & ~x259 & ~x291 & ~x420 & ~x604 & ~x616 & ~x673 & ~x686 & ~x704 & ~x726 & ~x737 & ~x764;
assign c9290 =  x245 &  x246 &  x247 &  x248 &  x330 &  x411 &  x500 &  x516 &  x542 &  x544 & ~x2 & ~x31 & ~x64 & ~x94 & ~x102 & ~x106 & ~x126 & ~x129 & ~x130 & ~x134 & ~x200 & ~x290 & ~x315 & ~x336 & ~x346 & ~x559 & ~x617 & ~x646 & ~x648 & ~x679 & ~x682 & ~x702 & ~x713 & ~x732 & ~x756 & ~x762 & ~x768 & ~x776;
assign c9292 =  x184 &  x185 &  x212 &  x271 &  x353 &  x463 &  x543 &  x626 & ~x11 & ~x29 & ~x36 & ~x59 & ~x93 & ~x119 & ~x204 & ~x258 & ~x281 & ~x308 & ~x341 & ~x420 & ~x616 & ~x730 & ~x759;
assign c9294 =  x247 &  x519 &  x572 & ~x66 & ~x93 & ~x101 & ~x126 & ~x342 & ~x429 & ~x455 & ~x746 & ~x767;
assign c9296 =  x546 &  x548 &  x652 &  x653 &  x655 &  x657 & ~x1 & ~x27 & ~x55 & ~x88 & ~x197 & ~x223 & ~x255 & ~x288 & ~x315 & ~x341 & ~x371 & ~x393 & ~x761;
assign c9298 =  x350 &  x482 & ~x55 & ~x115 & ~x130 & ~x132 & ~x168 & ~x185 & ~x227 & ~x283 & ~x549;
assign c9300 =  x158 &  x159 &  x160 & ~x63 & ~x340 & ~x761;
assign c9302 =  x581 & ~x34 & ~x202 & ~x431 & ~x455 & ~x456 & ~x457 & ~x482;
assign c9304 =  x328 &  x354 &  x358 &  x380 &  x383 &  x389 &  x569 &  x570 &  x573 &  x585 &  x586 & ~x27 & ~x28 & ~x56 & ~x59 & ~x72 & ~x81 & ~x97 & ~x122 & ~x136 & ~x153 & ~x167 & ~x174 & ~x226 & ~x648 & ~x703 & ~x707 & ~x717 & ~x720 & ~x743 & ~x773;
assign c9306 =  x323 &  x474 &  x586 & ~x179 & ~x185 & ~x311 & ~x606 & ~x617 & ~x687 & ~x695 & ~x703;
assign c9308 =  x247 &  x487 &  x507 &  x520 &  x608 &  x610 & ~x0 & ~x37 & ~x44 & ~x62 & ~x82 & ~x99 & ~x108 & ~x121 & ~x126 & ~x138 & ~x142 & ~x145 & ~x196 & ~x225 & ~x280 & ~x309 & ~x311 & ~x342 & ~x448 & ~x717 & ~x765 & ~x766 & ~x771 & ~x783;
assign c9310 =  x579 & ~x0 & ~x1 & ~x64 & ~x84 & ~x90 & ~x203 & ~x338 & ~x367 & ~x427 & ~x429 & ~x448 & ~x455 & ~x456 & ~x479 & ~x480 & ~x482 & ~x483 & ~x484 & ~x508 & ~x727 & ~x757;
assign c9312 = ~x16 & ~x18 & ~x24 & ~x88 & ~x154 & ~x207 & ~x225 & ~x257 & ~x262 & ~x307 & ~x366 & ~x392 & ~x433 & ~x455 & ~x742 & ~x765 & ~x775;
assign c9314 =  x194 &  x467 &  x500 &  x520 &  x523 &  x528 & ~x15 & ~x35 & ~x68 & ~x97 & ~x108 & ~x126 & ~x145 & ~x223 & ~x229 & ~x257 & ~x259 & ~x291 & ~x342 & ~x420 & ~x476 & ~x706 & ~x744 & ~x776;
assign c9316 =  x222 &  x385 &  x406 & ~x7 & ~x12 & ~x42 & ~x93 & ~x98 & ~x100 & ~x112 & ~x123 & ~x232 & ~x254 & ~x314 & ~x315 & ~x718 & ~x758;
assign c9318 =  x493 &  x573 & ~x6 & ~x56 & ~x59 & ~x62 & ~x66 & ~x67 & ~x87 & ~x97 & ~x102 & ~x106 & ~x122 & ~x123 & ~x140 & ~x148 & ~x223 & ~x291 & ~x345 & ~x392 & ~x429 & ~x453 & ~x455 & ~x476 & ~x617 & ~x748 & ~x753 & ~x770;
assign c9320 =  x239 &  x246 &  x450;
assign c9322 =  x301 &  x348 &  x387 &  x473 & ~x7 & ~x70 & ~x84 & ~x225 & ~x254 & ~x577 & ~x578 & ~x722 & ~x735 & ~x750 & ~x769;
assign c9324 =  x246 &  x274 &  x330 &  x331 &  x358 &  x666 & ~x67 & ~x112 & ~x122 & ~x141 & ~x199 & ~x280 & ~x317 & ~x338 & ~x341 & ~x760;
assign c9326 =  x579 & ~x27 & ~x38 & ~x95 & ~x112 & ~x118 & ~x173 & ~x232 & ~x431 & ~x588;
assign c9328 = ~x1 & ~x10 & ~x28 & ~x40 & ~x63 & ~x70 & ~x84 & ~x143 & ~x155 & ~x210 & ~x225 & ~x227 & ~x262 & ~x344 & ~x396 & ~x401 & ~x424 & ~x429 & ~x431 & ~x455 & ~x457 & ~x482 & ~x484 & ~x756 & ~x759;
assign c9330 =  x377 &  x521 &  x620 & ~x34 & ~x55 & ~x65 & ~x141 & ~x170 & ~x174 & ~x201 & ~x226 & ~x259 & ~x341 & ~x422 & ~x426 & ~x731 & ~x758;
assign c9332 =  x608 &  x609 &  x610 & ~x92 & ~x198 & ~x281 & ~x394 & ~x397 & ~x458 & ~x482;
assign c9334 =  x618 &  x654 &  x655 & ~x10 & ~x33 & ~x67 & ~x90 & ~x145 & ~x198 & ~x308 & ~x427 & ~x504 & ~x770;
assign c9336 = ~x83 & ~x97 & ~x123 & ~x214 & ~x282 & ~x393 & ~x401 & ~x617 & ~x640 & ~x668;
assign c9338 =  x388 &  x523 & ~x29 & ~x54 & ~x87 & ~x90 & ~x100 & ~x120 & ~x126 & ~x129 & ~x132 & ~x138 & ~x185 & ~x215 & ~x401 & ~x721 & ~x738 & ~x771;
assign c9340 = ~x82 & ~x108 & ~x131 & ~x136 & ~x140 & ~x144 & ~x150 & ~x167 & ~x170 & ~x206 & ~x226 & ~x234 & ~x318 & ~x427 & ~x449 & ~x455 & ~x480 & ~x483 & ~x484 & ~x508 & ~x509 & ~x510 & ~x511 & ~x773;
assign c9342 =  x493 & ~x8 & ~x185 & ~x214 & ~x599 & ~x634;
assign c9344 = ~x24 & ~x73 & ~x83 & ~x205 & ~x264 & ~x281 & ~x433 & ~x455 & ~x509;
assign c9346 =  x304 &  x383 &  x591 &  x624 & ~x58 & ~x59 & ~x125 & ~x150 & ~x284 & ~x634 & ~x716 & ~x780;
assign c9348 =  x300 &  x348 &  x358 &  x376 &  x417 &  x540 &  x542 &  x557 & ~x43 & ~x56 & ~x84 & ~x112 & ~x153 & ~x179 & ~x646 & ~x713;
assign c9350 = ~x3 & ~x123 & ~x129 & ~x183 & ~x209 & ~x291 & ~x345 & ~x391 & ~x508 & ~x510 & ~x511 & ~x690 & ~x703 & ~x712 & ~x719 & ~x772;
assign c9352 =  x664 & ~x23 & ~x79 & ~x149 & ~x173 & ~x179 & ~x308;
assign c9354 =  x478 &  x500 &  x534 &  x558 &  x575 & ~x34 & ~x71 & ~x97 & ~x98 & ~x229 & ~x257 & ~x315 & ~x392 & ~x588 & ~x690 & ~x695 & ~x713;
assign c9356 =  x441 &  x591 &  x626 & ~x60 & ~x119 & ~x226 & ~x311 & ~x362 & ~x448 & ~x644 & ~x776;
assign c9358 =  x184 &  x246 &  x247 &  x300 &  x304 &  x472 &  x520 &  x584 & ~x4 & ~x13 & ~x335 & ~x729 & ~x759;
assign c9360 = ~x26 & ~x61 & ~x117 & ~x169 & ~x170 & ~x199 & ~x309 & ~x446 & ~x452 & ~x480 & ~x482 & ~x540 & ~x690;
assign c9362 =  x376 &  x608 &  x610 &  x614 & ~x105 & ~x560 & ~x779;
assign c9364 =  x648 &  x678;
assign c9366 =  x451 &  x586;
assign c9368 =  x406 &  x409 &  x462 &  x499 &  x503 &  x531 & ~x36 & ~x58 & ~x99 & ~x141 & ~x144 & ~x197 & ~x207 & ~x231 & ~x392 & ~x737;
assign c9370 = ~x16 & ~x43 & ~x101 & ~x125 & ~x136 & ~x137 & ~x144 & ~x150 & ~x175 & ~x311 & ~x318 & ~x419 & ~x508 & ~x509 & ~x510 & ~x511 & ~x587;
assign c9372 =  x217 &  x244 &  x246 &  x247 &  x248 &  x275 &  x302 &  x325 &  x499 &  x541 &  x574 &  x584 & ~x1 & ~x5 & ~x79 & ~x87 & ~x96 & ~x148 & ~x149 & ~x307 & ~x312 & ~x363 & ~x364 & ~x707 & ~x763 & ~x776;
assign c9374 =  x293 &  x405 &  x466 &  x585 &  x586 & ~x39 & ~x40 & ~x47 & ~x68 & ~x80 & ~x93 & ~x150 & ~x176 & ~x196 & ~x252 & ~x313 & ~x677 & ~x721 & ~x773 & ~x774;
assign c9376 = ~x289 & ~x474 & ~x511 & ~x529;
assign c9378 =  x248 &  x295 &  x405 &  x543 & ~x59 & ~x172 & ~x563;
assign c9380 =  x333 &  x452 & ~x93 & ~x292 & ~x401 & ~x717;
assign c9382 = ~x8 & ~x34 & ~x56 & ~x112 & ~x176 & ~x193 & ~x225 & ~x259 & ~x342 & ~x400 & ~x486 & ~x510 & ~x511 & ~x513 & ~x736 & ~x775;
assign c9384 =  x266 &  x295 &  x303 &  x330 &  x377 &  x446 &  x480 & ~x98 & ~x136 & ~x587 & ~x658;
assign c9386 = ~x9 & ~x83 & ~x101 & ~x508 & ~x540 & ~x546 & ~x596;
assign c9388 =  x273 &  x302 &  x303 &  x330 &  x333 &  x383 &  x484 &  x497 & ~x42 & ~x68 & ~x106 & ~x140 & ~x144 & ~x153 & ~x174 & ~x176 & ~x179 & ~x185 & ~x191 & ~x207 & ~x288 & ~x504 & ~x594 & ~x603 & ~x613 & ~x713 & ~x765;
assign c9390 =  x212 &  x239 &  x246 &  x248 &  x460 &  x496 &  x500 & ~x1 & ~x2 & ~x10 & ~x54 & ~x57 & ~x99 & ~x173 & ~x227 & ~x424 & ~x588 & ~x615;
assign c9392 =  x579 & ~x318 & ~x429 & ~x455 & ~x457 & ~x479 & ~x482 & ~x510;
assign c9394 =  x158 &  x159 &  x160 & ~x339 & ~x482;
assign c9396 =  x250 & ~x9 & ~x578;
assign c9398 =  x475 &  x531;
assign c9400 =  x333 &  x478 &  x507 &  x558 &  x584 & ~x43 & ~x51 & ~x72 & ~x100 & ~x108 & ~x123 & ~x126 & ~x129 & ~x176 & ~x207 & ~x233 & ~x288 & ~x338 & ~x345 & ~x713 & ~x727 & ~x772;
assign c9402 =  x246 &  x387 &  x497 & ~x145 & ~x256 & ~x281 & ~x309 & ~x362 & ~x390 & ~x418 & ~x761;
assign c9404 =  x193 &  x216 &  x249;
assign c9406 =  x184 &  x212 &  x267 &  x294 &  x322 & ~x174 & ~x229 & ~x688;
assign c9408 =  x350 &  x378 &  x383 &  x386 &  x433 &  x490 &  x510 &  x517 & ~x27 & ~x93 & ~x126 & ~x136 & ~x146 & ~x185 & ~x191 & ~x214 & ~x368 & ~x563 & ~x604 & ~x695;
assign c9410 =  x271 &  x326 & ~x37 & ~x66 & ~x83 & ~x95 & ~x136 & ~x137 & ~x149 & ~x164 & ~x201 & ~x254 & ~x310 & ~x340 & ~x342 & ~x364 & ~x451 & ~x510 & ~x511 & ~x758;
assign c9412 =  x296 &  x300 &  x301 &  x303 &  x328 &  x382 &  x404 &  x477 &  x507 &  x513 &  x519 & ~x3 & ~x13 & ~x35 & ~x55 & ~x185 & ~x188 & ~x206 & ~x318 & ~x319 & ~x605 & ~x617 & ~x644 & ~x661 & ~x687 & ~x705 & ~x713 & ~x743 & ~x775 & ~x776 & ~x778;
assign c9414 =  x212 &  x246 &  x247 &  x248 &  x350 &  x376 &  x404 &  x456 & ~x56 & ~x112 & ~x204 & ~x232 & ~x677 & ~x736 & ~x739 & ~x744;
assign c9416 =  x267 &  x348 &  x380 &  x516 &  x571 &  x611 & ~x9 & ~x12 & ~x109 & ~x115 & ~x117 & ~x120 & ~x224 & ~x420 & ~x776;
assign c9418 =  x378 &  x655 &  x677;
assign c9420 =  x296 &  x326 &  x350 &  x380 &  x417 &  x494 &  x500 & ~x72 & ~x99 & ~x102 & ~x105 & ~x106 & ~x112 & ~x134 & ~x176 & ~x189 & ~x258 & ~x560 & ~x578 & ~x587 & ~x596 & ~x628 & ~x713 & ~x721 & ~x735;
assign c9422 =  x294 &  x385 & ~x550 & ~x567 & ~x578 & ~x596;
assign c9424 =  x276 &  x301 &  x302 &  x303 &  x328 &  x405 &  x457 &  x499 & ~x22 & ~x27 & ~x59 & ~x68 & ~x102 & ~x122 & ~x184 & ~x185 & ~x214 & ~x290 & ~x646 & ~x695 & ~x719 & ~x735 & ~x750;
assign c9426 =  x405 &  x458 &  x474 & ~x7 & ~x9 & ~x129 & ~x136 & ~x169 & ~x213 & ~x242 & ~x260 & ~x651 & ~x702 & ~x707;
assign c9428 = ~x10 & ~x152 & ~x291 & ~x453 & ~x454 & ~x460 & ~x483 & ~x699 & ~x727 & ~x776;
assign c9430 =  x735;
assign c9432 =  x608 &  x610 &  x611 & ~x1 & ~x3 & ~x12 & ~x17 & ~x29 & ~x39 & ~x43 & ~x72 & ~x85 & ~x95 & ~x101 & ~x134 & ~x145 & ~x150 & ~x179 & ~x199 & ~x229 & ~x259 & ~x315 & ~x342 & ~x362 & ~x390 & ~x423 & ~x424 & ~x560 & ~x617 & ~x730 & ~x742 & ~x744 & ~x758 & ~x776 & ~x779 & ~x780;
assign c9434 =  x72;
assign c9436 = ~x86 & ~x115 & ~x138 & ~x167 & ~x168 & ~x170 & ~x193 & ~x229 & ~x255 & ~x258 & ~x311 & ~x427 & ~x428 & ~x453 & ~x454 & ~x455 & ~x556 & ~x746 & ~x776;
assign c9438 =  x353 &  x462 &  x500 &  x548 &  x569 &  x584 & ~x17 & ~x135 & ~x151 & ~x196 & ~x200 & ~x229 & ~x372 & ~x395 & ~x419 & ~x429 & ~x454 & ~x455 & ~x762 & ~x773;
assign c9440 =  x247 &  x350 & ~x578 & ~x631 & ~x720;
assign c9442 =  x350 &  x376 &  x440 &  x450 &  x452 &  x467 & ~x9 & ~x25 & ~x61 & ~x68 & ~x136 & ~x174 & ~x284 & ~x345 & ~x655 & ~x703 & ~x770;
assign c9444 =  x376 &  x544 &  x619 &  x620 & ~x53 & ~x343 & ~x344;
assign c9446 =  x376 &  x488 &  x494 &  x533 &  x608 &  x610 &  x611 &  x614 & ~x29 & ~x44 & ~x71 & ~x79 & ~x84 & ~x97 & ~x126 & ~x144 & ~x336 & ~x727 & ~x767;
assign c9448 =  x618 &  x627 &  x629 &  x656;
assign c9450 =  x274 &  x296 &  x354 &  x450 &  x451 &  x452 &  x484 &  x497 &  x505 &  x506 &  x507 &  x517 &  x541 & ~x655 & ~x688 & ~x707;
assign c9452 =  x417 &  x462 &  x467 &  x620 &  x641 & ~x50 & ~x288 & ~x730;
assign c9454 =  x694 & ~x251 & ~x365;
assign c9456 =  x714 & ~x510;
assign c9458 =  x424 & ~x92 & ~x144 & ~x207 & ~x577 & ~x632;
assign c9460 =  x581 & ~x42 & ~x307 & ~x454 & ~x455 & ~x510;
assign c9462 = ~x103 & ~x104 & ~x205 & ~x206 & ~x397 & ~x401 & ~x487 & ~x514 & ~x537;
assign c9464 =  x329 &  x574 & ~x6 & ~x24 & ~x32 & ~x33 & ~x84 & ~x115 & ~x137 & ~x146 & ~x225 & ~x393 & ~x476 & ~x509 & ~x510 & ~x770 & ~x775;
assign c9466 =  x246 &  x247 &  x299 &  x304 &  x326 &  x354 &  x385 &  x461 &  x493 &  x520 &  x544 &  x574 & ~x0 & ~x27 & ~x30 & ~x33 & ~x34 & ~x65 & ~x112 & ~x114 & ~x120 & ~x139 & ~x168 & ~x169 & ~x171 & ~x223 & ~x309 & ~x317 & ~x344 & ~x449 & ~x450 & ~x453 & ~x454 & ~x475 & ~x720 & ~x772;
assign c9468 =  x266 &  x348 &  x436 &  x518 &  x543 & ~x34 & ~x61 & ~x112 & ~x177 & ~x229 & ~x342 & ~x531 & ~x587 & ~x722 & ~x730 & ~x776;
assign c9470 =  x214 &  x216 &  x218 &  x219 &  x244 &  x246 &  x247 &  x296 &  x301 &  x328 &  x416 &  x417 &  x434 &  x443 &  x464 &  x471 &  x514 & ~x25 & ~x43 & ~x58 & ~x68 & ~x70 & ~x81 & ~x84 & ~x93 & ~x149 & ~x170 & ~x175 & ~x315 & ~x338 & ~x504 & ~x688 & ~x709 & ~x720 & ~x721 & ~x726 & ~x727 & ~x728 & ~x735 & ~x758 & ~x780;
assign c9472 =  x249 &  x303 &  x304 &  x380 &  x469 &  x534 &  x545 & ~x11 & ~x108 & ~x179 & ~x223 & ~x291;
assign c9474 =  x249 &  x493 &  x584 &  x611 &  x612 &  x614 & ~x15 & ~x34 & ~x54 & ~x63 & ~x68 & ~x77 & ~x95 & ~x97 & ~x112 & ~x169 & ~x171 & ~x206 & ~x227 & ~x285 & ~x286 & ~x335 & ~x646 & ~x674 & ~x689 & ~x703 & ~x704 & ~x718 & ~x720 & ~x734 & ~x735 & ~x742 & ~x748 & ~x755 & ~x769 & ~x772 & ~x778;
assign c9476 =  x322 &  x656 & ~x81 & ~x201 & ~x205 & ~x223 & ~x232 & ~x369 & ~x398 & ~x727;
assign c9478 =  x302 &  x350 &  x353 &  x383 &  x387 &  x493 &  x526 &  x527 &  x553 & ~x58 & ~x59 & ~x93 & ~x112 & ~x129 & ~x136 & ~x137 & ~x179 & ~x206 & ~x226 & ~x374 & ~x427 & ~x617 & ~x630 & ~x634 & ~x713 & ~x718 & ~x765;
assign c9480 =  x350 &  x507 &  x519 &  x563 &  x614 & ~x23 & ~x62 & ~x167 & ~x226 & ~x364 & ~x678 & ~x709 & ~x726 & ~x756 & ~x772;
assign c9482 =  x411 &  x533 &  x534 &  x555 &  x556 &  x585 &  x586 & ~x6 & ~x35 & ~x136 & ~x654 & ~x657 & ~x720 & ~x740;
assign c9484 =  x422 & ~x225;
assign c9486 = ~x102 & ~x179 & ~x225 & ~x254 & ~x482 & ~x565;
assign c9488 = ~x174 & ~x179 & ~x429 & ~x454 & ~x482 & ~x485 & ~x513 & ~x537 & ~x538 & ~x540;
assign c9490 =  x302 &  x405 &  x502 & ~x6 & ~x43 & ~x54 & ~x125 & ~x129 & ~x223 & ~x292 & ~x318 & ~x400 & ~x628 & ~x664 & ~x735;
assign c9492 =  x608 & ~x84 & ~x224 & ~x230 & ~x252 & ~x373 & ~x390 & ~x482 & ~x745;
assign c9494 =  x98 &  x706;
assign c9496 =  x247 &  x266 &  x295 &  x322 &  x330 &  x358 &  x381 &  x493 &  x517 &  x545 & ~x33 & ~x112;
assign c9498 =  x184 &  x380 &  x387 &  x410 &  x737 & ~x198 & ~x307 & ~x315;
assign c91 =  x344;
assign c95 = ~x353 & ~x461;
assign c97 =  x445 & ~x377 & ~x403 & ~x579;
assign c99 =  x143;
assign c911 =  x191 & ~x353;
assign c913 =  x373 & ~x301;
assign c915 = ~x527;
assign c917 = ~x414;
assign c919 =  x399 & ~x301;
assign c921 = ~x410;
assign c923 =  x314;
assign c925 =  x112;
assign c927 = ~x299 & ~x612;
assign c929 =  x6;
assign c931 =  x230;
assign c933 =  x64;
assign c935 =  x92;
assign c937 =  x630 & ~x295;
assign c939 =  x144;
assign c941 =  x335;
assign c943 = ~x353 & ~x354 & ~x506;
assign c945 = ~x300 & ~x543 & ~x551 & ~x663;
assign c951 =  x85;
assign c953 =  x340;
assign c955 =  x339;
assign c957 =  x359 &  x381 & ~x301;
assign c959 =  x259;
assign c961 =  x410 &  x623 &  x634 &  x636 & ~x294;
assign c963 =  x372 &  x477 & ~x211;
assign c965 =  x232;
assign c967 =  x70;
assign c969 =  x24;
assign c971 =  x311;
assign c973 =  x242 &  x470 & ~x110 & ~x155 & ~x221 & ~x311 & ~x571 & ~x576 & ~x582 & ~x585 & ~x630 & ~x694;
assign c977 =  x334 & ~x211 & ~x294 & ~x348;
assign c979 =  x331 & ~x250 & ~x534 & ~x574 & ~x580 & ~x585;
assign c981 =  x745;
assign c983 =  x242 &  x331 &  x355 &  x359 &  x383 &  x410 & ~x15 & ~x22 & ~x36 & ~x56 & ~x58 & ~x65 & ~x82 & ~x93 & ~x113 & ~x159 & ~x182 & ~x189 & ~x212 & ~x221 & ~x232 & ~x237 & ~x308 & ~x311 & ~x318 & ~x584 & ~x585 & ~x587 & ~x616 & ~x620 & ~x647 & ~x745 & ~x752;
assign c985 =  x370;
assign c987 =  x466 &  x551 &  x578 & ~x220 & ~x221 & ~x294 & ~x425 & ~x698;
assign c989 = ~x130 & ~x246 & ~x277 & ~x396 & ~x447 & ~x585 & ~x591 & ~x652 & ~x667 & ~x779;
assign c991 =  x119;
assign c993 = ~x353;
assign c995 =  x728;
assign c997 = ~x211 & ~x377 & ~x669 & ~x695;
assign c999 =  x1;
assign c9101 =  x374 &  x403 &  x426 &  x427 &  x443 &  x505 &  x538 & ~x114 & ~x211 & ~x217 & ~x253 & ~x341 & ~x625 & ~x637 & ~x648 & ~x751 & ~x757;
assign c9103 =  x6;
assign c9105 = ~x304 & ~x541 & ~x580;
assign c9107 =  x284;
assign c9109 =  x374 &  x427 &  x552 & ~x278 & ~x612;
assign c9111 =  x305 &  x324 & ~x124 & ~x148 & ~x173 & ~x294 & ~x545;
assign c9113 =  x30;
assign c9115 =  x745;
assign c9117 =  x230;
assign c9119 =  x309;
assign c9121 =  x61;
assign c9123 =  x270 & ~x535 & ~x574 & ~x580 & ~x582 & ~x584 & ~x585 & ~x698 & ~x771;
assign c9125 =  x448;
assign c9127 =  x747;
assign c9129 = ~x274 & ~x301;
assign c9131 =  x149;
assign c9133 =  x760;
assign c9135 = ~x211 & ~x246 & ~x277 & ~x306 & ~x314;
assign c9137 =  x63;
assign c9139 =  x345;
assign c9141 = ~x356;
assign c9143 =  x257;
assign c9145 =  x426 &  x427 & ~x715;
assign c9147 = ~x90 & ~x221 & ~x294 & ~x376 & ~x477 & ~x644 & ~x704;
assign c9149 =  x630 &  x634 & ~x375;
assign c9151 =  x31;
assign c9153 =  x288 &  x314;
assign c9155 =  x30;
assign c9157 = ~x357 & ~x586;
assign c9159 =  x89;
assign c9161 =  x82;
assign c9163 =  x400 &  x402 &  x578;
assign c9165 = ~x403 & ~x523 & ~x580;
assign c9167 =  x363;
assign c9169 =  x92;
assign c9171 = ~x249 & ~x273 & ~x301;
assign c9173 =  x210 & ~x403;
assign c9175 =  x743;
assign c9177 =  x115;
assign c9179 =  x460 &  x470 &  x509 & ~x308 & ~x558 & ~x582 & ~x584 & ~x585 & ~x612;
assign c9181 = ~x489 & ~x580;
assign c9183 =  x481 & ~x249 & ~x263 & ~x278 & ~x294;
assign c9185 =  x368;
assign c9187 =  x12;
assign c9189 =  x729;
assign c9191 = ~x249 & ~x302 & ~x586 & ~x640;
assign c9193 =  x427 &  x487 &  x538 & ~x586 & ~x639;
assign c9195 =  x399 & ~x272;
assign c9197 = ~x489 & ~x642;
assign c9199 =  x119;
assign c9201 = ~x351 & ~x380;
assign c9203 = ~x250 & ~x351 & ~x352 & ~x615;
assign c9205 =  x252;
assign c9207 =  x373 & ~x560 & ~x586 & ~x601 & ~x613;
assign c9209 = ~x408 & ~x478;
assign c9211 =  x118;
assign c9213 =  x110;
assign c9215 = ~x408;
assign c9217 =  x427 &  x520;
assign c9219 = ~x245 & ~x300 & ~x586 & ~x639;
assign c9221 =  x370;
assign c9223 =  x257;
assign c9225 =  x594 & ~x518;
assign c9227 =  x4;
assign c9229 = ~x331 & ~x414;
assign c9231 =  x757;
assign c9233 =  x371;
assign c9235 =  x400 & ~x1 & ~x40 & ~x249 & ~x593;
assign c9237 = ~x435;
assign c9239 =  x439 & ~x294 & ~x535 & ~x571 & ~x572 & ~x575 & ~x580 & ~x581 & ~x593 & ~x656 & ~x670 & ~x695;
assign c9241 =  x228;
assign c9243 =  x291 & ~x388;
assign c9245 =  x286;
assign c9247 =  x398;
assign c9249 =  x346 & ~x250 & ~x312 & ~x668 & ~x734 & ~x736;
assign c9251 =  x346 &  x373 & ~x585;
assign c9253 = ~x278 & ~x320 & ~x552 & ~x561 & ~x635 & ~x638 & ~x769;
assign c9255 =  x400 & ~x160 & ~x187 & ~x273;
assign c9257 =  x498 & ~x408 & ~x606;
assign c9259 =  x215 &  x360 & ~x248 & ~x294;
assign c9261 = ~x249 & ~x323;
assign c9263 =  x11 &  x755;
assign c9265 = ~x333 & ~x525;
assign c9267 = ~x294 & ~x295 & ~x503;
assign c9269 = ~x353;
assign c9271 =  x297 &  x399;
assign c9273 =  x400 & ~x222 & ~x278 & ~x593 & ~x601 & ~x609 & ~x638 & ~x683;
assign c9275 = ~x249 & ~x276 & ~x277 & ~x582 & ~x590;
assign c9277 =  x360 & ~x211 & ~x267 & ~x294 & ~x348 & ~x505 & ~x561;
assign c9279 =  x358 & ~x379;
assign c9281 =  x346 &  x411 & ~x42 & ~x585;
assign c9283 =  x200;
assign c9285 = ~x357;
assign c9287 =  x345;
assign c9289 =  x427 &  x578 &  x605 & ~x183 & ~x194;
assign c9291 =  x363;
assign c9293 =  x368;
assign c9295 =  x145;
assign c9297 =  x93;
assign c9299 =  x773;
assign c9301 =  x271 &  x357 &  x439 & ~x51 & ~x79 & ~x194 & ~x206 & ~x287 & ~x320 & ~x534 & ~x573 & ~x574 & ~x635 & ~x721;
assign c9305 =  x345 &  x398;
assign c9307 =  x182 & ~x461;
assign c9309 =  x243 &  x331 &  x455 & ~x37 & ~x178 & ~x221 & ~x294 & ~x666 & ~x727;
assign c9311 =  x238 & ~x383;
assign c9313 =  x117;
assign c9315 =  x426;
assign c9317 =  x195;
assign c9319 =  x291;
assign c9321 =  x440 & ~x437;
assign c9323 = ~x356 & ~x607;
assign c9325 =  x171;
assign c9327 =  x362 &  x650 & ~x407;
assign c9329 =  x87;
assign c9331 = ~x14 & ~x146 & ~x199 & ~x249 & ~x286 & ~x476 & ~x534 & ~x570 & ~x580 & ~x581 & ~x591 & ~x607 & ~x620 & ~x645 & ~x650 & ~x696;
assign c9333 =  x281;
assign c9335 = ~x354;
assign c9337 =  x341;
assign c9339 =  x392 & ~x492;
assign c9341 = ~x494 & ~x573;
assign c9343 =  x773;
assign c9345 =  x344 &  x398;
assign c9347 =  x62;
assign c9349 =  x190 & ~x302 & ~x432;
assign c9351 =  x7;
assign c9353 =  x296 &  x427 &  x550 &  x556 & ~x158 & ~x278 & ~x290 & ~x422 & ~x589 & ~x620 & ~x667 & ~x694 & ~x746;
assign c9355 =  x745;
assign c9357 =  x242 & ~x304 & ~x378;
assign c9359 =  x281;
assign c9361 =  x400 & ~x301;
assign c9363 =  x746;
assign c9365 =  x233;
assign c9367 =  x92;
assign c9369 =  x400 & ~x59 & ~x163 & ~x250 & ~x263 & ~x273;
assign c9371 =  x154;
assign c9373 = ~x523;
assign c9375 =  x28;
assign c9377 =  x339;
assign c9379 =  x341;
assign c9381 =  x371;
assign c9383 =  x623 & ~x379 & ~x404;
assign c9385 =  x318 & ~x358;
assign c9387 =  x285;
assign c9389 =  x86;
assign c9391 =  x66;
assign c9393 = ~x414;
assign c9395 =  x600 &  x623 &  x630 &  x634 & ~x164 & ~x263 & ~x751;
assign c9397 =  x783;
assign c9399 =  x27;
assign c9401 =  x285;
assign c9403 =  x399 &  x476;
assign c9405 =  x400 & ~x300;
assign c9407 =  x89;
assign c9409 = ~x466;
assign c9411 =  x425 & ~x500;
assign c9413 =  x92;
assign c9415 = ~x408;
assign c9417 =  x744;
assign c9419 =  x426 & ~x378;
assign c9421 =  x90;
assign c9423 =  x761;
assign c9425 = ~x299 & ~x612;
assign c9427 =  x230;
assign c9429 = ~x379;
assign c9431 = ~x305 & ~x469;
assign c9433 =  x745;
assign c9435 = ~x356;
assign c9437 =  x400 &  x455 & ~x246 & ~x608;
assign c9439 =  x308;
assign c9441 =  x256;
assign c9443 =  x203;
assign c9445 =  x208;
assign c9447 = ~x351 & ~x352;
assign c9449 = ~x222 & ~x525 & ~x534 & ~x580;
assign c9451 =  x427 &  x605 & ~x644 & ~x691;
assign c9453 = ~x18 & ~x489 & ~x580;
assign c9455 =  x455 &  x460 &  x472 &  x508 & ~x249 & ~x593 & ~x778;
assign c9457 =  x191;
assign c9459 =  x141;
assign c9461 =  x756;
assign c9465 =  x556 & ~x490 & ~x694;
assign c9467 =  x64;
assign c9469 =  x91;
assign c9471 = ~x519 & ~x574;
assign c9473 = ~x435 & ~x505 & ~x608;
assign c9475 =  x443 &  x631 &  x633 & ~x221 & ~x712;
assign c9477 = ~x221 & ~x366 & ~x523 & ~x553 & ~x583;
assign c9479 =  x116;
assign c9481 =  x142;
assign c9483 = ~x437;
assign c9485 = ~x277 & ~x305 & ~x553;
assign c9487 =  x215 &  x541 &  x600 &  x605 &  x631 &  x634 & ~x116 & ~x294;
assign c9489 =  x344 &  x398;
assign c9491 =  x182 & ~x382;
assign c9493 = ~x523 & ~x543 & ~x552;
assign c9495 =  x399 & ~x74 & ~x585;
assign c9497 =  x400 & ~x273;
assign c9499 =  x85;

endmodule