module tm( x0,x1,x2,x3,x4,x5,x6,x7,x8,x9,x10,x11,x12,x13,x14,x15,x16,x17,x18,x19,x20,x21,x22,x23,x24,x25,x26,x27,x28,x29,x30,x31,x32,x33,x34,x35,x36,x37,x38,x39,x40,x41,x42,x43,x44,x45,x46,x47,x48,x49,x50,x51,x52,x53,x54,x55,x56,x57,x58,x59,x60,x61,x62,x63,x64,x65,x66,x67,x68,x69,x70,x71,x72,x73,x74,x75,x76,x77,x78,x79,x80,x81,x82,x83,x84,x85,x86,x87,x88,x89,x90,x91,x92,x93,x94,x95,x96,x97,x98,x99,x100,x101,x102,x103,x104,x105,x106,x107,x108,x109,x110,x111,x112,x113,x114,x115,x116,x117,x118,x119,x120,x121,x122,x123,x124,x125,x126,x127,x128,x129,x130,x131,x132,x133,x134,x135,x136,x137,x138,x139,x140,x141,x142,x143,x144,x145,x146,x147,x148,x149,x150,x151,x152,x153,x154,x155,x156,x157,x158,x159,x160,x161,x162,x163,x164,x165,x166,x167,x168,x169,x170,x171,x172,x173,x174,x175,x176,x177,x178,x179,x180,x181,x182,x183,x184,x185,x186,x187,x188,x189,x190,x191,x192,x193,x194,x195,x196,x197,x198,x199,x200,x201,x202,x203,x204,x205,x206,x207,x208,x209,x210,x211,x212,x213,x214,x215,x216,x217,x218,x219,x220,x221,x222,x223,x224,x225,x226,x227,x228,x229,x230,x231,x232,x233,x234,x235,x236,x237,x238,x239,x240,x241,x242,x243,x244,x245,x246,x247,x248,x249,x250,x251,x252,x253,x254,x255,x256,x257,x258,x259,x260,x261,x262,x263,x264,x265,x266,x267,x268,x269,x270,x271,x272,x273,x274,x275,x276,x277,x278,x279,x280,x281,x282,x283,x284,x285,x286,x287,x288,x289,x290,x291,x292,x293,x294,x295,x296,x297,x298,x299,x300,x301,x302,x303,x304,x305,x306,x307,x308,x309,x310,x311,x312,x313,x314,x315,x316,x317,x318,x319,x320,x321,x322,x323,x324,x325,x326,x327,x328,x329,x330,x331,x332,x333,x334,x335,x336,x337,x338,x339,x340,x341,x342,x343,x344,x345,x346,x347,x348,x349,x350,x351,x352,x353,x354,x355,x356,x357,x358,x359,x360,x361,x362,x363,x364,x365,x366,x367,x368,x369,x370,x371,x372,x373,x374,x375,x376,x377,x378,x379,x380,x381,x382,x383,x384,x385,x386,x387,x388,x389,x390,x391,x392,x393,x394,x395,x396,x397,x398,x399,x400,x401,x402,x403,x404,x405,x406,x407,x408,x409,x410,x411,x412,x413,x414,x415,x416,x417,x418,x419,x420,x421,x422,x423,x424,x425,x426,x427,x428,x429,x430,x431,x432,x433,x434,x435,x436,x437,x438,x439,x440,x441,x442,x443,x444,x445,x446,x447,x448,x449,x450,x451,x452,x453,x454,x455,x456,x457,x458,x459,x460,x461,x462,x463,x464,x465,x466,x467,x468,x469,x470,x471,x472,x473,x474,x475,x476,x477,x478,x479,x480,x481,x482,x483,x484,x485,x486,x487,x488,x489,x490,x491,x492,x493,x494,x495,x496,x497,x498,x499,x500,x501,x502,x503,x504,x505,x506,x507,x508,x509,x510,x511,x512,x513,x514,x515,x516,x517,x518,x519,x520,x521,x522,x523,x524,x525,x526,x527,x528,x529,x530,x531,x532,x533,x534,x535,x536,x537,x538,x539,x540,x541,x542,x543,x544,x545,x546,x547,x548,x549,x550,x551,x552,x553,x554,x555,x556,x557,x558,x559,x560,x561,x562,x563,x564,x565,x566,x567,x568,x569,x570,x571,x572,x573,x574,x575,x576,x577,x578,x579,x580,x581,x582,x583,x584,x585,x586,x587,x588,x589,x590,x591,x592,x593,x594,x595,x596,x597,x598,x599,x600,x601,x602,x603,x604,x605,x606,x607,x608,x609,x610,x611,x612,x613,x614,x615,x616,x617,x618,x619,x620,x621,x622,x623,x624,x625,x626,x627,x628,x629,x630,x631,x632,x633,x634,x635,x636,x637,x638,x639,x640,x641,x642,x643,x644,x645,x646,x647,x648,x649,x650,x651,x652,x653,x654,x655,x656,x657,x658,x659,x660,x661,x662,x663,x664,x665,x666,x667,x668,x669,x670,x671,x672,x673,x674,x675,x676,x677,x678,x679,x680,x681,x682,x683,x684,x685,x686,x687,x688,x689,x690,x691,x692,x693,x694,x695,x696,x697,x698,x699,x700,x701,x702,x703,x704,x705,x706,x707,x708,x709,x710,x711,x712,x713,x714,x715,x716,x717,x718,x719,x720,x721,x722,x723,x724,x725,x726,x727,x728,x729,x730,x731,x732,x733,x734,x735,x736,x737,x738,x739,x740,x741,x742,x743,x744,x745,x746,x747,x748,x749,x750,x751,x752,x753,x754,x755,x756,x757,x758,x759,x760,x761,x762,x763,x764,x765,x766,x767,x768,x769,x770,x771,x772,x773,x774,x775,x776,x777,x778,x779,x780,x781,x782,x783,c07,c615,c0273,c464,c011,c126,c439,c1125,c3286,c7146,c4276,c528,c5230,c1289,c9161,c7145,c359,c4144,c029,c680,c0219,c880,c6206,c925,c0150,c546,c9225,c0201,c0191,c5260,c6251,c4235,c967,c9141,c084,c1201,c7243,c8127,c587,c2283,c3210,c530,c934,c0199,c5160,c6105,c458,c5217,c4292,c21,c599,c6264,c736,c8188,c322,c3200,c9126,c7228,c6110,c6228,c388,c0181,c547,c492,c592,c295,c190,c6139,c88,c0141,c4125,c664,c9198,c5184,c090,c1133,c2289,c175,c4238,c1176,c4209,c0184,c5214,c525,c5127,c2236,c749,c8155,c1150,c0105,c6291,c974,c9142,c7209,c51,c9154,c3288,c5131,c4219,c0156,c214,c4229,c6278,c8170,c924,c0237,c366,c9183,c168,c9283,c9166,c964,c118,c1259,c6242,c293,c5235,c7211,c2190,c2233,c3148,c398,c1298,c259,c4180,c0161,c2250,c68,c7264,c7294,c9127,c1299,c1143,c3110,c9262,c0122,c25,c298,c328,c6118,c376,c864,c8112,c762,c6142,c0218,c245,c6103,c9185,c6231,c5225,c1117,c6114,c1197,c8251,c048,c6158,c5292,c1152,c2256,c2155,c8145,c7289,c710,c8246,c4163,c5118,c24,c7292,c088,c821,c223,c3293,c930,c396,c0265,c3218,c6208,c7116,c5255,c095,c7100,c3155,c621,c078,c249,c297,c5159,c1239,c4227,c2151,c5254,c3146,c537,c6165,c129,c4246,c665,c2213,c7299,c1100,c8288,c839,c580,c2220,c09,c757,c779,c1225,c8161,c0148,c211,c716,c6101,c6214,c798,c4241,c354,c8179,c9232,c65,c423,c4271,c7213,c4256,c631,c972,c844,c4143,c0228,c1128,c036,c0137,c794,c0206,c2242,c9205,c9137,c945,c53,c1156,c6104,c777,c0252,c367,c8254,c5170,c7274,c7262,c047,c0294,c7219,c6108,c2128,c6273,c987,c8243,c9231,c9218,c092,c4107,c0171,c043,c6217,c0276,c4199,c4228,c541,c8187,c393,c9147,c720,c1105,c1144,c427,c0144,c7120,c0288,c5247,c954,c1258,c9189,c0277,c69,c8174,c2116,c5136,c759,c614,c3240,c1180,c8122,c9148,c9259,c784,c4130,c2115,c6265,c2176,c2251,c763,c589,c699,c6136,c151,c8255,c5222,c4223,c596,c4245,c032,c3165,c5155,c6298,c7197,c848,c8196,c0165,c473,c566,c079,c6286,c782,c7202,c9214,c2211,c0239,c521,c221,c0153,c1267,c361,c075,c2154,c456,c241,c2244,c3291,c7154,c9263,c670,c2276,c2189,c1183,c3287,c072,c2225,c3184,c0207,c894,c9134,c9203,c8194,c8147,c498,c7251,c4178,c7183,c39,c3132,c1164,c3267,c9191,c116,c852,c742,c7180,c6195,c0159,c3254,c3177,c9224,c0270,c4160,c2142,c6156,c7204,c1122,c4288,c4265,c60,c7257,c1139,c7290,c1252,c522,c5271,c5224,c061,c115,c9292,c8191,c970,c9107,c9210,c419,c6146,c1135,c3233,c331,c831,c2241,c6187,c7248,c941,c063,c4259,c1238,c9213,c554,c918,c338,c861,c885,c2170,c1296,c1279,c2238,c2119,c3131,c3181,c5106,c575,c645,c7270,c4150,c985,c2185,c940,c616,c889,c545,c313,c0284,c5223,c5137,c8148,c320,c2265,c3180,c94,c937,c3142,c955,c0128,c8171,c0286,c7254,c451,c428,c1162,c5168,c7293,c3187,c185,c3284,c1169,c1234,c7143,c2194,c4218,c881,c3178,c7200,c40,c5203,c3271,c4298,c0167,c3169,c20,c590,c0204,c6258,c485,c7286,c1229,c025,c0197,c89,c8214,c6182,c6111,c6295,c30,c6266,c866,c6154,c261,c5280,c34,c466,c4106,c4149,c9228,c3183,c6173,c8181,c3281,c5252,c5122,c1281,c986,c7265,c890,c437,c12,c4112,c5185,c4258,c3292,c8263,c1188,c285,c379,c5130,c363,c454,c8208,c2161,c4172,c7110,c8257,c4250,c734,c049,c114,c0126,c7173,c6184,c7208,c5150,c6122,c1286,c4101,c951,c340,c181,c0215,c383,c141,c2124,c8225,c4239,c9230,c9242,c8294,c2150,c1126,c3258,c3265,c1295,c862,c4127,c1241,c778,c79,c6121,c018,c1193,c8121,c9162,c5153,c6289,c8242,c2181,c555,c582,c0187,c033,c1142,c7194,c2280,c77,c3108,c5147,c4167,c613,c915,c7214,c1290,c2262,c0119,c4277,c41,c9180,c7184,c7178,c7205,c069,c0229,c7157,c944,c2231,c9200,c874,c694,c7217,c2235,c8137,c9273,c729,c1190,c657,c1246,c5149,c6220,c543,c4214,c6175,c053,c3100,c7263,c836,c9254,c349,c8207,c6120,c337,c2222,c6180,c4204,c2199,c6210,c5250,c424,c042,c0248,c9247,c659,c7285,c264,c4187,c3138,c2273,c756,c766,c8205,c6283,c8266,c6163,c5205,c7210,c7170,c2297,c5105,c1219,c3243,c3127,c0236,c0113,c390,c9265,c3111,c4102,c2261,c476,c8227,c4152,c13,c6194,c4253,c5204,c642,c80,c461,c1111,c0140,c6128,c7241,c3241,c436,c8200,c172,c5236,c2180,c5288,c086,c284,c9105,c5296,c2131,c5278,c5287,c198,c0152,c1194,c1157,c6135,c5277,c2164,c558,c5213,c4222,c2138,c8163,c368,c369,c4110,c5157,c164,c5191,c4282,c443,c7164,c0182,c4224,c45,c4262,c0189,c4197,c19,c0102,c9184,c4115,c046,c0295,c627,c0160,c1216,c3221,c2224,c0151,c345,c4161,c3204,c563,c137,c226,c386,c690,c7207,c0287,c022,c5265,c8264,c7108,c6124,c3276,c9176,c2166,c3172,c5110,c045,c8219,c872,c0209,c1287,c0269,c3112,c4153,c5154,c6157,c4158,c6189,c7152,c7275,c1209,c9279,c8151,c938,c7297,c0106,c0123,c4168,c75,c362,c9167,c1160,c271,c559,c1231,c332,c2201,c9102,c655,c0101,c2253,c3153,c462,c7150,c3158,c935,c9174,c2218,c980,c8277,c8283,c2100,c6152,c429,c725,c6280,c72,c373,c10,c2249,c7189,c576,c2109,c6272,c247,c786,c7199,c816,c4296,c9135,c3299,c5234,c71,c968,c1269,c3122,c333,c9160,c7112,c629,c460,c572,c3277,c6239,c021,c0242,c3117,c4183,c1102,c8282,c1282,c425,c5263,c9112,c9156,c060,c136,c5100,c3248,c1154,c0147,c239,c1243,c6224,c3215,c845,c1173,c1113,c9115,c272,c2205,c5144,c1233,c270,c023,c6252,c83,c3168,c8185,c0155,c5228,c963,c319,c2139,c2247,c3216,c828,c9129,c9229,c1149,c134,c971,c188,c693,c58,c5108,c0142,c531,c5114,c721,c299,c7249,c49,c5129,c3198,c553,c5192,c232,c5197,c689,c7124,c99,c825,c1274,c4299,c6144,c0283,c752,c2195,c5146,c4138,c6192,c9204,c0175,c252,c040,c2208,c4192,c978,c9208,c3104,c3189,c165,c4182,c1112,c494,c8107,c9149,c5196,c167,c9216,c3217,c579,c1163,c213,c4131,c4135,c4207,c9234,c0115,c8285,c8235,c7172,c529,c121,c52,c1277,c347,c1236,c1202,c2254,c5257,c62,c098,c1250,c364,c7196,c1266,c3219,c184,c5282,c158,c6260,c931,c6193,c0253,c8197,c6293,c6150,c5261,c6190,c711,c5152,c1251,c074,c2165,c636,c6130,c569,c5209,c3234,c6100,c8212,c714,c4275,c3235,c8109,c9146,c5276,c7246,c316,c552,c495,c0235,c7291,c43,c5161,c571,c943,c3114,c3227,c2144,c076,c7279,c8111,c776,c2177,c5158,c671,c9240,c268,c6243,c5174,c5111,c859,c649,c887,c556,c5125,c235,c9159,c1212,c5264,c2196,c1245,c540,c33,c7118,c9296,c6166,c6170,c911,c0212,c8290,c2270,c161,c1124,c1232,c8274,c0136,c6285,c1170,c946,c526,c515,c2232,c5182,c5258,c399,c0198,c927,c479,c5166,c995,c942,c1148,c382,c2130,c4129,c9291,c1179,c9243,c4155,c0247,c1181,c174,c3296,c4252,c883,c92,c421,c1222,c446,c5132,c5206,c7162,c1214,c997,c171,c891,c8154,c0200,c920,c9118,c3209,c29,c2210,c1228,c0293,c489,c9139,c3255,c1254,c1177,c0272,c0281,c5269,c7121,c3174,c493,c750,c0192,c374,c577,c728,c7192,c6181,c8136,c0268,c2263,c8128,c6253,c5218,c981,c854,c7206,c414,c2198,c879,c7131,c2287,c4260,c1136,c7273,c868,c263,c6262,c027,c877,c1208,c1297,c342,c0254,c78,c135,c6137,c7187,c068,c644,c375,c667,c155,c8206,c9245,c1165,c142,c9257,c9144,c2160,c676,c066,c166,c336,c656,c739,c6117,c837,c6125,c2126,c2169,c5259,c583,c992,c775,c989,c5295,c70,c267,c27,c7101,c1168,c9297,c5299,c9235,c0221,c850,c2239,c3182,c1172,c8226,c6141,c4215,c5198,c0114,c0261,c6219,c138,c4170,c923,c523,c9271,c0203,c4272,c5109,c4132,c6234,c3214,c3253,c2277,c1270,c5220,c9207,c5102,c824,c8279,c1182,c3226,c5186,c684,c7171,c8265,c4251,c3145,c5128,c6249,c581,c9206,c7115,c0143,c9188,c3159,c256,c3263,c6126,c8166,c8271,c2125,c8275,c3270,c949,c1108,c8102,c910,c377,c052,c019,c3124,c9187,c397,c3207,c260,c9241,c8231,c378,c7168,c628,c119,c6237,c6199,c2135,c5162,c224,c6276,c6160,c197,c6267,c5212,c246,c497,c2132,c7161,c1213,c04,c7216,c6102,c4148,c95,c2117,c150,c8261,c6221,c8281,c9275,c5298,c669,c519,c274,c3290,c772,c4213,c5178,c7158,c510,c548,c430,c744,c0176,c4266,c3107,c2108,c457,c5231,c132,c832,c4123,c7151,c1263,c884,c3102,c8248,c2203,c028,c1175,c6223,c9299,c4166,c097,c567,c5294,c8220,c3154,c3197,c4165,c3245,c6248,c4226,c496,c1151,c0214,c966,c947,c0249,c818,c255,c7255,c3249,c2258,c830,c8278,c4139,c7137,c189,c4243,c594,c8291,c9249,c8286,c1280,c2294,c1247,c070,c3105,c7142,c4286,c624,c1226,c4174,c0230,c453,c654,c7256,c0132,c4255,c64,c0243,c1207,c6284,c6145,c9181,c5242,c8139,c3133,c686,c0193,c4237,c9136,c2186,c3128,c348,c849,c0133,c3190,c03,c465,c838,c6116,c156,c2200,c6241,c0205,c8125,c0223,c7156,c8141,c591,c1184,c2197,c916,c2259,c1271,c2192,c612,c7231,c2293,c730,c6168,c743,c8240,c9197,c0100,c4208,c2223,c0178,c8153,c0233,c8215,c4140,c3242,c6205,c5177,c7138,c6236,c3162,c5270,c6244,c6235,c6162,c486,c4133,c038,c7165,c4105,c1118,c1278,c5101,c8198,c9100,c8272,c448,c754,c467,c765,c131,c4291,c4195,c5244,c275,c244,c394,c2228,c2120,c4225,c564,c797,c6169,c8115,c8298,c5117,c2272,c4154,c5104,c9172,c7227,c851,c442,c2105,c3171,c8201,c0202,c9268,c6202,c145,c8292,c2129,c2163,c148,c9186,c0255,c3261,c3297,c1129,c0241,c0138,c5240,c0121,c9132,c3119,c0264,c2122,c2102,c6246,c9199,c077,c1155,c8195,c227,c6133,c3205,c2148,c8114,c7149,c218,c0274,c962,c9277,c2110,c0224,c2147,c1167,c7239,c9195,c9151,c4128,c248,c2295,c731,c7177,c5139,c9222,c0190,c633,c3199,c593,c912,c584,c1288,c4206,c288,c4297,c1198,c688,c173,c610,c8183,c2217,c993,c030,c8140,c194,c157,c1273,c640,c250,c9106,c8184,c5237,c1200,c4295,c86,c8268,c6177,c8221,c2106,c7193,c8160,c4114,c1265,c2214,c123,c5283,c8239,c2269,c9290,c16,c2267,c991,c7222,c5273,c3134,c799,c450,c4263,c7221,c2121,c751,c0134,c468,c2207,c3222,c7280,c8108,c0110,c3120,c7284,c1101,c0222,c1147,c0154,c93,c3201,c3272,c035,c472,c6127,c9261,c5135,c999,c8180,c820,c9294,c4171,c449,c389,c433,c0280,c1210,c483,c8204,c133,c191,c9212,c3274,c1211,c764,c1255,c7105,c220,c7136,c712,c792,c7266,c588,c3232,c733,c262,c4269,c8284,c3166,c4177,c2145,c8297,c010,c5285,c741,c4198,c0120,c094,c7195,c8172,c8164,c544,c746,c7133,c1221,c410,c0238,c176,c6176,c2298,c417,c1192,c3125,c678,c0245,c3163,c7117,c626,c785,c55,c888,c4254,c5175,c44,c1132,c9163,c9202,c1110,c562,c9168,c7122,c3140,c4279,c7181,c512,c7160,c330,c740,c7190,c899,c8262,c3152,c956,c7128,c3103,c0257,c422,c5227,c17,c9215,c1145,c1186,c323,c3206,c755,c698,c9253,c3231,c9211,c5290,c3279,c3275,c6149,c939,c243,c2174,c895,c9256,c7126,c933,c6174,c3160,c280,c994,c0263,c3257,c35,c8295,c26,c857,c998,c957,c0117,c961,c055,c5169,c5165,c344,c487,c392,c9280,c565,c6287,c758,c3208,c8133,c7258,c7191,c8256,c97,c9124,c117,c1230,c771,c8247,c660,c4261,c61,c3252,c153,c3236,c842,c8260,c7144,c713,c9175,c871,c0104,c7276,c7169,c619,c2282,c1185,c4120,c5208,c9272,c4210,c1260,c9286,c6153,c9196,c057,c3239,c535,c7212,c6203,c2246,c2193,c4124,c499,c9246,c1106,c9282,c4116,c4126,c9133,c8158,c237,c1141,c357,c4188,c1272,c1256,c3295,c183,c4249,c8103,c9178,c9113,c276,c455,c865,c0194,c7236,c814,c5239,c435,c6155,c286,c0282,c7139,c0211,c0289,c4242,c1161,c6263,c873,c9173,c7159,c3278,c732,c238,c8218,c9143,c416,c9258,c952,c2103,c4264,c7111,c3135,c863,c3237,c4184,c02,c215,c719,c0196,c5291,c1293,c7282,c913,c0244,c8237,c7252,c8287,c356,c1159,c3144,c973,c637,c897,c5246,c3246,c516,c8168,c723,c1285,c6288,c7153,c5142,c536,c0116,c56,c1220,c8224,c8126,c130,c6171,c5219,c598,c9217,c8202,c2187,c2127,c8252,c858,c0226,c2292,c4185,c159,c685,c326,c1114,c796,c7129,c892,c441,c0179,c4151,c265,c32,c738,c2162,c1174,c514,c6274,c3256,c6185,c8167,c234,c381,c8211,c371,c7188,c622,c635,c781,c0125,c9121,c4270,c4202,c2101,c9190,c5262,c9120,c9103,c2137,c46,c4111,c2264,c310,c5103,c5266,c0118,c2234,c4211,c557,c0124,c186,c666,c5124,c9264,c6164,c0260,c085,c160,c216,c5167,c4176,c5272,c8117,c7287,c2229,c7186,c0285,c788,c8250,c2281,c6196,c6292,c8105,c691,c1275,c3116,c149,c8216,c87,c3141,c432,c745,c6212,c661,c2290,c7220,c812,c856,c0173,c020,c5215,c8222,c4189,c081,c06,c351,c0290,c8192,c5183,c5274,c7245,c3170,c7223,c7296,c7247,c767,c8119,c289,c2167,c2156,c469,c822,c7277,c199,c380,c7167,c2158,c8165,c73,c4104,c641,c127,c0166,c840,c3244,c922,c1284,c7233,c5210,c9164,c0251,c054,c463,c5195,c9239,c4289,c8152,c1242,c6119,c5194,c8249,c8106,c6159,c9150,c632,c4201,c4196,c1127,c0213,c3143,c8176,c9295,c5253,c1204,c672,c236,c768,c5243,c484,c7203,c253,c9248,c726,c3230,c339,c652,c977,c0158,c724,c6218,c6255,c7135,c718,c254,c6179,c982,c841,c279,c1166,c8129,c026,c6222,c258,c5138,c2248,c9108,c3136,c242,c7259,c1119,c192,c4147,c780,c1109,c3106,c2279,c4273,c0162,c6147,c212,c5233,c3192,c1146,c2202,c9220,c481,c7106,c48,c7132,c2221,c2175,c6186,c90,c9170,c0135,c3101,c5141,c787,c080,c3280,c789,c7237,c4181,c74,c290,c9153,c8182,c140,c677,c31,c2299,c9193,c5216,c6167,c28,c5163,c9110,c9233,c0149,c452,c4136,c5279,c42,c8120,c067,c674,c0298,c8189,c3251,c7261,c976,c959,c4173,c2172,c4169,c6188,c3188,c0112,c2268,c4146,c96,c6238,c0109,c196,c1104,c819,c7260,c9219,c9223,c7147,c122,c511,c039,c761,c7179,c5115,c4267,c5248,c1235,c287,c3211,c5133,c2204,c8134,c542,c152,c7114,c3212,c8132,c6134,c7107,c513,c324,c1121,c8169,c210,c843,c5201,c936,c099,c2111,c00,c8203,c869,c3285,c2266,c57,c8241,c847,c8190,c1116,c9119,c9130,c550,c737,c1237,c3294,c5176,c2123,c2171,c870,c083,c4159,c2245,c459,c520,c4247,c7238,c0297,c1107,c2140,c896,c9194,c893,c7103,c8213,c3191,c1203,c0163,c8130,c2278,c9227,c0256,c6172,c8131,c735,c418,c3179,c412,c7295,c91,c63,c3196,c5200,c2209,c6198,c8293,c0231,c7229,c9201,c8162,c8149,c538,c620,c434,c6257,c0291,c4175,c8236,c5107,c1120,c7104,c8157,c7141,c1171,c1205,c05,c517,c791,c2257,c111,c8230,c0258,c929,c7253,c2134,c7250,c315,c0111,c2112,c647,c182,c1195,c6138,c447,c426,c9101,c041,c790,c8273,c3161,c8245,c663,c1294,c0131,c1283,c0266,c231,c5256,c5211,c1292,c0172,c4244,c7244,c6240,c9104,c5249,c1158,c662,c1264,c343,c650,c4230,c1268,c722,c3202,c8289,c6131,c5143,c988,c8280,c325,c3121,c5145,c311,c059,c990,c0208,c9260,c411,c618,c835,c6227,c277,c0278,c431,c6250,c9288,c0127,c4293,c179,c9171,c717,c813,c478,c490,c9278,c3109,c8156,c471,c3260,c3229,c3269,c673,c139,c4232,c8110,c016,c225,c8100,c6112,c327,c630,c8270,c6229,c534,c9276,c9109,c124,c2143,c8143,c9122,c2118,c524,c0145,c170,c195,c296,c4240,c3247,c6183,c4278,c7234,c7182,c2288,c6245,c8116,c0195,c1131,c193,c294,c3164,c1189,c876,c4109,c482,c8259,c6294,c7269,c5293,c37,c5297,c9274,c770,c2104,c475,c9289,c037,c9298,c2260,c8296,c2291,c3225,c4274,c2133,c7130,c950,c056,c8135,c0210,c867,c9145,c062,c01,c15,c2159,c9192,c66,c6230,c9165,c7123,c358,c3176,c4281,c7198,c8113,c0267,c1291,c3273,c6201,c9209,c783,c5164,c8217,c7224,c917,c8228,c7134,c3126,c586,c846,c9226,c826,c146,c14,c8144,c334,c2240,c087,c0108,c1240,c853,c4284,c969,c882,c318,c4156,c3139,c162,c5173,c2191,c5251,c7174,c9244,c1123,c8146,c415,c4231,c715,c7102,c5187,c1244,c643,c1178,c6211,c6148,c823,c4141,c1187,c539,c7215,c091,c0168,c4119,c570,c8199,c2152,c064,c125,c229,c4103,c065,c4285,c6297,c341,c960,c9182,c6270,c3250,c3259,c0180,c793,c7235,c8118,c384,c4234,c928,c0225,c67,c6161,c031,c7185,c8258,c350,c251,c76,c4194,c0107,c0220,c8244,c050,c0259,c4121,c2113,c291,c753,c3118,c6113,c8209,c0129,c8178,c6233,c4142,c1217,c6226,c3223,c5112,c7288,c658,c6178,c7230,c6268,c773,c9236,c6282,c59,c6197,c3298,c4191,c1261,c1115,c5171,c1257,c7148,c6254,c5151,c2296,c488,c257,c9138,c089,c8233,c269,c638,c8138,c0186,c3113,c9157,c7125,c4122,c7175,c230,c829,c4203,c0130,c4117,c6269,c0246,c5232,c491,c8223,c8124,c774,c266,c0157,c2230,c321,c7272,c2243,c898,c0216,c653,c98,c012,c0227,c2237,c9140,c0234,c143,c1199,c3264,c5238,c834,c6191,c352,c1130,c1223,c440,c7113,c815,c948,c0240,c5202,c4236,c8269,c096,c6225,c760,c4280,c9155,c533,c470,c3185,c7232,c3130,c574,c875,c6200,c480,c282,c2285,c391,c1206,c5121,c953,c921,c4268,c8276,c878,c697,c7218,c18,c6299,c438,c2153,c886,c2286,c395,c5120,c5134,c2178,c113,c5229,c178,c4290,c0139,c617,c560,c2274,c329,c47,c6107,c7226,c692,c0164,c4100,c7267,c1103,c9284,c8175,c6109,c682,c233,c8232,c9293,c312,c3123,c5199,c9158,c110,c2146,c8238,c5140,c4113,c2275,c860,c0262,c3151,c273,c8186,c695,c8210,c9252,c926,c177,c6281,c5245,c128,c0185,c595,c6247,c6275,c4179,c855,c8101,c6290,c017,c3147,c2284,c5119,c687,c84,c5189,c9250,c2184,c9285,c4205,c9152,c50,c4190,c9125,c3156,c013,c3150,c4233,c1276,c6207,c169,c549,c2212,c578,c0169,c573,c7281,c7283,c2227,c6123,c283,c360,c372,c82,c093,c180,c984,c5281,c2141,c7119,c965,c4217,c979,c387,c228,c675,c4145,c5190,c0217,c3289,c727,c6216,c1253,c474,c4193,c38,c0232,c217,c679,c6215,c2226,c9111,c2255,c748,c625,c747,c5172,c827,c8193,c278,c9267,c919,c3224,c681,c9179,c551,c163,c082,c3186,c073,c051,c696,c9266,c833,c5180,c6132,c112,c3262,c5284,c413,c034,c292,c975,c4212,c5193,c2183,c444,c668,c2271,c7155,c9237,c6143,c0275,c5226,c4220,c2173,c7163,c2114,c4164,c3195,c4283,c0174,c335,c6151,c518,c8234,c648,c4108,c9117,c651,c85,c9116,c9255,c0188,c3228,c4294,c9131,c1196,c2107,c0292,c3203,c4216,c014,c5221,c6256,c9269,c9251,c11,c7176,c8267,c355,c2157,c071,c3283,c5188,c5275,c9270,c4137,c2216,c6271,c3220,c385,c6209,c0250,c769,c7140,c983,c9169,c314,c222,c4221,c36,c6296,c9177,c1153,c187,c8159,c958,c6204,c1224,c4157,c147,c795,c54,c6140,c561,c5207,c4200,c634,c024,c8123,c1134,c044,c6279,c1227,c6106,c532,c7278,c08,c810,c0170,c3137,c527,c9221,c4287,c1248,c6277,c8177,c346,c3173,c7240,c477,c23,c353,c9238,c1137,c0183,c3115,c445,c015,c9128,c3282,c5289,c7166,c8253,c370,c8142,c5113,c2252,c5126,c9287,c4257,c6129,c22,c5116,c3175,c5268,c420,c5241,c6115,c5286,c2206,c6261,c0271,c0146,c7298,c9281,c7201,c1191,c5179,c1215,c2182,c6232,c8104,c683,c9114,c365,c0103,c0177,c3194,c4248,c3149,c639,c2168,c144,c811,c240,c4134,c2149,c7268,c996,c7225,c585,c1138,c058,c8173,c7242,c0296,c7127,c0299,c3157,c5267,c6213,c3266,c8150,c1262,c4162,c568,c817,c6259,c8229,c597,c5156,c932,c7109,c3238,c154,c5148,c5181,c3167,c1218,c2215,c3193,c0279,c2188,c623,c611,c8299,c2136,c914,c317,c3213,c3129,c1140,c2179,c4118,c3268,c4186,c646,c1249,c219,c120,c9123,c2219,c5123,c7271,c281,c81 );

input x0;
input x1;
input x2;
input x3;
input x4;
input x5;
input x6;
input x7;
input x8;
input x9;
input x10;
input x11;
input x12;
input x13;
input x14;
input x15;
input x16;
input x17;
input x18;
input x19;
input x20;
input x21;
input x22;
input x23;
input x24;
input x25;
input x26;
input x27;
input x28;
input x29;
input x30;
input x31;
input x32;
input x33;
input x34;
input x35;
input x36;
input x37;
input x38;
input x39;
input x40;
input x41;
input x42;
input x43;
input x44;
input x45;
input x46;
input x47;
input x48;
input x49;
input x50;
input x51;
input x52;
input x53;
input x54;
input x55;
input x56;
input x57;
input x58;
input x59;
input x60;
input x61;
input x62;
input x63;
input x64;
input x65;
input x66;
input x67;
input x68;
input x69;
input x70;
input x71;
input x72;
input x73;
input x74;
input x75;
input x76;
input x77;
input x78;
input x79;
input x80;
input x81;
input x82;
input x83;
input x84;
input x85;
input x86;
input x87;
input x88;
input x89;
input x90;
input x91;
input x92;
input x93;
input x94;
input x95;
input x96;
input x97;
input x98;
input x99;
input x100;
input x101;
input x102;
input x103;
input x104;
input x105;
input x106;
input x107;
input x108;
input x109;
input x110;
input x111;
input x112;
input x113;
input x114;
input x115;
input x116;
input x117;
input x118;
input x119;
input x120;
input x121;
input x122;
input x123;
input x124;
input x125;
input x126;
input x127;
input x128;
input x129;
input x130;
input x131;
input x132;
input x133;
input x134;
input x135;
input x136;
input x137;
input x138;
input x139;
input x140;
input x141;
input x142;
input x143;
input x144;
input x145;
input x146;
input x147;
input x148;
input x149;
input x150;
input x151;
input x152;
input x153;
input x154;
input x155;
input x156;
input x157;
input x158;
input x159;
input x160;
input x161;
input x162;
input x163;
input x164;
input x165;
input x166;
input x167;
input x168;
input x169;
input x170;
input x171;
input x172;
input x173;
input x174;
input x175;
input x176;
input x177;
input x178;
input x179;
input x180;
input x181;
input x182;
input x183;
input x184;
input x185;
input x186;
input x187;
input x188;
input x189;
input x190;
input x191;
input x192;
input x193;
input x194;
input x195;
input x196;
input x197;
input x198;
input x199;
input x200;
input x201;
input x202;
input x203;
input x204;
input x205;
input x206;
input x207;
input x208;
input x209;
input x210;
input x211;
input x212;
input x213;
input x214;
input x215;
input x216;
input x217;
input x218;
input x219;
input x220;
input x221;
input x222;
input x223;
input x224;
input x225;
input x226;
input x227;
input x228;
input x229;
input x230;
input x231;
input x232;
input x233;
input x234;
input x235;
input x236;
input x237;
input x238;
input x239;
input x240;
input x241;
input x242;
input x243;
input x244;
input x245;
input x246;
input x247;
input x248;
input x249;
input x250;
input x251;
input x252;
input x253;
input x254;
input x255;
input x256;
input x257;
input x258;
input x259;
input x260;
input x261;
input x262;
input x263;
input x264;
input x265;
input x266;
input x267;
input x268;
input x269;
input x270;
input x271;
input x272;
input x273;
input x274;
input x275;
input x276;
input x277;
input x278;
input x279;
input x280;
input x281;
input x282;
input x283;
input x284;
input x285;
input x286;
input x287;
input x288;
input x289;
input x290;
input x291;
input x292;
input x293;
input x294;
input x295;
input x296;
input x297;
input x298;
input x299;
input x300;
input x301;
input x302;
input x303;
input x304;
input x305;
input x306;
input x307;
input x308;
input x309;
input x310;
input x311;
input x312;
input x313;
input x314;
input x315;
input x316;
input x317;
input x318;
input x319;
input x320;
input x321;
input x322;
input x323;
input x324;
input x325;
input x326;
input x327;
input x328;
input x329;
input x330;
input x331;
input x332;
input x333;
input x334;
input x335;
input x336;
input x337;
input x338;
input x339;
input x340;
input x341;
input x342;
input x343;
input x344;
input x345;
input x346;
input x347;
input x348;
input x349;
input x350;
input x351;
input x352;
input x353;
input x354;
input x355;
input x356;
input x357;
input x358;
input x359;
input x360;
input x361;
input x362;
input x363;
input x364;
input x365;
input x366;
input x367;
input x368;
input x369;
input x370;
input x371;
input x372;
input x373;
input x374;
input x375;
input x376;
input x377;
input x378;
input x379;
input x380;
input x381;
input x382;
input x383;
input x384;
input x385;
input x386;
input x387;
input x388;
input x389;
input x390;
input x391;
input x392;
input x393;
input x394;
input x395;
input x396;
input x397;
input x398;
input x399;
input x400;
input x401;
input x402;
input x403;
input x404;
input x405;
input x406;
input x407;
input x408;
input x409;
input x410;
input x411;
input x412;
input x413;
input x414;
input x415;
input x416;
input x417;
input x418;
input x419;
input x420;
input x421;
input x422;
input x423;
input x424;
input x425;
input x426;
input x427;
input x428;
input x429;
input x430;
input x431;
input x432;
input x433;
input x434;
input x435;
input x436;
input x437;
input x438;
input x439;
input x440;
input x441;
input x442;
input x443;
input x444;
input x445;
input x446;
input x447;
input x448;
input x449;
input x450;
input x451;
input x452;
input x453;
input x454;
input x455;
input x456;
input x457;
input x458;
input x459;
input x460;
input x461;
input x462;
input x463;
input x464;
input x465;
input x466;
input x467;
input x468;
input x469;
input x470;
input x471;
input x472;
input x473;
input x474;
input x475;
input x476;
input x477;
input x478;
input x479;
input x480;
input x481;
input x482;
input x483;
input x484;
input x485;
input x486;
input x487;
input x488;
input x489;
input x490;
input x491;
input x492;
input x493;
input x494;
input x495;
input x496;
input x497;
input x498;
input x499;
input x500;
input x501;
input x502;
input x503;
input x504;
input x505;
input x506;
input x507;
input x508;
input x509;
input x510;
input x511;
input x512;
input x513;
input x514;
input x515;
input x516;
input x517;
input x518;
input x519;
input x520;
input x521;
input x522;
input x523;
input x524;
input x525;
input x526;
input x527;
input x528;
input x529;
input x530;
input x531;
input x532;
input x533;
input x534;
input x535;
input x536;
input x537;
input x538;
input x539;
input x540;
input x541;
input x542;
input x543;
input x544;
input x545;
input x546;
input x547;
input x548;
input x549;
input x550;
input x551;
input x552;
input x553;
input x554;
input x555;
input x556;
input x557;
input x558;
input x559;
input x560;
input x561;
input x562;
input x563;
input x564;
input x565;
input x566;
input x567;
input x568;
input x569;
input x570;
input x571;
input x572;
input x573;
input x574;
input x575;
input x576;
input x577;
input x578;
input x579;
input x580;
input x581;
input x582;
input x583;
input x584;
input x585;
input x586;
input x587;
input x588;
input x589;
input x590;
input x591;
input x592;
input x593;
input x594;
input x595;
input x596;
input x597;
input x598;
input x599;
input x600;
input x601;
input x602;
input x603;
input x604;
input x605;
input x606;
input x607;
input x608;
input x609;
input x610;
input x611;
input x612;
input x613;
input x614;
input x615;
input x616;
input x617;
input x618;
input x619;
input x620;
input x621;
input x622;
input x623;
input x624;
input x625;
input x626;
input x627;
input x628;
input x629;
input x630;
input x631;
input x632;
input x633;
input x634;
input x635;
input x636;
input x637;
input x638;
input x639;
input x640;
input x641;
input x642;
input x643;
input x644;
input x645;
input x646;
input x647;
input x648;
input x649;
input x650;
input x651;
input x652;
input x653;
input x654;
input x655;
input x656;
input x657;
input x658;
input x659;
input x660;
input x661;
input x662;
input x663;
input x664;
input x665;
input x666;
input x667;
input x668;
input x669;
input x670;
input x671;
input x672;
input x673;
input x674;
input x675;
input x676;
input x677;
input x678;
input x679;
input x680;
input x681;
input x682;
input x683;
input x684;
input x685;
input x686;
input x687;
input x688;
input x689;
input x690;
input x691;
input x692;
input x693;
input x694;
input x695;
input x696;
input x697;
input x698;
input x699;
input x700;
input x701;
input x702;
input x703;
input x704;
input x705;
input x706;
input x707;
input x708;
input x709;
input x710;
input x711;
input x712;
input x713;
input x714;
input x715;
input x716;
input x717;
input x718;
input x719;
input x720;
input x721;
input x722;
input x723;
input x724;
input x725;
input x726;
input x727;
input x728;
input x729;
input x730;
input x731;
input x732;
input x733;
input x734;
input x735;
input x736;
input x737;
input x738;
input x739;
input x740;
input x741;
input x742;
input x743;
input x744;
input x745;
input x746;
input x747;
input x748;
input x749;
input x750;
input x751;
input x752;
input x753;
input x754;
input x755;
input x756;
input x757;
input x758;
input x759;
input x760;
input x761;
input x762;
input x763;
input x764;
input x765;
input x766;
input x767;
input x768;
input x769;
input x770;
input x771;
input x772;
input x773;
input x774;
input x775;
input x776;
input x777;
input x778;
input x779;
input x780;
input x781;
input x782;
input x783;
output c07;
output c615;
output c0273;
output c464;
output c011;
output c126;
output c439;
output c1125;
output c3286;
output c7146;
output c4276;
output c528;
output c5230;
output c1289;
output c9161;
output c7145;
output c359;
output c4144;
output c029;
output c680;
output c0219;
output c880;
output c6206;
output c925;
output c0150;
output c546;
output c9225;
output c0201;
output c0191;
output c5260;
output c6251;
output c4235;
output c967;
output c9141;
output c084;
output c1201;
output c7243;
output c8127;
output c587;
output c2283;
output c3210;
output c530;
output c934;
output c0199;
output c5160;
output c6105;
output c458;
output c5217;
output c4292;
output c21;
output c599;
output c6264;
output c736;
output c8188;
output c322;
output c3200;
output c9126;
output c7228;
output c6110;
output c6228;
output c388;
output c0181;
output c547;
output c492;
output c592;
output c295;
output c190;
output c6139;
output c88;
output c0141;
output c4125;
output c664;
output c9198;
output c5184;
output c090;
output c1133;
output c2289;
output c175;
output c4238;
output c1176;
output c4209;
output c0184;
output c5214;
output c525;
output c5127;
output c2236;
output c749;
output c8155;
output c1150;
output c0105;
output c6291;
output c974;
output c9142;
output c7209;
output c51;
output c9154;
output c3288;
output c5131;
output c4219;
output c0156;
output c214;
output c4229;
output c6278;
output c8170;
output c924;
output c0237;
output c366;
output c9183;
output c168;
output c9283;
output c9166;
output c964;
output c118;
output c1259;
output c6242;
output c293;
output c5235;
output c7211;
output c2190;
output c2233;
output c3148;
output c398;
output c1298;
output c259;
output c4180;
output c0161;
output c2250;
output c68;
output c7264;
output c7294;
output c9127;
output c1299;
output c1143;
output c3110;
output c9262;
output c0122;
output c25;
output c298;
output c328;
output c6118;
output c376;
output c864;
output c8112;
output c762;
output c6142;
output c0218;
output c245;
output c6103;
output c9185;
output c6231;
output c5225;
output c1117;
output c6114;
output c1197;
output c8251;
output c048;
output c6158;
output c5292;
output c1152;
output c2256;
output c2155;
output c8145;
output c7289;
output c710;
output c8246;
output c4163;
output c5118;
output c24;
output c7292;
output c088;
output c821;
output c223;
output c3293;
output c930;
output c396;
output c0265;
output c3218;
output c6208;
output c7116;
output c5255;
output c095;
output c7100;
output c3155;
output c621;
output c078;
output c249;
output c297;
output c5159;
output c1239;
output c4227;
output c2151;
output c5254;
output c3146;
output c537;
output c6165;
output c129;
output c4246;
output c665;
output c2213;
output c7299;
output c1100;
output c8288;
output c839;
output c580;
output c2220;
output c09;
output c757;
output c779;
output c1225;
output c8161;
output c0148;
output c211;
output c716;
output c6101;
output c6214;
output c798;
output c4241;
output c354;
output c8179;
output c9232;
output c65;
output c423;
output c4271;
output c7213;
output c4256;
output c631;
output c972;
output c844;
output c4143;
output c0228;
output c1128;
output c036;
output c0137;
output c794;
output c0206;
output c2242;
output c9205;
output c9137;
output c945;
output c53;
output c1156;
output c6104;
output c777;
output c0252;
output c367;
output c8254;
output c5170;
output c7274;
output c7262;
output c047;
output c0294;
output c7219;
output c6108;
output c2128;
output c6273;
output c987;
output c8243;
output c9231;
output c9218;
output c092;
output c4107;
output c0171;
output c043;
output c6217;
output c0276;
output c4199;
output c4228;
output c541;
output c8187;
output c393;
output c9147;
output c720;
output c1105;
output c1144;
output c427;
output c0144;
output c7120;
output c0288;
output c5247;
output c954;
output c1258;
output c9189;
output c0277;
output c69;
output c8174;
output c2116;
output c5136;
output c759;
output c614;
output c3240;
output c1180;
output c8122;
output c9148;
output c9259;
output c784;
output c4130;
output c2115;
output c6265;
output c2176;
output c2251;
output c763;
output c589;
output c699;
output c6136;
output c151;
output c8255;
output c5222;
output c4223;
output c596;
output c4245;
output c032;
output c3165;
output c5155;
output c6298;
output c7197;
output c848;
output c8196;
output c0165;
output c473;
output c566;
output c079;
output c6286;
output c782;
output c7202;
output c9214;
output c2211;
output c0239;
output c521;
output c221;
output c0153;
output c1267;
output c361;
output c075;
output c2154;
output c456;
output c241;
output c2244;
output c3291;
output c7154;
output c9263;
output c670;
output c2276;
output c2189;
output c1183;
output c3287;
output c072;
output c2225;
output c3184;
output c0207;
output c894;
output c9134;
output c9203;
output c8194;
output c8147;
output c498;
output c7251;
output c4178;
output c7183;
output c39;
output c3132;
output c1164;
output c3267;
output c9191;
output c116;
output c852;
output c742;
output c7180;
output c6195;
output c0159;
output c3254;
output c3177;
output c9224;
output c0270;
output c4160;
output c2142;
output c6156;
output c7204;
output c1122;
output c4288;
output c4265;
output c60;
output c7257;
output c1139;
output c7290;
output c1252;
output c522;
output c5271;
output c5224;
output c061;
output c115;
output c9292;
output c8191;
output c970;
output c9107;
output c9210;
output c419;
output c6146;
output c1135;
output c3233;
output c331;
output c831;
output c2241;
output c6187;
output c7248;
output c941;
output c063;
output c4259;
output c1238;
output c9213;
output c554;
output c918;
output c338;
output c861;
output c885;
output c2170;
output c1296;
output c1279;
output c2238;
output c2119;
output c3131;
output c3181;
output c5106;
output c575;
output c645;
output c7270;
output c4150;
output c985;
output c2185;
output c940;
output c616;
output c889;
output c545;
output c313;
output c0284;
output c5223;
output c5137;
output c8148;
output c320;
output c2265;
output c3180;
output c94;
output c937;
output c3142;
output c955;
output c0128;
output c8171;
output c0286;
output c7254;
output c451;
output c428;
output c1162;
output c5168;
output c7293;
output c3187;
output c185;
output c3284;
output c1169;
output c1234;
output c7143;
output c2194;
output c4218;
output c881;
output c3178;
output c7200;
output c40;
output c5203;
output c3271;
output c4298;
output c0167;
output c3169;
output c20;
output c590;
output c0204;
output c6258;
output c485;
output c7286;
output c1229;
output c025;
output c0197;
output c89;
output c8214;
output c6182;
output c6111;
output c6295;
output c30;
output c6266;
output c866;
output c6154;
output c261;
output c5280;
output c34;
output c466;
output c4106;
output c4149;
output c9228;
output c3183;
output c6173;
output c8181;
output c3281;
output c5252;
output c5122;
output c1281;
output c986;
output c7265;
output c890;
output c437;
output c12;
output c4112;
output c5185;
output c4258;
output c3292;
output c8263;
output c1188;
output c285;
output c379;
output c5130;
output c363;
output c454;
output c8208;
output c2161;
output c4172;
output c7110;
output c8257;
output c4250;
output c734;
output c049;
output c114;
output c0126;
output c7173;
output c6184;
output c7208;
output c5150;
output c6122;
output c1286;
output c4101;
output c951;
output c340;
output c181;
output c0215;
output c383;
output c141;
output c2124;
output c8225;
output c4239;
output c9230;
output c9242;
output c8294;
output c2150;
output c1126;
output c3258;
output c3265;
output c1295;
output c862;
output c4127;
output c1241;
output c778;
output c79;
output c6121;
output c018;
output c1193;
output c8121;
output c9162;
output c5153;
output c6289;
output c8242;
output c2181;
output c555;
output c582;
output c0187;
output c033;
output c1142;
output c7194;
output c2280;
output c77;
output c3108;
output c5147;
output c4167;
output c613;
output c915;
output c7214;
output c1290;
output c2262;
output c0119;
output c4277;
output c41;
output c9180;
output c7184;
output c7178;
output c7205;
output c069;
output c0229;
output c7157;
output c944;
output c2231;
output c9200;
output c874;
output c694;
output c7217;
output c2235;
output c8137;
output c9273;
output c729;
output c1190;
output c657;
output c1246;
output c5149;
output c6220;
output c543;
output c4214;
output c6175;
output c053;
output c3100;
output c7263;
output c836;
output c9254;
output c349;
output c8207;
output c6120;
output c337;
output c2222;
output c6180;
output c4204;
output c2199;
output c6210;
output c5250;
output c424;
output c042;
output c0248;
output c9247;
output c659;
output c7285;
output c264;
output c4187;
output c3138;
output c2273;
output c756;
output c766;
output c8205;
output c6283;
output c8266;
output c6163;
output c5205;
output c7210;
output c7170;
output c2297;
output c5105;
output c1219;
output c3243;
output c3127;
output c0236;
output c0113;
output c390;
output c9265;
output c3111;
output c4102;
output c2261;
output c476;
output c8227;
output c4152;
output c13;
output c6194;
output c4253;
output c5204;
output c642;
output c80;
output c461;
output c1111;
output c0140;
output c6128;
output c7241;
output c3241;
output c436;
output c8200;
output c172;
output c5236;
output c2180;
output c5288;
output c086;
output c284;
output c9105;
output c5296;
output c2131;
output c5278;
output c5287;
output c198;
output c0152;
output c1194;
output c1157;
output c6135;
output c5277;
output c2164;
output c558;
output c5213;
output c4222;
output c2138;
output c8163;
output c368;
output c369;
output c4110;
output c5157;
output c164;
output c5191;
output c4282;
output c443;
output c7164;
output c0182;
output c4224;
output c45;
output c4262;
output c0189;
output c4197;
output c19;
output c0102;
output c9184;
output c4115;
output c046;
output c0295;
output c627;
output c0160;
output c1216;
output c3221;
output c2224;
output c0151;
output c345;
output c4161;
output c3204;
output c563;
output c137;
output c226;
output c386;
output c690;
output c7207;
output c0287;
output c022;
output c5265;
output c8264;
output c7108;
output c6124;
output c3276;
output c9176;
output c2166;
output c3172;
output c5110;
output c045;
output c8219;
output c872;
output c0209;
output c1287;
output c0269;
output c3112;
output c4153;
output c5154;
output c6157;
output c4158;
output c6189;
output c7152;
output c7275;
output c1209;
output c9279;
output c8151;
output c938;
output c7297;
output c0106;
output c0123;
output c4168;
output c75;
output c362;
output c9167;
output c1160;
output c271;
output c559;
output c1231;
output c332;
output c2201;
output c9102;
output c655;
output c0101;
output c2253;
output c3153;
output c462;
output c7150;
output c3158;
output c935;
output c9174;
output c2218;
output c980;
output c8277;
output c8283;
output c2100;
output c6152;
output c429;
output c725;
output c6280;
output c72;
output c373;
output c10;
output c2249;
output c7189;
output c576;
output c2109;
output c6272;
output c247;
output c786;
output c7199;
output c816;
output c4296;
output c9135;
output c3299;
output c5234;
output c71;
output c968;
output c1269;
output c3122;
output c333;
output c9160;
output c7112;
output c629;
output c460;
output c572;
output c3277;
output c6239;
output c021;
output c0242;
output c3117;
output c4183;
output c1102;
output c8282;
output c1282;
output c425;
output c5263;
output c9112;
output c9156;
output c060;
output c136;
output c5100;
output c3248;
output c1154;
output c0147;
output c239;
output c1243;
output c6224;
output c3215;
output c845;
output c1173;
output c1113;
output c9115;
output c272;
output c2205;
output c5144;
output c1233;
output c270;
output c023;
output c6252;
output c83;
output c3168;
output c8185;
output c0155;
output c5228;
output c963;
output c319;
output c2139;
output c2247;
output c3216;
output c828;
output c9129;
output c9229;
output c1149;
output c134;
output c971;
output c188;
output c693;
output c58;
output c5108;
output c0142;
output c531;
output c5114;
output c721;
output c299;
output c7249;
output c49;
output c5129;
output c3198;
output c553;
output c5192;
output c232;
output c5197;
output c689;
output c7124;
output c99;
output c825;
output c1274;
output c4299;
output c6144;
output c0283;
output c752;
output c2195;
output c5146;
output c4138;
output c6192;
output c9204;
output c0175;
output c252;
output c040;
output c2208;
output c4192;
output c978;
output c9208;
output c3104;
output c3189;
output c165;
output c4182;
output c1112;
output c494;
output c8107;
output c9149;
output c5196;
output c167;
output c9216;
output c3217;
output c579;
output c1163;
output c213;
output c4131;
output c4135;
output c4207;
output c9234;
output c0115;
output c8285;
output c8235;
output c7172;
output c529;
output c121;
output c52;
output c1277;
output c347;
output c1236;
output c1202;
output c2254;
output c5257;
output c62;
output c098;
output c1250;
output c364;
output c7196;
output c1266;
output c3219;
output c184;
output c5282;
output c158;
output c6260;
output c931;
output c6193;
output c0253;
output c8197;
output c6293;
output c6150;
output c5261;
output c6190;
output c711;
output c5152;
output c1251;
output c074;
output c2165;
output c636;
output c6130;
output c569;
output c5209;
output c3234;
output c6100;
output c8212;
output c714;
output c4275;
output c3235;
output c8109;
output c9146;
output c5276;
output c7246;
output c316;
output c552;
output c495;
output c0235;
output c7291;
output c43;
output c5161;
output c571;
output c943;
output c3114;
output c3227;
output c2144;
output c076;
output c7279;
output c8111;
output c776;
output c2177;
output c5158;
output c671;
output c9240;
output c268;
output c6243;
output c5174;
output c5111;
output c859;
output c649;
output c887;
output c556;
output c5125;
output c235;
output c9159;
output c1212;
output c5264;
output c2196;
output c1245;
output c540;
output c33;
output c7118;
output c9296;
output c6166;
output c6170;
output c911;
output c0212;
output c8290;
output c2270;
output c161;
output c1124;
output c1232;
output c8274;
output c0136;
output c6285;
output c1170;
output c946;
output c526;
output c515;
output c2232;
output c5182;
output c5258;
output c399;
output c0198;
output c927;
output c479;
output c5166;
output c995;
output c942;
output c1148;
output c382;
output c2130;
output c4129;
output c9291;
output c1179;
output c9243;
output c4155;
output c0247;
output c1181;
output c174;
output c3296;
output c4252;
output c883;
output c92;
output c421;
output c1222;
output c446;
output c5132;
output c5206;
output c7162;
output c1214;
output c997;
output c171;
output c891;
output c8154;
output c0200;
output c920;
output c9118;
output c3209;
output c29;
output c2210;
output c1228;
output c0293;
output c489;
output c9139;
output c3255;
output c1254;
output c1177;
output c0272;
output c0281;
output c5269;
output c7121;
output c3174;
output c493;
output c750;
output c0192;
output c374;
output c577;
output c728;
output c7192;
output c6181;
output c8136;
output c0268;
output c2263;
output c8128;
output c6253;
output c5218;
output c981;
output c854;
output c7206;
output c414;
output c2198;
output c879;
output c7131;
output c2287;
output c4260;
output c1136;
output c7273;
output c868;
output c263;
output c6262;
output c027;
output c877;
output c1208;
output c1297;
output c342;
output c0254;
output c78;
output c135;
output c6137;
output c7187;
output c068;
output c644;
output c375;
output c667;
output c155;
output c8206;
output c9245;
output c1165;
output c142;
output c9257;
output c9144;
output c2160;
output c676;
output c066;
output c166;
output c336;
output c656;
output c739;
output c6117;
output c837;
output c6125;
output c2126;
output c2169;
output c5259;
output c583;
output c992;
output c775;
output c989;
output c5295;
output c70;
output c267;
output c27;
output c7101;
output c1168;
output c9297;
output c5299;
output c9235;
output c0221;
output c850;
output c2239;
output c3182;
output c1172;
output c8226;
output c6141;
output c4215;
output c5198;
output c0114;
output c0261;
output c6219;
output c138;
output c4170;
output c923;
output c523;
output c9271;
output c0203;
output c4272;
output c5109;
output c4132;
output c6234;
output c3214;
output c3253;
output c2277;
output c1270;
output c5220;
output c9207;
output c5102;
output c824;
output c8279;
output c1182;
output c3226;
output c5186;
output c684;
output c7171;
output c8265;
output c4251;
output c3145;
output c5128;
output c6249;
output c581;
output c9206;
output c7115;
output c0143;
output c9188;
output c3159;
output c256;
output c3263;
output c6126;
output c8166;
output c8271;
output c2125;
output c8275;
output c3270;
output c949;
output c1108;
output c8102;
output c910;
output c377;
output c052;
output c019;
output c3124;
output c9187;
output c397;
output c3207;
output c260;
output c9241;
output c8231;
output c378;
output c7168;
output c628;
output c119;
output c6237;
output c6199;
output c2135;
output c5162;
output c224;
output c6276;
output c6160;
output c197;
output c6267;
output c5212;
output c246;
output c497;
output c2132;
output c7161;
output c1213;
output c04;
output c7216;
output c6102;
output c4148;
output c95;
output c2117;
output c150;
output c8261;
output c6221;
output c8281;
output c9275;
output c5298;
output c669;
output c519;
output c274;
output c3290;
output c772;
output c4213;
output c5178;
output c7158;
output c510;
output c548;
output c430;
output c744;
output c0176;
output c4266;
output c3107;
output c2108;
output c457;
output c5231;
output c132;
output c832;
output c4123;
output c7151;
output c1263;
output c884;
output c3102;
output c8248;
output c2203;
output c028;
output c1175;
output c6223;
output c9299;
output c4166;
output c097;
output c567;
output c5294;
output c8220;
output c3154;
output c3197;
output c4165;
output c3245;
output c6248;
output c4226;
output c496;
output c1151;
output c0214;
output c966;
output c947;
output c0249;
output c818;
output c255;
output c7255;
output c3249;
output c2258;
output c830;
output c8278;
output c4139;
output c7137;
output c189;
output c4243;
output c594;
output c8291;
output c9249;
output c8286;
output c1280;
output c2294;
output c1247;
output c070;
output c3105;
output c7142;
output c4286;
output c624;
output c1226;
output c4174;
output c0230;
output c453;
output c654;
output c7256;
output c0132;
output c4255;
output c64;
output c0243;
output c1207;
output c6284;
output c6145;
output c9181;
output c5242;
output c8139;
output c3133;
output c686;
output c0193;
output c4237;
output c9136;
output c2186;
output c3128;
output c348;
output c849;
output c0133;
output c3190;
output c03;
output c465;
output c838;
output c6116;
output c156;
output c2200;
output c6241;
output c0205;
output c8125;
output c0223;
output c7156;
output c8141;
output c591;
output c1184;
output c2197;
output c916;
output c2259;
output c1271;
output c2192;
output c612;
output c7231;
output c2293;
output c730;
output c6168;
output c743;
output c8240;
output c9197;
output c0100;
output c4208;
output c2223;
output c0178;
output c8153;
output c0233;
output c8215;
output c4140;
output c3242;
output c6205;
output c5177;
output c7138;
output c6236;
output c3162;
output c5270;
output c6244;
output c6235;
output c6162;
output c486;
output c4133;
output c038;
output c7165;
output c4105;
output c1118;
output c1278;
output c5101;
output c8198;
output c9100;
output c8272;
output c448;
output c754;
output c467;
output c765;
output c131;
output c4291;
output c4195;
output c5244;
output c275;
output c244;
output c394;
output c2228;
output c2120;
output c4225;
output c564;
output c797;
output c6169;
output c8115;
output c8298;
output c5117;
output c2272;
output c4154;
output c5104;
output c9172;
output c7227;
output c851;
output c442;
output c2105;
output c3171;
output c8201;
output c0202;
output c9268;
output c6202;
output c145;
output c8292;
output c2129;
output c2163;
output c148;
output c9186;
output c0255;
output c3261;
output c3297;
output c1129;
output c0241;
output c0138;
output c5240;
output c0121;
output c9132;
output c3119;
output c0264;
output c2122;
output c2102;
output c6246;
output c9199;
output c077;
output c1155;
output c8195;
output c227;
output c6133;
output c3205;
output c2148;
output c8114;
output c7149;
output c218;
output c0274;
output c962;
output c9277;
output c2110;
output c0224;
output c2147;
output c1167;
output c7239;
output c9195;
output c9151;
output c4128;
output c248;
output c2295;
output c731;
output c7177;
output c5139;
output c9222;
output c0190;
output c633;
output c3199;
output c593;
output c912;
output c584;
output c1288;
output c4206;
output c288;
output c4297;
output c1198;
output c688;
output c173;
output c610;
output c8183;
output c2217;
output c993;
output c030;
output c8140;
output c194;
output c157;
output c1273;
output c640;
output c250;
output c9106;
output c8184;
output c5237;
output c1200;
output c4295;
output c86;
output c8268;
output c6177;
output c8221;
output c2106;
output c7193;
output c8160;
output c4114;
output c1265;
output c2214;
output c123;
output c5283;
output c8239;
output c2269;
output c9290;
output c16;
output c2267;
output c991;
output c7222;
output c5273;
output c3134;
output c799;
output c450;
output c4263;
output c7221;
output c2121;
output c751;
output c0134;
output c468;
output c2207;
output c3222;
output c7280;
output c8108;
output c0110;
output c3120;
output c7284;
output c1101;
output c0222;
output c1147;
output c0154;
output c93;
output c3201;
output c3272;
output c035;
output c472;
output c6127;
output c9261;
output c5135;
output c999;
output c8180;
output c820;
output c9294;
output c4171;
output c449;
output c389;
output c433;
output c0280;
output c1210;
output c483;
output c8204;
output c133;
output c191;
output c9212;
output c3274;
output c1211;
output c764;
output c1255;
output c7105;
output c220;
output c7136;
output c712;
output c792;
output c7266;
output c588;
output c3232;
output c733;
output c262;
output c4269;
output c8284;
output c3166;
output c4177;
output c2145;
output c8297;
output c010;
output c5285;
output c741;
output c4198;
output c0120;
output c094;
output c7195;
output c8172;
output c8164;
output c544;
output c746;
output c7133;
output c1221;
output c410;
output c0238;
output c176;
output c6176;
output c2298;
output c417;
output c1192;
output c3125;
output c678;
output c0245;
output c3163;
output c7117;
output c626;
output c785;
output c55;
output c888;
output c4254;
output c5175;
output c44;
output c1132;
output c9163;
output c9202;
output c1110;
output c562;
output c9168;
output c7122;
output c3140;
output c4279;
output c7181;
output c512;
output c7160;
output c330;
output c740;
output c7190;
output c899;
output c8262;
output c3152;
output c956;
output c7128;
output c3103;
output c0257;
output c422;
output c5227;
output c17;
output c9215;
output c1145;
output c1186;
output c323;
output c3206;
output c755;
output c698;
output c9253;
output c3231;
output c9211;
output c5290;
output c3279;
output c3275;
output c6149;
output c939;
output c243;
output c2174;
output c895;
output c9256;
output c7126;
output c933;
output c6174;
output c3160;
output c280;
output c994;
output c0263;
output c3257;
output c35;
output c8295;
output c26;
output c857;
output c998;
output c957;
output c0117;
output c961;
output c055;
output c5169;
output c5165;
output c344;
output c487;
output c392;
output c9280;
output c565;
output c6287;
output c758;
output c3208;
output c8133;
output c7258;
output c7191;
output c8256;
output c97;
output c9124;
output c117;
output c1230;
output c771;
output c8247;
output c660;
output c4261;
output c61;
output c3252;
output c153;
output c3236;
output c842;
output c8260;
output c7144;
output c713;
output c9175;
output c871;
output c0104;
output c7276;
output c7169;
output c619;
output c2282;
output c1185;
output c4120;
output c5208;
output c9272;
output c4210;
output c1260;
output c9286;
output c6153;
output c9196;
output c057;
output c3239;
output c535;
output c7212;
output c6203;
output c2246;
output c2193;
output c4124;
output c499;
output c9246;
output c1106;
output c9282;
output c4116;
output c4126;
output c9133;
output c8158;
output c237;
output c1141;
output c357;
output c4188;
output c1272;
output c1256;
output c3295;
output c183;
output c4249;
output c8103;
output c9178;
output c9113;
output c276;
output c455;
output c865;
output c0194;
output c7236;
output c814;
output c5239;
output c435;
output c6155;
output c286;
output c0282;
output c7139;
output c0211;
output c0289;
output c4242;
output c1161;
output c6263;
output c873;
output c9173;
output c7159;
output c3278;
output c732;
output c238;
output c8218;
output c9143;
output c416;
output c9258;
output c952;
output c2103;
output c4264;
output c7111;
output c3135;
output c863;
output c3237;
output c4184;
output c02;
output c215;
output c719;
output c0196;
output c5291;
output c1293;
output c7282;
output c913;
output c0244;
output c8237;
output c7252;
output c8287;
output c356;
output c1159;
output c3144;
output c973;
output c637;
output c897;
output c5246;
output c3246;
output c516;
output c8168;
output c723;
output c1285;
output c6288;
output c7153;
output c5142;
output c536;
output c0116;
output c56;
output c1220;
output c8224;
output c8126;
output c130;
output c6171;
output c5219;
output c598;
output c9217;
output c8202;
output c2187;
output c2127;
output c8252;
output c858;
output c0226;
output c2292;
output c4185;
output c159;
output c685;
output c326;
output c1114;
output c796;
output c7129;
output c892;
output c441;
output c0179;
output c4151;
output c265;
output c32;
output c738;
output c2162;
output c1174;
output c514;
output c6274;
output c3256;
output c6185;
output c8167;
output c234;
output c381;
output c8211;
output c371;
output c7188;
output c622;
output c635;
output c781;
output c0125;
output c9121;
output c4270;
output c4202;
output c2101;
output c9190;
output c5262;
output c9120;
output c9103;
output c2137;
output c46;
output c4111;
output c2264;
output c310;
output c5103;
output c5266;
output c0118;
output c2234;
output c4211;
output c557;
output c0124;
output c186;
output c666;
output c5124;
output c9264;
output c6164;
output c0260;
output c085;
output c160;
output c216;
output c5167;
output c4176;
output c5272;
output c8117;
output c7287;
output c2229;
output c7186;
output c0285;
output c788;
output c8250;
output c2281;
output c6196;
output c6292;
output c8105;
output c691;
output c1275;
output c3116;
output c149;
output c8216;
output c87;
output c3141;
output c432;
output c745;
output c6212;
output c661;
output c2290;
output c7220;
output c812;
output c856;
output c0173;
output c020;
output c5215;
output c8222;
output c4189;
output c081;
output c06;
output c351;
output c0290;
output c8192;
output c5183;
output c5274;
output c7245;
output c3170;
output c7223;
output c7296;
output c7247;
output c767;
output c8119;
output c289;
output c2167;
output c2156;
output c469;
output c822;
output c7277;
output c199;
output c380;
output c7167;
output c2158;
output c8165;
output c73;
output c4104;
output c641;
output c127;
output c0166;
output c840;
output c3244;
output c922;
output c1284;
output c7233;
output c5210;
output c9164;
output c0251;
output c054;
output c463;
output c5195;
output c9239;
output c4289;
output c8152;
output c1242;
output c6119;
output c5194;
output c8249;
output c8106;
output c6159;
output c9150;
output c632;
output c4201;
output c4196;
output c1127;
output c0213;
output c3143;
output c8176;
output c9295;
output c5253;
output c1204;
output c672;
output c236;
output c768;
output c5243;
output c484;
output c7203;
output c253;
output c9248;
output c726;
output c3230;
output c339;
output c652;
output c977;
output c0158;
output c724;
output c6218;
output c6255;
output c7135;
output c718;
output c254;
output c6179;
output c982;
output c841;
output c279;
output c1166;
output c8129;
output c026;
output c6222;
output c258;
output c5138;
output c2248;
output c9108;
output c3136;
output c242;
output c7259;
output c1119;
output c192;
output c4147;
output c780;
output c1109;
output c3106;
output c2279;
output c4273;
output c0162;
output c6147;
output c212;
output c5233;
output c3192;
output c1146;
output c2202;
output c9220;
output c481;
output c7106;
output c48;
output c7132;
output c2221;
output c2175;
output c6186;
output c90;
output c9170;
output c0135;
output c3101;
output c5141;
output c787;
output c080;
output c3280;
output c789;
output c7237;
output c4181;
output c74;
output c290;
output c9153;
output c8182;
output c140;
output c677;
output c31;
output c2299;
output c9193;
output c5216;
output c6167;
output c28;
output c5163;
output c9110;
output c9233;
output c0149;
output c452;
output c4136;
output c5279;
output c42;
output c8120;
output c067;
output c674;
output c0298;
output c8189;
output c3251;
output c7261;
output c976;
output c959;
output c4173;
output c2172;
output c4169;
output c6188;
output c3188;
output c0112;
output c2268;
output c4146;
output c96;
output c6238;
output c0109;
output c196;
output c1104;
output c819;
output c7260;
output c9219;
output c9223;
output c7147;
output c122;
output c511;
output c039;
output c761;
output c7179;
output c5115;
output c4267;
output c5248;
output c1235;
output c287;
output c3211;
output c5133;
output c2204;
output c8134;
output c542;
output c152;
output c7114;
output c3212;
output c8132;
output c6134;
output c7107;
output c513;
output c324;
output c1121;
output c8169;
output c210;
output c843;
output c5201;
output c936;
output c099;
output c2111;
output c00;
output c8203;
output c869;
output c3285;
output c2266;
output c57;
output c8241;
output c847;
output c8190;
output c1116;
output c9119;
output c9130;
output c550;
output c737;
output c1237;
output c3294;
output c5176;
output c2123;
output c2171;
output c870;
output c083;
output c4159;
output c2245;
output c459;
output c520;
output c4247;
output c7238;
output c0297;
output c1107;
output c2140;
output c896;
output c9194;
output c893;
output c7103;
output c8213;
output c3191;
output c1203;
output c0163;
output c8130;
output c2278;
output c9227;
output c0256;
output c6172;
output c8131;
output c735;
output c418;
output c3179;
output c412;
output c7295;
output c91;
output c63;
output c3196;
output c5200;
output c2209;
output c6198;
output c8293;
output c0231;
output c7229;
output c9201;
output c8162;
output c8149;
output c538;
output c620;
output c434;
output c6257;
output c0291;
output c4175;
output c8236;
output c5107;
output c1120;
output c7104;
output c8157;
output c7141;
output c1171;
output c1205;
output c05;
output c517;
output c791;
output c2257;
output c111;
output c8230;
output c0258;
output c929;
output c7253;
output c2134;
output c7250;
output c315;
output c0111;
output c2112;
output c647;
output c182;
output c1195;
output c6138;
output c447;
output c426;
output c9101;
output c041;
output c790;
output c8273;
output c3161;
output c8245;
output c663;
output c1294;
output c0131;
output c1283;
output c0266;
output c231;
output c5256;
output c5211;
output c1292;
output c0172;
output c4244;
output c7244;
output c6240;
output c9104;
output c5249;
output c1158;
output c662;
output c1264;
output c343;
output c650;
output c4230;
output c1268;
output c722;
output c3202;
output c8289;
output c6131;
output c5143;
output c988;
output c8280;
output c325;
output c3121;
output c5145;
output c311;
output c059;
output c990;
output c0208;
output c9260;
output c411;
output c618;
output c835;
output c6227;
output c277;
output c0278;
output c431;
output c6250;
output c9288;
output c0127;
output c4293;
output c179;
output c9171;
output c717;
output c813;
output c478;
output c490;
output c9278;
output c3109;
output c8156;
output c471;
output c3260;
output c3229;
output c3269;
output c673;
output c139;
output c4232;
output c8110;
output c016;
output c225;
output c8100;
output c6112;
output c327;
output c630;
output c8270;
output c6229;
output c534;
output c9276;
output c9109;
output c124;
output c2143;
output c8143;
output c9122;
output c2118;
output c524;
output c0145;
output c170;
output c195;
output c296;
output c4240;
output c3247;
output c6183;
output c4278;
output c7234;
output c7182;
output c2288;
output c6245;
output c8116;
output c0195;
output c1131;
output c193;
output c294;
output c3164;
output c1189;
output c876;
output c4109;
output c482;
output c8259;
output c6294;
output c7269;
output c5293;
output c37;
output c5297;
output c9274;
output c770;
output c2104;
output c475;
output c9289;
output c037;
output c9298;
output c2260;
output c8296;
output c2291;
output c3225;
output c4274;
output c2133;
output c7130;
output c950;
output c056;
output c8135;
output c0210;
output c867;
output c9145;
output c062;
output c01;
output c15;
output c2159;
output c9192;
output c66;
output c6230;
output c9165;
output c7123;
output c358;
output c3176;
output c4281;
output c7198;
output c8113;
output c0267;
output c1291;
output c3273;
output c6201;
output c9209;
output c783;
output c5164;
output c8217;
output c7224;
output c917;
output c8228;
output c7134;
output c3126;
output c586;
output c846;
output c9226;
output c826;
output c146;
output c14;
output c8144;
output c334;
output c2240;
output c087;
output c0108;
output c1240;
output c853;
output c4284;
output c969;
output c882;
output c318;
output c4156;
output c3139;
output c162;
output c5173;
output c2191;
output c5251;
output c7174;
output c9244;
output c1123;
output c8146;
output c415;
output c4231;
output c715;
output c7102;
output c5187;
output c1244;
output c643;
output c1178;
output c6211;
output c6148;
output c823;
output c4141;
output c1187;
output c539;
output c7215;
output c091;
output c0168;
output c4119;
output c570;
output c8199;
output c2152;
output c064;
output c125;
output c229;
output c4103;
output c065;
output c4285;
output c6297;
output c341;
output c960;
output c9182;
output c6270;
output c3250;
output c3259;
output c0180;
output c793;
output c7235;
output c8118;
output c384;
output c4234;
output c928;
output c0225;
output c67;
output c6161;
output c031;
output c7185;
output c8258;
output c350;
output c251;
output c76;
output c4194;
output c0107;
output c0220;
output c8244;
output c050;
output c0259;
output c4121;
output c2113;
output c291;
output c753;
output c3118;
output c6113;
output c8209;
output c0129;
output c8178;
output c6233;
output c4142;
output c1217;
output c6226;
output c3223;
output c5112;
output c7288;
output c658;
output c6178;
output c7230;
output c6268;
output c773;
output c9236;
output c6282;
output c59;
output c6197;
output c3298;
output c4191;
output c1261;
output c1115;
output c5171;
output c1257;
output c7148;
output c6254;
output c5151;
output c2296;
output c488;
output c257;
output c9138;
output c089;
output c8233;
output c269;
output c638;
output c8138;
output c0186;
output c3113;
output c9157;
output c7125;
output c4122;
output c7175;
output c230;
output c829;
output c4203;
output c0130;
output c4117;
output c6269;
output c0246;
output c5232;
output c491;
output c8223;
output c8124;
output c774;
output c266;
output c0157;
output c2230;
output c321;
output c7272;
output c2243;
output c898;
output c0216;
output c653;
output c98;
output c012;
output c0227;
output c2237;
output c9140;
output c0234;
output c143;
output c1199;
output c3264;
output c5238;
output c834;
output c6191;
output c352;
output c1130;
output c1223;
output c440;
output c7113;
output c815;
output c948;
output c0240;
output c5202;
output c4236;
output c8269;
output c096;
output c6225;
output c760;
output c4280;
output c9155;
output c533;
output c470;
output c3185;
output c7232;
output c3130;
output c574;
output c875;
output c6200;
output c480;
output c282;
output c2285;
output c391;
output c1206;
output c5121;
output c953;
output c921;
output c4268;
output c8276;
output c878;
output c697;
output c7218;
output c18;
output c6299;
output c438;
output c2153;
output c886;
output c2286;
output c395;
output c5120;
output c5134;
output c2178;
output c113;
output c5229;
output c178;
output c4290;
output c0139;
output c617;
output c560;
output c2274;
output c329;
output c47;
output c6107;
output c7226;
output c692;
output c0164;
output c4100;
output c7267;
output c1103;
output c9284;
output c8175;
output c6109;
output c682;
output c233;
output c8232;
output c9293;
output c312;
output c3123;
output c5199;
output c9158;
output c110;
output c2146;
output c8238;
output c5140;
output c4113;
output c2275;
output c860;
output c0262;
output c3151;
output c273;
output c8186;
output c695;
output c8210;
output c9252;
output c926;
output c177;
output c6281;
output c5245;
output c128;
output c0185;
output c595;
output c6247;
output c6275;
output c4179;
output c855;
output c8101;
output c6290;
output c017;
output c3147;
output c2284;
output c5119;
output c687;
output c84;
output c5189;
output c9250;
output c2184;
output c9285;
output c4205;
output c9152;
output c50;
output c4190;
output c9125;
output c3156;
output c013;
output c3150;
output c4233;
output c1276;
output c6207;
output c169;
output c549;
output c2212;
output c578;
output c0169;
output c573;
output c7281;
output c7283;
output c2227;
output c6123;
output c283;
output c360;
output c372;
output c82;
output c093;
output c180;
output c984;
output c5281;
output c2141;
output c7119;
output c965;
output c4217;
output c979;
output c387;
output c228;
output c675;
output c4145;
output c5190;
output c0217;
output c3289;
output c727;
output c6216;
output c1253;
output c474;
output c4193;
output c38;
output c0232;
output c217;
output c679;
output c6215;
output c2226;
output c9111;
output c2255;
output c748;
output c625;
output c747;
output c5172;
output c827;
output c8193;
output c278;
output c9267;
output c919;
output c3224;
output c681;
output c9179;
output c551;
output c163;
output c082;
output c3186;
output c073;
output c051;
output c696;
output c9266;
output c833;
output c5180;
output c6132;
output c112;
output c3262;
output c5284;
output c413;
output c034;
output c292;
output c975;
output c4212;
output c5193;
output c2183;
output c444;
output c668;
output c2271;
output c7155;
output c9237;
output c6143;
output c0275;
output c5226;
output c4220;
output c2173;
output c7163;
output c2114;
output c4164;
output c3195;
output c4283;
output c0174;
output c335;
output c6151;
output c518;
output c8234;
output c648;
output c4108;
output c9117;
output c651;
output c85;
output c9116;
output c9255;
output c0188;
output c3228;
output c4294;
output c9131;
output c1196;
output c2107;
output c0292;
output c3203;
output c4216;
output c014;
output c5221;
output c6256;
output c9269;
output c9251;
output c11;
output c7176;
output c8267;
output c355;
output c2157;
output c071;
output c3283;
output c5188;
output c5275;
output c9270;
output c4137;
output c2216;
output c6271;
output c3220;
output c385;
output c6209;
output c0250;
output c769;
output c7140;
output c983;
output c9169;
output c314;
output c222;
output c4221;
output c36;
output c6296;
output c9177;
output c1153;
output c187;
output c8159;
output c958;
output c6204;
output c1224;
output c4157;
output c147;
output c795;
output c54;
output c6140;
output c561;
output c5207;
output c4200;
output c634;
output c024;
output c8123;
output c1134;
output c044;
output c6279;
output c1227;
output c6106;
output c532;
output c7278;
output c08;
output c810;
output c0170;
output c3137;
output c527;
output c9221;
output c4287;
output c1248;
output c6277;
output c8177;
output c346;
output c3173;
output c7240;
output c477;
output c23;
output c353;
output c9238;
output c1137;
output c0183;
output c3115;
output c445;
output c015;
output c9128;
output c3282;
output c5289;
output c7166;
output c8253;
output c370;
output c8142;
output c5113;
output c2252;
output c5126;
output c9287;
output c4257;
output c6129;
output c22;
output c5116;
output c3175;
output c5268;
output c420;
output c5241;
output c6115;
output c5286;
output c2206;
output c6261;
output c0271;
output c0146;
output c7298;
output c9281;
output c7201;
output c1191;
output c5179;
output c1215;
output c2182;
output c6232;
output c8104;
output c683;
output c9114;
output c365;
output c0103;
output c0177;
output c3194;
output c4248;
output c3149;
output c639;
output c2168;
output c144;
output c811;
output c240;
output c4134;
output c2149;
output c7268;
output c996;
output c7225;
output c585;
output c1138;
output c058;
output c8173;
output c7242;
output c0296;
output c7127;
output c0299;
output c3157;
output c5267;
output c6213;
output c3266;
output c8150;
output c1262;
output c4162;
output c568;
output c817;
output c6259;
output c8229;
output c597;
output c5156;
output c932;
output c7109;
output c3238;
output c154;
output c5148;
output c5181;
output c3167;
output c1218;
output c2215;
output c3193;
output c0279;
output c2188;
output c623;
output c611;
output c8299;
output c2136;
output c914;
output c317;
output c3213;
output c3129;
output c1140;
output c2179;
output c4118;
output c3268;
output c4186;
output c646;
output c1249;
output c219;
output c120;
output c9123;
output c2219;
output c5123;
output c7271;
output c281;
output c81;

assign c00 =  x270 &  x327 &  x347 &  x429 &  x457 &  x513;
assign c02 =  x294 &  x429 &  x430 &  x457 &  x512;
assign c04 =  x297 &  x325 &  x353 &  x375 &  x409 &  x486 & ~x50 & ~x83 & ~x95 & ~x100 & ~x123 & ~x148 & ~x162 & ~x192 & ~x231 & ~x483 & ~x753;
assign c06 =  x442 &  x453 & ~x408 & ~x494;
assign c08 =  x212 &  x440 &  x468 & ~x16 & ~x49 & ~x89 & ~x381 & ~x409 & ~x464 & ~x477 & ~x509 & ~x695 & ~x697 & ~x702 & ~x710 & ~x726 & ~x738 & ~x751;
assign c010 =  x427 &  x538 &  x566 & ~x180 & ~x203 & ~x502;
assign c012 =  x328 &  x375 &  x402 &  x429 &  x456 & ~x231 & ~x234 & ~x235;
assign c014 =  x261 &  x315 &  x316 &  x343 &  x455 & ~x39 & ~x67 & ~x78 & ~x97 & ~x109 & ~x140 & ~x142 & ~x279 & ~x337 & ~x680 & ~x738 & ~x760 & ~x774;
assign c016 =  x212 &  x430 &  x514 & ~x124 & ~x260 & ~x281 & ~x384 & ~x633;
assign c018 =  x327 &  x355 &  x402 &  x458 & ~x235 & ~x286;
assign c020 =  x506;
assign c022 =  x315 &  x370 &  x416;
assign c024 =  x468 &  x495 & ~x3 & ~x45 & ~x50 & ~x59 & ~x67 & ~x78 & ~x79 & ~x84 & ~x101 & ~x109 & ~x112 & ~x120 & ~x164 & ~x168 & ~x221 & ~x277 & ~x279 & ~x313 & ~x369 & ~x381 & ~x382 & ~x409 & ~x471 & ~x472 & ~x555 & ~x582 & ~x607 & ~x708 & ~x710 & ~x745;
assign c026 =  x274 &  x401 &  x511;
assign c028 =  x334 &  x618;
assign c030 =  x30;
assign c032 =  x385 & ~x70 & ~x222 & ~x304 & ~x326 & ~x408 & ~x410 & ~x466 & ~x708;
assign c034 =  x267 &  x327 &  x355 &  x512 &  x540 & ~x29 & ~x88 & ~x274 & ~x446;
assign c036 =  x425 & ~x411;
assign c038 =  x153 &  x207 &  x234 &  x262 &  x269 &  x318;
assign c040 =  x325 &  x409 &  x459 &  x486 &  x514 & ~x176 & ~x373 & ~x511;
assign c042 =  x213 &  x430 &  x486 &  x514 &  x626 & ~x234 & ~x373;
assign c044 =  x5;
assign c046 =  x23;
assign c048 =  x243 &  x387;
assign c050 =  x359 &  x482 & ~x354;
assign c052 =  x299 &  x327 &  x355 &  x375 &  x402 &  x438 &  x568 & ~x234 & ~x523 & ~x562;
assign c054 =  x429 &  x440 &  x457 &  x468 &  x485 &  x496 & ~x160 & ~x224 & ~x436 & ~x538 & ~x595 & ~x645 & ~x678;
assign c056 =  x374 &  x429 &  x456 &  x512 &  x540 &  x568 &  x596 & ~x176 & ~x313 & ~x675 & ~x707 & ~x755;
assign c058 =  x45;
assign c060 =  x401 &  x456 &  x652 & ~x234;
assign c062 =  x425 &  x442;
assign c064 =  x443 &  x498 & ~x438;
assign c066 =  x358 & ~x123 & ~x382 & ~x601;
assign c068 =  x427 &  x455 &  x511 &  x628 & ~x3 & ~x40 & ~x93 & ~x409 & ~x536;
assign c070 =  x275 &  x427 &  x509;
assign c072 =  x643;
assign c074 =  x328 &  x401 &  x511 & ~x203 & ~x632;
assign c076 =  x409 &  x430 & ~x263;
assign c078 =  x659 & ~x63 & ~x293 & ~x381 & ~x409 & ~x437 & ~x492 & ~x503 & ~x548 & ~x574 & ~x575 & ~x589;
assign c080 =  x169;
assign c082 =  x214 &  x372 &  x455 & ~x409 & ~x712 & ~x776;
assign c084 =  x400 &  x566 & ~x578;
assign c086 =  x327 &  x355 &  x430 & ~x176 & ~x234;
assign c088 =  x154 &  x207 &  x262 &  x412 &  x631;
assign c090 =  x346 &  x373 &  x374 &  x401 &  x429 &  x457 &  x513 & ~x21 & ~x46 & ~x123 & ~x162 & ~x176 & ~x204 & ~x259 & ~x313 & ~x408 & ~x537 & ~x580 & ~x758;
assign c092 =  x153 &  x234 &  x262 &  x290 &  x658;
assign c094 =  x510 &  x652 & ~x580;
assign c096 =  x210 &  x319 &  x347 &  x375 &  x459 &  x515 &  x631 & ~x504;
assign c098 =  x291 &  x319 &  x354 &  x355 &  x383 &  x438 &  x514;
assign c0100 =  x327 &  x373 &  x383 &  x401 &  x428 &  x456 &  x512 & ~x369 & ~x580 & ~x582;
assign c0102 =  x400 &  x428 & ~x403 & ~x548 & ~x601;
assign c0104 =  x344 &  x372 &  x400 &  x412 &  x428 &  x440 &  x468 &  x513;
assign c0106 =  x210 &  x383 &  x430 &  x486 &  x514 &  x630 & ~x302 & ~x613 & ~x764;
assign c0108 =  x213 &  x373 &  x400 &  x412 &  x427 &  x626;
assign c0110 =  x778;
assign c0112 =  x727;
assign c0114 =  x321 &  x375 &  x437 &  x438 & ~x0 & ~x46 & ~x83 & ~x114 & ~x137 & ~x204 & ~x234 & ~x235 & ~x248 & ~x260 & ~x284 & ~x290 & ~x342 & ~x366 & ~x420 & ~x469 & ~x580 & ~x609 & ~x641 & ~x686 & ~x708;
assign c0116 = ~x326 & ~x374 & ~x382 & ~x521 & ~x574;
assign c0118 =  x373 &  x427 &  x454 &  x537;
assign c0120 =  x207 &  x234 &  x262 & ~x382 & ~x409 & ~x438;
assign c0122 =  x9;
assign c0124 =  x214 &  x357 &  x385 & ~x69 & ~x111 & ~x123 & ~x193 & ~x326 & ~x381 & ~x396;
assign c0126 =  x372 &  x400 &  x427 &  x455 &  x540 &  x568 &  x597 & ~x230 & ~x375 & ~x708;
assign c0128 =  x359 &  x481;
assign c0130 =  x82;
assign c0132 =  x213 &  x375 &  x485 & ~x373 & ~x580 & ~x604;
assign c0134 =  x370 &  x398;
assign c0136 =  x299 &  x370 &  x441;
assign c0138 =  x399 &  x427 &  x566 & ~x204 & ~x258 & ~x462 & ~x607 & ~x663 & ~x766;
assign c0140 =  x374 &  x401 &  x456 &  x484 &  x511 &  x626 & ~x38 & ~x396 & ~x679 & ~x725;
assign c0142 =  x214 &  x358 &  x386 & ~x22 & ~x71 & ~x163 & ~x281 & ~x449 & ~x507 & ~x707 & ~x748 & ~x780;
assign c0144 =  x262 &  x429 &  x468 &  x486 &  x496 & ~x506 & ~x511;
assign c0146 =  x356 &  x384 &  x412 &  x440 &  x485 &  x513 & ~x105 & ~x286 & ~x381 & ~x621 & ~x708;
assign c0148 =  x214 &  x327 &  x402 &  x542 & ~x525 & ~x532 & ~x660 & ~x712;
assign c0150 =  x427 &  x455 &  x511 &  x567 & ~x135 & ~x204 & ~x375 & ~x415 & ~x475 & ~x535 & ~x582;
assign c0152 =  x347 &  x375 &  x383 &  x431 &  x486 & ~x16 & ~x86 & ~x96 & ~x343 & ~x563;
assign c0154 =  x617;
assign c0156 =  x425 & ~x176 & ~x285 & ~x411 & ~x610;
assign c0158 =  x214 &  x373 &  x428 &  x456 &  x484 &  x512 &  x540 & ~x14 & ~x57 & ~x142 & ~x145 & ~x166 & ~x203 & ~x368 & ~x618 & ~x757;
assign c0160 =  x20 &  x339;
assign c0162 =  x558;
assign c0164 =  x217 &  x303;
assign c0166 =  x444;
assign c0168 =  x328 &  x383 &  x401 &  x429 &  x512 &  x540 & ~x497 & ~x580 & ~x768;
assign c0170 =  x184 &  x375 &  x402 &  x457 &  x485 &  x513 &  x655 & ~x234 & ~x260 & ~x469 & ~x551 & ~x724 & ~x752;
assign c0172 =  x342 & ~x380 & ~x411 & ~x757 & ~x765 & ~x770;
assign c0174 =  x372 & ~x374 & ~x601;
assign c0176 =  x212 &  x215 &  x272 &  x347 &  x625 & ~x263;
assign c0178 =  x214 &  x236 &  x327 &  x630 & ~x76 & ~x463 & ~x667 & ~x712 & ~x716;
assign c0180 =  x401 &  x428 &  x538 & ~x207;
assign c0182 =  x282;
assign c0184 =  x207 &  x234 &  x467 &  x632 &  x657 &  x658 & ~x108 & ~x176 & ~x417 & ~x452 & ~x684 & ~x706 & ~x752 & ~x778;
assign c0186 =  x357 &  x385 &  x413 &  x428 &  x441 & ~x409 & ~x463;
assign c0188 =  x415 & ~x120 & ~x123 & ~x202 & ~x408;
assign c0190 =  x239 &  x294 &  x297 &  x375 &  x430 &  x458 &  x486 & ~x525 & ~x710;
assign c0192 =  x657 &  x658 &  x659 & ~x27 & ~x293 & ~x322 & ~x378 & ~x433 & ~x451 & ~x548 & ~x575 & ~x641;
assign c0194 =  x370 &  x471 & ~x409;
assign c0196 =  x154 &  x290 &  x468 &  x629 & ~x259 & ~x470;
assign c0198 =  x746;
assign c0200 =  x297 &  x325 &  x353 &  x354 &  x382 &  x430 &  x486 &  x514 & ~x11 & ~x123 & ~x189 & ~x230 & ~x274 & ~x286 & ~x334 & ~x370 & ~x386;
assign c0202 =  x560;
assign c0204 =  x213 &  x413 & ~x494;
assign c0206 =  x330 &  x358 &  x386 & ~x313 & ~x326 & ~x437;
assign c0208 =  x157 &  x185 &  x237 & ~x6 & ~x33 & ~x98 & ~x110 & ~x123 & ~x161 & ~x203 & ~x229 & ~x234 & ~x259 & ~x274 & ~x339 & ~x453 & ~x469 & ~x498 & ~x582 & ~x584 & ~x607 & ~x618 & ~x632 & ~x641 & ~x660;
assign c0210 =  x383 &  x401 &  x411 &  x429 &  x456 &  x457 &  x512 & ~x386 & ~x469 & ~x647 & ~x710 & ~x715 & ~x737;
assign c0212 =  x298 &  x375 &  x410 &  x458 &  x459;
assign c0214 =  x373 &  x401 &  x429 &  x457 &  x485 &  x513 &  x628 &  x657 & ~x26 & ~x108 & ~x204 & ~x221 & ~x312 & ~x446 & ~x472 & ~x538 & ~x560 & ~x616 & ~x666 & ~x703 & ~x706;
assign c0216 =  x158 &  x215 &  x328 & ~x354;
assign c0218 =  x302 &  x413 & ~x411;
assign c0220 =  x85;
assign c0222 =  x360;
assign c0224 =  x216 &  x329 &  x357 &  x385 &  x413 &  x541;
assign c0226 =  x374 &  x429 &  x457 &  x512 &  x624 & ~x235 & ~x259 & ~x343 & ~x647;
assign c0228 =  x319 &  x375 &  x601 &  x603 & ~x712;
assign c0230 =  x359 & ~x354;
assign c0232 =  x213 &  x316 &  x371;
assign c0234 =  x429 &  x513 &  x632 &  x658 & ~x652;
assign c0236 =  x298 &  x370 &  x385 &  x413;
assign c0238 =  x153 &  x291 &  x319 &  x347 &  x402 &  x430 &  x458 &  x486 &  x630 &  x631;
assign c0240 =  x316 &  x471 & ~x601;
assign c0242 =  x292 &  x400 &  x455;
assign c0244 =  x185 &  x486 &  x493 &  x514 &  x598 & ~x64 & ~x217 & ~x364 & ~x517;
assign c0246 =  x206 &  x233 &  x299 &  x632 & ~x348 & ~x520 & ~x752;
assign c0248 =  x439 &  x656 &  x657 &  x658 & ~x409 & ~x573;
assign c0250 =  x386 &  x510 & ~x354;
assign c0252 =  x326 &  x382 &  x402 &  x430 &  x486 &  x514 &  x629 & ~x132 & ~x475 & ~x509 & ~x616;
assign c0254 =  x291 &  x319 &  x402 &  x430 &  x439 &  x458 & ~x330 & ~x408 & ~x464;
assign c0256 =  x344 &  x399 &  x427 &  x455 & ~x17 & ~x164 & ~x346 & ~x404 & ~x405 & ~x419 & ~x424 & ~x432 & ~x506 & ~x695 & ~x705 & ~x744;
assign c0258 =  x428 &  x456 &  x539 & ~x123 & ~x549;
assign c0260 =  x302 &  x454 & ~x123 & ~x381 & ~x487 & ~x632 & ~x639 & ~x670;
assign c0262 =  x302 & ~x382;
assign c0264 =  x315 &  x539;
assign c0266 =  x188 &  x328 &  x493;
assign c0268 =  x11;
assign c0270 =  x334 &  x676;
assign c0272 =  x251 &  x530;
assign c0274 =  x297 &  x325 &  x371 &  x399 &  x400 &  x413;
assign c0276 =  x416;
assign c0278 =  x275 &  x453 &  x509;
assign c0280 =  x186 &  x214 &  x357 &  x626 & ~x223 & ~x289 & ~x563;
assign c0282 =  x477;
assign c0284 =  x270 &  x299 &  x327 &  x355 &  x402 &  x430 &  x486 &  x514 & ~x40 & ~x203 & ~x706;
assign c0286 =  x400 &  x428 &  x456 &  x484 & ~x256 & ~x286 & ~x403 & ~x471 & ~x520 & ~x556 & ~x617 & ~x665 & ~x750;
assign c0288 =  x344 &  x385 &  x441 &  x469 &  x496;
assign c0290 =  x370 &  x443 & ~x381 & ~x409;
assign c0292 =  x359 &  x387 & ~x176;
assign c0294 =  x154 &  x262 &  x522 &  x630 &  x657 & ~x652;
assign c0296 =  x414 &  x442 & ~x75 & ~x120 & ~x134 & ~x173 & ~x389 & ~x439 & ~x506 & ~x587 & ~x648 & ~x705 & ~x759 & ~x768;
assign c0298 =  x154 &  x265 &  x493 &  x631 & ~x535;
assign c01 =  x324 &  x350 &  x352;
assign c03 =  x408;
assign c05 =  x491 &  x518 &  x521 &  x547 & ~x656;
assign c07 =  x713;
assign c09 = ~x14 & ~x100 & ~x108 & ~x115 & ~x134 & ~x141 & ~x155 & ~x156 & ~x160 & ~x473 & ~x477 & ~x529 & ~x569 & ~x570 & ~x571 & ~x596 & ~x597 & ~x598 & ~x613 & ~x614 & ~x620 & ~x624 & ~x626 & ~x627 & ~x653 & ~x779;
assign c011 =  x551 &  x552 &  x579 & ~x237 & ~x238 & ~x264;
assign c013 =  x300 & ~x155 & ~x158 & ~x512 & ~x543 & ~x570 & ~x610;
assign c015 = ~x157 & ~x181 & ~x183 & ~x184 & ~x185 & ~x281 & ~x378 & ~x450 & ~x513 & ~x540 & ~x541 & ~x542 & ~x552 & ~x569 & ~x677 & ~x698;
assign c017 =  x461 & ~x27 & ~x36 & ~x49 & ~x50 & ~x62 & ~x77 & ~x89 & ~x114 & ~x115 & ~x117 & ~x225 & ~x229 & ~x279 & ~x331 & ~x345 & ~x351 & ~x352 & ~x365 & ~x397 & ~x445 & ~x561 & ~x588 & ~x620 & ~x664 & ~x671 & ~x677 & ~x685 & ~x691 & ~x693 & ~x704 & ~x721 & ~x734 & ~x743 & ~x767;
assign c019 =  x288 & ~x153 & ~x154 & ~x155 & ~x156 & ~x539 & ~x542 & ~x568 & ~x571;
assign c021 =  x653 & ~x388 & ~x395 & ~x456 & ~x457 & ~x512 & ~x513 & ~x514 & ~x539;
assign c023 =  x518 &  x548 &  x578 & ~x387 & ~x657;
assign c025 = ~x240 & ~x319 & ~x626 & ~x627 & ~x628 & ~x629 & ~x653 & ~x656;
assign c027 =  x516 &  x518 & ~x29 & ~x61 & ~x91 & ~x100 & ~x122 & ~x217 & ~x253 & ~x303 & ~x351 & ~x406 & ~x588 & ~x590 & ~x591 & ~x656;
assign c029 =  x317 & ~x71 & ~x88 & ~x338 & ~x351 & ~x361 & ~x561 & ~x568 & ~x570 & ~x596 & ~x624 & ~x672 & ~x754 & ~x780;
assign c031 =  x380 & ~x518;
assign c033 =  x379 & ~x268 & ~x295;
assign c035 = ~x11 & ~x214 & ~x222 & ~x241 & ~x242 & ~x246 & ~x268 & ~x269 & ~x271 & ~x272 & ~x503 & ~x624 & ~x712;
assign c037 =  x460 &  x489 &  x490 & ~x4 & ~x40 & ~x85 & ~x119 & ~x129 & ~x166 & ~x281 & ~x504 & ~x556 & ~x571 & ~x588 & ~x742;
assign c039 =  x405 &  x406 & ~x412;
assign c041 =  x378 &  x379 & ~x517;
assign c043 =  x377 &  x606;
assign c045 =  x436 &  x463 &  x464 &  x490 &  x491 &  x492 &  x517 &  x518 &  x545 & ~x29 & ~x94 & ~x140 & ~x280 & ~x350 & ~x590 & ~x620 & ~x669 & ~x691 & ~x721 & ~x724;
assign c047 =  x349 &  x350 &  x351 & ~x687;
assign c049 = ~x64 & ~x96 & ~x184 & ~x185 & ~x212 & ~x213 & ~x214 & ~x387 & ~x512 & ~x514 & ~x542;
assign c051 =  x433 &  x434 &  x462 &  x520 & ~x27 & ~x41 & ~x49 & ~x77 & ~x93 & ~x109 & ~x114 & ~x188 & ~x193 & ~x229 & ~x340 & ~x363 & ~x393 & ~x394 & ~x415 & ~x557 & ~x618 & ~x679 & ~x744 & ~x748 & ~x751;
assign c053 = ~x143 & ~x183 & ~x194 & ~x544 & ~x570 & ~x571 & ~x598 & ~x617 & ~x653 & ~x754 & ~x757;
assign c055 =  x460 &  x461 &  x463 &  x464 & ~x73 & ~x122 & ~x129 & ~x219 & ~x249 & ~x280 & ~x417 & ~x691 & ~x696 & ~x699;
assign c057 = ~x14 & ~x39 & ~x128 & ~x140 & ~x157 & ~x351 & ~x476 & ~x570 & ~x571 & ~x572 & ~x598 & ~x600 & ~x620 & ~x627 & ~x628 & ~x653;
assign c059 =  x323 & ~x246 & ~x272 & ~x300 & ~x457 & ~x460;
assign c061 =  x460 &  x461 &  x462 &  x463 &  x464 & ~x323;
assign c063 =  x518 &  x576 & ~x299;
assign c065 =  x211 & ~x10 & ~x12 & ~x83 & ~x245 & ~x269 & ~x271 & ~x272 & ~x283 & ~x298 & ~x299 & ~x394 & ~x482 & ~x692 & ~x704 & ~x750;
assign c067 =  x351 &  x352 & ~x457;
assign c069 =  x378 & ~x267;
assign c071 = ~x156 & ~x166 & ~x415 & ~x541 & ~x542 & ~x543 & ~x569 & ~x570 & ~x571 & ~x598 & ~x626;
assign c073 =  x128 &  x545 & ~x346 & ~x347;
assign c075 =  x209 &  x376 &  x378 & ~x544;
assign c077 =  x462 &  x463 &  x492 & ~x106 & ~x294 & ~x295;
assign c079 = ~x160 & ~x213 & ~x215 & ~x240 & ~x242 & ~x265 & ~x655 & ~x656 & ~x657;
assign c081 =  x460 &  x461 &  x462 & ~x56 & ~x72 & ~x84 & ~x145 & ~x351 & ~x378 & ~x380 & ~x419 & ~x535 & ~x613 & ~x689 & ~x703 & ~x726 & ~x727 & ~x732 & ~x751;
assign c083 =  x551 &  x552 &  x578 & ~x212 & ~x238 & ~x240;
assign c085 =  x405 &  x406 &  x407;
assign c087 =  x266 & ~x181 & ~x183 & ~x184 & ~x185 & ~x413 & ~x482 & ~x514 & ~x537 & ~x540 & ~x588 & ~x615 & ~x620 & ~x634;
assign c089 =  x320 & ~x202 & ~x242 & ~x244 & ~x269 & ~x270 & ~x272 & ~x297 & ~x299 & ~x300 & ~x314 & ~x332 & ~x536 & ~x588;
assign c091 =  x241 &  x243 & ~x4 & ~x36 & ~x51 & ~x52 & ~x62 & ~x71 & ~x90 & ~x91 & ~x114 & ~x126 & ~x129 & ~x143 & ~x147 & ~x157 & ~x171 & ~x233 & ~x287 & ~x303 & ~x329 & ~x341 & ~x356 & ~x387 & ~x389 & ~x393 & ~x440 & ~x484 & ~x499 & ~x615 & ~x617 & ~x635 & ~x693 & ~x726 & ~x732;
assign c093 =  x627 &  x653 & ~x64 & ~x106 & ~x115 & ~x117 & ~x302 & ~x303 & ~x340 & ~x388 & ~x450 & ~x455 & ~x484 & ~x744;
assign c095 =  x460 &  x461 &  x462 & ~x121 & ~x147 & ~x170 & ~x232 & ~x350 & ~x475;
assign c097 =  x634 & ~x570 & ~x600;
assign c099 =  x192;
assign c0101 =  x460 &  x461 &  x462 &  x488 &  x489 & ~x71 & ~x93 & ~x200 & ~x287 & ~x707;
assign c0103 =  x211 & ~x244 & ~x269 & ~x297 & ~x299 & ~x300;
assign c0105 =  x637;
assign c0107 =  x349 &  x350 & ~x239 & ~x276;
assign c0109 =  x516 &  x517 &  x518 & ~x17 & ~x49 & ~x64 & ~x79 & ~x83 & ~x86 & ~x98 & ~x166 & ~x253 & ~x284 & ~x319 & ~x346 & ~x351 & ~x364 & ~x387 & ~x444 & ~x532 & ~x590 & ~x613 & ~x658 & ~x680 & ~x698 & ~x753 & ~x769;
assign c0111 =  x179 &  x182 &  x653;
assign c0113 =  x295 & ~x14 & ~x24 & ~x29 & ~x32 & ~x33 & ~x41 & ~x61 & ~x66 & ~x74 & ~x86 & ~x92 & ~x106 & ~x114 & ~x115 & ~x119 & ~x161 & ~x190 & ~x200 & ~x281 & ~x336 & ~x388 & ~x406 & ~x418 & ~x427 & ~x457 & ~x458 & ~x461 & ~x484 & ~x499 & ~x505 & ~x506 & ~x561 & ~x613 & ~x618 & ~x620 & ~x650 & ~x668 & ~x689 & ~x690 & ~x701 & ~x729 & ~x733 & ~x754 & ~x756 & ~x761;
assign c0115 =  x489 &  x490 &  x576 & ~x74 & ~x167 & ~x174 & ~x333 & ~x335 & ~x613 & ~x646 & ~x656 & ~x720 & ~x744 & ~x755;
assign c0117 =  x461 &  x489 &  x490 & ~x14 & ~x15 & ~x65 & ~x102 & ~x178 & ~x351 & ~x367 & ~x446 & ~x448 & ~x645 & ~x759 & ~x771;
assign c0119 =  x351 &  x352 & ~x229 & ~x245 & ~x265;
assign c0121 =  x490 & ~x7 & ~x71 & ~x80 & ~x94 & ~x114 & ~x143 & ~x165 & ~x201 & ~x226 & ~x268 & ~x269 & ~x283 & ~x342 & ~x393 & ~x414 & ~x445 & ~x450 & ~x471 & ~x474 & ~x613 & ~x615 & ~x620 & ~x669 & ~x694 & ~x738 & ~x749 & ~x768 & ~x770 & ~x783;
assign c0123 =  x323 & ~x237 & ~x264 & ~x458 & ~x783;
assign c0125 =  x517 &  x518 & ~x303 & ~x401 & ~x455 & ~x458 & ~x619 & ~x657 & ~x743;
assign c0127 =  x489 &  x490 &  x517 &  x518 &  x519 & ~x1 & ~x24 & ~x29 & ~x111 & ~x166 & ~x400 & ~x406 & ~x421 & ~x746;
assign c0129 =  x434 &  x435 &  x436 & ~x18 & ~x30 & ~x39 & ~x42 & ~x97 & ~x113 & ~x280 & ~x282 & ~x283 & ~x339 & ~x418 & ~x450 & ~x475 & ~x559 & ~x615 & ~x699 & ~x739 & ~x748;
assign c0131 =  x432 &  x433 &  x434 & ~x27 & ~x188;
assign c0133 = ~x155 & ~x157 & ~x364 & ~x486 & ~x539 & ~x569 & ~x570 & ~x571 & ~x572 & ~x598 & ~x626 & ~x653;
assign c0135 =  x436 & ~x89 & ~x246 & ~x656;
assign c0137 =  x716;
assign c0139 =  x405 &  x633;
assign c0141 = ~x214 & ~x241 & ~x242 & ~x268 & ~x270 & ~x271 & ~x272 & ~x656;
assign c0143 =  x689;
assign c0145 =  x577 & ~x158 & ~x211 & ~x214 & ~x242 & ~x505;
assign c0147 =  x264 & ~x128 & ~x155 & ~x157 & ~x206 & ~x349 & ~x388 & ~x542 & ~x569 & ~x570;
assign c0149 =  x684 &  x712 & ~x158;
assign c0151 =  x406 &  x407 &  x408;
assign c0153 =  x435 &  x436 & ~x268;
assign c0155 = ~x136 & ~x166 & ~x412 & ~x443 & ~x512 & ~x513 & ~x571;
assign c0157 =  x545 &  x574 & ~x87 & ~x166 & ~x191 & ~x270 & ~x271 & ~x450 & ~x655 & ~x656 & ~x708;
assign c0159 =  x324 &  x350 &  x351;
assign c0161 = ~x213 & ~x214 & ~x265 & ~x269;
assign c0163 =  x551 &  x578 & ~x28 & ~x136 & ~x366 & ~x592 & ~x625 & ~x626 & ~x628 & ~x629 & ~x655 & ~x656 & ~x657 & ~x658 & ~x693;
assign c0165 =  x491 &  x492 &  x518 &  x521 &  x545 &  x546 & ~x14 & ~x31 & ~x111 & ~x253 & ~x282 & ~x334 & ~x361 & ~x478 & ~x531 & ~x565 & ~x613 & ~x752;
assign c0167 =  x491 & ~x321 & ~x340 & ~x376 & ~x542 & ~x569;
assign c0169 =  x406 & ~x412;
assign c0171 =  x408 & ~x213;
assign c0173 =  x235 &  x464 &  x492 &  x518 &  x546 & ~x41 & ~x82 & ~x92 & ~x323 & ~x350 & ~x351 & ~x613;
assign c0175 =  x461 &  x462 & ~x43 & ~x283 & ~x297 & ~x530 & ~x612 & ~x741;
assign c0177 =  x350 & ~x328 & ~x359 & ~x461 & ~x514;
assign c0179 =  x407 &  x408 & ~x297;
assign c0181 = ~x214 & ~x242 & ~x268 & ~x274 & ~x299 & ~x656 & ~x657;
assign c0183 =  x576 & ~x80 & ~x160 & ~x163 & ~x213 & ~x214 & ~x239 & ~x240 & ~x242 & ~x266 & ~x656;
assign c0185 =  x408 & ~x22 & ~x73 & ~x133 & ~x405 & ~x431 & ~x456 & ~x458;
assign c0187 =  x350 &  x351 &  x352 & ~x34 & ~x195 & ~x287 & ~x435 & ~x461 & ~x697 & ~x728 & ~x781;
assign c0189 =  x211 &  x462 &  x463 &  x464 &  x465 &  x489 &  x490 & ~x49 & ~x107 & ~x118 & ~x172 & ~x231 & ~x360 & ~x714 & ~x718 & ~x724 & ~x750 & ~x759;
assign c0191 =  x176 & ~x38 & ~x72 & ~x104 & ~x114 & ~x199 & ~x248 & ~x264 & ~x277 & ~x427 & ~x617 & ~x620 & ~x743 & ~x748;
assign c0193 =  x408 & ~x324;
assign c0195 =  x517 & ~x240 & ~x270;
assign c0197 =  x689 & ~x151;
assign c0199 =  x377 &  x378 &  x379 &  x380;
assign c0201 =  x490 &  x518 &  x521;
assign c0203 =  x491 & ~x14 & ~x42 & ~x58 & ~x94 & ~x166 & ~x333 & ~x570 & ~x571 & ~x597 & ~x598 & ~x688 & ~x778;
assign c0205 =  x323 & ~x406 & ~x458 & ~x459;
assign c0207 =  x349 &  x350 & ~x459;
assign c0209 =  x407 & ~x269;
assign c0211 =  x407 &  x408 & ~x295;
assign c0213 =  x379 &  x380 & ~x268;
assign c0215 =  x351 &  x378 & ~x266;
assign c0217 =  x351 &  x377 & ~x329;
assign c0219 =  x433 &  x434 & ~x199 & ~x273 & ~x360 & ~x729;
assign c0221 =  x460 & ~x166 & ~x291 & ~x361 & ~x629 & ~x656;
assign c0223 =  x436 &  x548 & ~x10 & ~x27 & ~x38 & ~x167 & ~x198 & ~x284 & ~x306 & ~x350 & ~x534 & ~x563 & ~x643 & ~x656 & ~x701 & ~x749 & ~x754 & ~x773 & ~x775;
assign c0225 =  x211 &  x432 &  x433 &  x434 & ~x58 & ~x337;
assign c0227 =  x434 &  x435 & ~x325;
assign c0229 =  x464 &  x520 & ~x22 & ~x172 & ~x320 & ~x336 & ~x629 & ~x656 & ~x773;
assign c0231 =  x350 &  x351 &  x352 & ~x518 & ~x544;
assign c0233 = ~x106 & ~x128 & ~x156 & ~x157 & ~x158 & ~x183 & ~x184 & ~x185 & ~x186 & ~x352 & ~x406 & ~x416 & ~x484 & ~x495 & ~x512 & ~x514 & ~x620;
assign c0235 =  x462 &  x463 &  x548 & ~x31 & ~x83 & ~x92 & ~x140 & ~x339 & ~x351 & ~x613 & ~x616 & ~x698 & ~x767;
assign c0237 = ~x14 & ~x73 & ~x129 & ~x152 & ~x154 & ~x155 & ~x156 & ~x194 & ~x378 & ~x542 & ~x543 & ~x544 & ~x568 & ~x569 & ~x570 & ~x571 & ~x597 & ~x598 & ~x599 & ~x626;
assign c0239 =  x407 &  x434 & ~x118 & ~x139 & ~x217;
assign c0241 =  x491 &  x518 &  x551 & ~x475 & ~x656;
assign c0243 =  x516 &  x518 &  x574 & ~x475 & ~x658;
assign c0245 =  x263 &  x264 & ~x153 & ~x155 & ~x156 & ~x182 & ~x183 & ~x184 & ~x190 & ~x542 & ~x568 & ~x569 & ~x570;
assign c0247 =  x179 &  x653 & ~x428 & ~x515;
assign c0249 = ~x214 & ~x295 & ~x628 & ~x629 & ~x653 & ~x656;
assign c0251 =  x322 & ~x237 & ~x238 & ~x405 & ~x513 & ~x514 & ~x650 & ~x738;
assign c0253 =  x377 &  x379 & ~x544;
assign c0255 =  x574 & ~x2 & ~x90 & ~x128 & ~x131 & ~x155 & ~x182 & ~x183 & ~x184 & ~x512 & ~x543;
assign c0257 = ~x155 & ~x156 & ~x352 & ~x569 & ~x570 & ~x571 & ~x598 & ~x627;
assign c0259 = ~x185 & ~x186 & ~x213 & ~x214 & ~x238 & ~x239 & ~x412 & ~x495;
assign c0261 =  x408 & ~x246 & ~x268 & ~x279 & ~x295;
assign c0263 =  x350 &  x351 & ~x238 & ~x239;
assign c0265 = ~x128 & ~x184 & ~x185 & ~x188 & ~x212 & ~x213 & ~x214 & ~x215 & ~x484;
assign c0267 =  x378 &  x379 &  x380;
assign c0269 = ~x2 & ~x27 & ~x29 & ~x47 & ~x85 & ~x118 & ~x156 & ~x157 & ~x168 & ~x179 & ~x181 & ~x183 & ~x184 & ~x185 & ~x226 & ~x228 & ~x280 & ~x417 & ~x482 & ~x495 & ~x498 & ~x504 & ~x512 & ~x524 & ~x554 & ~x556 & ~x558 & ~x559 & ~x565 & ~x620 & ~x698 & ~x704 & ~x721 & ~x733 & ~x751 & ~x769;
assign c0271 =  x232 & ~x29 & ~x119 & ~x190 & ~x429 & ~x433 & ~x455 & ~x617 & ~x743;
assign c0273 = ~x5 & ~x29 & ~x32 & ~x36 & ~x71 & ~x87 & ~x114 & ~x166 & ~x195 & ~x239 & ~x264 & ~x265 & ~x281 & ~x330 & ~x340 & ~x371 & ~x391 & ~x398 & ~x421 & ~x457 & ~x476 & ~x527 & ~x557 & ~x560 & ~x699 & ~x732 & ~x755 & ~x759 & ~x771 & ~x779;
assign c0275 = ~x2 & ~x4 & ~x118 & ~x169 & ~x244 & ~x246 & ~x269 & ~x270 & ~x271 & ~x272 & ~x298 & ~x360 & ~x417 & ~x453 & ~x592 & ~x624 & ~x653 & ~x709;
assign c0277 =  x490 &  x518 & ~x106 & ~x121 & ~x240 & ~x266 & ~x295 & ~x370 & ~x376;
assign c0279 =  x435 & ~x38 & ~x45 & ~x247 & ~x656;
assign c0281 =  x578 & ~x378 & ~x629 & ~x656;
assign c0283 =  x523 &  x551 & ~x72 & ~x166 & ~x472 & ~x629 & ~x630 & ~x655 & ~x656 & ~x658;
assign c0285 =  x211 & ~x242 & ~x272 & ~x656;
assign c0287 =  x380 &  x434 & ~x153;
assign c0289 =  x434 & ~x205 & ~x232 & ~x272 & ~x555 & ~x748;
assign c0291 =  x349 &  x380;
assign c0293 =  x433 &  x434 &  x461;
assign c0295 =  x405 &  x406 & ~x272 & ~x685 & ~x734 & ~x747;
assign c0297 =  x430 &  x434 &  x435 &  x436 & ~x476 & ~x502;
assign c0299 = ~x183 & ~x184 & ~x361 & ~x513 & ~x569 & ~x570 & ~x598;
assign c10 =  x576 &  x577 &  x605 & ~x25 & ~x28 & ~x35 & ~x54 & ~x56 & ~x58 & ~x62 & ~x76 & ~x78 & ~x86 & ~x88 & ~x142 & ~x160 & ~x215 & ~x222 & ~x224 & ~x226 & ~x243 & ~x244 & ~x270 & ~x298 & ~x300 & ~x367 & ~x373 & ~x382 & ~x391 & ~x418 & ~x423 & ~x448 & ~x452 & ~x459 & ~x504 & ~x505 & ~x509 & ~x514 & ~x536 & ~x537 & ~x540 & ~x544 & ~x562 & ~x567 & ~x585 & ~x589 & ~x620 & ~x641 & ~x657 & ~x674 & ~x676 & ~x685 & ~x699 & ~x725 & ~x759 & ~x764 & ~x765 & ~x781;
assign c12 =  x435 &  x575 &  x576 & ~x12 & ~x34 & ~x59 & ~x73 & ~x104 & ~x140 & ~x142 & ~x149 & ~x202 & ~x214 & ~x230 & ~x243 & ~x244 & ~x246 & ~x248 & ~x270 & ~x298 & ~x354 & ~x366 & ~x382 & ~x390 & ~x404 & ~x423 & ~x427 & ~x439 & ~x459 & ~x487 & ~x527 & ~x588 & ~x620 & ~x652 & ~x655 & ~x686 & ~x718 & ~x722 & ~x750;
assign c14 =  x266 &  x267 &  x293 &  x464 &  x575 &  x576 &  x604 & ~x93 & ~x113 & ~x146 & ~x149 & ~x150 & ~x159 & ~x160 & ~x214 & ~x223 & ~x225 & ~x229 & ~x247 & ~x270 & ~x280 & ~x298 & ~x299 & ~x336 & ~x357 & ~x365 & ~x370 & ~x469 & ~x537 & ~x568 & ~x587 & ~x619 & ~x621 & ~x678 & ~x681 & ~x706 & ~x718 & ~x778;
assign c16 =  x72;
assign c18 =  x196;
assign c110 =  x378 & ~x104 & ~x204 & ~x214 & ~x240 & ~x243 & ~x245 & ~x298 & ~x459 & ~x469 & ~x542 & ~x565 & ~x620 & ~x623 & ~x731 & ~x738 & ~x775;
assign c112 =  x186 &  x297 &  x377 &  x432 &  x571 & ~x8 & ~x17 & ~x26 & ~x62 & ~x65 & ~x180 & ~x193 & ~x287 & ~x400 & ~x416 & ~x440 & ~x499 & ~x508 & ~x526 & ~x552 & ~x639 & ~x696 & ~x731 & ~x768;
assign c114 =  x16;
assign c116 =  x544 &  x571 & ~x103 & ~x154 & ~x209 & ~x238 & ~x357 & ~x375 & ~x403 & ~x443 & ~x620 & ~x737;
assign c118 =  x72;
assign c120 =  x154 &  x155 & ~x110 & ~x148 & ~x169 & ~x187 & ~x214 & ~x242 & ~x298 & ~x301 & ~x326 & ~x390 & ~x404 & ~x438 & ~x451 & ~x454 & ~x486 & ~x487 & ~x515 & ~x668 & ~x677 & ~x727 & ~x773 & ~x776 & ~x783;
assign c124 =  x381 &  x432 & ~x211;
assign c126 =  x351 & ~x6 & ~x67 & ~x113 & ~x121 & ~x167 & ~x170 & ~x230 & ~x243 & ~x257 & ~x271 & ~x298 & ~x325 & ~x336 & ~x404 & ~x405 & ~x431 & ~x444 & ~x448 & ~x475 & ~x503 & ~x645 & ~x646 & ~x659 & ~x688 & ~x689 & ~x717 & ~x729 & ~x741;
assign c128 =  x86;
assign c130 =  x72;
assign c132 =  x241 &  x324 &  x379 &  x461 & ~x209 & ~x210 & ~x238 & ~x239 & ~x603 & ~x631 & ~x735;
assign c134 =  x186 &  x571 & ~x55 & ~x183 & ~x237 & ~x523 & ~x629 & ~x731;
assign c136 =  x520 &  x576 & ~x0 & ~x1 & ~x7 & ~x23 & ~x28 & ~x55 & ~x59 & ~x68 & ~x77 & ~x78 & ~x79 & ~x86 & ~x102 & ~x158 & ~x163 & ~x168 & ~x170 & ~x190 & ~x197 & ~x198 & ~x213 & ~x214 & ~x243 & ~x246 & ~x248 & ~x253 & ~x269 & ~x284 & ~x298 & ~x313 & ~x335 & ~x357 & ~x358 & ~x362 & ~x369 & ~x388 & ~x389 & ~x416 & ~x418 & ~x419 & ~x421 & ~x425 & ~x441 & ~x444 & ~x455 & ~x458 & ~x503 & ~x515 & ~x527 & ~x528 & ~x539 & ~x553 & ~x567 & ~x585 & ~x588 & ~x596 & ~x617 & ~x642 & ~x650 & ~x652 & ~x654 & ~x673 & ~x676 & ~x679 & ~x693 & ~x710 & ~x711 & ~x716 & ~x719 & ~x731 & ~x736 & ~x737 & ~x738 & ~x740 & ~x758 & ~x766 & ~x781;
assign c138 =  x85;
assign c140 =  x110;
assign c142 =  x433 & ~x23 & ~x59 & ~x138 & ~x214 & ~x243 & ~x281 & ~x289 & ~x296 & ~x298 & ~x324 & ~x325 & ~x326 & ~x352 & ~x380 & ~x514 & ~x623 & ~x728 & ~x774;
assign c144 =  x238 &  x295 &  x351 &  x378 &  x462 & ~x39 & ~x62 & ~x64 & ~x90 & ~x104 & ~x106 & ~x113 & ~x114 & ~x180 & ~x227 & ~x299 & ~x303 & ~x357 & ~x358 & ~x371 & ~x372 & ~x398 & ~x420 & ~x426 & ~x437 & ~x451 & ~x456 & ~x466 & ~x469 & ~x480 & ~x483 & ~x511 & ~x527 & ~x588 & ~x637 & ~x638 & ~x670 & ~x716 & ~x727 & ~x742 & ~x745 & ~x746 & ~x752;
assign c146 =  x295 &  x296 &  x323 &  x351 & ~x38 & ~x39 & ~x64 & ~x77 & ~x86 & ~x87 & ~x108 & ~x170 & ~x208 & ~x209 & ~x247 & ~x251 & ~x265 & ~x272 & ~x273 & ~x285 & ~x337 & ~x390 & ~x448 & ~x466 & ~x468 & ~x480 & ~x492 & ~x509 & ~x541 & ~x612 & ~x619 & ~x649 & ~x702 & ~x710 & ~x728 & ~x740 & ~x771 & ~x773 & ~x775;
assign c148 =  x649;
assign c150 =  x324 &  x461 &  x518 &  x519 &  x573 &  x574 & ~x147 & ~x163 & ~x232 & ~x343 & ~x421 & ~x500 & ~x523 & ~x626 & ~x682;
assign c152 =  x761;
assign c154 =  x323 &  x519 &  x545 &  x573 & ~x15 & ~x22 & ~x54 & ~x58 & ~x69 & ~x85 & ~x90 & ~x95 & ~x120 & ~x197 & ~x214 & ~x215 & ~x216 & ~x232 & ~x242 & ~x243 & ~x270 & ~x298 & ~x313 & ~x337 & ~x392 & ~x410 & ~x412 & ~x424 & ~x442 & ~x470 & ~x477 & ~x541 & ~x553 & ~x581 & ~x583 & ~x621 & ~x623 & ~x644 & ~x651 & ~x654 & ~x665 & ~x712 & ~x730 & ~x731 & ~x734 & ~x762 & ~x766 & ~x772 & ~x775 & ~x776 & ~x781;
assign c156 =  x161 &  x408 & ~x209 & ~x520;
assign c158 =  x460 & ~x209 & ~x212 & ~x239 & ~x600;
assign c160 = ~x30 & ~x48 & ~x107 & ~x113 & ~x214 & ~x225 & ~x243 & ~x258 & ~x270 & ~x271 & ~x308 & ~x316 & ~x340 & ~x352 & ~x361 & ~x380 & ~x408 & ~x452 & ~x485 & ~x512 & ~x554 & ~x556 & ~x565 & ~x626 & ~x638 & ~x705 & ~x740 & ~x755;
assign c162 =  x291 &  x521 &  x606 & ~x277 & ~x298 & ~x472 & ~x709;
assign c164 =  x297 & ~x107 & ~x152 & ~x156 & ~x179 & ~x183 & ~x209 & ~x211 & ~x347 & ~x348 & ~x357 & ~x577 & ~x629;
assign c166 =  x308;
assign c168 =  x184 &  x295 &  x324 &  x377 &  x461 &  x489 &  x545 &  x571 &  x600 & ~x32 & ~x39 & ~x59 & ~x63 & ~x76 & ~x140 & ~x145 & ~x152 & ~x175 & ~x200 & ~x207 & ~x221 & ~x253 & ~x417 & ~x428 & ~x448 & ~x457 & ~x513 & ~x554 & ~x595 & ~x623 & ~x680 & ~x681 & ~x743 & ~x750 & ~x780;
assign c170 = ~x70 & ~x79 & ~x170 & ~x175 & ~x214 & ~x215 & ~x233 & ~x241 & ~x242 & ~x273 & ~x275 & ~x288 & ~x289 & ~x298 & ~x387 & ~x402 & ~x427 & ~x440 & ~x444 & ~x487 & ~x510 & ~x515 & ~x523 & ~x528 & ~x529 & ~x553 & ~x583 & ~x671 & ~x677 & ~x716 & ~x737 & ~x742;
assign c174 =  x486 &  x624 &  x652 & ~x179 & ~x207 & ~x209;
assign c176 =  x489 & ~x209 & ~x210 & ~x514 & ~x568;
assign c178 =  x158 &  x270 &  x571 & ~x209 & ~x236;
assign c180 =  x405 & ~x53 & ~x134 & ~x135 & ~x145 & ~x242 & ~x243 & ~x271 & ~x287 & ~x298 & ~x312 & ~x325 & ~x346 & ~x380 & ~x397 & ~x487 & ~x497 & ~x514 & ~x532 & ~x556 & ~x562 & ~x582 & ~x587 & ~x651 & ~x710 & ~x730 & ~x761 & ~x767;
assign c182 = ~x214 & ~x228 & ~x243 & ~x289 & ~x298 & ~x308 & ~x315 & ~x340 & ~x380 & ~x393 & ~x421 & ~x436 & ~x439 & ~x494 & ~x495 & ~x506 & ~x640 & ~x717 & ~x737;
assign c184 =  x291 &  x577 & ~x49 & ~x104 & ~x137 & ~x160 & ~x161 & ~x213 & ~x214 & ~x246 & ~x256 & ~x270 & ~x298 & ~x362 & ~x393 & ~x554 & ~x563 & ~x565;
assign c188 =  x214 &  x242 &  x270 &  x571 & ~x180;
assign c190 =  x239 &  x267 &  x322 & ~x29 & ~x42 & ~x48 & ~x51 & ~x54 & ~x82 & ~x89 & ~x102 & ~x116 & ~x131 & ~x142 & ~x197 & ~x201 & ~x208 & ~x246 & ~x264 & ~x271 & ~x283 & ~x286 & ~x300 & ~x335 & ~x364 & ~x371 & ~x382 & ~x392 & ~x399 & ~x412 & ~x428 & ~x438 & ~x449 & ~x468 & ~x473 & ~x480 & ~x535 & ~x537 & ~x550 & ~x588 & ~x642 & ~x648 & ~x650 & ~x667 & ~x671 & ~x674 & ~x711 & ~x716 & ~x718 & ~x727 & ~x752 & ~x755 & ~x761 & ~x771;
assign c192 = ~x152 & ~x209 & ~x212 & ~x239 & ~x376 & ~x521 & ~x631 & ~x760;
assign c194 =  x155 &  x294 &  x547 & ~x62 & ~x147 & ~x214 & ~x216 & ~x243 & ~x259 & ~x298 & ~x456 & ~x558 & ~x607 & ~x638;
assign c196 =  x298 &  x460 & ~x28 & ~x38 & ~x147 & ~x207 & ~x209 & ~x211 & ~x266 & ~x293 & ~x375 & ~x521 & ~x600 & ~x605 & ~x628 & ~x638 & ~x716;
assign c198 =  x267 &  x294 &  x351 &  x378 &  x407 &  x545 &  x573 &  x601 &  x602 & ~x8 & ~x23 & ~x25 & ~x30 & ~x32 & ~x33 & ~x39 & ~x40 & ~x43 & ~x66 & ~x69 & ~x70 & ~x76 & ~x79 & ~x95 & ~x99 & ~x107 & ~x112 & ~x118 & ~x140 & ~x147 & ~x161 & ~x170 & ~x177 & ~x191 & ~x197 & ~x198 & ~x199 & ~x222 & ~x229 & ~x232 & ~x249 & ~x253 & ~x256 & ~x257 & ~x272 & ~x275 & ~x289 & ~x301 & ~x303 & ~x308 & ~x312 & ~x328 & ~x336 & ~x341 & ~x344 & ~x358 & ~x359 & ~x362 & ~x363 & ~x365 & ~x389 & ~x390 & ~x400 & ~x421 & ~x423 & ~x425 & ~x428 & ~x448 & ~x449 & ~x455 & ~x456 & ~x469 & ~x494 & ~x497 & ~x537 & ~x552 & ~x557 & ~x559 & ~x562 & ~x563 & ~x582 & ~x617 & ~x619 & ~x641 & ~x645 & ~x651 & ~x653 & ~x664 & ~x666 & ~x668 & ~x677 & ~x678 & ~x682 & ~x695 & ~x698 & ~x705 & ~x708 & ~x718 & ~x730 & ~x735 & ~x740 & ~x750 & ~x751 & ~x760 & ~x764 & ~x768 & ~x771 & ~x773 & ~x775 & ~x776 & ~x778 & ~x780 & ~x783;
assign c1100 =  x90;
assign c1102 =  x320 &  x519 &  x576 & ~x39 & ~x105 & ~x160 & ~x161 & ~x241 & ~x298 & ~x325 & ~x459 & ~x480 & ~x487 & ~x511;
assign c1106 =  x445;
assign c1108 =  x189 &  x651 & ~x237;
assign c1110 =  x616;
assign c1112 =  x571 &  x653 & ~x209 & ~x375;
assign c1114 =  x210 &  x238 &  x294 &  x351 &  x461 &  x575 & ~x20 & ~x55 & ~x59 & ~x95 & ~x164 & ~x233 & ~x243 & ~x261 & ~x287 & ~x298 & ~x312 & ~x372 & ~x416 & ~x424 & ~x439 & ~x449 & ~x453 & ~x458 & ~x473 & ~x484 & ~x498 & ~x523 & ~x526 & ~x594 & ~x640 & ~x641 & ~x712 & ~x773 & ~x774;
assign c1116 = ~x86 & ~x105 & ~x170 & ~x198 & ~x214 & ~x243 & ~x273 & ~x298 & ~x325 & ~x326 & ~x403 & ~x432 & ~x439 & ~x459 & ~x487 & ~x513 & ~x514 & ~x515 & ~x587 & ~x612 & ~x619 & ~x686 & ~x716 & ~x739 & ~x774;
assign c1118 =  x379 &  x544 & ~x1 & ~x26 & ~x32 & ~x62 & ~x73 & ~x111 & ~x113 & ~x179 & ~x180 & ~x200 & ~x209 & ~x229 & ~x232 & ~x234 & ~x265 & ~x279 & ~x301 & ~x312 & ~x318 & ~x326 & ~x329 & ~x355 & ~x382 & ~x430 & ~x436 & ~x492 & ~x547 & ~x588 & ~x638 & ~x688 & ~x742 & ~x750;
assign c1122 =  x623 & ~x209 & ~x211 & ~x293;
assign c1124 =  x568 &  x596 &  x623 & ~x183 & ~x372 & ~x600 & ~x631;
assign c1126 =  x155 &  x238 &  x267 & ~x15 & ~x31 & ~x47 & ~x71 & ~x86 & ~x102 & ~x105 & ~x119 & ~x142 & ~x158 & ~x163 & ~x171 & ~x177 & ~x188 & ~x193 & ~x214 & ~x247 & ~x248 & ~x284 & ~x285 & ~x298 & ~x336 & ~x370 & ~x383 & ~x416 & ~x421 & ~x443 & ~x468 & ~x500 & ~x525 & ~x539 & ~x563 & ~x585 & ~x588 & ~x651 & ~x653 & ~x681 & ~x682 & ~x699 & ~x713 & ~x716 & ~x739 & ~x760 & ~x769 & ~x780;
assign c1128 =  x695;
assign c1130 =  x585;
assign c1132 =  x139;
assign c1134 =  x189 & ~x184 & ~x212 & ~x574;
assign c1136 =  x112 &  x783;
assign c1138 =  x293 &  x321 & ~x43 & ~x77 & ~x84 & ~x185 & ~x214 & ~x232 & ~x242 & ~x243 & ~x244 & ~x254 & ~x271 & ~x283 & ~x288 & ~x298 & ~x337 & ~x382 & ~x393 & ~x410 & ~x414 & ~x476 & ~x482 & ~x532 & ~x544 & ~x600 & ~x619 & ~x624 & ~x626 & ~x627 & ~x628 & ~x649 & ~x656 & ~x681 & ~x693 & ~x720 & ~x736 & ~x759 & ~x767;
assign c1140 =  x617;
assign c1142 =  x139;
assign c1144 =  x722;
assign c1146 =  x155 &  x209 &  x239 &  x294 &  x547 & ~x214 & ~x243 & ~x298 & ~x303 & ~x456 & ~x609;
assign c1148 = ~x27 & ~x121 & ~x209 & ~x243 & ~x259 & ~x285 & ~x298 & ~x431 & ~x442 & ~x468 & ~x472 & ~x492 & ~x519 & ~x541;
assign c1150 =  x561;
assign c1152 =  x239 &  x295 &  x461 &  x515 &  x544 &  x571 & ~x58 & ~x85 & ~x87 & ~x94 & ~x95 & ~x178 & ~x191 & ~x235 & ~x247 & ~x288 & ~x310 & ~x438 & ~x520 & ~x638 & ~x726;
assign c1154 =  x239 & ~x126 & ~x179 & ~x209 & ~x403 & ~x492 & ~x554 & ~x568 & ~x576;
assign c1156 =  x532;
assign c1158 =  x773;
assign c1160 =  x69;
assign c1162 =  x239 &  x351 & ~x8 & ~x16 & ~x49 & ~x56 & ~x79 & ~x104 & ~x107 & ~x160 & ~x165 & ~x217 & ~x247 & ~x298 & ~x357 & ~x382 & ~x386 & ~x397 & ~x400 & ~x404 & ~x405 & ~x421 & ~x449 & ~x460 & ~x514 & ~x527 & ~x534 & ~x537 & ~x560 & ~x620 & ~x644 & ~x663 & ~x755 & ~x764 & ~x773;
assign c1166 =  x108;
assign c1168 =  x189 & ~x628;
assign c1170 =  x16;
assign c1172 =  x728;
assign c1174 =  x83;
assign c1176 =  x266 &  x294 & ~x0 & ~x87 & ~x147 & ~x187 & ~x213 & ~x214 & ~x215 & ~x244 & ~x325 & ~x342 & ~x384 & ~x404 & ~x411 & ~x432 & ~x471 & ~x476 & ~x480 & ~x643 & ~x754;
assign c1178 =  x63;
assign c1180 =  x702;
assign c1182 =  x488 & ~x82 & ~x127 & ~x152 & ~x209 & ~x243 & ~x298 & ~x341 & ~x347 & ~x390 & ~x437 & ~x505 & ~x577 & ~x681;
assign c1184 =  x238 &  x294 &  x518 &  x574 & ~x0 & ~x31 & ~x49 & ~x63 & ~x67 & ~x77 & ~x94 & ~x99 & ~x113 & ~x140 & ~x172 & ~x177 & ~x190 & ~x214 & ~x215 & ~x242 & ~x243 & ~x246 & ~x254 & ~x270 & ~x288 & ~x298 & ~x300 & ~x307 & ~x308 & ~x326 & ~x328 & ~x355 & ~x365 & ~x414 & ~x420 & ~x425 & ~x439 & ~x458 & ~x467 & ~x515 & ~x523 & ~x527 & ~x535 & ~x542 & ~x570 & ~x651 & ~x666 & ~x685 & ~x718 & ~x736 & ~x754;
assign c1186 =  x548 &  x604 & ~x0 & ~x13 & ~x28 & ~x45 & ~x130 & ~x145 & ~x167 & ~x214 & ~x242 & ~x243 & ~x259 & ~x270 & ~x275 & ~x298 & ~x307 & ~x339 & ~x356 & ~x449 & ~x451 & ~x456 & ~x513 & ~x515 & ~x532 & ~x558 & ~x582 & ~x626 & ~x639 & ~x641 & ~x648 & ~x666 & ~x695 & ~x716 & ~x751 & ~x760 & ~x764;
assign c1188 =  x238 &  x267 &  x545 &  x546 &  x600 & ~x106 & ~x142 & ~x178 & ~x205 & ~x246 & ~x484 & ~x512 & ~x522 & ~x619 & ~x638 & ~x661 & ~x698;
assign c1190 =  x239 &  x323 &  x461 &  x518 &  x545 &  x546 & ~x12 & ~x15 & ~x45 & ~x60 & ~x66 & ~x86 & ~x105 & ~x124 & ~x137 & ~x149 & ~x162 & ~x177 & ~x200 & ~x205 & ~x232 & ~x243 & ~x270 & ~x298 & ~x300 & ~x328 & ~x339 & ~x372 & ~x383 & ~x394 & ~x396 & ~x419 & ~x430 & ~x443 & ~x448 & ~x450 & ~x469 & ~x474 & ~x481 & ~x505 & ~x514 & ~x556 & ~x587 & ~x613 & ~x614 & ~x651 & ~x652 & ~x653 & ~x673 & ~x675 & ~x698 & ~x722 & ~x773;
assign c1192 =  x625 &  x652 & ~x209 & ~x602 & ~x656;
assign c1194 =  x781;
assign c1196 =  x297 & ~x9 & ~x62 & ~x94 & ~x117 & ~x118 & ~x180 & ~x209 & ~x211 & ~x238 & ~x247 & ~x251 & ~x266 & ~x289 & ~x314 & ~x347 & ~x395 & ~x439 & ~x499 & ~x521 & ~x547 & ~x559 & ~x574 & ~x577 & ~x584 & ~x631 & ~x667 & ~x748 & ~x770 & ~x780;
assign c1198 =  x211 &  x239 &  x267 &  x294 &  x323 &  x461 &  x489 & ~x18 & ~x51 & ~x61 & ~x62 & ~x77 & ~x111 & ~x132 & ~x149 & ~x161 & ~x169 & ~x190 & ~x214 & ~x221 & ~x243 & ~x257 & ~x270 & ~x271 & ~x283 & ~x298 & ~x327 & ~x358 & ~x362 & ~x368 & ~x369 & ~x416 & ~x418 & ~x500 & ~x507 & ~x532 & ~x568 & ~x588 & ~x612 & ~x690 & ~x698 & ~x705 & ~x708 & ~x716 & ~x731 & ~x778;
assign c1200 =  x239 &  x240 &  x296 &  x323 &  x571 &  x573 &  x600 &  x656 & ~x178 & ~x180 & ~x219 & ~x346 & ~x526 & ~x535 & ~x608;
assign c1202 =  x568 &  x594;
assign c1204 =  x641;
assign c1206 =  x350 & ~x2 & ~x3 & ~x4 & ~x12 & ~x39 & ~x40 & ~x42 & ~x47 & ~x62 & ~x67 & ~x70 & ~x78 & ~x88 & ~x92 & ~x93 & ~x97 & ~x102 & ~x142 & ~x145 & ~x150 & ~x152 & ~x162 & ~x177 & ~x178 & ~x193 & ~x197 & ~x208 & ~x209 & ~x218 & ~x235 & ~x246 & ~x252 & ~x253 & ~x264 & ~x275 & ~x287 & ~x291 & ~x292 & ~x306 & ~x319 & ~x346 & ~x385 & ~x391 & ~x401 & ~x420 & ~x426 & ~x427 & ~x428 & ~x446 & ~x453 & ~x468 & ~x471 & ~x492 & ~x494 & ~x498 & ~x507 & ~x511 & ~x512 & ~x519 & ~x521 & ~x522 & ~x575 & ~x581 & ~x590 & ~x591 & ~x603 & ~x613 & ~x631 & ~x651 & ~x664 & ~x665 & ~x672 & ~x678 & ~x680 & ~x703 & ~x718 & ~x741 & ~x771 & ~x776 & ~x781;
assign c1208 =  x154 &  x546 &  x574 & ~x28 & ~x38 & ~x91 & ~x139 & ~x145 & ~x174 & ~x193 & ~x213 & ~x214 & ~x244 & ~x252 & ~x298 & ~x311 & ~x427 & ~x486 & ~x487 & ~x497 & ~x501 & ~x513 & ~x536 & ~x538 & ~x563 & ~x719 & ~x725 & ~x740 & ~x781;
assign c1210 =  x321 & ~x193 & ~x213 & ~x214 & ~x242 & ~x243 & ~x298 & ~x325 & ~x352 & ~x380 & ~x414 & ~x439 & ~x588 & ~x747;
assign c1212 =  x22;
assign c1214 =  x561;
assign c1216 =  x351 &  x461 &  x518 & ~x56 & ~x81 & ~x107 & ~x108 & ~x178 & ~x209 & ~x293 & ~x372 & ~x389 & ~x492 & ~x575 & ~x639;
assign c1218 =  x545 & ~x243 & ~x256 & ~x298 & ~x319 & ~x325 & ~x408 & ~x577;
assign c1220 =  x591;
assign c1224 =  x463 &  x575 & ~x27 & ~x29 & ~x31 & ~x50 & ~x132 & ~x133 & ~x160 & ~x161 & ~x163 & ~x171 & ~x191 & ~x202 & ~x214 & ~x243 & ~x246 & ~x257 & ~x298 & ~x371 & ~x386 & ~x404 & ~x414 & ~x439 & ~x459 & ~x484 & ~x522 & ~x561 & ~x638 & ~x689 & ~x699 & ~x705 & ~x736 & ~x768;
assign c1226 =  x242 &  x324 &  x353 &  x570 & ~x7 & ~x124 & ~x153 & ~x154 & ~x193 & ~x223 & ~x236 & ~x283 & ~x338 & ~x357 & ~x368 & ~x537 & ~x730 & ~x750;
assign c1228 =  x294 &  x324 &  x460 &  x546 &  x571 &  x573 & ~x372 & ~x457 & ~x500;
assign c1230 =  x253;
assign c1232 =  x449;
assign c1234 =  x16;
assign c1236 =  x157 &  x408 &  x571 &  x600 & ~x148 & ~x512;
assign c1238 =  x32;
assign c1240 =  x239 &  x350 &  x600 & ~x113 & ~x243 & ~x247 & ~x464;
assign c1242 =  x621 & ~x209;
assign c1244 =  x48;
assign c1246 =  x367;
assign c1248 =  x574 & ~x18 & ~x32 & ~x58 & ~x214 & ~x245 & ~x297 & ~x326 & ~x404 & ~x443 & ~x654;
assign c1250 =  x590;
assign c1252 =  x267 &  x295 &  x323 &  x353 &  x571 & ~x50 & ~x152 & ~x219 & ~x301 & ~x357 & ~x780;
assign c1254 =  x362;
assign c1256 =  x136;
assign c1258 =  x12;
assign c1262 =  x520 &  x633 & ~x59 & ~x68 & ~x99 & ~x107 & ~x163 & ~x168 & ~x176 & ~x197 & ~x213 & ~x214 & ~x245 & ~x246 & ~x284 & ~x285 & ~x327 & ~x332 & ~x382 & ~x444 & ~x487 & ~x500 & ~x563 & ~x649 & ~x695 & ~x716;
assign c1264 =  x293 &  x350 &  x519 & ~x23 & ~x113 & ~x134 & ~x143 & ~x212 & ~x213 & ~x286 & ~x298 & ~x390 & ~x403 & ~x439 & ~x459 & ~x565 & ~x623 & ~x654 & ~x681 & ~x720 & ~x723;
assign c1266 =  x242 &  x381 & ~x209 & ~x210 & ~x211;
assign c1268 =  x159 & ~x403 & ~x603;
assign c1270 =  x154 &  x182 &  x266 &  x518 & ~x26 & ~x31 & ~x54 & ~x59 & ~x66 & ~x107 & ~x114 & ~x120 & ~x170 & ~x214 & ~x230 & ~x243 & ~x259 & ~x283 & ~x298 & ~x326 & ~x358 & ~x365 & ~x368 & ~x369 & ~x390 & ~x425 & ~x479 & ~x509 & ~x552 & ~x553 & ~x582 & ~x612 & ~x640 & ~x645 & ~x655 & ~x713 & ~x727 & ~x745 & ~x765;
assign c1272 =  x450;
assign c1274 =  x533;
assign c1276 =  x766;
assign c1278 =  x339;
assign c1280 =  x266 &  x294 &  x377 &  x462 &  x518 & ~x14 & ~x27 & ~x54 & ~x62 & ~x63 & ~x82 & ~x86 & ~x92 & ~x147 & ~x161 & ~x164 & ~x213 & ~x214 & ~x217 & ~x242 & ~x243 & ~x247 & ~x249 & ~x251 & ~x273 & ~x285 & ~x298 & ~x313 & ~x328 & ~x357 & ~x358 & ~x362 & ~x392 & ~x421 & ~x422 & ~x486 & ~x487 & ~x500 & ~x528 & ~x538 & ~x541 & ~x568 & ~x611 & ~x617 & ~x623 & ~x638 & ~x644 & ~x651 & ~x668 & ~x669 & ~x682 & ~x692 & ~x698 & ~x707 & ~x708 & ~x728 & ~x731 & ~x762 & ~x768 & ~x773 & ~x775;
assign c1282 =  x160 &  x297 &  x353;
assign c1284 =  x464 &  x576 &  x605 &  x606 & ~x25 & ~x147 & ~x170 & ~x193 & ~x245 & ~x417 & ~x459 & ~x461 & ~x504 & ~x764 & ~x778;
assign c1286 = ~x0 & ~x27 & ~x61 & ~x113 & ~x119 & ~x129 & ~x142 & ~x147 & ~x159 & ~x183 & ~x184 & ~x211 & ~x212 & ~x213 & ~x222 & ~x239 & ~x366 & ~x375 & ~x402 & ~x427 & ~x448 & ~x527 & ~x555 & ~x590 & ~x600 & ~x627 & ~x628 & ~x629 & ~x655 & ~x656 & ~x692 & ~x698 & ~x724 & ~x756 & ~x759 & ~x765 & ~x773 & ~x774;
assign c1288 =  x270 &  x297 &  x324 & ~x178 & ~x184 & ~x207 & ~x209 & ~x211 & ~x239 & ~x397 & ~x439 & ~x603 & ~x629 & ~x631 & ~x632;
assign c1290 =  x167;
assign c1292 = ~x213 & ~x270 & ~x352 & ~x355 & ~x429 & ~x487 & ~x600;
assign c1294 =  x405 & ~x213 & ~x214 & ~x325 & ~x352 & ~x459 & ~x542;
assign c1296 =  x291 &  x464 &  x491 &  x577 &  x606 & ~x6 & ~x28 & ~x39 & ~x46 & ~x106 & ~x111 & ~x130 & ~x138 & ~x192 & ~x199 & ~x200 & ~x256 & ~x273 & ~x301 & ~x311 & ~x328 & ~x412 & ~x417 & ~x449 & ~x475 & ~x511 & ~x515 & ~x527 & ~x532 & ~x535 & ~x563 & ~x587 & ~x644 & ~x668 & ~x671 & ~x676 & ~x694 & ~x699 & ~x709 & ~x711 & ~x728 & ~x731 & ~x738 & ~x740 & ~x742 & ~x746 & ~x750 & ~x773;
assign c1298 =  x324 & ~x183 & ~x184 & ~x212 & ~x239 & ~x521 & ~x600 & ~x742;
assign c11 =  x468;
assign c13 =  x317 & ~x523 & ~x524 & ~x597;
assign c15 =  x376 &  x465 & ~x462;
assign c17 =  x465 & ~x545 & ~x661;
assign c19 =  x468;
assign c111 =  x459 & ~x3 & ~x7 & ~x23 & ~x63 & ~x76 & ~x81 & ~x97 & ~x116 & ~x138 & ~x162 & ~x165 & ~x170 & ~x171 & ~x175 & ~x223 & ~x233 & ~x249 & ~x259 & ~x302 & ~x315 & ~x354 & ~x355 & ~x382 & ~x389 & ~x391 & ~x409 & ~x410 & ~x442 & ~x447 & ~x502 & ~x507 & ~x527 & ~x529 & ~x538 & ~x539 & ~x558 & ~x564 & ~x613 & ~x641 & ~x650 & ~x665 & ~x667 & ~x672 & ~x673 & ~x702 & ~x706 & ~x712 & ~x723 & ~x740 & ~x746 & ~x750 & ~x780;
assign c113 =  x375 &  x377 & ~x154 & ~x199 & ~x232 & ~x257 & ~x353 & ~x363 & ~x419 & ~x428 & ~x530 & ~x580 & ~x638 & ~x686 & ~x693 & ~x701 & ~x755;
assign c115 =  x374 &  x402;
assign c117 =  x521 &  x549 & ~x30 & ~x75 & ~x233 & ~x235 & ~x289 & ~x291 & ~x316 & ~x610;
assign c119 =  x235 &  x686;
assign c121 =  x207 &  x234 &  x352 & ~x349;
assign c123 =  x177 &  x632;
assign c125 =  x246 &  x293 & ~x558;
assign c127 =  x403 & ~x349;
assign c129 =  x461 &  x580;
assign c131 =  x207 & ~x17 & ~x30 & ~x102 & ~x109 & ~x267 & ~x294 & ~x307 & ~x471;
assign c133 =  x287;
assign c135 =  x487 &  x549 & ~x71 & ~x105 & ~x260 & ~x276 & ~x293 & ~x374 & ~x391 & ~x618 & ~x659;
assign c137 =  x511;
assign c139 =  x354 &  x355 & ~x161 & ~x309 & ~x693;
assign c141 =  x427;
assign c143 =  x150 &  x151 &  x152;
assign c145 =  x521 & ~x490 & ~x677;
assign c147 =  x152 &  x579 & ~x99;
assign c149 =  x205 & ~x72 & ~x167 & ~x173 & ~x199 & ~x504 & ~x524 & ~x723;
assign c151 =  x347 &  x375 & ~x295 & ~x636;
assign c153 =  x412;
assign c155 =  x319 &  x347 &  x404 & ~x120 & ~x151 & ~x422 & ~x449 & ~x537 & ~x754;
assign c157 =  x178 & ~x519;
assign c159 =  x273 & ~x95 & ~x282;
assign c161 =  x236 &  x380 &  x435 & ~x15 & ~x164 & ~x191 & ~x251 & ~x295 & ~x306 & ~x538 & ~x584 & ~x702;
assign c163 =  x236 & ~x15 & ~x86 & ~x93 & ~x105 & ~x115 & ~x174 & ~x194 & ~x295 & ~x308 & ~x412 & ~x413 & ~x509 & ~x580 & ~x610 & ~x632 & ~x722 & ~x749 & ~x782;
assign c165 =  x244 & ~x5 & ~x15 & ~x18 & ~x40 & ~x81 & ~x200 & ~x226 & ~x268 & ~x281 & ~x288 & ~x310 & ~x341 & ~x362 & ~x365 & ~x423 & ~x525 & ~x688 & ~x694 & ~x773;
assign c167 =  x347 &  x404 & ~x81 & ~x141 & ~x155 & ~x302 & ~x532 & ~x609 & ~x691 & ~x745 & ~x747 & ~x755;
assign c169 =  x488 &  x550 & ~x76 & ~x107 & ~x161 & ~x255 & ~x262 & ~x293 & ~x358 & ~x384 & ~x528 & ~x529 & ~x538 & ~x593 & ~x609 & ~x613 & ~x680 & ~x706 & ~x712 & ~x771;
assign c171 =  x233 & ~x736;
assign c173 =  x271 & ~x49 & ~x95 & ~x106 & ~x148 & ~x219 & ~x235 & ~x277 & ~x295 & ~x367 & ~x374 & ~x390 & ~x472 & ~x505 & ~x507 & ~x552 & ~x579 & ~x608 & ~x613 & ~x765;
assign c175 =  x685 & ~x350;
assign c177 =  x328 & ~x460;
assign c179 =  x350 & ~x295 & ~x323 & ~x330;
assign c181 =  x245 & ~x55 & ~x397 & ~x484;
assign c183 =  x461 &  x599 & ~x36 & ~x69 & ~x99 & ~x221 & ~x225 & ~x226 & ~x229 & ~x286 & ~x304 & ~x351 & ~x474 & ~x578 & ~x585 & ~x614 & ~x677 & ~x684 & ~x712 & ~x744;
assign c185 =  x148;
assign c187 =  x436 & ~x8 & ~x20 & ~x32 & ~x63 & ~x64 & ~x78 & ~x119 & ~x161 & ~x257 & ~x282 & ~x304 & ~x350 & ~x356 & ~x359 & ~x371 & ~x420 & ~x471 & ~x577 & ~x610 & ~x615 & ~x646 & ~x651 & ~x746 & ~x748 & ~x777;
assign c189 =  x264 &  x683 &  x684 & ~x73 & ~x230 & ~x444 & ~x507 & ~x538 & ~x616 & ~x637 & ~x669 & ~x724;
assign c191 =  x458;
assign c193 = ~x378 & ~x379 & ~x606 & ~x634;
assign c195 =  x375 & ~x350;
assign c197 =  x374 & ~x267;
assign c199 =  x260;
assign c1101 =  x121;
assign c1103 =  x319 &  x347 &  x348 &  x376 & ~x322;
assign c1105 =  x510;
assign c1107 =  x319 & ~x25 & ~x61 & ~x86 & ~x205 & ~x276 & ~x496 & ~x544 & ~x550 & ~x572 & ~x619 & ~x632 & ~x649 & ~x707;
assign c1109 =  x411;
assign c1111 =  x409 & ~x463;
assign c1113 =  x129 &  x540 &  x567;
assign c1117 =  x660 &  x687;
assign c1119 =  x203;
assign c1121 =  x289 & ~x101 & ~x624;
assign c1123 =  x711;
assign c1125 =  x204;
assign c1127 =  x150 &  x151 & ~x320 & ~x383;
assign c1129 =  x237 & ~x349 & ~x350 & ~x391 & ~x428 & ~x529;
assign c1131 =  x497;
assign c1133 =  x437 &  x438 & ~x260 & ~x498 & ~x635;
assign c1135 =  x429 &  x461 & ~x147 & ~x162;
assign c1137 =  x510;
assign c1139 =  x537;
assign c1141 =  x374 &  x402 &  x403;
assign c1143 = ~x350 & ~x351 & ~x602 & ~x631;
assign c1145 =  x657 &  x658 & ~x164 & ~x220 & ~x282 & ~x410 & ~x448 & ~x472 & ~x578 & ~x634 & ~x732;
assign c1147 =  x153 &  x378 & ~x490;
assign c1149 =  x521 & ~x490;
assign c1151 =  x436 & ~x102 & ~x219 & ~x351 & ~x390 & ~x441 & ~x443 & ~x727 & ~x733 & ~x738;
assign c1153 =  x399;
assign c1155 =  x318 &  x319 & ~x8 & ~x226 & ~x444 & ~x578 & ~x635;
assign c1157 =  x410;
assign c1159 =  x510;
assign c1161 =  x467;
assign c1163 = ~x102 & ~x129 & ~x176 & ~x220 & ~x226 & ~x249 & ~x261 & ~x349 & ~x350 & ~x363 & ~x378 & ~x717 & ~x719 & ~x751 & ~x755;
assign c1165 =  x511;
assign c1167 =  x186 &  x434 &  x626 & ~x24 & ~x64 & ~x114 & ~x145 & ~x225 & ~x288 & ~x338 & ~x366 & ~x426 & ~x467 & ~x474 & ~x511 & ~x517 & ~x544 & ~x674 & ~x702 & ~x706 & ~x723 & ~x732 & ~x754 & ~x764;
assign c1169 =  x382 &  x383;
assign c1171 =  x317 & ~x342;
assign c1173 =  x238 &  x245 & ~x7 & ~x26 & ~x34 & ~x168 & ~x199 & ~x505 & ~x697;
assign c1175 =  x215 & ~x19 & ~x67 & ~x151 & ~x203 & ~x232 & ~x261 & ~x307 & ~x323 & ~x401 & ~x418 & ~x454 & ~x606 & ~x618 & ~x638 & ~x649 & ~x774;
assign c1177 =  x157 &  x459 & ~x20 & ~x192 & ~x200 & ~x371 & ~x373 & ~x389 & ~x399 & ~x443 & ~x448 & ~x476 & ~x508 & ~x538 & ~x545 & ~x671 & ~x679 & ~x694 & ~x719 & ~x724;
assign c1179 =  x235 &  x686;
assign c1181 =  x465 &  x466;
assign c1183 =  x710;
assign c1185 =  x151 &  x152;
assign c1187 =  x211 &  x409 & ~x495 & ~x533 & ~x571 & ~x575 & ~x608 & ~x670;
assign c1189 =  x655 & ~x47 & ~x75 & ~x138 & ~x142 & ~x147 & ~x161 & ~x177 & ~x229 & ~x268 & ~x358 & ~x421 & ~x428 & ~x445 & ~x551 & ~x558 & ~x619 & ~x632 & ~x637 & ~x687 & ~x692 & ~x694 & ~x730;
assign c1191 =  x402 & ~x44 & ~x193 & ~x362 & ~x471 & ~x586 & ~x589 & ~x604 & ~x611 & ~x636 & ~x756;
assign c1193 =  x234 & ~x122 & ~x282 & ~x320 & ~x339 & ~x615 & ~x634;
assign c1195 =  x495;
assign c1197 =  x235 &  x712;
assign c1199 =  x686 &  x687 & ~x128 & ~x623;
assign c1201 =  x549 & ~x41 & ~x55 & ~x121 & ~x166 & ~x225 & ~x290 & ~x336 & ~x363 & ~x397 & ~x446 & ~x450 & ~x475 & ~x481 & ~x490 & ~x497 & ~x505 & ~x608 & ~x732 & ~x779;
assign c1203 =  x300 &  x301;
assign c1205 =  x521 & ~x323;
assign c1207 =  x346 &  x374;
assign c1209 =  x206 & ~x88 & ~x349;
assign c1211 =  x348 &  x404 & ~x36 & ~x457 & ~x517 & ~x564 & ~x621 & ~x635 & ~x688 & ~x694;
assign c1213 =  x439;
assign c1215 =  x152 &  x580 & ~x102 & ~x114;
assign c1217 =  x274;
assign c1219 =  x207 &  x379 &  x517 & ~x31 & ~x65 & ~x113 & ~x167 & ~x196 & ~x247 & ~x332 & ~x347 & ~x349 & ~x457 & ~x506 & ~x510 & ~x595 & ~x610;
assign c1221 =  x466;
assign c1223 =  x315;
assign c1225 =  x402 &  x403 &  x404 & ~x458 & ~x502 & ~x555 & ~x605;
assign c1227 =  x345 & ~x80;
assign c1229 =  x458 & ~x137 & ~x144 & ~x262 & ~x298 & ~x424 & ~x450 & ~x585 & ~x645 & ~x653 & ~x730;
assign c1231 =  x598 &  x628 &  x658 & ~x10 & ~x17 & ~x19 & ~x38 & ~x41 & ~x43 & ~x57 & ~x58 & ~x80 & ~x87 & ~x134 & ~x163 & ~x164 & ~x178 & ~x191 & ~x197 & ~x202 & ~x221 & ~x229 & ~x247 & ~x257 & ~x312 & ~x343 & ~x365 & ~x393 & ~x414 & ~x446 & ~x455 & ~x526 & ~x537 & ~x572 & ~x613 & ~x669 & ~x701 & ~x705 & ~x710 & ~x718 & ~x720 & ~x759 & ~x767;
assign c1233 = ~x295 & ~x545 & ~x550 & ~x726;
assign c1235 =  x430 & ~x9 & ~x15 & ~x18 & ~x28 & ~x54 & ~x60 & ~x67 & ~x72 & ~x109 & ~x169 & ~x312 & ~x325 & ~x368 & ~x386 & ~x418 & ~x424 & ~x477 & ~x479 & ~x500 & ~x557 & ~x698 & ~x703 & ~x709 & ~x733 & ~x745 & ~x762 & ~x771;
assign c1237 =  x494 & ~x278 & ~x290 & ~x481;
assign c1239 =  x207 &  x325 & ~x17 & ~x21 & ~x65 & ~x86 & ~x114 & ~x193 & ~x230 & ~x287 & ~x293 & ~x308 & ~x366 & ~x367 & ~x375 & ~x474 & ~x510 & ~x512 & ~x557 & ~x587 & ~x668 & ~x671 & ~x700 & ~x704 & ~x738 & ~x745 & ~x752 & ~x754 & ~x768 & ~x772 & ~x781;
assign c1241 =  x437 & ~x490 & ~x719;
assign c1243 =  x404 & ~x350;
assign c1245 =  x237 &  x244 &  x298 & ~x136 & ~x588 & ~x613 & ~x725 & ~x746;
assign c1247 =  x234 & ~x65 & ~x222 & ~x291 & ~x308 & ~x349 & ~x368 & ~x370 & ~x507 & ~x747;
assign c1249 =  x494;
assign c1251 =  x409 & ~x434;
assign c1253 =  x301;
assign c1255 =  x457;
assign c1257 =  x150 &  x151 &  x152 & ~x669;
assign c1259 =  x150 &  x151 &  x152;
assign c1261 =  x289 & ~x128 & ~x147 & ~x199 & ~x663;
assign c1263 =  x511 &  x539;
assign c1265 =  x459 &  x549 & ~x43 & ~x705;
assign c1267 = ~x236 & ~x378 & ~x379;
assign c1269 = ~x406 & ~x407 & ~x505;
assign c1271 =  x375;
assign c1273 =  x236 & ~x48 & ~x72 & ~x171 & ~x332 & ~x349 & ~x367 & ~x467 & ~x571 & ~x595;
assign c1275 =  x437 & ~x579;
assign c1277 =  x182 &  x209 &  x658 &  x685;
assign c1279 =  x399;
assign c1281 =  x459 &  x521 & ~x25 & ~x29 & ~x108 & ~x135 & ~x392 & ~x423 & ~x665 & ~x729 & ~x754 & ~x773;
assign c1283 =  x157 &  x354 & ~x295 & ~x477 & ~x594;
assign c1285 =  x234 &  x269 & ~x125 & ~x148 & ~x163 & ~x361 & ~x468 & ~x473 & ~x506 & ~x568 & ~x635 & ~x700 & ~x704 & ~x767;
assign c1287 =  x459 & ~x123 & ~x131 & ~x176 & ~x221 & ~x323 & ~x696 & ~x732 & ~x756 & ~x774;
assign c1289 =  x628 & ~x434 & ~x435 & ~x462;
assign c1291 =  x514 &  x580;
assign c1293 =  x234 & ~x560 & ~x569 & ~x606;
assign c1295 =  x550 & ~x170 & ~x334 & ~x583 & ~x635 & ~x730 & ~x753;
assign c1297 = ~x350 & ~x351 & ~x575 & ~x635;
assign c1299 = ~x189 & ~x377 & ~x378 & ~x379;
assign c20 =  x180 &  x488 &  x515 &  x626 & ~x91 & ~x106 & ~x315 & ~x368 & ~x493 & ~x710;
assign c22 =  x528;
assign c24 =  x460 & ~x409 & ~x490 & ~x492 & ~x493;
assign c26 =  x431 &  x512 & ~x266 & ~x301 & ~x313 & ~x334;
assign c28 =  x613;
assign c210 =  x59;
assign c212 =  x500;
assign c214 =  x761;
assign c216 =  x65;
assign c218 =  x207 &  x516 &  x543 & ~x383 & ~x494 & ~x521 & ~x619;
assign c220 =  x155 &  x156 & ~x19 & ~x51 & ~x239 & ~x352 & ~x369 & ~x506 & ~x685 & ~x711;
assign c222 =  x667;
assign c224 =  x464 &  x488 &  x537;
assign c226 =  x477;
assign c228 =  x584;
assign c230 =  x88;
assign c232 =  x527 & ~x601;
assign c234 =  x153 &  x297 & ~x289 & ~x409 & ~x412 & ~x465 & ~x492 & ~x667;
assign c236 =  x296 &  x514 &  x542 & ~x215 & ~x299;
assign c238 =  x501;
assign c240 = ~x39 & ~x45 & ~x132 & ~x214 & ~x299 & ~x327 & ~x366 & ~x575 & ~x601 & ~x602 & ~x604 & ~x607 & ~x628 & ~x629 & ~x657 & ~x689 & ~x694 & ~x720 & ~x737 & ~x779;
assign c242 =  x294 & ~x154 & ~x213 & ~x326 & ~x354 & ~x631;
assign c244 =  x634 &  x635 & ~x66 & ~x96 & ~x275 & ~x301 & ~x346 & ~x356 & ~x373 & ~x448 & ~x584;
assign c246 =  x209 &  x298 &  x326 &  x599 &  x600 &  x602 & ~x8 & ~x56 & ~x112 & ~x276 & ~x301 & ~x333 & ~x420 & ~x424 & ~x482 & ~x504 & ~x645 & ~x721 & ~x748 & ~x757 & ~x759;
assign c248 =  x30;
assign c250 =  x390;
assign c252 =  x521 &  x554 & ~x443;
assign c254 =  x528;
assign c256 =  x353 &  x381 &  x491 &  x545 & ~x383 & ~x630 & ~x657;
assign c258 =  x464 &  x482 & ~x5 & ~x59 & ~x78 & ~x121 & ~x143 & ~x147 & ~x195 & ~x229 & ~x288 & ~x340 & ~x601 & ~x631 & ~x635 & ~x644 & ~x684 & ~x717 & ~x724;
assign c260 =  x122 & ~x319 & ~x497;
assign c262 =  x7;
assign c264 =  x517 &  x576 &  x604 &  x626 & ~x768;
assign c266 =  x122 & ~x206 & ~x350;
assign c268 =  x465 &  x537 & ~x325;
assign c270 =  x531;
assign c272 =  x486 &  x570 & ~x292 & ~x301 & ~x384;
assign c274 =  x530;
assign c276 =  x127 &  x485 & ~x428;
assign c278 =  x584;
assign c280 =  x432 &  x485 & ~x382 & ~x579 & ~x602 & ~x628 & ~x689;
assign c282 =  x432 &  x467 &  x469 & ~x381;
assign c284 =  x403 &  x483 & ~x135 & ~x266 & ~x283 & ~x294 & ~x314 & ~x681 & ~x778;
assign c286 =  x153 &  x327 & ~x10 & ~x25 & ~x31 & ~x34 & ~x36 & ~x294 & ~x352 & ~x365 & ~x380 & ~x390 & ~x472 & ~x726 & ~x740;
assign c288 =  x297 &  x488 &  x515 &  x605 & ~x426 & ~x438 & ~x492;
assign c290 =  x526 & ~x604 & ~x658;
assign c292 =  x488 &  x515 &  x629 &  x630 & ~x81 & ~x292 & ~x373 & ~x494;
assign c294 =  x583;
assign c296 =  x56;
assign c298 =  x151 &  x153 &  x326 & ~x187 & ~x216 & ~x351 & ~x441;
assign c2100 =  x536;
assign c2102 =  x581 & ~x469 & ~x498;
assign c2104 =  x354 &  x491 &  x518 &  x569 & ~x351;
assign c2106 =  x155 &  x431 &  x457;
assign c2108 =  x473;
assign c2110 =  x390;
assign c2112 =  x472 & ~x604;
assign c2114 =  x465 &  x537 & ~x324 & ~x352;
assign c2116 =  x156 &  x353 &  x381 &  x436 &  x518 &  x545 & ~x6 & ~x34 & ~x73 & ~x80 & ~x118 & ~x120 & ~x172 & ~x332 & ~x360 & ~x391 & ~x424 & ~x495 & ~x645 & ~x678 & ~x702 & ~x709 & ~x716;
assign c2118 =  x184 &  x436 &  x463 &  x518 &  x545 &  x569 &  x597 & ~x412 & ~x658;
assign c2120 =  x355 &  x546 &  x600 & ~x310 & ~x352 & ~x380 & ~x428;
assign c2122 =  x182 &  x209 &  x210 &  x516 &  x517 &  x543 &  x571 & ~x75 & ~x128 & ~x193 & ~x275 & ~x306 & ~x308 & ~x309 & ~x335 & ~x360 & ~x374 & ~x385 & ~x402 & ~x642 & ~x700 & ~x726 & ~x736 & ~x749;
assign c2124 =  x532;
assign c2126 =  x336;
assign c2128 =  x472 &  x493;
assign c2130 = ~x274 & ~x299 & ~x326 & ~x601 & ~x603 & ~x631;
assign c2132 =  x459 &  x577 & ~x371 & ~x399 & ~x409 & ~x683;
assign c2134 =  x641;
assign c2136 =  x127 &  x128 & ~x211 & ~x237 & ~x239 & ~x295 & ~x344 & ~x656;
assign c2138 =  x543 &  x605 &  x624;
assign c2140 =  x526 & ~x180;
assign c2142 =  x29;
assign c2144 =  x12;
assign c2146 =  x472;
assign c2148 =  x484 &  x539 & ~x103;
assign c2150 =  x483 & ~x574 & ~x600;
assign c2152 =  x268 &  x601 &  x605 & ~x314 & ~x409 & ~x437;
assign c2154 =  x404 &  x429 &  x483 & ~x40 & ~x64 & ~x133 & ~x192 & ~x231 & ~x281 & ~x739;
assign c2156 =  x755;
assign c2158 =  x157 &  x158 &  x515 & ~x37 & ~x295 & ~x349 & ~x375 & ~x401 & ~x403;
assign c2160 =  x26;
assign c2162 =  x283;
assign c2164 =  x184 &  x299 &  x327 &  x355 &  x463 & ~x324 & ~x352 & ~x684 & ~x771;
assign c2166 =  x46;
assign c2168 =  x151 &  x152 & ~x157 & ~x221 & ~x236 & ~x245 & ~x370 & ~x481 & ~x563 & ~x580 & ~x617;
assign c2170 =  x599 &  x600 &  x634 & ~x59 & ~x278 & ~x308 & ~x321 & ~x403 & ~x430 & ~x528 & ~x670;
assign c2172 =  x446;
assign c2174 =  x297 &  x353 &  x381 &  x436 &  x491 &  x518 &  x546 &  x573 &  x600 & ~x39 & ~x63 & ~x93 & ~x132 & ~x159 & ~x190 & ~x216 & ~x248 & ~x251 & ~x275 & ~x391 & ~x503 & ~x723 & ~x736;
assign c2176 =  x576 &  x578 & ~x275 & ~x429 & ~x438 & ~x493 & ~x761;
assign c2178 =  x155 &  x158 &  x460 &  x567 & ~x292;
assign c2180 =  x546 &  x606 & ~x430 & ~x483;
assign c2182 =  x584;
assign c2184 =  x511 & ~x111 & ~x136 & ~x143 & ~x200 & ~x205 & ~x256 & ~x276 & ~x304 & ~x601 & ~x602 & ~x628 & ~x672 & ~x688 & ~x722;
assign c2186 =  x154 &  x184 &  x516 & ~x3 & ~x5 & ~x8 & ~x9 & ~x11 & ~x28 & ~x48 & ~x49 & ~x52 & ~x60 & ~x61 & ~x88 & ~x90 & ~x102 & ~x103 & ~x104 & ~x110 & ~x136 & ~x140 & ~x143 & ~x163 & ~x165 & ~x198 & ~x224 & ~x253 & ~x256 & ~x257 & ~x276 & ~x306 & ~x310 & ~x313 & ~x367 & ~x372 & ~x376 & ~x387 & ~x391 & ~x397 & ~x403 & ~x419 & ~x445 & ~x452 & ~x456 & ~x457 & ~x470 & ~x471 & ~x473 & ~x477 & ~x480 & ~x506 & ~x527 & ~x557 & ~x643 & ~x669 & ~x726 & ~x727 & ~x742 & ~x743 & ~x745 & ~x749 & ~x752 & ~x759 & ~x776;
assign c2188 =  x155 &  x184 &  x326 &  x353 &  x381 &  x491 &  x546 &  x599 & ~x245 & ~x301;
assign c2190 =  x210 &  x516 &  x629 & ~x403 & ~x521;
assign c2192 =  x43 &  x670;
assign c2194 =  x153 &  x154 &  x212 &  x268 & ~x77 & ~x81 & ~x104 & ~x145 & ~x159 & ~x166 & ~x174 & ~x189 & ~x196 & ~x245 & ~x250 & ~x252 & ~x275 & ~x321 & ~x330 & ~x364 & ~x367 & ~x444 & ~x450 & ~x483 & ~x501 & ~x560 & ~x620 & ~x674 & ~x700 & ~x701 & ~x722 & ~x751;
assign c2196 =  x179 &  x180 &  x208 & ~x185 & ~x214 & ~x373 & ~x711 & ~x713;
assign c2198 =  x726;
assign c2200 =  x266 &  x473;
assign c2202 =  x488 &  x489 &  x491 &  x518 &  x519 & ~x28 & ~x107 & ~x120 & ~x133 & ~x223 & ~x602 & ~x628 & ~x629 & ~x631 & ~x656 & ~x714 & ~x738 & ~x771;
assign c2204 =  x184 &  x212 &  x464 &  x597 & ~x323 & ~x379;
assign c2206 =  x268 &  x487 &  x514 &  x541 &  x542;
assign c2208 =  x527 & ~x633;
assign c2210 =  x355 &  x463 &  x566 & ~x656 & ~x684;
assign c2212 =  x459 &  x510 & ~x657;
assign c2214 =  x155 &  x353 &  x489 &  x516 &  x543 & ~x70 & ~x113 & ~x383 & ~x430 & ~x449 & ~x493 & ~x494 & ~x529;
assign c2216 =  x389;
assign c2218 =  x520 &  x547 &  x600 &  x626 & ~x276 & ~x352 & ~x380 & ~x427;
assign c2220 =  x156 &  x457 & ~x235 & ~x320 & ~x321 & ~x346;
assign c2222 =  x124 & ~x353 & ~x409 & ~x414;
assign c2224 =  x120;
assign c2226 =  x554;
assign c2228 =  x210 &  x353 &  x489 &  x517 &  x571 & ~x58 & ~x245 & ~x254 & ~x328;
assign c2230 =  x431 &  x457 &  x484 &  x512 & ~x318;
assign c2232 =  x153 &  x493 &  x547 & ~x32 & ~x352;
assign c2234 =  x634 & ~x383 & ~x413 & ~x494 & ~x578;
assign c2236 =  x609 & ~x456 & ~x496;
assign c2238 =  x328 &  x438 &  x567 & ~x352;
assign c2240 =  x263 & ~x181 & ~x382 & ~x602;
assign c2242 = ~x29 & ~x126 & ~x183 & ~x185 & ~x187 & ~x199 & ~x212 & ~x214 & ~x215 & ~x242 & ~x246 & ~x249 & ~x272 & ~x298 & ~x299 & ~x326 & ~x354 & ~x447 & ~x530 & ~x656 & ~x660 & ~x748 & ~x755;
assign c2244 =  x581 & ~x259;
assign c2248 =  x128 &  x129 &  x158 &  x186 & ~x39 & ~x136 & ~x211 & ~x310 & ~x657;
assign c2250 =  x458 &  x484 &  x511 & ~x385 & ~x586 & ~x681 & ~x682 & ~x691 & ~x722 & ~x731;
assign c2252 =  x460 & ~x181 & ~x383 & ~x575 & ~x629 & ~x655 & ~x660;
assign c2254 =  x93;
assign c2256 =  x617;
assign c2258 =  x432 &  x512 & ~x601 & ~x628 & ~x629;
assign c2260 =  x158 &  x159 &  x244 & ~x18 & ~x116 & ~x172 & ~x223 & ~x251 & ~x286 & ~x324 & ~x387 & ~x584 & ~x586 & ~x706 & ~x723 & ~x751;
assign c2262 =  x136;
assign c2264 =  x63;
assign c2266 =  x156 &  x465 &  x520 & ~x324 & ~x352;
assign c2268 =  x24;
assign c2270 =  x296 & ~x242 & ~x438;
assign c2272 =  x473;
assign c2274 =  x463 &  x536;
assign c2276 =  x501;
assign c2278 =  x389;
assign c2280 =  x520 &  x553 & ~x644 & ~x662;
assign c2282 = ~x214 & ~x297 & ~x299 & ~x354 & ~x381 & ~x601 & ~x602 & ~x608 & ~x632;
assign c2284 =  x336;
assign c2286 =  x97;
assign c2288 =  x125 & ~x354 & ~x409;
assign c2290 =  x408 &  x546 & ~x185 & ~x245 & ~x271 & ~x354 & ~x455;
assign c2292 =  x640;
assign c2294 =  x490 &  x493 & ~x356 & ~x438 & ~x602 & ~x632 & ~x660;
assign c2296 =  x179 &  x487 & ~x409 & ~x464 & ~x491;
assign c21 =  x318 &  x346 &  x374 &  x402 & ~x38 & ~x41 & ~x84 & ~x199 & ~x201 & ~x278 & ~x323 & ~x341 & ~x423 & ~x453 & ~x502 & ~x528 & ~x565 & ~x666 & ~x671 & ~x696 & ~x723 & ~x735 & ~x760;
assign c23 =  x219;
assign c25 =  x379 &  x380 & ~x55 & ~x115 & ~x308 & ~x313 & ~x358 & ~x399 & ~x453 & ~x503 & ~x513 & ~x515 & ~x543 & ~x614 & ~x646 & ~x667 & ~x691 & ~x693 & ~x745 & ~x748 & ~x768 & ~x783;
assign c27 =  x323 &  x350 & ~x333 & ~x487 & ~x488 & ~x489 & ~x704;
assign c29 =  x185 &  x407 &  x434 &  x435 &  x655 & ~x124 & ~x145 & ~x168 & ~x497 & ~x664;
assign c211 = ~x13 & ~x33 & ~x162 & ~x251 & ~x309 & ~x487 & ~x488 & ~x489 & ~x514 & ~x517 & ~x518 & ~x546 & ~x547 & ~x589 & ~x748;
assign c213 =  x378 &  x379 &  x407 & ~x6 & ~x8 & ~x11 & ~x19 & ~x26 & ~x28 & ~x44 & ~x49 & ~x50 & ~x52 & ~x62 & ~x86 & ~x99 & ~x111 & ~x121 & ~x124 & ~x137 & ~x150 & ~x166 & ~x176 & ~x196 & ~x198 & ~x230 & ~x260 & ~x276 & ~x278 & ~x334 & ~x428 & ~x453 & ~x498 & ~x500 & ~x524 & ~x557 & ~x579 & ~x585 & ~x642 & ~x662 & ~x692 & ~x705 & ~x750 & ~x755 & ~x761 & ~x774 & ~x779;
assign c215 = ~x23 & ~x33 & ~x110 & ~x134 & ~x142 & ~x147 & ~x158 & ~x160 & ~x162 & ~x168 & ~x175 & ~x186 & ~x217 & ~x222 & ~x240 & ~x241 & ~x258 & ~x260 & ~x270 & ~x285 & ~x287 & ~x307 & ~x341 & ~x417 & ~x447 & ~x564 & ~x585 & ~x589 & ~x623 & ~x649 & ~x666 & ~x676 & ~x681 & ~x698 & ~x714 & ~x738 & ~x741 & ~x747 & ~x770;
assign c217 =  x710;
assign c219 =  x318 &  x346 &  x374 & ~x2 & ~x6 & ~x21 & ~x27 & ~x49 & ~x65 & ~x83 & ~x84 & ~x141 & ~x149 & ~x164 & ~x174 & ~x191 & ~x196 & ~x222 & ~x223 & ~x250 & ~x255 & ~x282 & ~x312 & ~x315 & ~x322 & ~x339 & ~x362 & ~x364 & ~x366 & ~x367 & ~x426 & ~x447 & ~x508 & ~x611 & ~x612 & ~x614 & ~x617 & ~x620 & ~x636 & ~x637 & ~x666 & ~x676 & ~x679 & ~x700 & ~x714 & ~x715 & ~x725 & ~x729 & ~x753 & ~x754 & ~x764;
assign c221 = ~x13 & ~x27 & ~x34 & ~x44 & ~x47 & ~x48 & ~x63 & ~x66 & ~x78 & ~x93 & ~x98 & ~x106 & ~x112 & ~x125 & ~x128 & ~x147 & ~x149 & ~x152 & ~x156 & ~x167 & ~x168 & ~x171 & ~x173 & ~x174 & ~x175 & ~x196 & ~x198 & ~x252 & ~x253 & ~x334 & ~x335 & ~x338 & ~x340 & ~x342 & ~x366 & ~x416 & ~x424 & ~x443 & ~x480 & ~x505 & ~x523 & ~x525 & ~x529 & ~x534 & ~x535 & ~x540 & ~x554 & ~x561 & ~x579 & ~x581 & ~x591 & ~x616 & ~x637 & ~x664 & ~x671 & ~x704 & ~x715 & ~x722 & ~x755 & ~x768 & ~x769 & ~x772 & ~x773;
assign c223 =  x347 &  x375 & ~x26 & ~x71 & ~x97 & ~x124 & ~x125 & ~x142 & ~x249 & ~x359 & ~x398 & ~x417 & ~x448 & ~x469 & ~x471 & ~x508 & ~x552 & ~x553 & ~x607 & ~x609 & ~x611 & ~x617 & ~x646 & ~x648 & ~x666 & ~x667 & ~x716 & ~x727 & ~x750 & ~x775;
assign c225 =  x347 & ~x99 & ~x124 & ~x125 & ~x171 & ~x257 & ~x372 & ~x395 & ~x398 & ~x472 & ~x561 & ~x675 & ~x699;
assign c227 =  x320 &  x348 & ~x5 & ~x29 & ~x91 & ~x146 & ~x150 & ~x178 & ~x286 & ~x289 & ~x300 & ~x309 & ~x335 & ~x392 & ~x417 & ~x479 & ~x562 & ~x608 & ~x716 & ~x750 & ~x753;
assign c229 =  x289 &  x317 &  x345 & ~x34 & ~x109 & ~x110 & ~x168 & ~x197 & ~x224 & ~x229 & ~x286 & ~x313 & ~x389 & ~x557 & ~x624 & ~x638 & ~x665 & ~x667 & ~x705;
assign c231 =  x259 &  x343;
assign c233 =  x376 &  x657 &  x658 & ~x21 & ~x31 & ~x44 & ~x55 & ~x105 & ~x142 & ~x307 & ~x362 & ~x395 & ~x447 & ~x449 & ~x540 & ~x559 & ~x586 & ~x668 & ~x669 & ~x698 & ~x742;
assign c235 =  x316 &  x344 &  x372 &  x400;
assign c237 =  x321 &  x349 & ~x9 & ~x17 & ~x33 & ~x38 & ~x39 & ~x54 & ~x67 & ~x81 & ~x94 & ~x109 & ~x110 & ~x122 & ~x141 & ~x202 & ~x220 & ~x227 & ~x251 & ~x286 & ~x308 & ~x317 & ~x334 & ~x337 & ~x345 & ~x361 & ~x364 & ~x389 & ~x421 & ~x447 & ~x448 & ~x500 & ~x503 & ~x524 & ~x530 & ~x588 & ~x614 & ~x639 & ~x646 & ~x650 & ~x666 & ~x669 & ~x670 & ~x671 & ~x699 & ~x704 & ~x706 & ~x713 & ~x715 & ~x717 & ~x741 & ~x755 & ~x756 & ~x761 & ~x770;
assign c239 =  x343 & ~x37 & ~x546;
assign c241 = ~x2 & ~x15 & ~x37 & ~x41 & ~x53 & ~x56 & ~x58 & ~x59 & ~x81 & ~x84 & ~x134 & ~x147 & ~x162 & ~x176 & ~x311 & ~x313 & ~x337 & ~x393 & ~x400 & ~x421 & ~x425 & ~x449 & ~x453 & ~x458 & ~x472 & ~x475 & ~x511 & ~x513 & ~x523 & ~x531 & ~x540 & ~x552 & ~x569 & ~x585 & ~x612 & ~x637 & ~x661 & ~x689 & ~x694 & ~x727 & ~x749;
assign c243 =  x318 &  x345 &  x373 &  x401 & ~x58 & ~x60 & ~x170 & ~x171 & ~x284 & ~x350 & ~x376 & ~x638 & ~x649 & ~x667 & ~x691 & ~x755 & ~x771 & ~x779;
assign c245 =  x185 &  x322 &  x350 & ~x13 & ~x77 & ~x88 & ~x97 & ~x145 & ~x168 & ~x170 & ~x175 & ~x286 & ~x312 & ~x339 & ~x364 & ~x475 & ~x479 & ~x582 & ~x614 & ~x668 & ~x692 & ~x729 & ~x750;
assign c247 =  x342 &  x426;
assign c249 =  x442 &  x525;
assign c251 =  x214 &  x407 &  x433 &  x434 & ~x64 & ~x97 & ~x118 & ~x147 & ~x176 & ~x196 & ~x280 & ~x471 & ~x503 & ~x553 & ~x738 & ~x750;
assign c253 =  x318 &  x346 &  x374 & ~x1 & ~x17 & ~x34 & ~x38 & ~x54 & ~x55 & ~x63 & ~x74 & ~x88 & ~x89 & ~x91 & ~x92 & ~x94 & ~x110 & ~x118 & ~x144 & ~x145 & ~x149 & ~x163 & ~x166 & ~x171 & ~x174 & ~x175 & ~x176 & ~x199 & ~x222 & ~x227 & ~x231 & ~x252 & ~x280 & ~x307 & ~x309 & ~x313 & ~x315 & ~x337 & ~x343 & ~x360 & ~x362 & ~x366 & ~x370 & ~x422 & ~x447 & ~x471 & ~x478 & ~x505 & ~x529 & ~x530 & ~x531 & ~x534 & ~x562 & ~x563 & ~x583 & ~x585 & ~x612 & ~x617 & ~x636 & ~x639 & ~x641 & ~x646 & ~x664 & ~x665 & ~x666 & ~x675 & ~x676 & ~x713 & ~x717 & ~x718 & ~x721 & ~x724 & ~x732 & ~x738 & ~x745 & ~x747 & ~x748 & ~x755 & ~x762 & ~x764 & ~x771 & ~x781;
assign c255 =  x411 &  x440 &  x552 & ~x20 & ~x142 & ~x165 & ~x477 & ~x479 & ~x530 & ~x643 & ~x684 & ~x707 & ~x746 & ~x750;
assign c257 =  x375 &  x658 &  x659;
assign c259 =  x317 &  x345 &  x372 &  x400 & ~x1 & ~x18 & ~x58 & ~x105 & ~x115 & ~x172 & ~x249 & ~x305 & ~x310 & ~x363 & ~x364 & ~x530 & ~x585 & ~x591 & ~x640 & ~x647 & ~x648 & ~x667 & ~x698 & ~x716 & ~x733 & ~x742 & ~x754 & ~x769;
assign c261 =  x406 &  x434 & ~x2 & ~x28 & ~x58 & ~x60 & ~x97 & ~x110 & ~x144 & ~x197 & ~x228 & ~x442 & ~x449 & ~x472 & ~x475 & ~x548 & ~x552 & ~x563 & ~x576 & ~x610 & ~x635 & ~x674 & ~x691 & ~x699 & ~x717 & ~x738 & ~x749 & ~x776;
assign c263 =  x291 &  x319 &  x346 &  x347 &  x374 &  x402 & ~x21 & ~x200 & ~x260 & ~x316 & ~x528 & ~x664;
assign c265 =  x315 &  x399;
assign c267 =  x377 &  x405 & ~x23 & ~x51 & ~x74 & ~x84 & ~x110 & ~x167 & ~x334 & ~x337 & ~x364 & ~x389 & ~x487 & ~x502 & ~x513 & ~x514 & ~x638 & ~x643 & ~x745 & ~x771;
assign c269 =  x552 &  x580 & ~x10 & ~x17 & ~x58 & ~x64 & ~x82 & ~x110 & ~x118 & ~x164 & ~x167 & ~x191 & ~x199 & ~x279 & ~x280 & ~x309 & ~x338 & ~x364 & ~x507 & ~x517 & ~x528 & ~x536 & ~x547 & ~x548 & ~x587 & ~x615 & ~x695 & ~x702 & ~x705 & ~x712 & ~x725 & ~x745 & ~x748 & ~x749 & ~x751 & ~x772 & ~x776;
assign c271 =  x315 &  x371 &  x399 & ~x643;
assign c273 =  x321 &  x348 &  x349 &  x376 & ~x97 & ~x107 & ~x176 & ~x262 & ~x453 & ~x554 & ~x559 & ~x664 & ~x722 & ~x723 & ~x762;
assign c275 =  x291 &  x319 &  x347 & ~x0 & ~x14 & ~x16 & ~x40 & ~x59 & ~x65 & ~x82 & ~x86 & ~x110 & ~x168 & ~x173 & ~x175 & ~x192 & ~x194 & ~x200 & ~x203 & ~x224 & ~x269 & ~x284 & ~x315 & ~x316 & ~x366 & ~x390 & ~x417 & ~x506 & ~x528 & ~x563 & ~x590 & ~x593 & ~x615 & ~x636 & ~x645 & ~x646 & ~x691 & ~x693 & ~x721 & ~x726 & ~x744 & ~x771;
assign c277 =  x434 &  x462 & ~x106 & ~x515 & ~x543 & ~x568 & ~x570 & ~x581;
assign c279 = ~x122 & ~x162 & ~x176 & ~x286 & ~x402 & ~x421 & ~x449 & ~x459 & ~x485 & ~x487 & ~x512 & ~x513 & ~x515 & ~x530 & ~x553 & ~x641 & ~x694 & ~x749 & ~x750 & ~x759 & ~x762 & ~x766;
assign c281 = ~x60 & ~x125 & ~x128 & ~x161 & ~x389 & ~x513 & ~x540 & ~x541 & ~x542 & ~x543 & ~x555 & ~x566 & ~x568 & ~x569 & ~x570 & ~x595 & ~x649;
assign c283 =  x379 & ~x1 & ~x32 & ~x33 & ~x65 & ~x70 & ~x90 & ~x193 & ~x221 & ~x253 & ~x334 & ~x364 & ~x389 & ~x399 & ~x422 & ~x426 & ~x443 & ~x450 & ~x483 & ~x485 & ~x487 & ~x515 & ~x517 & ~x644 & ~x698 & ~x727 & ~x741 & ~x767 & ~x769 & ~x774;
assign c285 =  x323 &  x350 &  x351 & ~x0 & ~x1 & ~x16 & ~x21 & ~x53 & ~x55 & ~x58 & ~x94 & ~x99 & ~x100 & ~x106 & ~x141 & ~x226 & ~x228 & ~x231 & ~x238 & ~x289 & ~x331 & ~x339 & ~x449 & ~x469 & ~x505 & ~x529 & ~x562 & ~x611 & ~x613 & ~x614 & ~x636 & ~x640 & ~x664 & ~x666;
assign c287 =  x315 &  x426;
assign c289 =  x291 &  x319 &  x346 &  x374 &  x402 & ~x24 & ~x53 & ~x55 & ~x85 & ~x139 & ~x145 & ~x178 & ~x201 & ~x311 & ~x314 & ~x340 & ~x447 & ~x448 & ~x474 & ~x563 & ~x618 & ~x671 & ~x688 & ~x721 & ~x780 & ~x781;
assign c291 =  x442 &  x525 & ~x26 & ~x616 & ~x670 & ~x733 & ~x748;
assign c293 =  x292 &  x320 &  x347 &  x375 & ~x17 & ~x27 & ~x31 & ~x53 & ~x92 & ~x96 & ~x121 & ~x142 & ~x150 & ~x166 & ~x171 & ~x176 & ~x195 & ~x204 & ~x232 & ~x289 & ~x309 & ~x315 & ~x338 & ~x341 & ~x361 & ~x370 & ~x390 & ~x397 & ~x422 & ~x424 & ~x446 & ~x471 & ~x474 & ~x553 & ~x555 & ~x589 & ~x607 & ~x609 & ~x614 & ~x638 & ~x643 & ~x673 & ~x676 & ~x678 & ~x692 & ~x694 & ~x706 & ~x710 & ~x714 & ~x717 & ~x720 & ~x723 & ~x736 & ~x756 & ~x762 & ~x765 & ~x767 & ~x771 & ~x779;
assign c295 =  x290 &  x318 &  x346 & ~x10 & ~x11 & ~x54 & ~x117 & ~x144 & ~x196 & ~x265 & ~x672 & ~x704 & ~x711;
assign c297 =  x319 &  x347 & ~x4 & ~x21 & ~x41 & ~x224 & ~x229 & ~x240 & ~x269 & ~x280 & ~x426 & ~x453 & ~x534 & ~x558 & ~x564 & ~x646 & ~x666 & ~x667 & ~x704 & ~x755;
assign c299 =  x344 &  x372 &  x400 & ~x59 & ~x160 & ~x198 & ~x250 & ~x256 & ~x348 & ~x536 & ~x652 & ~x714;
assign c2101 =  x236 &  x437 & ~x4 & ~x128 & ~x150 & ~x156 & ~x569 & ~x570 & ~x610;
assign c2103 =  x345 &  x413 & ~x32;
assign c2105 =  x320 &  x548 & ~x1 & ~x29 & ~x41 & ~x53 & ~x56 & ~x96 & ~x113 & ~x138 & ~x148 & ~x176 & ~x202 & ~x220 & ~x228 & ~x281 & ~x289 & ~x370 & ~x393 & ~x398 & ~x470 & ~x476 & ~x500 & ~x502 & ~x527 & ~x555 & ~x585 & ~x646 & ~x651 & ~x704 & ~x771 & ~x772;
assign c2107 =  x435 &  x682 & ~x130 & ~x423 & ~x717 & ~x762;
assign c2109 =  x377 &  x378 &  x433 & ~x8 & ~x97 & ~x150 & ~x176 & ~x523 & ~x607 & ~x666;
assign c2111 =  x237 & ~x9 & ~x39 & ~x56 & ~x59 & ~x149 & ~x150 & ~x515 & ~x542 & ~x571 & ~x583 & ~x669 & ~x699;
assign c2113 =  x320 &  x321 &  x348 & ~x2 & ~x20 & ~x27 & ~x66 & ~x93 & ~x117 & ~x167 & ~x176 & ~x207 & ~x228 & ~x290 & ~x333 & ~x414 & ~x444 & ~x475 & ~x582 & ~x608 & ~x614 & ~x640 & ~x660 & ~x664 & ~x671 & ~x674 & ~x690 & ~x702 & ~x721 & ~x726 & ~x772;
assign c2115 =  x523 &  x632 & ~x23 & ~x66 & ~x84 & ~x162 & ~x251 & ~x337 & ~x364 & ~x421 & ~x423 & ~x449 & ~x506 & ~x563 & ~x583 & ~x610 & ~x617 & ~x646 & ~x766;
assign c2117 =  x348 &  x376 &  x377 &  x434 & ~x39 & ~x56 & ~x427 & ~x498 & ~x501 & ~x639 & ~x643;
assign c2119 =  x289 &  x317 &  x345 &  x373 & ~x30 & ~x616 & ~x667 & ~x707;
assign c2121 = ~x33 & ~x42 & ~x46 & ~x63 & ~x85 & ~x124 & ~x156 & ~x191 & ~x196 & ~x280 & ~x285 & ~x286 & ~x334 & ~x389 & ~x392 & ~x427 & ~x503 & ~x512 & ~x530 & ~x536 & ~x540 & ~x541 & ~x568 & ~x581 & ~x584 & ~x637 & ~x674 & ~x689 & ~x690 & ~x781;
assign c2123 =  x378 & ~x12 & ~x13 & ~x21 & ~x88 & ~x97 & ~x168 & ~x235 & ~x236 & ~x263 & ~x371 & ~x385 & ~x417 & ~x448 & ~x479;
assign c2125 =  x317 &  x345 &  x373 & ~x8 & ~x27 & ~x53 & ~x56 & ~x60 & ~x106 & ~x110 & ~x134 & ~x219 & ~x252 & ~x256 & ~x309 & ~x348 & ~x395 & ~x419 & ~x586 & ~x639 & ~x643 & ~x646 & ~x653 & ~x666 & ~x671 & ~x672 & ~x704 & ~x715 & ~x718 & ~x721 & ~x732 & ~x733 & ~x739 & ~x743 & ~x756 & ~x761 & ~x763 & ~x766 & ~x776;
assign c2127 =  x350 &  x351 &  x378 & ~x41 & ~x150 & ~x170 & ~x177 & ~x470 & ~x523 & ~x552;
assign c2129 =  x349 &  x350 &  x658 & ~x8 & ~x39 & ~x87 & ~x91 & ~x93 & ~x137 & ~x195 & ~x360 & ~x732 & ~x735;
assign c2131 =  x287 &  x398 & ~x623;
assign c2133 =  x233 &  x260 &  x288 &  x316 & ~x52 & ~x313 & ~x337 & ~x616 & ~x646 & ~x681 & ~x706 & ~x783;
assign c2135 =  x434 & ~x0 & ~x8 & ~x10 & ~x24 & ~x57 & ~x58 & ~x96 & ~x97 & ~x125 & ~x145 & ~x150 & ~x168 & ~x198 & ~x232 & ~x260 & ~x280 & ~x289 & ~x338 & ~x389 & ~x391 & ~x398 & ~x448 & ~x454 & ~x507 & ~x510 & ~x523 & ~x524 & ~x532 & ~x534 & ~x577 & ~x583 & ~x632 & ~x633 & ~x637 & ~x639 & ~x690 & ~x704 & ~x727 & ~x735 & ~x737 & ~x741 & ~x752 & ~x755 & ~x759 & ~x776;
assign c2137 =  x264 & ~x96 & ~x198 & ~x201 & ~x434 & ~x461 & ~x462 & ~x488 & ~x489 & ~x503 & ~x582 & ~x611 & ~x639 & ~x667 & ~x759;
assign c2139 = ~x250 & ~x336 & ~x459 & ~x462 & ~x487 & ~x488 & ~x489 & ~x545 & ~x546 & ~x547 & ~x617 & ~x669 & ~x721;
assign c2141 =  x290 &  x345 &  x373 &  x401 &  x429 & ~x3 & ~x255 & ~x321 & ~x693;
assign c2143 =  x346 &  x374 & ~x1 & ~x8 & ~x9 & ~x22 & ~x51 & ~x52 & ~x53 & ~x55 & ~x81 & ~x84 & ~x95 & ~x107 & ~x110 & ~x114 & ~x123 & ~x140 & ~x146 & ~x189 & ~x243 & ~x280 & ~x286 & ~x300 & ~x308 & ~x309 & ~x313 & ~x341 & ~x362 & ~x394 & ~x398 & ~x416 & ~x417 & ~x418 & ~x422 & ~x447 & ~x507 & ~x528 & ~x562 & ~x582 & ~x585 & ~x589 & ~x609 & ~x610 & ~x612 & ~x614 & ~x674 & ~x697 & ~x708 & ~x721 & ~x738 & ~x741 & ~x745 & ~x755 & ~x757 & ~x762 & ~x765 & ~x766 & ~x772 & ~x773 & ~x776;
assign c2145 =  x319 &  x347 &  x375 & ~x1 & ~x2 & ~x8 & ~x9 & ~x30 & ~x33 & ~x39 & ~x51 & ~x52 & ~x60 & ~x74 & ~x76 & ~x85 & ~x94 & ~x97 & ~x144 & ~x147 & ~x168 & ~x174 & ~x257 & ~x309 & ~x334 & ~x371 & ~x390 & ~x395 & ~x396 & ~x417 & ~x422 & ~x450 & ~x506 & ~x531 & ~x561 & ~x581 & ~x582 & ~x583 & ~x614 & ~x636 & ~x644 & ~x666 & ~x670 & ~x695 & ~x699 & ~x705 & ~x737 & ~x755 & ~x763 & ~x771 & ~x774;
assign c2147 =  x344 &  x372 &  x400 & ~x9 & ~x51 & ~x52 & ~x59 & ~x72 & ~x137 & ~x171 & ~x199 & ~x306 & ~x313 & ~x348 & ~x424 & ~x449 & ~x450 & ~x479 & ~x532 & ~x587 & ~x591 & ~x616 & ~x619 & ~x643 & ~x646 & ~x650 & ~x666 & ~x671 & ~x707 & ~x729 & ~x737 & ~x741 & ~x748 & ~x750 & ~x761 & ~x766;
assign c2149 =  x348 & ~x0 & ~x20 & ~x59 & ~x64 & ~x95 & ~x358 & ~x456 & ~x484 & ~x501 & ~x508 & ~x517 & ~x545 & ~x585 & ~x718 & ~x746;
assign c2151 =  x233 &  x261 & ~x41 & ~x52 & ~x169 & ~x599 & ~x614 & ~x619 & ~x639 & ~x706 & ~x724 & ~x749 & ~x766;
assign c2153 = ~x4 & ~x71 & ~x111 & ~x472 & ~x513 & ~x517 & ~x543 & ~x545 & ~x573 & ~x585 & ~x610;
assign c2155 =  x342 &  x370 &  x426;
assign c2157 =  x351 & ~x41 & ~x72 & ~x77 & ~x139 & ~x223 & ~x358 & ~x486 & ~x487 & ~x488 & ~x489 & ~x515 & ~x743;
assign c2159 = ~x11 & ~x76 & ~x199 & ~x278 & ~x311 & ~x337 & ~x448 & ~x449 & ~x459 & ~x460 & ~x461 & ~x462 & ~x463 & ~x487 & ~x488 & ~x489 & ~x515 & ~x516 & ~x517 & ~x518 & ~x519 & ~x616 & ~x667 & ~x668 & ~x730 & ~x739;
assign c2161 =  x433 &  x656 &  x657 & ~x4 & ~x50 & ~x52 & ~x56 & ~x59 & ~x74 & ~x83 & ~x84 & ~x86 & ~x94 & ~x109 & ~x117 & ~x123 & ~x137 & ~x251 & ~x308 & ~x311 & ~x412 & ~x424 & ~x452 & ~x479 & ~x480 & ~x532 & ~x536 & ~x557 & ~x588 & ~x611 & ~x614 & ~x619 & ~x646 & ~x674 & ~x692 & ~x694 & ~x696 & ~x701 & ~x706 & ~x727 & ~x749;
assign c2163 =  x267 & ~x96 & ~x123 & ~x124 & ~x168 & ~x453 & ~x542 & ~x568 & ~x694 & ~x747 & ~x762;
assign c2165 =  x660 & ~x7 & ~x8 & ~x30 & ~x33 & ~x37 & ~x52 & ~x56 & ~x80 & ~x88 & ~x89 & ~x94 & ~x96 & ~x110 & ~x130 & ~x146 & ~x190 & ~x198 & ~x221 & ~x251 & ~x340 & ~x390 & ~x394 & ~x418 & ~x422 & ~x448 & ~x476 & ~x479 & ~x532 & ~x535 & ~x545 & ~x546 & ~x596 & ~x613 & ~x614 & ~x682 & ~x711 & ~x751 & ~x756 & ~x761 & ~x767 & ~x775 & ~x776;
assign c2167 =  x319 &  x320 &  x347 &  x348 & ~x14 & ~x45 & ~x48 & ~x195 & ~x199 & ~x336 & ~x344 & ~x399 & ~x471 & ~x582 & ~x665 & ~x689 & ~x719 & ~x748;
assign c2169 =  x316 &  x371 &  x399 & ~x109 & ~x530 & ~x651 & ~x766;
assign c2171 =  x288 &  x400;
assign c2173 =  x406 &  x433 &  x434 &  x435 & ~x4 & ~x10 & ~x39 & ~x59 & ~x87 & ~x93 & ~x123 & ~x124 & ~x167 & ~x168 & ~x176 & ~x194 & ~x199 & ~x250 & ~x309 & ~x417 & ~x505 & ~x509 & ~x510 & ~x524 & ~x539 & ~x552 & ~x563 & ~x704 & ~x732 & ~x733 & ~x737 & ~x770 & ~x771 & ~x776;
assign c2175 = ~x3 & ~x9 & ~x33 & ~x48 & ~x52 & ~x84 & ~x87 & ~x97 & ~x111 & ~x121 & ~x125 & ~x141 & ~x150 & ~x151 & ~x152 & ~x156 & ~x173 & ~x202 & ~x276 & ~x285 & ~x309 & ~x315 & ~x332 & ~x343 & ~x387 & ~x396 & ~x472 & ~x478 & ~x479 & ~x509 & ~x523 & ~x550 & ~x552 & ~x554 & ~x576 & ~x644 & ~x646 & ~x660 & ~x664 & ~x716 & ~x750 & ~x762;
assign c2177 =  x437 & ~x97 & ~x304 & ~x350 & ~x508 & ~x540 & ~x542 & ~x543 & ~x568 & ~x569 & ~x570 & ~x755;
assign c2179 =  x319 &  x347 &  x548 & ~x41 & ~x75 & ~x89 & ~x91 & ~x178 & ~x281 & ~x423 & ~x552 & ~x580 & ~x636 & ~x735;
assign c2181 =  x243 &  x271 & ~x20 & ~x33 & ~x34 & ~x39 & ~x41 & ~x52 & ~x97 & ~x158 & ~x167 & ~x176 & ~x198 & ~x199 & ~x282 & ~x334 & ~x337 & ~x480 & ~x532 & ~x566 & ~x674 & ~x745 & ~x749;
assign c2183 =  x318 &  x346 &  x374 & ~x1 & ~x10 & ~x17 & ~x29 & ~x31 & ~x53 & ~x56 & ~x61 & ~x86 & ~x110 & ~x137 & ~x168 & ~x222 & ~x251 & ~x256 & ~x294 & ~x313 & ~x390 & ~x419 & ~x424 & ~x557 & ~x562 & ~x592 & ~x622 & ~x639 & ~x654 & ~x675 & ~x700 & ~x727 & ~x770;
assign c2185 =  x350 &  x351 &  x379 &  x407 & ~x59 & ~x96 & ~x97 & ~x99 & ~x111 & ~x119 & ~x165 & ~x176 & ~x289 & ~x314 & ~x372 & ~x447 & ~x582 & ~x608 & ~x664 & ~x754 & ~x775;
assign c2187 =  x411 & ~x538 & ~x568 & ~x570 & ~x595 & ~x614 & ~x755;
assign c2189 = ~x2 & ~x250 & ~x457 & ~x487 & ~x514 & ~x515 & ~x517 & ~x543 & ~x545 & ~x678 & ~x722;
assign c2191 =  x321 &  x349 & ~x3 & ~x16 & ~x25 & ~x43 & ~x81 & ~x89 & ~x97 & ~x114 & ~x143 & ~x166 & ~x168 & ~x176 & ~x204 & ~x230 & ~x232 & ~x258 & ~x260 & ~x442 & ~x451 & ~x480 & ~x524 & ~x526 & ~x532 & ~x533 & ~x583 & ~x609 & ~x622 & ~x637 & ~x650 & ~x666 & ~x720 & ~x738 & ~x747 & ~x755 & ~x771;
assign c2193 =  x372 &  x400 &  x428 & ~x2 & ~x8 & ~x16 & ~x28 & ~x48 & ~x51 & ~x63 & ~x80 & ~x90 & ~x106 & ~x141 & ~x144 & ~x168 & ~x254 & ~x276 & ~x309 & ~x338 & ~x366 & ~x375 & ~x378 & ~x392 & ~x477 & ~x532 & ~x640 & ~x649 & ~x666 & ~x677 & ~x731 & ~x741 & ~x747 & ~x750 & ~x779;
assign c2195 =  x261 &  x659 & ~x18 & ~x56 & ~x93 & ~x117 & ~x134 & ~x139 & ~x223 & ~x246 & ~x280 & ~x641 & ~x651 & ~x693 & ~x717 & ~x745 & ~x759;
assign c2197 =  x320 &  x348 &  x376 & ~x58 & ~x91 & ~x96 & ~x151 & ~x168 & ~x251 & ~x256 & ~x280 & ~x336 & ~x370 & ~x393 & ~x442 & ~x445 & ~x470 & ~x500 & ~x505 & ~x536 & ~x553 & ~x554 & ~x563 & ~x581 & ~x665 & ~x691 & ~x705 & ~x750 & ~x752 & ~x760;
assign c2199 = ~x23 & ~x24 & ~x76 & ~x86 & ~x91 & ~x123 & ~x126 & ~x127 & ~x168 & ~x177 & ~x197 & ~x198 & ~x204 & ~x207 & ~x209 & ~x210 & ~x278 & ~x280 & ~x288 & ~x341 & ~x440 & ~x480 & ~x533 & ~x607 & ~x619 & ~x639 & ~x646 & ~x673 & ~x674 & ~x691 & ~x708 & ~x745 & ~x749 & ~x761;
assign c2201 =  x375 &  x376 & ~x6 & ~x34 & ~x37 & ~x45 & ~x58 & ~x198 & ~x199 & ~x255 & ~x280 & ~x361 & ~x424 & ~x480 & ~x485 & ~x510 & ~x588 & ~x718 & ~x733 & ~x775;
assign c2203 = ~x2 & ~x10 & ~x66 & ~x121 & ~x128 & ~x158 & ~x168 & ~x251 & ~x280 & ~x309 & ~x367 & ~x389 & ~x446 & ~x449 & ~x506 & ~x510 & ~x533 & ~x541 & ~x542 & ~x543 & ~x552 & ~x568 & ~x569 & ~x570 & ~x664 & ~x699 & ~x727 & ~x782;
assign c2205 =  x317 &  x345 & ~x240 & ~x267 & ~x423 & ~x595 & ~x667;
assign c2207 =  x321 &  x348 &  x376 & ~x3 & ~x4 & ~x9 & ~x10 & ~x23 & ~x47 & ~x54 & ~x70 & ~x83 & ~x96 & ~x110 & ~x168 & ~x198 & ~x201 & ~x207 & ~x230 & ~x252 & ~x260 & ~x289 & ~x309 & ~x388 & ~x415 & ~x416 & ~x424 & ~x471 & ~x472 & ~x553 & ~x617 & ~x636 & ~x666 & ~x690 & ~x692 & ~x697 & ~x698 & ~x732 & ~x741 & ~x751 & ~x764 & ~x765 & ~x774;
assign c2209 =  x270 & ~x26 & ~x55 & ~x74 & ~x87 & ~x94 & ~x97 & ~x127 & ~x146 & ~x148 & ~x309 & ~x333 & ~x342 & ~x399 & ~x414 & ~x453 & ~x530 & ~x540 & ~x588 & ~x664 & ~x694 & ~x714 & ~x720;
assign c2211 =  x344 &  x372 &  x400 &  x428 & ~x375;
assign c2213 =  x373 &  x401 &  x430 & ~x8 & ~x16 & ~x22 & ~x24 & ~x32 & ~x69 & ~x71 & ~x83 & ~x89 & ~x97 & ~x139 & ~x167 & ~x168 & ~x171 & ~x174 & ~x196 & ~x221 & ~x277 & ~x280 & ~x308 & ~x362 & ~x366 & ~x389 & ~x399 & ~x505 & ~x506 & ~x614 & ~x644 & ~x666 & ~x694 & ~x697 & ~x701 & ~x702 & ~x717 & ~x718 & ~x720 & ~x724 & ~x727 & ~x738 & ~x741 & ~x746 & ~x749 & ~x755 & ~x764 & ~x771 & ~x777;
assign c2215 =  x350 &  x351 &  x379 & ~x53 & ~x89 & ~x97 & ~x100 & ~x150 & ~x167 & ~x309 & ~x421 & ~x588 & ~x632;
assign c2217 =  x342 &  x426;
assign c2219 =  x523 & ~x10 & ~x68 & ~x89 & ~x221 & ~x251 & ~x308 & ~x389 & ~x390 & ~x517 & ~x532 & ~x545 & ~x546 & ~x547 & ~x548 & ~x557 & ~x589 & ~x617 & ~x646 & ~x755;
assign c2221 = ~x3 & ~x15 & ~x28 & ~x37 & ~x92 & ~x95 & ~x97 & ~x99 & ~x124 & ~x156 & ~x168 & ~x170 & ~x286 & ~x495 & ~x511 & ~x548 & ~x564 & ~x592 & ~x619 & ~x633 & ~x634 & ~x647 & ~x688 & ~x721 & ~x722 & ~x754 & ~x756 & ~x769 & ~x770;
assign c2223 =  x347 &  x375 &  x376 & ~x0 & ~x4 & ~x9 & ~x12 & ~x17 & ~x33 & ~x37 & ~x39 & ~x41 & ~x74 & ~x84 & ~x85 & ~x110 & ~x117 & ~x118 & ~x144 & ~x145 & ~x146 & ~x150 & ~x167 & ~x194 & ~x201 & ~x222 & ~x224 & ~x248 & ~x249 & ~x252 & ~x253 & ~x254 & ~x286 & ~x287 & ~x334 & ~x340 & ~x366 & ~x389 & ~x391 & ~x416 & ~x425 & ~x427 & ~x443 & ~x445 & ~x474 & ~x476 & ~x477 & ~x480 & ~x505 & ~x534 & ~x553 & ~x583 & ~x589 & ~x611 & ~x612 & ~x614 & ~x616 & ~x618 & ~x636 & ~x637 & ~x643 & ~x646 & ~x675 & ~x700 & ~x701 & ~x702 & ~x721 & ~x722 & ~x729 & ~x740 & ~x748 & ~x749 & ~x750 & ~x761 & ~x767 & ~x770 & ~x771 & ~x773 & ~x775 & ~x776;
assign c2225 =  x267 & ~x0 & ~x9 & ~x61 & ~x69 & ~x79 & ~x87 & ~x88 & ~x94 & ~x96 & ~x105 & ~x106 & ~x117 & ~x140 & ~x149 & ~x150 & ~x195 & ~x198 & ~x226 & ~x250 & ~x278 & ~x307 & ~x308 & ~x335 & ~x341 & ~x362 & ~x418 & ~x471 & ~x474 & ~x487 & ~x488 & ~x582 & ~x589 & ~x606 & ~x611 & ~x634 & ~x639 & ~x641 & ~x643 & ~x670 & ~x672 & ~x674 & ~x693 & ~x700 & ~x723 & ~x754 & ~x757 & ~x771;
assign c2227 =  x260 & ~x156 & ~x168 & ~x569 & ~x570 & ~x571;
assign c2229 =  x240 & ~x36 & ~x175 & ~x337 & ~x417 & ~x513 & ~x536 & ~x541 & ~x577 & ~x640 & ~x646 & ~x674 & ~x782;
assign c2231 =  x320 &  x348 & ~x1 & ~x36 & ~x68 & ~x93 & ~x139 & ~x149 & ~x150 & ~x259 & ~x386 & ~x393 & ~x554 & ~x555 & ~x583 & ~x639 & ~x653 & ~x654 & ~x664 & ~x717 & ~x733 & ~x748 & ~x753 & ~x768;
assign c2233 =  x370 &  x398;
assign c2235 =  x303 & ~x121 & ~x123;
assign c2237 =  x319 & ~x30 & ~x44 & ~x70 & ~x96 & ~x118 & ~x151 & ~x198 & ~x283 & ~x339 & ~x367 & ~x370 & ~x416 & ~x417 & ~x422 & ~x452 & ~x488 & ~x528 & ~x588 & ~x589 & ~x674 & ~x700 & ~x704 & ~x707 & ~x724 & ~x757 & ~x768;
assign c2239 =  x407 &  x435 &  x464 &  x659 & ~x137 & ~x545;
assign c2241 =  x233 &  x261 &  x289 &  x317 & ~x168 & ~x338 & ~x417 & ~x666 & ~x714;
assign c2243 =  x323 &  x350 &  x351 & ~x4 & ~x9 & ~x10 & ~x11 & ~x16 & ~x55 & ~x84 & ~x89 & ~x121 & ~x168 & ~x170 & ~x174 & ~x175 & ~x252 & ~x289 & ~x310 & ~x364 & ~x389 & ~x393 & ~x421 & ~x423 & ~x428 & ~x503 & ~x505 & ~x552 & ~x564 & ~x583 & ~x606 & ~x619 & ~x639 & ~x664 & ~x678 & ~x707 & ~x716 & ~x717 & ~x745 & ~x752 & ~x770 & ~x775;
assign c2245 =  x411 & ~x27 & ~x85 & ~x108 & ~x388 & ~x444 & ~x449 & ~x503 & ~x510 & ~x540 & ~x566 & ~x568 & ~x570 & ~x625 & ~x670 & ~x727 & ~x761;
assign c2247 =  x271 & ~x16 & ~x23 & ~x25 & ~x27 & ~x28 & ~x30 & ~x41 & ~x47 & ~x59 & ~x60 & ~x94 & ~x119 & ~x124 & ~x125 & ~x130 & ~x131 & ~x139 & ~x156 & ~x165 & ~x176 & ~x198 & ~x224 & ~x337 & ~x365 & ~x389 & ~x394 & ~x414 & ~x427 & ~x443 & ~x446 & ~x477 & ~x502 & ~x529 & ~x532 & ~x536 & ~x537 & ~x563 & ~x581 & ~x590 & ~x609 & ~x637 & ~x639 & ~x643 & ~x662 & ~x663 & ~x666 & ~x697 & ~x700 & ~x717 & ~x720 & ~x725 & ~x726 & ~x745;
assign c2249 = ~x6 & ~x56 & ~x60 & ~x89 & ~x97 & ~x144 & ~x162 & ~x194 & ~x282 & ~x334 & ~x432 & ~x433 & ~x459 & ~x461 & ~x488 & ~x489 & ~x517 & ~x545;
assign c2251 =  x291 &  x319 &  x346 &  x374 &  x402 & ~x6 & ~x11 & ~x18 & ~x19 & ~x20 & ~x33 & ~x42 & ~x47 & ~x54 & ~x61 & ~x110 & ~x111 & ~x118 & ~x137 & ~x173 & ~x176 & ~x195 & ~x231 & ~x255 & ~x259 & ~x280 & ~x286 & ~x307 & ~x341 & ~x369 & ~x370 & ~x391 & ~x394 & ~x420 & ~x556 & ~x562 & ~x613 & ~x615 & ~x643 & ~x663 & ~x664 & ~x677 & ~x700 & ~x708 & ~x710 & ~x729 & ~x734 & ~x740 & ~x744 & ~x745 & ~x750 & ~x753 & ~x756 & ~x771 & ~x774 & ~x775 & ~x779;
assign c2253 =  x190 & ~x131;
assign c2255 =  x455 & ~x0 & ~x10 & ~x16 & ~x18 & ~x28 & ~x40 & ~x46 & ~x47 & ~x49 & ~x51 & ~x53 & ~x57 & ~x64 & ~x66 & ~x84 & ~x88 & ~x91 & ~x117 & ~x120 & ~x167 & ~x198 & ~x222 & ~x228 & ~x251 & ~x256 & ~x277 & ~x279 & ~x281 & ~x393 & ~x394 & ~x403 & ~x405 & ~x407 & ~x418 & ~x422 & ~x433 & ~x434 & ~x477 & ~x507 & ~x534 & ~x558 & ~x563 & ~x612 & ~x614 & ~x640 & ~x641 & ~x646 & ~x668 & ~x681 & ~x682 & ~x698 & ~x705 & ~x706 & ~x707 & ~x708 & ~x724 & ~x738 & ~x740 & ~x746 & ~x749 & ~x756 & ~x761 & ~x765 & ~x771;
assign c2257 =  x350 &  x434 & ~x96 & ~x167 & ~x168 & ~x176 & ~x178 & ~x337 & ~x364 & ~x427 & ~x496 & ~x762;
assign c2259 =  x442 &  x525;
assign c2261 =  x378 &  x379 &  x380 &  x407 & ~x0 & ~x4 & ~x85 & ~x143 & ~x167 & ~x280 & ~x335 & ~x448 & ~x500 & ~x515 & ~x516 & ~x517 & ~x588 & ~x611 & ~x677 & ~x696 & ~x707 & ~x727 & ~x762;
assign c2263 =  x287 &  x315 & ~x60 & ~x620 & ~x671 & ~x782;
assign c2265 =  x321 &  x348 &  x376 & ~x148 & ~x198 & ~x228 & ~x229 & ~x343 & ~x393 & ~x420 & ~x427 & ~x454 & ~x472 & ~x530 & ~x554 & ~x622 & ~x650 & ~x705 & ~x737 & ~x741 & ~x765 & ~x771;
assign c2269 =  x349 &  x350 &  x351 & ~x28 & ~x88 & ~x145 & ~x194 & ~x199 & ~x250 & ~x341 & ~x389 & ~x421 & ~x425 & ~x427 & ~x485 & ~x585 & ~x615 & ~x641 & ~x706;
assign c2271 =  x357 & ~x12 & ~x30 & ~x72 & ~x132 & ~x170 & ~x224 & ~x451 & ~x505 & ~x537 & ~x560 & ~x566 & ~x593 & ~x636 & ~x760 & ~x776 & ~x777;
assign c2273 =  x343 &  x371 &  x427 &  x455;
assign c2275 =  x217 &  x407 & ~x63 & ~x152 & ~x194 & ~x338 & ~x475 & ~x537 & ~x552 & ~x565 & ~x612;
assign c2277 =  x239 &  x240 & ~x50 & ~x56 & ~x97 & ~x106 & ~x124 & ~x511 & ~x555 & ~x568 & ~x580 & ~x588 & ~x608 & ~x614 & ~x636 & ~x689 & ~x719 & ~x771;
assign c2279 =  x350 &  x378 &  x379 & ~x4 & ~x11 & ~x47 & ~x76 & ~x167 & ~x168 & ~x175 & ~x178 & ~x196 & ~x198 & ~x256 & ~x286 & ~x309 & ~x341 & ~x359 & ~x364 & ~x415 & ~x419 & ~x425 & ~x427 & ~x478 & ~x497 & ~x552 & ~x611 & ~x632 & ~x638 & ~x664 & ~x728 & ~x738 & ~x760 & ~x771;
assign c2281 = ~x3 & ~x8 & ~x162 & ~x167 & ~x309 & ~x514 & ~x515 & ~x516 & ~x517 & ~x518 & ~x543 & ~x545 & ~x546 & ~x547 & ~x646 & ~x650 & ~x747 & ~x755;
assign c2283 =  x319 &  x320 &  x347 & ~x8 & ~x89 & ~x168 & ~x243 & ~x283 & ~x370 & ~x389 & ~x530 & ~x558 & ~x614 & ~x651 & ~x749 & ~x755 & ~x762 & ~x771;
assign c2285 =  x377 &  x433 & ~x78 & ~x79 & ~x97 & ~x123 & ~x144 & ~x168 & ~x334 & ~x427 & ~x442 & ~x458 & ~x553 & ~x614 & ~x643 & ~x696;
assign c2287 =  x321 &  x349 & ~x8 & ~x63 & ~x66 & ~x97 & ~x124 & ~x145 & ~x150 & ~x168 & ~x176 & ~x250 & ~x260 & ~x290 & ~x333 & ~x370 & ~x390 & ~x454 & ~x563 & ~x646 & ~x670 & ~x674 & ~x704 & ~x717 & ~x731 & ~x736 & ~x750;
assign c2289 =  x322 &  x349 &  x350 &  x351 &  x379 &  x380 & ~x109 & ~x362 & ~x751 & ~x771 & ~x777;
assign c2291 = ~x21 & ~x51 & ~x58 & ~x59 & ~x69 & ~x128 & ~x141 & ~x152 & ~x160 & ~x224 & ~x252 & ~x331 & ~x361 & ~x362 & ~x479 & ~x510 & ~x542 & ~x543 & ~x566 & ~x569 & ~x570 & ~x591 & ~x611 & ~x617 & ~x619 & ~x646 & ~x701 & ~x707 & ~x749 & ~x755 & ~x761;
assign c2293 = ~x28 & ~x39 & ~x86 & ~x91 & ~x137 & ~x150 & ~x158 & ~x164 & ~x340 & ~x503 & ~x540 & ~x541 & ~x543 & ~x555 & ~x569 & ~x570 & ~x624 & ~x643 & ~x762;
assign c2295 =  x350 &  x378 &  x658 & ~x4 & ~x18 & ~x30 & ~x48 & ~x59 & ~x60 & ~x88 & ~x95 & ~x111 & ~x143 & ~x162 & ~x167 & ~x168 & ~x190 & ~x198 & ~x251 & ~x276 & ~x304 & ~x329 & ~x423 & ~x453 & ~x454 & ~x472 & ~x477 & ~x504 & ~x557 & ~x591 & ~x643 & ~x646 & ~x648 & ~x666 & ~x669 & ~x674 & ~x700 & ~x718 & ~x719 & ~x722 & ~x753 & ~x755 & ~x763 & ~x766 & ~x771 & ~x773;
assign c2297 = ~x8 & ~x56 & ~x59 & ~x72 & ~x93 & ~x111 & ~x167 & ~x221 & ~x253 & ~x256 & ~x308 & ~x389 & ~x434 & ~x435 & ~x458 & ~x459 & ~x460 & ~x461 & ~x462 & ~x463 & ~x487 & ~x488 & ~x489 & ~x491 & ~x515 & ~x516 & ~x518 & ~x610 & ~x643 & ~x646 & ~x665 & ~x666 & ~x699 & ~x761;
assign c2299 =  x317 &  x345 &  x372 &  x400 &  x428 & ~x37 & ~x42 & ~x47 & ~x108 & ~x194 & ~x226 & ~x252 & ~x283 & ~x337 & ~x338 & ~x364 & ~x639 & ~x648 & ~x679 & ~x697 & ~x719;
assign c30 =  x183 &  x434 &  x460 & ~x320 & ~x346;
assign c34 =  x145;
assign c36 =  x90;
assign c38 =  x156 &  x626 & ~x136 & ~x236 & ~x288 & ~x458;
assign c310 =  x207 &  x208 &  x209 &  x268 &  x295 &  x322 & ~x13 & ~x49 & ~x65 & ~x272 & ~x300 & ~x369 & ~x416 & ~x703;
assign c312 =  x380 &  x536 & ~x400;
assign c314 =  x154 &  x240 &  x322 & ~x158 & ~x244 & ~x459 & ~x461;
assign c316 =  x591;
assign c318 =  x759;
assign c320 =  x28;
assign c322 =  x507;
assign c324 =  x150 &  x265;
assign c328 =  x57;
assign c330 =  x211 & ~x190 & ~x228 & ~x301 & ~x319 & ~x484 & ~x573 & ~x600 & ~x602;
assign c332 =  x212 &  x213 &  x404 &  x405 & ~x94 & ~x122 & ~x198 & ~x315 & ~x321 & ~x347 & ~x373 & ~x374 & ~x423 & ~x483 & ~x619 & ~x767;
assign c334 =  x177 &  x264 &  x552;
assign c336 =  x298 &  x378 &  x601 & ~x26 & ~x198 & ~x248 & ~x255 & ~x290 & ~x292 & ~x451 & ~x502 & ~x503 & ~x586 & ~x617 & ~x691;
assign c338 =  x756;
assign c340 =  x434 &  x657 & ~x191 & ~x249 & ~x320 & ~x572 & ~x573 & ~x612;
assign c342 =  x626 &  x628 & ~x263 & ~x366 & ~x431 & ~x441 & ~x458 & ~x462 & ~x475 & ~x645 & ~x691;
assign c344 =  x198;
assign c346 =  x272 &  x299 &  x353 &  x381 &  x595 & ~x458;
assign c348 =  x636;
assign c350 =  x265 &  x553;
assign c352 =  x293 &  x526;
assign c354 =  x211 &  x212 &  x213 &  x297 &  x378 &  x406 &  x438 &  x467 & ~x370;
assign c356 =  x575 &  x601 &  x627 &  x628 &  x629 & ~x37 & ~x83 & ~x191 & ~x203 & ~x220 & ~x301 & ~x371 & ~x373 & ~x458 & ~x543;
assign c358 =  x325 &  x596 &  x599 &  x601 &  x602 &  x627 & ~x710;
assign c360 =  x267 &  x496 &  x579 & ~x371;
assign c362 =  x298 &  x377 & ~x47 & ~x228 & ~x319 & ~x320 & ~x484 & ~x561;
assign c364 =  x685 & ~x215 & ~x571 & ~x573 & ~x574 & ~x627;
assign c366 =  x589;
assign c368 =  x180 & ~x81 & ~x87 & ~x263 & ~x264 & ~x265 & ~x344 & ~x413 & ~x502 & ~x571 & ~x572 & ~x581 & ~x664;
assign c370 =  x123 &  x629 & ~x234 & ~x244;
assign c372 =  x418;
assign c374 =  x86;
assign c376 =  x95;
assign c378 =  x256;
assign c380 =  x126 &  x321 & ~x433;
assign c382 =  x178 &  x238 &  x292 & ~x189;
assign c384 =  x184 &  x297 &  x323 &  x547 & ~x289 & ~x609 & ~x659;
assign c386 =  x154 &  x654 & ~x236 & ~x263;
assign c388 =  x298 &  x323 &  x325 &  x596 &  x597 & ~x290 & ~x431;
assign c390 =  x209 &  x213 &  x268 &  x295 &  x322 &  x628 & ~x244 & ~x272;
assign c392 =  x678;
assign c394 =  x504;
assign c396 =  x560;
assign c398 =  x533;
assign c3100 =  x52;
assign c3102 =  x684 & ~x317 & ~x628;
assign c3104 =  x209 &  x211 &  x405 & ~x88 & ~x120 & ~x122 & ~x217 & ~x248 & ~x293 & ~x320 & ~x347 & ~x374 & ~x399 & ~x400 & ~x611;
assign c3106 =  x686 & ~x373 & ~x573 & ~x600 & ~x601 & ~x602 & ~x628;
assign c3108 =  x536;
assign c3110 =  x561;
assign c3112 =  x56;
assign c3114 =  x229 &  x293;
assign c3116 =  x778;
assign c3118 =  x266 &  x606 &  x632 & ~x214;
assign c3120 =  x208 &  x209 &  x235 & ~x71 & ~x319 & ~x320 & ~x347 & ~x374 & ~x572;
assign c3122 =  x648;
assign c3124 =  x297 &  x322 &  x323 & ~x264 & ~x289;
assign c3126 =  x78;
assign c3128 =  x209 &  x629 &  x653 & ~x347 & ~x371 & ~x540;
assign c3130 =  x140;
assign c3132 =  x212 &  x244 &  x381 &  x405 & ~x320 & ~x399;
assign c3134 =  x241 &  x377 &  x381 &  x409 &  x552 & ~x492;
assign c3136 =  x173;
assign c3138 =  x156 &  x270 &  x297 &  x322 &  x599;
assign c3140 =  x393;
assign c3142 =  x177 &  x178 &  x293 & ~x158 & ~x214 & ~x244;
assign c3144 =  x632 & ~x262 & ~x263 & ~x318 & ~x573 & ~x670;
assign c3146 =  x178 &  x686 & ~x185 & ~x272 & ~x327 & ~x571;
assign c3148 =  x124 &  x321 & ~x207;
assign c3150 =  x656 & ~x215 & ~x262 & ~x289 & ~x299 & ~x546;
assign c3152 =  x308;
assign c3154 =  x336;
assign c3156 =  x152 &  x576 &  x631 & ~x290 & ~x517 & ~x518;
assign c3158 =  x175 &  x293;
assign c3160 =  x378 &  x548 &  x575 & ~x40 & ~x81 & ~x174 & ~x233 & ~x287 & ~x289 & ~x319 & ~x320 & ~x335 & ~x497 & ~x662 & ~x719;
assign c3162 =  x326 &  x404 &  x405 &  x406 &  x655 & ~x320;
assign c3164 =  x151 &  x294 & ~x207;
assign c3166 =  x750;
assign c3168 =  x116;
assign c3170 =  x223;
assign c3172 =  x126 &  x240 &  x294 & ~x209 & ~x217;
assign c3174 =  x323 &  x378 &  x548 &  x628 & ~x32;
assign c3176 =  x326 &  x564;
assign c3178 =  x591;
assign c3180 =  x152 & ~x61 & ~x230 & ~x235 & ~x236 & ~x259 & ~x301 & ~x316 & ~x458 & ~x459 & ~x486 & ~x554 & ~x610 & ~x757;
assign c3182 =  x267 &  x627 & ~x301;
assign c3184 =  x208 &  x685 & ~x187 & ~x217 & ~x218 & ~x220 & ~x469 & ~x599 & ~x628;
assign c3186 =  x128 &  x323 & ~x236;
assign c3188 =  x245 &  x327 &  x353 & ~x554 & ~x634 & ~x635 & ~x661 & ~x764;
assign c3190 =  x209 &  x682 & ~x217 & ~x218 & ~x346 & ~x347;
assign c3192 =  x299 &  x326 &  x353 &  x575 & ~x91 & ~x232 & ~x249 & ~x358 & ~x390 & ~x499 & ~x556 & ~x607;
assign c3194 =  x200;
assign c3196 =  x592;
assign c3198 =  x506;
assign c3200 =  x272 &  x327 &  x378 &  x380 & ~x289 & ~x292 & ~x294;
assign c3202 =  x268 &  x323 &  x626 & ~x244 & ~x431 & ~x462;
assign c3204 =  x478;
assign c3206 =  x201;
assign c3208 =  x653 &  x654 & ~x136 & ~x292 & ~x318 & ~x319 & ~x543;
assign c3210 =  x44;
assign c3212 =  x753;
assign c3214 =  x579 &  x635 &  x689;
assign c3216 =  x562;
assign c3218 =  x405 &  x409 &  x551 &  x578 &  x603 &  x604 &  x605 & ~x133;
assign c3220 =  x657 & ~x189 & ~x244 & ~x299 & ~x319 & ~x573;
assign c3222 =  x209 &  x239 &  x295 &  x376 &  x405;
assign c3224 =  x377 &  x435 &  x496 &  x606;
assign c3226 =  x206 & ~x289 & ~x343 & ~x547 & ~x628;
assign c3230 =  x223;
assign c3232 =  x184 &  x235 & ~x319 & ~x320 & ~x374 & ~x545;
assign c3234 =  x228 &  x470;
assign c3236 =  x706;
assign c3238 =  x713;
assign c3240 =  x531;
assign c3242 =  x205 &  x206 &  x578 & ~x289 & ~x312 & ~x335 & ~x340 & ~x344 & ~x511 & ~x694;
assign c3244 =  x657 & ~x262 & ~x263 & ~x288 & ~x573 & ~x599 & ~x600;
assign c3246 =  x180 &  x295 & ~x237 & ~x263 & ~x289 & ~x341;
assign c3248 =  x677;
assign c3250 =  x126 &  x240 &  x293 & ~x431;
assign c3252 =  x657 & ~x160 & ~x191 & ~x219 & ~x263 & ~x264 & ~x510 & ~x567 & ~x571 & ~x573 & ~x610 & ~x716;
assign c3254 =  x11;
assign c3256 =  x196;
assign c3258 =  x377 &  x630 &  x656 & ~x320 & ~x346;
assign c3260 =  x178 &  x659 & ~x102 & ~x263 & ~x287 & ~x506 & ~x637 & ~x721;
assign c3262 =  x214 &  x245 &  x327 &  x379;
assign c3264 =  x216 &  x327 &  x379 &  x380 & ~x486;
assign c3266 =  x215 &  x270 &  x325 &  x548 &  x575 & ~x250 & ~x284 & ~x345 & ~x580 & ~x611;
assign c3268 =  x156 &  x184 &  x521 &  x573 &  x603 &  x628 & ~x161 & ~x688;
assign c3270 =  x243 &  x298 &  x410 &  x628 & ~x492;
assign c3272 =  x122 &  x265;
assign c3274 =  x244 &  x272 &  x299 &  x300 &  x326 &  x353 &  x378 & ~x94 & ~x146 & ~x319 & ~x560;
assign c3276 =  x155 &  x242 &  x269 &  x324 &  x601 & ~x470 & ~x581 & ~x716;
assign c3278 =  x266 &  x411 &  x580 & ~x300;
assign c3280 =  x422;
assign c3282 =  x209 &  x235 &  x240 &  x462 & ~x319 & ~x374 & ~x401 & ~x600;
assign c3284 =  x322 &  x323 & ~x319 & ~x545 & ~x691;
assign c3286 = ~x28 & ~x158 & ~x186 & ~x215 & ~x219 & ~x272 & ~x344 & ~x371 & ~x373 & ~x469 & ~x545 & ~x546 & ~x547 & ~x571 & ~x572 & ~x573 & ~x574 & ~x737;
assign c3288 =  x107;
assign c3290 =  x156 &  x297 &  x323 &  x547 & ~x534 & ~x739;
assign c3292 =  x675;
assign c3294 =  x377 &  x439 &  x497 & ~x244;
assign c3296 =  x658 & ~x32 & ~x237 & ~x263 & ~x290 & ~x487 & ~x573;
assign c3298 =  x194;
assign c31 = ~x2 & ~x17 & ~x19 & ~x20 & ~x31 & ~x40 & ~x45 & ~x101 & ~x144 & ~x148 & ~x172 & ~x222 & ~x269 & ~x280 & ~x337 & ~x394 & ~x409 & ~x425 & ~x437 & ~x465 & ~x475 & ~x592 & ~x644 & ~x649 & ~x678 & ~x710 & ~x717 & ~x726 & ~x730 & ~x734 & ~x747 & ~x763 & ~x780 & ~x781;
assign c33 =  x514 &  x542 & ~x10 & ~x410;
assign c35 =  x516 &  x544 &  x572 & ~x6 & ~x17 & ~x21 & ~x36 & ~x38 & ~x39 & ~x49 & ~x70 & ~x90 & ~x101 & ~x107 & ~x112 & ~x138 & ~x167 & ~x169 & ~x171 & ~x192 & ~x195 & ~x227 & ~x248 & ~x304 & ~x306 & ~x308 & ~x311 & ~x313 & ~x330 & ~x338 & ~x365 & ~x367 & ~x370 & ~x390 & ~x395 & ~x412 & ~x416 & ~x423 & ~x445 & ~x446 & ~x447 & ~x448 & ~x449 & ~x476 & ~x480 & ~x509 & ~x538 & ~x539 & ~x567 & ~x586 & ~x587 & ~x589 & ~x591 & ~x615 & ~x619 & ~x641 & ~x675 & ~x691 & ~x694 & ~x730 & ~x732 & ~x750 & ~x751 & ~x759 & ~x760 & ~x765 & ~x769 & ~x778 & ~x781;
assign c37 =  x489 &  x517 & ~x4 & ~x7 & ~x11 & ~x21 & ~x26 & ~x33 & ~x49 & ~x52 & ~x54 & ~x55 & ~x62 & ~x72 & ~x79 & ~x80 & ~x94 & ~x108 & ~x112 & ~x118 & ~x137 & ~x146 & ~x167 & ~x171 & ~x224 & ~x311 & ~x361 & ~x365 & ~x388 & ~x391 & ~x424 & ~x501 & ~x505 & ~x530 & ~x531 & ~x549 & ~x562 & ~x576 & ~x585 & ~x589 & ~x616 & ~x642 & ~x647 & ~x648 & ~x677 & ~x693 & ~x694 & ~x695 & ~x697 & ~x745 & ~x750 & ~x755 & ~x759 & ~x761 & ~x770;
assign c39 = ~x22 & ~x25 & ~x33 & ~x47 & ~x54 & ~x60 & ~x80 & ~x89 & ~x117 & ~x143 & ~x151 & ~x170 & ~x205 & ~x226 & ~x230 & ~x296 & ~x323 & ~x324 & ~x337 & ~x362 & ~x391 & ~x418 & ~x427 & ~x504 & ~x562 & ~x642 & ~x678 & ~x689 & ~x692 & ~x711 & ~x738 & ~x753 & ~x757 & ~x781;
assign c311 =  x263 &  x291 &  x346 & ~x0 & ~x2 & ~x16 & ~x20 & ~x48 & ~x57 & ~x70 & ~x76 & ~x101 & ~x112 & ~x117 & ~x167 & ~x168 & ~x174 & ~x177 & ~x205 & ~x231 & ~x253 & ~x258 & ~x283 & ~x308 & ~x361 & ~x362 & ~x365 & ~x396 & ~x397 & ~x446 & ~x448 & ~x471 & ~x489 & ~x529 & ~x531 & ~x591 & ~x614 & ~x619 & ~x671 & ~x672 & ~x676 & ~x705 & ~x721 & ~x756 & ~x770 & ~x775;
assign c313 =  x429 &  x430 &  x456 &  x457 & ~x4 & ~x7 & ~x8 & ~x9 & ~x14 & ~x24 & ~x26 & ~x31 & ~x36 & ~x60 & ~x67 & ~x83 & ~x106 & ~x116 & ~x253 & ~x281 & ~x283 & ~x336 & ~x474 & ~x478 & ~x534 & ~x557 & ~x589 & ~x615 & ~x616 & ~x617 & ~x618 & ~x647 & ~x649 & ~x665 & ~x672 & ~x678 & ~x680 & ~x681 & ~x684 & ~x694 & ~x710 & ~x737 & ~x739 & ~x757 & ~x768 & ~x779;
assign c315 =  x437 &  x492 & ~x23 & ~x31 & ~x100 & ~x101 & ~x125 & ~x141 & ~x152 & ~x153 & ~x154 & ~x156 & ~x162 & ~x171 & ~x194 & ~x338 & ~x364 & ~x417 & ~x524 & ~x592 & ~x650 & ~x651 & ~x653 & ~x705 & ~x709 & ~x731 & ~x769 & ~x777 & ~x779;
assign c317 =  x288 &  x372 & ~x489 & ~x620 & ~x751;
assign c319 =  x463 &  x518 &  x572 & ~x221 & ~x336 & ~x348 & ~x376;
assign c321 =  x288 &  x344 &  x373;
assign c323 =  x463 &  x491 &  x518 & ~x5 & ~x7 & ~x14 & ~x18 & ~x22 & ~x25 & ~x44 & ~x48 & ~x54 & ~x59 & ~x70 & ~x80 & ~x81 & ~x87 & ~x90 & ~x111 & ~x144 & ~x160 & ~x173 & ~x218 & ~x221 & ~x222 & ~x249 & ~x277 & ~x279 & ~x283 & ~x302 & ~x331 & ~x333 & ~x357 & ~x362 & ~x387 & ~x449 & ~x476 & ~x527 & ~x587 & ~x593 & ~x620 & ~x623 & ~x624 & ~x651 & ~x652 & ~x654 & ~x672 & ~x678 & ~x681 & ~x705 & ~x709 & ~x715 & ~x723 & ~x725 & ~x728 & ~x745 & ~x747 & ~x756 & ~x769 & ~x771 & ~x783;
assign c325 =  x398 & ~x309;
assign c327 =  x259 &  x314 & ~x112 & ~x393 & ~x677;
assign c329 = ~x100 & ~x165 & ~x353 & ~x380 & ~x408 & ~x409 & ~x436 & ~x465 & ~x616 & ~x725 & ~x732;
assign c331 =  x374 & ~x8 & ~x52 & ~x67 & ~x176 & ~x177 & ~x253 & ~x323 & ~x365 & ~x670 & ~x678 & ~x719;
assign c333 =  x275;
assign c335 = ~x324 & ~x380 & ~x435;
assign c337 =  x431 &  x486 &  x513 &  x514 &  x541 & ~x111 & ~x477 & ~x689 & ~x708 & ~x715;
assign c339 =  x487 &  x515 &  x543 & ~x6 & ~x52 & ~x167 & ~x338 & ~x365 & ~x426 & ~x427 & ~x451 & ~x558 & ~x691 & ~x713 & ~x715 & ~x716 & ~x718 & ~x738 & ~x770;
assign c341 =  x382 &  x437 &  x465 & ~x43 & ~x152 & ~x153 & ~x281 & ~x336 & ~x406 & ~x418 & ~x446 & ~x448 & ~x528 & ~x534 & ~x612 & ~x678 & ~x703 & ~x733;
assign c343 =  x383 & ~x1 & ~x19 & ~x26 & ~x98 & ~x378 & ~x379 & ~x406 & ~x407 & ~x416 & ~x449 & ~x562 & ~x616 & ~x623 & ~x641 & ~x652 & ~x666 & ~x671 & ~x708;
assign c345 = ~x0 & ~x37 & ~x39 & ~x44 & ~x56 & ~x59 & ~x105 & ~x108 & ~x116 & ~x147 & ~x148 & ~x197 & ~x267 & ~x268 & ~x296 & ~x302 & ~x324 & ~x334 & ~x353 & ~x361 & ~x391 & ~x420 & ~x448 & ~x471 & ~x501 & ~x589 & ~x611 & ~x620 & ~x678 & ~x710 & ~x763;
assign c347 =  x320 &  x624 & ~x101 & ~x148 & ~x152 & ~x153 & ~x178 & ~x229 & ~x311 & ~x418 & ~x504 & ~x672 & ~x764;
assign c349 = ~x11 & ~x17 & ~x25 & ~x101 & ~x125 & ~x132 & ~x153 & ~x155 & ~x165 & ~x177 & ~x180 & ~x181 & ~x182 & ~x192 & ~x281 & ~x342 & ~x525 & ~x550 & ~x578 & ~x593 & ~x605 & ~x649 & ~x669 & ~x689 & ~x750 & ~x781;
assign c351 =  x187 & ~x6 & ~x12 & ~x20 & ~x23 & ~x31 & ~x51 & ~x59 & ~x72 & ~x82 & ~x83 & ~x85 & ~x100 & ~x101 & ~x107 & ~x108 & ~x227 & ~x256 & ~x280 & ~x297 & ~x336 & ~x355 & ~x364 & ~x528 & ~x529 & ~x556 & ~x591 & ~x678 & ~x731 & ~x743 & ~x744 & ~x751;
assign c353 =  x218 & ~x20 & ~x98 & ~x311 & ~x361 & ~x449 & ~x589 & ~x644;
assign c355 =  x263 &  x290 &  x318 &  x346 & ~x1 & ~x2 & ~x6 & ~x16 & ~x18 & ~x20 & ~x24 & ~x37 & ~x40 & ~x47 & ~x70 & ~x77 & ~x82 & ~x86 & ~x92 & ~x98 & ~x99 & ~x102 & ~x109 & ~x122 & ~x136 & ~x142 & ~x143 & ~x144 & ~x145 & ~x146 & ~x169 & ~x172 & ~x199 & ~x221 & ~x227 & ~x255 & ~x259 & ~x277 & ~x279 & ~x304 & ~x305 & ~x307 & ~x312 & ~x336 & ~x361 & ~x363 & ~x365 & ~x392 & ~x414 & ~x415 & ~x424 & ~x471 & ~x473 & ~x489 & ~x528 & ~x532 & ~x560 & ~x586 & ~x611 & ~x617 & ~x642 & ~x647 & ~x648 & ~x666 & ~x668 & ~x672 & ~x678 & ~x701 & ~x703 & ~x728 & ~x737 & ~x749 & ~x773 & ~x776;
assign c357 =  x464 &  x492 & ~x10 & ~x45 & ~x46 & ~x51 & ~x73 & ~x100 & ~x107 & ~x126 & ~x133 & ~x225 & ~x256 & ~x279 & ~x365 & ~x392 & ~x397 & ~x507 & ~x551 & ~x565 & ~x592 & ~x595 & ~x624 & ~x644 & ~x655 & ~x678 & ~x679 & ~x681 & ~x703 & ~x710 & ~x724 & ~x740 & ~x749 & ~x763 & ~x765 & ~x781;
assign c359 = ~x14 & ~x26 & ~x80 & ~x141 & ~x143 & ~x170 & ~x280 & ~x308 & ~x323 & ~x336 & ~x350 & ~x351 & ~x376 & ~x377 & ~x378 & ~x392 & ~x404 & ~x405 & ~x406 & ~x559 & ~x589 & ~x668 & ~x669 & ~x671 & ~x672 & ~x703 & ~x712 & ~x719 & ~x754 & ~x776;
assign c361 =  x487 &  x514 &  x542 &  x570;
assign c363 =  x462 &  x518 & ~x31 & ~x113 & ~x146 & ~x170 & ~x325 & ~x391 & ~x424 & ~x534 & ~x653 & ~x678 & ~x679 & ~x687 & ~x692 & ~x712 & ~x731 & ~x738 & ~x766;
assign c365 = ~x9 & ~x108 & ~x153 & ~x156 & ~x182 & ~x377 & ~x378 & ~x642 & ~x757;
assign c367 =  x287 &  x315 &  x343 & ~x2 & ~x7 & ~x21 & ~x31 & ~x36 & ~x45 & ~x48 & ~x54 & ~x60 & ~x75 & ~x86 & ~x89 & ~x108 & ~x123 & ~x307 & ~x335 & ~x336 & ~x364 & ~x389 & ~x418 & ~x446 & ~x447 & ~x560 & ~x593 & ~x614 & ~x620 & ~x622 & ~x641 & ~x678 & ~x679 & ~x702 & ~x721 & ~x730 & ~x750 & ~x759;
assign c369 = ~x60 & ~x131 & ~x152 & ~x153 & ~x154 & ~x156 & ~x181 & ~x182 & ~x210 & ~x395 & ~x418 & ~x559 & ~x578 & ~x692 & ~x728 & ~x765 & ~x783;
assign c371 =  x315 &  x343 &  x371 & ~x224 & ~x781;
assign c373 =  x458 &  x485 &  x512 &  x539 & ~x370;
assign c375 =  x232 & ~x142 & ~x376 & ~x377 & ~x378 & ~x404 & ~x406 & ~x477 & ~x589 & ~x620;
assign c377 = ~x124 & ~x176 & ~x177 & ~x205 & ~x252 & ~x296 & ~x297 & ~x324 & ~x325 & ~x354 & ~x355 & ~x449 & ~x589 & ~x707;
assign c379 = ~x24 & ~x98 & ~x281 & ~x350 & ~x352 & ~x379 & ~x380 & ~x408 & ~x699 & ~x781;
assign c381 = ~x4 & ~x7 & ~x20 & ~x49 & ~x77 & ~x143 & ~x172 & ~x252 & ~x280 & ~x354 & ~x381 & ~x409 & ~x410 & ~x437 & ~x449 & ~x465 & ~x493 & ~x495 & ~x536 & ~x587 & ~x616 & ~x620 & ~x621 & ~x649 & ~x675 & ~x683 & ~x760;
assign c383 =  x372 &  x400 & ~x6 & ~x8 & ~x10 & ~x54 & ~x60 & ~x85 & ~x118 & ~x165 & ~x278 & ~x280 & ~x308 & ~x338 & ~x418 & ~x444 & ~x472 & ~x503 & ~x516 & ~x589 & ~x620 & ~x640 & ~x646 & ~x647 & ~x668 & ~x674 & ~x731 & ~x746 & ~x768 & ~x770 & ~x772 & ~x775;
assign c385 =  x403 &  x431 &  x458 &  x485 &  x513 & ~x22 & ~x36 & ~x169 & ~x196 & ~x340 & ~x424 & ~x452 & ~x587 & ~x644 & ~x731 & ~x736 & ~x738 & ~x745 & ~x754;
assign c387 =  x160 & ~x1 & ~x15 & ~x17 & ~x32 & ~x51 & ~x60 & ~x80 & ~x83 & ~x113 & ~x138 & ~x170 & ~x227 & ~x275 & ~x284 & ~x296 & ~x309 & ~x335 & ~x337 & ~x562 & ~x588 & ~x589 & ~x647 & ~x678 & ~x698 & ~x732 & ~x754 & ~x768 & ~x769;
assign c389 =  x288 &  x316 &  x344 &  x373 & ~x33 & ~x101 & ~x620 & ~x747;
assign c391 =  x153 &  x262 &  x290 & ~x12 & ~x14 & ~x24 & ~x25 & ~x37 & ~x45 & ~x88 & ~x98 & ~x107 & ~x108 & ~x114 & ~x116 & ~x138 & ~x141 & ~x144 & ~x146 & ~x190 & ~x226 & ~x229 & ~x238 & ~x279 & ~x336 & ~x337 & ~x340 & ~x364 & ~x391 & ~x449 & ~x452 & ~x505 & ~x557 & ~x559 & ~x562 & ~x587 & ~x589 & ~x592 & ~x612 & ~x672 & ~x676 & ~x693 & ~x702 & ~x703 & ~x710 & ~x727 & ~x767;
assign c393 =  x345 & ~x8 & ~x17 & ~x22 & ~x116 & ~x267 & ~x268 & ~x269 & ~x279 & ~x302 & ~x393 & ~x395 & ~x424 & ~x449 & ~x534 & ~x678 & ~x754;
assign c395 =  x374 & ~x10 & ~x17 & ~x26 & ~x27 & ~x29 & ~x37 & ~x41 & ~x57 & ~x60 & ~x79 & ~x83 & ~x105 & ~x112 & ~x116 & ~x124 & ~x125 & ~x138 & ~x146 & ~x148 & ~x152 & ~x153 & ~x166 & ~x180 & ~x204 & ~x205 & ~x224 & ~x250 & ~x336 & ~x365 & ~x499 & ~x504 & ~x532 & ~x588 & ~x613 & ~x620 & ~x644 & ~x668 & ~x671 & ~x677 & ~x678 & ~x712 & ~x719 & ~x726 & ~x731 & ~x749 & ~x754 & ~x758 & ~x775 & ~x776;
assign c397 =  x182 & ~x52 & ~x77 & ~x110 & ~x146 & ~x267 & ~x279 & ~x296 & ~x324 & ~x325 & ~x465 & ~x493 & ~x615 & ~x671 & ~x738 & ~x772;
assign c399 =  x436 &  x463 &  x464 &  x491 & ~x26 & ~x64 & ~x192 & ~x279 & ~x280 & ~x350 & ~x361 & ~x378 & ~x590 & ~x649 & ~x682;
assign c3101 =  x517 &  x545 & ~x8 & ~x20 & ~x131 & ~x199 & ~x355 & ~x505 & ~x562 & ~x615 & ~x621 & ~x622 & ~x681 & ~x712;
assign c3103 = ~x0 & ~x8 & ~x26 & ~x59 & ~x79 & ~x89 & ~x98 & ~x146 & ~x152 & ~x153 & ~x172 & ~x193 & ~x205 & ~x228 & ~x279 & ~x336 & ~x361 & ~x391 & ~x395 & ~x420 & ~x494 & ~x495 & ~x496 & ~x524 & ~x534 & ~x550 & ~x551 & ~x578 & ~x590 & ~x591 & ~x592 & ~x593 & ~x620 & ~x647 & ~x649 & ~x651 & ~x691 & ~x749;
assign c3105 =  x460 &  x487 &  x514 &  x542 &  x570 & ~x84 & ~x509;
assign c3107 =  x237 & ~x27 & ~x59 & ~x89 & ~x149 & ~x204 & ~x205 & ~x232 & ~x269 & ~x274 & ~x297 & ~x304 & ~x325 & ~x335 & ~x474 & ~x620 & ~x621 & ~x689 & ~x734;
assign c3109 =  x431 &  x458 &  x486 & ~x170 & ~x226 & ~x286 & ~x424 & ~x660 & ~x707;
assign c3111 =  x436 &  x464 &  x491 & ~x72 & ~x130 & ~x192 & ~x197 & ~x350 & ~x391 & ~x417 & ~x449 & ~x477 & ~x562 & ~x589 & ~x593 & ~x622 & ~x679 & ~x701 & ~x726 & ~x740 & ~x757;
assign c3113 =  x157 & ~x15 & ~x20 & ~x31 & ~x73 & ~x79 & ~x88 & ~x107 & ~x229 & ~x269 & ~x285 & ~x297 & ~x361 & ~x420 & ~x535 & ~x589 & ~x614 & ~x620 & ~x678 & ~x679 & ~x681 & ~x682 & ~x710 & ~x756 & ~x757 & ~x767 & ~x779;
assign c3115 =  x261 &  x289 &  x317 &  x318 & ~x49 & ~x93 & ~x98 & ~x100 & ~x122 & ~x138 & ~x141 & ~x332 & ~x336 & ~x338 & ~x366 & ~x391 & ~x424 & ~x448 & ~x449 & ~x531 & ~x589 & ~x620 & ~x622 & ~x651 & ~x679 & ~x710 & ~x726 & ~x735 & ~x763 & ~x767 & ~x778 & ~x781;
assign c3117 =  x261 &  x289 &  x290 &  x317 & ~x17 & ~x24 & ~x27 & ~x29 & ~x36 & ~x38 & ~x40 & ~x43 & ~x45 & ~x48 & ~x55 & ~x57 & ~x65 & ~x67 & ~x68 & ~x81 & ~x93 & ~x98 & ~x101 & ~x111 & ~x116 & ~x141 & ~x171 & ~x172 & ~x223 & ~x226 & ~x245 & ~x254 & ~x278 & ~x312 & ~x333 & ~x338 & ~x361 & ~x389 & ~x390 & ~x391 & ~x394 & ~x416 & ~x447 & ~x502 & ~x562 & ~x589 & ~x610 & ~x612 & ~x619 & ~x641 & ~x649 & ~x669 & ~x670 & ~x679 & ~x705 & ~x716 & ~x726 & ~x731 & ~x748 & ~x754 & ~x757 & ~x760 & ~x763 & ~x771 & ~x778 & ~x781;
assign c3119 = ~x324 & ~x352 & ~x435;
assign c3121 =  x329 &  x357 & ~x4 & ~x6 & ~x24 & ~x27 & ~x31 & ~x33 & ~x37 & ~x43 & ~x51 & ~x54 & ~x56 & ~x67 & ~x69 & ~x70 & ~x77 & ~x78 & ~x90 & ~x91 & ~x107 & ~x114 & ~x138 & ~x163 & ~x193 & ~x248 & ~x276 & ~x306 & ~x307 & ~x336 & ~x361 & ~x445 & ~x449 & ~x473 & ~x478 & ~x557 & ~x559 & ~x588 & ~x616 & ~x618 & ~x670 & ~x723 & ~x726 & ~x727 & ~x734 & ~x755 & ~x769 & ~x772;
assign c3123 = ~x323 & ~x348 & ~x350 & ~x351 & ~x375 & ~x376 & ~x377 & ~x378 & ~x379 & ~x403 & ~x404 & ~x406 & ~x432 & ~x706;
assign c3125 =  x408 &  x436 &  x464 &  x492 & ~x0 & ~x6 & ~x9 & ~x17 & ~x29 & ~x43 & ~x46 & ~x54 & ~x55 & ~x57 & ~x103 & ~x108 & ~x114 & ~x115 & ~x144 & ~x163 & ~x216 & ~x220 & ~x250 & ~x277 & ~x312 & ~x336 & ~x387 & ~x472 & ~x502 & ~x523 & ~x524 & ~x525 & ~x532 & ~x562 & ~x565 & ~x620 & ~x624 & ~x652 & ~x654 & ~x678 & ~x679 & ~x681 & ~x682 & ~x683 & ~x693 & ~x721 & ~x724 & ~x727 & ~x757 & ~x765;
assign c3127 =  x186 &  x347 & ~x1 & ~x8 & ~x10 & ~x17 & ~x25 & ~x30 & ~x32 & ~x44 & ~x49 & ~x59 & ~x60 & ~x69 & ~x77 & ~x87 & ~x110 & ~x123 & ~x144 & ~x171 & ~x172 & ~x202 & ~x252 & ~x267 & ~x296 & ~x336 & ~x370 & ~x391 & ~x396 & ~x451 & ~x502 & ~x562 & ~x583 & ~x585 & ~x593 & ~x612 & ~x617 & ~x619 & ~x620 & ~x637 & ~x647 & ~x648 & ~x650 & ~x668 & ~x672 & ~x678 & ~x679 & ~x695 & ~x700 & ~x703 & ~x706 & ~x708 & ~x715 & ~x723 & ~x735 & ~x749 & ~x757 & ~x766 & ~x768 & ~x771 & ~x777 & ~x778;
assign c3129 = ~x28 & ~x31 & ~x98 & ~x116 & ~x125 & ~x131 & ~x152 & ~x193 & ~x306 & ~x366 & ~x391 & ~x495 & ~x524 & ~x525 & ~x551 & ~x562 & ~x592 & ~x622 & ~x623 & ~x626 & ~x648 & ~x672 & ~x681 & ~x683 & ~x710 & ~x750 & ~x757 & ~x782;
assign c3131 =  x262 &  x290 &  x318 & ~x1 & ~x7 & ~x17 & ~x22 & ~x26 & ~x41 & ~x48 & ~x60 & ~x66 & ~x83 & ~x107 & ~x108 & ~x119 & ~x120 & ~x141 & ~x146 & ~x171 & ~x172 & ~x197 & ~x223 & ~x225 & ~x226 & ~x251 & ~x268 & ~x279 & ~x280 & ~x281 & ~x283 & ~x286 & ~x337 & ~x338 & ~x361 & ~x370 & ~x392 & ~x398 & ~x421 & ~x424 & ~x426 & ~x446 & ~x449 & ~x583 & ~x590 & ~x592 & ~x615 & ~x619 & ~x637 & ~x643 & ~x664 & ~x671 & ~x672 & ~x691 & ~x712 & ~x725 & ~x744 & ~x747 & ~x754 & ~x757 & ~x759 & ~x773 & ~x775;
assign c3133 =  x431 &  x458 &  x485 &  x486 &  x513 & ~x11 & ~x19 & ~x29 & ~x31 & ~x113 & ~x118 & ~x165 & ~x284 & ~x285 & ~x309 & ~x393 & ~x397 & ~x644 & ~x698 & ~x704 & ~x707 & ~x708 & ~x711;
assign c3135 =  x459 &  x514 &  x570 & ~x37 & ~x59 & ~x138 & ~x426 & ~x616 & ~x771 & ~x776;
assign c3137 =  x486 &  x514 &  x541 & ~x516 & ~x689 & ~x726;
assign c3139 =  x346 &  x402 &  x403 & ~x17 & ~x31 & ~x39 & ~x118 & ~x144 & ~x152 & ~x153 & ~x166 & ~x309 & ~x528 & ~x534;
assign c3141 =  x399 & ~x7 & ~x10 & ~x12 & ~x17 & ~x25 & ~x49 & ~x60 & ~x90 & ~x120 & ~x133 & ~x199 & ~x225 & ~x279 & ~x335 & ~x365 & ~x478 & ~x517 & ~x557 & ~x562 & ~x584 & ~x592 & ~x618 & ~x620 & ~x647 & ~x672 & ~x678 & ~x680 & ~x683 & ~x710 & ~x726 & ~x738 & ~x765 & ~x781;
assign c3143 =  x517 &  x544 &  x572 & ~x8 & ~x22 & ~x32 & ~x38 & ~x43 & ~x77 & ~x90 & ~x100 & ~x101 & ~x108 & ~x116 & ~x219 & ~x251 & ~x278 & ~x337 & ~x338 & ~x387 & ~x392 & ~x393 & ~x418 & ~x424 & ~x441 & ~x444 & ~x502 & ~x505 & ~x507 & ~x535 & ~x586 & ~x592 & ~x596 & ~x621 & ~x670 & ~x675 & ~x678 & ~x695 & ~x706 & ~x717 & ~x747 & ~x761;
assign c3145 =  x488 &  x516 &  x572 & ~x131 & ~x309 & ~x311 & ~x337 & ~x338 & ~x420 & ~x671 & ~x681;
assign c3147 =  x460 &  x487 &  x515 &  x542 & ~x17 & ~x20 & ~x72 & ~x311 & ~x452 & ~x457 & ~x506 & ~x615 & ~x715 & ~x718 & ~x751 & ~x761;
assign c3149 =  x431 &  x485 &  x512 & ~x4 & ~x9 & ~x11 & ~x53 & ~x106 & ~x253 & ~x286 & ~x534 & ~x560 & ~x562 & ~x644 & ~x703 & ~x741 & ~x757 & ~x759;
assign c3151 =  x379 &  x463 &  x518 & ~x1 & ~x2 & ~x17 & ~x33 & ~x50 & ~x53 & ~x56 & ~x79 & ~x91 & ~x106 & ~x116 & ~x171 & ~x193 & ~x200 & ~x227 & ~x248 & ~x255 & ~x278 & ~x279 & ~x281 & ~x304 & ~x336 & ~x338 & ~x365 & ~x395 & ~x416 & ~x449 & ~x474 & ~x509 & ~x535 & ~x557 & ~x565 & ~x566 & ~x569 & ~x584 & ~x587 & ~x593 & ~x595 & ~x616 & ~x619 & ~x620 & ~x623 & ~x641 & ~x642 & ~x649 & ~x672 & ~x678 & ~x679 & ~x689 & ~x694 & ~x699 & ~x716 & ~x726 & ~x727 & ~x744 & ~x757 & ~x760 & ~x763 & ~x767 & ~x769 & ~x781;
assign c3153 =  x358;
assign c3155 = ~x31 & ~x41 & ~x90 & ~x98 & ~x101 & ~x193 & ~x350 & ~x361 & ~x376 & ~x377 & ~x378 & ~x404 & ~x474 & ~x559 & ~x655 & ~x672 & ~x678 & ~x682 & ~x703 & ~x711;
assign c3157 =  x409 &  x437 &  x464 &  x465 &  x492 & ~x10 & ~x17 & ~x20 & ~x29 & ~x48 & ~x64 & ~x71 & ~x76 & ~x77 & ~x100 & ~x109 & ~x112 & ~x132 & ~x139 & ~x143 & ~x167 & ~x169 & ~x197 & ~x199 & ~x221 & ~x247 & ~x276 & ~x280 & ~x308 & ~x338 & ~x350 & ~x385 & ~x395 & ~x416 & ~x417 & ~x418 & ~x419 & ~x420 & ~x423 & ~x448 & ~x449 & ~x500 & ~x504 & ~x592 & ~x595 & ~x623 & ~x624 & ~x668 & ~x672 & ~x678 & ~x697 & ~x707 & ~x709 & ~x751 & ~x752 & ~x755 & ~x759 & ~x776;
assign c3159 =  x488 &  x543 &  x570 & ~x20 & ~x73 & ~x119 & ~x166 & ~x365 & ~x392 & ~x425 & ~x439 & ~x693;
assign c3161 = ~x6 & ~x12 & ~x20 & ~x43 & ~x44 & ~x48 & ~x49 & ~x90 & ~x108 & ~x142 & ~x173 & ~x213 & ~x216 & ~x225 & ~x238 & ~x239 & ~x240 & ~x241 & ~x248 & ~x268 & ~x269 & ~x275 & ~x333 & ~x336 & ~x392 & ~x418 & ~x421 & ~x424 & ~x530 & ~x531 & ~x562 & ~x590 & ~x617 & ~x620 & ~x623 & ~x647 & ~x650 & ~x652 & ~x667 & ~x672 & ~x679 & ~x766 & ~x770;
assign c3163 =  x491 &  x546 & ~x79 & ~x133 & ~x156 & ~x197 & ~x305 & ~x366 & ~x395 & ~x420 & ~x449 & ~x534 & ~x592 & ~x616 & ~x621 & ~x624 & ~x634 & ~x651 & ~x681 & ~x703 & ~x722 & ~x726;
assign c3165 =  x454 &  x455 & ~x14 & ~x26 & ~x78 & ~x80 & ~x90 & ~x146 & ~x164 & ~x200 & ~x219 & ~x220 & ~x228 & ~x254 & ~x306 & ~x337 & ~x367 & ~x392 & ~x449 & ~x450 & ~x589 & ~x644 & ~x671 & ~x672 & ~x703 & ~x710 & ~x711 & ~x732 & ~x744 & ~x776;
assign c3167 = ~x6 & ~x116 & ~x349 & ~x350 & ~x376 & ~x377 & ~x378 & ~x403 & ~x404 & ~x406 & ~x434 & ~x535 & ~x595 & ~x622 & ~x678;
assign c3169 =  x431 &  x458 &  x485 &  x513 &  x540;
assign c3171 =  x517 &  x544 & ~x8 & ~x14 & ~x24 & ~x32 & ~x60 & ~x73 & ~x101 & ~x110 & ~x144 & ~x228 & ~x280 & ~x365 & ~x391 & ~x424 & ~x447 & ~x449 & ~x534 & ~x589 & ~x590 & ~x591 & ~x615 & ~x631 & ~x633 & ~x646 & ~x672 & ~x691 & ~x740 & ~x751 & ~x762;
assign c3173 =  x543 &  x570 & ~x170 & ~x350 & ~x419 & ~x557 & ~x672 & ~x726 & ~x729;
assign c3175 =  x259 &  x287 &  x315 & ~x247 & ~x279 & ~x365 & ~x391 & ~x564 & ~x589 & ~x675 & ~x678 & ~x726 & ~x781;
assign c3177 =  x464 &  x492 & ~x17 & ~x19 & ~x20 & ~x45 & ~x61 & ~x89 & ~x98 & ~x125 & ~x143 & ~x166 & ~x176 & ~x223 & ~x307 & ~x365 & ~x525 & ~x551 & ~x555 & ~x565 & ~x619 & ~x620 & ~x624 & ~x644 & ~x650 & ~x652 & ~x654 & ~x655 & ~x670 & ~x678 & ~x679 & ~x683 & ~x709 & ~x747 & ~x780;
assign c3179 =  x291 &  x346 &  x374 &  x402 &  x403 & ~x205 & ~x418 & ~x674;
assign c3181 =  x491 &  x518 &  x546 & ~x19 & ~x31 & ~x33 & ~x34 & ~x39 & ~x47 & ~x54 & ~x77 & ~x131 & ~x132 & ~x170 & ~x172 & ~x197 & ~x215 & ~x223 & ~x226 & ~x305 & ~x334 & ~x424 & ~x453 & ~x472 & ~x505 & ~x510 & ~x534 & ~x586 & ~x590 & ~x606 & ~x620 & ~x623 & ~x634 & ~x636 & ~x649 & ~x651 & ~x668 & ~x672 & ~x678 & ~x693 & ~x694 & ~x722 & ~x726 & ~x744 & ~x766 & ~x771;
assign c3183 =  x431 &  x458 &  x485 &  x540;
assign c3185 =  x427 &  x455 & ~x6 & ~x7 & ~x22 & ~x24 & ~x47 & ~x72 & ~x73 & ~x105 & ~x116 & ~x139 & ~x193 & ~x279 & ~x282 & ~x309 & ~x335 & ~x338 & ~x390 & ~x391 & ~x392 & ~x395 & ~x418 & ~x452 & ~x531 & ~x557 & ~x562 & ~x590 & ~x617 & ~x731 & ~x744 & ~x757 & ~x763 & ~x765 & ~x766;
assign c3187 =  x461 &  x488 &  x516 &  x543 &  x570 & ~x63 & ~x588;
assign c3189 = ~x11 & ~x25 & ~x43 & ~x64 & ~x96 & ~x144 & ~x148 & ~x170 & ~x195 & ~x225 & ~x266 & ~x278 & ~x280 & ~x296 & ~x297 & ~x323 & ~x324 & ~x367 & ~x424 & ~x502 & ~x589 & ~x591 & ~x615 & ~x616 & ~x620 & ~x622 & ~x647 & ~x651 & ~x667 & ~x672 & ~x678 & ~x679 & ~x713 & ~x726 & ~x731 & ~x734 & ~x759 & ~x763;
assign c3191 =  x263 &  x291 & ~x0 & ~x4 & ~x7 & ~x10 & ~x12 & ~x14 & ~x17 & ~x20 & ~x22 & ~x24 & ~x27 & ~x31 & ~x34 & ~x40 & ~x41 & ~x43 & ~x47 & ~x54 & ~x57 & ~x60 & ~x67 & ~x70 & ~x79 & ~x82 & ~x86 & ~x91 & ~x93 & ~x98 & ~x102 & ~x103 & ~x107 & ~x113 & ~x116 & ~x118 & ~x120 & ~x132 & ~x148 & ~x164 & ~x166 & ~x171 & ~x177 & ~x192 & ~x193 & ~x223 & ~x224 & ~x228 & ~x230 & ~x248 & ~x250 & ~x279 & ~x283 & ~x284 & ~x309 & ~x312 & ~x332 & ~x335 & ~x336 & ~x340 & ~x343 & ~x361 & ~x365 & ~x366 & ~x367 & ~x384 & ~x386 & ~x388 & ~x391 & ~x392 & ~x396 & ~x397 & ~x418 & ~x421 & ~x424 & ~x426 & ~x445 & ~x449 & ~x450 & ~x474 & ~x499 & ~x509 & ~x525 & ~x528 & ~x552 & ~x588 & ~x593 & ~x608 & ~x610 & ~x614 & ~x620 & ~x622 & ~x649 & ~x663 & ~x666 & ~x667 & ~x668 & ~x671 & ~x672 & ~x674 & ~x678 & ~x679 & ~x694 & ~x699 & ~x701 & ~x703 & ~x719 & ~x733 & ~x735 & ~x746 & ~x750 & ~x751 & ~x755 & ~x757 & ~x759 & ~x760 & ~x763 & ~x765 & ~x767 & ~x769 & ~x776 & ~x780 & ~x782;
assign c3193 =  x461 &  x516 &  x544 &  x572 & ~x37 & ~x89 & ~x107 & ~x192 & ~x198 & ~x221 & ~x343 & ~x412 & ~x535 & ~x592 & ~x649 & ~x727 & ~x752 & ~x758;
assign c3195 =  x459 &  x486 &  x513 & ~x2 & ~x7 & ~x13 & ~x19 & ~x21 & ~x24 & ~x26 & ~x28 & ~x38 & ~x44 & ~x45 & ~x47 & ~x57 & ~x59 & ~x62 & ~x69 & ~x73 & ~x79 & ~x81 & ~x86 & ~x87 & ~x105 & ~x136 & ~x193 & ~x194 & ~x225 & ~x253 & ~x278 & ~x280 & ~x284 & ~x305 & ~x308 & ~x310 & ~x334 & ~x335 & ~x343 & ~x361 & ~x363 & ~x365 & ~x367 & ~x369 & ~x393 & ~x418 & ~x421 & ~x423 & ~x447 & ~x448 & ~x449 & ~x475 & ~x506 & ~x532 & ~x534 & ~x560 & ~x562 & ~x587 & ~x588 & ~x589 & ~x590 & ~x613 & ~x617 & ~x667 & ~x668 & ~x674 & ~x675 & ~x687 & ~x688 & ~x689 & ~x693 & ~x702 & ~x705 & ~x710 & ~x719 & ~x725 & ~x726 & ~x734 & ~x735 & ~x744 & ~x745 & ~x755 & ~x779;
assign c3197 =  x344 &  x372 &  x400 & ~x7 & ~x10 & ~x14 & ~x22 & ~x31 & ~x43 & ~x60 & ~x138 & ~x166 & ~x200 & ~x391 & ~x416 & ~x449 & ~x474 & ~x726 & ~x765 & ~x782;
assign c3199 =  x517 &  x544 &  x572 & ~x7 & ~x8 & ~x11 & ~x21 & ~x46 & ~x57 & ~x64 & ~x79 & ~x85 & ~x89 & ~x109 & ~x118 & ~x135 & ~x141 & ~x146 & ~x172 & ~x195 & ~x226 & ~x227 & ~x278 & ~x283 & ~x307 & ~x335 & ~x340 & ~x361 & ~x391 & ~x397 & ~x418 & ~x422 & ~x424 & ~x444 & ~x448 & ~x449 & ~x502 & ~x509 & ~x535 & ~x565 & ~x585 & ~x590 & ~x591 & ~x593 & ~x649 & ~x678 & ~x703 & ~x725 & ~x726 & ~x738 & ~x744 & ~x746 & ~x751 & ~x763;
assign c3201 =  x248;
assign c3203 =  x358;
assign c3205 =  x233 & ~x27 & ~x81 & ~x82 & ~x168 & ~x280 & ~x350 & ~x376 & ~x377 & ~x402 & ~x404 & ~x406 & ~x420 & ~x776;
assign c3207 =  x289 & ~x117 & ~x152 & ~x183;
assign c3209 =  x489 &  x517 &  x544 &  x572 & ~x0 & ~x4 & ~x7 & ~x17 & ~x24 & ~x25 & ~x37 & ~x43 & ~x79 & ~x89 & ~x90 & ~x104 & ~x107 & ~x111 & ~x115 & ~x121 & ~x142 & ~x193 & ~x228 & ~x248 & ~x283 & ~x314 & ~x336 & ~x361 & ~x366 & ~x370 & ~x392 & ~x416 & ~x423 & ~x505 & ~x509 & ~x532 & ~x535 & ~x536 & ~x589 & ~x591 & ~x648 & ~x726 & ~x730 & ~x744 & ~x745 & ~x749 & ~x763 & ~x764 & ~x769;
assign c3211 =  x516 &  x571 & ~x6 & ~x8 & ~x41 & ~x59 & ~x281 & ~x457 & ~x467 & ~x567 & ~x729 & ~x743;
assign c3213 =  x435 & ~x98 & ~x155 & ~x493 & ~x550 & ~x576 & ~x577 & ~x674 & ~x687 & ~x703;
assign c3215 =  x290 &  x345 &  x373 &  x401 & ~x672;
assign c3217 =  x369;
assign c3219 =  x461 &  x488 &  x516 &  x543 &  x571 & ~x79 & ~x448 & ~x468 & ~x700 & ~x770;
assign c3221 =  x486 &  x514 &  x541 & ~x19 & ~x24 & ~x89 & ~x107 & ~x227 & ~x282 & ~x365 & ~x420 & ~x428 & ~x439 & ~x589 & ~x643 & ~x690 & ~x692 & ~x701 & ~x751 & ~x773 & ~x774;
assign c3225 =  x263 &  x290 &  x291 &  x318 &  x346 &  x347 & ~x0 & ~x4 & ~x11 & ~x14 & ~x20 & ~x35 & ~x45 & ~x63 & ~x95 & ~x100 & ~x121 & ~x143 & ~x146 & ~x171 & ~x172 & ~x226 & ~x231 & ~x259 & ~x280 & ~x281 & ~x283 & ~x304 & ~x330 & ~x390 & ~x442 & ~x561 & ~x591 & ~x609 & ~x615 & ~x616 & ~x643 & ~x647 & ~x672 & ~x713 & ~x745 & ~x748 & ~x755 & ~x778;
assign c3227 = ~x20 & ~x24 & ~x26 & ~x28 & ~x54 & ~x57 & ~x90 & ~x146 & ~x194 & ~x223 & ~x248 & ~x268 & ~x296 & ~x306 & ~x307 & ~x311 & ~x340 & ~x352 & ~x380 & ~x478 & ~x532 & ~x590 & ~x615 & ~x644 & ~x645 & ~x678 & ~x704 & ~x714 & ~x727 & ~x732 & ~x746 & ~x750 & ~x757 & ~x761 & ~x762 & ~x781;
assign c3229 =  x490 & ~x297 & ~x353 & ~x361 & ~x381 & ~x437 & ~x533 & ~x679 & ~x680 & ~x682 & ~x707 & ~x708 & ~x745 & ~x746;
assign c3231 =  x429 &  x430 &  x457 &  x485 & ~x33 & ~x61 & ~x75 & ~x108 & ~x169 & ~x195 & ~x228 & ~x506 & ~x650 & ~x693 & ~x699 & ~x710 & ~x762;
assign c3233 =  x487 &  x542 & ~x0 & ~x2 & ~x9 & ~x22 & ~x25 & ~x26 & ~x29 & ~x33 & ~x49 & ~x66 & ~x84 & ~x141 & ~x192 & ~x226 & ~x250 & ~x276 & ~x278 & ~x302 & ~x304 & ~x305 & ~x336 & ~x340 & ~x361 & ~x364 & ~x392 & ~x393 & ~x425 & ~x448 & ~x531 & ~x589 & ~x642 & ~x666 & ~x667 & ~x668 & ~x672 & ~x687 & ~x690 & ~x712 & ~x716 & ~x718 & ~x726 & ~x734 & ~x744 & ~x751 & ~x762 & ~x777 & ~x781;
assign c3235 =  x407 &  x433 &  x461 &  x488 &  x516 &  x543 & ~x2 & ~x22 & ~x27 & ~x29 & ~x34 & ~x37 & ~x39 & ~x43 & ~x45 & ~x57 & ~x61 & ~x81 & ~x82 & ~x105 & ~x114 & ~x135 & ~x137 & ~x143 & ~x146 & ~x172 & ~x195 & ~x247 & ~x279 & ~x335 & ~x356 & ~x361 & ~x363 & ~x448 & ~x449 & ~x452 & ~x617 & ~x619 & ~x641 & ~x644 & ~x669 & ~x672 & ~x705 & ~x708 & ~x719 & ~x722 & ~x748 & ~x753 & ~x766 & ~x773 & ~x781;
assign c3237 =  x457 &  x484 &  x567 & ~x397;
assign c3239 =  x487 &  x515 &  x542 & ~x24 & ~x61 & ~x410 & ~x412 & ~x757;
assign c3241 = ~x14 & ~x24 & ~x102 & ~x168 & ~x281 & ~x353 & ~x381 & ~x409 & ~x436 & ~x464 & ~x465 & ~x615 & ~x671 & ~x697 & ~x698 & ~x703 & ~x715;
assign c3243 = ~x2 & ~x5 & ~x7 & ~x9 & ~x10 & ~x15 & ~x30 & ~x31 & ~x32 & ~x37 & ~x39 & ~x43 & ~x51 & ~x57 & ~x60 & ~x68 & ~x74 & ~x108 & ~x113 & ~x117 & ~x138 & ~x163 & ~x167 & ~x171 & ~x172 & ~x193 & ~x199 & ~x223 & ~x225 & ~x249 & ~x283 & ~x304 & ~x307 & ~x309 & ~x320 & ~x334 & ~x340 & ~x348 & ~x349 & ~x350 & ~x365 & ~x376 & ~x377 & ~x378 & ~x387 & ~x391 & ~x421 & ~x422 & ~x449 & ~x472 & ~x502 & ~x504 & ~x505 & ~x534 & ~x560 & ~x589 & ~x591 & ~x640 & ~x642 & ~x643 & ~x647 & ~x668 & ~x682 & ~x686 & ~x687 & ~x689 & ~x694 & ~x695 & ~x699 & ~x709 & ~x711 & ~x718 & ~x729 & ~x730 & ~x731 & ~x734 & ~x748 & ~x751 & ~x763 & ~x764 & ~x780;
assign c3245 =  x461 &  x515 &  x570 & ~x54 & ~x60 & ~x446 & ~x452 & ~x715;
assign c3247 = ~x24 & ~x75 & ~x94 & ~x97 & ~x152 & ~x153 & ~x180 & ~x181 & ~x408 & ~x502 & ~x507 & ~x516 & ~x531 & ~x699 & ~x756;
assign c3249 =  x315 &  x372 & ~x14 & ~x37 & ~x141 & ~x279 & ~x417 & ~x449 & ~x532 & ~x592 & ~x644 & ~x672 & ~x751 & ~x753 & ~x765;
assign c3251 =  x261 &  x289 &  x317 &  x345 &  x374 & ~x10 & ~x12 & ~x20 & ~x38 & ~x75 & ~x79 & ~x100 & ~x117 & ~x146 & ~x167 & ~x172 & ~x199 & ~x225 & ~x228 & ~x257 & ~x279 & ~x307 & ~x391 & ~x447 & ~x557 & ~x559 & ~x562 & ~x591 & ~x670 & ~x678 & ~x726 & ~x729 & ~x740 & ~x776;
assign c3253 =  x607 &  x608 &  x609 & ~x256 & ~x364 & ~x648 & ~x737;
assign c3255 =  x288 &  x316 & ~x28 & ~x34 & ~x48 & ~x70 & ~x78 & ~x79 & ~x98 & ~x102 & ~x105 & ~x141 & ~x142 & ~x143 & ~x167 & ~x192 & ~x223 & ~x225 & ~x280 & ~x336 & ~x390 & ~x393 & ~x423 & ~x488 & ~x489 & ~x490 & ~x534 & ~x584 & ~x614 & ~x619 & ~x649 & ~x672 & ~x697 & ~x703 & ~x725 & ~x731 & ~x760;
assign c3257 = ~x100 & ~x251 & ~x354 & ~x403 & ~x409 & ~x412 & ~x437 & ~x465 & ~x466 & ~x496 & ~x522 & ~x678 & ~x775 & ~x781;
assign c3259 =  x347 & ~x4 & ~x11 & ~x114 & ~x132 & ~x152 & ~x205 & ~x278 & ~x284 & ~x307 & ~x336 & ~x340 & ~x361 & ~x416 & ~x418 & ~x448 & ~x495 & ~x525 & ~x551 & ~x562 & ~x620 & ~x720 & ~x752 & ~x769;
assign c3261 = ~x20 & ~x89 & ~x96 & ~x103 & ~x116 & ~x241 & ~x253 & ~x269 & ~x392 & ~x437 & ~x438 & ~x440 & ~x465 & ~x477 & ~x617 & ~x667 & ~x712 & ~x714 & ~x717 & ~x719 & ~x725 & ~x746;
assign c3263 =  x522 & ~x16 & ~x19 & ~x20 & ~x24 & ~x36 & ~x49 & ~x64 & ~x79 & ~x91 & ~x115 & ~x143 & ~x193 & ~x194 & ~x281 & ~x323 & ~x324 & ~x351 & ~x352 & ~x361 & ~x389 & ~x391 & ~x418 & ~x503 & ~x534 & ~x679 & ~x681 & ~x732 & ~x734 & ~x738 & ~x750 & ~x762 & ~x763;
assign c3265 = ~x7 & ~x8 & ~x29 & ~x49 & ~x53 & ~x96 & ~x98 & ~x100 & ~x112 & ~x137 & ~x146 & ~x152 & ~x170 & ~x180 & ~x339 & ~x495 & ~x496 & ~x500 & ~x504 & ~x524 & ~x538 & ~x550 & ~x566 & ~x577 & ~x578 & ~x580 & ~x587 & ~x593 & ~x605 & ~x615 & ~x621 & ~x622 & ~x623 & ~x708 & ~x719 & ~x732 & ~x733 & ~x776;
assign c3267 =  x288 &  x316 &  x344 &  x373 & ~x87 & ~x449;
assign c3269 =  x426 & ~x2 & ~x33 & ~x38 & ~x40 & ~x59 & ~x66 & ~x78 & ~x116 & ~x137 & ~x143 & ~x170 & ~x336 & ~x364 & ~x394 & ~x473 & ~x531 & ~x616 & ~x672 & ~x678 & ~x679 & ~x711 & ~x763 & ~x781;
assign c3271 =  x260 & ~x7 & ~x19 & ~x20 & ~x31 & ~x54 & ~x77 & ~x78 & ~x104 & ~x113 & ~x119 & ~x139 & ~x144 & ~x146 & ~x166 & ~x210 & ~x249 & ~x362 & ~x392 & ~x477 & ~x504 & ~x508 & ~x557 & ~x620 & ~x645 & ~x703 & ~x722 & ~x729 & ~x732;
assign c3273 =  x437 &  x465 &  x492 & ~x15 & ~x70 & ~x109 & ~x182 & ~x334 & ~x499 & ~x593 & ~x594 & ~x679 & ~x763;
assign c3275 = ~x0 & ~x7 & ~x10 & ~x20 & ~x27 & ~x40 & ~x47 & ~x77 & ~x78 & ~x80 & ~x83 & ~x86 & ~x95 & ~x96 & ~x110 & ~x115 & ~x166 & ~x167 & ~x170 & ~x172 & ~x173 & ~x197 & ~x200 & ~x278 & ~x279 & ~x280 & ~x284 & ~x294 & ~x303 & ~x312 & ~x323 & ~x334 & ~x336 & ~x338 & ~x351 & ~x360 & ~x369 & ~x391 & ~x392 & ~x393 & ~x424 & ~x448 & ~x449 & ~x502 & ~x534 & ~x562 & ~x589 & ~x591 & ~x592 & ~x619 & ~x620 & ~x647 & ~x648 & ~x649 & ~x660 & ~x661 & ~x668 & ~x672 & ~x674 & ~x675 & ~x678 & ~x679 & ~x689 & ~x694 & ~x695 & ~x698 & ~x699 & ~x705 & ~x707 & ~x716 & ~x732 & ~x735 & ~x744 & ~x748 & ~x750 & ~x751 & ~x778;
assign c3277 =  x487 &  x542 & ~x0 & ~x18 & ~x31 & ~x55 & ~x80 & ~x104 & ~x110 & ~x114 & ~x280 & ~x307 & ~x412 & ~x427 & ~x453 & ~x561 & ~x589 & ~x702 & ~x705 & ~x717 & ~x743 & ~x766;
assign c3279 = ~x86 & ~x91 & ~x103 & ~x132 & ~x152 & ~x176 & ~x177 & ~x279 & ~x308 & ~x381 & ~x382 & ~x409 & ~x410 & ~x437 & ~x642 & ~x672 & ~x782;
assign c3281 =  x317 &  x345 &  x373 &  x401 & ~x107 & ~x121 & ~x228 & ~x336 & ~x669 & ~x747 & ~x771;
assign c3283 =  x492 &  x546 & ~x3 & ~x11 & ~x12 & ~x20 & ~x31 & ~x76 & ~x101 & ~x323 & ~x351 & ~x388 & ~x557 & ~x562 & ~x589 & ~x612 & ~x616 & ~x617 & ~x646 & ~x687 & ~x695 & ~x754 & ~x777;
assign c3285 =  x436 &  x463 &  x464 &  x491 & ~x10 & ~x59 & ~x109 & ~x116 & ~x131 & ~x133 & ~x247 & ~x312 & ~x314 & ~x370 & ~x451 & ~x481 & ~x524 & ~x537 & ~x540 & ~x550 & ~x562 & ~x622 & ~x623 & ~x624 & ~x652 & ~x693 & ~x751 & ~x775;
assign c3287 = ~x0 & ~x4 & ~x6 & ~x10 & ~x20 & ~x26 & ~x36 & ~x43 & ~x45 & ~x49 & ~x90 & ~x112 & ~x148 & ~x164 & ~x173 & ~x198 & ~x200 & ~x202 & ~x217 & ~x220 & ~x239 & ~x240 & ~x254 & ~x267 & ~x268 & ~x269 & ~x278 & ~x280 & ~x281 & ~x309 & ~x363 & ~x418 & ~x421 & ~x565 & ~x592 & ~x619 & ~x620 & ~x622 & ~x640 & ~x652 & ~x672 & ~x681 & ~x682 & ~x707 & ~x726 & ~x771;
assign c3289 =  x428 &  x429 & ~x3 & ~x20 & ~x25 & ~x26 & ~x59 & ~x113 & ~x169 & ~x172 & ~x228 & ~x312 & ~x392 & ~x424 & ~x448 & ~x505 & ~x530 & ~x535 & ~x562 & ~x586 & ~x589 & ~x614 & ~x619 & ~x642 & ~x649 & ~x650 & ~x652 & ~x655 & ~x656 & ~x668 & ~x672 & ~x673 & ~x678 & ~x681 & ~x682 & ~x724 & ~x781 & ~x782;
assign c3291 =  x431 &  x459 &  x486 & ~x18 & ~x25 & ~x32 & ~x40 & ~x62 & ~x72 & ~x77 & ~x107 & ~x116 & ~x165 & ~x225 & ~x306 & ~x340 & ~x393 & ~x395 & ~x419 & ~x474 & ~x477 & ~x478 & ~x516 & ~x534 & ~x536 & ~x650 & ~x674 & ~x678 & ~x692 & ~x708 & ~x709 & ~x725 & ~x726 & ~x741;
assign c3293 =  x317 &  x318 &  x345 &  x346 &  x374 & ~x8 & ~x12 & ~x14 & ~x19 & ~x20 & ~x66 & ~x74 & ~x90 & ~x98 & ~x103 & ~x106 & ~x113 & ~x117 & ~x123 & ~x125 & ~x148 & ~x229 & ~x278 & ~x279 & ~x284 & ~x306 & ~x307 & ~x310 & ~x332 & ~x336 & ~x338 & ~x361 & ~x365 & ~x366 & ~x474 & ~x477 & ~x505 & ~x557 & ~x619 & ~x648 & ~x669 & ~x670 & ~x675 & ~x703 & ~x726 & ~x732 & ~x745 & ~x751 & ~x757 & ~x763 & ~x775 & ~x777;
assign c3295 =  x463 &  x491 &  x518 &  x546 & ~x6 & ~x20 & ~x25 & ~x60 & ~x130 & ~x301 & ~x306 & ~x338 & ~x414 & ~x509 & ~x560 & ~x586 & ~x620 & ~x622 & ~x623 & ~x626 & ~x654 & ~x673 & ~x678 & ~x702 & ~x773 & ~x778;
assign c3297 =  x182 & ~x10 & ~x11 & ~x82 & ~x98 & ~x121 & ~x140 & ~x172 & ~x228 & ~x267 & ~x268 & ~x269 & ~x277 & ~x296 & ~x297 & ~x304 & ~x324 & ~x325 & ~x328 & ~x360 & ~x562 & ~x617 & ~x672 & ~x746 & ~x751;
assign c3299 =  x463 &  x518 & ~x24 & ~x152 & ~x225 & ~x281 & ~x451 & ~x550 & ~x577 & ~x592 & ~x605 & ~x622 & ~x635 & ~x668 & ~x678 & ~x769;
assign c40 =  x411 & ~x209 & ~x238 & ~x548 & ~x562 & ~x575 & ~x602 & ~x603;
assign c42 =  x777;
assign c44 =  x490 &  x491 & ~x139 & ~x155 & ~x237 & ~x507 & ~x548 & ~x550 & ~x576 & ~x577 & ~x625 & ~x766;
assign c46 =  x381 &  x465 & ~x224 & ~x236 & ~x327 & ~x516 & ~x598;
assign c48 =  x534;
assign c410 =  x409 &  x432 &  x436 & ~x208 & ~x236 & ~x328 & ~x595 & ~x602;
assign c412 =  x300 &  x383 &  x411 & ~x212 & ~x224 & ~x307 & ~x352;
assign c414 =  x431 &  x432 & ~x100 & ~x211 & ~x351 & ~x378 & ~x379 & ~x514 & ~x544 & ~x621 & ~x627;
assign c416 =  x344 &  x372 &  x401 & ~x153 & ~x236 & ~x384;
assign c418 =  x642;
assign c420 =  x140;
assign c422 =  x296 &  x324 &  x380 &  x408 & ~x118 & ~x208 & ~x247 & ~x281 & ~x327 & ~x337 & ~x369 & ~x394 & ~x481 & ~x500 & ~x551 & ~x623 & ~x655 & ~x775;
assign c424 =  x478;
assign c426 =  x326 &  x381 &  x402 &  x403 &  x464 & ~x157 & ~x267 & ~x481 & ~x550;
assign c428 =  x352 &  x380 &  x463 &  x491 & ~x62 & ~x76 & ~x127 & ~x143 & ~x196 & ~x239 & ~x327 & ~x515 & ~x539 & ~x543 & ~x549 & ~x598 & ~x759 & ~x781;
assign c430 =  x399 & ~x27 & ~x208 & ~x236 & ~x377 & ~x572 & ~x575 & ~x602;
assign c432 =  x17;
assign c434 =  x438 & ~x209 & ~x351 & ~x519 & ~x547 & ~x602 & ~x713;
assign c436 =  x299 &  x327 &  x383 & ~x56 & ~x69 & ~x82 & ~x105 & ~x240 & ~x268 & ~x294 & ~x324 & ~x479 & ~x567 & ~x598 & ~x680 & ~x725 & ~x746 & ~x758 & ~x775;
assign c438 =  x354 &  x381 &  x437 & ~x38 & ~x83 & ~x119 & ~x184 & ~x224 & ~x258 & ~x268 & ~x389 & ~x445 & ~x541 & ~x571 & ~x586 & ~x613 & ~x628 & ~x708 & ~x716 & ~x719 & ~x721 & ~x746 & ~x777;
assign c440 =  x431 &  x432 &  x437 &  x438 &  x439 & ~x486;
assign c442 =  x768;
assign c444 =  x300 &  x327 &  x354 &  x355 &  x382 &  x437 & ~x1 & ~x7 & ~x24 & ~x40 & ~x52 & ~x58 & ~x88 & ~x90 & ~x114 & ~x124 & ~x125 & ~x128 & ~x137 & ~x186 & ~x241 & ~x253 & ~x284 & ~x296 & ~x313 & ~x332 & ~x359 & ~x420 & ~x422 & ~x473 & ~x475 & ~x478 & ~x506 & ~x508 & ~x528 & ~x537 & ~x556 & ~x564 & ~x615 & ~x635 & ~x637 & ~x640 & ~x670 & ~x690 & ~x708 & ~x721 & ~x734 & ~x745 & ~x748 & ~x754 & ~x759 & ~x776;
assign c446 =  x320 &  x354 &  x376 &  x518 & ~x127 & ~x388;
assign c448 =  x319 &  x352 &  x428 & ~x327;
assign c450 =  x271 &  x353 &  x354 &  x381 & ~x241 & ~x577;
assign c452 =  x372 &  x494 & ~x237 & ~x267 & ~x293 & ~x320 & ~x378 & ~x656;
assign c454 =  x487 &  x488 &  x490 &  x491 &  x494 &  x520 & ~x46 & ~x82 & ~x107 & ~x378 & ~x406 & ~x418 & ~x621 & ~x648 & ~x714 & ~x719;
assign c456 =  x292 &  x320 &  x324 &  x352 &  x407 & ~x288 & ~x354;
assign c458 =  x320 &  x347 &  x490 & ~x548 & ~x576;
assign c460 =  x29;
assign c462 =  x300 &  x355 &  x410 & ~x214 & ~x298 & ~x352 & ~x568;
assign c464 =  x46 &  x168;
assign c466 =  x346 &  x405 &  x465 &  x492 & ~x213 & ~x269 & ~x511 & ~x577 & ~x606;
assign c468 =  x347 &  x352 &  x461 & ~x575;
assign c470 =  x397 &  x425 & ~x359;
assign c472 =  x459 &  x460 & ~x324 & ~x352 & ~x379 & ~x514 & ~x544 & ~x626 & ~x747;
assign c474 =  x456 &  x487 &  x488 &  x490 & ~x171 & ~x433 & ~x627;
assign c476 =  x338;
assign c478 =  x296 &  x324 &  x352 &  x408 &  x491 &  x519 &  x520 & ~x63 & ~x204 & ~x216 & ~x259 & ~x309 & ~x327 & ~x585;
assign c480 =  x401 &  x402 &  x411 &  x429 &  x431 &  x432 &  x437 & ~x12 & ~x88 & ~x139 & ~x175 & ~x220 & ~x285 & ~x311 & ~x390 & ~x421 & ~x445 & ~x469 & ~x510 & ~x514 & ~x590 & ~x621 & ~x647 & ~x650 & ~x692 & ~x697 & ~x722 & ~x758;
assign c482 =  x399 &  x427 &  x432 &  x439 & ~x192 & ~x514 & ~x654 & ~x655 & ~x744 & ~x752;
assign c484 =  x345 &  x401 &  x490 & ~x577;
assign c486 =  x375 &  x404 &  x491 & ~x215 & ~x515 & ~x521;
assign c488 =  x325 &  x375 &  x381 &  x404 &  x437 & ~x199;
assign c490 =  x451 &  x730;
assign c492 =  x245 &  x383 & ~x213 & ~x215;
assign c494 =  x346 &  x400 &  x429 & ~x259 & ~x333 & ~x576 & ~x577 & ~x587 & ~x764;
assign c496 =  x320 &  x352 &  x462 & ~x575;
assign c498 =  x381 &  x437 &  x465 & ~x208 & ~x236 & ~x247 & ~x602;
assign c4100 =  x490 & ~x129 & ~x213 & ~x294 & ~x359 & ~x392 & ~x541 & ~x548 & ~x549 & ~x576 & ~x605;
assign c4102 =  x456 &  x466 & ~x212 & ~x268 & ~x352 & ~x406;
assign c4104 =  x246 & ~x95 & ~x188 & ~x269 & ~x295 & ~x337 & ~x688;
assign c4106 =  x325 &  x381 &  x484 &  x491 & ~x179 & ~x623 & ~x680 & ~x705 & ~x710 & ~x752 & ~x773;
assign c4110 =  x320 &  x348 &  x375 &  x465 &  x490 & ~x175 & ~x261 & ~x313 & ~x342 & ~x443 & ~x478 & ~x571 & ~x621 & ~x642 & ~x770;
assign c4112 =  x379 &  x402 &  x490 & ~x247 & ~x327 & ~x577;
assign c4114 =  x326 &  x354 &  x374 &  x402 &  x456 & ~x329 & ~x378;
assign c4116 =  x320 &  x325 &  x381 &  x403 &  x431 & ~x262 & ~x599;
assign c4118 =  x317 &  x372 &  x400 &  x401 & ~x185 & ~x286;
assign c4120 =  x346 &  x354 &  x374 &  x401 &  x429 &  x437 & ~x602;
assign c4122 =  x484 &  x513 &  x516 &  x517 & ~x130 & ~x367 & ~x393 & ~x404 & ~x406 & ~x433;
assign c4124 =  x7 &  x139;
assign c4126 =  x455 &  x483 &  x484 &  x485 & ~x209 & ~x405 & ~x559 & ~x565 & ~x626 & ~x671 & ~x711;
assign c4128 =  x325 &  x381 &  x437 &  x520 & ~x41 & ~x50 & ~x105 & ~x237 & ~x285 & ~x311 & ~x526 & ~x567 & ~x568 & ~x572 & ~x580 & ~x591 & ~x598 & ~x600 & ~x627 & ~x655 & ~x767;
assign c4130 =  x516 &  x599 &  x654;
assign c4132 =  x398 & ~x236 & ~x295;
assign c4134 =  x435 & ~x107 & ~x210 & ~x220 & ~x258 & ~x272 & ~x486 & ~x487 & ~x493 & ~x521 & ~x523 & ~x541 & ~x549;
assign c4136 =  x347 &  x429 &  x437 &  x458 &  x459 &  x463 & ~x40 & ~x46 & ~x106 & ~x260 & ~x315 & ~x587 & ~x588 & ~x598 & ~x701 & ~x728 & ~x741 & ~x768;
assign c4138 =  x516 &  x599 & ~x157;
assign c4140 =  x667;
assign c4142 =  x326 &  x381 &  x430 &  x431 &  x437 & ~x24 & ~x197 & ~x210 & ~x396 & ~x497 & ~x510 & ~x513 & ~x585 & ~x740;
assign c4144 =  x382 &  x403 &  x405 &  x406 &  x409 &  x548 & ~x75 & ~x150 & ~x202 & ~x231 & ~x387 & ~x388 & ~x485 & ~x500 & ~x513 & ~x514 & ~x528 & ~x618 & ~x709 & ~x744;
assign c4146 =  x365;
assign c4148 =  x327 &  x382 &  x430 &  x431 & ~x241 & ~x626;
assign c4150 =  x319 &  x374 &  x400 &  x429 &  x491 & ~x288 & ~x328 & ~x378;
assign c4152 =  x403 &  x408 & ~x186 & ~x485 & ~x575 & ~x602;
assign c4154 =  x113;
assign c4156 =  x487 & ~x81 & ~x111 & ~x207 & ~x405 & ~x406 & ~x433 & ~x602 & ~x740;
assign c4158 =  x326 &  x520 &  x521 & ~x231 & ~x288 & ~x379 & ~x406 & ~x625;
assign c4160 =  x404 &  x408 & ~x208 & ~x236 & ~x515 & ~x550 & ~x566 & ~x622;
assign c4162 =  x766;
assign c4164 =  x703;
assign c4166 =  x434 &  x438 & ~x259 & ~x260 & ~x326 & ~x521;
assign c4168 =  x475;
assign c4170 =  x671;
assign c4174 =  x381 &  x491 & ~x2 & ~x53 & ~x107 & ~x172 & ~x213 & ~x239 & ~x252 & ~x268 & ~x445 & ~x452 & ~x508 & ~x511 & ~x521 & ~x577 & ~x585 & ~x592;
assign c4176 =  x344 &  x454;
assign c4178 =  x279;
assign c4180 =  x11;
assign c4182 =  x484 & ~x261 & ~x405 & ~x406 & ~x433 & ~x727;
assign c4184 =  x295 &  x351 &  x379 &  x434 &  x463 &  x491 &  x547 & ~x99 & ~x326 & ~x580 & ~x749 & ~x783;
assign c4186 =  x494 &  x578 & ~x210 & ~x237 & ~x602 & ~x629 & ~x657;
assign c4188 =  x318 &  x374 &  x405 &  x438 &  x492 & ~x74 & ~x83 & ~x514;
assign c4190 =  x324 &  x352 &  x491 & ~x167 & ~x181 & ~x218 & ~x237 & ~x247 & ~x303 & ~x327 & ~x529 & ~x541 & ~x606 & ~x655;
assign c4192 =  x296 &  x352 &  x430 & ~x300 & ~x326 & ~x329;
assign c4194 =  x346 &  x354 &  x381 &  x403 & ~x351;
assign c4196 =  x224;
assign c4198 =  x396;
assign c4200 =  x301 & ~x214 & ~x298;
assign c4202 =  x113;
assign c4204 =  x33;
assign c4206 =  x348 &  x375 &  x464 &  x465 &  x491 &  x492 &  x520 &  x548 & ~x103 & ~x140 & ~x206 & ~x246 & ~x332 & ~x775;
assign c4208 =  x465 &  x520 &  x661 & ~x206 & ~x327;
assign c4210 =  x345 &  x399 & ~x81 & ~x327 & ~x391 & ~x509 & ~x571 & ~x597 & ~x626 & ~x710;
assign c4212 =  x406 & ~x519 & ~x521 & ~x548 & ~x575;
assign c4214 =  x324 &  x347 &  x352 &  x380 &  x407 & ~x140 & ~x300 & ~x568;
assign c4216 =  x49;
assign c4218 =  x216 &  x299 & ~x140 & ~x184 & ~x199 & ~x268 & ~x294 & ~x359 & ~x626 & ~x680;
assign c4220 =  x398 &  x454 &  x459;
assign c4222 =  x728;
assign c4224 =  x700;
assign c4226 =  x491 &  x494 &  x631 & ~x327 & ~x598;
assign c4228 =  x379 &  x459 &  x462 &  x490 & ~x150 & ~x286 & ~x299 & ~x326;
assign c4230 =  x344 &  x352 &  x373 &  x488 &  x490 & ~x95 & ~x302;
assign c4232 =  x430 &  x431 &  x432 & ~x56 & ~x65 & ~x139 & ~x229 & ~x255 & ~x259 & ~x420 & ~x472 & ~x481 & ~x515 & ~x573 & ~x627 & ~x665 & ~x673 & ~x683 & ~x741 & ~x760 & ~x766;
assign c4234 =  x346 &  x374 &  x402 & ~x66 & ~x109 & ~x121 & ~x140 & ~x501 & ~x575 & ~x602 & ~x684 & ~x687 & ~x708 & ~x722;
assign c4236 =  x343 &  x371 &  x399 &  x465 & ~x141 & ~x236 & ~x443 & ~x508 & ~x526 & ~x626 & ~x720 & ~x721 & ~x781;
assign c4238 =  x344 &  x371 &  x430 &  x431 & ~x61 & ~x336;
assign c4240 =  x520 &  x662;
assign c4242 =  x429 &  x491 &  x517 & ~x260 & ~x405 & ~x433 & ~x584;
assign c4244 =  x375 &  x382 &  x402 &  x429 & ~x379;
assign c4246 =  x115;
assign c4248 =  x381 &  x490 &  x517 & ~x576;
assign c4250 =  x381 &  x400 &  x401 &  x429 & ~x53 & ~x209 & ~x541 & ~x572 & ~x598;
assign c4252 =  x246 &  x456 & ~x187;
assign c4254 =  x325 &  x456 & ~x218 & ~x327;
assign c4256 =  x673;
assign c4258 =  x324 &  x345 &  x352 &  x408 & ~x65 & ~x92 & ~x96 & ~x124 & ~x182 & ~x183 & ~x209 & ~x224 & ~x237 & ~x256 & ~x453 & ~x474 & ~x476 & ~x540 & ~x542 & ~x553 & ~x710 & ~x720 & ~x725 & ~x773 & ~x775;
assign c4260 =  x189 & ~x405;
assign c4262 =  x381 &  x402 & ~x572 & ~x599 & ~x602 & ~x658;
assign c4264 =  x589;
assign c4266 =  x163;
assign c4268 =  x320 &  x352 &  x375 &  x403 &  x490 &  x491 & ~x606;
assign c4270 =  x345 &  x352 & ~x327;
assign c4272 =  x352 &  x380 &  x464 &  x465 &  x520 & ~x31 & ~x57 & ~x60 & ~x72 & ~x84 & ~x98 & ~x111 & ~x131 & ~x162 & ~x168 & ~x275 & ~x307 & ~x364 & ~x383 & ~x423 & ~x523 & ~x525 & ~x555 & ~x597 & ~x688 & ~x745;
assign c4274 =  x488 &  x494 &  x518 &  x520 & ~x56 & ~x365 & ~x405 & ~x571 & ~x639 & ~x740;
assign c4276 =  x318 &  x377 & ~x127 & ~x128 & ~x521 & ~x525 & ~x603 & ~x633 & ~x688;
assign c4278 =  x327 &  x410 &  x465 & ~x185 & ~x240 & ~x268 & ~x341 & ~x352 & ~x477 & ~x706;
assign c4280 =  x352 &  x463 &  x464 &  x491 & ~x1 & ~x14 & ~x88 & ~x140 & ~x148 & ~x272 & ~x326 & ~x327 & ~x510 & ~x541 & ~x543 & ~x568 & ~x597 & ~x601 & ~x714 & ~x742;
assign c4282 =  x346 &  x401 &  x460 &  x465 &  x489 &  x490 &  x491 & ~x259 & ~x541;
assign c4284 =  x320 &  x347 &  x402 &  x457 & ~x331 & ~x405;
assign c4286 =  x347 &  x381 & ~x324 & ~x542 & ~x577;
assign c4288 =  x351 &  x374 &  x402 &  x434 &  x490 & ~x188 & ~x204 & ~x215 & ~x244 & ~x272 & ~x550;
assign c4290 =  x438 & ~x209 & ~x357 & ~x377 & ~x405 & ~x602 & ~x626;
assign c4292 =  x318 &  x346 &  x352 & ~x209 & ~x237 & ~x257 & ~x550;
assign c4296 =  x562;
assign c4298 =  x323 &  x375 &  x379 &  x406 & ~x327 & ~x424;
assign c41 =  x153 &  x154 & ~x21 & ~x674;
assign c43 =  x210 &  x211 &  x212 &  x236 & ~x5 & ~x8 & ~x10 & ~x12 & ~x18 & ~x40 & ~x43 & ~x51 & ~x57 & ~x58 & ~x59 & ~x60 & ~x81 & ~x82 & ~x97 & ~x106 & ~x121 & ~x125 & ~x144 & ~x166 & ~x167 & ~x168 & ~x202 & ~x220 & ~x226 & ~x246 & ~x257 & ~x340 & ~x362 & ~x386 & ~x413 & ~x426 & ~x445 & ~x454 & ~x468 & ~x478 & ~x527 & ~x580 & ~x596 & ~x614 & ~x620 & ~x637 & ~x674 & ~x681 & ~x701 & ~x726 & ~x747 & ~x776;
assign c45 = ~x408 & ~x410 & ~x437 & ~x619 & ~x665;
assign c47 =  x97;
assign c49 =  x183 &  x184 &  x656 &  x657 & ~x43 & ~x97 & ~x100 & ~x194 & ~x284 & ~x529;
assign c411 =  x209 &  x211 &  x212 &  x235 & ~x20 & ~x199 & ~x225 & ~x307 & ~x310 & ~x594 & ~x650;
assign c413 =  x182 &  x183 &  x184 &  x208 & ~x0 & ~x82 & ~x199 & ~x292 & ~x310 & ~x477 & ~x735;
assign c415 =  x542 &  x570 &  x571 & ~x273 & ~x368 & ~x421 & ~x659 & ~x735;
assign c417 =  x625 &  x626 & ~x488 & ~x668;
assign c419 =  x125 &  x544;
assign c421 =  x128;
assign c423 =  x266 &  x269 & ~x65 & ~x94 & ~x100 & ~x102 & ~x104 & ~x187 & ~x367 & ~x388 & ~x449 & ~x460 & ~x532 & ~x641 & ~x720 & ~x724 & ~x777;
assign c425 =  x235 &  x236 &  x238 &  x239 & ~x3 & ~x16 & ~x21 & ~x43 & ~x48 & ~x57 & ~x58 & ~x59 & ~x65 & ~x89 & ~x126 & ~x135 & ~x153 & ~x228 & ~x281 & ~x421 & ~x449 & ~x499 & ~x562 & ~x565 & ~x591 & ~x613 & ~x615 & ~x619 & ~x651 & ~x677 & ~x681 & ~x730 & ~x740 & ~x782;
assign c427 =  x151;
assign c429 =  x294 & ~x3 & ~x20 & ~x52 & ~x118 & ~x160 & ~x169 & ~x173 & ~x283 & ~x334 & ~x364 & ~x416 & ~x435 & ~x480 & ~x504 & ~x535 & ~x584 & ~x670 & ~x707 & ~x733 & ~x739 & ~x763 & ~x779;
assign c431 =  x180 &  x181 &  x182 &  x183 & ~x21 & ~x36 & ~x42 & ~x130 & ~x138 & ~x192 & ~x279 & ~x292 & ~x532;
assign c433 =  x567 & ~x263;
assign c435 =  x542 &  x543 &  x544 &  x570 & ~x271;
assign c437 =  x127 &  x154 & ~x49 & ~x106 & ~x144 & ~x363 & ~x682 & ~x709 & ~x783;
assign c439 = ~x75 & ~x132 & ~x137 & ~x168 & ~x225 & ~x284 & ~x311 & ~x365 & ~x409 & ~x410 & ~x436 & ~x437 & ~x438 & ~x465 & ~x529 & ~x559 & ~x586 & ~x641 & ~x698 & ~x703 & ~x706 & ~x781;
assign c441 =  x238 &  x239 &  x240 & ~x20 & ~x22 & ~x68 & ~x119 & ~x126 & ~x153 & ~x155 & ~x160 & ~x227 & ~x307 & ~x336 & ~x348 & ~x442 & ~x571 & ~x641 & ~x642 & ~x725 & ~x756 & ~x758 & ~x764;
assign c443 =  x541 &  x570 &  x571 & ~x160 & ~x251 & ~x332 & ~x421 & ~x587;
assign c445 =  x265 &  x266 &  x291 & ~x6 & ~x29 & ~x54 & ~x103 & ~x106 & ~x134 & ~x164 & ~x169 & ~x175 & ~x179 & ~x184 & ~x199 & ~x204 & ~x305 & ~x335 & ~x370 & ~x388 & ~x412 & ~x413 & ~x480 & ~x496 & ~x561 & ~x569 & ~x586 & ~x595 & ~x610 & ~x640 & ~x644 & ~x664 & ~x701 & ~x733 & ~x763 & ~x773;
assign c447 = ~x18 & ~x36 & ~x84 & ~x192 & ~x221 & ~x283 & ~x310 & ~x425 & ~x462 & ~x463 & ~x480 & ~x492 & ~x512 & ~x567 & ~x614 & ~x615 & ~x639 & ~x691 & ~x719 & ~x754;
assign c449 =  x211 &  x235 &  x236 & ~x284 & ~x292 & ~x415 & ~x571 & ~x701;
assign c451 =  x595;
assign c453 =  x542 &  x543 &  x545 &  x571 & ~x297 & ~x308 & ~x311;
assign c455 =  x238 &  x239 &  x240 &  x241 &  x242 & ~x88 & ~x280;
assign c457 =  x236 &  x238 &  x239 &  x240 & ~x32 & ~x96 & ~x251 & ~x276 & ~x312 & ~x362 & ~x397 & ~x413 & ~x425 & ~x477 & ~x497 & ~x499 & ~x559 & ~x589 & ~x668 & ~x760;
assign c459 =  x184 &  x185 &  x214 &  x215 & ~x37 & ~x60 & ~x81 & ~x196 & ~x268 & ~x281 & ~x314 & ~x446 & ~x502 & ~x503 & ~x611 & ~x669 & ~x727 & ~x753;
assign c461 =  x207 &  x208 &  x211 & ~x18 & ~x69 & ~x84 & ~x123 & ~x191 & ~x251 & ~x281 & ~x307 & ~x320 & ~x532 & ~x562 & ~x619 & ~x761;
assign c463 =  x123;
assign c465 =  x539 & ~x263 & ~x308 & ~x316 & ~x344;
assign c467 = ~x144 & ~x372 & ~x373 & ~x376 & ~x400 & ~x401 & ~x402 & ~x429 & ~x752;
assign c469 = ~x372 & ~x401 & ~x402 & ~x412 & ~x492;
assign c471 =  x294 & ~x106 & ~x155 & ~x159 & ~x176 & ~x187 & ~x228 & ~x308 & ~x333 & ~x420 & ~x421 & ~x429 & ~x430 & ~x476 & ~x532 & ~x559 & ~x590 & ~x619 & ~x644 & ~x694 & ~x774;
assign c473 =  x567 & ~x287;
assign c475 =  x235 &  x236 &  x238 &  x262 & ~x6 & ~x56 & ~x67 & ~x83 & ~x99 & ~x251 & ~x333 & ~x504 & ~x556 & ~x763;
assign c477 =  x239 &  x241 &  x265 &  x291 & ~x496;
assign c479 =  x241 &  x266 &  x267 & ~x153 & ~x161 & ~x308 & ~x310 & ~x333 & ~x415 & ~x442 & ~x503 & ~x504 & ~x532 & ~x589 & ~x615 & ~x619 & ~x637 & ~x664 & ~x777;
assign c481 =  x235 &  x236 &  x237 &  x238 &  x239 & ~x53 & ~x419 & ~x559 & ~x595;
assign c483 =  x187 &  x625;
assign c485 =  x211 &  x212 & ~x22 & ~x320 & ~x375 & ~x397 & ~x414 & ~x415 & ~x586 & ~x619;
assign c487 =  x322 & ~x18 & ~x33 & ~x59 & ~x61 & ~x76 & ~x91 & ~x111 & ~x139 & ~x222 & ~x335 & ~x392 & ~x435 & ~x504 & ~x529 & ~x560 & ~x589 & ~x614 & ~x615 & ~x637 & ~x643 & ~x673 & ~x694 & ~x701 & ~x760 & ~x777;
assign c489 = ~x69 & ~x373 & ~x376 & ~x400 & ~x401 & ~x402 & ~x403 & ~x430;
assign c491 =  x433 & ~x144 & ~x202 & ~x335 & ~x341 & ~x344 & ~x382 & ~x409 & ~x410 & ~x438 & ~x639 & ~x647 & ~x693;
assign c493 =  x266 &  x267 & ~x15 & ~x19 & ~x22 & ~x40 & ~x85 & ~x112 & ~x116 & ~x118 & ~x122 & ~x127 & ~x129 & ~x143 & ~x155 & ~x161 & ~x196 & ~x221 & ~x280 & ~x308 & ~x335 & ~x338 & ~x375 & ~x387 & ~x424 & ~x498 & ~x502 & ~x508 & ~x586 & ~x589 & ~x593 & ~x610 & ~x617 & ~x637 & ~x640 & ~x672 & ~x677 & ~x693 & ~x695 & ~x703 & ~x722 & ~x750 & ~x761 & ~x762 & ~x764 & ~x769 & ~x770 & ~x782;
assign c495 =  x515 &  x543 &  x544 &  x545 &  x573 & ~x186 & ~x270 & ~x283 & ~x659 & ~x701;
assign c497 =  x441 &  x544 & ~x49 & ~x144 & ~x161 & ~x256 & ~x615 & ~x628 & ~x637 & ~x659 & ~x777;
assign c499 =  x211 &  x212 & ~x61 & ~x109 & ~x135 & ~x151 & ~x153 & ~x163 & ~x206 & ~x316 & ~x343 & ~x362 & ~x438 & ~x498 & ~x532 & ~x725 & ~x732;
assign c4101 =  x183 &  x184 &  x628 &  x629 & ~x3 & ~x24 & ~x450 & ~x507 & ~x649;
assign c4103 =  x212 &  x214 &  x238 & ~x25 & ~x31 & ~x34 & ~x36 & ~x41 & ~x43 & ~x138 & ~x363 & ~x525 & ~x617 & ~x619 & ~x659 & ~x730 & ~x768;
assign c4105 =  x525 & ~x43 & ~x160 & ~x161 & ~x164 & ~x218 & ~x476 & ~x643 & ~x723;
assign c4107 =  x209 &  x211 &  x235 &  x236 &  x240 & ~x504;
assign c4109 =  x433 & ~x230 & ~x252 & ~x357 & ~x409 & ~x410 & ~x437 & ~x438;
assign c4111 =  x205 &  x206 &  x207 & ~x3 & ~x13 & ~x81 & ~x161 & ~x274 & ~x310 & ~x318 & ~x346 & ~x566 & ~x649 & ~x735 & ~x749 & ~x765;
assign c4113 =  x233 &  x498 & ~x226 & ~x702;
assign c4115 =  x211 &  x214 &  x236 & ~x153 & ~x169 & ~x415 & ~x770;
assign c4117 =  x265 &  x266 &  x290 &  x291 & ~x88 & ~x106 & ~x159 & ~x183 & ~x192 & ~x202 & ~x251 & ~x566;
assign c4119 =  x294 &  x297 & ~x363 & ~x459 & ~x460 & ~x694 & ~x749;
assign c4121 =  x573 & ~x22 & ~x59 & ~x286 & ~x334 & ~x341 & ~x353 & ~x381 & ~x419 & ~x448 & ~x657 & ~x686 & ~x687;
assign c4123 =  x238 &  x239 & ~x3 & ~x23 & ~x32 & ~x85 & ~x86 & ~x148 & ~x387 & ~x421 & ~x462 & ~x479 & ~x488 & ~x586 & ~x732;
assign c4125 =  x100;
assign c4127 =  x657 &  x660 & ~x574;
assign c4129 =  x97;
assign c4131 =  x262 &  x293 &  x294;
assign c4133 =  x240 &  x241 &  x266 &  x291 & ~x115 & ~x162 & ~x182 & ~x476 & ~x557 & ~x698 & ~x701 & ~x756 & ~x762;
assign c4135 =  x265 &  x266 &  x268 & ~x5 & ~x79 & ~x157 & ~x251 & ~x337 & ~x460 & ~x613 & ~x754;
assign c4137 =  x602 &  x604 & ~x381;
assign c4139 =  x128 & ~x69 & ~x86 & ~x141 & ~x143 & ~x250 & ~x268 & ~x305 & ~x306 & ~x310 & ~x333 & ~x369 & ~x418 & ~x420 & ~x447 & ~x476 & ~x477 & ~x530 & ~x559 & ~x561 & ~x610 & ~x640 & ~x644 & ~x673 & ~x701 & ~x712 & ~x763;
assign c4141 =  x210 &  x211 &  x236 &  x263 & ~x3 & ~x10 & ~x14 & ~x17 & ~x24 & ~x43 & ~x46 & ~x49 & ~x84 & ~x87 & ~x93 & ~x97 & ~x116 & ~x117 & ~x120 & ~x132 & ~x136 & ~x138 & ~x142 & ~x150 & ~x153 & ~x159 & ~x160 & ~x190 & ~x294 & ~x322 & ~x332 & ~x363 & ~x367 & ~x369 & ~x370 & ~x391 & ~x395 & ~x412 & ~x440 & ~x473 & ~x476 & ~x480 & ~x496 & ~x506 & ~x511 & ~x527 & ~x559 & ~x563 & ~x580 & ~x595 & ~x598 & ~x614 & ~x615 & ~x620 & ~x644 & ~x677 & ~x738 & ~x750 & ~x767 & ~x773 & ~x781;
assign c4143 =  x213 &  x214 &  x215 &  x238 &  x239 & ~x251 & ~x469;
assign c4145 =  x567;
assign c4147 = ~x88 & ~x92 & ~x100 & ~x222 & ~x375 & ~x402 & ~x428 & ~x429 & ~x448 & ~x454 & ~x694 & ~x699 & ~x727;
assign c4149 =  x214 &  x215 &  x239 &  x240 & ~x152;
assign c4151 =  x604 & ~x3 & ~x16 & ~x49 & ~x88 & ~x144 & ~x171 & ~x251 & ~x335 & ~x338 & ~x454 & ~x492 & ~x563 & ~x610 & ~x620 & ~x674 & ~x725;
assign c4153 =  x180 &  x181 &  x182 &  x183 & ~x0 & ~x82 & ~x88 & ~x97 & ~x132 & ~x165 & ~x171 & ~x201 & ~x202 & ~x219 & ~x292 & ~x308 & ~x499 & ~x532 & ~x589 & ~x640 & ~x723 & ~x730 & ~x757 & ~x775;
assign c4155 =  x657 & ~x8 & ~x16 & ~x84 & ~x281 & ~x397 & ~x398 & ~x414 & ~x483 & ~x490 & ~x644 & ~x672 & ~x730 & ~x750 & ~x754 & ~x757 & ~x778;
assign c4157 =  x266 &  x291 & ~x16 & ~x24 & ~x30 & ~x42 & ~x43 & ~x44 & ~x91 & ~x99 & ~x104 & ~x138 & ~x155 & ~x184 & ~x190 & ~x308 & ~x310 & ~x362 & ~x389 & ~x415 & ~x475 & ~x476 & ~x500 & ~x530 & ~x589 & ~x640 & ~x644 & ~x662 & ~x668 & ~x693 & ~x702 & ~x717 & ~x778 & ~x782;
assign c4159 =  x632 & ~x36 & ~x97 & ~x251 & ~x363 & ~x492 & ~x520 & ~x585 & ~x757;
assign c4161 = ~x21 & ~x283 & ~x374 & ~x375 & ~x402 & ~x430 & ~x431 & ~x459 & ~x488 & ~x581 & ~x610 & ~x698;
assign c4163 = ~x5 & ~x9 & ~x13 & ~x24 & ~x34 & ~x35 & ~x57 & ~x70 & ~x103 & ~x137 & ~x162 & ~x313 & ~x318 & ~x356 & ~x367 & ~x372 & ~x385 & ~x420 & ~x429 & ~x430 & ~x431 & ~x458 & ~x593 & ~x644 & ~x648 & ~x668 & ~x760;
assign c4165 =  x543 &  x571 &  x573 & ~x246 & ~x270;
assign c4167 =  x182 &  x183 &  x184 &  x185 & ~x5 & ~x6 & ~x22 & ~x58 & ~x76 & ~x88 & ~x142 & ~x173 & ~x201 & ~x219 & ~x251 & ~x256 & ~x308 & ~x321 & ~x421 & ~x446 & ~x448 & ~x525 & ~x638 & ~x672 & ~x696 & ~x697 & ~x751 & ~x761;
assign c4169 =  x597 &  x598 & ~x7 & ~x235 & ~x415 & ~x679;
assign c4171 = ~x44 & ~x55 & ~x77 & ~x164 & ~x195 & ~x203 & ~x219 & ~x229 & ~x277 & ~x318 & ~x344 & ~x345 & ~x372 & ~x373 & ~x421 & ~x430 & ~x648 & ~x701 & ~x729 & ~x731 & ~x761 & ~x778 & ~x779;
assign c4173 =  x622;
assign c4175 =  x571 &  x572 &  x573 & ~x35 & ~x192 & ~x270 & ~x283 & ~x335 & ~x418 & ~x561 & ~x644 & ~x677 & ~x701 & ~x770 & ~x782;
assign c4177 =  x542 &  x570 & ~x400 & ~x652 & ~x730;
assign c4179 =  x211 &  x628 & ~x730;
assign c4181 = ~x408 & ~x409 & ~x410 & ~x437;
assign c4183 =  x628 & ~x7 & ~x16 & ~x18 & ~x169 & ~x248 & ~x364 & ~x476 & ~x490 & ~x508 & ~x641 & ~x668 & ~x706 & ~x708 & ~x722 & ~x730;
assign c4185 =  x573 &  x574 & ~x13 & ~x77 & ~x91 & ~x107 & ~x177 & ~x231 & ~x301 & ~x308 & ~x314 & ~x316 & ~x317 & ~x331 & ~x338 & ~x343 & ~x344 & ~x359 & ~x372 & ~x387 & ~x389 & ~x400 & ~x428 & ~x448 & ~x503 & ~x659 & ~x674 & ~x694 & ~x702 & ~x721 & ~x739 & ~x749 & ~x779;
assign c4187 =  x238 &  x239 &  x240 &  x241 &  x242 & ~x13 & ~x15 & ~x64 & ~x68 & ~x138 & ~x172 & ~x255 & ~x421 & ~x533 & ~x560 & ~x564 & ~x588 & ~x619 & ~x673 & ~x729 & ~x756;
assign c4189 =  x153 &  x154 &  x179 & ~x192 & ~x760;
assign c4191 =  x208 &  x211 &  x212 &  x235 &  x236;
assign c4193 =  x542 & ~x344 & ~x637 & ~x754;
assign c4195 =  x239 &  x240 &  x241 &  x265 & ~x415 & ~x468 & ~x619;
assign c4197 =  x543 & ~x11 & ~x40 & ~x57 & ~x88 & ~x173 & ~x194 & ~x219 & ~x226 & ~x251 & ~x284 & ~x338 & ~x362 & ~x372 & ~x398 & ~x399 & ~x400 & ~x415 & ~x532 & ~x615 & ~x640 & ~x659 & ~x682 & ~x701 & ~x730;
assign c4199 =  x183 &  x184 &  x185 &  x186 & ~x20 & ~x45 & ~x64 & ~x68 & ~x73 & ~x79 & ~x82 & ~x90 & ~x93 & ~x115 & ~x137 & ~x283 & ~x284 & ~x309 & ~x310 & ~x334 & ~x342 & ~x363 & ~x395 & ~x414 & ~x415 & ~x477 & ~x482 & ~x525 & ~x557 & ~x610 & ~x639 & ~x640 & ~x644 & ~x671 & ~x691 & ~x725 & ~x735 & ~x751 & ~x763 & ~x778;
assign c4201 =  x180 &  x181 &  x182 &  x183 & ~x3 & ~x17 & ~x18 & ~x35 & ~x50 & ~x69 & ~x75 & ~x82 & ~x106 & ~x108 & ~x109 & ~x144 & ~x169 & ~x198 & ~x226 & ~x252 & ~x276 & ~x283 & ~x306 & ~x307 & ~x336 & ~x356 & ~x362 & ~x363 & ~x483 & ~x511 & ~x532 & ~x557 & ~x561 & ~x617 & ~x644 & ~x711 & ~x730 & ~x749 & ~x774;
assign c4203 =  x211 &  x236 &  x263 & ~x69 & ~x279 & ~x305 & ~x342 & ~x348 & ~x385 & ~x439 & ~x440 & ~x467 & ~x483 & ~x499 & ~x525 & ~x723 & ~x730 & ~x775;
assign c4205 = ~x408 & ~x409 & ~x437 & ~x438;
assign c4207 =  x209 &  x211 &  x212 &  x325 & ~x15 & ~x34 & ~x43 & ~x47 & ~x54 & ~x81 & ~x84 & ~x96 & ~x98 & ~x106 & ~x115 & ~x129 & ~x152 & ~x157 & ~x162 & ~x164 & ~x178 & ~x199 & ~x228 & ~x308 & ~x310 & ~x313 & ~x329 & ~x337 & ~x363 & ~x393 & ~x397 & ~x398 & ~x399 & ~x439 & ~x446 & ~x455 & ~x467 & ~x480 & ~x495 & ~x529 & ~x555 & ~x557 & ~x564 & ~x571 & ~x581 & ~x589 & ~x596 & ~x642 & ~x643 & ~x663 & ~x668 & ~x691 & ~x700 & ~x720 & ~x726 & ~x770;
assign c4209 =  x568 &  x569 & ~x284 & ~x335 & ~x633;
assign c4211 =  x628 &  x629 & ~x18 & ~x138 & ~x363 & ~x462;
assign c4213 =  x181 &  x182 &  x183 & ~x0 & ~x51 & ~x60 & ~x68 & ~x85 & ~x86 & ~x96 & ~x97 & ~x110 & ~x128 & ~x145 & ~x164 & ~x165 & ~x167 & ~x197 & ~x199 & ~x228 & ~x278 & ~x282 & ~x302 & ~x305 & ~x313 & ~x332 & ~x335 & ~x336 & ~x357 & ~x358 & ~x365 & ~x367 & ~x369 & ~x384 & ~x385 & ~x391 & ~x455 & ~x476 & ~x481 & ~x484 & ~x503 & ~x510 & ~x526 & ~x538 & ~x560 & ~x563 & ~x567 & ~x618 & ~x639 & ~x640 & ~x696 & ~x700 & ~x716 & ~x728 & ~x744 & ~x745 & ~x754 & ~x755 & ~x757 & ~x758 & ~x763 & ~x777;
assign c4215 =  x738;
assign c4217 =  x544 &  x545 &  x573 &  x574 & ~x271 & ~x631 & ~x753;
assign c4219 =  x717;
assign c4221 =  x182 &  x183 &  x184 & ~x3 & ~x64 & ~x84 & ~x220 & ~x226 & ~x228 & ~x321 & ~x362 & ~x392 & ~x399 & ~x421 & ~x483 & ~x506 & ~x589 & ~x592 & ~x619 & ~x638 & ~x649 & ~x669 & ~x738 & ~x753 & ~x754 & ~x763 & ~x783;
assign c4223 =  x571 &  x572 &  x573 &  x601 & ~x3 & ~x34 & ~x193 & ~x199 & ~x277 & ~x398 & ~x420 & ~x619 & ~x637 & ~x668 & ~x683 & ~x715;
assign c4225 =  x571 &  x601 & ~x9 & ~x10 & ~x13 & ~x36 & ~x41 & ~x42 & ~x83 & ~x159 & ~x197 & ~x415 & ~x473 & ~x528 & ~x560 & ~x640 & ~x643 & ~x675 & ~x716 & ~x726 & ~x753 & ~x754 & ~x761 & ~x773 & ~x774;
assign c4227 =  x240 &  x241 &  x242 &  x244 &  x266 & ~x157 & ~x160;
assign c4229 =  x656 &  x657 &  x659 & ~x48 & ~x310 & ~x564 & ~x588 & ~x644 & ~x775;
assign c4231 =  x211 &  x236 & ~x3 & ~x24 & ~x31 & ~x61 & ~x66 & ~x74 & ~x82 & ~x100 & ~x143 & ~x152 & ~x153 & ~x154 & ~x179 & ~x199 & ~x201 & ~x283 & ~x307 & ~x358 & ~x383 & ~x391 & ~x399 & ~x439 & ~x454 & ~x483 & ~x500 & ~x512 & ~x522 & ~x537 & ~x539 & ~x614 & ~x619 & ~x638 & ~x674 & ~x692 & ~x752;
assign c4233 =  x543 &  x544 &  x549 & ~x162;
assign c4235 =  x574 & ~x3 & ~x72 & ~x194 & ~x463 & ~x632 & ~x670 & ~x746;
assign c4237 =  x628 & ~x6 & ~x36 & ~x49 & ~x55 & ~x61 & ~x105 & ~x137 & ~x284 & ~x304 & ~x333 & ~x338 & ~x365 & ~x470 & ~x488 & ~x502 & ~x517 & ~x558 & ~x690 & ~x751 & ~x771;
assign c4239 = ~x372 & ~x414 & ~x426 & ~x427 & ~x462 & ~x463 & ~x490 & ~x491 & ~x668 & ~x754 & ~x773;
assign c4241 =  x596 &  x597 &  x598 & ~x422 & ~x730;
assign c4243 =  x156 &  x157 & ~x5 & ~x10 & ~x108 & ~x267 & ~x344 & ~x668 & ~x701;
assign c4245 =  x211 &  x212 &  x236 &  x263 & ~x14 & ~x18 & ~x33 & ~x107 & ~x316 & ~x339 & ~x399 & ~x448;
assign c4247 =  x570 & ~x16 & ~x21 & ~x57 & ~x76 & ~x79 & ~x84 & ~x92 & ~x106 & ~x136 & ~x141 & ~x145 & ~x149 & ~x205 & ~x226 & ~x308 & ~x339 & ~x344 & ~x370 & ~x395 & ~x423 & ~x424 & ~x476 & ~x528 & ~x557 & ~x618 & ~x619 & ~x632 & ~x635 & ~x640 & ~x669 & ~x671 & ~x728 & ~x743 & ~x751 & ~x777;
assign c4249 = ~x252 & ~x320 & ~x368 & ~x372 & ~x373 & ~x374 & ~x394 & ~x400 & ~x402 & ~x453;
assign c4251 =  x211 &  x212 &  x214 & ~x228 & ~x251 & ~x321 & ~x369 & ~x397 & ~x414 & ~x499 & ~x638 & ~x648 & ~x649 & ~x672 & ~x701 & ~x718 & ~x752 & ~x754 & ~x766;
assign c4255 =  x208 &  x209 &  x210 &  x211 & ~x34 & ~x43 & ~x78 & ~x84 & ~x112 & ~x133 & ~x137 & ~x153 & ~x162 & ~x279 & ~x337 & ~x348 & ~x386 & ~x421 & ~x423 & ~x444 & ~x477 & ~x561 & ~x588 & ~x601 & ~x619 & ~x644 & ~x673 & ~x702 & ~x740 & ~x745;
assign c4257 =  x241 &  x242 &  x243 & ~x8 & ~x9 & ~x24 & ~x113 & ~x121 & ~x157 & ~x159 & ~x196 & ~x222 & ~x366 & ~x415 & ~x480 & ~x528 & ~x588 & ~x633 & ~x659 & ~x753;
assign c4259 = ~x36 & ~x313 & ~x319 & ~x342 & ~x344 & ~x345 & ~x347 & ~x372 & ~x373 & ~x374 & ~x376;
assign c4261 =  x244 &  x266 & ~x84 & ~x284 & ~x637 & ~x677 & ~x701 & ~x723;
assign c4263 =  x181 &  x182 &  x183 & ~x9 & ~x25 & ~x30 & ~x69 & ~x144 & ~x192 & ~x199 & ~x225 & ~x251 & ~x292 & ~x310 & ~x332 & ~x333 & ~x335 & ~x339 & ~x363 & ~x384 & ~x413 & ~x503 & ~x561 & ~x586 & ~x615 & ~x620 & ~x647 & ~x675 & ~x701 & ~x706 & ~x763;
assign c4265 =  x207 &  x211 & ~x8 & ~x162 & ~x222 & ~x251 & ~x386 & ~x395 & ~x615 & ~x654 & ~x694 & ~x734 & ~x754;
assign c4267 =  x543 &  x549 & ~x31 & ~x36 & ~x53 & ~x197 & ~x270 & ~x271 & ~x280 & ~x284 & ~x533 & ~x557 & ~x640 & ~x644 & ~x649 & ~x657 & ~x695 & ~x754 & ~x775 & ~x781;
assign c4269 = ~x8 & ~x167 & ~x256 & ~x277 & ~x306 & ~x309 & ~x318 & ~x330 & ~x336 & ~x368 & ~x399 & ~x400 & ~x409 & ~x459 & ~x590 & ~x723 & ~x770;
assign c4271 =  x206 &  x208 &  x232 & ~x69 & ~x76 & ~x87 & ~x100 & ~x137 & ~x144 & ~x164 & ~x226 & ~x421 & ~x682 & ~x725;
assign c4273 =  x234 &  x235 &  x236 &  x238 & ~x134 & ~x137 & ~x161 & ~x201 & ~x228 & ~x246 & ~x278 & ~x415 & ~x676;
assign c4275 = ~x46 & ~x250 & ~x344 & ~x345 & ~x348 & ~x371 & ~x373 & ~x374 & ~x375 & ~x708;
assign c4277 =  x238 &  x239 &  x240 & ~x36 & ~x152 & ~x184 & ~x251 & ~x480 & ~x483 & ~x619 & ~x701 & ~x730;
assign c4279 =  x571 &  x572 &  x573 & ~x1 & ~x16 & ~x53 & ~x61 & ~x84 & ~x113 & ~x120 & ~x138 & ~x145 & ~x166 & ~x171 & ~x196 & ~x201 & ~x225 & ~x251 & ~x283 & ~x451 & ~x611 & ~x616 & ~x633 & ~x653 & ~x657 & ~x659 & ~x696 & ~x720 & ~x734 & ~x745 & ~x769 & ~x775;
assign c4281 =  x210 &  x211 &  x212 &  x236 & ~x47 & ~x57 & ~x116 & ~x267 & ~x293 & ~x305 & ~x307 & ~x386 & ~x421 & ~x446 & ~x468 & ~x564 & ~x581 & ~x694 & ~x721;
assign c4283 =  x266 &  x290 &  x297 & ~x99 & ~x144 & ~x196 & ~x397 & ~x564 & ~x694 & ~x774;
assign c4285 = ~x0 & ~x4 & ~x34 & ~x35 & ~x36 & ~x37 & ~x68 & ~x70 & ~x72 & ~x80 & ~x85 & ~x143 & ~x194 & ~x333 & ~x342 & ~x343 & ~x370 & ~x372 & ~x373 & ~x374 & ~x375 & ~x399 & ~x424 & ~x425 & ~x478 & ~x668 & ~x680 & ~x705 & ~x735 & ~x754 & ~x756;
assign c4287 =  x152 &  x153 &  x179 & ~x192;
assign c4289 =  x206 &  x207 &  x208 & ~x24 & ~x40 & ~x56 & ~x162 & ~x283 & ~x318 & ~x319 & ~x561 & ~x614 & ~x619 & ~x667 & ~x709;
assign c4291 =  x236 &  x632 & ~x18 & ~x98 & ~x280 & ~x335 & ~x439 & ~x446 & ~x524;
assign c4293 =  x571 & ~x3 & ~x43 & ~x115 & ~x311 & ~x335 & ~x339 & ~x353 & ~x560 & ~x682 & ~x761 & ~x770;
assign c4295 =  x265 &  x266 &  x267 &  x269 & ~x6 & ~x27 & ~x42 & ~x43 & ~x52 & ~x69 & ~x100 & ~x102 & ~x155 & ~x171 & ~x172 & ~x175 & ~x195 & ~x201 & ~x212 & ~x222 & ~x253 & ~x282 & ~x363 & ~x367 & ~x424 & ~x476 & ~x524 & ~x559 & ~x584 & ~x589 & ~x610 & ~x642 & ~x700 & ~x725 & ~x727 & ~x750 & ~x754 & ~x761 & ~x783;
assign c4297 =  x293 &  x294 & ~x184 & ~x408 & ~x701;
assign c4299 =  x234 &  x235 &  x236 &  x261 &  x549 & ~x480;
assign c50 =  x275 & ~x153;
assign c52 =  x333;
assign c54 =  x291 & ~x48 & ~x150 & ~x204 & ~x224 & ~x232 & ~x286 & ~x334 & ~x367 & ~x409 & ~x440 & ~x446 & ~x511 & ~x515 & ~x525 & ~x539 & ~x542 & ~x554 & ~x566 & ~x573;
assign c56 =  x239 &  x242 &  x245 &  x266 &  x268 & ~x18 & ~x90 & ~x176 & ~x253 & ~x355 & ~x385 & ~x395 & ~x496 & ~x558 & ~x559 & ~x666 & ~x756;
assign c58 =  x290 &  x318 &  x346 &  x375 &  x406 &  x550 &  x577 & ~x516 & ~x714;
assign c510 =  x247 &  x268 & ~x85 & ~x107 & ~x154 & ~x186 & ~x367 & ~x588 & ~x739 & ~x779;
assign c512 = ~x74 & ~x184 & ~x208 & ~x210 & ~x211 & ~x438 & ~x578 & ~x649;
assign c514 =  x275 & ~x125 & ~x157 & ~x184 & ~x205 & ~x366 & ~x440 & ~x498 & ~x529;
assign c516 =  x188 &  x189 &  x190 &  x213 & ~x247 & ~x333 & ~x394 & ~x416;
assign c518 =  x206 &  x234 &  x290 &  x318 & ~x163 & ~x270 & ~x276 & ~x368 & ~x398 & ~x714;
assign c520 =  x136;
assign c522 =  x182 & ~x237 & ~x238 & ~x239 & ~x240 & ~x243 & ~x463;
assign c524 =  x343 &  x583;
assign c526 =  x154 &  x155 & ~x50 & ~x108 & ~x238 & ~x239 & ~x240 & ~x269 & ~x272 & ~x486 & ~x700;
assign c528 = ~x10 & ~x14 & ~x57 & ~x69 & ~x77 & ~x85 & ~x122 & ~x131 & ~x134 & ~x138 & ~x148 & ~x165 & ~x173 & ~x200 & ~x244 & ~x248 & ~x251 & ~x252 & ~x268 & ~x269 & ~x271 & ~x301 & ~x336 & ~x357 & ~x385 & ~x387 & ~x424 & ~x446 & ~x452 & ~x484 & ~x503 & ~x505 & ~x511 & ~x553 & ~x556 & ~x561 & ~x573 & ~x574 & ~x582 & ~x592 & ~x594 & ~x611 & ~x679 & ~x712 & ~x714 & ~x719 & ~x774 & ~x778;
assign c530 =  x220;
assign c532 =  x278;
assign c534 =  x217 &  x218 &  x239 & ~x330 & ~x357 & ~x703;
assign c536 =  x233 &  x261 &  x289 &  x346 & ~x492;
assign c538 =  x207 & ~x58 & ~x68 & ~x106 & ~x145 & ~x163 & ~x175 & ~x243 & ~x269 & ~x273 & ~x360 & ~x368 & ~x422 & ~x511 & ~x573 & ~x574 & ~x645 & ~x749;
assign c540 =  x155 &  x631 & ~x21 & ~x239 & ~x240 & ~x269 & ~x299 & ~x301 & ~x400 & ~x463;
assign c542 =  x155 &  x178 & ~x60 & ~x89 & ~x164 & ~x237 & ~x239 & ~x241 & ~x244 & ~x272 & ~x519 & ~x560 & ~x591 & ~x700 & ~x743 & ~x765 & ~x772;
assign c544 =  x233 &  x261 &  x346 & ~x297 & ~x546;
assign c546 =  x217 &  x218 &  x240 & ~x7 & ~x46 & ~x129 & ~x198 & ~x333 & ~x423 & ~x453 & ~x612;
assign c548 =  x287 &  x315 &  x373 &  x554 & ~x460;
assign c550 =  x263 &  x291 &  x319 &  x347 &  x375 &  x405 &  x549 &  x550 &  x577 & ~x2 & ~x7 & ~x125 & ~x386 & ~x425 & ~x613;
assign c552 =  x539 & ~x523 & ~x605;
assign c556 =  x233 &  x633 &  x634 & ~x269 & ~x521;
assign c558 =  x217 &  x239 & ~x6 & ~x39 & ~x51 & ~x54 & ~x59 & ~x62 & ~x77 & ~x89 & ~x94 & ~x96 & ~x99 & ~x164 & ~x172 & ~x196 & ~x258 & ~x276 & ~x309 & ~x328 & ~x340 & ~x391 & ~x418 & ~x420 & ~x424 & ~x440 & ~x442 & ~x497 & ~x505 & ~x562 & ~x584 & ~x587 & ~x609 & ~x618 & ~x645 & ~x663 & ~x696 & ~x738 & ~x749 & ~x759 & ~x777 & ~x782;
assign c560 =  x777;
assign c562 =  x247 & ~x183 & ~x186 & ~x656;
assign c564 =  x204 &  x344 & ~x272;
assign c566 =  x210 &  x289 &  x317 &  x345 &  x401 &  x402 & ~x67 & ~x101 & ~x510;
assign c568 =  x335;
assign c570 =  x371;
assign c572 =  x320 & ~x73 & ~x197 & ~x355 & ~x411 & ~x458 & ~x468 & ~x486 & ~x551 & ~x578 & ~x606 & ~x662 & ~x757;
assign c574 = ~x9 & ~x38 & ~x92 & ~x142 & ~x208 & ~x209 & ~x210 & ~x211 & ~x288 & ~x412 & ~x448 & ~x473 & ~x479 & ~x522 & ~x662 & ~x719 & ~x724 & ~x759 & ~x765;
assign c576 =  x236 &  x264 &  x265 &  x352 &  x598 & ~x457 & ~x489;
assign c578 =  x209 &  x210 &  x211 &  x213 &  x236 &  x237 & ~x194 & ~x270 & ~x273 & ~x515 & ~x773;
assign c580 = ~x54 & ~x134 & ~x156 & ~x162 & ~x169 & ~x178 & ~x181 & ~x182 & ~x183 & ~x211 & ~x258 & ~x287 & ~x411 & ~x438 & ~x440 & ~x468 & ~x496 & ~x524 & ~x525 & ~x582 & ~x606 & ~x663 & ~x768;
assign c582 =  x137;
assign c584 =  x161 & ~x142 & ~x244 & ~x272 & ~x483;
assign c586 =  x209 &  x263 &  x291 &  x377 &  x522 &  x577 & ~x256;
assign c588 =  x511 & ~x98 & ~x181 & ~x385 & ~x656;
assign c590 =  x162 & ~x244;
assign c592 =  x232 &  x260 &  x663;
assign c594 =  x212 &  x686 & ~x352 & ~x382;
assign c596 =  x260 &  x373 & ~x20 & ~x165 & ~x167 & ~x244 & ~x420 & ~x517 & ~x546 & ~x592 & ~x678 & ~x758;
assign c598 =  x305;
assign c5100 =  x316 &  x660 & ~x576;
assign c5102 =  x242 &  x245 & ~x42 & ~x54 & ~x65 & ~x68 & ~x74 & ~x125 & ~x159 & ~x307 & ~x309 & ~x342 & ~x356 & ~x390 & ~x394 & ~x440 & ~x449 & ~x505 & ~x532 & ~x585 & ~x636 & ~x641 & ~x679 & ~x729 & ~x751;
assign c5104 =  x305;
assign c5106 =  x628 & ~x30 & ~x34 & ~x72 & ~x98 & ~x111 & ~x120 & ~x143 & ~x171 & ~x173 & ~x216 & ~x239 & ~x240 & ~x242 & ~x244 & ~x251 & ~x269 & ~x270 & ~x271 & ~x273 & ~x301 & ~x329 & ~x335 & ~x359 & ~x361 & ~x367 & ~x398 & ~x417 & ~x425 & ~x450 & ~x457 & ~x463 & ~x472 & ~x486 & ~x584 & ~x667 & ~x685 & ~x689 & ~x693 & ~x725 & ~x744 & ~x747;
assign c5108 =  x276;
assign c5110 =  x304 & ~x184;
assign c5112 =  x208 &  x235 &  x263 &  x291 &  x320 & ~x275 & ~x460 & ~x486 & ~x661;
assign c5114 =  x465 & ~x89 & ~x365 & ~x439 & ~x496 & ~x523 & ~x551 & ~x606 & ~x632 & ~x659;
assign c5116 = ~x129 & ~x156 & ~x180 & ~x181 & ~x409 & ~x438 & ~x468 & ~x522 & ~x551 & ~x578 & ~x605 & ~x606;
assign c5118 =  x287 &  x372 & ~x521;
assign c5120 =  x155 &  x628 &  x629 & ~x26 & ~x28 & ~x40 & ~x82 & ~x120 & ~x162 & ~x191 & ~x217 & ~x239 & ~x240 & ~x244 & ~x271 & ~x458 & ~x501 & ~x516 & ~x674 & ~x700 & ~x702 & ~x710 & ~x731 & ~x744;
assign c5122 =  x305;
assign c5124 =  x40;
assign c5126 =  x237 &  x319 &  x347 &  x375 &  x376 &  x493 & ~x544;
assign c5128 =  x317 &  x633 &  x685 & ~x256 & ~x484 & ~x543;
assign c5130 =  x237 &  x291 &  x347 &  x375 & ~x56 & ~x68 & ~x191 & ~x389 & ~x398 & ~x427 & ~x458 & ~x497;
assign c5132 =  x275;
assign c5134 =  x211 &  x214 &  x236 &  x239 &  x660 & ~x155;
assign c5136 =  x403 & ~x159 & ~x182 & ~x208 & ~x210 & ~x551;
assign c5138 =  x207 &  x235 &  x263 &  x291 &  x319 &  x347 &  x522 & ~x66 & ~x135 & ~x400;
assign c5140 =  x8;
assign c5142 =  x206 &  x262 &  x290 &  x318 &  x578 & ~x455;
assign c5144 =  x155 & ~x54 & ~x217 & ~x239 & ~x240 & ~x247 & ~x269 & ~x288 & ~x329 & ~x391 & ~x424 & ~x446 & ~x458 & ~x487 & ~x501 & ~x615 & ~x662 & ~x670 & ~x697 & ~x700 & ~x718 & ~x746 & ~x749 & ~x765 & ~x774;
assign c5146 =  x188 &  x238 &  x239 & ~x80 & ~x193 & ~x244;
assign c5148 =  x167;
assign c5150 =  x707;
assign c5152 =  x320 &  x627 & ~x239 & ~x240 & ~x269 & ~x462;
assign c5154 =  x304 & ~x525;
assign c5156 =  x323 & ~x157 & ~x183 & ~x208 & ~x211 & ~x467 & ~x578;
assign c5158 =  x235 &  x290 &  x318 &  x579 &  x632 & ~x173 & ~x343 & ~x514 & ~x520;
assign c5160 =  x264 &  x292 &  x375 &  x376 &  x404 &  x405 &  x521 &  x548 & ~x12 & ~x99 & ~x167 & ~x253 & ~x760;
assign c5162 =  x209 &  x210 &  x213 &  x214 &  x237 &  x632 &  x659 & ~x134 & ~x279 & ~x330 & ~x331 & ~x625;
assign c5164 = ~x211 & ~x606 & ~x632;
assign c5166 =  x192;
assign c5168 =  x206 &  x234 &  x262 &  x524 & ~x269 & ~x301 & ~x398;
assign c5170 =  x181 &  x182 &  x209 &  x347 & ~x56 & ~x269 & ~x486;
assign c5172 =  x188 &  x210 &  x211 &  x238 &  x239 & ~x3 & ~x52 & ~x203 & ~x328 & ~x334 & ~x443 & ~x650;
assign c5174 =  x189 &  x213 &  x239 & ~x17 & ~x61 & ~x300 & ~x364 & ~x498 & ~x593 & ~x719;
assign c5176 = ~x69 & ~x124 & ~x156 & ~x172 & ~x180 & ~x255 & ~x261 & ~x379 & ~x409 & ~x410 & ~x438 & ~x522 & ~x551 & ~x578 & ~x605 & ~x606 & ~x633 & ~x661 & ~x667 & ~x753;
assign c5178 =  x403 & ~x240 & ~x630;
assign c5180 =  x511 & ~x186;
assign c5182 =  x217 &  x242 & ~x300 & ~x327 & ~x356 & ~x387;
assign c5184 =  x209 &  x210 &  x213 &  x214 &  x237 &  x238 &  x239 & ~x0 & ~x5 & ~x22 & ~x23 & ~x31 & ~x57 & ~x68 & ~x77 & ~x87 & ~x102 & ~x148 & ~x149 & ~x162 & ~x226 & ~x229 & ~x252 & ~x258 & ~x278 & ~x296 & ~x298 & ~x308 & ~x312 & ~x329 & ~x331 & ~x335 & ~x422 & ~x424 & ~x426 & ~x473 & ~x500 & ~x526 & ~x646 & ~x675 & ~x699 & ~x702 & ~x703 & ~x729 & ~x750 & ~x767;
assign c5186 =  x263 &  x291 &  x466 &  x494 &  x522 &  x550 &  x577;
assign c5188 =  x259 &  x314 &  x555;
assign c5190 =  x301 & ~x183 & ~x213 & ~x411;
assign c5192 =  x157 & ~x25 & ~x164 & ~x239 & ~x240 & ~x245 & ~x269 & ~x369 & ~x486 & ~x505 & ~x710 & ~x738;
assign c5194 =  x375 & ~x97 & ~x378 & ~x380 & ~x409 & ~x411 & ~x438 & ~x551 & ~x610;
assign c5196 =  x403 & ~x181 & ~x554 & ~x575 & ~x602;
assign c5198 =  x206 &  x234 & ~x269 & ~x329 & ~x492 & ~x520 & ~x547;
assign c5200 =  x422;
assign c5202 =  x192;
assign c5204 = ~x18 & ~x53 & ~x73 & ~x75 & ~x82 & ~x99 & ~x112 & ~x139 & ~x173 & ~x215 & ~x237 & ~x238 & ~x239 & ~x240 & ~x244 & ~x267 & ~x269 & ~x271 & ~x298 & ~x308 & ~x334 & ~x335 & ~x365 & ~x397 & ~x443 & ~x623 & ~x714 & ~x745 & ~x765;
assign c5206 = ~x11 & ~x42 & ~x43 & ~x80 & ~x170 & ~x237 & ~x238 & ~x239 & ~x240 & ~x269 & ~x276 & ~x310 & ~x311 & ~x334 & ~x370 & ~x486 & ~x520 & ~x651 & ~x666 & ~x677 & ~x679 & ~x694 & ~x760;
assign c5208 =  x556;
assign c5210 =  x188 &  x211 & ~x244 & ~x269 & ~x270;
assign c5212 = ~x238 & ~x239 & ~x240 & ~x269 & ~x400 & ~x432 & ~x434;
assign c5214 =  x238 &  x265 &  x294 &  x547 & ~x152 & ~x261 & ~x487 & ~x606 & ~x618 & ~x712 & ~x714;
assign c5216 =  x265 &  x293 &  x376 &  x548 & ~x203 & ~x205 & ~x312 & ~x486 & ~x551 & ~x606 & ~x611;
assign c5218 = ~x10 & ~x49 & ~x153 & ~x407 & ~x409 & ~x410 & ~x419 & ~x437 & ~x521 & ~x522 & ~x551 & ~x578 & ~x783;
assign c5220 =  x176 &  x608;
assign c5222 =  x249;
assign c5224 =  x277;
assign c5226 =  x217 &  x219 & ~x327;
assign c5228 =  x248 & ~x355;
assign c5230 =  x249;
assign c5232 =  x293 &  x538 & ~x41 & ~x146 & ~x198 & ~x329 & ~x372 & ~x400 & ~x444 & ~x506 & ~x677 & ~x686 & ~x727 & ~x781;
assign c5234 =  x301 &  x304;
assign c5236 =  x264 &  x292 &  x493 &  x628 & ~x145 & ~x382 & ~x421 & ~x440 & ~x515 & ~x586 & ~x729;
assign c5238 =  x158 &  x159 &  x160 & ~x429;
assign c5240 =  x136;
assign c5242 =  x292 &  x403 &  x577 & ~x46 & ~x260 & ~x287 & ~x777;
assign c5244 =  x133 &  x156;
assign c5246 =  x213 &  x236 &  x237 &  x238 & ~x11 & ~x114 & ~x513 & ~x516 & ~x517 & ~x547 & ~x650 & ~x764 & ~x771;
assign c5248 = ~x186;
assign c5250 =  x210 &  x238 &  x293 &  x547 &  x598 & ~x429;
assign c5252 =  x209 &  x210 &  x237 &  x264 &  x293 &  x548 &  x627 &  x628 & ~x283 & ~x345;
assign c5254 =  x206 &  x207 &  x235 &  x290 &  x318 &  x495;
assign c5256 =  x191 & ~x248;
assign c5258 =  x184 &  x207 &  x208 &  x209 &  x210 &  x375 & ~x269 & ~x298;
assign c5260 =  x550 &  x577 & ~x243 & ~x266 & ~x343 & ~x446 & ~x514 & ~x587;
assign c5262 =  x158 &  x159 & ~x242 & ~x246 & ~x272 & ~x486;
assign c5264 =  x713;
assign c5266 =  x263 &  x264 & ~x96 & ~x125 & ~x141 & ~x172 & ~x205 & ~x380 & ~x385 & ~x409 & ~x438 & ~x505;
assign c5268 =  x131 &  x158 &  x210 & ~x245;
assign c5270 =  x375 & ~x382 & ~x410 & ~x576 & ~x602 & ~x630;
assign c5272 =  x232 &  x316 &  x372 & ~x329 & ~x547;
assign c5274 =  x304;
assign c5276 =  x245 &  x247 &  x268 & ~x677;
assign c5278 =  x182 &  x208 & ~x238 & ~x239 & ~x243 & ~x269 & ~x299 & ~x515 & ~x516 & ~x557;
assign c5280 =  x190 &  x214 & ~x298;
assign c5282 =  x159 &  x160 &  x210 & ~x23 & ~x269;
assign c5284 =  x155 & ~x85 & ~x101 & ~x218 & ~x239 & ~x240 & ~x269 & ~x298 & ~x300 & ~x471 & ~x490 & ~x512 & ~x556 & ~x704 & ~x771;
assign c5286 =  x289 &  x346 &  x633 & ~x520;
assign c5288 =  x206 &  x208 &  x262 &  x290 &  x318 &  x319 & ~x99 & ~x272;
assign c5290 =  x511 & ~x156 & ~x183 & ~x603;
assign c5292 =  x235 &  x290 &  x318 &  x375 &  x495;
assign c5294 = ~x98 & ~x181 & ~x184 & ~x208 & ~x209 & ~x210 & ~x211 & ~x261 & ~x411 & ~x551 & ~x553 & ~x578;
assign c5296 =  x192;
assign c5298 =  x162 & ~x244;
assign c51 =  x330 &  x358;
assign c53 =  x329 &  x412 &  x440;
assign c55 =  x426 &  x454 & ~x353;
assign c57 =  x325 &  x406 &  x433 &  x434;
assign c59 =  x243 &  x298 &  x325 & ~x24 & ~x30 & ~x83 & ~x139 & ~x175 & ~x219 & ~x226 & ~x230 & ~x259 & ~x340 & ~x357 & ~x389 & ~x417 & ~x559 & ~x562 & ~x741 & ~x765 & ~x776 & ~x781;
assign c511 =  x328 &  x355 & ~x9 & ~x21 & ~x30 & ~x33 & ~x38 & ~x57 & ~x63 & ~x87 & ~x106 & ~x137 & ~x174 & ~x203 & ~x283 & ~x306 & ~x307 & ~x323 & ~x333 & ~x362 & ~x391 & ~x449 & ~x451 & ~x535 & ~x559 & ~x664 & ~x675 & ~x742 & ~x754 & ~x772;
assign c513 =  x325 &  x435;
assign c515 =  x323 &  x351 &  x406 & ~x62 & ~x219 & ~x226 & ~x280 & ~x356 & ~x421 & ~x424 & ~x497 & ~x511 & ~x592 & ~x594 & ~x710 & ~x758 & ~x759;
assign c517 =  x328 &  x355 & ~x12 & ~x16 & ~x22 & ~x35 & ~x65 & ~x67 & ~x79 & ~x106 & ~x107 & ~x139 & ~x166 & ~x173 & ~x194 & ~x203 & ~x226 & ~x256 & ~x305 & ~x359 & ~x368 & ~x395 & ~x441 & ~x445 & ~x447 & ~x449 & ~x469 & ~x478 & ~x535 & ~x563 & ~x590 & ~x614 & ~x615 & ~x675 & ~x704 & ~x726 & ~x735 & ~x742 & ~x760;
assign c519 =  x329 & ~x739;
assign c521 =  x297 &  x325 &  x380 & ~x571;
assign c523 =  x430 &  x458 &  x485 &  x486 &  x513 &  x541 & ~x254 & ~x506 & ~x536 & ~x676 & ~x731 & ~x769 & ~x778;
assign c525 =  x243 &  x325 & ~x374;
assign c527 =  x455 &  x625 & ~x391;
assign c529 =  x380 &  x408 &  x435 & ~x128 & ~x194 & ~x572 & ~x752;
assign c531 =  x152 &  x267 & ~x678;
assign c533 = ~x11 & ~x122 & ~x128 & ~x185 & ~x317 & ~x346 & ~x448 & ~x599 & ~x627 & ~x654;
assign c535 = ~x292 & ~x319 & ~x320 & ~x347 & ~x348 & ~x375 & ~x376 & ~x403 & ~x431 & ~x706;
assign c537 =  x324 & ~x15 & ~x28 & ~x128 & ~x226 & ~x249 & ~x332 & ~x511 & ~x561 & ~x621 & ~x627;
assign c539 =  x357 &  x384;
assign c541 =  x434 &  x461 &  x488 &  x516 & ~x61 & ~x590 & ~x669 & ~x739;
assign c543 =  x328 & ~x320;
assign c545 =  x430 &  x457 &  x458 &  x485 &  x513 &  x541 & ~x28 & ~x81 & ~x488 & ~x645 & ~x745 & ~x767;
assign c547 =  x464 & ~x377 & ~x405 & ~x756;
assign c549 =  x413 & ~x352;
assign c551 =  x325 & ~x4 & ~x38 & ~x40 & ~x50 & ~x81 & ~x88 & ~x137 & ~x139 & ~x148 & ~x164 & ~x166 & ~x171 & ~x191 & ~x293 & ~x341 & ~x365 & ~x421 & ~x425 & ~x445 & ~x448 & ~x450 & ~x563 & ~x586 & ~x638 & ~x664 & ~x665 & ~x699 & ~x746 & ~x758 & ~x759 & ~x761 & ~x780;
assign c553 =  x435 &  x491 & ~x321;
assign c555 =  x433 &  x488 &  x515 & ~x16 & ~x31 & ~x254 & ~x275 & ~x301 & ~x467 & ~x473 & ~x556 & ~x564 & ~x586 & ~x727 & ~x777;
assign c557 =  x274 &  x626;
assign c559 =  x325 &  x379 &  x407 & ~x3 & ~x16 & ~x31 & ~x37 & ~x46 & ~x67 & ~x77 & ~x82 & ~x112 & ~x117 & ~x137 & ~x150 & ~x163 & ~x248 & ~x276 & ~x277 & ~x472 & ~x543 & ~x699 & ~x704 & ~x769;
assign c561 =  x458 &  x486 &  x514 & ~x0 & ~x1 & ~x9 & ~x64 & ~x79 & ~x87 & ~x88 & ~x106 & ~x110 & ~x113 & ~x114 & ~x173 & ~x194 & ~x305 & ~x341 & ~x424 & ~x426 & ~x448 & ~x455 & ~x476 & ~x566 & ~x585 & ~x589 & ~x592 & ~x622 & ~x652 & ~x669 & ~x673 & ~x678 & ~x684 & ~x692 & ~x711 & ~x723 & ~x737 & ~x743 & ~x772 & ~x778;
assign c563 =  x331;
assign c565 =  x354 &  x381 &  x409 & ~x85 & ~x91 & ~x105 & ~x323 & ~x421 & ~x589 & ~x614 & ~x766;
assign c567 =  x484 &  x596 &  x625 & ~x50 & ~x117 & ~x202 & ~x336 & ~x448 & ~x732 & ~x780;
assign c569 =  x464 & ~x377 & ~x626;
assign c573 =  x436 & ~x132 & ~x156 & ~x715;
assign c575 =  x379 &  x406 &  x434 &  x461 & ~x15 & ~x25 & ~x30 & ~x35 & ~x76 & ~x80 & ~x146 & ~x309 & ~x360 & ~x391 & ~x420 & ~x421 & ~x447 & ~x482 & ~x511 & ~x539 & ~x560 & ~x564 & ~x567 & ~x587 & ~x648 & ~x672 & ~x681 & ~x698 & ~x716 & ~x726 & ~x730 & ~x732 & ~x733 & ~x760 & ~x767;
assign c577 =  x459 &  x486 &  x487 &  x514 & ~x6 & ~x23 & ~x40 & ~x88 & ~x90 & ~x107 & ~x246 & ~x257 & ~x275 & ~x334 & ~x336 & ~x339 & ~x361 & ~x369 & ~x371 & ~x386 & ~x412 & ~x527 & ~x536 & ~x558 & ~x640 & ~x645 & ~x646 & ~x694 & ~x711 & ~x735 & ~x749 & ~x767;
assign c579 =  x325 &  x405 &  x406 & ~x54 & ~x60 & ~x79 & ~x137 & ~x166 & ~x167 & ~x199 & ~x276 & ~x277 & ~x302 & ~x357 & ~x365 & ~x366 & ~x397 & ~x418 & ~x482 & ~x508 & ~x530 & ~x538 & ~x592 & ~x642 & ~x672 & ~x731 & ~x742 & ~x745 & ~x760 & ~x771;
assign c581 =  x354 & ~x223 & ~x322 & ~x350 & ~x413 & ~x476 & ~x619;
assign c583 = ~x42 & ~x69 & ~x89 & ~x141 & ~x242 & ~x269 & ~x285 & ~x357 & ~x366 & ~x399 & ~x420 & ~x470 & ~x507 & ~x538 & ~x592 & ~x598 & ~x624 & ~x627 & ~x647 & ~x653 & ~x654 & ~x657 & ~x687;
assign c585 =  x385 & ~x661 & ~x781;
assign c587 =  x455 &  x483 &  x597 & ~x408;
assign c589 =  x435 &  x489 &  x517 & ~x1 & ~x12 & ~x24 & ~x26 & ~x96 & ~x115 & ~x116 & ~x229 & ~x368 & ~x450 & ~x477 & ~x583 & ~x620 & ~x699 & ~x704 & ~x780 & ~x781;
assign c591 =  x456 &  x457 &  x484 &  x540 & ~x664;
assign c593 =  x330 &  x626;
assign c595 =  x458 &  x572 & ~x19 & ~x115 & ~x202 & ~x244 & ~x254 & ~x389 & ~x563 & ~x567 & ~x624 & ~x654 & ~x718;
assign c597 = ~x103 & ~x319 & ~x320 & ~x347 & ~x348 & ~x376 & ~x403 & ~x435;
assign c599 =  x409 &  x463 &  x464 & ~x352;
assign c5101 =  x357 & ~x499;
assign c5103 =  x435 &  x463 &  x518 & ~x445 & ~x509 & ~x541 & ~x542;
assign c5105 =  x458 &  x486 &  x514 &  x542 &  x599 & ~x38 & ~x42 & ~x53 & ~x77 & ~x115 & ~x192 & ~x202 & ~x233 & ~x302 & ~x308 & ~x453 & ~x478 & ~x528 & ~x564 & ~x624 & ~x690 & ~x741 & ~x755 & ~x771;
assign c5107 =  x354 &  x436 &  x463;
assign c5109 =  x269 & ~x57 & ~x60 & ~x85 & ~x108 & ~x218 & ~x292 & ~x302 & ~x356 & ~x398 & ~x415 & ~x425 & ~x505 & ~x518 & ~x545 & ~x615 & ~x704 & ~x740 & ~x759 & ~x769;
assign c5111 =  x382 & ~x132 & ~x158 & ~x159 & ~x323 & ~x349 & ~x377 & ~x422 & ~x567 & ~x594;
assign c5113 =  x430 &  x458 &  x485 &  x486 &  x513 &  x541 & ~x1 & ~x16 & ~x18 & ~x21 & ~x30 & ~x40 & ~x42 & ~x52 & ~x64 & ~x65 & ~x80 & ~x83 & ~x87 & ~x121 & ~x137 & ~x173 & ~x176 & ~x192 & ~x197 & ~x221 & ~x223 & ~x278 & ~x286 & ~x334 & ~x338 & ~x339 & ~x363 & ~x369 & ~x370 & ~x414 & ~x421 & ~x444 & ~x448 & ~x531 & ~x592 & ~x612 & ~x615 & ~x621 & ~x672 & ~x678 & ~x691 & ~x722 & ~x738 & ~x758 & ~x763 & ~x768 & ~x778;
assign c5115 = ~x320 & ~x347 & ~x348 & ~x375 & ~x376 & ~x403 & ~x404 & ~x430;
assign c5117 =  x459 &  x486 &  x514 &  x571 & ~x474;
assign c5119 =  x324 &  x406 & ~x24 & ~x69 & ~x275 & ~x292 & ~x395 & ~x414 & ~x752 & ~x780;
assign c5121 =  x121;
assign c5123 =  x386 & ~x326 & ~x353;
assign c5125 =  x269;
assign c5127 =  x325 &  x379 &  x405 & ~x150 & ~x221 & ~x382 & ~x707;
assign c5129 =  x406 &  x433 &  x434 &  x460 & ~x52 & ~x58 & ~x60 & ~x65 & ~x114 & ~x115 & ~x150 & ~x167 & ~x206 & ~x226 & ~x314 & ~x372 & ~x386 & ~x448 & ~x478 & ~x561 & ~x612 & ~x613 & ~x649 & ~x709 & ~x737 & ~x767 & ~x781;
assign c5131 =  x456 &  x484;
assign c5133 =  x459 &  x460 &  x487 &  x515 &  x543 & ~x46 & ~x60 & ~x106 & ~x117 & ~x448 & ~x619 & ~x718 & ~x731;
assign c5135 =  x328 & ~x17 & ~x109 & ~x120 & ~x253 & ~x323 & ~x472 & ~x504 & ~x505 & ~x586 & ~x620 & ~x707 & ~x740 & ~x780;
assign c5137 =  x296 &  x323 &  x604 &  x624 & ~x519;
assign c5139 =  x379 & ~x20 & ~x31 & ~x37 & ~x43 & ~x73 & ~x110 & ~x119 & ~x158 & ~x173 & ~x186 & ~x214 & ~x277 & ~x333 & ~x359 & ~x386 & ~x392 & ~x415 & ~x417 & ~x418 & ~x452 & ~x477 & ~x479 & ~x514 & ~x528 & ~x539 & ~x571 & ~x599 & ~x618 & ~x624 & ~x654 & ~x694 & ~x698 & ~x699 & ~x766 & ~x777;
assign c5141 =  x460 &  x488 & ~x91 & ~x164 & ~x169 & ~x249 & ~x289 & ~x318;
assign c5143 =  x491 &  x546 & ~x448 & ~x652 & ~x655;
assign c5145 =  x295 &  x322 &  x655 & ~x7 & ~x63 & ~x265 & ~x780;
assign c5147 =  x151 &  x152 & ~x83 & ~x91 & ~x109 & ~x114 & ~x140 & ~x168 & ~x235 & ~x262 & ~x343 & ~x415 & ~x424 & ~x441 & ~x445 & ~x500 & ~x589 & ~x703;
assign c5149 =  x354 &  x408 & ~x413;
assign c5151 =  x460 &  x488 &  x515 &  x543 & ~x11 & ~x14 & ~x32 & ~x48 & ~x147 & ~x164 & ~x195 & ~x391 & ~x402 & ~x477 & ~x509 & ~x512 & ~x587 & ~x594 & ~x609 & ~x678 & ~x741;
assign c5153 =  x271 &  x325 &  x379 & ~x117 & ~x252 & ~x527 & ~x555 & ~x590 & ~x744 & ~x759 & ~x781;
assign c5155 =  x517 &  x545 &  x573 & ~x16 & ~x276 & ~x303 & ~x414 & ~x418 & ~x423 & ~x625 & ~x652 & ~x668 & ~x781;
assign c5157 =  x228;
assign c5159 =  x329 & ~x117 & ~x223 & ~x323 & ~x562 & ~x693;
assign c5161 =  x152 &  x295 & ~x236 & ~x290 & ~x317 & ~x739;
assign c5163 =  x457 &  x496 & ~x55 & ~x476;
assign c5165 = ~x206 & ~x374 & ~x375 & ~x403 & ~x586 & ~x598;
assign c5167 =  x324 & ~x20 & ~x30 & ~x55 & ~x102 & ~x104 & ~x265 & ~x273 & ~x277 & ~x281 & ~x343 & ~x370 & ~x371 & ~x485 & ~x565 & ~x692 & ~x704 & ~x757;
assign c5169 =  x380 &  x461 &  x462;
assign c5171 =  x400 &  x455 & ~x12 & ~x16 & ~x20 & ~x28 & ~x37 & ~x38 & ~x46 & ~x50 & ~x116 & ~x250 & ~x378 & ~x406 & ~x451 & ~x531 & ~x585 & ~x587 & ~x644 & ~x713 & ~x752 & ~x758 & ~x765;
assign c5173 =  x328 &  x356 &  x383 & ~x16 & ~x21 & ~x22 & ~x42 & ~x64 & ~x72 & ~x81 & ~x87 & ~x107 & ~x108 & ~x115 & ~x121 & ~x142 & ~x145 & ~x147 & ~x148 & ~x170 & ~x280 & ~x335 & ~x360 & ~x415 & ~x420 & ~x422 & ~x450 & ~x476 & ~x501 & ~x530 & ~x561 & ~x583 & ~x585 & ~x638 & ~x640 & ~x642 & ~x643 & ~x644 & ~x646 & ~x671 & ~x706 & ~x724 & ~x737 & ~x739 & ~x743 & ~x770 & ~x772;
assign c5175 =  x327 &  x355 &  x382 & ~x0 & ~x7 & ~x12 & ~x20 & ~x38 & ~x60 & ~x81 & ~x117 & ~x194 & ~x201 & ~x277 & ~x331 & ~x341 & ~x360 & ~x560 & ~x765 & ~x769;
assign c5177 =  x382 &  x437 & ~x1 & ~x2 & ~x7 & ~x35 & ~x77 & ~x127 & ~x128 & ~x133 & ~x139 & ~x193 & ~x249 & ~x252 & ~x338 & ~x421 & ~x472 & ~x479 & ~x527 & ~x555 & ~x568 & ~x589 & ~x599 & ~x610 & ~x626 & ~x653 & ~x753 & ~x780;
assign c5179 =  x328 & ~x24 & ~x62 & ~x118 & ~x172 & ~x322 & ~x323 & ~x360 & ~x448 & ~x476 & ~x564 & ~x666 & ~x673 & ~x740 & ~x749 & ~x765;
assign c5181 = ~x241 & ~x296 & ~x318 & ~x447 & ~x482 & ~x510 & ~x627 & ~x628;
assign c5183 =  x380 &  x407 & ~x1 & ~x68 & ~x94 & ~x98 & ~x151 & ~x276 & ~x295 & ~x371 & ~x413 & ~x427 & ~x452 & ~x500 & ~x504 & ~x510 & ~x551 & ~x571 & ~x639 & ~x703 & ~x718 & ~x722 & ~x728 & ~x752;
assign c5185 =  x411 & ~x64 & ~x90 & ~x91 & ~x107 & ~x115 & ~x154 & ~x191 & ~x197 & ~x248 & ~x277 & ~x281 & ~x331 & ~x335 & ~x366 & ~x448 & ~x471 & ~x481 & ~x500 & ~x508 & ~x558 & ~x566 & ~x585 & ~x587 & ~x594 & ~x612 & ~x624 & ~x627 & ~x669 & ~x671 & ~x682 & ~x720 & ~x722 & ~x742 & ~x753 & ~x777 & ~x780;
assign c5187 =  x455 &  x567 & ~x379;
assign c5189 =  x327 &  x354 &  x409 & ~x20 & ~x43 & ~x63 & ~x104 & ~x111 & ~x414 & ~x421 & ~x501 & ~x672 & ~x732 & ~x758;
assign c5191 =  x269 &  x325 &  x381 & ~x4 & ~x36 & ~x91 & ~x119 & ~x144 & ~x195 & ~x572 & ~x599 & ~x722;
assign c5193 =  x152 &  x295 &  x322 & ~x1 & ~x40 & ~x104 & ~x290 & ~x356 & ~x386 & ~x715 & ~x764;
assign c5195 =  x462 & ~x14 & ~x111 & ~x169 & ~x222 & ~x230 & ~x272 & ~x393 & ~x509 & ~x537 & ~x540 & ~x657 & ~x658 & ~x738 & ~x741 & ~x775;
assign c5197 =  x437 & ~x377 & ~x406 & ~x570 & ~x627;
assign c5199 =  x455 &  x483 & ~x32 & ~x35 & ~x338 & ~x377;
assign c5201 =  x459 &  x486 &  x514 &  x541;
assign c5203 =  x243 &  x299 &  x326 & ~x20 & ~x62 & ~x104 & ~x194 & ~x418 & ~x688 & ~x709;
assign c5205 =  x603 & ~x4 & ~x21 & ~x27 & ~x64 & ~x77 & ~x79 & ~x82 & ~x83 & ~x104 & ~x106 & ~x120 & ~x143 & ~x149 & ~x163 & ~x171 & ~x172 & ~x174 & ~x197 & ~x198 & ~x199 & ~x215 & ~x216 & ~x221 & ~x224 & ~x225 & ~x249 & ~x275 & ~x299 & ~x357 & ~x385 & ~x424 & ~x446 & ~x504 & ~x508 & ~x511 & ~x527 & ~x538 & ~x568 & ~x584 & ~x624 & ~x625 & ~x637 & ~x644 & ~x657 & ~x691 & ~x699 & ~x705 & ~x709 & ~x714 & ~x717 & ~x736 & ~x766 & ~x778 & ~x781;
assign c5207 =  x742;
assign c5209 =  x327 &  x355 & ~x23 & ~x26 & ~x40 & ~x83 & ~x91 & ~x103 & ~x111 & ~x114 & ~x121 & ~x137 & ~x173 & ~x249 & ~x283 & ~x322 & ~x473 & ~x499 & ~x532 & ~x560 & ~x564 & ~x586 & ~x673 & ~x675 & ~x694 & ~x704 & ~x719 & ~x720 & ~x767;
assign c5211 =  x325 &  x407 &  x434 &  x435;
assign c5213 =  x295 &  x322 &  x379 &  x656 & ~x30 & ~x221 & ~x279 & ~x280 & ~x311 & ~x333 & ~x341 & ~x452 & ~x731 & ~x763;
assign c5215 =  x485 &  x512 &  x540 &  x596 & ~x27 & ~x55 & ~x120 & ~x166 & ~x307 & ~x559 & ~x619 & ~x744;
assign c5217 =  x412 & ~x175 & ~x205 & ~x406;
assign c5219 = ~x165 & ~x264 & ~x290 & ~x292 & ~x318 & ~x319 & ~x346 & ~x400 & ~x482 & ~x555;
assign c5221 =  x518 &  x546 & ~x110 & ~x455 & ~x540 & ~x592 & ~x597 & ~x654 & ~x707 & ~x713 & ~x765;
assign c5223 =  x229;
assign c5225 =  x460 &  x488 &  x516 &  x544 & ~x54 & ~x119 & ~x280 & ~x302 & ~x566 & ~x622 & ~x710;
assign c5227 =  x354 &  x409 & ~x0 & ~x7 & ~x33 & ~x37 & ~x105 & ~x122 & ~x132 & ~x230 & ~x393 & ~x441 & ~x649 & ~x663 & ~x779;
assign c5229 =  x297 &  x407 & ~x20 & ~x101 & ~x391 & ~x540 & ~x555 & ~x563 & ~x586 & ~x645 & ~x777;
assign c5231 =  x439 &  x440 & ~x79 & ~x110 & ~x115 & ~x138 & ~x235 & ~x389 & ~x451 & ~x501 & ~x666 & ~x688 & ~x743;
assign c5233 =  x323 & ~x8 & ~x20 & ~x28 & ~x33 & ~x44 & ~x58 & ~x68 & ~x82 & ~x99 & ~x110 & ~x112 & ~x121 & ~x134 & ~x172 & ~x199 & ~x225 & ~x228 & ~x245 & ~x250 & ~x253 & ~x271 & ~x274 & ~x309 & ~x312 & ~x314 & ~x326 & ~x359 & ~x365 & ~x368 & ~x390 & ~x420 & ~x448 & ~x456 & ~x475 & ~x477 & ~x481 & ~x510 & ~x533 & ~x557 & ~x562 & ~x567 & ~x587 & ~x592 & ~x594 & ~x614 & ~x621 & ~x641 & ~x652 & ~x670 & ~x671 & ~x677 & ~x695 & ~x704 & ~x707 & ~x720 & ~x731 & ~x755 & ~x762 & ~x783;
assign c5235 =  x359;
assign c5237 =  x426 &  x454;
assign c5239 =  x457 &  x485 &  x572 &  x600 &  x601 & ~x93 & ~x164 & ~x191 & ~x337 & ~x424 & ~x448 & ~x586 & ~x670 & ~x687 & ~x690 & ~x700 & ~x712 & ~x716 & ~x737 & ~x746 & ~x749;
assign c5241 =  x322 &  x406 & ~x13 & ~x75 & ~x85 & ~x95 & ~x111 & ~x128 & ~x129 & ~x133 & ~x169 & ~x225 & ~x248 & ~x249 & ~x276 & ~x279 & ~x448 & ~x529 & ~x539 & ~x675 & ~x682 & ~x772;
assign c5243 =  x326 &  x354 &  x382 & ~x0 & ~x6 & ~x14 & ~x31 & ~x76 & ~x104 & ~x117 & ~x127 & ~x202 & ~x307 & ~x386 & ~x395 & ~x477 & ~x614 & ~x692 & ~x723 & ~x759;
assign c5245 =  x152 &  x349 & ~x2 & ~x76 & ~x168 & ~x262 & ~x290 & ~x316 & ~x614 & ~x722 & ~x755;
assign c5247 =  x327 &  x355 & ~x14 & ~x34 & ~x104 & ~x116 & ~x121 & ~x123 & ~x151 & ~x202 & ~x350 & ~x421 & ~x424 & ~x472 & ~x527 & ~x560 & ~x634 & ~x729 & ~x744;
assign c5249 =  x326 &  x408 & ~x96 & ~x249 & ~x418 & ~x426 & ~x500 & ~x527 & ~x530 & ~x693 & ~x697 & ~x703;
assign c5251 = ~x46 & ~x292 & ~x319 & ~x347 & ~x348 & ~x374 & ~x375 & ~x403 & ~x464;
assign c5253 =  x414;
assign c5255 =  x257 &  x295 &  x495;
assign c5257 =  x429 &  x484 &  x512 &  x540 &  x597 & ~x23 & ~x31 & ~x81 & ~x83 & ~x85 & ~x169 & ~x277 & ~x279 & ~x367 & ~x390 & ~x528 & ~x739 & ~x744;
assign c5259 =  x462 &  x517 & ~x20 & ~x115 & ~x164 & ~x371 & ~x387 & ~x445 & ~x555 & ~x592 & ~x594 & ~x692 & ~x693 & ~x780;
assign c5261 = ~x4 & ~x5 & ~x22 & ~x30 & ~x36 & ~x37 & ~x57 & ~x79 & ~x85 & ~x86 & ~x90 & ~x91 & ~x115 & ~x140 & ~x145 & ~x191 & ~x213 & ~x222 & ~x280 & ~x301 & ~x367 & ~x418 & ~x425 & ~x504 & ~x512 & ~x538 & ~x555 & ~x570 & ~x571 & ~x582 & ~x596 & ~x620 & ~x627 & ~x651 & ~x654 & ~x655 & ~x657 & ~x678 & ~x684 & ~x693 & ~x706 & ~x707 & ~x765;
assign c5263 = ~x128 & ~x218 & ~x375 & ~x376 & ~x403 & ~x404 & ~x652 & ~x682;
assign c5265 =  x386;
assign c5267 = ~x51 & ~x79 & ~x102 & ~x114 & ~x128 & ~x134 & ~x144 & ~x159 & ~x165 & ~x168 & ~x169 & ~x215 & ~x224 & ~x226 & ~x280 & ~x281 & ~x312 & ~x334 & ~x385 & ~x448 & ~x455 & ~x456 & ~x482 & ~x485 & ~x512 & ~x538 & ~x542 & ~x590 & ~x592 & ~x617 & ~x624 & ~x627 & ~x637 & ~x654 & ~x655 & ~x683 & ~x693 & ~x698 & ~x711 & ~x712 & ~x724 & ~x735 & ~x744 & ~x762 & ~x764 & ~x767 & ~x770 & ~x776 & ~x777 & ~x779 & ~x782;
assign c5269 =  x429 &  x456 &  x457 &  x484 &  x540 & ~x77 & ~x194 & ~x752 & ~x767;
assign c5271 =  x295 &  x378 & ~x18 & ~x49 & ~x162 & ~x167 & ~x252 & ~x276 & ~x293 & ~x304 & ~x398 & ~x416 & ~x454 & ~x477 & ~x568 & ~x587 & ~x707 & ~x727;
assign c5273 =  x458 &  x486 &  x514 &  x571 & ~x169;
assign c5275 =  x387;
assign c5277 =  x431 &  x458 &  x486 &  x514 & ~x6 & ~x10 & ~x45 & ~x49 & ~x67 & ~x70 & ~x91 & ~x112 & ~x140 & ~x197 & ~x230 & ~x277 & ~x361 & ~x393 & ~x450 & ~x476 & ~x506 & ~x534 & ~x561 & ~x585 & ~x613 & ~x620 & ~x651 & ~x723 & ~x733 & ~x744 & ~x753 & ~x776 & ~x780;
assign c5279 =  x325 &  x408 & ~x20 & ~x25 & ~x42 & ~x91 & ~x102 & ~x106 & ~x142 & ~x169 & ~x254 & ~x305 & ~x341 & ~x386 & ~x445 & ~x483 & ~x665 & ~x671 & ~x699 & ~x750 & ~x755 & ~x760 & ~x763 & ~x772;
assign c5281 =  x358 & ~x378;
assign c5283 =  x358 & ~x353;
assign c5285 =  x325 &  x326 &  x380 & ~x1 & ~x19 & ~x277 & ~x305 & ~x309 & ~x400 & ~x416 & ~x422 & ~x424 & ~x581 & ~x693 & ~x764 & ~x772 & ~x780;
assign c5287 =  x353 &  x434 &  x462;
assign c5289 =  x269 &  x295 &  x348 &  x522 & ~x20 & ~x56 & ~x59 & ~x60 & ~x62 & ~x72 & ~x76 & ~x78 & ~x82 & ~x83 & ~x103 & ~x109 & ~x116 & ~x117 & ~x134 & ~x145 & ~x195 & ~x224 & ~x283 & ~x305 & ~x312 & ~x313 & ~x338 & ~x366 & ~x370 & ~x421 & ~x423 & ~x504 & ~x539 & ~x618 & ~x670 & ~x737 & ~x740 & ~x759 & ~x780;
assign c5291 =  x357 & ~x78 & ~x148 & ~x749;
assign c5293 =  x152 &  x295 & ~x20 & ~x57 & ~x112 & ~x114 & ~x139 & ~x144 & ~x219 & ~x262 & ~x263 & ~x394 & ~x417 & ~x491 & ~x555 & ~x648 & ~x689 & ~x772;
assign c5295 =  x326 &  x407 & ~x40 & ~x413 & ~x418 & ~x455 & ~x537;
assign c5297 =  x125 & ~x194 & ~x264;
assign c5299 =  x381 &  x409 & ~x111 & ~x157 & ~x452 & ~x502 & ~x540 & ~x542 & ~x568 & ~x582 & ~x599 & ~x626 & ~x680 & ~x709 & ~x750;
assign c60 =  x156 &  x265 & ~x162 & ~x263;
assign c62 =  x403 &  x431 & ~x147 & ~x204 & ~x214 & ~x240 & ~x241 & ~x267 & ~x268 & ~x299 & ~x315 & ~x392 & ~x420 & ~x451 & ~x583 & ~x625 & ~x729;
assign c64 =  x316 & ~x211 & ~x238 & ~x239 & ~x402 & ~x687;
assign c66 =  x317 &  x372 &  x428 &  x456 &  x457 &  x605 & ~x272 & ~x362;
assign c68 =  x156 &  x236 &  x291 &  x346 &  x373 &  x374 &  x496 &  x524 & ~x105 & ~x500 & ~x735;
assign c610 =  x549 &  x574 & ~x42 & ~x185 & ~x190 & ~x211 & ~x212 & ~x239 & ~x266 & ~x267;
assign c612 =  x126 &  x288 &  x399 & ~x162 & ~x211 & ~x239;
assign c614 = ~x127 & ~x157 & ~x183 & ~x184 & ~x185 & ~x186 & ~x211 & ~x212 & ~x214 & ~x215 & ~x238 & ~x239 & ~x240 & ~x266 & ~x267 & ~x274 & ~x654 & ~x656 & ~x684;
assign c616 =  x601 & ~x127 & ~x158 & ~x159 & ~x183 & ~x184 & ~x188 & ~x211 & ~x212 & ~x213 & ~x238 & ~x265 & ~x450 & ~x619 & ~x661 & ~x748;
assign c620 =  x237 &  x291 &  x318 &  x428 &  x630 & ~x151 & ~x196 & ~x334 & ~x364 & ~x588;
assign c622 =  x155 &  x290 &  x317 &  x318 &  x345 &  x401 &  x515 &  x631 & ~x147 & ~x190 & ~x426;
assign c624 =  x235 &  x262 &  x289 &  x290 &  x317 &  x318 &  x345 &  x401 & ~x211 & ~x238 & ~x239 & ~x240 & ~x241 & ~x266 & ~x654;
assign c626 =  x133 & ~x130;
assign c628 =  x320 &  x403 & ~x180 & ~x207 & ~x290 & ~x427;
assign c630 =  x237 &  x264 & ~x111 & ~x161 & ~x206 & ~x212 & ~x239 & ~x240 & ~x243 & ~x247 & ~x257 & ~x266 & ~x315 & ~x472 & ~x558 & ~x625 & ~x680;
assign c632 =  x415 & ~x184 & ~x212 & ~x264 & ~x290;
assign c634 =  x321 &  x404 &  x432 & ~x180 & ~x207 & ~x215 & ~x235 & ~x242 & ~x263 & ~x269 & ~x290 & ~x291 & ~x326 & ~x389 & ~x633;
assign c636 =  x89;
assign c638 =  x387 & ~x186 & ~x290;
assign c640 =  x359 & ~x346;
assign c642 = ~x17 & ~x156 & ~x184 & ~x185 & ~x186 & ~x211 & ~x212 & ~x213 & ~x214 & ~x215 & ~x216 & ~x238 & ~x239 & ~x240 & ~x265 & ~x349 & ~x376 & ~x655 & ~x657;
assign c644 =  x92;
assign c646 =  x211 &  x265 &  x402 & ~x13 & ~x41 & ~x54 & ~x154 & ~x208 & ~x269 & ~x307 & ~x337 & ~x528 & ~x594 & ~x636 & ~x652 & ~x687 & ~x693;
assign c648 =  x321 &  x456 & ~x209 & ~x301;
assign c650 =  x478;
assign c652 =  x387 & ~x240 & ~x292;
assign c654 =  x132 &  x159 &  x213 & ~x208 & ~x209;
assign c656 =  x415 & ~x212;
assign c658 =  x574 &  x605 & ~x60 & ~x63 & ~x184 & ~x185 & ~x186 & ~x188 & ~x202 & ~x212 & ~x239 & ~x312 & ~x508 & ~x623 & ~x625 & ~x638 & ~x664;
assign c660 =  x187 &  x214 &  x321 & ~x152 & ~x182 & ~x207 & ~x289 & ~x752;
assign c662 = ~x51 & ~x55 & ~x158 & ~x171 & ~x183 & ~x184 & ~x185 & ~x187 & ~x211 & ~x212 & ~x237 & ~x238 & ~x239 & ~x265 & ~x266 & ~x293 & ~x320 & ~x376 & ~x389 & ~x620 & ~x637 & ~x656 & ~x687;
assign c664 =  x441 &  x545 & ~x131 & ~x157 & ~x212 & ~x624;
assign c666 =  x375 &  x403 & ~x93 & ~x187 & ~x213 & ~x267 & ~x268 & ~x294 & ~x530 & ~x567 & ~x568 & ~x583 & ~x586 & ~x596 & ~x609 & ~x751;
assign c668 =  x487 & ~x65 & ~x184 & ~x186 & ~x212 & ~x238 & ~x239 & ~x478 & ~x589 & ~x628 & ~x686 & ~x687;
assign c670 =  x574 & ~x184 & ~x211 & ~x212 & ~x237 & ~x239 & ~x264 & ~x292 & ~x656;
assign c672 =  x105 & ~x181;
assign c674 =  x413 &  x440 &  x521 &  x547 & ~x241;
assign c676 =  x104 & ~x154;
assign c678 = ~x212 & ~x239;
assign c680 =  x401 &  x485 & ~x28 & ~x55 & ~x76 & ~x82 & ~x107 & ~x162 & ~x174 & ~x214 & ~x216 & ~x217 & ~x240 & ~x241 & ~x242 & ~x268 & ~x362 & ~x369 & ~x422 & ~x451 & ~x509 & ~x566 & ~x592 & ~x656 & ~x664 & ~x688 & ~x697 & ~x738 & ~x748;
assign c682 =  x387 & ~x292 & ~x320 & ~x459;
assign c684 =  x75;
assign c686 =  x316 &  x426 & ~x241;
assign c688 = ~x16 & ~x45 & ~x158 & ~x164 & ~x185 & ~x188 & ~x212 & ~x214 & ~x226 & ~x238 & ~x239 & ~x241 & ~x242 & ~x266 & ~x267 & ~x293 & ~x294 & ~x295 & ~x311 & ~x321 & ~x335 & ~x360 & ~x389 & ~x405 & ~x449 & ~x480 & ~x561 & ~x566 & ~x655 & ~x656 & ~x687 & ~x741 & ~x747 & ~x760;
assign c690 =  x371;
assign c692 =  x320 &  x428 &  x456 &  x568 &  x597 & ~x125 & ~x207 & ~x587;
assign c694 =  x574 & ~x99 & ~x157 & ~x208 & ~x211 & ~x236 & ~x264 & ~x292 & ~x347;
assign c698 =  x78;
assign c6100 = ~x147 & ~x188 & ~x212 & ~x215 & ~x242 & ~x266 & ~x599 & ~x659 & ~x693;
assign c6102 =  x156 &  x290 &  x317 &  x372 &  x400 &  x428 & ~x143 & ~x331 & ~x586;
assign c6104 =  x750;
assign c6106 =  x127 & ~x131 & ~x186 & ~x212 & ~x214 & ~x239 & ~x241;
assign c6108 =  x321 &  x376 &  x403 & ~x237 & ~x264 & ~x291 & ~x327 & ~x583;
assign c6110 =  x320 &  x494 & ~x47 & ~x240 & ~x267;
assign c6112 =  x132 &  x213 & ~x207 & ~x208 & ~x263;
assign c6114 =  x107;
assign c6116 =  x415 & ~x134 & ~x266 & ~x347 & ~x661;
assign c6118 =  x132 &  x267 & ~x61 & ~x115 & ~x180 & ~x207 & ~x301;
assign c6120 =  x101 &  x156;
assign c6122 =  x266 &  x293 & ~x152 & ~x153 & ~x180 & ~x190 & ~x205 & ~x207 & ~x236 & ~x269 & ~x297 & ~x299 & ~x318 & ~x661;
assign c6124 =  x102 &  x266;
assign c6126 =  x237 &  x403 & ~x207 & ~x239 & ~x242;
assign c6128 =  x126 & ~x63 & ~x105 & ~x129 & ~x162 & ~x186 & ~x187 & ~x188 & ~x190 & ~x200 & ~x213 & ~x214 & ~x216 & ~x217 & ~x240 & ~x241 & ~x242 & ~x329 & ~x331 & ~x479 & ~x534 & ~x596 & ~x648 & ~x715;
assign c6130 =  x291 &  x402 &  x431 &  x515 & ~x135 & ~x242 & ~x609 & ~x626 & ~x751;
assign c6132 =  x156 &  x291 &  x318 &  x373 &  x401 &  x551 & ~x123 & ~x269 & ~x756;
assign c6134 =  x101 & ~x215 & ~x216;
assign c6136 = ~x158 & ~x185 & ~x187 & ~x188 & ~x212 & ~x214 & ~x238 & ~x239 & ~x240 & ~x266 & ~x293 & ~x294 & ~x346 & ~x375 & ~x431 & ~x620;
assign c6138 =  x266 &  x293 &  x321 &  x515 & ~x207 & ~x242 & ~x269;
assign c6140 =  x552 & ~x239 & ~x241 & ~x266 & ~x267 & ~x268 & ~x271 & ~x294 & ~x320 & ~x375 & ~x559 & ~x637;
assign c6142 =  x408 &  x414 & ~x656;
assign c6144 =  x106 &  x374 &  x456 &  x484;
assign c6146 =  x108;
assign c6148 =  x104;
assign c6150 =  x116;
assign c6152 =  x359 &  x370 & ~x263 & ~x402;
assign c6154 =  x83;
assign c6156 =  x402 &  x467 & ~x151 & ~x207 & ~x242 & ~x261;
assign c6158 =  x267 &  x321 &  x431 &  x459 &  x547 & ~x153 & ~x154 & ~x207 & ~x209 & ~x234 & ~x263 & ~x278 & ~x335 & ~x760 & ~x773;
assign c6160 =  x413 &  x456 &  x547 & ~x186 & ~x187 & ~x214 & ~x215 & ~x241 & ~x243 & ~x275 & ~x641 & ~x656 & ~x660 & ~x694 & ~x760;
assign c6162 =  x75;
assign c6164 =  x343 &  x427 &  x499 & ~x659;
assign c6166 =  x63;
assign c6168 =  x320 &  x374 &  x431 &  x599 &  x631 & ~x38 & ~x152 & ~x327;
assign c6170 =  x290 &  x440 & ~x144 & ~x187 & ~x265 & ~x266 & ~x293 & ~x362 & ~x376 & ~x656 & ~x724 & ~x725;
assign c6172 =  x605 &  x606 & ~x162 & ~x184 & ~x185 & ~x200 & ~x211 & ~x212 & ~x239 & ~x241 & ~x266;
assign c6174 =  x129 &  x291 &  x318 &  x345 &  x630;
assign c6176 =  x494 &  x521 &  x574 & ~x187 & ~x212 & ~x266;
assign c6178 =  x186 & ~x182 & ~x209;
assign c6180 =  x574 & ~x184 & ~x212 & ~x215 & ~x216 & ~x239 & ~x266 & ~x320;
assign c6182 =  x94;
assign c6184 =  x399 &  x511 & ~x242 & ~x347;
assign c6186 =  x128 &  x318 &  x345 &  x401 & ~x232 & ~x287 & ~x656;
assign c6188 =  x359;
assign c6190 =  x159 &  x293 &  x403 & ~x207 & ~x290;
assign c6192 =  x431 &  x516 &  x574 & ~x242 & ~x268 & ~x389;
assign c6194 =  x404 &  x516 &  x544 & ~x136 & ~x215 & ~x221 & ~x262 & ~x268 & ~x298;
assign c6196 =  x545 & ~x24 & ~x37 & ~x184 & ~x185 & ~x189 & ~x212 & ~x213 & ~x214 & ~x215 & ~x221 & ~x239 & ~x266 & ~x267 & ~x294 & ~x333 & ~x450 & ~x656 & ~x692 & ~x747;
assign c6198 =  x402 &  x485 &  x597 & ~x207 & ~x453;
assign c6200 =  x238 &  x265 &  x320 & ~x112 & ~x167 & ~x180 & ~x188 & ~x205 & ~x208 & ~x245 & ~x268 & ~x502 & ~x640 & ~x651 & ~x740;
assign c6202 =  x321 &  x431 &  x460 & ~x208 & ~x290 & ~x291 & ~x318 & ~x325;
assign c6204 =  x321 &  x376 &  x574 & ~x117 & ~x196 & ~x205 & ~x207 & ~x209 & ~x235 & ~x261 & ~x263 & ~x299 & ~x307 & ~x310 & ~x329 & ~x443 & ~x477 & ~x501 & ~x674 & ~x706;
assign c6206 =  x237 &  x320 &  x571 & ~x34 & ~x190 & ~x207 & ~x235 & ~x242 & ~x250 & ~x368 & ~x502 & ~x562 & ~x583 & ~x624 & ~x704 & ~x776;
assign c6208 =  x320 &  x431 &  x515 & ~x134 & ~x151 & ~x269;
assign c6210 =  x410 &  x411 &  x440 &  x467 &  x468 & ~x245 & ~x300 & ~x327;
assign c6212 =  x262 &  x289 &  x317 &  x572 &  x574 & ~x186 & ~x215 & ~x216 & ~x265 & ~x304;
assign c6214 =  x103 & ~x126;
assign c6216 =  x459 &  x460 &  x487 & ~x151 & ~x242 & ~x243 & ~x268 & ~x288 & ~x470 & ~x719;
assign c6218 =  x676;
assign c6220 =  x321 &  x574 & ~x237 & ~x264 & ~x265 & ~x620 & ~x657 & ~x658;
assign c6222 =  x263 &  x318 &  x372 &  x598 & ~x241 & ~x507;
assign c6224 =  x320 &  x403 & ~x215 & ~x240 & ~x242 & ~x267;
assign c6226 =  x92;
assign c6228 =  x131 &  x158 & ~x152 & ~x188 & ~x208;
assign c6230 =  x403 &  x431 &  x488 &  x516 &  x521 & ~x202 & ~x215 & ~x222 & ~x230 & ~x241;
assign c6232 = ~x185 & ~x209 & ~x211 & ~x212 & ~x237 & ~x239 & ~x264 & ~x266;
assign c6234 =  x322 &  x404 &  x431 &  x574 & ~x151 & ~x264 & ~x265 & ~x420;
assign c6236 =  x293 &  x321 & ~x187 & ~x190 & ~x208 & ~x235 & ~x241 & ~x296 & ~x318 & ~x346 & ~x480 & ~x672;
assign c6238 =  x290 &  x345 &  x483 &  x511 &  x569 & ~x204 & ~x271 & ~x673 & ~x781;
assign c6240 =  x441 & ~x187 & ~x211 & ~x212 & ~x266 & ~x292;
assign c6242 =  x122 &  x329 & ~x184 & ~x211;
assign c6244 =  x267 &  x294 &  x403 &  x404 &  x431 &  x487 &  x574 & ~x207 & ~x261 & ~x289;
assign c6246 =  x186 &  x240 &  x294 &  x322 & ~x180 & ~x192 & ~x208 & ~x260 & ~x273 & ~x297 & ~x389 & ~x479;
assign c6248 =  x317 &  x400 &  x484 & ~x21 & ~x51 & ~x188 & ~x195 & ~x214 & ~x215 & ~x230 & ~x240 & ~x241 & ~x336 & ~x503 & ~x622 & ~x719 & ~x764;
assign c6250 =  x576 & ~x188 & ~x211 & ~x212 & ~x214 & ~x238 & ~x239 & ~x241 & ~x266 & ~x267 & ~x655;
assign c6252 =  x290 &  x318 &  x346 &  x374 &  x485 &  x606 &  x632 &  x633 & ~x271;
assign c6254 =  x77;
assign c6256 =  x574 & ~x132 & ~x184 & ~x185 & ~x211 & ~x212 & ~x237 & ~x239 & ~x265 & ~x266 & ~x292 & ~x624;
assign c6258 =  x133 &  x160 &  x456;
assign c6260 =  x294 &  x431 &  x515 & ~x77 & ~x137 & ~x179 & ~x208 & ~x291 & ~x417;
assign c6262 =  x321 &  x404 & ~x152 & ~x208 & ~x242 & ~x264 & ~x346 & ~x612 & ~x687;
assign c6264 =  x291 &  x319 &  x346 &  x429 &  x485 & ~x32 & ~x43 & ~x50 & ~x122 & ~x214 & ~x232 & ~x242 & ~x270 & ~x272 & ~x276 & ~x537 & ~x693 & ~x717 & ~x742;
assign c6266 =  x400 &  x522 &  x568 & ~x152;
assign c6268 =  x98 &  x126 & ~x177 & ~x212;
assign c6270 =  x574 & ~x131 & ~x184 & ~x188 & ~x212 & ~x214 & ~x239 & ~x265 & ~x266 & ~x320 & ~x656 & ~x659;
assign c6272 =  x316 &  x399 &  x455 &  x483 &  x552 & ~x271 & ~x331 & ~x474 & ~x686;
assign c6274 =  x102 & ~x299;
assign c6276 =  x100 & ~x65 & ~x88 & ~x188 & ~x214 & ~x269 & ~x295 & ~x314;
assign c6278 =  x496 &  x576 & ~x158 & ~x183 & ~x188 & ~x212 & ~x238 & ~x239;
assign c6280 =  x291 &  x319 &  x403 &  x431 &  x459 & ~x177 & ~x244 & ~x294 & ~x655;
assign c6282 =  x163 & ~x236;
assign c6284 =  x75;
assign c6286 =  x322 &  x404 &  x431 & ~x70 & ~x154 & ~x176 & ~x207 & ~x208 & ~x209 & ~x230 & ~x235 & ~x264 & ~x289 & ~x306 & ~x383 & ~x392 & ~x479 & ~x591 & ~x743;
assign c6288 =  x291 &  x374 &  x375 &  x401 &  x514 & ~x178 & ~x241 & ~x267 & ~x268 & ~x343 & ~x507 & ~x652;
assign c6290 =  x458 &  x574 & ~x184 & ~x185 & ~x238 & ~x264;
assign c6292 =  x291 &  x319 &  x347 &  x431 &  x458 &  x459 &  x600 &  x631 & ~x3 & ~x145 & ~x177 & ~x298 & ~x329 & ~x480 & ~x596 & ~x685 & ~x775;
assign c6294 =  x129 & ~x162 & ~x207 & ~x208 & ~x241 & ~x392 & ~x624 & ~x721;
assign c6296 =  x320 &  x514 & ~x207 & ~x230 & ~x260 & ~x261 & ~x269 & ~x271 & ~x299 & ~x331 & ~x397 & ~x424 & ~x480 & ~x595 & ~x596 & ~x620 & ~x686 & ~x688 & ~x704 & ~x724;
assign c6298 =  x127 &  x289 &  x400 &  x606 & ~x266;
assign c61 =  x217 & ~x38 & ~x120 & ~x362 & ~x388 & ~x584 & ~x631 & ~x643 & ~x691 & ~x782;
assign c63 = ~x129 & ~x226 & ~x313 & ~x521 & ~x575 & ~x602 & ~x603 & ~x630;
assign c65 =  x658 & ~x67 & ~x101 & ~x199 & ~x245 & ~x421 & ~x429 & ~x467 & ~x531 & ~x667;
assign c67 =  x350 & ~x20 & ~x430 & ~x461;
assign c69 =  x242 & ~x30 & ~x95 & ~x406 & ~x461 & ~x463 & ~x490 & ~x752;
assign c611 =  x270 &  x297 &  x298 &  x326 & ~x653;
assign c613 =  x518 &  x540 & ~x356 & ~x601;
assign c615 =  x684;
assign c617 =  x206 &  x658 & ~x12 & ~x32 & ~x57 & ~x73 & ~x94 & ~x96 & ~x100 & ~x101 & ~x175 & ~x337 & ~x388 & ~x484 & ~x526 & ~x642 & ~x666 & ~x733 & ~x780;
assign c619 =  x270 &  x325 & ~x0 & ~x7 & ~x15 & ~x29 & ~x33 & ~x45 & ~x49 & ~x75 & ~x80 & ~x85 & ~x91 & ~x106 & ~x112 & ~x114 & ~x115 & ~x170 & ~x367 & ~x394 & ~x442 & ~x502 & ~x504 & ~x531 & ~x589 & ~x619 & ~x651 & ~x677 & ~x698 & ~x703 & ~x705 & ~x717 & ~x722 & ~x730 & ~x739 & ~x759 & ~x767;
assign c621 = ~x92 & ~x223 & ~x514 & ~x515 & ~x516 & ~x541 & ~x542;
assign c623 = ~x541 & ~x542 & ~x543 & ~x544 & ~x545;
assign c625 =  x657 & ~x3 & ~x10 & ~x59 & ~x112 & ~x140 & ~x167 & ~x191 & ~x243 & ~x274 & ~x283 & ~x310 & ~x362 & ~x389 & ~x390 & ~x423 & ~x457 & ~x472 & ~x474 & ~x483 & ~x485 & ~x506 & ~x511 & ~x555 & ~x564 & ~x638 & ~x646 & ~x670 & ~x695 & ~x713 & ~x714 & ~x744 & ~x753 & ~x757 & ~x759 & ~x763 & ~x764 & ~x771 & ~x777;
assign c627 = ~x515 & ~x516 & ~x541 & ~x542 & ~x543 & ~x563 & ~x614;
assign c629 = ~x492 & ~x520 & ~x576 & ~x631;
assign c631 =  x301 &  x302 & ~x379 & ~x380 & ~x418;
assign c633 =  x216 &  x301;
assign c635 =  x178 &  x181 & ~x15 & ~x47 & ~x65 & ~x87 & ~x95 & ~x96 & ~x101 & ~x244 & ~x253 & ~x448 & ~x450 & ~x454 & ~x646 & ~x671 & ~x693 & ~x717 & ~x743;
assign c637 = ~x492 & ~x494 & ~x504 & ~x520 & ~x522 & ~x524 & ~x549 & ~x605;
assign c639 =  x462 & ~x424 & ~x520 & ~x521 & ~x550 & ~x604 & ~x633;
assign c641 = ~x72 & ~x370 & ~x388 & ~x485 & ~x489 & ~x514 & ~x515 & ~x516 & ~x517 & ~x518 & ~x620;
assign c643 =  x239 &  x296 &  x378 & ~x88 & ~x159 & ~x364 & ~x422 & ~x439;
assign c645 =  x269 &  x352 &  x380 &  x409 &  x436 &  x437 & ~x328 & ~x329;
assign c647 =  x243 &  x271 &  x299 & ~x147 & ~x176 & ~x688 & ~x750;
assign c649 =  x242 &  x270 & ~x7 & ~x10 & ~x19 & ~x25 & ~x26 & ~x38 & ~x46 & ~x47 & ~x59 & ~x60 & ~x74 & ~x106 & ~x118 & ~x121 & ~x141 & ~x194 & ~x224 & ~x231 & ~x248 & ~x257 & ~x285 & ~x332 & ~x340 & ~x341 & ~x369 & ~x393 & ~x473 & ~x480 & ~x501 & ~x530 & ~x563 & ~x565 & ~x584 & ~x618 & ~x640 & ~x691 & ~x716 & ~x728 & ~x753 & ~x764;
assign c651 =  x538 &  x542 & ~x373;
assign c653 =  x303 & ~x606;
assign c655 =  x462 & ~x332 & ~x543 & ~x570 & ~x571;
assign c657 =  x247;
assign c659 = ~x158 & ~x541 & ~x542 & ~x543 & ~x549;
assign c661 =  x216 &  x355;
assign c663 =  x325 & ~x8 & ~x12 & ~x37 & ~x38 & ~x48 & ~x75 & ~x77 & ~x121 & ~x200 & ~x250 & ~x343 & ~x369 & ~x411 & ~x418 & ~x467 & ~x468 & ~x475 & ~x533 & ~x557 & ~x590 & ~x685 & ~x737 & ~x742;
assign c665 = ~x96 & ~x108 & ~x116 & ~x122 & ~x251 & ~x279 & ~x308 & ~x369 & ~x458 & ~x483 & ~x484 & ~x485 & ~x487 & ~x514 & ~x563 & ~x737 & ~x773;
assign c667 = ~x494 & ~x541 & ~x542 & ~x576 & ~x606;
assign c669 =  x154 &  x406 &  x435 & ~x411 & ~x466 & ~x467 & ~x476 & ~x498 & ~x591 & ~x608;
assign c671 =  x245 &  x273 &  x301 & ~x379;
assign c673 = ~x513 & ~x517 & ~x543 & ~x544;
assign c675 =  x352 &  x380 &  x407 & ~x5 & ~x17 & ~x20 & ~x50 & ~x65 & ~x67 & ~x75 & ~x77 & ~x83 & ~x108 & ~x141 & ~x144 & ~x146 & ~x150 & ~x167 & ~x231 & ~x308 & ~x309 & ~x359 & ~x441 & ~x445 & ~x530 & ~x565 & ~x640 & ~x644 & ~x710 & ~x736 & ~x760 & ~x779 & ~x783;
assign c677 = ~x408 & ~x433 & ~x434 & ~x463;
assign c679 =  x436 &  x437 & ~x100 & ~x522 & ~x570;
assign c681 = ~x12 & ~x114 & ~x253 & ~x305 & ~x338 & ~x339 & ~x547 & ~x575 & ~x576 & ~x603 & ~x604 & ~x631 & ~x697 & ~x757 & ~x777;
assign c683 =  x242 & ~x11 & ~x14 & ~x16 & ~x23 & ~x42 & ~x82 & ~x89 & ~x108 & ~x115 & ~x150 & ~x176 & ~x177 & ~x227 & ~x313 & ~x338 & ~x339 & ~x479 & ~x486 & ~x563 & ~x666 & ~x691 & ~x694 & ~x704 & ~x770;
assign c685 =  x245 & ~x378 & ~x379 & ~x631;
assign c687 =  x355 &  x383 & ~x14 & ~x67 & ~x142 & ~x352 & ~x379 & ~x380 & ~x441 & ~x767;
assign c689 =  x274 & ~x379;
assign c691 =  x653 & ~x2 & ~x94 & ~x101 & ~x250 & ~x370 & ~x695 & ~x775;
assign c693 =  x177 &  x178 & ~x1 & ~x5 & ~x26 & ~x32 & ~x42 & ~x47 & ~x49 & ~x69 & ~x228 & ~x251 & ~x273 & ~x333 & ~x341 & ~x356 & ~x359 & ~x423 & ~x446 & ~x480 & ~x504 & ~x651 & ~x652;
assign c695 = ~x406 & ~x407 & ~x408 & ~x433 & ~x434 & ~x435 & ~x461 & ~x462 & ~x463 & ~x489 & ~x492 & ~x506;
assign c697 =  x356 & ~x199 & ~x381 & ~x405 & ~x406 & ~x407 & ~x408 & ~x409 & ~x433;
assign c699 =  x510 & ~x340 & ~x382 & ~x435 & ~x436 & ~x462 & ~x752;
assign c6101 =  x429 & ~x540 & ~x544 & ~x571;
assign c6103 =  x151 &  x178 &  x179 &  x183 & ~x385;
assign c6105 =  x566 & ~x429;
assign c6107 =  x246 &  x274;
assign c6109 = ~x545 & ~x571 & ~x600;
assign c6111 =  x149 &  x151 & ~x287 & ~x397;
assign c6113 = ~x350 & ~x379 & ~x380 & ~x381 & ~x406 & ~x407 & ~x433 & ~x434 & ~x435 & ~x461 & ~x462 & ~x463 & ~x489 & ~x491;
assign c6115 =  x243 &  x271 &  x409;
assign c6117 =  x123 &  x124 & ~x330 & ~x358 & ~x363 & ~x413;
assign c6119 =  x603 &  x655;
assign c6121 =  x206 &  x349 &  x350 & ~x2 & ~x96;
assign c6123 =  x464 & ~x570 & ~x605;
assign c6125 =  x323 & ~x520 & ~x575 & ~x576;
assign c6127 =  x217 &  x245 & ~x352;
assign c6129 =  x577 & ~x2 & ~x231 & ~x385 & ~x411 & ~x430 & ~x445 & ~x709;
assign c6131 =  x215 &  x243 &  x327 & ~x350 & ~x351;
assign c6133 =  x657 &  x658 &  x685;
assign c6135 = ~x353 & ~x433 & ~x436 & ~x461 & ~x462 & ~x463 & ~x489 & ~x492 & ~x493 & ~x517 & ~x518;
assign c6137 =  x270 &  x298 &  x325 & ~x30 & ~x31 & ~x32 & ~x53 & ~x68 & ~x77 & ~x82 & ~x91 & ~x93 & ~x96 & ~x114 & ~x145 & ~x192 & ~x196 & ~x219 & ~x227 & ~x283 & ~x306 & ~x309 & ~x357 & ~x358 & ~x365 & ~x395 & ~x591 & ~x617 & ~x622 & ~x667 & ~x691 & ~x724 & ~x733 & ~x741 & ~x773 & ~x775;
assign c6139 =  x684;
assign c6141 = ~x511 & ~x514 & ~x515 & ~x516 & ~x541 & ~x542 & ~x543 & ~x708;
assign c6143 = ~x97 & ~x108 & ~x118 & ~x169 & ~x246 & ~x251 & ~x309 & ~x551 & ~x570 & ~x571 & ~x572 & ~x638;
assign c6145 =  x652;
assign c6147 =  x461 & ~x72 & ~x339 & ~x520 & ~x552 & ~x576 & ~x577 & ~x579 & ~x604 & ~x716;
assign c6149 =  x622;
assign c6151 =  x271 &  x299 &  x382 & ~x350;
assign c6153 =  x206 &  x208 &  x233 & ~x408 & ~x584 & ~x712 & ~x734;
assign c6155 =  x242 &  x548 & ~x108 & ~x476 & ~x489;
assign c6157 = ~x430 & ~x433 & ~x434 & ~x435 & ~x461 & ~x462 & ~x463 & ~x489 & ~x492;
assign c6159 =  x299 &  x437 &  x438 & ~x172 & ~x251 & ~x279 & ~x311;
assign c6161 =  x178 &  x206 & ~x358 & ~x372;
assign c6163 =  x188 & ~x362 & ~x365 & ~x367 & ~x562 & ~x630 & ~x631 & ~x711;
assign c6165 =  x323 &  x406 & ~x136 & ~x189 & ~x357 & ~x410 & ~x437 & ~x465 & ~x466 & ~x467 & ~x484 & ~x584 & ~x593 & ~x777;
assign c6167 =  x593;
assign c6169 =  x433 &  x462 & ~x486 & ~x496 & ~x522;
assign c6171 = ~x94 & ~x351 & ~x379 & ~x381 & ~x407 & ~x408 & ~x433 & ~x434 & ~x435 & ~x461 & ~x462 & ~x463 & ~x487 & ~x491 & ~x648;
assign c6173 =  x217 &  x245 &  x273;
assign c6175 = ~x540 & ~x543 & ~x544 & ~x570 & ~x571;
assign c6177 =  x270 &  x298 &  x381 & ~x12 & ~x37 & ~x166 & ~x737;
assign c6179 = ~x67 & ~x228 & ~x280 & ~x357 & ~x396 & ~x430 & ~x489 & ~x776;
assign c6181 =  x622;
assign c6183 =  x296 & ~x396 & ~x601 & ~x602;
assign c6185 =  x462 &  x518 & ~x91 & ~x495 & ~x542 & ~x578;
assign c6187 =  x269 & ~x573 & ~x749;
assign c6189 =  x301 & ~x353 & ~x380 & ~x462;
assign c6191 =  x268 &  x296 &  x352 &  x380 & ~x357;
assign c6193 = ~x227 & ~x408 & ~x486 & ~x489 & ~x515 & ~x516 & ~x517;
assign c6195 =  x300 &  x409 &  x436 &  x437 & ~x120 & ~x541;
assign c6197 =  x406 &  x407 & ~x44 & ~x112 & ~x356 & ~x383 & ~x394 & ~x484 & ~x485 & ~x486 & ~x487;
assign c6199 =  x325 &  x463 & ~x572;
assign c6201 = ~x67 & ~x547 & ~x601 & ~x630;
assign c6203 = ~x105 & ~x118 & ~x408 & ~x409 & ~x436 & ~x467 & ~x493 & ~x494 & ~x495 & ~x520 & ~x522 & ~x591 & ~x699 & ~x750 & ~x757 & ~x764 & ~x779;
assign c6205 = ~x381 & ~x575 & ~x601 & ~x602 & ~x603 & ~x604;
assign c6207 =  x491 & ~x571 & ~x572 & ~x598;
assign c6209 = ~x337 & ~x454 & ~x461 & ~x462 & ~x489 & ~x515 & ~x516 & ~x517 & ~x526 & ~x608 & ~x746;
assign c6211 = ~x545 & ~x572 & ~x573 & ~x628;
assign c6213 = ~x20 & ~x146 & ~x170 & ~x355 & ~x362 & ~x411 & ~x600 & ~x601 & ~x757 & ~x766;
assign c6215 =  x125 &  x152 &  x154 &  x183 & ~x0 & ~x66 & ~x104 & ~x255 & ~x444 & ~x471 & ~x527 & ~x641 & ~x673 & ~x683;
assign c6217 =  x596 &  x625 & ~x428 & ~x457 & ~x497 & ~x706;
assign c6219 =  x566 &  x567 &  x595 &  x596 & ~x62 & ~x193 & ~x309 & ~x370 & ~x442 & ~x652 & ~x754;
assign c6221 =  x298 &  x353 & ~x356 & ~x413;
assign c6223 = ~x49 & ~x361 & ~x436 & ~x462 & ~x463 & ~x489 & ~x491 & ~x515 & ~x516 & ~x517 & ~x518 & ~x740;
assign c6225 =  x326 &  x435 &  x490 & ~x494 & ~x512 & ~x605;
assign c6227 =  x215 &  x300 &  x328;
assign c6229 =  x302 & ~x407 & ~x408;
assign c6231 =  x301 &  x302 & ~x352;
assign c6233 = ~x101 & ~x103 & ~x521 & ~x531 & ~x541 & ~x575 & ~x576 & ~x603 & ~x663 & ~x774;
assign c6235 =  x271 &  x299 &  x381;
assign c6237 =  x244 &  x300 &  x328 & ~x379;
assign c6239 =  x380 &  x596 & ~x385;
assign c6241 =  x178 &  x179 &  x203;
assign c6243 = ~x422 & ~x511 & ~x515 & ~x541 & ~x542 & ~x694;
assign c6245 =  x626 &  x627 & ~x429 & ~x456 & ~x483 & ~x545 & ~x667;
assign c6247 =  x624 & ~x425 & ~x517;
assign c6249 =  x270 &  x326 &  x354 & ~x16 & ~x32 & ~x44 & ~x144 & ~x197 & ~x224 & ~x251 & ~x341 & ~x417 & ~x533 & ~x565 & ~x640 & ~x678 & ~x780;
assign c6251 =  x300 &  x328 &  x355 & ~x73 & ~x253 & ~x352 & ~x423 & ~x527 & ~x584 & ~x651 & ~x672 & ~x737 & ~x762;
assign c6253 =  x123 &  x124 &  x125 &  x570 & ~x109 & ~x313 & ~x478 & ~x621 & ~x667 & ~x712;
assign c6255 =  x323 &  x380 &  x435 & ~x136;
assign c6257 =  x491 & ~x544 & ~x571;
assign c6259 =  x380 & ~x313 & ~x344 & ~x358 & ~x439;
assign c6261 = ~x52 & ~x75 & ~x78 & ~x99 & ~x308 & ~x313 & ~x388 & ~x397 & ~x461 & ~x462 & ~x485 & ~x489 & ~x515 & ~x517 & ~x589 & ~x706 & ~x733 & ~x767;
assign c6263 =  x298 &  x326 &  x354 &  x437 & ~x1 & ~x350 & ~x390 & ~x422 & ~x650;
assign c6265 =  x210 &  x323 & ~x21 & ~x38 & ~x75 & ~x99 & ~x104 & ~x107 & ~x328 & ~x356 & ~x357 & ~x382 & ~x584 & ~x675 & ~x677 & ~x709 & ~x754;
assign c6267 =  x300 &  x328 & ~x253 & ~x351 & ~x379 & ~x380;
assign c6269 =  x246 &  x274 & ~x43 & ~x446 & ~x714 & ~x744;
assign c6271 = ~x544 & ~x545 & ~x628;
assign c6273 =  x405 &  x407 & ~x487 & ~x515 & ~x541;
assign c6275 =  x154 &  x268 &  x297;
assign c6277 =  x184 &  x625 & ~x397;
assign c6279 =  x349 &  x378 &  x406 & ~x74 & ~x83 & ~x85 & ~x94 & ~x112 & ~x146 & ~x165 & ~x277 & ~x338 & ~x363 & ~x370 & ~x429 & ~x439 & ~x441 & ~x484 & ~x485 & ~x497 & ~x565 & ~x640 & ~x646 & ~x706 & ~x712 & ~x776;
assign c6281 =  x178 &  x179 & ~x93 & ~x218 & ~x363 & ~x388 & ~x546 & ~x619 & ~x701 & ~x731;
assign c6283 = ~x96 & ~x131 & ~x544 & ~x570 & ~x571;
assign c6285 =  x625 &  x626 &  x628 &  x654 & ~x2 & ~x220 & ~x565 & ~x584 & ~x737 & ~x757 & ~x780;
assign c6287 =  x570 & ~x1 & ~x33 & ~x38 & ~x56 & ~x96 & ~x100 & ~x112 & ~x120 & ~x369 & ~x397 & ~x440 & ~x441 & ~x457 & ~x458 & ~x468 & ~x485 & ~x486 & ~x497 & ~x533 & ~x669 & ~x699 & ~x728 & ~x745 & ~x782;
assign c6289 = ~x33 & ~x96 & ~x384 & ~x388 & ~x411 & ~x437 & ~x441 & ~x493 & ~x494 & ~x495 & ~x496 & ~x497 & ~x522 & ~x757;
assign c6291 =  x380 & ~x148 & ~x329 & ~x332 & ~x357 & ~x369 & ~x410 & ~x413 & ~x439 & ~x536;
assign c6293 =  x573 & ~x33 & ~x430 & ~x461 & ~x462 & ~x489 & ~x491 & ~x668;
assign c6295 =  x178 &  x179 &  x208 &  x209 & ~x477 & ~x646;
assign c6297 =  x274 & ~x631;
assign c6299 =  x299 &  x355 & ~x350 & ~x351 & ~x377 & ~x406 & ~x407 & ~x777;
assign c70 =  x297 &  x298 &  x407 &  x435 &  x462 & ~x18 & ~x42 & ~x60 & ~x114 & ~x122 & ~x138 & ~x150 & ~x151 & ~x158 & ~x160 & ~x193 & ~x220 & ~x249 & ~x254 & ~x275 & ~x361 & ~x366 & ~x371 & ~x390 & ~x391 & ~x397 & ~x412 & ~x415 & ~x416 & ~x450 & ~x497 & ~x520 & ~x521 & ~x522 & ~x524 & ~x549 & ~x551 & ~x555 & ~x558 & ~x563 & ~x575 & ~x576 & ~x589 & ~x602 & ~x603 & ~x604 & ~x634 & ~x646 & ~x667 & ~x694;
assign c72 =  x180 &  x185 &  x212 &  x489 &  x573 & ~x316 & ~x690;
assign c74 =  x236 &  x238 &  x240 &  x406 &  x489 &  x544 & ~x549 & ~x582 & ~x604 & ~x634;
assign c76 =  x233 &  x261 &  x264 &  x266 &  x267 &  x464 & ~x156;
assign c78 =  x668;
assign c710 =  x235 &  x517 & ~x159 & ~x316 & ~x319 & ~x332 & ~x348 & ~x454 & ~x575 & ~x576 & ~x630 & ~x662 & ~x775;
assign c712 = ~x406 & ~x434 & ~x436 & ~x488 & ~x571 & ~x598 & ~x624;
assign c714 =  x717;
assign c716 =  x270 &  x545 &  x684 &  x712 & ~x61 & ~x529 & ~x580 & ~x621 & ~x645;
assign c718 =  x321 &  x355 & ~x629;
assign c720 =  x239 &  x407 &  x411 & ~x315 & ~x550 & ~x635;
assign c722 =  x210 &  x214 &  x243 &  x244 &  x270 & ~x576 & ~x580;
assign c724 =  x235 &  x238 &  x240 &  x324 &  x462 &  x489 & ~x522 & ~x527 & ~x607;
assign c726 =  x271 &  x299 &  x382 &  x464 & ~x33 & ~x190 & ~x406 & ~x433 & ~x434 & ~x489 & ~x570;
assign c728 =  x285;
assign c730 =  x213 &  x235 &  x236 &  x238 &  x269 &  x489 & ~x345 & ~x588;
assign c732 =  x438 &  x493 & ~x157 & ~x365 & ~x417 & ~x433 & ~x435 & ~x477 & ~x487 & ~x568 & ~x594 & ~x595 & ~x642;
assign c734 =  x518 &  x519 &  x574 &  x658 &  x686 & ~x14 & ~x77 & ~x89 & ~x99 & ~x102 & ~x108 & ~x116 & ~x122 & ~x140 & ~x172 & ~x193 & ~x215 & ~x219 & ~x227 & ~x243 & ~x271 & ~x285 & ~x306 & ~x361 & ~x391 & ~x395 & ~x400 & ~x418 & ~x452 & ~x505 & ~x508 & ~x527 & ~x531 & ~x571 & ~x582 & ~x609 & ~x625 & ~x636 & ~x651 & ~x681 & ~x718 & ~x739 & ~x742;
assign c736 =  x236 &  x239 &  x240 & ~x58 & ~x253 & ~x349 & ~x404 & ~x406 & ~x433 & ~x488 & ~x531 & ~x559 & ~x571 & ~x586 & ~x653 & ~x668 & ~x748;
assign c738 =  x270 &  x517 &  x544 &  x681 & ~x160;
assign c740 =  x338;
assign c742 =  x775;
assign c744 =  x62;
assign c746 = ~x153 & ~x160 & ~x183 & ~x230 & ~x358 & ~x406 & ~x433 & ~x434 & ~x439 & ~x488 & ~x522 & ~x540 & ~x549 & ~x597;
assign c748 = ~x60 & ~x147 & ~x157 & ~x183 & ~x184 & ~x226 & ~x275 & ~x334 & ~x433 & ~x434 & ~x441 & ~x488 & ~x522 & ~x542 & ~x571 & ~x595 & ~x606 & ~x614 & ~x623 & ~x625 & ~x705 & ~x708;
assign c750 =  x407 &  x489 &  x544 & ~x35 & ~x46 & ~x376 & ~x419 & ~x500 & ~x508 & ~x522 & ~x551 & ~x564 & ~x575 & ~x576 & ~x582 & ~x629 & ~x685 & ~x740 & ~x777;
assign c752 =  x209 &  x214 & ~x0 & ~x9 & ~x220 & ~x251 & ~x314 & ~x320 & ~x371 & ~x375 & ~x522 & ~x548 & ~x550 & ~x576 & ~x577 & ~x603 & ~x635 & ~x643 & ~x697 & ~x782;
assign c754 = ~x154 & ~x181 & ~x184 & ~x363 & ~x433 & ~x491 & ~x546;
assign c756 =  x715 & ~x119 & ~x155 & ~x404;
assign c758 =  x205 &  x206 &  x207 &  x464 &  x519 & ~x315 & ~x571 & ~x572 & ~x645 & ~x662;
assign c762 =  x205 &  x206 &  x519 & ~x0 & ~x219 & ~x284 & ~x315 & ~x319 & ~x414 & ~x445 & ~x533 & ~x554 & ~x571 & ~x623 & ~x655 & ~x700 & ~x741;
assign c764 =  x715 & ~x433;
assign c768 =  x269 &  x546 &  x574 &  x601 & ~x85 & ~x157 & ~x188 & ~x191 & ~x216 & ~x272 & ~x349 & ~x374 & ~x396 & ~x418 & ~x427 & ~x444 & ~x478 & ~x563 & ~x577 & ~x583 & ~x594 & ~x597 & ~x646 & ~x750 & ~x780;
assign c770 =  x288 &  x293 & ~x5 & ~x544 & ~x597;
assign c772 =  x185 &  x207 &  x545 & ~x80 & ~x161 & ~x292 & ~x310 & ~x320;
assign c774 =  x441 & ~x17 & ~x160 & ~x570 & ~x571 & ~x624 & ~x645;
assign c776 =  x438 &  x462 & ~x114 & ~x219 & ~x224 & ~x315 & ~x345 & ~x371 & ~x375 & ~x400 & ~x523 & ~x551 & ~x554;
assign c778 =  x7;
assign c780 =  x202 &  x548;
assign c782 =  x240 &  x489 & ~x72 & ~x80 & ~x116 & ~x117 & ~x130 & ~x134 & ~x172 & ~x174 & ~x287 & ~x316 & ~x320 & ~x321 & ~x332 & ~x371 & ~x419 & ~x510 & ~x522 & ~x523 & ~x537 & ~x549 & ~x575 & ~x576 & ~x592 & ~x596 & ~x603 & ~x604 & ~x662 & ~x666 & ~x690 & ~x769;
assign c784 =  x261 &  x264 &  x266 & ~x315 & ~x571 & ~x626;
assign c786 =  x321 & ~x183 & ~x211 & ~x237;
assign c788 =  x5;
assign c790 =  x710 & ~x602 & ~x603;
assign c792 =  x179 &  x242 &  x517 & ~x426 & ~x659;
assign c794 =  x493 &  x521 & ~x16 & ~x21 & ~x31 & ~x37 & ~x43 & ~x52 & ~x54 & ~x58 & ~x69 & ~x72 & ~x76 & ~x80 & ~x93 & ~x94 & ~x100 & ~x111 & ~x114 & ~x118 & ~x127 & ~x135 & ~x137 & ~x153 & ~x155 & ~x162 & ~x164 & ~x171 & ~x197 & ~x225 & ~x247 & ~x304 & ~x305 & ~x336 & ~x362 & ~x396 & ~x406 & ~x433 & ~x434 & ~x444 & ~x478 & ~x488 & ~x502 & ~x503 & ~x538 & ~x564 & ~x565 & ~x571 & ~x597 & ~x620 & ~x624 & ~x639 & ~x643 & ~x647 & ~x654 & ~x692 & ~x729 & ~x733 & ~x737 & ~x748 & ~x774 & ~x776 & ~x779;
assign c796 = ~x333 & ~x379 & ~x407 & ~x433 & ~x435 & ~x489 & ~x506 & ~x517 & ~x565 & ~x571 & ~x654 & ~x742;
assign c798 =  x242 &  x269 &  x491 & ~x81 & ~x99 & ~x109 & ~x217 & ~x330 & ~x418 & ~x433 & ~x542 & ~x569 & ~x576 & ~x592 & ~x640 & ~x670 & ~x690 & ~x731;
assign c7100 =  x260 &  x294 &  x519;
assign c7102 =  x742;
assign c7104 =  x169;
assign c7106 =  x214 &  x236 &  x240 & ~x292 & ~x575 & ~x603;
assign c7108 =  x272 & ~x406 & ~x418 & ~x433 & ~x445 & ~x488 & ~x597;
assign c7110 =  x677;
assign c7112 =  x293 &  x316 & ~x191 & ~x509 & ~x542 & ~x570 & ~x597 & ~x730;
assign c7114 =  x238 &  x239 &  x240 &  x435 &  x462 &  x463 & ~x89 & ~x218 & ~x243 & ~x280 & ~x299 & ~x326 & ~x327 & ~x333 & ~x555 & ~x565 & ~x598 & ~x624 & ~x625 & ~x681;
assign c7116 =  x235 &  x239 &  x240 &  x489 &  x517 &  x545 & ~x43 & ~x117 & ~x140 & ~x157 & ~x163 & ~x193 & ~x315 & ~x371 & ~x756;
assign c7118 =  x61;
assign c7120 = ~x351 & ~x433 & ~x435 & ~x488 & ~x573;
assign c7122 =  x18;
assign c7124 = ~x178 & ~x183 & ~x184 & ~x185 & ~x433 & ~x542 & ~x597;
assign c7126 =  x178 & ~x54 & ~x123 & ~x146 & ~x272 & ~x273 & ~x283 & ~x291 & ~x315 & ~x359 & ~x363 & ~x445 & ~x512 & ~x549 & ~x557 & ~x568 & ~x663 & ~x691;
assign c7128 =  x233 &  x240 &  x266 &  x462 & ~x5 & ~x28 & ~x337 & ~x371 & ~x503 & ~x594;
assign c7130 =  x462 &  x624 & ~x601;
assign c7132 =  x232 &  x233 &  x234 &  x235 &  x261 & ~x130 & ~x154 & ~x349 & ~x377 & ~x667 & ~x723 & ~x739 & ~x772;
assign c7134 = ~x82 & ~x184 & ~x406 & ~x433 & ~x488 & ~x517 & ~x518 & ~x571 & ~x597;
assign c7136 =  x271 &  x293 &  x295 &  x298 &  x325 & ~x80 & ~x183;
assign c7138 =  x704;
assign c7140 = ~x183 & ~x184 & ~x214 & ~x244 & ~x462 & ~x625;
assign c7142 =  x316 &  x320 & ~x651;
assign c7144 = ~x152 & ~x406 & ~x408 & ~x433 & ~x463 & ~x517 & ~x571 & ~x625;
assign c7146 =  x573 & ~x5 & ~x38 & ~x73 & ~x87 & ~x101 & ~x167 & ~x221 & ~x259 & ~x312 & ~x376 & ~x406 & ~x418 & ~x420 & ~x433 & ~x461 & ~x488 & ~x566 & ~x567 & ~x576 & ~x591 & ~x592 & ~x594 & ~x596 & ~x603 & ~x636 & ~x644 & ~x659 & ~x721 & ~x745 & ~x748 & ~x783;
assign c7148 =  x677;
assign c7152 =  x238 &  x266 &  x295 &  x323 &  x491 &  x547 &  x659 & ~x55 & ~x244 & ~x271 & ~x452 & ~x532 & ~x597 & ~x598 & ~x625 & ~x774;
assign c7154 = ~x186 & ~x349 & ~x379 & ~x406 & ~x435 & ~x489 & ~x570 & ~x624 & ~x781;
assign c7156 =  x321 &  x340;
assign c7158 =  x597 &  x624 & ~x602 & ~x631;
assign c7160 =  x185 &  x574 &  x602 & ~x320 & ~x400 & ~x404 & ~x598;
assign c7162 =  x736;
assign c7164 =  x772;
assign c7166 =  x231 &  x520 &  x604;
assign c7168 =  x239 &  x240 &  x267 &  x295 &  x324 &  x462 & ~x72 & ~x347 & ~x371 & ~x564 & ~x571 & ~x627;
assign c7170 =  x316;
assign c7172 =  x231 & ~x153 & ~x625 & ~x654;
assign c7174 =  x676;
assign c7176 =  x205 &  x206 &  x238 &  x520 &  x548 & ~x151 & ~x190 & ~x215 & ~x681 & ~x731;
assign c7178 =  x367;
assign c7180 =  x269 &  x713 & ~x34 & ~x67 & ~x101 & ~x127 & ~x153 & ~x160 & ~x221 & ~x224 & ~x330 & ~x362 & ~x363 & ~x391 & ~x399 & ~x400 & ~x444 & ~x509 & ~x527 & ~x593 & ~x645 & ~x654 & ~x705 & ~x718 & ~x738 & ~x770 & ~x775;
assign c7182 =  x267 &  x293 & ~x152 & ~x160 & ~x183 & ~x211 & ~x255 & ~x624 & ~x763;
assign c7184 =  x328 &  x355 &  x383 & ~x434 & ~x488 & ~x623 & ~x624;
assign c7186 =  x704;
assign c7188 =  x570 &  x679;
assign c7190 =  x717;
assign c7192 =  x240 &  x464 &  x491 &  x575 &  x687 & ~x299 & ~x597 & ~x598 & ~x599;
assign c7194 =  x167;
assign c7196 =  x238 &  x240 &  x489 &  x516 &  x517 & ~x75 & ~x344 & ~x521 & ~x550 & ~x575 & ~x576 & ~x603 & ~x698;
assign c7198 =  x321 &  x322 & ~x142 & ~x151 & ~x178 & ~x183 & ~x209 & ~x624;
assign c7200 =  x259 &  x262 &  x266 &  x267 & ~x151 & ~x571;
assign c7202 =  x284;
assign c7204 =  x238 & ~x349 & ~x434 & ~x435 & ~x490;
assign c7206 =  x266 &  x632 &  x660 &  x688;
assign c7208 =  x573 &  x601 &  x628 &  x683 &  x711 & ~x406 & ~x532;
assign c7210 =  x208 &  x462 &  x489 &  x517 & ~x82 & ~x163 & ~x277 & ~x292 & ~x300 & ~x314 & ~x414 & ~x522 & ~x575 & ~x576 & ~x633;
assign c7212 =  x439 &  x440 & ~x183 & ~x571;
assign c7214 = ~x177 & ~x183 & ~x433 & ~x488 & ~x490 & ~x517 & ~x573 & ~x599 & ~x654;
assign c7216 =  x339;
assign c7218 =  x517 &  x544 &  x599 &  x600 &  x682 & ~x46 & ~x49 & ~x54 & ~x78 & ~x100 & ~x164 & ~x337 & ~x387 & ~x401 & ~x418 & ~x421 & ~x528 & ~x557 & ~x576 & ~x591 & ~x594 & ~x603 & ~x631 & ~x634 & ~x659 & ~x661 & ~x675 & ~x687 & ~x700 & ~x771 & ~x776;
assign c7220 = ~x183 & ~x435 & ~x488 & ~x491 & ~x573 & ~x629;
assign c7222 =  x244 &  x263 &  x267 &  x269 & ~x185;
assign c7226 =  x243 &  x271 &  x299 &  x327 &  x462 & ~x75 & ~x123 & ~x134 & ~x250 & ~x333 & ~x450 & ~x521 & ~x522 & ~x560 & ~x576 & ~x578 & ~x591 & ~x603 & ~x609 & ~x614 & ~x619 & ~x665 & ~x672 & ~x763;
assign c7228 =  x440 &  x441 & ~x571 & ~x596 & ~x599 & ~x622 & ~x653;
assign c7230 =  x42;
assign c7232 =  x630 &  x713 & ~x433 & ~x597;
assign c7234 =  x32;
assign c7236 =  x207 &  x489 & ~x59 & ~x153 & ~x190 & ~x320 & ~x397 & ~x522 & ~x525 & ~x554 & ~x576 & ~x634;
assign c7238 =  x300 & ~x184 & ~x185 & ~x191 & ~x575;
assign c7242 =  x207 &  x239 &  x240 &  x462 & ~x52 & ~x108 & ~x189 & ~x272 & ~x291 & ~x292 & ~x339 & ~x345 & ~x371 & ~x523 & ~x550 & ~x595 & ~x695;
assign c7244 =  x263 &  x266 &  x269 &  x271 &  x298 &  x382 & ~x331 & ~x396 & ~x477 & ~x740;
assign c7246 =  x238 &  x242 &  x297 &  x407 &  x462 & ~x157 & ~x221 & ~x277 & ~x342 & ~x371 & ~x551 & ~x575 & ~x576 & ~x664 & ~x687 & ~x770;
assign c7248 =  x207 &  x517 & ~x9 & ~x57 & ~x60 & ~x61 & ~x81 & ~x142 & ~x193 & ~x225 & ~x283 & ~x286 & ~x314 & ~x315 & ~x319 & ~x356 & ~x372 & ~x426 & ~x445 & ~x498 & ~x499 & ~x500 & ~x506 & ~x525 & ~x539 & ~x553 & ~x566 & ~x567 & ~x576 & ~x578 & ~x634 & ~x635 & ~x662 & ~x703 & ~x720;
assign c7250 =  x678;
assign c7252 =  x435 &  x517 &  x600 & ~x101 & ~x157 & ~x197 & ~x248 & ~x315 & ~x319 & ~x320 & ~x400 & ~x522 & ~x549 & ~x576 & ~x603 & ~x637 & ~x662 & ~x701 & ~x718 & ~x769;
assign c7254 =  x293 &  x294 & ~x183 & ~x210 & ~x211 & ~x212 & ~x238;
assign c7256 =  x10;
assign c7258 = ~x210 & ~x211 & ~x239 & ~x434;
assign c7260 =  x299 & ~x36 & ~x106 & ~x120 & ~x160 & ~x260 & ~x288 & ~x349 & ~x510 & ~x575 & ~x576 & ~x629 & ~x635 & ~x659 & ~x722;
assign c7262 =  x207 &  x208 &  x209 &  x267 &  x545 &  x600 & ~x576 & ~x634 & ~x662;
assign c7266 =  x256;
assign c7268 =  x464 &  x491 &  x519 &  x574 & ~x29 & ~x73 & ~x78 & ~x90 & ~x99 & ~x139 & ~x151 & ~x170 & ~x188 & ~x191 & ~x229 & ~x286 & ~x331 & ~x419 & ~x433 & ~x439 & ~x488 & ~x489 & ~x522 & ~x523 & ~x526 & ~x550 & ~x551 & ~x587 & ~x597 & ~x598 & ~x614 & ~x634 & ~x637 & ~x679 & ~x699 & ~x742 & ~x744 & ~x770 & ~x777;
assign c7270 =  x195;
assign c7272 =  x269 &  x464 &  x546 &  x574 & ~x75 & ~x156 & ~x186 & ~x345 & ~x374 & ~x423 & ~x597;
assign c7274 =  x227;
assign c7276 =  x463 &  x545 &  x573 &  x600 &  x627 &  x628 &  x683 & ~x37 & ~x58 & ~x76 & ~x78 & ~x79 & ~x88 & ~x101 & ~x106 & ~x114 & ~x120 & ~x123 & ~x137 & ~x189 & ~x219 & ~x225 & ~x277 & ~x281 & ~x341 & ~x365 & ~x367 & ~x423 & ~x426 & ~x450 & ~x498 & ~x525 & ~x556 & ~x603 & ~x604 & ~x606 & ~x620 & ~x641 & ~x659 & ~x689 & ~x692 & ~x725 & ~x728 & ~x730 & ~x735 & ~x742 & ~x743 & ~x774;
assign c7278 =  x167;
assign c7280 =  x235 &  x655 & ~x603;
assign c7282 =  x232 &  x233 &  x235 &  x236 &  x464 &  x519 &  x603 & ~x279 & ~x391;
assign c7284 =  x739;
assign c7286 =  x269 &  x352 &  x574 &  x630 &  x686 & ~x2 & ~x19 & ~x39 & ~x44 & ~x65 & ~x67 & ~x75 & ~x94 & ~x102 & ~x124 & ~x145 & ~x165 & ~x167 & ~x188 & ~x219 & ~x301 & ~x330 & ~x336 & ~x342 & ~x346 & ~x418 & ~x425 & ~x426 & ~x452 & ~x477 & ~x559 & ~x586 & ~x593 & ~x594 & ~x597 & ~x599 & ~x636 & ~x650 & ~x652 & ~x655 & ~x682 & ~x697 & ~x701 & ~x758 & ~x771;
assign c7288 =  x231 &  x260 &  x266 &  x267 & ~x181 & ~x223 & ~x564 & ~x667;
assign c7290 =  x624 &  x678;
assign c7292 =  x241 &  x574 & ~x96 & ~x166 & ~x188 & ~x385 & ~x403 & ~x432 & ~x433 & ~x459 & ~x559 & ~x570 & ~x571 & ~x635 & ~x642 & ~x682;
assign c7294 =  x77;
assign c7296 =  x312;
assign c7298 = ~x154 & ~x405 & ~x435 & ~x517 & ~x545 & ~x546 & ~x572 & ~x629;
assign c71 =  x349 &  x376 &  x377 &  x378 & ~x36 & ~x37 & ~x86 & ~x90 & ~x94 & ~x95 & ~x118 & ~x121 & ~x189 & ~x311 & ~x336 & ~x358 & ~x366 & ~x420 & ~x426 & ~x672 & ~x735 & ~x748 & ~x771;
assign c73 =  x541 &  x542 & ~x3 & ~x79 & ~x127 & ~x176 & ~x505 & ~x615 & ~x652 & ~x658 & ~x674 & ~x687 & ~x729 & ~x753;
assign c75 =  x158;
assign c77 =  x348 &  x376 &  x377 & ~x42 & ~x60 & ~x61 & ~x64 & ~x94 & ~x95 & ~x109 & ~x159 & ~x160 & ~x193 & ~x198 & ~x311 & ~x335 & ~x336 & ~x422 & ~x445 & ~x448 & ~x456 & ~x457 & ~x478 & ~x479 & ~x480 & ~x484 & ~x507 & ~x558 & ~x561 & ~x568 & ~x590 & ~x615 & ~x618 & ~x646 & ~x690 & ~x733 & ~x767;
assign c79 =  x345 &  x458 &  x460 & ~x124;
assign c711 =  x555;
assign c713 =  x376 &  x377 &  x404 &  x405 & ~x16 & ~x21 & ~x59 & ~x87 & ~x90 & ~x146 & ~x153 & ~x255 & ~x307 & ~x386 & ~x394 & ~x414 & ~x427 & ~x446 & ~x560 & ~x611 & ~x673 & ~x728 & ~x735 & ~x743 & ~x744 & ~x780;
assign c715 =  x428 &  x457 &  x486 &  x487 & ~x91 & ~x110 & ~x112 & ~x113 & ~x146 & ~x169 & ~x174 & ~x228 & ~x306 & ~x474 & ~x477 & ~x648 & ~x675 & ~x749;
assign c717 =  x488 & ~x232 & ~x245 & ~x324 & ~x748;
assign c719 = ~x39 & ~x74 & ~x83 & ~x114 & ~x176 & ~x206 & ~x353 & ~x369 & ~x381 & ~x391 & ~x409 & ~x437 & ~x465 & ~x714 & ~x741 & ~x745 & ~x755;
assign c721 = ~x232 & ~x236 & ~x263 & ~x289 & ~x382 & ~x466;
assign c723 =  x554;
assign c725 =  x607 & ~x37 & ~x446;
assign c727 = ~x208 & ~x325 & ~x437 & ~x465;
assign c729 =  x351 & ~x62 & ~x151 & ~x180 & ~x204 & ~x206 & ~x235 & ~x311 & ~x358 & ~x371 & ~x419 & ~x456 & ~x457 & ~x465 & ~x711 & ~x731 & ~x757;
assign c731 =  x526;
assign c733 =  x510;
assign c735 =  x455 &  x484 & ~x711 & ~x712;
assign c737 =  x157 & ~x252 & ~x336 & ~x703 & ~x712 & ~x747;
assign c739 =  x158;
assign c741 = ~x59 & ~x146 & ~x167 & ~x184 & ~x198 & ~x240 & ~x241 & ~x268 & ~x269 & ~x276 & ~x296 & ~x323 & ~x336 & ~x395 & ~x669;
assign c743 =  x211 &  x577 & ~x9 & ~x160 & ~x164 & ~x232 & ~x389 & ~x496 & ~x712 & ~x735 & ~x748;
assign c745 =  x400 &  x458 &  x459;
assign c747 =  x577 &  x605 & ~x197 & ~x259;
assign c749 =  x158;
assign c751 =  x581;
assign c753 =  x663 & ~x265;
assign c755 =  x553;
assign c757 =  x580 & ~x165 & ~x732;
assign c759 =  x347 &  x432;
assign c761 =  x401 &  x429 & ~x267 & ~x323;
assign c763 =  x404 &  x405 & ~x3 & ~x5 & ~x32 & ~x93 & ~x109 & ~x138 & ~x149 & ~x176 & ~x469 & ~x496 & ~x510 & ~x615 & ~x668 & ~x748;
assign c765 = ~x206 & ~x233 & ~x353 & ~x381 & ~x409 & ~x464 & ~x685;
assign c767 =  x372 &  x400 &  x486 & ~x7 & ~x322 & ~x443 & ~x651;
assign c769 =  x608;
assign c771 =  x374 &  x403 &  x405 & ~x39 & ~x457;
assign c773 =  x577 &  x629 & ~x164 & ~x306 & ~x422 & ~x503 & ~x713;
assign c775 =  x607 & ~x138 & ~x143 & ~x166 & ~x329;
assign c777 =  x577 &  x605 & ~x4 & ~x43 & ~x44 & ~x88 & ~x143 & ~x167 & ~x197 & ~x257 & ~x395 & ~x499 & ~x505 & ~x574 & ~x697 & ~x738 & ~x759 & ~x760 & ~x779 & ~x782;
assign c779 =  x402 &  x403 & ~x37 & ~x136 & ~x141 & ~x148 & ~x231 & ~x254 & ~x282 & ~x322 & ~x441 & ~x456 & ~x470 & ~x586 & ~x701 & ~x748;
assign c781 =  x351 &  x377 & ~x95 & ~x106 & ~x110 & ~x310 & ~x382 & ~x410 & ~x448 & ~x588 & ~x672 & ~x675 & ~x697 & ~x701;
assign c783 =  x291 &  x404 &  x405;
assign c785 =  x375 &  x403 & ~x232 & ~x466;
assign c787 =  x378 &  x576 & ~x14 & ~x24 & ~x99 & ~x116 & ~x124 & ~x133 & ~x172 & ~x281 & ~x283 & ~x314 & ~x394 & ~x440 & ~x480 & ~x489 & ~x702 & ~x723 & ~x746;
assign c789 =  x371 &  x460 & ~x59 & ~x85 & ~x86 & ~x106 & ~x143 & ~x145 & ~x148 & ~x420 & ~x443 & ~x587 & ~x588;
assign c791 =  x605 &  x606 & ~x329 & ~x492;
assign c793 =  x514 &  x542 & ~x95 & ~x186 & ~x509 & ~x656 & ~x658 & ~x687 & ~x737 & ~x779;
assign c795 =  x401 &  x429 &  x458 &  x487;
assign c797 =  x155 & ~x106 & ~x289;
assign c799 =  x378 & ~x77 & ~x152 & ~x263 & ~x410 & ~x711;
assign c7101 =  x378 & ~x53 & ~x177 & ~x182 & ~x264 & ~x385 & ~x388 & ~x466 & ~x741 & ~x767;
assign c7103 =  x540 &  x541 & ~x2 & ~x35 & ~x61 & ~x67 & ~x109 & ~x136 & ~x146 & ~x280 & ~x306 & ~x310 & ~x333 & ~x338 & ~x366 & ~x390 & ~x559 & ~x619 & ~x622 & ~x649 & ~x673 & ~x676 & ~x687 & ~x712 & ~x713 & ~x715 & ~x746 & ~x748 & ~x752 & ~x776;
assign c7105 =  x348 &  x350 & ~x21 & ~x37 & ~x58 & ~x78 & ~x92 & ~x94 & ~x106 & ~x133 & ~x138 & ~x166 & ~x196 & ~x222 & ~x254 & ~x306 & ~x332 & ~x333 & ~x421 & ~x430 & ~x431 & ~x446 & ~x448 & ~x453 & ~x481 & ~x482 & ~x483 & ~x617 & ~x642 & ~x665 & ~x703 & ~x740 & ~x763;
assign c7107 =  x290 &  x404 & ~x28 & ~x61 & ~x470 & ~x496 & ~x585;
assign c7109 =  x374 &  x402 &  x460 & ~x393 & ~x449;
assign c7111 =  x485 &  x513 &  x514;
assign c7113 = ~x38 & ~x50 & ~x67 & ~x69 & ~x108 & ~x114 & ~x136 & ~x151 & ~x152 & ~x153 & ~x208 & ~x226 & ~x338 & ~x357 & ~x381 & ~x382 & ~x396 & ~x409 & ~x410 & ~x451 & ~x465 & ~x479 & ~x501 & ~x533 & ~x636 & ~x658 & ~x694 & ~x705 & ~x743 & ~x761 & ~x777;
assign c7115 = ~x12 & ~x37 & ~x42 & ~x66 & ~x149 & ~x241 & ~x267 & ~x268 & ~x269 & ~x295 & ~x296 & ~x388 & ~x534 & ~x646 & ~x667 & ~x699 & ~x780 & ~x782;
assign c7117 =  x429 &  x487 & ~x67 & ~x71 & ~x220 & ~x256 & ~x259 & ~x432 & ~x444;
assign c7119 =  x405 &  x406 & ~x62 & ~x194 & ~x383 & ~x421 & ~x437 & ~x456 & ~x465;
assign c7121 =  x538 & ~x715;
assign c7123 =  x608 & ~x273;
assign c7125 =  x566;
assign c7127 =  x578 &  x605 & ~x20 & ~x61 & ~x114 & ~x279 & ~x281 & ~x364 & ~x531 & ~x687 & ~x758;
assign c7129 =  x606 &  x657;
assign c7131 =  x400 &  x460;
assign c7133 =  x595 & ~x7 & ~x45 & ~x101 & ~x501 & ~x588 & ~x589 & ~x591 & ~x679;
assign c7135 = ~x35 & ~x203 & ~x204 & ~x263 & ~x297 & ~x298 & ~x353 & ~x381 & ~x615;
assign c7137 =  x402 &  x431 & ~x204 & ~x323 & ~x756;
assign c7139 =  x513 & ~x267 & ~x675;
assign c7141 =  x430 &  x458 &  x460 & ~x204 & ~x279;
assign c7143 =  x456 &  x486 & ~x255 & ~x479;
assign c7145 =  x539;
assign c7147 =  x126;
assign c7149 =  x372 &  x432 & ~x55 & ~x203;
assign c7151 =  x399 &  x458;
assign c7153 =  x405 & ~x131 & ~x176 & ~x202 & ~x206 & ~x394 & ~x420 & ~x494 & ~x509 & ~x634 & ~x703;
assign c7155 =  x120;
assign c7157 =  x401 &  x458 &  x459 &  x460 & ~x311 & ~x558;
assign c7159 =  x378 & ~x383 & ~x437 & ~x465 & ~x685;
assign c7161 =  x317 &  x431 &  x432 & ~x202 & ~x440 & ~x496;
assign c7163 =  x184 &  x348 & ~x304 & ~x696 & ~x782;
assign c7165 =  x291 &  x405 & ~x12 & ~x30 & ~x41 & ~x58 & ~x81 & ~x136 & ~x158 & ~x160 & ~x232 & ~x260 & ~x281 & ~x310 & ~x334 & ~x340 & ~x442 & ~x469 & ~x579 & ~x661 & ~x662 & ~x664 & ~x666 & ~x722 & ~x744 & ~x772;
assign c7167 =  x577 & ~x9 & ~x360 & ~x464 & ~x483 & ~x615 & ~x736;
assign c7169 =  x155 & ~x142 & ~x445 & ~x561;
assign c7171 = ~x146 & ~x262 & ~x289 & ~x341 & ~x353 & ~x354 & ~x365 & ~x381 & ~x426 & ~x479 & ~x503 & ~x708;
assign c7173 =  x156 & ~x685;
assign c7175 = ~x36 & ~x61 & ~x268 & ~x269 & ~x270 & ~x297 & ~x325 & ~x352 & ~x395 & ~x627;
assign c7177 =  x577 & ~x21 & ~x30 & ~x35 & ~x37 & ~x146 & ~x194 & ~x232 & ~x311 & ~x384 & ~x393 & ~x423 & ~x558 & ~x639 & ~x641 & ~x642 & ~x664 & ~x712 & ~x773;
assign c7179 =  x401 &  x402 &  x434 & ~x443 & ~x480;
assign c7181 = ~x36 & ~x51 & ~x106 & ~x145 & ~x157 & ~x241 & ~x268 & ~x269 & ~x277 & ~x283 & ~x295 & ~x296 & ~x339 & ~x496 & ~x497 & ~x560 & ~x608 & ~x775;
assign c7183 = ~x115 & ~x241 & ~x269 & ~x289 & ~x297 & ~x368 & ~x381 & ~x383 & ~x410 & ~x428 & ~x698 & ~x763;
assign c7185 =  x569 &  x572 &  x598 & ~x584 & ~x712;
assign c7187 =  x159;
assign c7189 =  x405 &  x464 &  x520 & ~x21 & ~x93 & ~x94 & ~x174 & ~x175 & ~x202 & ~x258 & ~x280 & ~x281 & ~x283 & ~x306 & ~x385 & ~x424 & ~x457 & ~x468 & ~x496 & ~x622 & ~x674 & ~x780;
assign c7191 =  x426 & ~x202 & ~x295;
assign c7193 =  x378 & ~x236 & ~x263 & ~x382 & ~x466;
assign c7195 =  x349 &  x376 &  x377 & ~x138 & ~x252 & ~x304 & ~x330 & ~x355 & ~x392 & ~x417 & ~x421 & ~x424 & ~x456 & ~x470 & ~x503 & ~x513 & ~x517 & ~x529;
assign c7197 =  x153 &  x154 &  x576 & ~x1 & ~x46 & ~x106 & ~x364 & ~x447 & ~x507 & ~x641 & ~x670;
assign c7199 =  x184 &  x349 & ~x306;
assign c7201 =  x351 &  x378 & ~x311 & ~x412 & ~x457 & ~x466 & ~x686;
assign c7203 =  x350 &  x377 &  x378 & ~x6 & ~x46 & ~x53 & ~x91 & ~x94 & ~x95 & ~x113 & ~x117 & ~x122 & ~x136 & ~x151 & ~x357 & ~x385 & ~x411 & ~x419 & ~x427 & ~x456 & ~x470 & ~x476 & ~x483 & ~x484 & ~x509 & ~x538 & ~x582 & ~x640 & ~x641 & ~x728 & ~x751 & ~x776;
assign c7205 =  x401 &  x429 & ~x1 & ~x64 & ~x73 & ~x115 & ~x169 & ~x223 & ~x251 & ~x257 & ~x267 & ~x306 & ~x322 & ~x388 & ~x420 & ~x479 & ~x670 & ~x671 & ~x709 & ~x779;
assign c7207 = ~x83 & ~x171 & ~x223 & ~x242 & ~x267 & ~x269 & ~x297 & ~x338 & ~x539 & ~x646 & ~x673 & ~x677 & ~x757;
assign c7209 =  x404 & ~x438 & ~x466;
assign c7211 =  x606 &  x657;
assign c7213 =  x432 & ~x66 & ~x384 & ~x437;
assign c7215 =  x402 &  x431 & ~x43 & ~x148 & ~x169 & ~x322 & ~x440 & ~x470 & ~x592 & ~x620;
assign c7217 =  x551 & ~x4 & ~x17 & ~x35 & ~x65 & ~x82 & ~x131 & ~x142 & ~x227 & ~x229 & ~x252 & ~x257 & ~x308 & ~x335 & ~x336 & ~x366 & ~x641 & ~x687 & ~x708 & ~x714 & ~x740;
assign c7219 =  x405 & ~x466 & ~x711;
assign c7221 =  x455;
assign c7223 =  x401 &  x430 &  x458;
assign c7225 =  x511 & ~x176 & ~x558 & ~x687;
assign c7227 =  x159;
assign c7229 =  x539;
assign c7231 =  x372 &  x401 &  x403 & ~x470;
assign c7233 =  x377 &  x404 &  x405 & ~x202 & ~x322 & ~x336 & ~x390 & ~x586;
assign c7235 =  x576 & ~x34 & ~x55 & ~x101 & ~x115 & ~x147 & ~x192 & ~x232 & ~x233 & ~x249 & ~x307 & ~x309 & ~x333 & ~x421 & ~x466 & ~x508 & ~x560 & ~x697;
assign c7237 =  x578 & ~x17 & ~x32 & ~x42 & ~x57 & ~x116 & ~x149 & ~x171 & ~x225 & ~x254 & ~x281 & ~x310 & ~x337 & ~x369 & ~x504 & ~x547 & ~x745;
assign c7239 =  x595 & ~x250;
assign c7241 =  x485 &  x514 & ~x30 & ~x39 & ~x44 & ~x56 & ~x70 & ~x74 & ~x88 & ~x117 & ~x144 & ~x278 & ~x338 & ~x364 & ~x448 & ~x452 & ~x474 & ~x533 & ~x618 & ~x623 & ~x694 & ~x698 & ~x711 & ~x730 & ~x749 & ~x754 & ~x755 & ~x757 & ~x759 & ~x770 & ~x782;
assign c7243 =  x430 &  x432 & ~x470;
assign c7245 =  x405 &  x407 & ~x22 & ~x23 & ~x90 & ~x266 & ~x267 & ~x393 & ~x416 & ~x457 & ~x504 & ~x697 & ~x701 & ~x776;
assign c7247 =  x375 &  x404 &  x405 & ~x62 & ~x145 & ~x192 & ~x249 & ~x422 & ~x428 & ~x478 & ~x611 & ~x696 & ~x702 & ~x705;
assign c7249 =  x404 &  x405 & ~x296;
assign c7251 =  x348 &  x349 &  x350 & ~x3 & ~x5 & ~x9 & ~x37 & ~x44 & ~x58 & ~x91 & ~x99 & ~x106 & ~x109 & ~x128 & ~x146 & ~x149 & ~x171 & ~x199 & ~x201 & ~x228 & ~x229 & ~x250 & ~x254 & ~x255 & ~x256 & ~x257 & ~x280 & ~x304 & ~x333 & ~x362 & ~x369 & ~x370 & ~x387 & ~x394 & ~x418 & ~x419 & ~x428 & ~x445 & ~x451 & ~x457 & ~x473 & ~x498 & ~x504 & ~x530 & ~x611 & ~x613 & ~x617 & ~x691 & ~x718 & ~x724 & ~x729 & ~x734 & ~x735 & ~x755 & ~x757 & ~x760 & ~x764 & ~x770 & ~x777 & ~x780;
assign c7253 =  x607 & ~x42 & ~x329;
assign c7255 =  x598 & ~x15 & ~x16 & ~x28 & ~x30 & ~x44 & ~x62 & ~x64 & ~x66 & ~x81 & ~x86 & ~x98 & ~x102 & ~x111 & ~x113 & ~x136 & ~x159 & ~x168 & ~x171 & ~x172 & ~x222 & ~x229 & ~x250 & ~x258 & ~x275 & ~x281 & ~x282 & ~x302 & ~x336 & ~x342 & ~x394 & ~x395 & ~x502 & ~x527 & ~x530 & ~x533 & ~x554 & ~x555 & ~x556 & ~x558 & ~x561 & ~x608 & ~x615 & ~x620 & ~x640 & ~x684 & ~x685 & ~x699 & ~x713 & ~x715 & ~x721 & ~x723 & ~x760 & ~x764 & ~x766 & ~x769 & ~x776 & ~x779 & ~x780 & ~x782 & ~x783;
assign c7257 =  x125;
assign c7259 =  x376 &  x377 &  x378 & ~x22 & ~x35 & ~x39 & ~x101 & ~x198 & ~x283 & ~x305 & ~x311 & ~x312 & ~x388 & ~x394 & ~x418 & ~x423 & ~x454 & ~x460 & ~x461 & ~x568 & ~x586 & ~x642 & ~x750 & ~x755 & ~x780 & ~x782;
assign c7261 =  x495 &  x542 & ~x9 & ~x29 & ~x48 & ~x53 & ~x76 & ~x133 & ~x146 & ~x170 & ~x199 & ~x281 & ~x311 & ~x332 & ~x533 & ~x562 & ~x611 & ~x651 & ~x673 & ~x687 & ~x711 & ~x741 & ~x762;
assign c7263 =  x568 & ~x352 & ~x677 & ~x751;
assign c7265 =  x568 & ~x19 & ~x35 & ~x75 & ~x81 & ~x99 & ~x352 & ~x393 & ~x683 & ~x685 & ~x725 & ~x740 & ~x757;
assign c7267 =  x372 &  x400 &  x429 &  x433 & ~x176;
assign c7269 =  x374 &  x432 & ~x99 & ~x441;
assign c7271 =  x428 &  x458 &  x488;
assign c7273 =  x430 &  x459 & ~x33 & ~x37 & ~x42 & ~x65 & ~x72 & ~x125 & ~x140 & ~x141 & ~x174 & ~x176 & ~x203 & ~x303 & ~x322 & ~x337 & ~x368 & ~x395 & ~x451 & ~x468 & ~x483 & ~x496 & ~x587 & ~x635 & ~x672 & ~x724;
assign c7275 =  x374 &  x403 &  x432 & ~x440;
assign c7277 =  x400 &  x458;
assign c7279 =  x431 & ~x232 & ~x296 & ~x324;
assign c7281 =  x656 &  x657 & ~x0 & ~x15 & ~x17 & ~x42 & ~x86 & ~x121 & ~x195 & ~x253 & ~x254 & ~x255 & ~x279 & ~x305 & ~x338 & ~x340 & ~x368 & ~x396 & ~x464 & ~x474 & ~x477 & ~x531 & ~x556 & ~x558 & ~x611 & ~x672 & ~x694 & ~x697 & ~x711 & ~x714 & ~x735 & ~x745 & ~x768 & ~x782;
assign c7283 =  x399 &  x428 &  x460;
assign c7285 =  x483 &  x514;
assign c7287 =  x429 &  x458 &  x459 & ~x129 & ~x175 & ~x323 & ~x468 & ~x509 & ~x674 & ~x739 & ~x769 & ~x777 & ~x778;
assign c7289 =  x430 & ~x13 & ~x37 & ~x195 & ~x232 & ~x322 & ~x335 & ~x438 & ~x466 & ~x556;
assign c7291 =  x467 &  x496 &  x524 & ~x10 & ~x78 & ~x90 & ~x162 & ~x223 & ~x304 & ~x358 & ~x452 & ~x476 & ~x643;
assign c7293 =  x514 & ~x353;
assign c7297 =  x377 &  x378 &  x380 & ~x16 & ~x113 & ~x149 & ~x166 & ~x222 & ~x249 & ~x281 & ~x383 & ~x385 & ~x411 & ~x421 & ~x440 & ~x470 & ~x513 & ~x766 & ~x776;
assign c7299 =  x405 & ~x437 & ~x628;
assign c80 =  x179 &  x288 &  x317 &  x347 &  x376 & ~x188 & ~x311 & ~x562 & ~x681;
assign c82 =  x404 &  x485 &  x540 & ~x148 & ~x175 & ~x223 & ~x331 & ~x384 & ~x515 & ~x545 & ~x556 & ~x637 & ~x644 & ~x649 & ~x676 & ~x741;
assign c84 =  x406 &  x432 &  x459 &  x486 &  x513 &  x655 & ~x203 & ~x389;
assign c86 =  x502;
assign c88 =  x380 &  x459 &  x513 &  x541 &  x656 & ~x544 & ~x743;
assign c810 =  x502;
assign c812 =  x513 &  x569 &  x656 & ~x131 & ~x572;
assign c814 =  x156 &  x349 &  x485 & ~x543;
assign c816 =  x325 &  x376 &  x457 &  x540 & ~x444 & ~x583 & ~x611;
assign c818 =  x460 &  x515 &  x657 & ~x266;
assign c820 =  x460 &  x515 &  x657 & ~x573;
assign c822 =  x487 &  x595 & ~x208 & ~x429;
assign c824 =  x187 &  x265 &  x293 & ~x400 & ~x521;
assign c826 =  x572 &  x600 &  x659 & ~x45 & ~x52 & ~x54 & ~x63 & ~x104 & ~x172 & ~x176 & ~x198 & ~x278 & ~x391 & ~x439 & ~x497 & ~x511 & ~x557 & ~x569 & ~x583 & ~x584 & ~x592 & ~x596 & ~x597 & ~x639 & ~x673 & ~x681 & ~x724 & ~x745;
assign c828 =  x327 &  x488 & ~x123 & ~x228 & ~x296 & ~x411 & ~x553 & ~x564 & ~x583;
assign c830 =  x567 & ~x296 & ~x520;
assign c832 =  x311;
assign c834 =  x574 &  x662;
assign c836 =  x290 &  x376 &  x488 & ~x401;
assign c838 =  x544 &  x600 & ~x195 & ~x200 & ~x390 & ~x470 & ~x513 & ~x574 & ~x598 & ~x626 & ~x677 & ~x690;
assign c840 =  x489 &  x544 &  x687;
assign c842 =  x290 &  x348 &  x377 & ~x84 & ~x225 & ~x373 & ~x400 & ~x667;
assign c844 =  x316 &  x545 &  x660;
assign c846 =  x16;
assign c848 =  x352 &  x380 &  x404 &  x511 &  x539 & ~x35 & ~x225 & ~x453 & ~x665;
assign c850 =  x13;
assign c852 =  x332;
assign c854 =  x461 &  x569 &  x657 & ~x106 & ~x205 & ~x341 & ~x678 & ~x780;
assign c856 =  x377 &  x379 &  x380 &  x458 &  x485 &  x539 &  x625;
assign c858 =  x318 &  x376 &  x461 & ~x400 & ~x625;
assign c860 =  x732;
assign c862 =  x286 &  x372;
assign c864 =  x152 &  x286 &  x373;
assign c866 =  x153 &  x292 &  x321 &  x379;
assign c868 =  x325 &  x350 &  x457 &  x597;
assign c870 =  x24;
assign c872 =  x514 &  x542 &  x570 & ~x6 & ~x69 & ~x159 & ~x161 & ~x191 & ~x309 & ~x389 & ~x483 & ~x511 & ~x567 & ~x573 & ~x678 & ~x703 & ~x713 & ~x774;
assign c874 =  x289 &  x318 &  x376 & ~x0 & ~x21 & ~x44 & ~x71 & ~x120 & ~x134 & ~x252 & ~x285 & ~x303 & ~x312 & ~x369 & ~x400 & ~x420 & ~x443 & ~x510 & ~x511 & ~x537 & ~x673;
assign c876 =  x318 &  x488 &  x516 & ~x18 & ~x66 & ~x126 & ~x136 & ~x226 & ~x420 & ~x440 & ~x456 & ~x474 & ~x480 & ~x509 & ~x510 & ~x511 & ~x525 & ~x529 & ~x588 & ~x590 & ~x638 & ~x731 & ~x743 & ~x744 & ~x751 & ~x754 & ~x769 & ~x770;
assign c878 =  x110;
assign c880 =  x263 &  x517 &  x658 & ~x225 & ~x284 & ~x384 & ~x456 & ~x511 & ~x540 & ~x596 & ~x680 & ~x704;
assign c882 =  x265 &  x515 &  x569 &  x654 & ~x742;
assign c884 =  x516 &  x544 &  x633 &  x660 & ~x597;
assign c886 =  x154 &  x348 &  x485;
assign c888 =  x87;
assign c890 =  x403 &  x540 &  x656 & ~x572;
assign c892 =  x488 &  x543 &  x657 & ~x400;
assign c894 =  x461 &  x488 &  x515 &  x542 &  x574 & ~x549;
assign c896 =  x234 &  x462 &  x660 & ~x626;
assign c898 =  x477;
assign c8100 =  x357 & ~x494 & ~x497;
assign c8102 =  x302 &  x458 & ~x385;
assign c8104 =  x154 &  x292 & ~x238 & ~x553;
assign c8106 =  x20;
assign c8108 =  x478;
assign c8110 =  x328 &  x460 & ~x352 & ~x494 & ~x521;
assign c8112 =  x292 &  x460 &  x487 & ~x288 & ~x447 & ~x456 & ~x494 & ~x521;
assign c8114 =  x165;
assign c8116 =  x514 &  x542 & ~x80 & ~x516 & ~x573 & ~x600;
assign c8118 =  x20;
assign c8120 =  x405 &  x432 &  x567 & ~x52 & ~x414 & ~x529 & ~x571 & ~x649;
assign c8122 =  x153 &  x154 &  x377 & ~x574 & ~x596 & ~x653 & ~x748;
assign c8124 =  x26;
assign c8126 =  x767;
assign c8128 =  x206 &  x299 &  x343 &  x432;
assign c8130 =  x317 &  x345 &  x461 &  x516 & ~x0 & ~x56 & ~x91 & ~x133 & ~x162 & ~x218 & ~x224 & ~x249 & ~x282 & ~x390 & ~x442 & ~x525 & ~x567 & ~x568 & ~x728;
assign c8132 =  x720;
assign c8134 =  x376 &  x379 &  x457 &  x484 & ~x547;
assign c8136 =  x474;
assign c8138 =  x168;
assign c8140 =  x783;
assign c8142 =  x331;
assign c8144 =  x405 &  x458 &  x539 & ~x542;
assign c8146 =  x153 & ~x128 & ~x175 & ~x209 & ~x479 & ~x547;
assign c8148 =  x331 &  x384;
assign c8150 =  x663 & ~x598;
assign c8152 =  x334;
assign c8154 =  x153 &  x233 &  x261 &  x376;
assign c8156 =  x207 &  x234 &  x261 &  x659;
assign c8158 =  x159 &  x488;
assign c8160 =  x699;
assign c8162 =  x515 &  x543 &  x571 &  x686 & ~x485 & ~x573;
assign c8164 =  x110;
assign c8166 =  x356 & ~x326 & ~x467 & ~x521 & ~x526;
assign c8168 =  x487 &  x514 &  x542 &  x656 & ~x149 & ~x572;
assign c8170 =  x690;
assign c8172 =  x290 &  x517 &  x544 &  x545 & ~x140 & ~x596;
assign c8174 =  x384 &  x595 & ~x520;
assign c8176 =  x359 &  x384;
assign c8178 =  x516 &  x659 & ~x602;
assign c8180 =  x245 &  x349 & ~x374 & ~x521;
assign c8182 =  x574 &  x634 & ~x311 & ~x597 & ~x625;
assign c8184 =  x276;
assign c8186 =  x61;
assign c8188 =  x233 &  x320 & ~x315;
assign c8190 =  x58;
assign c8192 =  x334;
assign c8194 =  x350 &  x485 &  x512 & ~x108 & ~x175 & ~x230 & ~x282 & ~x514 & ~x527 & ~x583;
assign c8196 =  x393;
assign c8198 =  x544 &  x658 & ~x33 & ~x51 & ~x146 & ~x176 & ~x218 & ~x511 & ~x513 & ~x530 & ~x574 & ~x582 & ~x781;
assign c8200 =  x404 &  x601 &  x633 &  x660 & ~x13 & ~x202 & ~x339 & ~x619 & ~x626 & ~x701;
assign c8202 =  x205 &  x286 & ~x262;
assign c8204 =  x315 &  x461 &  x607;
assign c8206 =  x316 &  x517 &  x660;
assign c8208 =  x186 & ~x152 & ~x189 & ~x200 & ~x268 & ~x296 & ~x363 & ~x401 & ~x427 & ~x467;
assign c8210 =  x515 &  x547 &  x598 & ~x107 & ~x440 & ~x540;
assign c8212 =  x236 &  x515 &  x570 &  x598 & ~x232;
assign c8214 =  x343 &  x634;
assign c8216 =  x261 &  x347 &  x375 &  x376 & ~x220 & ~x372;
assign c8218 =  x372 &  x517 &  x634;
assign c8220 =  x544 &  x686 & ~x202 & ~x567;
assign c8222 =  x459 &  x514 &  x657 & ~x500 & ~x573;
assign c8224 =  x515 &  x654 & ~x296;
assign c8226 =  x515 &  x543 &  x657 & ~x23 & ~x384 & ~x545 & ~x676 & ~x679;
assign c8228 =  x403 &  x569 & ~x93 & ~x102 & ~x188 & ~x399 & ~x443;
assign c8230 =  x65;
assign c8232 =  x405 &  x515 &  x658;
assign c8234 =  x544 &  x659 & ~x574 & ~x597;
assign c8236 =  x460 &  x515 &  x542 &  x570 & ~x572;
assign c8238 =  x459 &  x486 &  x540 &  x653;
assign c8240 =  x116;
assign c8242 =  x335;
assign c8244 =  x196 &  x727;
assign c8246 =  x237 &  x488 &  x543 &  x570 &  x656;
assign c8248 =  x312;
assign c8252 =  x290 &  x319 &  x348 &  x349 & ~x482 & ~x563 & ~x680 & ~x681 & ~x711 & ~x741 & ~x776;
assign c8254 =  x290 &  x348 & ~x238;
assign c8256 =  x299 &  x655 & ~x206 & ~x572;
assign c8258 =  x186 &  x320 &  x488 & ~x466 & ~x578 & ~x733;
assign c8260 =  x254;
assign c8262 =  x301 &  x328 &  x460 & ~x411 & ~x468 & ~x620;
assign c8264 =  x404 &  x405 &  x544 &  x631 & ~x43 & ~x201 & ~x513 & ~x567;
assign c8266 =  x186 &  x461 & ~x207 & ~x402;
assign c8268 =  x574 &  x634 & ~x599;
assign c8270 =  x331;
assign c8272 =  x265 &  x461 &  x514 &  x568;
assign c8274 =  x236 &  x542 & ~x100 & ~x205 & ~x226 & ~x467 & ~x537 & ~x552 & ~x582 & ~x587;
assign c8276 =  x459 &  x541 & ~x41 & ~x51 & ~x86 & ~x104 & ~x145 & ~x174 & ~x247 & ~x259 & ~x411 & ~x413 & ~x428 & ~x456 & ~x482 & ~x533 & ~x590 & ~x607 & ~x612 & ~x678 & ~x708 & ~x712 & ~x714 & ~x716 & ~x717 & ~x752;
assign c8278 =  x302 &  x460 & ~x152;
assign c8280 =  x421;
assign c8282 =  x154 &  x288 &  x345 &  x404 & ~x190 & ~x264;
assign c8284 =  x278;
assign c8286 =  x376 &  x378 &  x485 & ~x573;
assign c8288 =  x516 & ~x149 & ~x178 & ~x428 & ~x563 & ~x573;
assign c8290 =  x383 & ~x271 & ~x296 & ~x426;
assign c8292 =  x302 & ~x296;
assign c8294 =  x378 &  x458 &  x624 & ~x44 & ~x195 & ~x307 & ~x400 & ~x515;
assign c8296 =  x291 &  x320 &  x348 &  x406 & ~x26 & ~x116 & ~x120 & ~x201 & ~x226 & ~x288 & ~x413 & ~x690;
assign c8298 =  x153 &  x154 &  x292 &  x321 & ~x239;
assign c81 = ~x8 & ~x40 & ~x51 & ~x93 & ~x169 & ~x223 & ~x246 & ~x273 & ~x302 & ~x309 & ~x331 & ~x341 & ~x477 & ~x603 & ~x616 & ~x629 & ~x630 & ~x631 & ~x657 & ~x658 & ~x659 & ~x665 & ~x669 & ~x698 & ~x711 & ~x751 & ~x753;
assign c83 =  x346 &  x374 &  x601 & ~x1 & ~x35 & ~x44 & ~x260 & ~x306 & ~x460 & ~x461 & ~x639 & ~x729 & ~x734 & ~x749 & ~x779;
assign c85 =  x427 &  x428 & ~x154 & ~x420;
assign c87 =  x239 &  x266 &  x267 &  x629 & ~x270 & ~x326;
assign c89 = ~x6 & ~x248 & ~x316 & ~x474 & ~x615 & ~x628 & ~x629 & ~x630 & ~x631 & ~x656 & ~x657 & ~x658 & ~x666 & ~x710 & ~x719;
assign c811 =  x148;
assign c813 = ~x235 & ~x244 & ~x248 & ~x260 & ~x291 & ~x302 & ~x317 & ~x319 & ~x345 & ~x354 & ~x450 & ~x455;
assign c815 =  x181 &  x208 &  x209 &  x575 &  x576 &  x577 &  x601 &  x604 &  x629 &  x630 & ~x91 & ~x316 & ~x391 & ~x392;
assign c817 =  x401 &  x429 &  x430 & ~x28 & ~x33 & ~x34 & ~x47 & ~x64 & ~x83 & ~x117 & ~x125 & ~x217 & ~x246 & ~x273 & ~x274 & ~x275 & ~x285 & ~x294 & ~x309 & ~x329 & ~x361 & ~x418 & ~x420 & ~x449 & ~x472 & ~x555 & ~x558 & ~x614 & ~x636 & ~x644 & ~x649 & ~x669 & ~x675 & ~x680 & ~x690 & ~x707 & ~x720 & ~x724 & ~x727 & ~x728 & ~x731 & ~x747 & ~x750 & ~x762 & ~x766;
assign c819 =  x408 &  x437 &  x438 &  x465 &  x492 & ~x7 & ~x8 & ~x9 & ~x35 & ~x37 & ~x39 & ~x41 & ~x63 & ~x79 & ~x80 & ~x86 & ~x89 & ~x122 & ~x144 & ~x147 & ~x153 & ~x154 & ~x198 & ~x220 & ~x223 & ~x250 & ~x251 & ~x304 & ~x338 & ~x389 & ~x392 & ~x416 & ~x417 & ~x420 & ~x504 & ~x526 & ~x530 & ~x560 & ~x587 & ~x638 & ~x673 & ~x694 & ~x707 & ~x744 & ~x752;
assign c821 =  x267 &  x294 &  x295 & ~x130 & ~x185 & ~x215 & ~x371;
assign c823 =  x298 &  x354 &  x381 &  x437 & ~x1 & ~x75 & ~x81 & ~x156 & ~x221 & ~x254 & ~x338 & ~x394 & ~x500 & ~x587 & ~x595 & ~x638 & ~x690 & ~x780;
assign c825 = ~x1 & ~x72 & ~x217 & ~x230 & ~x235 & ~x236 & ~x244 & ~x263 & ~x299 & ~x326;
assign c827 =  x679 & ~x486;
assign c829 = ~x35 & ~x47 & ~x193 & ~x249 & ~x378 & ~x402 & ~x403 & ~x404 & ~x405 & ~x428 & ~x479 & ~x500 & ~x696 & ~x731 & ~x762;
assign c831 = ~x158 & ~x165 & ~x185 & ~x186 & ~x187 & ~x215 & ~x216 & ~x477 & ~x628 & ~x629 & ~x656 & ~x657 & ~x669 & ~x753;
assign c833 =  x436 & ~x25 & ~x28 & ~x51 & ~x71 & ~x92 & ~x105 & ~x126 & ~x130 & ~x137 & ~x143 & ~x154 & ~x155 & ~x156 & ~x157 & ~x161 & ~x273 & ~x276 & ~x280 & ~x287 & ~x313 & ~x385 & ~x450 & ~x563 & ~x568 & ~x615 & ~x621 & ~x626 & ~x669 & ~x694 & ~x727;
assign c835 = ~x156 & ~x184 & ~x601 & ~x628 & ~x657 & ~x753;
assign c837 = ~x0 & ~x6 & ~x48 & ~x267 & ~x280 & ~x294 & ~x319 & ~x321 & ~x345 & ~x348 & ~x349 & ~x376 & ~x689 & ~x690 & ~x722 & ~x753;
assign c839 =  x544 &  x599 & ~x302 & ~x306 & ~x472 & ~x475 & ~x535 & ~x576 & ~x595 & ~x603 & ~x611 & ~x630 & ~x631 & ~x649 & ~x658 & ~x674 & ~x715;
assign c841 =  x466 &  x467 &  x494 &  x495 &  x522 &  x550 & ~x68 & ~x78 & ~x95 & ~x134 & ~x333 & ~x475 & ~x490 & ~x560 & ~x640 & ~x669 & ~x751 & ~x753 & ~x774;
assign c843 =  x182 &  x185 &  x209 &  x211 &  x212 &  x606 & ~x25 & ~x316 & ~x502;
assign c845 =  x549 &  x576 &  x577 &  x603 &  x604 &  x605 & ~x43 & ~x53 & ~x64 & ~x119 & ~x143 & ~x251 & ~x286 & ~x302 & ~x304 & ~x329 & ~x330 & ~x361 & ~x516 & ~x586 & ~x610 & ~x669 & ~x709 & ~x711 & ~x777;
assign c847 =  x182 &  x209 & ~x29 & ~x41 & ~x48 & ~x63 & ~x66 & ~x142 & ~x171 & ~x196 & ~x241 & ~x242 & ~x243 & ~x244 & ~x245 & ~x271 & ~x272 & ~x273 & ~x277 & ~x280 & ~x285 & ~x301 & ~x327 & ~x328 & ~x330 & ~x339 & ~x357 & ~x359 & ~x501 & ~x502 & ~x563 & ~x585 & ~x586 & ~x640 & ~x669 & ~x693 & ~x719 & ~x731 & ~x778;
assign c849 =  x353 &  x381 & ~x5 & ~x15 & ~x80 & ~x81 & ~x82 & ~x84 & ~x140 & ~x172 & ~x194 & ~x230 & ~x249 & ~x278 & ~x280 & ~x302 & ~x338 & ~x361 & ~x388 & ~x416 & ~x420 & ~x447 & ~x477 & ~x503 & ~x506 & ~x560 & ~x612 & ~x628 & ~x655 & ~x656 & ~x670 & ~x680 & ~x711 & ~x751 & ~x753 & ~x756 & ~x760 & ~x762;
assign c851 =  x413 &  x441 &  x469 & ~x3 & ~x41 & ~x85 & ~x115 & ~x141 & ~x197 & ~x227 & ~x277 & ~x283 & ~x366 & ~x476 & ~x555 & ~x560 & ~x611 & ~x617 & ~x641 & ~x645 & ~x691 & ~x727 & ~x759 & ~x763 & ~x779;
assign c853 =  x603 &  x629 &  x630 & ~x298 & ~x300 & ~x326 & ~x354 & ~x364 & ~x530;
assign c855 =  x437 & ~x17 & ~x48 & ~x199 & ~x273 & ~x274 & ~x328 & ~x329 & ~x331 & ~x359 & ~x476 & ~x487 & ~x499 & ~x517 & ~x650 & ~x669 & ~x705 & ~x716 & ~x753 & ~x762;
assign c857 =  x440 &  x468 &  x495 &  x496 &  x523 & ~x246 & ~x311;
assign c859 = ~x406 & ~x430 & ~x432 & ~x433;
assign c861 = ~x112 & ~x366 & ~x431 & ~x432 & ~x433 & ~x455 & ~x459 & ~x460 & ~x461 & ~x517 & ~x586 & ~x613 & ~x617 & ~x644 & ~x749 & ~x753;
assign c863 = ~x13 & ~x26 & ~x29 & ~x35 & ~x41 & ~x63 & ~x64 & ~x78 & ~x92 & ~x97 & ~x105 & ~x121 & ~x195 & ~x198 & ~x251 & ~x253 & ~x322 & ~x323 & ~x349 & ~x350 & ~x376 & ~x377 & ~x378 & ~x395 & ~x404 & ~x417 & ~x420 & ~x445 & ~x502 & ~x503 & ~x535 & ~x585 & ~x620 & ~x640 & ~x690 & ~x696 & ~x722 & ~x723 & ~x731 & ~x770 & ~x774;
assign c865 =  x436 &  x519 & ~x6 & ~x16 & ~x24 & ~x40 & ~x73 & ~x86 & ~x91 & ~x92 & ~x100 & ~x105 & ~x118 & ~x124 & ~x129 & ~x148 & ~x156 & ~x157 & ~x167 & ~x203 & ~x230 & ~x231 & ~x286 & ~x302 & ~x341 & ~x360 & ~x361 & ~x364 & ~x417 & ~x448 & ~x474 & ~x512 & ~x513 & ~x558 & ~x563 & ~x577 & ~x582 & ~x587 & ~x605 & ~x639 & ~x676 & ~x690 & ~x695 & ~x702 & ~x722 & ~x727 & ~x753 & ~x777 & ~x778;
assign c867 = ~x24 & ~x34 & ~x48 & ~x105 & ~x111 & ~x119 & ~x369 & ~x502 & ~x626 & ~x628 & ~x629 & ~x630 & ~x631 & ~x656 & ~x657 & ~x658 & ~x659 & ~x666 & ~x669;
assign c869 = ~x41 & ~x380 & ~x381 & ~x408 & ~x435 & ~x463 & ~x464;
assign c871 = ~x70 & ~x321 & ~x348 & ~x375 & ~x656 & ~x657 & ~x658;
assign c873 =  x269 &  x296 &  x297 & ~x66 & ~x76 & ~x110 & ~x220 & ~x223 & ~x291 & ~x294 & ~x319 & ~x320 & ~x321 & ~x341 & ~x345 & ~x454 & ~x669 & ~x775;
assign c875 = ~x103 & ~x109 & ~x251 & ~x335 & ~x336 & ~x378 & ~x379 & ~x380 & ~x391 & ~x408 & ~x410 & ~x508 & ~x535 & ~x560 & ~x561 & ~x587 & ~x705 & ~x764 & ~x768;
assign c877 = ~x154 & ~x182 & ~x183 & ~x628 & ~x656 & ~x711;
assign c879 = ~x3 & ~x28 & ~x58 & ~x69 & ~x91 & ~x96 & ~x109 & ~x138 & ~x142 & ~x227 & ~x251 & ~x302 & ~x330 & ~x367 & ~x446 & ~x455 & ~x459 & ~x460 & ~x461 & ~x462 & ~x486 & ~x490 & ~x499 & ~x530 & ~x531 & ~x620 & ~x692 & ~x705 & ~x709 & ~x719 & ~x737 & ~x746 & ~x752 & ~x753 & ~x757 & ~x773;
assign c881 =  x576 &  x577 &  x578 &  x579 &  x603 &  x604 & ~x33 & ~x88 & ~x105 & ~x115 & ~x199 & ~x312 & ~x418 & ~x493 & ~x503 & ~x615 & ~x731 & ~x766;
assign c883 = ~x3 & ~x41 & ~x81 & ~x83 & ~x111 & ~x329 & ~x333 & ~x336 & ~x340 & ~x350 & ~x352 & ~x353 & ~x354 & ~x355 & ~x358 & ~x359 & ~x380 & ~x381 & ~x382 & ~x445 & ~x474 & ~x587 & ~x640 & ~x669 & ~x671 & ~x716;
assign c885 =  x466 &  x522 & ~x73 & ~x379;
assign c887 =  x98;
assign c889 =  x127 & ~x295 & ~x657 & ~x658;
assign c891 = ~x12 & ~x431 & ~x432 & ~x433 & ~x434 & ~x455 & ~x459 & ~x460 & ~x752;
assign c893 =  x426;
assign c895 = ~x8 & ~x24 & ~x49 & ~x56 & ~x64 & ~x70 & ~x78 & ~x88 & ~x92 & ~x101 & ~x104 & ~x107 & ~x119 & ~x145 & ~x166 & ~x170 & ~x249 & ~x332 & ~x333 & ~x349 & ~x359 & ~x375 & ~x376 & ~x393 & ~x402 & ~x404 & ~x431 & ~x503 & ~x561 & ~x613 & ~x670 & ~x695 & ~x696 & ~x712 & ~x726 & ~x753 & ~x762 & ~x773;
assign c897 =  x209 &  x629 & ~x24 & ~x34 & ~x83 & ~x96 & ~x459 & ~x460 & ~x461 & ~x735 & ~x761 & ~x778;
assign c899 =  x381 &  x437 &  x491 & ~x29 & ~x44 & ~x46 & ~x93 & ~x151 & ~x157 & ~x179 & ~x416 & ~x424 & ~x447 & ~x500 & ~x509 & ~x527 & ~x592 & ~x596 & ~x615 & ~x663 & ~x719 & ~x749;
assign c8101 =  x150 & ~x251 & ~x264 & ~x291 & ~x319 & ~x345 & ~x719 & ~x724 & ~x738;
assign c8103 =  x125 & ~x658;
assign c8105 =  x455 & ~x309 & ~x322;
assign c8107 =  x239 &  x267 &  x294 &  x295 & ~x244 & ~x382 & ~x688 & ~x769;
assign c8109 = ~x16 & ~x147 & ~x154 & ~x155 & ~x569 & ~x594 & ~x603 & ~x633 & ~x638 & ~x659 & ~x662 & ~x702 & ~x726 & ~x767;
assign c8111 =  x296 &  x297 &  x713 & ~x155 & ~x156;
assign c8113 =  x203 & ~x291;
assign c8115 =  x294 & ~x235 & ~x242 & ~x354;
assign c8117 = ~x4 & ~x42 & ~x50 & ~x58 & ~x99 & ~x123 & ~x125 & ~x128 & ~x139 & ~x154 & ~x155 & ~x156 & ~x157 & ~x158 & ~x182 & ~x183 & ~x184 & ~x185 & ~x186 & ~x251 & ~x257 & ~x330 & ~x361 & ~x396 & ~x414 & ~x504 & ~x528 & ~x585 & ~x586 & ~x649 & ~x669 & ~x719 & ~x731 & ~x765;
assign c8119 =  x437 &  x438 &  x465 &  x466 &  x492 &  x493 &  x520 &  x521 & ~x2 & ~x9 & ~x66 & ~x74 & ~x82 & ~x106 & ~x109 & ~x112 & ~x126 & ~x137 & ~x138 & ~x141 & ~x143 & ~x177 & ~x199 & ~x228 & ~x250 & ~x255 & ~x280 & ~x304 & ~x307 & ~x335 & ~x367 & ~x390 & ~x418 & ~x446 & ~x449 & ~x477 & ~x559 & ~x581 & ~x615 & ~x620 & ~x639 & ~x640 & ~x669 & ~x671 & ~x700 & ~x728 & ~x739 & ~x749 & ~x750 & ~x753 & ~x767 & ~x780;
assign c8121 = ~x366 & ~x378 & ~x379 & ~x406 & ~x433 & ~x449 & ~x563 & ~x641 & ~x720;
assign c8123 = ~x47 & ~x155 & ~x156 & ~x460 & ~x631;
assign c8125 =  x491 & ~x9 & ~x47 & ~x206 & ~x366 & ~x378 & ~x446 & ~x659 & ~x690 & ~x751 & ~x753 & ~x769 & ~x773;
assign c8127 = ~x12 & ~x28 & ~x220 & ~x295 & ~x321 & ~x348 & ~x349 & ~x350 & ~x375 & ~x376 & ~x377 & ~x447 & ~x534 & ~x559 & ~x687 & ~x690 & ~x692 & ~x698 & ~x757;
assign c8129 = ~x0 & ~x6 & ~x17 & ~x22 & ~x33 & ~x34 & ~x35 & ~x48 & ~x60 & ~x70 & ~x82 & ~x100 & ~x118 & ~x119 & ~x165 & ~x222 & ~x223 & ~x248 & ~x273 & ~x274 & ~x276 & ~x300 & ~x302 & ~x304 & ~x331 & ~x332 & ~x338 & ~x359 & ~x361 & ~x388 & ~x389 & ~x390 & ~x445 & ~x461 & ~x462 & ~x463 & ~x477 & ~x487 & ~x488 & ~x502 & ~x503 & ~x533 & ~x613 & ~x643 & ~x647 & ~x669 & ~x695 & ~x698 & ~x718 & ~x739;
assign c8131 =  x439 &  x466 &  x494 &  x521 & ~x6 & ~x27 & ~x33 & ~x54 & ~x85 & ~x93 & ~x109 & ~x126 & ~x139 & ~x152 & ~x163 & ~x169 & ~x171 & ~x173 & ~x228 & ~x248 & ~x251 & ~x253 & ~x283 & ~x304 & ~x332 & ~x341 & ~x360 & ~x396 & ~x418 & ~x422 & ~x474 & ~x476 & ~x477 & ~x526 & ~x532 & ~x554 & ~x641 & ~x669 & ~x675 & ~x692 & ~x705 & ~x730 & ~x731 & ~x745 & ~x749 & ~x762;
assign c8133 =  x267 & ~x244 & ~x260 & ~x262 & ~x354 & ~x577;
assign c8135 =  x408 &  x437 & ~x18 & ~x20 & ~x29 & ~x41 & ~x48 & ~x90 & ~x98 & ~x110 & ~x119 & ~x126 & ~x138 & ~x140 & ~x171 & ~x199 & ~x275 & ~x300 & ~x301 & ~x304 & ~x328 & ~x331 & ~x356 & ~x359 & ~x487 & ~x490 & ~x505 & ~x507 & ~x541 & ~x639 & ~x640 & ~x696 & ~x705 & ~x707 & ~x733 & ~x736;
assign c8137 =  x269 &  x297 & ~x21 & ~x22 & ~x36 & ~x41 & ~x42 & ~x73 & ~x77 & ~x85 & ~x90 & ~x100 & ~x105 & ~x137 & ~x171 & ~x195 & ~x218 & ~x219 & ~x250 & ~x283 & ~x293 & ~x294 & ~x302 & ~x304 & ~x312 & ~x318 & ~x319 & ~x321 & ~x332 & ~x334 & ~x336 & ~x338 & ~x388 & ~x400 & ~x417 & ~x424 & ~x479 & ~x613 & ~x615 & ~x617 & ~x620 & ~x675 & ~x693 & ~x706 & ~x737 & ~x778 & ~x782;
assign c8139 =  x436 &  x437 &  x465 &  x492 & ~x34 & ~x41 & ~x92 & ~x136 & ~x152 & ~x308 & ~x363 & ~x450 & ~x630 & ~x657;
assign c8141 =  x123 & ~x291;
assign c8143 =  x413 &  x468 & ~x556 & ~x745;
assign c8145 =  x602 & ~x90 & ~x215 & ~x242 & ~x243 & ~x244 & ~x272 & ~x299 & ~x326 & ~x354 & ~x356 & ~x359;
assign c8147 = ~x18 & ~x27 & ~x28 & ~x60 & ~x86 & ~x141 & ~x143 & ~x302 & ~x359 & ~x364 & ~x367 & ~x417 & ~x456 & ~x458 & ~x459 & ~x460 & ~x461 & ~x462 & ~x474 & ~x502 & ~x527 & ~x586 & ~x617 & ~x638 & ~x650 & ~x721 & ~x753 & ~x762;
assign c8149 = ~x196 & ~x215 & ~x242 & ~x243 & ~x244 & ~x260 & ~x272 & ~x273 & ~x302 & ~x331 & ~x656 & ~x657;
assign c8151 =  x264 &  x491 & ~x1 & ~x13 & ~x24 & ~x30 & ~x51 & ~x54 & ~x71 & ~x91 & ~x100 & ~x135 & ~x155 & ~x156 & ~x157 & ~x176 & ~x196 & ~x199 & ~x204 & ~x225 & ~x228 & ~x231 & ~x260 & ~x285 & ~x312 & ~x341 & ~x359 & ~x364 & ~x395 & ~x418 & ~x475 & ~x498 & ~x515 & ~x552 & ~x584 & ~x609 & ~x638 & ~x640 & ~x666 & ~x672 & ~x721 & ~x726 & ~x727 & ~x753 & ~x773;
assign c8153 =  x629 &  x630 & ~x242 & ~x243 & ~x244 & ~x302 & ~x304 & ~x354 & ~x361 & ~x718;
assign c8155 =  x436 &  x491 &  x519 & ~x8 & ~x37 & ~x45 & ~x65 & ~x99 & ~x113 & ~x116 & ~x131 & ~x155 & ~x156 & ~x157 & ~x166 & ~x253 & ~x257 & ~x284 & ~x414 & ~x480 & ~x496 & ~x500 & ~x550 & ~x569 & ~x589 & ~x596 & ~x606 & ~x691 & ~x697 & ~x706 & ~x719 & ~x776;
assign c8157 =  x353 &  x381 &  x436 & ~x122 & ~x575 & ~x630 & ~x631 & ~x658;
assign c8159 =  x408 &  x436 &  x437 & ~x24 & ~x41 & ~x65 & ~x116 & ~x166 & ~x310 & ~x419 & ~x603 & ~x630 & ~x631 & ~x657 & ~x658 & ~x659 & ~x693 & ~x722 & ~x766;
assign c8161 =  x468 &  x496 &  x522 &  x550 & ~x5 & ~x20 & ~x86 & ~x137 & ~x223 & ~x392 & ~x418 & ~x448 & ~x502 & ~x617 & ~x638 & ~x643 & ~x670 & ~x738 & ~x775 & ~x783;
assign c8163 = ~x1 & ~x9 & ~x19 & ~x27 & ~x28 & ~x29 & ~x34 & ~x66 & ~x71 & ~x89 & ~x143 & ~x277 & ~x278 & ~x330 & ~x331 & ~x357 & ~x392 & ~x420 & ~x458 & ~x459 & ~x460 & ~x461 & ~x462 & ~x500 & ~x517 & ~x518 & ~x642 & ~x697 & ~x704 & ~x749 & ~x765 & ~x778 & ~x779 & ~x782;
assign c8165 =  x182 &  x209 &  x578 &  x579 &  x606 & ~x53 & ~x56 & ~x134 & ~x143 & ~x171 & ~x246 & ~x250 & ~x273 & ~x275 & ~x279 & ~x303 & ~x313 & ~x331 & ~x366 & ~x391 & ~x451 & ~x491 & ~x507 & ~x510 & ~x641 & ~x696 & ~x757 & ~x772 & ~x776;
assign c8167 =  x438 &  x439 &  x466 &  x493 &  x494 & ~x16 & ~x17 & ~x23 & ~x43 & ~x51 & ~x88 & ~x104 & ~x114 & ~x165 & ~x196 & ~x226 & ~x279 & ~x341 & ~x447 & ~x451 & ~x477 & ~x617 & ~x640 & ~x641 & ~x670 & ~x703 & ~x706 & ~x729 & ~x731 & ~x741 & ~x747 & ~x768 & ~x769 & ~x774 & ~x778 & ~x783;
assign c8169 = ~x249 & ~x261 & ~x274 & ~x283 & ~x286 & ~x316 & ~x336 & ~x447 & ~x628 & ~x629 & ~x656 & ~x657 & ~x669 & ~x729 & ~x737 & ~x755 & ~x759;
assign c8171 = ~x184 & ~x185 & ~x211 & ~x214 & ~x628;
assign c8173 = ~x24 & ~x34 & ~x107 & ~x326 & ~x352 & ~x354 & ~x380 & ~x381 & ~x410 & ~x459 & ~x487 & ~x530 & ~x646 & ~x669 & ~x727 & ~x742 & ~x773;
assign c8175 = ~x2 & ~x5 & ~x21 & ~x51 & ~x59 & ~x69 & ~x71 & ~x74 & ~x76 & ~x77 & ~x83 & ~x86 & ~x96 & ~x126 & ~x127 & ~x137 & ~x153 & ~x154 & ~x155 & ~x156 & ~x157 & ~x182 & ~x183 & ~x184 & ~x185 & ~x191 & ~x197 & ~x250 & ~x448 & ~x499 & ~x555 & ~x565 & ~x581 & ~x593 & ~x608 & ~x614 & ~x617 & ~x618 & ~x634 & ~x635 & ~x669 & ~x689 & ~x702 & ~x728 & ~x731 & ~x733 & ~x783;
assign c8177 =  x264 &  x346 &  x491 & ~x9 & ~x18 & ~x41 & ~x47 & ~x93 & ~x106 & ~x121 & ~x156 & ~x157 & ~x177 & ~x359 & ~x369 & ~x421 & ~x475 & ~x501 & ~x514 & ~x582 & ~x593 & ~x640 & ~x642 & ~x676 & ~x702 & ~x722 & ~x753 & ~x757 & ~x770 & ~x776;
assign c8179 =  x468 &  x496 & ~x459 & ~x639 & ~x702;
assign c8181 =  x438 &  x466 & ~x243 & ~x272 & ~x518;
assign c8183 =  x353 &  x381 &  x436 &  x437 &  x465 & ~x128 & ~x155 & ~x156 & ~x157 & ~x702 & ~x751 & ~x776 & ~x780;
assign c8185 = ~x406 & ~x407 & ~x408 & ~x769;
assign c8187 =  x296 & ~x237 & ~x263 & ~x264 & ~x291 & ~x320 & ~x356 & ~x753;
assign c8189 =  x268 &  x296 &  x297 & ~x8 & ~x68 & ~x77 & ~x87 & ~x249 & ~x265 & ~x273 & ~x318 & ~x319 & ~x371 & ~x622 & ~x716 & ~x753;
assign c8191 = ~x46 & ~x89 & ~x307 & ~x320 & ~x321 & ~x348 & ~x367 & ~x376 & ~x402 & ~x464 & ~x474;
assign c8193 =  x353 &  x381 &  x491 & ~x35 & ~x40 & ~x115 & ~x118 & ~x155 & ~x156 & ~x190 & ~x359 & ~x510 & ~x538 & ~x577 & ~x646 & ~x770;
assign c8195 =  x401 &  x431 & ~x6 & ~x8 & ~x51 & ~x52 & ~x54 & ~x60 & ~x70 & ~x82 & ~x89 & ~x91 & ~x117 & ~x118 & ~x148 & ~x198 & ~x250 & ~x251 & ~x282 & ~x285 & ~x308 & ~x314 & ~x331 & ~x333 & ~x337 & ~x342 & ~x392 & ~x417 & ~x445 & ~x446 & ~x447 & ~x449 & ~x451 & ~x502 & ~x557 & ~x560 & ~x587 & ~x589 & ~x642 & ~x650 & ~x657 & ~x658 & ~x668 & ~x708 & ~x715 & ~x724 & ~x729 & ~x743 & ~x753 & ~x756 & ~x760 & ~x768 & ~x780;
assign c8197 =  x552 &  x553 &  x578 &  x579 &  x580 & ~x329;
assign c8199 =  x208 &  x209 &  x210 &  x211 &  x212 & ~x20 & ~x25 & ~x53 & ~x64 & ~x165 & ~x169 & ~x197 & ~x293 & ~x367 & ~x486 & ~x490 & ~x762;
assign c8201 =  x429 & ~x260 & ~x286 & ~x330 & ~x331 & ~x378 & ~x379 & ~x640;
assign c8203 =  x466 &  x493 &  x494 &  x521 &  x522 &  x549 & ~x8 & ~x9 & ~x11 & ~x21 & ~x28 & ~x38 & ~x44 & ~x54 & ~x57 & ~x59 & ~x80 & ~x96 & ~x98 & ~x105 & ~x113 & ~x119 & ~x122 & ~x162 & ~x165 & ~x168 & ~x170 & ~x196 & ~x198 & ~x227 & ~x251 & ~x277 & ~x286 & ~x310 & ~x339 & ~x364 & ~x368 & ~x396 & ~x416 & ~x418 & ~x452 & ~x471 & ~x474 & ~x554 & ~x561 & ~x564 & ~x585 & ~x586 & ~x592 & ~x608 & ~x622 & ~x640 & ~x669 & ~x675 & ~x709 & ~x725 & ~x727 & ~x739 & ~x740 & ~x743 & ~x753 & ~x777;
assign c8205 =  x439 &  x466 &  x467 &  x494 &  x495 &  x522 & ~x4 & ~x21 & ~x24 & ~x47 & ~x62 & ~x76 & ~x83 & ~x86 & ~x122 & ~x126 & ~x172 & ~x201 & ~x221 & ~x250 & ~x336 & ~x364 & ~x558 & ~x589 & ~x619 & ~x620 & ~x668 & ~x679 & ~x693 & ~x696 & ~x700 & ~x727 & ~x739 & ~x751 & ~x779;
assign c8207 =  x212 &  x240 &  x267 &  x268 &  x295 &  x296 & ~x107 & ~x244 & ~x274 & ~x307 & ~x319 & ~x340 & ~x382 & ~x640 & ~x671 & ~x719;
assign c8209 = ~x13 & ~x87 & ~x117 & ~x225 & ~x270 & ~x271 & ~x274 & ~x327 & ~x328 & ~x451 & ~x461 & ~x477 & ~x486 & ~x487 & ~x640 & ~x745 & ~x749;
assign c8211 =  x212 &  x213 &  x215 &  x626 &  x630 &  x655 & ~x0 & ~x13 & ~x14 & ~x16 & ~x19 & ~x24 & ~x26 & ~x36 & ~x47 & ~x53 & ~x74 & ~x98 & ~x99 & ~x101 & ~x118 & ~x120 & ~x121 & ~x122 & ~x137 & ~x138 & ~x141 & ~x170 & ~x199 & ~x222 & ~x223 & ~x251 & ~x254 & ~x302 & ~x305 & ~x310 & ~x331 & ~x336 & ~x338 & ~x364 & ~x367 & ~x369 & ~x386 & ~x387 & ~x420 & ~x421 & ~x444 & ~x448 & ~x471 & ~x474 & ~x476 & ~x517 & ~x527 & ~x586 & ~x667 & ~x668 & ~x676 & ~x677 & ~x704 & ~x727 & ~x742 & ~x745 & ~x758 & ~x773 & ~x774;
assign c8213 =  x434 & ~x49 & ~x88 & ~x105 & ~x173 & ~x249 & ~x250 & ~x320 & ~x321 & ~x348 & ~x376 & ~x397 & ~x402 & ~x404 & ~x449 & ~x647 & ~x740;
assign c8215 =  x212 &  x213 &  x215 &  x238 &  x239 &  x240 &  x241 &  x242 &  x243 &  x244 & ~x2 & ~x16 & ~x24 & ~x35 & ~x60 & ~x88 & ~x111 & ~x284 & ~x366 & ~x391 & ~x395 & ~x474 & ~x543 & ~x644 & ~x648 & ~x666 & ~x709 & ~x718 & ~x727 & ~x735 & ~x750;
assign c8217 = ~x378 & ~x379 & ~x380 & ~x381 & ~x408 & ~x418 & ~x437 & ~x781;
assign c8219 = ~x41 & ~x88 & ~x142 & ~x169 & ~x286 & ~x474 & ~x614 & ~x628 & ~x629 & ~x630 & ~x631 & ~x638 & ~x656 & ~x657 & ~x658 & ~x659 & ~x669 & ~x687 & ~x720 & ~x722 & ~x759;
assign c8221 =  x412 &  x468 &  x523 & ~x474;
assign c8223 =  x508;
assign c8225 =  x239 &  x267 &  x268 &  x294 &  x296 & ~x41 & ~x244 & ~x302 & ~x355;
assign c8227 =  x182 &  x209 & ~x22 & ~x119 & ~x169 & ~x171 & ~x272 & ~x273 & ~x274 & ~x281 & ~x298 & ~x303 & ~x325 & ~x326 & ~x332 & ~x343 & ~x354 & ~x355 & ~x371 & ~x448 & ~x502 & ~x508 & ~x534 & ~x560 & ~x590 & ~x694 & ~x716 & ~x718 & ~x757 & ~x778;
assign c8229 =  x214 &  x242 &  x269 &  x297 &  x325 &  x352 &  x406 & ~x27 & ~x67 & ~x77 & ~x81 & ~x85 & ~x90 & ~x94 & ~x115 & ~x136 & ~x193 & ~x253 & ~x286 & ~x308 & ~x313 & ~x319 & ~x320 & ~x330 & ~x364 & ~x444 & ~x446 & ~x448 & ~x452 & ~x479 & ~x502 & ~x593 & ~x643 & ~x673 & ~x690 & ~x712 & ~x728 & ~x738 & ~x742 & ~x748 & ~x753 & ~x767 & ~x775;
assign c8231 =  x630 & ~x403 & ~x404 & ~x405 & ~x432;
assign c8233 = ~x11 & ~x275 & ~x321 & ~x364 & ~x479 & ~x614 & ~x628 & ~x630 & ~x631 & ~x656 & ~x657 & ~x658 & ~x683 & ~x731;
assign c8235 =  x439 &  x466 &  x467 &  x494 &  x522 &  x549;
assign c8237 =  x102;
assign c8239 =  x411 &  x439 &  x466 &  x467 &  x494 &  x521 & ~x1 & ~x169 & ~x196 & ~x415 & ~x638 & ~x675 & ~x732 & ~x764 & ~x783;
assign c8241 = ~x216 & ~x244 & ~x261 & ~x291 & ~x326 & ~x330 & ~x354 & ~x437 & ~x665 & ~x724;
assign c8243 =  x268 &  x269 &  x296 &  x297 &  x298 & ~x155 & ~x182;
assign c8245 =  x214 &  x215 &  x216 & ~x13 & ~x20 & ~x28 & ~x32 & ~x34 & ~x44 & ~x50 & ~x64 & ~x79 & ~x87 & ~x104 & ~x106 & ~x118 & ~x143 & ~x253 & ~x305 & ~x339 & ~x353 & ~x361 & ~x366 & ~x381 & ~x382 & ~x421 & ~x477 & ~x517 & ~x529 & ~x530 & ~x534 & ~x585 & ~x614 & ~x669 & ~x700 & ~x711 & ~x731 & ~x745 & ~x746 & ~x762 & ~x780 & ~x782;
assign c8247 = ~x405 & ~x434 & ~x436 & ~x464;
assign c8249 =  x268 &  x296 & ~x2 & ~x12 & ~x16 & ~x56 & ~x264 & ~x286 & ~x290 & ~x308 & ~x318 & ~x319 & ~x320 & ~x399 & ~x590 & ~x591 & ~x614 & ~x641 & ~x706 & ~x753;
assign c8251 =  x296 & ~x51 & ~x235 & ~x236 & ~x248 & ~x275 & ~x289 & ~x291 & ~x300 & ~x319 & ~x343 & ~x373 & ~x665;
assign c8253 =  x629 &  x630 & ~x170 & ~x280 & ~x455 & ~x457 & ~x459 & ~x460 & ~x461 & ~x474 & ~x477 & ~x487 & ~x490 & ~x502 & ~x504 & ~x514 & ~x640 & ~x718 & ~x744 & ~x757 & ~x763 & ~x769;
assign c8255 =  x426;
assign c8257 =  x436 & ~x34 & ~x127 & ~x151 & ~x154 & ~x155 & ~x156 & ~x157 & ~x250 & ~x392 & ~x486 & ~x585 & ~x622 & ~x640 & ~x649 & ~x669 & ~x690;
assign c8259 =  x381 & ~x248 & ~x339 & ~x350 & ~x376 & ~x378 & ~x404 & ~x644;
assign c8261 = ~x1 & ~x47 & ~x72 & ~x85 & ~x88 & ~x283 & ~x341 & ~x354 & ~x378 & ~x379 & ~x380 & ~x381 & ~x668;
assign c8263 =  x437 &  x465 &  x466 &  x493 &  x519 & ~x2 & ~x12 & ~x14 & ~x28 & ~x29 & ~x41 & ~x60 & ~x66 & ~x69 & ~x71 & ~x82 & ~x86 & ~x88 & ~x119 & ~x141 & ~x164 & ~x176 & ~x198 & ~x202 & ~x257 & ~x331 & ~x341 & ~x359 & ~x364 & ~x366 & ~x389 & ~x416 & ~x445 & ~x478 & ~x560 & ~x587 & ~x620 & ~x636 & ~x641 & ~x668 & ~x697 & ~x716 & ~x733 & ~x742 & ~x753 & ~x756 & ~x771 & ~x778;
assign c8265 = ~x380 & ~x406 & ~x407 & ~x436;
assign c8267 =  x433 & ~x6 & ~x35 & ~x53 & ~x116 & ~x136 & ~x167 & ~x295 & ~x316 & ~x321 & ~x322 & ~x348 & ~x349 & ~x376 & ~x476 & ~x503 & ~x643 & ~x754;
assign c8269 =  x266 & ~x28 & ~x48 & ~x77 & ~x135 & ~x186 & ~x215 & ~x216 & ~x242 & ~x244 & ~x449 & ~x609 & ~x633 & ~x634 & ~x663 & ~x707;
assign c8271 =  x381 & ~x295 & ~x321 & ~x348 & ~x349 & ~x376 & ~x402 & ~x690;
assign c8273 =  x437 &  x438 & ~x5 & ~x7 & ~x25 & ~x29 & ~x82 & ~x111 & ~x125 & ~x274 & ~x294 & ~x301 & ~x359 & ~x392 & ~x448 & ~x474 & ~x475 & ~x490 & ~x532 & ~x666 & ~x720 & ~x746 & ~x765 & ~x774 & ~x782;
assign c8275 =  x400 &  x428 & ~x73 & ~x203 & ~x230 & ~x278 & ~x339 & ~x349 & ~x350 & ~x507 & ~x562 & ~x615 & ~x651 & ~x722 & ~x766;
assign c8277 = ~x12 & ~x29 & ~x44 & ~x51 & ~x99 & ~x102 & ~x117 & ~x171 & ~x272 & ~x274 & ~x300 & ~x301 & ~x302 & ~x459 & ~x460 & ~x461 & ~x474 & ~x481 & ~x518 & ~x585 & ~x592 & ~x614 & ~x644 & ~x648 & ~x650 & ~x715 & ~x728 & ~x736 & ~x753;
assign c8279 =  x525 &  x552 &  x578 &  x579 & ~x2 & ~x18 & ~x164 & ~x278 & ~x340 & ~x423 & ~x562 & ~x678 & ~x716 & ~x739 & ~x748 & ~x757;
assign c8281 =  x601 & ~x243 & ~x260 & ~x271 & ~x326;
assign c8283 = ~x14 & ~x51 & ~x89 & ~x113 & ~x278 & ~x354 & ~x362 & ~x380 & ~x381 & ~x408 & ~x436 & ~x464 & ~x592 & ~x727 & ~x733;
assign c8285 =  x296 &  x297 & ~x182 & ~x631 & ~x659;
assign c8287 = ~x66 & ~x74 & ~x88 & ~x101 & ~x110 & ~x119 & ~x121 & ~x138 & ~x198 & ~x199 & ~x379 & ~x389 & ~x435 & ~x436 & ~x447 & ~x452 & ~x474 & ~x502 & ~x530 & ~x586 & ~x592 & ~x617 & ~x649 & ~x716 & ~x742 & ~x753 & ~x757 & ~x778;
assign c8289 = ~x216 & ~x244 & ~x261 & ~x271 & ~x272 & ~x273 & ~x328 & ~x657 & ~x658;
assign c8291 =  x271 &  x621;
assign c8293 = ~x141 & ~x294 & ~x340 & ~x349 & ~x367 & ~x376 & ~x404 & ~x431 & ~x451 & ~x641 & ~x702 & ~x733 & ~x773 & ~x781;
assign c8295 =  x381 &  x437 &  x491 &  x492 & ~x1 & ~x6 & ~x20 & ~x64 & ~x69 & ~x79 & ~x81 & ~x132 & ~x136 & ~x138 & ~x143 & ~x145 & ~x171 & ~x174 & ~x193 & ~x201 & ~x224 & ~x227 & ~x251 & ~x275 & ~x311 & ~x334 & ~x336 & ~x338 & ~x366 & ~x367 & ~x390 & ~x396 & ~x418 & ~x473 & ~x474 & ~x479 & ~x501 & ~x506 & ~x530 & ~x534 & ~x559 & ~x562 & ~x577 & ~x615 & ~x635 & ~x663 & ~x669 & ~x689 & ~x717 & ~x729 & ~x737 & ~x742 & ~x753 & ~x761;
assign c8297 =  x354 &  x381 &  x382 &  x409 &  x437 &  x465 &  x491 &  x519 &  x546 & ~x37 & ~x41 & ~x81 & ~x97 & ~x100 & ~x251 & ~x361 & ~x559 & ~x586 & ~x645 & ~x675 & ~x690 & ~x720 & ~x742 & ~x769;
assign c8299 = ~x121 & ~x155 & ~x156 & ~x157 & ~x182 & ~x183 & ~x184 & ~x185 & ~x210 & ~x211 & ~x212 & ~x721 & ~x731;
assign c90 =  x392;
assign c92 =  x210 &  x343 &  x411 &  x439 & ~x653;
assign c94 =  x340;
assign c96 =  x378 & ~x304 & ~x466 & ~x486 & ~x540 & ~x551 & ~x593 & ~x605 & ~x629;
assign c98 =  x432 &  x518 & ~x95 & ~x134 & ~x191 & ~x200 & ~x222 & ~x324 & ~x448 & ~x495 & ~x522 & ~x549 & ~x576 & ~x577 & ~x632 & ~x635 & ~x659 & ~x660 & ~x756;
assign c910 =  x209 &  x235 &  x317 &  x345 & ~x73 & ~x145 & ~x202 & ~x246 & ~x511 & ~x568 & ~x571 & ~x572 & ~x600 & ~x622 & ~x626 & ~x627 & ~x628;
assign c912 =  x368;
assign c914 =  x208 &  x343 & ~x602 & ~x650 & ~x684;
assign c916 =  x292 &  x380 & ~x6 & ~x25 & ~x38 & ~x53 & ~x57 & ~x58 & ~x67 & ~x73 & ~x89 & ~x112 & ~x122 & ~x125 & ~x138 & ~x146 & ~x166 & ~x171 & ~x201 & ~x231 & ~x234 & ~x248 & ~x253 & ~x256 & ~x288 & ~x304 & ~x316 & ~x332 & ~x370 & ~x372 & ~x397 & ~x411 & ~x422 & ~x439 & ~x440 & ~x446 & ~x451 & ~x467 & ~x479 & ~x484 & ~x493 & ~x494 & ~x496 & ~x500 & ~x503 & ~x514 & ~x521 & ~x523 & ~x534 & ~x549 & ~x550 & ~x551 & ~x558 & ~x577 & ~x591 & ~x596 & ~x605 & ~x615 & ~x618 & ~x633 & ~x636 & ~x663 & ~x673 & ~x676 & ~x689 & ~x722 & ~x734 & ~x737 & ~x759 & ~x769 & ~x774 & ~x776 & ~x779;
assign c918 =  x717 & ~x580 & ~x658;
assign c920 =  x238 & ~x65 & ~x169 & ~x496 & ~x525 & ~x546 & ~x552 & ~x573 & ~x602 & ~x630 & ~x657 & ~x658 & ~x684 & ~x686 & ~x701;
assign c922 =  x705;
assign c924 =  x236 &  x343 & ~x7 & ~x13 & ~x26 & ~x61 & ~x78 & ~x126 & ~x137 & ~x170 & ~x217 & ~x227 & ~x303 & ~x444 & ~x480 & ~x543 & ~x559 & ~x571 & ~x608 & ~x668 & ~x678 & ~x706;
assign c926 =  x352 &  x380 & ~x57 & ~x71 & ~x84 & ~x109 & ~x186 & ~x466 & ~x476 & ~x510 & ~x514 & ~x522 & ~x550 & ~x572 & ~x581 & ~x653;
assign c928 =  x205 &  x341;
assign c930 =  x209 &  x212 &  x317 &  x410 & ~x206 & ~x223 & ~x294;
assign c932 =  x214 &  x317 &  x410 &  x438 &  x465 &  x493 & ~x256 & ~x498 & ~x734;
assign c934 =  x209 &  x213 &  x317 &  x373 &  x492 & ~x479 & ~x523 & ~x596 & ~x605;
assign c936 =  x180 &  x316 & ~x11 & ~x96 & ~x138 & ~x277 & ~x303 & ~x366 & ~x560 & ~x571 & ~x572 & ~x764;
assign c938 =  x714 & ~x132 & ~x158 & ~x233 & ~x234 & ~x288 & ~x570 & ~x572 & ~x599 & ~x600 & ~x626 & ~x627 & ~x628 & ~x653 & ~x767;
assign c940 =  x213 &  x353 & ~x46 & ~x48 & ~x50 & ~x67 & ~x74 & ~x94 & ~x112 & ~x117 & ~x153 & ~x160 & ~x170 & ~x220 & ~x228 & ~x233 & ~x234 & ~x252 & ~x258 & ~x286 & ~x336 & ~x425 & ~x439 & ~x441 & ~x445 & ~x448 & ~x469 & ~x480 & ~x521 & ~x522 & ~x525 & ~x533 & ~x549 & ~x552 & ~x553 & ~x555 & ~x558 & ~x560 & ~x567 & ~x577 & ~x578 & ~x580 & ~x605 & ~x611 & ~x613 & ~x617 & ~x618 & ~x635 & ~x664 & ~x665 & ~x667 & ~x706 & ~x751 & ~x769 & ~x776;
assign c942 =  x465 &  x492 &  x520 &  x548 &  x576 &  x603 &  x631 & ~x17 & ~x38 & ~x91 & ~x104 & ~x145 & ~x156 & ~x158 & ~x159 & ~x175 & ~x189 & ~x199 & ~x247 & ~x251 & ~x304 & ~x334 & ~x358 & ~x364 & ~x385 & ~x426 & ~x439 & ~x440 & ~x450 & ~x472 & ~x497 & ~x526 & ~x557 & ~x560 & ~x571 & ~x572 & ~x578 & ~x600 & ~x623 & ~x650 & ~x651 & ~x653 & ~x654 & ~x664 & ~x681 & ~x682 & ~x723;
assign c944 =  x185 &  x214 &  x410 &  x438 &  x492 &  x493 &  x520 & ~x9 & ~x13 & ~x75 & ~x510 & ~x552 & ~x553 & ~x563 & ~x662 & ~x723;
assign c946 =  x352 & ~x27 & ~x98 & ~x158 & ~x214 & ~x463 & ~x543 & ~x572 & ~x573 & ~x653 & ~x681;
assign c948 =  x353 &  x519 & ~x18 & ~x28 & ~x94 & ~x124 & ~x151 & ~x153 & ~x197 & ~x233 & ~x276 & ~x280 & ~x313 & ~x343 & ~x398 & ~x450 & ~x467 & ~x497 & ~x524 & ~x533 & ~x536 & ~x549 & ~x576 & ~x577 & ~x589 & ~x604 & ~x631 & ~x632 & ~x661 & ~x686 & ~x743;
assign c950 =  x639;
assign c952 =  x214 &  x238 &  x409 & ~x207 & ~x232 & ~x387 & ~x601 & ~x628 & ~x629 & ~x657;
assign c954 =  x385 &  x396;
assign c956 = ~x187 & ~x234 & ~x493 & ~x520 & ~x548 & ~x627;
assign c958 =  x356 &  x383 &  x411 &  x438 &  x439 &  x466 & ~x572 & ~x661;
assign c960 =  x210 &  x316 &  x411 &  x439 &  x466;
assign c962 =  x693;
assign c964 =  x491 & ~x54 & ~x86 & ~x144 & ~x158 & ~x159 & ~x234 & ~x247 & ~x254 & ~x286 & ~x315 & ~x439 & ~x477 & ~x499 & ~x521 & ~x549 & ~x576 & ~x577 & ~x578 & ~x604 & ~x605 & ~x632 & ~x661 & ~x673 & ~x687 & ~x716 & ~x737 & ~x767;
assign c966 =  x236 &  x372 &  x438 &  x465 &  x493 & ~x202 & ~x205 & ~x306 & ~x330 & ~x426 & ~x501 & ~x664;
assign c968 =  x263 & ~x187 & ~x232 & ~x233 & ~x462 & ~x468 & ~x523 & ~x572 & ~x699 & ~x719 & ~x759;
assign c970 =  x181 &  x385 &  x496;
assign c972 =  x368 &  x426 &  x455 & ~x347;
assign c974 =  x719;
assign c976 =  x342 & ~x344;
assign c978 =  x263 &  x317 &  x372 &  x410 & ~x15 & ~x68 & ~x110 & ~x314 & ~x320 & ~x663 & ~x674 & ~x728;
assign c980 =  x212 &  x319 & ~x11 & ~x25 & ~x26 & ~x61 & ~x67 & ~x70 & ~x93 & ~x149 & ~x175 & ~x204 & ~x217 & ~x220 & ~x222 & ~x233 & ~x247 & ~x261 & ~x287 & ~x289 & ~x306 & ~x307 & ~x310 & ~x365 & ~x371 & ~x394 & ~x412 & ~x414 & ~x427 & ~x439 & ~x443 & ~x452 & ~x470 & ~x477 & ~x502 & ~x503 & ~x507 & ~x536 & ~x541 & ~x549 & ~x554 & ~x560 & ~x563 & ~x577 & ~x585 & ~x632 & ~x653 & ~x676 & ~x689 & ~x693 & ~x719 & ~x721 & ~x749 & ~x751 & ~x762;
assign c982 =  x688 &  x716 & ~x599 & ~x685;
assign c984 =  x662 &  x719 & ~x687;
assign c986 =  x180 &  x383 &  x411 & ~x236 & ~x525;
assign c988 =  x182 &  x263 & ~x17 & ~x165 & ~x204 & ~x205 & ~x233 & ~x629 & ~x730 & ~x781;
assign c990 =  x209 &  x436 & ~x188 & ~x205 & ~x222 & ~x249 & ~x276 & ~x307 & ~x466 & ~x526 & ~x531 & ~x541 & ~x549 & ~x554 & ~x557 & ~x576 & ~x577 & ~x626 & ~x632;
assign c992 =  x710 & ~x190 & ~x207 & ~x365 & ~x631 & ~x632 & ~x658 & ~x685;
assign c994 =  x342 &  x439 & ~x346 & ~x660;
assign c996 =  x328 &  x407 &  x438;
assign c998 =  x722;
assign c9100 =  x211 &  x317 &  x345 &  x407 &  x464 &  x492 & ~x72 & ~x112 & ~x160 & ~x258 & ~x331 & ~x342 & ~x425 & ~x479 & ~x522 & ~x567 & ~x605 & ~x642 & ~x723 & ~x734 & ~x736;
assign c9102 =  x369;
assign c9104 = ~x204 & ~x404 & ~x519 & ~x546 & ~x573 & ~x574 & ~x575 & ~x602 & ~x628 & ~x629 & ~x630 & ~x657 & ~x658 & ~x686;
assign c9106 =  x208 &  x343 &  x371 & ~x628 & ~x683;
assign c9108 =  x23;
assign c9110 =  x185 &  x215 & ~x206 & ~x603 & ~x630 & ~x658 & ~x686;
assign c9112 =  x242 &  x376 & ~x493 & ~x576 & ~x658;
assign c9114 =  x292 &  x319 & ~x19 & ~x57 & ~x59 & ~x65 & ~x90 & ~x102 & ~x132 & ~x190 & ~x208 & ~x234 & ~x235 & ~x236 & ~x275 & ~x280 & ~x286 & ~x310 & ~x316 & ~x336 & ~x338 & ~x451 & ~x504 & ~x522 & ~x549 & ~x550 & ~x560 & ~x563 & ~x576 & ~x577 & ~x586 & ~x604 & ~x624 & ~x659 & ~x660 & ~x673 & ~x691 & ~x696;
assign c9116 =  x546 &  x712 & ~x232 & ~x571 & ~x605 & ~x632;
assign c9118 =  x186 &  x292 & ~x549 & ~x603 & ~x631 & ~x658;
assign c9120 =  x693;
assign c9122 =  x236 &  x492 &  x575 & ~x89 & ~x105 & ~x109 & ~x166 & ~x174 & ~x201 & ~x202 & ~x217 & ~x283 & ~x312 & ~x388 & ~x496 & ~x572 & ~x578 & ~x583 & ~x599 & ~x600 & ~x626 & ~x627 & ~x655 & ~x663 & ~x674 & ~x683;
assign c9124 =  x721;
assign c9126 =  x186 & ~x137 & ~x426 & ~x538 & ~x568 & ~x575 & ~x629 & ~x645 & ~x685 & ~x724;
assign c9128 =  x206 &  x413 &  x441 &  x496;
assign c9130 =  x328 &  x681;
assign c9132 =  x355 &  x410 & ~x205 & ~x232 & ~x549 & ~x604 & ~x631;
assign c9134 =  x545 & ~x235 & ~x541;
assign c9136 =  x323 &  x347 &  x350 & ~x15 & ~x98 & ~x133 & ~x158 & ~x160 & ~x187 & ~x218 & ~x245 & ~x302 & ~x385 & ~x423 & ~x425 & ~x439 & ~x469 & ~x515 & ~x592 & ~x663 & ~x766;
assign c9138 =  x181 &  x353 &  x465 & ~x123 & ~x243 & ~x571 & ~x572 & ~x583;
assign c9140 =  x766;
assign c9142 =  x721;
assign c9144 =  x371 &  x399 &  x485 & ~x442 & ~x623;
assign c9146 =  x737;
assign c9148 =  x263 &  x465 &  x493 &  x520 &  x548 & ~x89 & ~x219 & ~x247 & ~x441 & ~x504 & ~x527 & ~x573 & ~x600 & ~x681;
assign c9150 =  x378 & ~x295 & ~x438 & ~x604;
assign c9152 =  x643;
assign c9154 =  x319 &  x352 &  x380 &  x435 & ~x3 & ~x4 & ~x56 & ~x70 & ~x82 & ~x125 & ~x159 & ~x172 & ~x194 & ~x198 & ~x232 & ~x233 & ~x250 & ~x260 & ~x304 & ~x331 & ~x342 & ~x356 & ~x391 & ~x410 & ~x417 & ~x447 & ~x448 & ~x511 & ~x522 & ~x577 & ~x646 & ~x702 & ~x718 & ~x720 & ~x734 & ~x738 & ~x764 & ~x765 & ~x767;
assign c9156 =  x214 &  x263 &  x408 &  x410 &  x437 &  x465 &  x492 & ~x1 & ~x81 & ~x137 & ~x149 & ~x205 & ~x222 & ~x233 & ~x388 & ~x416 & ~x470 & ~x534 & ~x590 & ~x606 & ~x653 & ~x662 & ~x671;
assign c9158 = ~x6 & ~x7 & ~x78 & ~x94 & ~x115 & ~x118 & ~x144 & ~x189 & ~x195 & ~x213 & ~x244 & ~x245 & ~x256 & ~x275 & ~x329 & ~x336 & ~x449 & ~x471 & ~x503 & ~x540 & ~x571 & ~x572 & ~x573 & ~x600 & ~x601 & ~x602 & ~x626 & ~x628 & ~x629 & ~x630 & ~x657 & ~x658 & ~x671 & ~x686 & ~x705 & ~x713;
assign c9160 =  x292 & ~x235 & ~x344 & ~x495 & ~x548 & ~x575 & ~x658;
assign c9162 =  x319 &  x383 & ~x208 & ~x233;
assign c9164 =  x710;
assign c9166 =  x292 &  x383 &  x410 &  x437 & ~x49 & ~x88 & ~x140 & ~x202 & ~x234 & ~x338 & ~x613 & ~x726;
assign c9168 =  x180 &  x315 &  x410 & ~x218;
assign c9170 =  x215 &  x329 &  x357 &  x385;
assign c9172 =  x463 & ~x12 & ~x78 & ~x99 & ~x105 & ~x126 & ~x160 & ~x206 & ~x229 & ~x260 & ~x304 & ~x420 & ~x467 & ~x468 & ~x484 & ~x496 & ~x508 & ~x520 & ~x536 & ~x548 & ~x569 & ~x575 & ~x577 & ~x596 & ~x623 & ~x631 & ~x632 & ~x647 & ~x658 & ~x688 & ~x689;
assign c9174 =  x341 & ~x319;
assign c9176 =  x342 & ~x575;
assign c9178 =  x235 &  x409 &  x493 &  x521 & ~x40 & ~x106 & ~x108 & ~x138 & ~x145 & ~x222 & ~x245 & ~x387 & ~x453 & ~x519 & ~x601 & ~x667;
assign c9180 =  x238 &  x515 & ~x42 & ~x572;
assign c9182 =  x719;
assign c9184 =  x111;
assign c9186 =  x380 &  x493 & ~x5 & ~x57 & ~x129 & ~x159 & ~x187 & ~x205 & ~x256 & ~x257 & ~x330 & ~x397 & ~x425 & ~x511 & ~x563 & ~x572 & ~x573 & ~x653 & ~x663 & ~x696 & ~x707 & ~x730;
assign c9188 =  x408 &  x409 &  x492 &  x547 & ~x16 & ~x34 & ~x49 & ~x119 & ~x121 & ~x153 & ~x189 & ~x217 & ~x232 & ~x308 & ~x439 & ~x522 & ~x523 & ~x571 & ~x572 & ~x577 & ~x593 & ~x600 & ~x605 & ~x699;
assign c9190 =  x343 &  x371 &  x399 &  x410 & ~x6 & ~x347 & ~x536 & ~x626;
assign c9192 =  x237 &  x329 &  x466 &  x521;
assign c9194 =  x208 &  x316 & ~x28 & ~x109 & ~x246 & ~x572 & ~x573 & ~x599 & ~x626 & ~x627 & ~x653 & ~x655;
assign c9196 =  x373 &  x378 & ~x341 & ~x572 & ~x627 & ~x645 & ~x724 & ~x775;
assign c9198 =  x178 &  x691;
assign c9200 =  x403 &  x629 &  x712 & ~x205;
assign c9202 =  x209 &  x548 &  x576 &  x603 & ~x601;
assign c9204 =  x720;
assign c9206 =  x209 &  x288 & ~x51 & ~x165 & ~x215 & ~x218 & ~x419 & ~x500 & ~x531 & ~x601 & ~x626;
assign c9208 =  x209 & ~x243 & ~x546 & ~x572 & ~x573 & ~x600 & ~x601 & ~x602 & ~x628 & ~x629 & ~x683;
assign c9210 =  x342 & ~x145;
assign c9212 =  x342 & ~x73 & ~x145 & ~x290 & ~x317 & ~x347;
assign c9214 =  x179 &  x410 & ~x236 & ~x292;
assign c9216 = ~x50 & ~x60 & ~x72 & ~x102 & ~x131 & ~x152 & ~x158 & ~x189 & ~x201 & ~x205 & ~x215 & ~x220 & ~x233 & ~x247 & ~x253 & ~x257 & ~x303 & ~x313 & ~x339 & ~x386 & ~x419 & ~x439 & ~x446 & ~x474 & ~x494 & ~x509 & ~x511 & ~x521 & ~x522 & ~x539 & ~x549 & ~x553 & ~x572 & ~x577 & ~x586 & ~x599 & ~x600 & ~x605 & ~x624 & ~x627 & ~x671 & ~x703 & ~x728 & ~x736;
assign c9218 =  x180 & ~x7 & ~x39 & ~x75 & ~x215 & ~x217 & ~x245 & ~x302 & ~x385 & ~x542 & ~x568 & ~x572 & ~x573 & ~x601 & ~x624 & ~x653 & ~x681 & ~x705 & ~x708 & ~x738 & ~x748;
assign c9220 =  x407 &  x546 & ~x216 & ~x233 & ~x495 & ~x521 & ~x549 & ~x572 & ~x576 & ~x604 & ~x632 & ~x653;
assign c9222 =  x180 &  x353 &  x437 & ~x32 & ~x34 & ~x215 & ~x265 & ~x385 & ~x447 & ~x513 & ~x517 & ~x676;
assign c9224 =  x763;
assign c9226 =  x185 &  x328 &  x356 &  x384 &  x411 & ~x756;
assign c9228 =  x212 &  x213 &  x404 & ~x521 & ~x548 & ~x549 & ~x576 & ~x604 & ~x631;
assign c9230 =  x181 &  x207 &  x317 & ~x70 & ~x171 & ~x187 & ~x244 & ~x600;
assign c9232 =  x240 &  x319 & ~x208 & ~x412 & ~x549 & ~x582 & ~x604 & ~x631;
assign c9234 =  x356 &  x357 &  x385 &  x439 & ~x295 & ~x322;
assign c9236 =  x325 &  x380 &  x436 & ~x2 & ~x48 & ~x57 & ~x91 & ~x103 & ~x168 & ~x169 & ~x176 & ~x193 & ~x202 & ~x204 & ~x216 & ~x226 & ~x242 & ~x247 & ~x284 & ~x341 & ~x426 & ~x439 & ~x442 & ~x482 & ~x487 & ~x505 & ~x514 & ~x572 & ~x698 & ~x733 & ~x752 & ~x767;
assign c9238 =  x212 &  x240 &  x319 &  x380 & ~x3 & ~x8 & ~x9 & ~x12 & ~x14 & ~x17 & ~x40 & ~x42 & ~x53 & ~x57 & ~x59 & ~x64 & ~x74 & ~x79 & ~x87 & ~x90 & ~x94 & ~x103 & ~x106 & ~x114 & ~x118 & ~x127 & ~x145 & ~x149 & ~x150 & ~x152 & ~x156 & ~x158 & ~x161 & ~x162 & ~x178 & ~x187 & ~x188 & ~x200 & ~x205 & ~x218 & ~x233 & ~x245 & ~x248 & ~x275 & ~x276 & ~x277 & ~x281 & ~x282 & ~x284 & ~x285 & ~x286 & ~x287 & ~x301 & ~x311 & ~x312 & ~x330 & ~x331 & ~x332 & ~x341 & ~x386 & ~x387 & ~x394 & ~x395 & ~x426 & ~x439 & ~x440 & ~x450 & ~x468 & ~x470 & ~x472 & ~x474 & ~x477 & ~x483 & ~x495 & ~x498 & ~x524 & ~x537 & ~x551 & ~x557 & ~x560 & ~x578 & ~x583 & ~x596 & ~x607 & ~x619 & ~x648 & ~x664 & ~x672 & ~x673 & ~x678 & ~x679 & ~x691 & ~x705 & ~x719 & ~x731 & ~x737 & ~x753 & ~x757 & ~x761 & ~x763 & ~x770 & ~x771 & ~x777 & ~x783;
assign c9240 =  x112;
assign c9242 =  x212 &  x238 &  x355 &  x383 &  x410 &  x437 &  x464 &  x465 & ~x7 & ~x31 & ~x49 & ~x144 & ~x145 & ~x179 & ~x206 & ~x257 & ~x367 & ~x470 & ~x496 & ~x636 & ~x664 & ~x692 & ~x706;
assign c9244 =  x214 &  x319 & ~x36 & ~x99 & ~x121 & ~x148 & ~x149 & ~x160 & ~x192 & ~x196 & ~x207 & ~x208 & ~x224 & ~x235 & ~x258 & ~x262 & ~x288 & ~x305 & ~x312 & ~x337 & ~x413 & ~x441 & ~x508 & ~x522 & ~x535 & ~x549 & ~x578 & ~x604 & ~x632 & ~x644 & ~x750;
assign c9246 =  x438 &  x466 &  x493 &  x520 &  x684;
assign c9248 =  x236 & ~x78 & ~x111 & ~x131 & ~x149 & ~x152 & ~x158 & ~x159 & ~x195 & ~x215 & ~x245 & ~x256 & ~x283 & ~x304 & ~x331 & ~x501 & ~x506 & ~x561 & ~x572 & ~x599 & ~x602 & ~x624 & ~x628 & ~x629 & ~x685 & ~x686 & ~x764 & ~x783;
assign c9250 =  x236 & ~x5 & ~x14 & ~x34 & ~x47 & ~x48 & ~x52 & ~x58 & ~x109 & ~x135 & ~x143 & ~x150 & ~x196 & ~x204 & ~x205 & ~x215 & ~x244 & ~x247 & ~x253 & ~x259 & ~x284 & ~x315 & ~x330 & ~x355 & ~x357 & ~x366 & ~x387 & ~x410 & ~x438 & ~x439 & ~x495 & ~x499 & ~x514 & ~x554 & ~x565 & ~x592 & ~x606 & ~x607 & ~x637 & ~x741 & ~x753 & ~x754 & ~x766;
assign c9252 =  x369 & ~x575;
assign c9254 =  x207 &  x208 &  x288 & ~x215 & ~x219 & ~x507 & ~x572 & ~x599 & ~x601 & ~x627;
assign c9256 =  x343 & ~x603 & ~x626 & ~x631 & ~x658;
assign c9258 =  x209 &  x373 & ~x347 & ~x601 & ~x627 & ~x653 & ~x683;
assign c9260 =  x210 &  x211 &  x212 &  x319 & ~x28 & ~x54 & ~x94 & ~x101 & ~x116 & ~x118 & ~x204 & ~x282 & ~x288 & ~x335 & ~x339 & ~x357 & ~x386 & ~x438 & ~x441 & ~x498 & ~x521 & ~x532 & ~x540 & ~x549 & ~x552 & ~x565 & ~x567 & ~x577 & ~x581 & ~x607 & ~x651 & ~x653 & ~x663 & ~x748 & ~x751 & ~x769;
assign c9262 =  x706;
assign c9264 =  x263 &  x492 & ~x204 & ~x234 & ~x247 & ~x257 & ~x522 & ~x586 & ~x599 & ~x600 & ~x622 & ~x628 & ~x653;
assign c9266 =  x185 & ~x439 & ~x548 & ~x549 & ~x566 & ~x575 & ~x603 & ~x604 & ~x658;
assign c9268 =  x345 &  x373 &  x410 &  x437 &  x465 &  x492 &  x493 &  x520 &  x548 & ~x578;
assign c9270 =  x186 &  x237 &  x399;
assign c9272 =  x345 &  x373 & ~x46 & ~x48 & ~x62 & ~x83 & ~x102 & ~x129 & ~x132 & ~x137 & ~x158 & ~x191 & ~x233 & ~x247 & ~x385 & ~x440 & ~x450 & ~x470 & ~x477 & ~x495 & ~x499 & ~x571 & ~x572 & ~x592 & ~x600 & ~x627 & ~x628 & ~x637 & ~x663;
assign c9274 =  x182 &  x208 &  x352 & ~x158 & ~x171 & ~x201 & ~x204 & ~x221 & ~x433 & ~x514 & ~x550 & ~x622;
assign c9276 =  x207 &  x317 &  x409 & ~x215 & ~x363 & ~x764;
assign c9278 =  x263 &  x376 & ~x549 & ~x631;
assign c9280 =  x353 &  x378 & ~x233 & ~x549 & ~x604 & ~x659;
assign c9284 =  x182 &  x235 &  x317 &  x465 &  x493 & ~x217 & ~x342 & ~x571;
assign c9286 =  x234 &  x350 & ~x185;
assign c9288 =  x180 &  x288 &  x410 &  x438 & ~x114 & ~x145 & ~x218 & ~x680;
assign c9290 =  x209 &  x214 &  x372 & ~x415 & ~x599 & ~x627 & ~x636;
assign c9292 =  x212 &  x317 & ~x495 & ~x581 & ~x632;
assign c9294 =  x378 &  x404 & ~x76 & ~x103 & ~x133 & ~x158 & ~x253 & ~x357 & ~x385 & ~x440 & ~x441 & ~x488 & ~x511 & ~x549 & ~x589 & ~x677 & ~x703 & ~x745 & ~x780;
assign c9296 =  x235 & ~x22 & ~x33 & ~x73 & ~x150 & ~x153 & ~x187 & ~x191 & ~x205 & ~x215 & ~x497 & ~x571 & ~x573 & ~x599 & ~x601 & ~x616 & ~x627 & ~x629 & ~x656 & ~x685;
assign c9298 =  x371 & ~x204 & ~x346 & ~x453 & ~x572 & ~x635;
assign c91 = ~x298 & ~x325 & ~x360 & ~x389 & ~x451 & ~x491 & ~x492 & ~x723 & ~x740 & ~x742;
assign c93 =  x127;
assign c95 = ~x26 & ~x39 & ~x51 & ~x56 & ~x85 & ~x86 & ~x94 & ~x124 & ~x125 & ~x126 & ~x127 & ~x155 & ~x182 & ~x183 & ~x196 & ~x210 & ~x225 & ~x238 & ~x304 & ~x367 & ~x447 & ~x477 & ~x501 & ~x528 & ~x536 & ~x595 & ~x614 & ~x623 & ~x640 & ~x676 & ~x721 & ~x757 & ~x781;
assign c97 =  x202;
assign c99 =  x568 & ~x16 & ~x51 & ~x114 & ~x139 & ~x146 & ~x177 & ~x368 & ~x371 & ~x618 & ~x718;
assign c911 =  x543 &  x571 &  x599 &  x600 & ~x12 & ~x54 & ~x146 & ~x444 & ~x447 & ~x709 & ~x756;
assign c913 =  x685 & ~x328 & ~x491;
assign c915 =  x240 &  x463 & ~x377 & ~x403 & ~x429 & ~x430 & ~x529;
assign c917 =  x149;
assign c919 =  x267 &  x463 & ~x270 & ~x271 & ~x326 & ~x327;
assign c921 =  x436 & ~x89 & ~x181 & ~x210 & ~x211 & ~x239 & ~x266 & ~x533;
assign c923 =  x266 &  x267 &  x268 & ~x26 & ~x54 & ~x99 & ~x114 & ~x129 & ~x150 & ~x155 & ~x156 & ~x183 & ~x334 & ~x365 & ~x430 & ~x431 & ~x441 & ~x459 & ~x535 & ~x542 & ~x543 & ~x639 & ~x699 & ~x749 & ~x752 & ~x766 & ~x775;
assign c925 =  x660 & ~x160 & ~x169 & ~x353 & ~x413 & ~x743;
assign c927 =  x405 & ~x12 & ~x70 & ~x74 & ~x123 & ~x129 & ~x139 & ~x282 & ~x283 & ~x284 & ~x306 & ~x395 & ~x409 & ~x555 & ~x562 & ~x621 & ~x714 & ~x716 & ~x723 & ~x726 & ~x738 & ~x742 & ~x744 & ~x773 & ~x779;
assign c929 = ~x15 & ~x76 & ~x149 & ~x168 & ~x310 & ~x348 & ~x377 & ~x378 & ~x429 & ~x430 & ~x433 & ~x457 & ~x459 & ~x468 & ~x487 & ~x500 & ~x588 & ~x690 & ~x758;
assign c931 =  x519 & ~x184 & ~x211 & ~x240 & ~x267 & ~x284 & ~x761;
assign c933 =  x191;
assign c935 = ~x39 & ~x156 & ~x183 & ~x184 & ~x185 & ~x204 & ~x212 & ~x221 & ~x239 & ~x240 & ~x252 & ~x267 & ~x268 & ~x582 & ~x639 & ~x677;
assign c937 =  x461 &  x516 &  x658;
assign c939 =  x266 &  x267 &  x268 & ~x2 & ~x10 & ~x33 & ~x51 & ~x54 & ~x104 & ~x141 & ~x146 & ~x155 & ~x182 & ~x201 & ~x249 & ~x280 & ~x377 & ~x430 & ~x486 & ~x533 & ~x561 & ~x674 & ~x705 & ~x720 & ~x727;
assign c941 = ~x0 & ~x10 & ~x23 & ~x24 & ~x32 & ~x55 & ~x66 & ~x68 & ~x73 & ~x82 & ~x104 & ~x106 & ~x110 & ~x119 & ~x122 & ~x127 & ~x128 & ~x129 & ~x132 & ~x135 & ~x140 & ~x155 & ~x171 & ~x183 & ~x193 & ~x199 & ~x201 & ~x203 & ~x211 & ~x221 & ~x222 & ~x230 & ~x232 & ~x239 & ~x256 & ~x267 & ~x278 & ~x310 & ~x362 & ~x363 & ~x390 & ~x394 & ~x418 & ~x421 & ~x508 & ~x541 & ~x584 & ~x593 & ~x594 & ~x597 & ~x609 & ~x614 & ~x622 & ~x648 & ~x666 & ~x670 & ~x681 & ~x697 & ~x698 & ~x704 & ~x719 & ~x725 & ~x747 & ~x752 & ~x761 & ~x766 & ~x769 & ~x774 & ~x777;
assign c943 =  x463 & ~x9 & ~x98 & ~x146 & ~x170 & ~x184 & ~x211 & ~x212 & ~x239 & ~x340 & ~x417 & ~x423 & ~x499 & ~x530 & ~x555 & ~x558 & ~x696 & ~x707 & ~x708 & ~x737;
assign c945 = ~x290 & ~x326 & ~x327 & ~x381;
assign c947 =  x567 &  x568;
assign c949 =  x632 & ~x182 & ~x430;
assign c951 =  x267 &  x268 &  x270 & ~x123 & ~x378 & ~x405 & ~x432 & ~x459 & ~x460 & ~x503 & ~x512 & ~x557;
assign c953 =  x513 &  x625 &  x654 & ~x11 & ~x40 & ~x51 & ~x66 & ~x137 & ~x146 & ~x202 & ~x279 & ~x640;
assign c955 =  x543 &  x571 &  x599 &  x627 & ~x7 & ~x39 & ~x84 & ~x109 & ~x142 & ~x176 & ~x277 & ~x283 & ~x311 & ~x312 & ~x642 & ~x743;
assign c957 =  x519 & ~x2 & ~x9 & ~x10 & ~x14 & ~x42 & ~x61 & ~x65 & ~x96 & ~x199 & ~x212 & ~x225 & ~x240 & ~x250 & ~x268 & ~x269 & ~x284 & ~x363 & ~x418 & ~x532 & ~x612 & ~x623 & ~x624 & ~x665 & ~x764;
assign c959 =  x267 &  x270 &  x318 & ~x64 & ~x77 & ~x157 & ~x183 & ~x202 & ~x338 & ~x377 & ~x378 & ~x389 & ~x405 & ~x444 & ~x453 & ~x503 & ~x553 & ~x615 & ~x640;
assign c961 =  x458 &  x512 & ~x48 & ~x74 & ~x83 & ~x85 & ~x92 & ~x129 & ~x135 & ~x363 & ~x445 & ~x477 & ~x616 & ~x645 & ~x718 & ~x719 & ~x749 & ~x781;
assign c963 =  x570 & ~x437;
assign c965 =  x622;
assign c967 =  x656 &  x658 &  x659 &  x660 &  x685 &  x686 & ~x429 & ~x503 & ~x557 & ~x561 & ~x614 & ~x726;
assign c969 =  x188 & ~x3 & ~x16 & ~x34 & ~x36 & ~x60 & ~x70 & ~x76 & ~x96 & ~x102 & ~x116 & ~x119 & ~x121 & ~x142 & ~x143 & ~x168 & ~x170 & ~x200 & ~x227 & ~x253 & ~x329 & ~x338 & ~x339 & ~x360 & ~x363 & ~x390 & ~x394 & ~x446 & ~x450 & ~x479 & ~x482 & ~x484 & ~x640 & ~x649 & ~x677 & ~x695 & ~x721 & ~x729 & ~x730 & ~x735 & ~x742 & ~x744;
assign c971 =  x375 &  x402 &  x403 &  x429 & ~x41 & ~x141 & ~x162 & ~x198 & ~x327 & ~x328 & ~x706 & ~x742 & ~x780;
assign c973 =  x406 & ~x45 & ~x46 & ~x84 & ~x114 & ~x117 & ~x138 & ~x225 & ~x298 & ~x299 & ~x325 & ~x326 & ~x327 & ~x353 & ~x357 & ~x360 & ~x362 & ~x444 & ~x663;
assign c975 =  x487 &  x543 &  x570;
assign c977 =  x296 & ~x86 & ~x111 & ~x161 & ~x181 & ~x182 & ~x209 & ~x210 & ~x237 & ~x238 & ~x304 & ~x531 & ~x570 & ~x617 & ~x783;
assign c979 =  x295 &  x435 &  x462 & ~x327 & ~x641 & ~x714 & ~x753;
assign c981 =  x260;
assign c983 =  x176;
assign c985 =  x621;
assign c987 =  x593;
assign c989 =  x487 &  x542 &  x570 & ~x780;
assign c991 =  x462 &  x517 & ~x3 & ~x5 & ~x18 & ~x33 & ~x70 & ~x98 & ~x116 & ~x121 & ~x193 & ~x198 & ~x201 & ~x312 & ~x402 & ~x418 & ~x451 & ~x452 & ~x457 & ~x469 & ~x524 & ~x551 & ~x553 & ~x565 & ~x608 & ~x708 & ~x759 & ~x761;
assign c993 = ~x55 & ~x84 & ~x115 & ~x118 & ~x298 & ~x326 & ~x327 & ~x352 & ~x353 & ~x364 & ~x382 & ~x415 & ~x506;
assign c995 =  x161;
assign c997 =  x602 &  x630 & ~x95 & ~x138 & ~x139 & ~x168 & ~x366 & ~x375 & ~x393 & ~x429 & ~x485 & ~x500 & ~x502 & ~x671 & ~x757 & ~x761;
assign c999 =  x244 &  x654 &  x655 & ~x67 & ~x77 & ~x85 & ~x94 & ~x97 & ~x138 & ~x227 & ~x440 & ~x560 & ~x584 & ~x698 & ~x699 & ~x705 & ~x708 & ~x723 & ~x743;
assign c9101 = ~x1 & ~x5 & ~x8 & ~x14 & ~x22 & ~x25 & ~x31 & ~x44 & ~x49 & ~x73 & ~x81 & ~x82 & ~x83 & ~x129 & ~x133 & ~x144 & ~x146 & ~x154 & ~x163 & ~x182 & ~x198 & ~x210 & ~x218 & ~x225 & ~x238 & ~x247 & ~x252 & ~x265 & ~x266 & ~x303 & ~x306 & ~x308 & ~x309 & ~x333 & ~x338 & ~x388 & ~x393 & ~x417 & ~x419 & ~x473 & ~x498 & ~x504 & ~x505 & ~x534 & ~x556 & ~x563 & ~x564 & ~x589 & ~x590 & ~x591 & ~x594 & ~x620 & ~x627 & ~x640 & ~x642 & ~x669 & ~x671 & ~x675 & ~x677 & ~x680 & ~x682 & ~x696 & ~x698 & ~x702 & ~x707 & ~x720 & ~x727 & ~x734 & ~x745 & ~x765 & ~x767 & ~x768 & ~x776 & ~x779;
assign c9103 =  x159 & ~x385;
assign c9105 =  x122;
assign c9107 =  x375 &  x376 &  x402 &  x403 &  x429 & ~x1 & ~x4 & ~x17 & ~x23 & ~x27 & ~x29 & ~x38 & ~x49 & ~x57 & ~x58 & ~x63 & ~x94 & ~x98 & ~x102 & ~x110 & ~x111 & ~x117 & ~x118 & ~x121 & ~x123 & ~x134 & ~x137 & ~x145 & ~x147 & ~x163 & ~x169 & ~x172 & ~x196 & ~x197 & ~x225 & ~x247 & ~x276 & ~x330 & ~x333 & ~x338 & ~x342 & ~x395 & ~x445 & ~x452 & ~x499 & ~x501 & ~x503 & ~x531 & ~x561 & ~x585 & ~x619 & ~x622 & ~x642 & ~x645 & ~x650 & ~x677 & ~x704 & ~x707 & ~x714 & ~x715 & ~x716 & ~x722 & ~x740 & ~x742 & ~x746 & ~x766 & ~x767 & ~x768 & ~x773 & ~x775 & ~x782;
assign c9109 =  x626 & ~x323 & ~x378 & ~x379;
assign c9111 =  x569 & ~x39 & ~x65 & ~x68 & ~x139 & ~x170 & ~x287 & ~x453 & ~x587 & ~x617 & ~x633 & ~x673 & ~x742 & ~x744 & ~x766;
assign c9113 =  x519 &  x523 &  x549;
assign c9115 =  x262 & ~x84 & ~x138 & ~x304 & ~x373 & ~x403 & ~x429 & ~x430 & ~x457 & ~x670;
assign c9117 =  x436 & ~x182 & ~x210 & ~x211 & ~x238 & ~x266 & ~x360 & ~x555 & ~x557 & ~x640 & ~x736 & ~x742;
assign c9119 =  x349 & ~x270 & ~x298 & ~x325;
assign c9121 =  x269 & ~x39 & ~x81 & ~x99 & ~x115 & ~x183 & ~x376 & ~x377 & ~x405 & ~x432 & ~x447 & ~x459 & ~x502 & ~x513 & ~x516;
assign c9123 =  x177 & ~x138;
assign c9125 =  x218 & ~x1 & ~x338 & ~x648 & ~x750;
assign c9127 =  x266 &  x267 &  x268 & ~x12 & ~x31 & ~x41 & ~x91 & ~x100 & ~x103 & ~x139 & ~x142 & ~x151 & ~x182 & ~x331 & ~x367 & ~x377 & ~x405 & ~x421 & ~x458 & ~x516 & ~x564 & ~x615 & ~x666 & ~x672 & ~x677 & ~x723 & ~x753 & ~x770 & ~x772 & ~x774;
assign c9129 =  x231 & ~x102 & ~x114 & ~x179 & ~x338 & ~x386 & ~x754;
assign c9131 = ~x8 & ~x21 & ~x27 & ~x40 & ~x93 & ~x95 & ~x113 & ~x114 & ~x115 & ~x117 & ~x120 & ~x124 & ~x183 & ~x211 & ~x212 & ~x239 & ~x240 & ~x267 & ~x295 & ~x388 & ~x539 & ~x554 & ~x556 & ~x559 & ~x583 & ~x610 & ~x670 & ~x769;
assign c9133 =  x129;
assign c9135 =  x269 &  x270 & ~x182 & ~x209 & ~x210 & ~x459;
assign c9137 =  x154 &  x462 & ~x4 & ~x73 & ~x194 & ~x312 & ~x371 & ~x415 & ~x536 & ~x748;
assign c9139 =  x266 &  x269 &  x270 & ~x85 & ~x249 & ~x377 & ~x378 & ~x405 & ~x424 & ~x433 & ~x514 & ~x584;
assign c9141 =  x322 & ~x263;
assign c9143 =  x268 &  x296 &  x463 & ~x209 & ~x327 & ~x357 & ~x766;
assign c9145 =  x567 & ~x691;
assign c9147 =  x299 &  x327 & ~x115 & ~x183 & ~x184 & ~x211 & ~x240 & ~x593 & ~x611 & ~x755;
assign c9149 =  x604 &  x605 & ~x5 & ~x136 & ~x246 & ~x298 & ~x326 & ~x327 & ~x716 & ~x717;
assign c9151 = ~x84 & ~x141 & ~x263 & ~x290 & ~x315 & ~x326 & ~x327 & ~x329 & ~x354 & ~x678 & ~x748;
assign c9153 =  x469 & ~x6 & ~x82 & ~x111 & ~x255 & ~x271 & ~x337 & ~x386 & ~x392 & ~x449 & ~x504 & ~x533 & ~x584 & ~x616 & ~x639 & ~x713 & ~x723 & ~x762 & ~x781;
assign c9155 =  x240 &  x270 & ~x22 & ~x36 & ~x39 & ~x53 & ~x82 & ~x84 & ~x140 & ~x362 & ~x364 & ~x377 & ~x378 & ~x389 & ~x394 & ~x430 & ~x433 & ~x448 & ~x458 & ~x459 & ~x477 & ~x486 & ~x496 & ~x542 & ~x609 & ~x621 & ~x677;
assign c9157 =  x241 &  x436 &  x463 & ~x30 & ~x33 & ~x37 & ~x40 & ~x60 & ~x123 & ~x162 & ~x252 & ~x304 & ~x310 & ~x350 & ~x370 & ~x371 & ~x401 & ~x402 & ~x444 & ~x476 & ~x510 & ~x531 & ~x553 & ~x612 & ~x728 & ~x729 & ~x782;
assign c9159 =  x442 & ~x312;
assign c9161 =  x541 &  x569 & ~x66 & ~x88 & ~x120 & ~x139 & ~x162 & ~x228 & ~x250 & ~x323 & ~x390 & ~x418 & ~x614 & ~x715 & ~x766;
assign c9163 =  x286;
assign c9167 =  x156 & ~x274 & ~x326 & ~x327;
assign c9169 =  x267 &  x517 & ~x225 & ~x402 & ~x427 & ~x429 & ~x639;
assign c9171 =  x204 &  x235 &  x240;
assign c9173 = ~x12 & ~x43 & ~x62 & ~x94 & ~x116 & ~x193 & ~x305 & ~x306 & ~x314 & ~x327 & ~x372 & ~x382 & ~x385 & ~x416 & ~x428 & ~x477 & ~x500 & ~x582 & ~x633 & ~x704 & ~x731 & ~x732 & ~x741 & ~x742 & ~x748 & ~x751 & ~x753;
assign c9175 =  x436 & ~x182 & ~x211 & ~x238 & ~x239 & ~x266;
assign c9177 =  x467 & ~x121 & ~x327 & ~x332 & ~x412 & ~x677 & ~x749 & ~x772;
assign c9179 =  x191;
assign c9181 =  x99;
assign c9183 =  x154 & ~x290 & ~x372 & ~x731;
assign c9185 =  x595;
assign c9187 = ~x174 & ~x182 & ~x210 & ~x211 & ~x238 & ~x239 & ~x266 & ~x393 & ~x554 & ~x780 & ~x783;
assign c9189 =  x542 &  x570 &  x598 & ~x12 & ~x17 & ~x36 & ~x65 & ~x84 & ~x115 & ~x137 & ~x141 & ~x142 & ~x150 & ~x169 & ~x194 & ~x196 & ~x223 & ~x225 & ~x226 & ~x227 & ~x257 & ~x276 & ~x285 & ~x334 & ~x338 & ~x361 & ~x421 & ~x526 & ~x556 & ~x557 & ~x584 & ~x593 & ~x614 & ~x637 & ~x677 & ~x723 & ~x732 & ~x735 & ~x742 & ~x743 & ~x744 & ~x747 & ~x752 & ~x764 & ~x781;
assign c9191 =  x159;
assign c9193 =  x238 & ~x30 & ~x39 & ~x55 & ~x62 & ~x66 & ~x78 & ~x104 & ~x107 & ~x124 & ~x133 & ~x162 & ~x179 & ~x195 & ~x254 & ~x333 & ~x334 & ~x338 & ~x349 & ~x351 & ~x360 & ~x365 & ~x378 & ~x379 & ~x389 & ~x407 & ~x446 & ~x449 & ~x461 & ~x474 & ~x500 & ~x503 & ~x514 & ~x530 & ~x536 & ~x585 & ~x645 & ~x667 & ~x672 & ~x733 & ~x750 & ~x751 & ~x756 & ~x776;
assign c9195 =  x241 & ~x14 & ~x130 & ~x352 & ~x379 & ~x380 & ~x408 & ~x482 & ~x484 & ~x756;
assign c9197 =  x229;
assign c9199 =  x174;
assign c9201 =  x568 &  x596 & ~x23 & ~x30 & ~x49 & ~x60 & ~x81 & ~x102 & ~x107 & ~x112 & ~x154 & ~x171 & ~x281 & ~x616 & ~x666 & ~x720 & ~x725;
assign c9203 =  x220;
assign c9205 =  x516 &  x626 & ~x429;
assign c9207 =  x240 &  x436 & ~x183 & ~x377 & ~x378 & ~x405 & ~x430 & ~x513;
assign c9209 =  x156 & ~x9 & ~x70 & ~x92 & ~x111 & ~x290 & ~x393 & ~x397 & ~x536 & ~x613 & ~x668 & ~x715 & ~x723 & ~x761 & ~x762 & ~x770;
assign c9211 = ~x13 & ~x341 & ~x408 & ~x437 & ~x499 & ~x689 & ~x742;
assign c9213 =  x267 &  x268 &  x270 & ~x38 & ~x73 & ~x126 & ~x198 & ~x255 & ~x304 & ~x378 & ~x433 & ~x752;
assign c9215 =  x402 & ~x182 & ~x210 & ~x266 & ~x294;
assign c9217 =  x432 &  x487 &  x542 & ~x2 & ~x4 & ~x21 & ~x48 & ~x65 & ~x84 & ~x85 & ~x112 & ~x138 & ~x168 & ~x169 & ~x170 & ~x198 & ~x200 & ~x203 & ~x283 & ~x391 & ~x421 & ~x474 & ~x477 & ~x587 & ~x613 & ~x614 & ~x615 & ~x616 & ~x640 & ~x671 & ~x694 & ~x699 & ~x722 & ~x730 & ~x749 & ~x772 & ~x774;
assign c9219 =  x231 &  x435 & ~x9 & ~x22 & ~x56 & ~x59 & ~x60 & ~x71 & ~x76 & ~x89 & ~x123 & ~x143 & ~x164 & ~x225 & ~x310 & ~x392 & ~x393 & ~x473 & ~x475 & ~x507 & ~x584 & ~x648 & ~x671 & ~x672 & ~x696 & ~x697 & ~x734 & ~x735;
assign c9221 = ~x12 & ~x42 & ~x108 & ~x182 & ~x210 & ~x211 & ~x223 & ~x238 & ~x266 & ~x565 & ~x646 & ~x717;
assign c9223 =  x458 &  x511;
assign c9225 = ~x54 & ~x93 & ~x95 & ~x137 & ~x156 & ~x183 & ~x211 & ~x212 & ~x224 & ~x239 & ~x240 & ~x251 & ~x266 & ~x267 & ~x285 & ~x323 & ~x422 & ~x451 & ~x477 & ~x701 & ~x741 & ~x776;
assign c9227 = ~x104 & ~x156 & ~x212 & ~x233 & ~x240 & ~x260 & ~x268 & ~x269 & ~x276 & ~x689 & ~x714 & ~x778;
assign c9229 = ~x92 & ~x153 & ~x182 & ~x375 & ~x401 & ~x402 & ~x403 & ~x404 & ~x429 & ~x453 & ~x457;
assign c9231 =  x570 &  x598 &  x599 &  x627 &  x628 & ~x443 & ~x476 & ~x530 & ~x615 & ~x726 & ~x736 & ~x737 & ~x744;
assign c9233 =  x176;
assign c9235 =  x257;
assign c9237 = ~x74 & ~x181 & ~x182 & ~x210 & ~x211 & ~x238 & ~x239 & ~x250 & ~x266 & ~x267 & ~x475 & ~x652;
assign c9239 =  x443;
assign c9241 =  x581 & ~x695;
assign c9243 =  x128;
assign c9245 = ~x5 & ~x40 & ~x62 & ~x68 & ~x74 & ~x81 & ~x97 & ~x114 & ~x126 & ~x128 & ~x138 & ~x151 & ~x284 & ~x323 & ~x359 & ~x362 & ~x377 & ~x378 & ~x385 & ~x387 & ~x405 & ~x418 & ~x427 & ~x429 & ~x430 & ~x446 & ~x458 & ~x503 & ~x526 & ~x569 & ~x589 & ~x622 & ~x623 & ~x642 & ~x662 & ~x671 & ~x702 & ~x757;
assign c9247 =  x461 &  x489 & ~x3 & ~x5 & ~x22 & ~x38 & ~x43 & ~x83 & ~x89 & ~x119 & ~x120 & ~x139 & ~x146 & ~x162 & ~x169 & ~x223 & ~x255 & ~x283 & ~x301 & ~x360 & ~x383 & ~x384 & ~x394 & ~x402 & ~x512 & ~x639 & ~x640 & ~x647 & ~x677 & ~x699 & ~x704 & ~x705 & ~x712 & ~x732 & ~x739 & ~x766 & ~x781;
assign c9249 =  x566;
assign c9251 =  x524 & ~x268 & ~x285;
assign c9253 =  x148;
assign c9255 =  x201;
assign c9257 =  x623;
assign c9259 =  x270 &  x271 &  x299 & ~x114 & ~x139 & ~x351 & ~x378 & ~x379 & ~x433 & ~x457 & ~x484 & ~x485;
assign c9261 =  x299 &  x626 & ~x377;
assign c9263 = ~x23 & ~x38 & ~x43 & ~x56 & ~x99 & ~x123 & ~x371 & ~x436 & ~x437 & ~x465 & ~x535 & ~x615 & ~x742;
assign c9265 =  x246 &  x299;
assign c9267 = ~x100 & ~x110 & ~x199 & ~x253 & ~x379 & ~x380 & ~x408 & ~x409 & ~x517 & ~x545 & ~x619 & ~x742;
assign c9269 =  x382 & ~x156 & ~x211 & ~x239 & ~x240 & ~x268 & ~x323 & ~x503;
assign c9271 =  x318 & ~x73 & ~x195 & ~x211 & ~x212 & ~x222 & ~x239 & ~x286 & ~x531 & ~x560 & ~x719;
assign c9273 =  x498;
assign c9275 =  x160;
assign c9277 =  x627 &  x655 &  x656 & ~x198 & ~x290 & ~x311 & ~x496 & ~x500 & ~x582 & ~x750;
assign c9279 =  x129;
assign c9281 =  x157 & ~x327;
assign c9283 = ~x130 & ~x280 & ~x360 & ~x406 & ~x407 & ~x408 & ~x435 & ~x436 & ~x446 & ~x464 & ~x478 & ~x491 & ~x517 & ~x777;
assign c9285 =  x266 &  x268 & ~x164 & ~x167 & ~x375 & ~x430 & ~x455 & ~x512;
assign c9287 =  x484 &  x511 & ~x7 & ~x21 & ~x715 & ~x716 & ~x745 & ~x780;
assign c9289 =  x128;
assign c9291 =  x318 & ~x184 & ~x206 & ~x212 & ~x240 & ~x558 & ~x718 & ~x725;
assign c9293 =  x240 &  x270 & ~x148 & ~x150 & ~x323 & ~x378 & ~x431 & ~x516 & ~x581 & ~x748;
assign c9295 =  x658 & ~x327 & ~x353 & ~x355 & ~x484;
assign c9297 =  x268 &  x269 & ~x14 & ~x85 & ~x105 & ~x121 & ~x156 & ~x182 & ~x191 & ~x378 & ~x405 & ~x456 & ~x489;
assign c9299 =  x241 & ~x1 & ~x2 & ~x32 & ~x34 & ~x53 & ~x68 & ~x76 & ~x77 & ~x93 & ~x121 & ~x129 & ~x133 & ~x138 & ~x143 & ~x161 & ~x175 & ~x200 & ~x202 & ~x221 & ~x227 & ~x278 & ~x306 & ~x311 & ~x331 & ~x338 & ~x350 & ~x377 & ~x390 & ~x392 & ~x394 & ~x395 & ~x403 & ~x405 & ~x419 & ~x421 & ~x430 & ~x443 & ~x457 & ~x468 & ~x472 & ~x484 & ~x498 & ~x505 & ~x513 & ~x529 & ~x534 & ~x541 & ~x564 & ~x586 & ~x589 & ~x595 & ~x607 & ~x636 & ~x665 & ~x668 & ~x677 & ~x690 & ~x699 & ~x706 & ~x725 & ~x730 & ~x747 & ~x752 & ~x753 & ~x758 & ~x772 & ~x775 & ~x777;

endmodule