module tm( x0,x1,x2,x3,x4,x5,x6,x7,x8,x9,x10,x11,x12,x13,x14,x15,x16,x17,x18,x19,x20,x21,x22,x23,x24,x25,x26,x27,x28,x29,x30,x31,x32,x33,x34,x35,x36,x37,x38,x39,x40,x41,x42,x43,x44,x45,x46,x47,x48,x49,x50,x51,x52,x53,x54,x55,x56,x57,x58,x59,x60,x61,x62,x63,x64,x65,x66,x67,x68,x69,x70,x71,x72,x73,x74,x75,x76,x77,x78,x79,x80,x81,x82,x83,x84,x85,x86,x87,x88,x89,x90,x91,x92,x93,x94,x95,c2218,c4384,c1456,c3279,c283,c2319,c4328,c11,c5266,c476,c0315,c5451,c3418,c2156,c5463,c1237,c0207,c449,c6376,c0250,c1434,c6462,c3164,c084,c3469,c197,c1402,c6131,c364,c5284,c159,c2101,c2341,c6357,c1348,c259,c0273,c597,c3424,c1119,c3131,c4102,c681,c1443,c6343,c4391,c6465,c1191,c3466,c6403,c4176,c4416,c5362,c0156,c5193,c41,c5239,c0254,c0391,c3440,c075,c359,c3307,c3276,c043,c1215,c0137,c2247,c4383,c6333,c2231,c4177,c652,c4403,c3364,c0189,c1483,c2144,c524,c0302,c0445,c4117,c627,c5145,c1480,c244,c4474,c2475,c6418,c4456,c1482,c4388,c0277,c2451,c40,c6456,c3481,c666,c6424,c357,c4168,c2143,c5338,c32,c5352,c3267,c6426,c5167,c0271,c1317,c189,c5408,c4441,c427,c4475,c1415,c1249,c594,c4346,c6275,c3121,c174,c6380,c5357,c3208,c0181,c3187,c0195,c2347,c6353,c1289,c5115,c2259,c0395,c3423,c2108,c3227,c3323,c4374,c224,c3356,c1374,c0496,c4207,c5448,c4135,c0176,c157,c4345,c6249,c1241,c599,c0414,c3295,c6409,c486,c421,c1417,c2492,c1438,c2373,c689,c2121,c214,c0438,c3454,c2169,c269,c5331,c2103,c0152,c0386,c4387,c1171,c4364,c240,c2489,c3247,c6197,c0209,c1104,c2130,c2278,c4439,c528,c5429,c5403,c217,c684,c2327,c1189,c2459,c6435,c2482,c0121,c459,c0347,c3216,c5120,c5443,c6388,c5340,c6180,c676,c4309,c6490,c0263,c2336,c3464,c6305,c1256,c1280,c2316,c5102,c130,c365,c4128,c1158,c6201,c3403,c6208,c0381,c3475,c034,c6276,c4186,c072,c3292,c4376,c2412,c6261,c1496,c0472,c1295,c4165,c4216,c116,c1433,c479,c010,c0451,c3490,c3492,c1377,c6367,c6284,c1184,c0359,c5492,c464,c05,c1216,c1305,c260,c6302,c2281,c2481,c590,c0336,c3431,c2265,c5333,c2348,c4213,c3488,c2390,c1488,c4212,c6105,c3405,c5150,c6262,c2282,c5327,c6245,c0420,c4464,c216,c0487,c2163,c426,c4339,c1275,c5351,c2225,c6464,c1476,c0394,c461,c5416,c1197,c5217,c0404,c0477,c6369,c0368,c4283,c0217,c5202,c5414,c4118,c44,c4162,c2193,c5142,c4420,c1153,c0133,c2126,c4243,c122,c2277,c6159,c0313,c4264,c1164,c319,c6419,c0427,c0411,c1174,c2355,c3495,c6303,c451,c2398,c1234,c0310,c6117,c4362,c3102,c312,c2456,c39,c046,c3209,c5111,c5179,c0272,c566,c5330,c2138,c237,c4438,c266,c0214,c280,c3174,c331,c195,c4154,c026,c0291,c0125,c4113,c1327,c114,c3184,c0282,c0443,c1293,c4326,c3413,c428,c4200,c5222,c20,c0498,c1458,c2215,c0247,c142,c016,c168,c1245,c2164,c3463,c5267,c5364,c4467,c0415,c1328,c1462,c62,c0396,c4378,c6452,c0374,c612,c5358,c0371,c1387,c1395,c329,c5227,c012,c4394,c5295,c4231,c4191,c6347,c1366,c5130,c5458,c1351,c1236,c6454,c6103,c4144,c6281,c3368,c1141,c08,c258,c0481,c581,c6216,c2109,c2363,c4494,c2228,c4385,c5436,c63,c1440,c3123,c6188,c3260,c2279,c6277,c5268,c057,c1435,c52,c2137,c0122,c0325,c053,c2146,c3433,c0304,c0266,c1226,c0312,c415,c0221,c3139,c0348,c480,c6162,c6172,c1465,c0229,c2212,c4256,c2467,c0154,c2186,c3313,c5380,c5204,c432,c1136,c3176,c465,c565,c6332,c5312,c412,c123,c6113,c6315,c1178,c5322,c6268,c6161,c2180,c616,c6423,c3272,c3372,c0377,c1350,c4120,c5140,c6483,c0105,c553,c552,c330,c2350,c1130,c4305,c5353,c2424,c5418,c0252,c1331,c1263,c6398,c4214,c450,c6115,c560,c664,c6241,c3225,c336,c0466,c4194,c173,c0455,c0465,c376,c5164,c6346,c1375,c6381,c2132,c4413,c5134,c3180,c3248,c3218,c5343,c0123,c5132,c4227,c4334,c013,c3265,c2113,c494,c6273,c5275,c3402,c4298,c5444,c0492,c3115,c5305,c3204,c6179,c054,c1269,c4315,c6106,c6441,c323,c2375,c4238,c24,c1355,c523,c0106,c1436,c2127,c2148,c4111,c1262,c5214,c2176,c0190,c5394,c4314,c5170,c521,c1365,c649,c2188,c516,c6167,c0168,c0429,c3330,c6470,c4291,c170,c6393,c3261,c5240,c425,c4304,c6233,c1105,c6210,c0488,c483,c574,c00,c5432,c674,c568,c4344,c4255,c6394,c3312,c0180,c513,c2365,c5470,c6484,c4386,c4481,c6256,c1492,c5430,c2266,c4142,c5194,c2294,c2498,c6363,c4114,c5439,c10,c4197,c4311,c5241,c2241,c325,c378,c0403,c272,c3274,c5456,c0167,c080,c186,c1151,c4461,c3280,c592,c0295,c1279,c5196,c5223,c5431,c6207,c6431,c4262,c2414,c0144,c0224,c5246,c4218,c4410,c1475,c6242,c1219,c1329,c3494,c6174,c1270,c5162,c3322,c5411,c3191,c1131,c2426,c6360,c3378,c3443,c422,c5231,c4297,c587,c6330,c619,c6119,c356,c4427,c6355,c6127,c1335,c225,c3314,c3430,c5300,c6163,c0241,c2151,c1144,c3203,c6327,c6450,c0286,c1179,c6126,c0148,c0283,c4280,c3181,c0215,c179,c2449,c1165,c5288,c5390,c6324,c2383,c5291,c424,c5387,c1401,c6364,c6183,c2116,c352,c4104,c4300,c530,c079,c4215,c6181,c436,c6336,c2447,c082,c1251,c3285,c1315,c0475,c0183,c2486,c1123,c1453,c2323,c349,c3388,c2484,c411,c1425,c2381,c6266,c178,c648,c6459,c4463,c1420,c2464,c5110,c326,c3242,c0275,c1344,c060,c5230,c6402,c077,c4101,c3256,c5149,c2395,c2255,c1134,c3379,c3381,c635,c6202,c110,c4308,c0300,c5206,c50,c5335,c6236,c0288,c6143,c2441,c0177,c1232,c548,c2312,c3376,c1391,c4437,c0467,c0170,c4204,c1252,c0324,c2290,c3214,c4247,c1286,c4358,c341,c3141,c5449,c0355,c2499,c4396,c5491,c6265,c437,c3459,c1261,c5348,c431,c3344,c5211,c096,c2222,c3207,c6267,c270,c6123,c099,c6250,c1356,c6466,c6135,c6153,c4320,c4155,c6102,c5171,c1324,c5392,c3396,c158,c4381,c642,c6370,c6294,c5349,c218,c5498,c5106,c4312,c067,c2457,c2182,c4159,c0108,c0473,c1410,c6495,c4459,c5114,c2275,c2309,c5283,c3155,c6178,c1211,c2334,c1460,c6144,c0428,c6325,c044,c48,c6352,c5341,c3107,c1116,c5158,c3186,c3485,c4217,c3293,c5185,c1129,c366,c1148,c247,c2253,c6209,c193,c5128,c1446,c6175,c1137,c4445,c4125,c617,c0284,c0196,c0184,c6218,c3194,c514,c5313,c6482,c2269,c5481,c3199,c2234,c580,c2159,c2402,c321,c6366,c3136,c268,c6390,c1294,c5437,c0200,c0151,c4251,c1468,c3104,c3110,c5494,c0204,c2133,c3220,c3238,c5285,c6270,c0193,c6391,c3226,c2224,c696,c036,c6192,c1362,c5455,c5127,c1203,c2288,c290,c3254,c3346,c5379,c4136,c030,c6491,c5163,c5224,c256,c5365,c2468,c0150,c13,c4476,c1147,c5397,c5286,c539,c598,c0188,c236,c389,c257,c5287,c4143,c3221,c467,c3168,c0212,c370,c4103,c3437,c1162,c673,c1310,c4100,c398,c6227,c6194,c1322,c5182,c3268,c43,c342,c3338,c1448,c228,c3306,c5125,c5405,c1228,c1429,c0157,c6311,c274,c5235,c6182,c1347,c5465,c049,c6316,c4237,c0328,c5190,c6372,c2419,c45,c3389,c0236,c2487,c2439,c2251,c2232,c3200,c2488,c5374,c0439,c2473,c399,c5303,c299,c2173,c4257,c1495,c2476,c0318,c6361,c49,c4121,c670,c4436,c5329,c5176,c2140,c2364,c1132,c4306,c6314,c0128,c4190,c3320,c6479,c5178,c1484,c583,c5401,c6164,c6252,c440,c6328,c5460,c5271,c6436,c4355,c3117,c6322,c5136,c2134,c1100,c0131,c5304,c6239,c4115,c0301,c0116,c1384,c6146,c3382,c4409,c0424,c0425,c555,c3112,c3253,c3193,c1299,c6453,c5367,c3415,c0491,c0162,c1115,c255,c3229,c384,c6351,c1209,c6138,c0103,c315,c1161,c0419,c6255,c0142,c613,c324,c2118,c5175,c2387,c1244,c3395,c2142,c1250,c5301,c6382,c143,c320,c4296,c3124,c6350,c6358,c1212,c2293,c078,c3219,c1430,c4284,c6300,c5438,c4465,c546,c1332,c0384,c2434,c2285,c061,c6331,c0238,c2371,c6282,c611,c6226,c4370,c190,c2466,c022,c2129,c3441,c289,c1175,c675,c2401,c0448,c4453,c0191,c1399,c3277,c5213,c493,c54,c6341,c5315,c698,c1491,c3233,c3215,c1357,c3497,c64,c6145,c1173,c3188,c2359,c2368,c374,c3491,c278,c0174,c3499,c1303,c2149,c1308,c6246,c1302,c6433,c6445,c176,c5412,c61,c4484,c2252,c0141,c690,c0308,c6354,c2314,c3406,c6203,c1349,c3334,c2154,c285,c5219,c695,c2430,c4367,c4492,c434,c4278,c0178,c117,c2393,c2254,c1113,c671,c444,c543,c6299,c6147,c4199,c372,c5378,c5148,c3310,c6116,c6170,c0290,c1222,c1330,c2287,c4321,c1264,c6272,c4405,c144,c1321,c6280,c4130,c232,c2406,c4246,c2208,c6118,c3245,c5477,c1202,c0124,c1360,c361,c5314,c5233,c4303,c6287,c5197,c4158,c5104,c2260,c1152,c418,c1477,c297,c3134,c251,c3154,c4323,c148,c2425,c2298,c0192,c0149,c3428,c4139,c1254,c2472,c4225,c3409,c0342,c2442,c1230,c0129,c4286,c1287,c37,c4127,c59,c5425,c1160,c588,c5489,c4285,c1213,c2302,c4351,c537,c056,c068,c3133,c6321,c0232,c5346,c468,c161,c6240,c267,c4249,c6100,c1421,c5113,c6359,c6235,c6438,c6389,c496,c2239,c2403,c1479,c131,c0486,c0219,c0337,c1112,c151,c2306,c2227,c4274,c6121,c1273,c5342,c498,c5375,c088,c2493,c4397,c1193,c1390,c4489,c4477,c139,c2382,c2354,c5318,c5141,c2335,c3489,c4195,c1288,c1283,c5126,c2305,c1157,c5325,c5203,c1354,c687,c0421,c5165,c3429,c6230,c6399,c4234,c0338,c6422,c2410,c3347,c3471,c5187,c2195,c5272,c3365,c339,c3342,c0331,c1314,c2307,c0226,c5199,c4172,c0213,c6476,c1411,c595,c090,c3175,c571,c413,c0454,c60,c125,c3426,c469,c2453,c252,c0405,c1200,c6442,c4380,c1296,c6478,c4174,c2171,c2202,c1472,c2158,c0433,c4147,c6263,c4279,c2150,c3398,c0228,c1442,c4341,c4471,c083,c0109,c348,c6395,c4166,c661,c511,c287,c2361,c1325,c2471,c4288,c6186,c4210,c4330,c2386,c276,c6406,c5336,c050,c5143,c1383,c0161,c5131,c213,c692,c5399,c6386,c0485,c4377,c2374,c4479,c313,c2396,c554,c5105,c334,c025,c1466,c3425,c0317,c0471,c2211,c0499,c2276,c2105,c2157,c2199,c697,c2345,c1214,c1386,c0298,c4140,c2460,c1255,c1208,c296,c0289,c1370,c3445,c2183,c294,c0119,c3359,c5221,c2233,c2479,c570,c3325,c5493,c2450,c3150,c4472,c1290,c6134,c628,c6413,c0440,c6337,c0197,c3457,c5415,c165,c1372,c3317,c0101,c1110,c095,c2376,c1334,c4209,c3192,c5434,c6415,c0389,c383,c5228,c646,c6140,c1463,c2284,c242,c169,c6253,c1169,c5157,c6283,c5251,c2220,c4411,c430,c4106,c4123,c532,c6248,c0199,c4451,c30,c166,c371,c4379,c0497,c0171,c3303,c2192,c0255,c3182,c3282,c6404,c5116,c5151,c097,c3370,c0307,c2417,c3452,c027,c453,c4372,c065,c1247,c286,c5388,c037,c2470,c0450,c18,c4244,c3240,c6259,c076,c4448,c087,c1451,c098,c196,c4241,c3422,c1124,c5361,c6379,c4219,c2198,c2184,c0139,c4265,c3416,c6198,c3239,c0278,c0446,c1457,c0117,c5317,c2324,c4193,c0436,c3472,c0385,c4307,c4301,c2117,c145,c017,c485,c0360,c2203,c5243,c5201,c4281,c6461,c0269,c1300,c4175,c249,c6231,c4417,c381,c3270,c6411,c435,c593,c654,c5135,c1341,c510,c5297,c2342,c3408,c1364,c6247,c3266,c4167,c3250,c092,c229,c1437,c3177,c149,c3479,c2311,c243,c1337,c1282,c5270,c1405,c4222,c577,c0132,c2461,c3449,c433,c6169,c6225,c0120,c5417,c5218,c3399,c446,c5245,c1265,c223,c0285,c350,c0281,c0235,c4156,c1346,c4310,c4496,c4112,c0380,c3284,c452,c0303,c073,c2427,c3183,c167,c3332,c3394,c3255,c0367,c3249,c5409,c6362,c1109,c3190,c4208,c2268,c564,c0185,c1367,c3390,c3417,c5410,c2349,c5382,c118,c693,c6443,c6497,c0457,c5488,c1146,c6342,c3252,c4418,c2185,c0469,c6449,c3251,c3421,c5319,c5253,c6458,c2445,c3162,c1225,c0182,c484,c4149,c660,c3296,c4248,c442,c1336,c2339,c5328,c3167,c2370,c5247,c1318,c4498,c3108,c517,c0169,c4319,c153,c630,c672,c1187,c4455,c0340,c6487,c2422,c6173,c0135,c6200,c355,c5472,c12,c2111,c2207,c6166,c1181,c4354,c345,c5280,c09,c5469,c4452,c2165,c6345,c066,c2358,c2145,c3271,c3473,c134,c2310,c0412,c36,c495,c6238,c343,c113,c691,c3196,c4357,c0393,c1388,c3223,c3432,c3327,c3290,c5289,c6489,c6295,c569,c4119,c6499,c4485,c2344,c1101,c4317,c3434,c3205,c0268,c3166,c1248,c4151,c5166,c0339,c3468,c2340,c344,c2286,c4371,c5107,c4415,c3264,c6187,c2352,c2139,c160,c5236,c3447,c191,c6177,c6368,c1156,c625,c1159,c1276,c0251,c128,c3318,c314,c579,c221,c121,c219,c4169,c4270,c563,c147,c5370,c5407,c3297,c417,c5153,c2346,c6396,c4495,c5138,c35,c65,c140,c4421,c3358,c6122,c4449,c1127,c475,c621,c0246,c0260,c0493,c6112,c4134,c4224,c3197,c3329,c273,c1185,c2299,c182,c1176,c3142,c2409,c0240,c2343,c3122,c3137,c3460,c0453,c4340,c1389,c2333,c589,c0245,c1418,c062,c3170,c0130,c5413,c024,c3369,c4375,c31,c6110,c6141,c429,c5433,c443,c3210,c6191,c2496,c2178,c0444,c1102,c1235,c6421,c041,c3206,c3278,c497,c5363,c5344,c56,c610,c33,c2214,c0476,c1373,c386,c5316,c254,c2431,c6237,c4373,c0230,c1339,c2120,c3480,c1285,c4268,c5497,c1217,c1284,c6290,c1108,c0358,c4348,c0356,c0410,c2378,c6356,c141,c680,c5323,c0198,c6214,c3385,c439,c638,c499,c5256,c5292,c0265,c2321,c6292,c5447,c3300,c3158,c6229,c1313,c3147,c3152,c2240,c368,c0458,c0326,c0293,c1419,c1447,c0470,c230,c231,c318,c385,c4343,c0323,c392,c490,c3185,c6109,c5377,c3289,c0392,c2196,c2274,c3326,c6335,c1393,c3410,c1229,c6288,c1201,c2315,c3333,c1198,c5459,c2366,c5306,c5356,c5147,c538,c6444,c3397,c5321,c6124,c6468,c363,c215,c4327,c388,c1371,c2166,c3331,c6171,c2235,c5281,c0480,c0407,c0408,c0459,c0296,c3273,c639,c5208,c0249,c1199,c3435,c4356,c1307,c6348,c653,c1240,c0482,c66,c5212,c5391,c3224,c2107,c6271,c0343,c3298,c1459,c3484,c2429,c4254,c4189,c4361,c395,c0175,c3383,c488,c5129,c6212,c6492,c1172,c2125,c6204,c0113,c048,c0341,c2112,c332,c1196,c3138,c1103,c4316,c4457,c6414,c5468,c2440,c5478,c120,c322,c4302,c086,c4399,c0346,c3476,c5103,c3125,c1206,c1277,c561,c5252,c4450,c1218,c4276,c2261,c622,c4163,c1297,c0126,c3305,c5294,c1381,c1396,c5216,c2152,c380,c3393,c53,c111,c3262,c1398,c0210,c2491,c4109,c4153,c4202,c4447,c353,c559,c0306,c3140,c375,c591,c6446,c4182,c67,c633,c1382,c3106,c2304,c6494,c180,c4423,c5453,c2175,c4178,c5172,c6349,c064,c1227,c4110,c1271,c4490,c460,c1470,c2174,c6279,c6317,c5100,c549,c311,c3316,c150,c2465,c3145,c4407,c5452,c3287,c4185,c2320,c2313,c5473,c69,c5400,c058,c0430,c0329,c2435,c651,c1121,c3478,c6384,c2219,c5248,c4338,c6365,c1278,c5276,c5257,c2191,c0305,c647,c1192,c0211,c558,c4480,c5154,c4325,c0431,c618,c2380,c5479,c6339,c3160,c3116,c1133,c2421,c414,c463,c4360,c4295,c5471,c3228,c4138,c6114,c641,c6157,c445,c3257,c0158,c3113,c615,c678,c5188,c2405,c0146,c233,c572,c46,c0463,c2474,c5195,c2197,c6108,c3201,c6467,c4294,c0160,c4313,c4425,c5440,c0299,c1450,c584,c6234,c5137,c6264,c1469,c5480,c2135,c3127,c3353,c337,c4491,c410,c5101,c6304,c279,c6430,c0287,c632,c3458,c1311,c6155,c0294,c187,c631,c3496,c1243,c2436,c1340,c6326,c2438,c2204,c4180,c1306,c5326,c2318,c2454,c011,c481,c3241,c1407,c6460,c4318,c5298,c456,c1353,c5355,c0248,c1489,c0242,c146,c2292,c3308,c5457,c3235,c3148,c2325,c2416,c1224,c1428,c4446,c6374,c6477,c3109,c0179,c4273,c4369,c3444,c6392,c0353,c462,c4290,c5234,c250,c2168,c2236,c5112,c2177,c5238,c624,c3319,c0399,c4271,c3450,c4122,c373,c2124,c3341,c16,c2128,c0390,c4430,c4466,c2469,c2205,c6463,c1342,c4266,c6306,c6329,c5389,c5189,c310,c0166,c261,c3178,c4272,c582,c1239,c57,c1454,c039,c0461,c4382,c0322,c3367,c263,c4198,c2338,c3165,c2248,c4133,c1163,c58,c2495,c2155,c1126,c133,c2362,c0376,c2179,c5226,c585,c5146,c6133,c0409,c557,c6301,c4499,c5200,c1464,c0143,c6160,c3132,c3455,c2200,c0239,c4366,c0205,c4275,c5359,c0460,c2263,c0434,c298,c5464,c3301,c6309,c1257,c575,c3135,c4332,c23,c5435,c4221,c1326,c2418,c6168,c3234,c1445,c4292,c5250,c0201,c4390,c2160,c6260,c5174,c1485,c6416,c1467,c0435,c519,c2141,c4164,c2170,c0227,c2331,c5302,c0165,c175,c019,c0173,c1397,c2245,c3439,c4299,c644,c3151,c3483,c4245,c38,c4392,c1140,c253,c5168,c059,c527,c6385,c6107,c0261,c1149,c5308,c2329,c5395,c0397,c3340,c0456,c0417,c6137,c070,c1168,c6220,c4203,c2229,c416,c0363,c4470,c623,c4365,c6205,c4230,c3453,c1481,c4460,c1135,c6420,c5232,c4287,c1368,c346,c3401,c3302,c6312,c2201,c6432,c47,c5160,c6439,c4250,c6298,c0332,c2303,c4431,c535,c1343,c3391,c6196,c6308,c1292,c0474,c1408,c2322,c1404,c0321,c379,c5446,c2360,c1155,c2480,c293,c4414,c6148,c3392,c6498,c3195,c0233,c0118,c562,c2190,c265,c264,c1427,c0413,c1210,c2432,c3349,c27,c0364,c1345,c1452,c4395,c0237,c2328,c2478,c474,c2272,c19,c387,c1180,c5180,c6111,c1274,c5366,c0140,c4205,c1403,c4486,c0104,c5152,c4259,c3474,c659,c5274,c1441,c5265,c4433,c0206,c0344,c2385,c071,c2262,c1128,c2477,c3336,c2249,c4422,c2448,c5161,c281,c0267,c2490,c2291,c4160,c3232,c3387,c643,c4132,c3477,c1183,c282,c2119,c0276,c1166,c5173,c2379,c3363,c020,c1272,c4404,c5487,c6323,c2408,c423,c2404,c668,c51,c154,c5445,c2106,c5386,c5474,c0452,c1423,c0382,c1167,c3169,c3411,c15,c5225,c172,c5385,c4488,c5123,c1392,c6440,c227,c1499,c369,c6184,c0253,c3328,c2483,c0334,c045,c645,c1486,c6193,c2332,c6149,c089,c351,c4408,c472,c5406,c6104,c4260,c038,c473,c686,c4226,c1106,c5441,c0379,c127,c1281,c2308,c2301,c4232,c0100,c4150,c4398,c135,c5320,c2147,c5108,c1107,c2356,c3153,c3442,c2391,c6221,c5279,c0110,c0388,c0270,c0490,c3461,c4235,c3362,c4468,c1471,c5205,c6156,c394,c5484,c2407,c5402,c6130,c0297,c1145,c210,c3172,c0280,c4482,c518,c2455,c0483,c192,c2242,c0234,c4342,c2413,c4483,c466,c5262,c4293,c1188,c2131,c1439,c4401,c5119,c358,c3436,c5192,c5475,c550,c1494,c470,c5290,c4393,c5209,c198,c2246,c3118,c0292,c0354,c0114,c1358,c3366,c2102,c578,c573,c3236,c0222,c5169,c2216,c4469,c512,c3246,c5124,c6258,c4129,c0279,c2115,c4406,c0423,c1413,c4236,c4242,c3361,c2161,c0441,c688,c07,c636,c0112,c3337,c284,c0187,c4108,c6320,c3128,c248,c162,c4454,c291,c34,c4335,c5354,c0163,c3163,c491,c5269,c5450,c0373,c667,c6101,c5499,c1186,c2428,c1143,c2400,c382,c3486,c3335,c4184,c1246,c2420,c4233,c5261,c547,c6378,c1238,c5220,c6412,c3237,c295,c4349,c3161,c4324,c454,c032,c5263,c040,c390,c6244,c6448,c2372,c6434,c6120,c2213,c156,c1182,c1426,c4337,c245,c3159,c55,c2458,c1412,c3243,c2221,c1268,c3130,c6286,c25,c3294,c262,c5181,c2433,c420,c2377,c0400,c3448,c1320,c4173,c2122,c4444,c5118,c699,c4400,c2443,c3304,c1207,c3173,c3355,c5144,c238,c3380,c5466,c6455,c5454,c4363,c360,c0274,c4336,c5121,c0398,c0449,c637,c2388,c3189,c3100,c1385,c5372,c6189,c3149,c3230,c5244,c5309,c6257,c6291,c2389,c2497,c6338,c2485,c0345,c3120,c4240,c665,c6222,c6425,c2267,c212,c4269,c2437,c5381,c397,c1194,c1154,c1432,c1233,c3202,c0468,c1253,c22,c4282,c0426,c5184,c525,c14,c2367,c6152,c3493,c6293,c3384,c2296,c3386,c3309,c063,c0145,c0370,c3288,c4440,c2300,c2494,c477,c4211,c5155,c6488,c0375,c28,c029,c3414,c6475,c1400,c3258,c4105,c5368,c06,c277,c6334,c0262,c1120,c626,c0418,c0115,c4196,c4267,c534,c1298,c5278,c0361,c3498,c3269,c5419,c0220,c01,c3373,c6451,c5260,c028,c1312,c5422,c4131,c335,c2415,c1378,c6340,c5337,c3101,c447,c0351,c2446,c3179,c0327,c3311,c0107,c6469,c4261,c5310,c5133,c4141,c3482,c4116,c5476,c1376,c5249,c6377,c4171,c5198,c5393,c669,c136,c656,c541,c5122,c393,c663,c4148,c5307,c5207,c396,c4424,c0357,c5183,c655,c3291,c6471,c288,c5311,c1490,c2206,c441,c3315,c2271,c0216,c1220,c0489,c3420,c2189,c2462,c2230,c3299,c03,c155,c6307,c6158,c2104,c2256,c3286,c682,c1424,c3462,c2237,c3129,c1142,c0134,c047,c3321,c522,c586,c4181,c551,c6310,c6232,c657,c2351,c4493,c5242,c6485,c2172,c1291,c2114,c4458,c033,c2330,c6481,c3371,c4107,c5421,c6486,c6136,c0111,c4497,c338,c018,c5485,c2411,c4402,c6480,c2223,c0350,c3103,c6428,c5186,c1117,c2295,c1444,c124,c222,c6151,c2187,c3263,c3213,c6150,c3111,c4389,c0223,c4353,c6387,c091,c6285,c051,c340,c4426,c0147,c5273,c1416,c0416,c6269,c023,c1461,c4228,c2369,c4192,c4329,c1150,c4277,c4443,c3357,c081,c1493,c126,c1369,c074,c567,c5293,c2384,c5324,c5264,c2264,c0365,c6297,c163,c6213,c194,c482,c596,c5404,c5467,c2238,c015,c5210,c679,c2210,c68,c362,c1319,c3275,c0442,c0256,c0225,c2153,c3211,c6319,c6375,c0330,c0218,c0422,c6224,c2280,c177,c2444,c6289,c3212,c6427,c1352,c455,c5462,c0464,c5347,c171,c1478,c556,c4161,c5373,c2209,c3281,c526,c4223,c1361,c0202,c2452,c4478,c0136,c1497,c2392,c0335,c1259,c5442,c377,c152,c6493,c3350,c1309,c1122,c6129,c0203,c0264,c1498,c199,c0257,c2162,c0462,c2243,c0437,c1449,c3375,c536,c3352,c29,c6243,c0172,c6437,c5427,c042,c5277,c2217,c6278,c2136,c6228,c1170,c478,c4170,c115,c055,c2297,c3283,c094,c02,c2273,c0479,c4434,c5424,c3427,c3222,c6128,c3404,c6383,c1316,c1422,c4289,c1304,c5334,c6142,c5258,c241,c0378,c2357,c3114,c5376,c271,c0362,c529,c6496,c683,c184,c1190,c4145,c4183,c3146,c1333,c6154,c6400,c2399,c662,c629,c1359,c5482,c0447,c4412,c4368,c1231,c2423,c1258,c0406,c2337,c6457,c0159,c5360,c035,c138,c3244,c4229,c6199,c5109,c0316,c093,c576,c0186,c0258,c5229,c1177,c4220,c6125,c6407,c0320,c4206,c3419,c4352,c471,c5339,c545,c6132,c3231,c0314,c542,c129,c3171,c275,c2257,c6408,c0372,c650,c6401,c4252,c4263,c4462,c3217,c5396,c3198,c1338,c0369,c2283,c052,c0138,c246,c4428,c4435,c6417,c2226,c1242,c489,c620,c42,c1394,c164,c458,c6185,c0208,c3324,c3105,c1221,c3119,c5332,c1455,c5215,c3360,c1301,c438,c211,c4126,c0352,c2100,c3259,c119,c5428,c658,c3126,c6195,c3143,c0231,c6139,c4188,c4124,c317,c6274,c185,c6313,c2110,c3157,c021,c3438,c1114,c04,c2326,c1138,c3374,c6206,c1118,c5117,c6405,c0333,c4152,c4350,c0155,c6410,c614,c487,c677,c2194,c6223,c4333,c4146,c1363,c085,c448,c2250,c685,c220,c2394,c2167,c367,c0319,c391,c5139,c0387,c2181,c069,c5191,c0127,c6472,c5369,c5423,c1414,c4487,c0311,c0244,c354,c6215,c0309,c6219,c0243,c0402,c6474,c515,c1260,c0494,c492,c4429,c0153,c5461,c4322,c239,c234,c5490,c112,c5259,c6296,c014,c5345,c5384,c5299,c2244,c0194,c1379,c1125,c2289,c1473,c188,c1487,c3465,c0102,c5156,c1267,c6344,c3467,c333,c2397,c6371,c3412,c328,c2463,c4347,c316,c3343,c5426,c5282,c3377,c183,c5496,c4179,c3156,c3456,c3487,c4359,c2123,c5177,c0432,c6211,c0478,c4201,c640,c4258,c347,c0401,c0349,c0383,c235,c4419,c5350,c292,c520,c6254,c6447,c0366,c031,c1205,c1204,c1139,c3144,c3354,c3345,c6190,c1223,c3470,c5237,c6217,c1266,c1474,c5254,c5495,c137,c0164,c544,c1380,c6397,c2258,c0484,c0259,c4331,c4442,c3348,c531,c6373,c226,c533,c457,c6165,c5398,c4473,c634,c1111,c3407,c6318,c17,c181,c4432,c3446,c5383,c4253,c3451,c1431,c6176,c5420,c132,c21,c0495,c1323,c4137,c5486,c5483,c3351,c5296,c419,c5159,c26,c694,c6473,c1409,c4157,c5371,c2270,c3400,c3339,c4187,c540,c1406,c327,c6429,c2353,c6251,c2317,c4239,c1195,c5255 );

input x0;
input x1;
input x2;
input x3;
input x4;
input x5;
input x6;
input x7;
input x8;
input x9;
input x10;
input x11;
input x12;
input x13;
input x14;
input x15;
input x16;
input x17;
input x18;
input x19;
input x20;
input x21;
input x22;
input x23;
input x24;
input x25;
input x26;
input x27;
input x28;
input x29;
input x30;
input x31;
input x32;
input x33;
input x34;
input x35;
input x36;
input x37;
input x38;
input x39;
input x40;
input x41;
input x42;
input x43;
input x44;
input x45;
input x46;
input x47;
input x48;
input x49;
input x50;
input x51;
input x52;
input x53;
input x54;
input x55;
input x56;
input x57;
input x58;
input x59;
input x60;
input x61;
input x62;
input x63;
input x64;
input x65;
input x66;
input x67;
input x68;
input x69;
input x70;
input x71;
input x72;
input x73;
input x74;
input x75;
input x76;
input x77;
input x78;
input x79;
input x80;
input x81;
input x82;
input x83;
input x84;
input x85;
input x86;
input x87;
input x88;
input x89;
input x90;
input x91;
input x92;
input x93;
input x94;
input x95;
output c2218;
output c4384;
output c1456;
output c3279;
output c283;
output c2319;
output c4328;
output c11;
output c5266;
output c476;
output c0315;
output c5451;
output c3418;
output c2156;
output c5463;
output c1237;
output c0207;
output c449;
output c6376;
output c0250;
output c1434;
output c6462;
output c3164;
output c084;
output c3469;
output c197;
output c1402;
output c6131;
output c364;
output c5284;
output c159;
output c2101;
output c2341;
output c6357;
output c1348;
output c259;
output c0273;
output c597;
output c3424;
output c1119;
output c3131;
output c4102;
output c681;
output c1443;
output c6343;
output c4391;
output c6465;
output c1191;
output c3466;
output c6403;
output c4176;
output c4416;
output c5362;
output c0156;
output c5193;
output c41;
output c5239;
output c0254;
output c0391;
output c3440;
output c075;
output c359;
output c3307;
output c3276;
output c043;
output c1215;
output c0137;
output c2247;
output c4383;
output c6333;
output c2231;
output c4177;
output c652;
output c4403;
output c3364;
output c0189;
output c1483;
output c2144;
output c524;
output c0302;
output c0445;
output c4117;
output c627;
output c5145;
output c1480;
output c244;
output c4474;
output c2475;
output c6418;
output c4456;
output c1482;
output c4388;
output c0277;
output c2451;
output c40;
output c6456;
output c3481;
output c666;
output c6424;
output c357;
output c4168;
output c2143;
output c5338;
output c32;
output c5352;
output c3267;
output c6426;
output c5167;
output c0271;
output c1317;
output c189;
output c5408;
output c4441;
output c427;
output c4475;
output c1415;
output c1249;
output c594;
output c4346;
output c6275;
output c3121;
output c174;
output c6380;
output c5357;
output c3208;
output c0181;
output c3187;
output c0195;
output c2347;
output c6353;
output c1289;
output c5115;
output c2259;
output c0395;
output c3423;
output c2108;
output c3227;
output c3323;
output c4374;
output c224;
output c3356;
output c1374;
output c0496;
output c4207;
output c5448;
output c4135;
output c0176;
output c157;
output c4345;
output c6249;
output c1241;
output c599;
output c0414;
output c3295;
output c6409;
output c486;
output c421;
output c1417;
output c2492;
output c1438;
output c2373;
output c689;
output c2121;
output c214;
output c0438;
output c3454;
output c2169;
output c269;
output c5331;
output c2103;
output c0152;
output c0386;
output c4387;
output c1171;
output c4364;
output c240;
output c2489;
output c3247;
output c6197;
output c0209;
output c1104;
output c2130;
output c2278;
output c4439;
output c528;
output c5429;
output c5403;
output c217;
output c684;
output c2327;
output c1189;
output c2459;
output c6435;
output c2482;
output c0121;
output c459;
output c0347;
output c3216;
output c5120;
output c5443;
output c6388;
output c5340;
output c6180;
output c676;
output c4309;
output c6490;
output c0263;
output c2336;
output c3464;
output c6305;
output c1256;
output c1280;
output c2316;
output c5102;
output c130;
output c365;
output c4128;
output c1158;
output c6201;
output c3403;
output c6208;
output c0381;
output c3475;
output c034;
output c6276;
output c4186;
output c072;
output c3292;
output c4376;
output c2412;
output c6261;
output c1496;
output c0472;
output c1295;
output c4165;
output c4216;
output c116;
output c1433;
output c479;
output c010;
output c0451;
output c3490;
output c3492;
output c1377;
output c6367;
output c6284;
output c1184;
output c0359;
output c5492;
output c464;
output c05;
output c1216;
output c1305;
output c260;
output c6302;
output c2281;
output c2481;
output c590;
output c0336;
output c3431;
output c2265;
output c5333;
output c2348;
output c4213;
output c3488;
output c2390;
output c1488;
output c4212;
output c6105;
output c3405;
output c5150;
output c6262;
output c2282;
output c5327;
output c6245;
output c0420;
output c4464;
output c216;
output c0487;
output c2163;
output c426;
output c4339;
output c1275;
output c5351;
output c2225;
output c6464;
output c1476;
output c0394;
output c461;
output c5416;
output c1197;
output c5217;
output c0404;
output c0477;
output c6369;
output c0368;
output c4283;
output c0217;
output c5202;
output c5414;
output c4118;
output c44;
output c4162;
output c2193;
output c5142;
output c4420;
output c1153;
output c0133;
output c2126;
output c4243;
output c122;
output c2277;
output c6159;
output c0313;
output c4264;
output c1164;
output c319;
output c6419;
output c0427;
output c0411;
output c1174;
output c2355;
output c3495;
output c6303;
output c451;
output c2398;
output c1234;
output c0310;
output c6117;
output c4362;
output c3102;
output c312;
output c2456;
output c39;
output c046;
output c3209;
output c5111;
output c5179;
output c0272;
output c566;
output c5330;
output c2138;
output c237;
output c4438;
output c266;
output c0214;
output c280;
output c3174;
output c331;
output c195;
output c4154;
output c026;
output c0291;
output c0125;
output c4113;
output c1327;
output c114;
output c3184;
output c0282;
output c0443;
output c1293;
output c4326;
output c3413;
output c428;
output c4200;
output c5222;
output c20;
output c0498;
output c1458;
output c2215;
output c0247;
output c142;
output c016;
output c168;
output c1245;
output c2164;
output c3463;
output c5267;
output c5364;
output c4467;
output c0415;
output c1328;
output c1462;
output c62;
output c0396;
output c4378;
output c6452;
output c0374;
output c612;
output c5358;
output c0371;
output c1387;
output c1395;
output c329;
output c5227;
output c012;
output c4394;
output c5295;
output c4231;
output c4191;
output c6347;
output c1366;
output c5130;
output c5458;
output c1351;
output c1236;
output c6454;
output c6103;
output c4144;
output c6281;
output c3368;
output c1141;
output c08;
output c258;
output c0481;
output c581;
output c6216;
output c2109;
output c2363;
output c4494;
output c2228;
output c4385;
output c5436;
output c63;
output c1440;
output c3123;
output c6188;
output c3260;
output c2279;
output c6277;
output c5268;
output c057;
output c1435;
output c52;
output c2137;
output c0122;
output c0325;
output c053;
output c2146;
output c3433;
output c0304;
output c0266;
output c1226;
output c0312;
output c415;
output c0221;
output c3139;
output c0348;
output c480;
output c6162;
output c6172;
output c1465;
output c0229;
output c2212;
output c4256;
output c2467;
output c0154;
output c2186;
output c3313;
output c5380;
output c5204;
output c432;
output c1136;
output c3176;
output c465;
output c565;
output c6332;
output c5312;
output c412;
output c123;
output c6113;
output c6315;
output c1178;
output c5322;
output c6268;
output c6161;
output c2180;
output c616;
output c6423;
output c3272;
output c3372;
output c0377;
output c1350;
output c4120;
output c5140;
output c6483;
output c0105;
output c553;
output c552;
output c330;
output c2350;
output c1130;
output c4305;
output c5353;
output c2424;
output c5418;
output c0252;
output c1331;
output c1263;
output c6398;
output c4214;
output c450;
output c6115;
output c560;
output c664;
output c6241;
output c3225;
output c336;
output c0466;
output c4194;
output c173;
output c0455;
output c0465;
output c376;
output c5164;
output c6346;
output c1375;
output c6381;
output c2132;
output c4413;
output c5134;
output c3180;
output c3248;
output c3218;
output c5343;
output c0123;
output c5132;
output c4227;
output c4334;
output c013;
output c3265;
output c2113;
output c494;
output c6273;
output c5275;
output c3402;
output c4298;
output c5444;
output c0492;
output c3115;
output c5305;
output c3204;
output c6179;
output c054;
output c1269;
output c4315;
output c6106;
output c6441;
output c323;
output c2375;
output c4238;
output c24;
output c1355;
output c523;
output c0106;
output c1436;
output c2127;
output c2148;
output c4111;
output c1262;
output c5214;
output c2176;
output c0190;
output c5394;
output c4314;
output c5170;
output c521;
output c1365;
output c649;
output c2188;
output c516;
output c6167;
output c0168;
output c0429;
output c3330;
output c6470;
output c4291;
output c170;
output c6393;
output c3261;
output c5240;
output c425;
output c4304;
output c6233;
output c1105;
output c6210;
output c0488;
output c483;
output c574;
output c00;
output c5432;
output c674;
output c568;
output c4344;
output c4255;
output c6394;
output c3312;
output c0180;
output c513;
output c2365;
output c5470;
output c6484;
output c4386;
output c4481;
output c6256;
output c1492;
output c5430;
output c2266;
output c4142;
output c5194;
output c2294;
output c2498;
output c6363;
output c4114;
output c5439;
output c10;
output c4197;
output c4311;
output c5241;
output c2241;
output c325;
output c378;
output c0403;
output c272;
output c3274;
output c5456;
output c0167;
output c080;
output c186;
output c1151;
output c4461;
output c3280;
output c592;
output c0295;
output c1279;
output c5196;
output c5223;
output c5431;
output c6207;
output c6431;
output c4262;
output c2414;
output c0144;
output c0224;
output c5246;
output c4218;
output c4410;
output c1475;
output c6242;
output c1219;
output c1329;
output c3494;
output c6174;
output c1270;
output c5162;
output c3322;
output c5411;
output c3191;
output c1131;
output c2426;
output c6360;
output c3378;
output c3443;
output c422;
output c5231;
output c4297;
output c587;
output c6330;
output c619;
output c6119;
output c356;
output c4427;
output c6355;
output c6127;
output c1335;
output c225;
output c3314;
output c3430;
output c5300;
output c6163;
output c0241;
output c2151;
output c1144;
output c3203;
output c6327;
output c6450;
output c0286;
output c1179;
output c6126;
output c0148;
output c0283;
output c4280;
output c3181;
output c0215;
output c179;
output c2449;
output c1165;
output c5288;
output c5390;
output c6324;
output c2383;
output c5291;
output c424;
output c5387;
output c1401;
output c6364;
output c6183;
output c2116;
output c352;
output c4104;
output c4300;
output c530;
output c079;
output c4215;
output c6181;
output c436;
output c6336;
output c2447;
output c082;
output c1251;
output c3285;
output c1315;
output c0475;
output c0183;
output c2486;
output c1123;
output c1453;
output c2323;
output c349;
output c3388;
output c2484;
output c411;
output c1425;
output c2381;
output c6266;
output c178;
output c648;
output c6459;
output c4463;
output c1420;
output c2464;
output c5110;
output c326;
output c3242;
output c0275;
output c1344;
output c060;
output c5230;
output c6402;
output c077;
output c4101;
output c3256;
output c5149;
output c2395;
output c2255;
output c1134;
output c3379;
output c3381;
output c635;
output c6202;
output c110;
output c4308;
output c0300;
output c5206;
output c50;
output c5335;
output c6236;
output c0288;
output c6143;
output c2441;
output c0177;
output c1232;
output c548;
output c2312;
output c3376;
output c1391;
output c4437;
output c0467;
output c0170;
output c4204;
output c1252;
output c0324;
output c2290;
output c3214;
output c4247;
output c1286;
output c4358;
output c341;
output c3141;
output c5449;
output c0355;
output c2499;
output c4396;
output c5491;
output c6265;
output c437;
output c3459;
output c1261;
output c5348;
output c431;
output c3344;
output c5211;
output c096;
output c2222;
output c3207;
output c6267;
output c270;
output c6123;
output c099;
output c6250;
output c1356;
output c6466;
output c6135;
output c6153;
output c4320;
output c4155;
output c6102;
output c5171;
output c1324;
output c5392;
output c3396;
output c158;
output c4381;
output c642;
output c6370;
output c6294;
output c5349;
output c218;
output c5498;
output c5106;
output c4312;
output c067;
output c2457;
output c2182;
output c4159;
output c0108;
output c0473;
output c1410;
output c6495;
output c4459;
output c5114;
output c2275;
output c2309;
output c5283;
output c3155;
output c6178;
output c1211;
output c2334;
output c1460;
output c6144;
output c0428;
output c6325;
output c044;
output c48;
output c6352;
output c5341;
output c3107;
output c1116;
output c5158;
output c3186;
output c3485;
output c4217;
output c3293;
output c5185;
output c1129;
output c366;
output c1148;
output c247;
output c2253;
output c6209;
output c193;
output c5128;
output c1446;
output c6175;
output c1137;
output c4445;
output c4125;
output c617;
output c0284;
output c0196;
output c0184;
output c6218;
output c3194;
output c514;
output c5313;
output c6482;
output c2269;
output c5481;
output c3199;
output c2234;
output c580;
output c2159;
output c2402;
output c321;
output c6366;
output c3136;
output c268;
output c6390;
output c1294;
output c5437;
output c0200;
output c0151;
output c4251;
output c1468;
output c3104;
output c3110;
output c5494;
output c0204;
output c2133;
output c3220;
output c3238;
output c5285;
output c6270;
output c0193;
output c6391;
output c3226;
output c2224;
output c696;
output c036;
output c6192;
output c1362;
output c5455;
output c5127;
output c1203;
output c2288;
output c290;
output c3254;
output c3346;
output c5379;
output c4136;
output c030;
output c6491;
output c5163;
output c5224;
output c256;
output c5365;
output c2468;
output c0150;
output c13;
output c4476;
output c1147;
output c5397;
output c5286;
output c539;
output c598;
output c0188;
output c236;
output c389;
output c257;
output c5287;
output c4143;
output c3221;
output c467;
output c3168;
output c0212;
output c370;
output c4103;
output c3437;
output c1162;
output c673;
output c1310;
output c4100;
output c398;
output c6227;
output c6194;
output c1322;
output c5182;
output c3268;
output c43;
output c342;
output c3338;
output c1448;
output c228;
output c3306;
output c5125;
output c5405;
output c1228;
output c1429;
output c0157;
output c6311;
output c274;
output c5235;
output c6182;
output c1347;
output c5465;
output c049;
output c6316;
output c4237;
output c0328;
output c5190;
output c6372;
output c2419;
output c45;
output c3389;
output c0236;
output c2487;
output c2439;
output c2251;
output c2232;
output c3200;
output c2488;
output c5374;
output c0439;
output c2473;
output c399;
output c5303;
output c299;
output c2173;
output c4257;
output c1495;
output c2476;
output c0318;
output c6361;
output c49;
output c4121;
output c670;
output c4436;
output c5329;
output c5176;
output c2140;
output c2364;
output c1132;
output c4306;
output c6314;
output c0128;
output c4190;
output c3320;
output c6479;
output c5178;
output c1484;
output c583;
output c5401;
output c6164;
output c6252;
output c440;
output c6328;
output c5460;
output c5271;
output c6436;
output c4355;
output c3117;
output c6322;
output c5136;
output c2134;
output c1100;
output c0131;
output c5304;
output c6239;
output c4115;
output c0301;
output c0116;
output c1384;
output c6146;
output c3382;
output c4409;
output c0424;
output c0425;
output c555;
output c3112;
output c3253;
output c3193;
output c1299;
output c6453;
output c5367;
output c3415;
output c0491;
output c0162;
output c1115;
output c255;
output c3229;
output c384;
output c6351;
output c1209;
output c6138;
output c0103;
output c315;
output c1161;
output c0419;
output c6255;
output c0142;
output c613;
output c324;
output c2118;
output c5175;
output c2387;
output c1244;
output c3395;
output c2142;
output c1250;
output c5301;
output c6382;
output c143;
output c320;
output c4296;
output c3124;
output c6350;
output c6358;
output c1212;
output c2293;
output c078;
output c3219;
output c1430;
output c4284;
output c6300;
output c5438;
output c4465;
output c546;
output c1332;
output c0384;
output c2434;
output c2285;
output c061;
output c6331;
output c0238;
output c2371;
output c6282;
output c611;
output c6226;
output c4370;
output c190;
output c2466;
output c022;
output c2129;
output c3441;
output c289;
output c1175;
output c675;
output c2401;
output c0448;
output c4453;
output c0191;
output c1399;
output c3277;
output c5213;
output c493;
output c54;
output c6341;
output c5315;
output c698;
output c1491;
output c3233;
output c3215;
output c1357;
output c3497;
output c64;
output c6145;
output c1173;
output c3188;
output c2359;
output c2368;
output c374;
output c3491;
output c278;
output c0174;
output c3499;
output c1303;
output c2149;
output c1308;
output c6246;
output c1302;
output c6433;
output c6445;
output c176;
output c5412;
output c61;
output c4484;
output c2252;
output c0141;
output c690;
output c0308;
output c6354;
output c2314;
output c3406;
output c6203;
output c1349;
output c3334;
output c2154;
output c285;
output c5219;
output c695;
output c2430;
output c4367;
output c4492;
output c434;
output c4278;
output c0178;
output c117;
output c2393;
output c2254;
output c1113;
output c671;
output c444;
output c543;
output c6299;
output c6147;
output c4199;
output c372;
output c5378;
output c5148;
output c3310;
output c6116;
output c6170;
output c0290;
output c1222;
output c1330;
output c2287;
output c4321;
output c1264;
output c6272;
output c4405;
output c144;
output c1321;
output c6280;
output c4130;
output c232;
output c2406;
output c4246;
output c2208;
output c6118;
output c3245;
output c5477;
output c1202;
output c0124;
output c1360;
output c361;
output c5314;
output c5233;
output c4303;
output c6287;
output c5197;
output c4158;
output c5104;
output c2260;
output c1152;
output c418;
output c1477;
output c297;
output c3134;
output c251;
output c3154;
output c4323;
output c148;
output c2425;
output c2298;
output c0192;
output c0149;
output c3428;
output c4139;
output c1254;
output c2472;
output c4225;
output c3409;
output c0342;
output c2442;
output c1230;
output c0129;
output c4286;
output c1287;
output c37;
output c4127;
output c59;
output c5425;
output c1160;
output c588;
output c5489;
output c4285;
output c1213;
output c2302;
output c4351;
output c537;
output c056;
output c068;
output c3133;
output c6321;
output c0232;
output c5346;
output c468;
output c161;
output c6240;
output c267;
output c4249;
output c6100;
output c1421;
output c5113;
output c6359;
output c6235;
output c6438;
output c6389;
output c496;
output c2239;
output c2403;
output c1479;
output c131;
output c0486;
output c0219;
output c0337;
output c1112;
output c151;
output c2306;
output c2227;
output c4274;
output c6121;
output c1273;
output c5342;
output c498;
output c5375;
output c088;
output c2493;
output c4397;
output c1193;
output c1390;
output c4489;
output c4477;
output c139;
output c2382;
output c2354;
output c5318;
output c5141;
output c2335;
output c3489;
output c4195;
output c1288;
output c1283;
output c5126;
output c2305;
output c1157;
output c5325;
output c5203;
output c1354;
output c687;
output c0421;
output c5165;
output c3429;
output c6230;
output c6399;
output c4234;
output c0338;
output c6422;
output c2410;
output c3347;
output c3471;
output c5187;
output c2195;
output c5272;
output c3365;
output c339;
output c3342;
output c0331;
output c1314;
output c2307;
output c0226;
output c5199;
output c4172;
output c0213;
output c6476;
output c1411;
output c595;
output c090;
output c3175;
output c571;
output c413;
output c0454;
output c60;
output c125;
output c3426;
output c469;
output c2453;
output c252;
output c0405;
output c1200;
output c6442;
output c4380;
output c1296;
output c6478;
output c4174;
output c2171;
output c2202;
output c1472;
output c2158;
output c0433;
output c4147;
output c6263;
output c4279;
output c2150;
output c3398;
output c0228;
output c1442;
output c4341;
output c4471;
output c083;
output c0109;
output c348;
output c6395;
output c4166;
output c661;
output c511;
output c287;
output c2361;
output c1325;
output c2471;
output c4288;
output c6186;
output c4210;
output c4330;
output c2386;
output c276;
output c6406;
output c5336;
output c050;
output c5143;
output c1383;
output c0161;
output c5131;
output c213;
output c692;
output c5399;
output c6386;
output c0485;
output c4377;
output c2374;
output c4479;
output c313;
output c2396;
output c554;
output c5105;
output c334;
output c025;
output c1466;
output c3425;
output c0317;
output c0471;
output c2211;
output c0499;
output c2276;
output c2105;
output c2157;
output c2199;
output c697;
output c2345;
output c1214;
output c1386;
output c0298;
output c4140;
output c2460;
output c1255;
output c1208;
output c296;
output c0289;
output c1370;
output c3445;
output c2183;
output c294;
output c0119;
output c3359;
output c5221;
output c2233;
output c2479;
output c570;
output c3325;
output c5493;
output c2450;
output c3150;
output c4472;
output c1290;
output c6134;
output c628;
output c6413;
output c0440;
output c6337;
output c0197;
output c3457;
output c5415;
output c165;
output c1372;
output c3317;
output c0101;
output c1110;
output c095;
output c2376;
output c1334;
output c4209;
output c3192;
output c5434;
output c6415;
output c0389;
output c383;
output c5228;
output c646;
output c6140;
output c1463;
output c2284;
output c242;
output c169;
output c6253;
output c1169;
output c5157;
output c6283;
output c5251;
output c2220;
output c4411;
output c430;
output c4106;
output c4123;
output c532;
output c6248;
output c0199;
output c4451;
output c30;
output c166;
output c371;
output c4379;
output c0497;
output c0171;
output c3303;
output c2192;
output c0255;
output c3182;
output c3282;
output c6404;
output c5116;
output c5151;
output c097;
output c3370;
output c0307;
output c2417;
output c3452;
output c027;
output c453;
output c4372;
output c065;
output c1247;
output c286;
output c5388;
output c037;
output c2470;
output c0450;
output c18;
output c4244;
output c3240;
output c6259;
output c076;
output c4448;
output c087;
output c1451;
output c098;
output c196;
output c4241;
output c3422;
output c1124;
output c5361;
output c6379;
output c4219;
output c2198;
output c2184;
output c0139;
output c4265;
output c3416;
output c6198;
output c3239;
output c0278;
output c0446;
output c1457;
output c0117;
output c5317;
output c2324;
output c4193;
output c0436;
output c3472;
output c0385;
output c4307;
output c4301;
output c2117;
output c145;
output c017;
output c485;
output c0360;
output c2203;
output c5243;
output c5201;
output c4281;
output c6461;
output c0269;
output c1300;
output c4175;
output c249;
output c6231;
output c4417;
output c381;
output c3270;
output c6411;
output c435;
output c593;
output c654;
output c5135;
output c1341;
output c510;
output c5297;
output c2342;
output c3408;
output c1364;
output c6247;
output c3266;
output c4167;
output c3250;
output c092;
output c229;
output c1437;
output c3177;
output c149;
output c3479;
output c2311;
output c243;
output c1337;
output c1282;
output c5270;
output c1405;
output c4222;
output c577;
output c0132;
output c2461;
output c3449;
output c433;
output c6169;
output c6225;
output c0120;
output c5417;
output c5218;
output c3399;
output c446;
output c5245;
output c1265;
output c223;
output c0285;
output c350;
output c0281;
output c0235;
output c4156;
output c1346;
output c4310;
output c4496;
output c4112;
output c0380;
output c3284;
output c452;
output c0303;
output c073;
output c2427;
output c3183;
output c167;
output c3332;
output c3394;
output c3255;
output c0367;
output c3249;
output c5409;
output c6362;
output c1109;
output c3190;
output c4208;
output c2268;
output c564;
output c0185;
output c1367;
output c3390;
output c3417;
output c5410;
output c2349;
output c5382;
output c118;
output c693;
output c6443;
output c6497;
output c0457;
output c5488;
output c1146;
output c6342;
output c3252;
output c4418;
output c2185;
output c0469;
output c6449;
output c3251;
output c3421;
output c5319;
output c5253;
output c6458;
output c2445;
output c3162;
output c1225;
output c0182;
output c484;
output c4149;
output c660;
output c3296;
output c4248;
output c442;
output c1336;
output c2339;
output c5328;
output c3167;
output c2370;
output c5247;
output c1318;
output c4498;
output c3108;
output c517;
output c0169;
output c4319;
output c153;
output c630;
output c672;
output c1187;
output c4455;
output c0340;
output c6487;
output c2422;
output c6173;
output c0135;
output c6200;
output c355;
output c5472;
output c12;
output c2111;
output c2207;
output c6166;
output c1181;
output c4354;
output c345;
output c5280;
output c09;
output c5469;
output c4452;
output c2165;
output c6345;
output c066;
output c2358;
output c2145;
output c3271;
output c3473;
output c134;
output c2310;
output c0412;
output c36;
output c495;
output c6238;
output c343;
output c113;
output c691;
output c3196;
output c4357;
output c0393;
output c1388;
output c3223;
output c3432;
output c3327;
output c3290;
output c5289;
output c6489;
output c6295;
output c569;
output c4119;
output c6499;
output c4485;
output c2344;
output c1101;
output c4317;
output c3434;
output c3205;
output c0268;
output c3166;
output c1248;
output c4151;
output c5166;
output c0339;
output c3468;
output c2340;
output c344;
output c2286;
output c4371;
output c5107;
output c4415;
output c3264;
output c6187;
output c2352;
output c2139;
output c160;
output c5236;
output c3447;
output c191;
output c6177;
output c6368;
output c1156;
output c625;
output c1159;
output c1276;
output c0251;
output c128;
output c3318;
output c314;
output c579;
output c221;
output c121;
output c219;
output c4169;
output c4270;
output c563;
output c147;
output c5370;
output c5407;
output c3297;
output c417;
output c5153;
output c2346;
output c6396;
output c4495;
output c5138;
output c35;
output c65;
output c140;
output c4421;
output c3358;
output c6122;
output c4449;
output c1127;
output c475;
output c621;
output c0246;
output c0260;
output c0493;
output c6112;
output c4134;
output c4224;
output c3197;
output c3329;
output c273;
output c1185;
output c2299;
output c182;
output c1176;
output c3142;
output c2409;
output c0240;
output c2343;
output c3122;
output c3137;
output c3460;
output c0453;
output c4340;
output c1389;
output c2333;
output c589;
output c0245;
output c1418;
output c062;
output c3170;
output c0130;
output c5413;
output c024;
output c3369;
output c4375;
output c31;
output c6110;
output c6141;
output c429;
output c5433;
output c443;
output c3210;
output c6191;
output c2496;
output c2178;
output c0444;
output c1102;
output c1235;
output c6421;
output c041;
output c3206;
output c3278;
output c497;
output c5363;
output c5344;
output c56;
output c610;
output c33;
output c2214;
output c0476;
output c1373;
output c386;
output c5316;
output c254;
output c2431;
output c6237;
output c4373;
output c0230;
output c1339;
output c2120;
output c3480;
output c1285;
output c4268;
output c5497;
output c1217;
output c1284;
output c6290;
output c1108;
output c0358;
output c4348;
output c0356;
output c0410;
output c2378;
output c6356;
output c141;
output c680;
output c5323;
output c0198;
output c6214;
output c3385;
output c439;
output c638;
output c499;
output c5256;
output c5292;
output c0265;
output c2321;
output c6292;
output c5447;
output c3300;
output c3158;
output c6229;
output c1313;
output c3147;
output c3152;
output c2240;
output c368;
output c0458;
output c0326;
output c0293;
output c1419;
output c1447;
output c0470;
output c230;
output c231;
output c318;
output c385;
output c4343;
output c0323;
output c392;
output c490;
output c3185;
output c6109;
output c5377;
output c3289;
output c0392;
output c2196;
output c2274;
output c3326;
output c6335;
output c1393;
output c3410;
output c1229;
output c6288;
output c1201;
output c2315;
output c3333;
output c1198;
output c5459;
output c2366;
output c5306;
output c5356;
output c5147;
output c538;
output c6444;
output c3397;
output c5321;
output c6124;
output c6468;
output c363;
output c215;
output c4327;
output c388;
output c1371;
output c2166;
output c3331;
output c6171;
output c2235;
output c5281;
output c0480;
output c0407;
output c0408;
output c0459;
output c0296;
output c3273;
output c639;
output c5208;
output c0249;
output c1199;
output c3435;
output c4356;
output c1307;
output c6348;
output c653;
output c1240;
output c0482;
output c66;
output c5212;
output c5391;
output c3224;
output c2107;
output c6271;
output c0343;
output c3298;
output c1459;
output c3484;
output c2429;
output c4254;
output c4189;
output c4361;
output c395;
output c0175;
output c3383;
output c488;
output c5129;
output c6212;
output c6492;
output c1172;
output c2125;
output c6204;
output c0113;
output c048;
output c0341;
output c2112;
output c332;
output c1196;
output c3138;
output c1103;
output c4316;
output c4457;
output c6414;
output c5468;
output c2440;
output c5478;
output c120;
output c322;
output c4302;
output c086;
output c4399;
output c0346;
output c3476;
output c5103;
output c3125;
output c1206;
output c1277;
output c561;
output c5252;
output c4450;
output c1218;
output c4276;
output c2261;
output c622;
output c4163;
output c1297;
output c0126;
output c3305;
output c5294;
output c1381;
output c1396;
output c5216;
output c2152;
output c380;
output c3393;
output c53;
output c111;
output c3262;
output c1398;
output c0210;
output c2491;
output c4109;
output c4153;
output c4202;
output c4447;
output c353;
output c559;
output c0306;
output c3140;
output c375;
output c591;
output c6446;
output c4182;
output c67;
output c633;
output c1382;
output c3106;
output c2304;
output c6494;
output c180;
output c4423;
output c5453;
output c2175;
output c4178;
output c5172;
output c6349;
output c064;
output c1227;
output c4110;
output c1271;
output c4490;
output c460;
output c1470;
output c2174;
output c6279;
output c6317;
output c5100;
output c549;
output c311;
output c3316;
output c150;
output c2465;
output c3145;
output c4407;
output c5452;
output c3287;
output c4185;
output c2320;
output c2313;
output c5473;
output c69;
output c5400;
output c058;
output c0430;
output c0329;
output c2435;
output c651;
output c1121;
output c3478;
output c6384;
output c2219;
output c5248;
output c4338;
output c6365;
output c1278;
output c5276;
output c5257;
output c2191;
output c0305;
output c647;
output c1192;
output c0211;
output c558;
output c4480;
output c5154;
output c4325;
output c0431;
output c618;
output c2380;
output c5479;
output c6339;
output c3160;
output c3116;
output c1133;
output c2421;
output c414;
output c463;
output c4360;
output c4295;
output c5471;
output c3228;
output c4138;
output c6114;
output c641;
output c6157;
output c445;
output c3257;
output c0158;
output c3113;
output c615;
output c678;
output c5188;
output c2405;
output c0146;
output c233;
output c572;
output c46;
output c0463;
output c2474;
output c5195;
output c2197;
output c6108;
output c3201;
output c6467;
output c4294;
output c0160;
output c4313;
output c4425;
output c5440;
output c0299;
output c1450;
output c584;
output c6234;
output c5137;
output c6264;
output c1469;
output c5480;
output c2135;
output c3127;
output c3353;
output c337;
output c4491;
output c410;
output c5101;
output c6304;
output c279;
output c6430;
output c0287;
output c632;
output c3458;
output c1311;
output c6155;
output c0294;
output c187;
output c631;
output c3496;
output c1243;
output c2436;
output c1340;
output c6326;
output c2438;
output c2204;
output c4180;
output c1306;
output c5326;
output c2318;
output c2454;
output c011;
output c481;
output c3241;
output c1407;
output c6460;
output c4318;
output c5298;
output c456;
output c1353;
output c5355;
output c0248;
output c1489;
output c0242;
output c146;
output c2292;
output c3308;
output c5457;
output c3235;
output c3148;
output c2325;
output c2416;
output c1224;
output c1428;
output c4446;
output c6374;
output c6477;
output c3109;
output c0179;
output c4273;
output c4369;
output c3444;
output c6392;
output c0353;
output c462;
output c4290;
output c5234;
output c250;
output c2168;
output c2236;
output c5112;
output c2177;
output c5238;
output c624;
output c3319;
output c0399;
output c4271;
output c3450;
output c4122;
output c373;
output c2124;
output c3341;
output c16;
output c2128;
output c0390;
output c4430;
output c4466;
output c2469;
output c2205;
output c6463;
output c1342;
output c4266;
output c6306;
output c6329;
output c5389;
output c5189;
output c310;
output c0166;
output c261;
output c3178;
output c4272;
output c582;
output c1239;
output c57;
output c1454;
output c039;
output c0461;
output c4382;
output c0322;
output c3367;
output c263;
output c4198;
output c2338;
output c3165;
output c2248;
output c4133;
output c1163;
output c58;
output c2495;
output c2155;
output c1126;
output c133;
output c2362;
output c0376;
output c2179;
output c5226;
output c585;
output c5146;
output c6133;
output c0409;
output c557;
output c6301;
output c4499;
output c5200;
output c1464;
output c0143;
output c6160;
output c3132;
output c3455;
output c2200;
output c0239;
output c4366;
output c0205;
output c4275;
output c5359;
output c0460;
output c2263;
output c0434;
output c298;
output c5464;
output c3301;
output c6309;
output c1257;
output c575;
output c3135;
output c4332;
output c23;
output c5435;
output c4221;
output c1326;
output c2418;
output c6168;
output c3234;
output c1445;
output c4292;
output c5250;
output c0201;
output c4390;
output c2160;
output c6260;
output c5174;
output c1485;
output c6416;
output c1467;
output c0435;
output c519;
output c2141;
output c4164;
output c2170;
output c0227;
output c2331;
output c5302;
output c0165;
output c175;
output c019;
output c0173;
output c1397;
output c2245;
output c3439;
output c4299;
output c644;
output c3151;
output c3483;
output c4245;
output c38;
output c4392;
output c1140;
output c253;
output c5168;
output c059;
output c527;
output c6385;
output c6107;
output c0261;
output c1149;
output c5308;
output c2329;
output c5395;
output c0397;
output c3340;
output c0456;
output c0417;
output c6137;
output c070;
output c1168;
output c6220;
output c4203;
output c2229;
output c416;
output c0363;
output c4470;
output c623;
output c4365;
output c6205;
output c4230;
output c3453;
output c1481;
output c4460;
output c1135;
output c6420;
output c5232;
output c4287;
output c1368;
output c346;
output c3401;
output c3302;
output c6312;
output c2201;
output c6432;
output c47;
output c5160;
output c6439;
output c4250;
output c6298;
output c0332;
output c2303;
output c4431;
output c535;
output c1343;
output c3391;
output c6196;
output c6308;
output c1292;
output c0474;
output c1408;
output c2322;
output c1404;
output c0321;
output c379;
output c5446;
output c2360;
output c1155;
output c2480;
output c293;
output c4414;
output c6148;
output c3392;
output c6498;
output c3195;
output c0233;
output c0118;
output c562;
output c2190;
output c265;
output c264;
output c1427;
output c0413;
output c1210;
output c2432;
output c3349;
output c27;
output c0364;
output c1345;
output c1452;
output c4395;
output c0237;
output c2328;
output c2478;
output c474;
output c2272;
output c19;
output c387;
output c1180;
output c5180;
output c6111;
output c1274;
output c5366;
output c0140;
output c4205;
output c1403;
output c4486;
output c0104;
output c5152;
output c4259;
output c3474;
output c659;
output c5274;
output c1441;
output c5265;
output c4433;
output c0206;
output c0344;
output c2385;
output c071;
output c2262;
output c1128;
output c2477;
output c3336;
output c2249;
output c4422;
output c2448;
output c5161;
output c281;
output c0267;
output c2490;
output c2291;
output c4160;
output c3232;
output c3387;
output c643;
output c4132;
output c3477;
output c1183;
output c282;
output c2119;
output c0276;
output c1166;
output c5173;
output c2379;
output c3363;
output c020;
output c1272;
output c4404;
output c5487;
output c6323;
output c2408;
output c423;
output c2404;
output c668;
output c51;
output c154;
output c5445;
output c2106;
output c5386;
output c5474;
output c0452;
output c1423;
output c0382;
output c1167;
output c3169;
output c3411;
output c15;
output c5225;
output c172;
output c5385;
output c4488;
output c5123;
output c1392;
output c6440;
output c227;
output c1499;
output c369;
output c6184;
output c0253;
output c3328;
output c2483;
output c0334;
output c045;
output c645;
output c1486;
output c6193;
output c2332;
output c6149;
output c089;
output c351;
output c4408;
output c472;
output c5406;
output c6104;
output c4260;
output c038;
output c473;
output c686;
output c4226;
output c1106;
output c5441;
output c0379;
output c127;
output c1281;
output c2308;
output c2301;
output c4232;
output c0100;
output c4150;
output c4398;
output c135;
output c5320;
output c2147;
output c5108;
output c1107;
output c2356;
output c3153;
output c3442;
output c2391;
output c6221;
output c5279;
output c0110;
output c0388;
output c0270;
output c0490;
output c3461;
output c4235;
output c3362;
output c4468;
output c1471;
output c5205;
output c6156;
output c394;
output c5484;
output c2407;
output c5402;
output c6130;
output c0297;
output c1145;
output c210;
output c3172;
output c0280;
output c4482;
output c518;
output c2455;
output c0483;
output c192;
output c2242;
output c0234;
output c4342;
output c2413;
output c4483;
output c466;
output c5262;
output c4293;
output c1188;
output c2131;
output c1439;
output c4401;
output c5119;
output c358;
output c3436;
output c5192;
output c5475;
output c550;
output c1494;
output c470;
output c5290;
output c4393;
output c5209;
output c198;
output c2246;
output c3118;
output c0292;
output c0354;
output c0114;
output c1358;
output c3366;
output c2102;
output c578;
output c573;
output c3236;
output c0222;
output c5169;
output c2216;
output c4469;
output c512;
output c3246;
output c5124;
output c6258;
output c4129;
output c0279;
output c2115;
output c4406;
output c0423;
output c1413;
output c4236;
output c4242;
output c3361;
output c2161;
output c0441;
output c688;
output c07;
output c636;
output c0112;
output c3337;
output c284;
output c0187;
output c4108;
output c6320;
output c3128;
output c248;
output c162;
output c4454;
output c291;
output c34;
output c4335;
output c5354;
output c0163;
output c3163;
output c491;
output c5269;
output c5450;
output c0373;
output c667;
output c6101;
output c5499;
output c1186;
output c2428;
output c1143;
output c2400;
output c382;
output c3486;
output c3335;
output c4184;
output c1246;
output c2420;
output c4233;
output c5261;
output c547;
output c6378;
output c1238;
output c5220;
output c6412;
output c3237;
output c295;
output c4349;
output c3161;
output c4324;
output c454;
output c032;
output c5263;
output c040;
output c390;
output c6244;
output c6448;
output c2372;
output c6434;
output c6120;
output c2213;
output c156;
output c1182;
output c1426;
output c4337;
output c245;
output c3159;
output c55;
output c2458;
output c1412;
output c3243;
output c2221;
output c1268;
output c3130;
output c6286;
output c25;
output c3294;
output c262;
output c5181;
output c2433;
output c420;
output c2377;
output c0400;
output c3448;
output c1320;
output c4173;
output c2122;
output c4444;
output c5118;
output c699;
output c4400;
output c2443;
output c3304;
output c1207;
output c3173;
output c3355;
output c5144;
output c238;
output c3380;
output c5466;
output c6455;
output c5454;
output c4363;
output c360;
output c0274;
output c4336;
output c5121;
output c0398;
output c0449;
output c637;
output c2388;
output c3189;
output c3100;
output c1385;
output c5372;
output c6189;
output c3149;
output c3230;
output c5244;
output c5309;
output c6257;
output c6291;
output c2389;
output c2497;
output c6338;
output c2485;
output c0345;
output c3120;
output c4240;
output c665;
output c6222;
output c6425;
output c2267;
output c212;
output c4269;
output c2437;
output c5381;
output c397;
output c1194;
output c1154;
output c1432;
output c1233;
output c3202;
output c0468;
output c1253;
output c22;
output c4282;
output c0426;
output c5184;
output c525;
output c14;
output c2367;
output c6152;
output c3493;
output c6293;
output c3384;
output c2296;
output c3386;
output c3309;
output c063;
output c0145;
output c0370;
output c3288;
output c4440;
output c2300;
output c2494;
output c477;
output c4211;
output c5155;
output c6488;
output c0375;
output c28;
output c029;
output c3414;
output c6475;
output c1400;
output c3258;
output c4105;
output c5368;
output c06;
output c277;
output c6334;
output c0262;
output c1120;
output c626;
output c0418;
output c0115;
output c4196;
output c4267;
output c534;
output c1298;
output c5278;
output c0361;
output c3498;
output c3269;
output c5419;
output c0220;
output c01;
output c3373;
output c6451;
output c5260;
output c028;
output c1312;
output c5422;
output c4131;
output c335;
output c2415;
output c1378;
output c6340;
output c5337;
output c3101;
output c447;
output c0351;
output c2446;
output c3179;
output c0327;
output c3311;
output c0107;
output c6469;
output c4261;
output c5310;
output c5133;
output c4141;
output c3482;
output c4116;
output c5476;
output c1376;
output c5249;
output c6377;
output c4171;
output c5198;
output c5393;
output c669;
output c136;
output c656;
output c541;
output c5122;
output c393;
output c663;
output c4148;
output c5307;
output c5207;
output c396;
output c4424;
output c0357;
output c5183;
output c655;
output c3291;
output c6471;
output c288;
output c5311;
output c1490;
output c2206;
output c441;
output c3315;
output c2271;
output c0216;
output c1220;
output c0489;
output c3420;
output c2189;
output c2462;
output c2230;
output c3299;
output c03;
output c155;
output c6307;
output c6158;
output c2104;
output c2256;
output c3286;
output c682;
output c1424;
output c3462;
output c2237;
output c3129;
output c1142;
output c0134;
output c047;
output c3321;
output c522;
output c586;
output c4181;
output c551;
output c6310;
output c6232;
output c657;
output c2351;
output c4493;
output c5242;
output c6485;
output c2172;
output c1291;
output c2114;
output c4458;
output c033;
output c2330;
output c6481;
output c3371;
output c4107;
output c5421;
output c6486;
output c6136;
output c0111;
output c4497;
output c338;
output c018;
output c5485;
output c2411;
output c4402;
output c6480;
output c2223;
output c0350;
output c3103;
output c6428;
output c5186;
output c1117;
output c2295;
output c1444;
output c124;
output c222;
output c6151;
output c2187;
output c3263;
output c3213;
output c6150;
output c3111;
output c4389;
output c0223;
output c4353;
output c6387;
output c091;
output c6285;
output c051;
output c340;
output c4426;
output c0147;
output c5273;
output c1416;
output c0416;
output c6269;
output c023;
output c1461;
output c4228;
output c2369;
output c4192;
output c4329;
output c1150;
output c4277;
output c4443;
output c3357;
output c081;
output c1493;
output c126;
output c1369;
output c074;
output c567;
output c5293;
output c2384;
output c5324;
output c5264;
output c2264;
output c0365;
output c6297;
output c163;
output c6213;
output c194;
output c482;
output c596;
output c5404;
output c5467;
output c2238;
output c015;
output c5210;
output c679;
output c2210;
output c68;
output c362;
output c1319;
output c3275;
output c0442;
output c0256;
output c0225;
output c2153;
output c3211;
output c6319;
output c6375;
output c0330;
output c0218;
output c0422;
output c6224;
output c2280;
output c177;
output c2444;
output c6289;
output c3212;
output c6427;
output c1352;
output c455;
output c5462;
output c0464;
output c5347;
output c171;
output c1478;
output c556;
output c4161;
output c5373;
output c2209;
output c3281;
output c526;
output c4223;
output c1361;
output c0202;
output c2452;
output c4478;
output c0136;
output c1497;
output c2392;
output c0335;
output c1259;
output c5442;
output c377;
output c152;
output c6493;
output c3350;
output c1309;
output c1122;
output c6129;
output c0203;
output c0264;
output c1498;
output c199;
output c0257;
output c2162;
output c0462;
output c2243;
output c0437;
output c1449;
output c3375;
output c536;
output c3352;
output c29;
output c6243;
output c0172;
output c6437;
output c5427;
output c042;
output c5277;
output c2217;
output c6278;
output c2136;
output c6228;
output c1170;
output c478;
output c4170;
output c115;
output c055;
output c2297;
output c3283;
output c094;
output c02;
output c2273;
output c0479;
output c4434;
output c5424;
output c3427;
output c3222;
output c6128;
output c3404;
output c6383;
output c1316;
output c1422;
output c4289;
output c1304;
output c5334;
output c6142;
output c5258;
output c241;
output c0378;
output c2357;
output c3114;
output c5376;
output c271;
output c0362;
output c529;
output c6496;
output c683;
output c184;
output c1190;
output c4145;
output c4183;
output c3146;
output c1333;
output c6154;
output c6400;
output c2399;
output c662;
output c629;
output c1359;
output c5482;
output c0447;
output c4412;
output c4368;
output c1231;
output c2423;
output c1258;
output c0406;
output c2337;
output c6457;
output c0159;
output c5360;
output c035;
output c138;
output c3244;
output c4229;
output c6199;
output c5109;
output c0316;
output c093;
output c576;
output c0186;
output c0258;
output c5229;
output c1177;
output c4220;
output c6125;
output c6407;
output c0320;
output c4206;
output c3419;
output c4352;
output c471;
output c5339;
output c545;
output c6132;
output c3231;
output c0314;
output c542;
output c129;
output c3171;
output c275;
output c2257;
output c6408;
output c0372;
output c650;
output c6401;
output c4252;
output c4263;
output c4462;
output c3217;
output c5396;
output c3198;
output c1338;
output c0369;
output c2283;
output c052;
output c0138;
output c246;
output c4428;
output c4435;
output c6417;
output c2226;
output c1242;
output c489;
output c620;
output c42;
output c1394;
output c164;
output c458;
output c6185;
output c0208;
output c3324;
output c3105;
output c1221;
output c3119;
output c5332;
output c1455;
output c5215;
output c3360;
output c1301;
output c438;
output c211;
output c4126;
output c0352;
output c2100;
output c3259;
output c119;
output c5428;
output c658;
output c3126;
output c6195;
output c3143;
output c0231;
output c6139;
output c4188;
output c4124;
output c317;
output c6274;
output c185;
output c6313;
output c2110;
output c3157;
output c021;
output c3438;
output c1114;
output c04;
output c2326;
output c1138;
output c3374;
output c6206;
output c1118;
output c5117;
output c6405;
output c0333;
output c4152;
output c4350;
output c0155;
output c6410;
output c614;
output c487;
output c677;
output c2194;
output c6223;
output c4333;
output c4146;
output c1363;
output c085;
output c448;
output c2250;
output c685;
output c220;
output c2394;
output c2167;
output c367;
output c0319;
output c391;
output c5139;
output c0387;
output c2181;
output c069;
output c5191;
output c0127;
output c6472;
output c5369;
output c5423;
output c1414;
output c4487;
output c0311;
output c0244;
output c354;
output c6215;
output c0309;
output c6219;
output c0243;
output c0402;
output c6474;
output c515;
output c1260;
output c0494;
output c492;
output c4429;
output c0153;
output c5461;
output c4322;
output c239;
output c234;
output c5490;
output c112;
output c5259;
output c6296;
output c014;
output c5345;
output c5384;
output c5299;
output c2244;
output c0194;
output c1379;
output c1125;
output c2289;
output c1473;
output c188;
output c1487;
output c3465;
output c0102;
output c5156;
output c1267;
output c6344;
output c3467;
output c333;
output c2397;
output c6371;
output c3412;
output c328;
output c2463;
output c4347;
output c316;
output c3343;
output c5426;
output c5282;
output c3377;
output c183;
output c5496;
output c4179;
output c3156;
output c3456;
output c3487;
output c4359;
output c2123;
output c5177;
output c0432;
output c6211;
output c0478;
output c4201;
output c640;
output c4258;
output c347;
output c0401;
output c0349;
output c0383;
output c235;
output c4419;
output c5350;
output c292;
output c520;
output c6254;
output c6447;
output c0366;
output c031;
output c1205;
output c1204;
output c1139;
output c3144;
output c3354;
output c3345;
output c6190;
output c1223;
output c3470;
output c5237;
output c6217;
output c1266;
output c1474;
output c5254;
output c5495;
output c137;
output c0164;
output c544;
output c1380;
output c6397;
output c2258;
output c0484;
output c0259;
output c4331;
output c4442;
output c3348;
output c531;
output c6373;
output c226;
output c533;
output c457;
output c6165;
output c5398;
output c4473;
output c634;
output c1111;
output c3407;
output c6318;
output c17;
output c181;
output c4432;
output c3446;
output c5383;
output c4253;
output c3451;
output c1431;
output c6176;
output c5420;
output c132;
output c21;
output c0495;
output c1323;
output c4137;
output c5486;
output c5483;
output c3351;
output c5296;
output c419;
output c5159;
output c26;
output c694;
output c6473;
output c1409;
output c4157;
output c5371;
output c2270;
output c3400;
output c3339;
output c4187;
output c540;
output c1406;
output c327;
output c6429;
output c2353;
output c6251;
output c2317;
output c4239;
output c1195;
output c5255;

assign c00 = ~x68;
assign c02 =  x54;
assign c04 =  x3 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c06 =  x44;
assign c08 =  x64;
assign c010 =  x85;
assign c012 = ~x88;
assign c014 = ~x68;
assign c016 =  x2 &  x6 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c018 =  x34;
assign c020 =  x14 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c022 =  x24;
assign c024 = ~x87;
assign c026 =  x83;
assign c028 =  x25;
assign c030 = ~x67;
assign c032 =  x74;
assign c034 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c036 =  x24;
assign c038 =  x0 &  x17 &  x18 &  x19 &  x20 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x39 &  x40 &  x47 &  x48 &  x49 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x70 &  x76 &  x77 &  x79 &  x80 &  x86 &  x88 &  x90 & ~x2 & ~x4 & ~x22 & ~x23 & ~x24 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x53 & ~x54 & ~x62 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c040 = ~x68;
assign c042 =  x74;
assign c044 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c046 = ~x40;
assign c048 = ~x68;
assign c050 =  x74;
assign c052 = ~x49;
assign c054 =  x54;
assign c056 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x14 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c058 =  x24;
assign c060 = ~x67;
assign c062 =  x6 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c064 = ~x47;
assign c066 =  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x95;
assign c068 =  x74;
assign c070 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c072 =  x35;
assign c074 =  x74;
assign c076 = ~x36;
assign c078 =  x84;
assign c080 = ~x19;
assign c082 =  x75;
assign c084 =  x83;
assign c086 = ~x18;
assign c088 = ~x36;
assign c090 =  x54;
assign c092 = ~x67;
assign c094 = ~x18;
assign c096 = ~x57;
assign c098 = ~x87;
assign c0100 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c0102 =  x3 &  x17 &  x18 &  x19 &  x26 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x48 &  x49 &  x50 &  x51 &  x56 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x82 & ~x83 & ~x92 & ~x93 & ~x95;
assign c0104 =  x24;
assign c0106 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x61 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c0108 =  x94;
assign c0110 =  x54;
assign c0112 =  x43;
assign c0114 =  x65;
assign c0116 = ~x49;
assign c0118 = ~x76;
assign c0120 =  x23;
assign c0122 =  x83;
assign c0124 =  x54;
assign c0126 = ~x18;
assign c0128 = ~x47;
assign c0130 = ~x47;
assign c0132 =  x23;
assign c0134 = ~x49;
assign c0136 = ~x28;
assign c0138 =  x33;
assign c0140 = ~x40;
assign c0142 = ~x88;
assign c0144 =  x74;
assign c0146 =  x95;
assign c0148 = ~x27;
assign c0150 =  x25;
assign c0152 =  x84;
assign c0154 =  x43;
assign c0156 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x4 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c0158 =  x44;
assign c0160 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x8 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x61 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c0162 =  x75;
assign c0164 =  x16 &  x17 &  x18 &  x19 &  x20 &  x21 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c0166 = ~x36;
assign c0168 =  x8 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x28 &  x29 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x69 &  x70 &  x71 &  x76 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x90 &  x91 & ~x22 & ~x24 & ~x25 & ~x32 & ~x35 & ~x43 & ~x45 & ~x52 & ~x62 & ~x63 & ~x64 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x83 & ~x84 & ~x92 & ~x93 & ~x94 & ~x95;
assign c0170 = ~x18;
assign c0172 = ~x39;
assign c0174 = ~x47;
assign c0176 = ~x87;
assign c0178 = ~x87;
assign c0180 =  x25;
assign c0182 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x9 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c0184 = ~x47;
assign c0186 =  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c0188 =  x75;
assign c0190 = ~x47;
assign c0192 = ~x68;
assign c0194 =  x2 &  x16 &  x19 &  x26 &  x27 &  x30 &  x36 &  x37 &  x46 &  x48 &  x56 &  x57 &  x59 &  x60 &  x66 &  x67 &  x68 &  x70 &  x76 &  x77 &  x78 &  x79 &  x88 &  x90 & ~x0 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x35 & ~x44 & ~x52 & ~x54 & ~x55 & ~x62 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x95;
assign c0196 = ~x69;
assign c0198 =  x24;
assign c0200 = ~x49;
assign c0202 =  x23;
assign c0204 = ~x19;
assign c0206 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c0208 =  x0 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c0210 =  x0 &  x3 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c0212 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c0214 =  x43;
assign c0216 = ~x57;
assign c0218 =  x43;
assign c0220 =  x94;
assign c0222 = ~x17;
assign c0224 = ~x49;
assign c0226 = ~x19;
assign c0228 = ~x88;
assign c0230 = ~x67;
assign c0232 = ~x88;
assign c0234 =  x84;
assign c0236 = ~x36;
assign c0238 = ~x68;
assign c0240 = ~x17;
assign c0242 = ~x20;
assign c0244 =  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c0246 =  x54;
assign c0248 =  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x15 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c0250 = ~x78;
assign c0252 =  x94 &  x95;
assign c0254 =  x43;
assign c0256 =  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x1 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c0258 =  x64;
assign c0260 = ~x58;
assign c0262 = ~x57;
assign c0264 =  x25;
assign c0266 = ~x47;
assign c0268 = ~x49;
assign c0270 = ~x28;
assign c0272 =  x0 &  x3 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x70 &  x77 &  x78 &  x88 &  x90 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x62 & ~x63 & ~x64 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94;
assign c0274 =  x23;
assign c0276 = ~x29;
assign c0278 = ~x29;
assign c0280 = ~x40;
assign c0282 = ~x18;
assign c0284 =  x54;
assign c0286 =  x85;
assign c0288 = ~x18;
assign c0290 =  x3 &  x6 &  x16 &  x18 &  x19 &  x26 &  x27 &  x28 &  x37 &  x38 &  x39 &  x40 &  x48 &  x49 &  x56 &  x60 &  x66 &  x67 &  x69 &  x77 &  x78 &  x79 &  x86 &  x88 & ~x5 & ~x24 & ~x25 & ~x35 & ~x44 & ~x53 & ~x55 & ~x64 & ~x65 & ~x74 & ~x84 & ~x85 & ~x93 & ~x95;
assign c0292 = ~x68;
assign c0294 = ~x40;
assign c0296 =  x84;
assign c0298 =  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c0300 = ~x57;
assign c0302 =  x74;
assign c0304 =  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c0306 =  x74;
assign c0308 = ~x49;
assign c0310 =  x44;
assign c0312 = ~x18;
assign c0314 = ~x49;
assign c0316 =  x3 &  x6 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c0318 =  x34;
assign c0320 =  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c0322 = ~x67;
assign c0324 =  x24;
assign c0326 =  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c0328 =  x43;
assign c0330 =  x44;
assign c0332 = ~x79;
assign c0334 = ~x40;
assign c0336 =  x44;
assign c0338 =  x44;
assign c0340 = ~x89;
assign c0342 =  x23;
assign c0344 =  x24;
assign c0346 = ~x67;
assign c0348 = ~x40;
assign c0350 =  x54;
assign c0352 =  x75;
assign c0354 =  x3 &  x8 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c0356 = ~x88;
assign c0358 =  x24;
assign c0360 = ~x67;
assign c0362 = ~x36;
assign c0364 = ~x18;
assign c0366 =  x3 &  x16 &  x17 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x50 &  x51 &  x56 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x80 &  x86 &  x87 &  x89 &  x90 &  x91 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x44 & ~x45 & ~x52 & ~x53 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x74 & ~x75 & ~x83 & ~x84 & ~x92 & ~x94;
assign c0368 = ~x57;
assign c0370 = ~x78;
assign c0372 =  x23;
assign c0374 =  x16 &  x17 &  x19 &  x20 &  x26 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x60 &  x67 &  x68 &  x70 &  x76 &  x78 &  x79 &  x80 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x4 & ~x10 & ~x22 & ~x23 & ~x25 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x53 & ~x55 & ~x62 & ~x64 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x92 & ~x94 & ~x95;
assign c0376 =  x25;
assign c0378 = ~x69;
assign c0380 = ~x78;
assign c0382 = ~x68;
assign c0384 =  x23;
assign c0386 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x10 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c0388 =  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c0390 = ~x69;
assign c0392 =  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c0394 = ~x47;
assign c0396 =  x54;
assign c0398 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c0400 = ~x59;
assign c0402 = ~x17;
assign c0404 =  x24;
assign c0406 = ~x78;
assign c0408 =  x43;
assign c0410 = ~x17;
assign c0412 = ~x68;
assign c0414 = ~x37;
assign c0416 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c0418 =  x16 &  x17 &  x18 &  x19 &  x20 &  x21 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x14 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c0420 =  x3 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c0422 = ~x28;
assign c0424 = ~x18;
assign c0426 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c0428 =  x54;
assign c0430 = ~x17;
assign c0432 =  x65;
assign c0434 =  x75;
assign c0436 = ~x18;
assign c0438 =  x24;
assign c0440 = ~x88;
assign c0442 =  x34;
assign c0444 = ~x88;
assign c0446 =  x84;
assign c0448 =  x74;
assign c0450 = ~x57;
assign c0452 =  x6 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c0454 =  x94;
assign c0456 =  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c0458 = ~x48;
assign c0460 = ~x88;
assign c0462 =  x35;
assign c0464 =  x84;
assign c0466 =  x6 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c0468 =  x74;
assign c0470 =  x44;
assign c0472 = ~x38;
assign c0474 = ~x39;
assign c0476 =  x54;
assign c0478 =  x95;
assign c0480 =  x74;
assign c0482 =  x1 &  x17 &  x18 &  x26 &  x27 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x47 &  x48 &  x50 &  x57 &  x58 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x87 &  x89 &  x90 &  x91 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x34 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x72 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x94;
assign c0484 = ~x19;
assign c0486 =  x24;
assign c0488 =  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c0490 = ~x68;
assign c0492 =  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c0494 = ~x50;
assign c0496 = ~x18;
assign c0498 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c01 = ~x28;
assign c03 = ~x37;
assign c05 =  x22;
assign c07 = ~x76;
assign c09 =  x92;
assign c011 = ~x46;
assign c013 =  x25;
assign c015 = ~x76;
assign c017 =  x35;
assign c019 = ~x67;
assign c021 = ~x46;
assign c023 = ~x76;
assign c025 = ~x26;
assign c027 = ~x16;
assign c029 = ~x36;
assign c033 =  x22;
assign c035 = ~x77;
assign c037 = ~x77;
assign c039 = ~x36;
assign c043 = ~x78;
assign c045 = ~x29;
assign c047 = ~x57;
assign c049 = ~x58;
assign c051 = ~x47;
assign c053 = ~x56;
assign c055 = ~x66;
assign c057 = ~x16;
assign c059 = ~x66;
assign c061 = ~x77;
assign c063 = ~x66;
assign c065 = ~x56;
assign c067 = ~x26;
assign c069 =  x22;
assign c071 = ~x26;
assign c073 = ~x38;
assign c077 = ~x38;
assign c079 = ~x28;
assign c081 = ~x76;
assign c083 = ~x78;
assign c085 = ~x39;
assign c087 = ~x36;
assign c089 =  x55;
assign c091 = ~x56;
assign c093 =  x74 & ~x78;
assign c095 =  x55;
assign c097 = ~x26;
assign c099 = ~x48;
assign c0101 =  x75;
assign c0103 = ~x76;
assign c0107 = ~x66;
assign c0109 = ~x46;
assign c0111 = ~x27;
assign c0113 =  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x3 & ~x23 & ~x25 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x71 & ~x72 & ~x73 & ~x74 & ~x83 & ~x84 & ~x93 & ~x94 & ~x95;
assign c0115 = ~x16;
assign c0117 =  x75;
assign c0119 = ~x76;
assign c0121 =  x25 & ~x67;
assign c0123 =  x45;
assign c0127 =  x84;
assign c0129 = ~x6 & ~x60;
assign c0131 = ~x87;
assign c0133 =  x5 & ~x80;
assign c0135 = ~x76;
assign c0137 =  x45;
assign c0139 = ~x78;
assign c0141 =  x62;
assign c0143 = ~x76;
assign c0145 = ~x88;
assign c0147 = ~x16;
assign c0149 =  x85;
assign c0151 =  x54;
assign c0153 = ~x76;
assign c0155 = ~x26;
assign c0157 = ~x56;
assign c0159 = ~x26;
assign c0161 = ~x19;
assign c0169 = ~x37 & ~x66;
assign c0171 = ~x38;
assign c0173 = ~x46;
assign c0175 =  x62;
assign c0177 =  x44;
assign c0179 =  x35;
assign c0181 = ~x78;
assign c0183 = ~x36;
assign c0185 = ~x37 & ~x87;
assign c0187 = ~x38;
assign c0189 = ~x26;
assign c0191 = ~x86;
assign c0193 = ~x47;
assign c0195 = ~x58;
assign c0197 = ~x87;
assign c0199 = ~x76;
assign c0201 = ~x16;
assign c0203 = ~x76;
assign c0205 = ~x56;
assign c0207 = ~x26;
assign c0211 =  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c0213 =  x45;
assign c0217 = ~x56;
assign c0219 =  x64;
assign c0221 = ~x56;
assign c0223 = ~x48;
assign c0227 = ~x86;
assign c0229 = ~x17;
assign c0231 = ~x46;
assign c0233 =  x62;
assign c0235 = ~x16;
assign c0237 = ~x30;
assign c0241 = ~x38;
assign c0245 =  x95;
assign c0247 = ~x77;
assign c0249 =  x62;
assign c0251 = ~x38;
assign c0253 = ~x26;
assign c0255 =  x25;
assign c0257 = ~x38;
assign c0259 =  x35;
assign c0263 = ~x26;
assign c0265 =  x24;
assign c0267 = ~x66;
assign c0271 = ~x69;
assign c0273 = ~x58;
assign c0275 = ~x86;
assign c0277 = ~x28;
assign c0279 = ~x26;
assign c0281 = ~x16;
assign c0283 = ~x58;
assign c0285 = ~x20;
assign c0287 = ~x66;
assign c0289 = ~x26;
assign c0291 = ~x26;
assign c0293 =  x45;
assign c0295 = ~x58;
assign c0297 =  x25;
assign c0299 =  x85;
assign c0301 =  x24;
assign c0303 = ~x56;
assign c0309 = ~x16;
assign c0311 = ~x6 & ~x60;
assign c0315 =  x55;
assign c0317 =  x23;
assign c0319 =  x55;
assign c0321 = ~x87;
assign c0323 = ~x56;
assign c0325 = ~x16;
assign c0327 = ~x76;
assign c0331 = ~x16;
assign c0333 = ~x47;
assign c0335 =  x16 &  x17 &  x18 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x76 &  x77 &  x78 &  x79 &  x80 &  x81 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x94 & ~x95;
assign c0337 = ~x58;
assign c0339 = ~x76;
assign c0341 = ~x90;
assign c0343 =  x92;
assign c0345 = ~x46;
assign c0347 = ~x58;
assign c0349 = ~x76;
assign c0353 =  x51 & ~x80;
assign c0355 = ~x78;
assign c0357 = ~x28;
assign c0359 = ~x56;
assign c0361 = ~x27;
assign c0363 = ~x58;
assign c0365 =  x75;
assign c0367 = ~x46;
assign c0369 = ~x66;
assign c0371 = ~x77;
assign c0373 = ~x18;
assign c0375 =  x22;
assign c0377 = ~x77;
assign c0379 = ~x36;
assign c0381 = ~x29;
assign c0383 =  x35;
assign c0385 =  x35;
assign c0387 =  x55;
assign c0389 =  x0 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x3 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c0391 = ~x16;
assign c0393 = ~x30;
assign c0395 =  x55;
assign c0397 = ~x26;
assign c0399 = ~x86;
assign c0401 = ~x76;
assign c0403 = ~x86;
assign c0405 = ~x26;
assign c0407 = ~x27;
assign c0409 =  x23;
assign c0411 = ~x36;
assign c0413 = ~x36;
assign c0415 =  x45;
assign c0417 = ~x76;
assign c0419 = ~x60;
assign c0421 = ~x26;
assign c0423 = ~x76;
assign c0427 = ~x86;
assign c0429 = ~x18;
assign c0431 =  x24;
assign c0435 = ~x66;
assign c0437 = ~x17;
assign c0439 =  x54;
assign c0441 = ~x37;
assign c0443 = ~x26;
assign c0445 = ~x66;
assign c0447 = ~x26;
assign c0449 = ~x37;
assign c0457 = ~x66;
assign c0459 = ~x76;
assign c0461 = ~x86;
assign c0463 =  x73;
assign c0465 = ~x66;
assign c0467 = ~x87;
assign c0469 = ~x76;
assign c0471 = ~x47;
assign c0473 = ~x56;
assign c0475 = ~x28;
assign c0477 = ~x37;
assign c0479 = ~x26;
assign c0481 = ~x76;
assign c0483 = ~x66;
assign c0485 =  x35;
assign c0487 =  x25;
assign c0489 = ~x18;
assign c0491 = ~x26;
assign c0493 = ~x77;
assign c0495 = ~x66;
assign c0497 = ~x27;
assign c0499 = ~x48;
assign c10 =  x55;
assign c12 = ~x37;
assign c14 = ~x26;
assign c16 = ~x76;
assign c18 =  x44;
assign c110 =  x85;
assign c112 = ~x46;
assign c114 = ~x26;
assign c116 = ~x46;
assign c118 = ~x77;
assign c120 = ~x16;
assign c122 = ~x16;
assign c124 = ~x67;
assign c126 = ~x66;
assign c128 = ~x46;
assign c132 = ~x46;
assign c134 = ~x46;
assign c136 =  x55;
assign c138 =  x35;
assign c140 = ~x58;
assign c142 =  x12 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x2 & ~x3 & ~x14 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c146 = ~x56;
assign c148 =  x75;
assign c150 =  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x21 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x0 & ~x1 & ~x2 & ~x3 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c152 = ~x16;
assign c154 = ~x17;
assign c156 = ~x76;
assign c158 = ~x86;
assign c160 = ~x76;
assign c162 = ~x66;
assign c164 = ~x56;
assign c166 =  x44;
assign c168 =  x44;
assign c170 = ~x76;
assign c172 =  x45;
assign c174 = ~x66;
assign c176 = ~x76;
assign c178 = ~x67;
assign c180 = ~x67;
assign c182 = ~x36;
assign c184 = ~x57;
assign c188 = ~x66;
assign c190 = ~x48;
assign c192 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x1 & ~x2 & ~x3 & ~x5 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x61 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c194 = ~x68;
assign c196 = ~x56;
assign c198 =  x65;
assign c1100 = ~x26;
assign c1102 =  x65;
assign c1104 = ~x86;
assign c1106 =  x34;
assign c1108 = ~x36;
assign c1110 = ~x26;
assign c1112 = ~x77;
assign c1114 =  x85;
assign c1116 = ~x46;
assign c1120 = ~x56;
assign c1122 = ~x66;
assign c1124 = ~x66;
assign c1126 = ~x26;
assign c1128 = ~x36;
assign c1130 = ~x26;
assign c1132 =  x16 &  x17 &  x18 &  x19 &  x20 &  x21 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x61 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x1 & ~x2 & ~x3 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c1134 =  x35;
assign c1136 =  x85;
assign c1138 =  x53 & ~x26;
assign c1140 =  x74;
assign c1142 = ~x17;
assign c1144 = ~x76;
assign c1146 = ~x26;
assign c1148 =  x55;
assign c1150 = ~x66;
assign c1152 = ~x26;
assign c1154 =  x45;
assign c1156 =  x45;
assign c1158 = ~x76;
assign c1160 = ~x67;
assign c1162 = ~x76;
assign c1164 = ~x26;
assign c1166 =  x65;
assign c1168 = ~x76;
assign c1170 =  x9 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x1 & ~x2 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x61 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c1172 =  x83;
assign c1174 = ~x86;
assign c1176 = ~x76;
assign c1178 = ~x86;
assign c1180 = ~x76;
assign c1184 = ~x26;
assign c1186 = ~x67;
assign c1188 = ~x37;
assign c1190 = ~x56;
assign c1192 = ~x36;
assign c1194 = ~x39;
assign c1196 = ~x77;
assign c1200 = ~x36;
assign c1202 =  x55 & ~x46;
assign c1204 = ~x76;
assign c1206 = ~x56;
assign c1208 = ~x17;
assign c1210 = ~x26;
assign c1214 = ~x26;
assign c1216 = ~x26;
assign c1218 =  x45;
assign c1220 =  x45;
assign c1222 = ~x26;
assign c1224 = ~x26;
assign c1226 = ~x89;
assign c1228 = ~x66;
assign c1230 =  x75 & ~x36;
assign c1232 = ~x26;
assign c1234 = ~x90;
assign c1236 = ~x56;
assign c1238 =  x16 &  x17 &  x18 &  x19 &  x20 &  x21 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x0 & ~x1 & ~x2 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x61 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c1240 = ~x27;
assign c1242 = ~x87;
assign c1244 =  x95;
assign c1246 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x2 & ~x3 & ~x10 & ~x12 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c1248 =  x35;
assign c1250 =  x85;
assign c1252 = ~x16;
assign c1254 =  x45;
assign c1256 = ~x17;
assign c1258 = ~x77;
assign c1260 = ~x86;
assign c1262 =  x45;
assign c1264 =  x1 &  x2 &  x3 &  x4 &  x5 &  x16 &  x17 &  x18 &  x19 &  x20 &  x21 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x0 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c1268 =  x65;
assign c1270 = ~x26;
assign c1272 =  x45;
assign c1274 = ~x46;
assign c1276 =  x54;
assign c1278 = ~x17;
assign c1280 =  x55;
assign c1282 =  x55;
assign c1284 =  x75;
assign c1286 = ~x76;
assign c1288 = ~x26;
assign c1290 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x1 & ~x2 & ~x3 & ~x5 & ~x6 & ~x13 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c1292 = ~x37;
assign c1294 = ~x46;
assign c1296 = ~x16;
assign c1298 = ~x87;
assign c1300 =  x74 & ~x19;
assign c1302 = ~x76;
assign c1306 = ~x76;
assign c1308 = ~x26;
assign c1310 = ~x16;
assign c1312 = ~x66;
assign c1314 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x2 & ~x3 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x61 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c1316 =  x44;
assign c1318 = ~x76;
assign c1320 = ~x26;
assign c1322 = ~x86;
assign c1324 = ~x16;
assign c1326 = ~x26;
assign c1328 = ~x76;
assign c1330 = ~x16;
assign c1332 = ~x36;
assign c1334 = ~x56;
assign c1336 = ~x66;
assign c1338 = ~x26;
assign c1340 = ~x47;
assign c1342 =  x65;
assign c1344 =  x85;
assign c1346 = ~x77;
assign c1348 = ~x26;
assign c1350 = ~x66;
assign c1352 = ~x26;
assign c1354 = ~x56;
assign c1356 = ~x26;
assign c1358 = ~x38;
assign c1360 =  x1 &  x2 &  x3 &  x4 &  x5 &  x16 &  x17 &  x18 &  x19 &  x20 &  x21 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x0 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c1362 =  x24;
assign c1364 = ~x26;
assign c1366 = ~x76;
assign c1370 =  x1 &  x2 &  x3 &  x4 &  x5 &  x16 &  x17 &  x18 &  x19 &  x20 &  x21 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x0 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c1372 = ~x16;
assign c1374 = ~x57;
assign c1376 = ~x76;
assign c1378 = ~x77;
assign c1380 =  x25;
assign c1382 = ~x56;
assign c1384 = ~x66;
assign c1386 = ~x46;
assign c1388 =  x44;
assign c1390 =  x54;
assign c1392 =  x25;
assign c1394 = ~x76;
assign c1396 = ~x38;
assign c1398 = ~x86;
assign c1400 = ~x16;
assign c1404 =  x83;
assign c1408 = ~x86;
assign c1410 = ~x86;
assign c1412 = ~x87;
assign c1414 = ~x56;
assign c1416 =  x24;
assign c1418 = ~x28;
assign c1420 = ~x76;
assign c1422 =  x65;
assign c1424 = ~x26;
assign c1426 =  x1 &  x2 &  x3 &  x4 &  x5 &  x16 &  x17 &  x18 &  x19 &  x20 &  x21 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x0 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c1428 = ~x76;
assign c1430 = ~x67;
assign c1432 =  x35;
assign c1434 =  x45 &  x95;
assign c1436 =  x4 &  x13 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x2 & ~x3 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c1438 =  x45;
assign c1440 =  x74;
assign c1442 =  x24;
assign c1444 = ~x36;
assign c1446 = ~x29;
assign c1450 = ~x76;
assign c1452 = ~x36;
assign c1456 = ~x76;
assign c1458 =  x85;
assign c1460 =  x25;
assign c1462 = ~x66;
assign c1464 =  x35;
assign c1466 = ~x66;
assign c1468 = ~x46;
assign c1470 = ~x16;
assign c1472 =  x75;
assign c1474 =  x55;
assign c1476 =  x9 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x1 & ~x2 & ~x3 & ~x11 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c1478 = ~x56;
assign c1480 = ~x46;
assign c1482 = ~x66;
assign c1484 = ~x89;
assign c1486 = ~x18;
assign c1488 =  x45;
assign c1490 = ~x16;
assign c1492 =  x65 & ~x36;
assign c1494 = ~x36;
assign c1496 =  x45;
assign c1498 = ~x36;
assign c11 = ~x70;
assign c13 =  x0 &  x5 &  x16 &  x26 &  x46 &  x86 & ~x43 & ~x44 & ~x75;
assign c15 =  x2 &  x17 &  x18 &  x20 &  x26 &  x27 &  x36 &  x37 &  x39 &  x47 &  x50 &  x56 &  x57 &  x59 &  x60 &  x67 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x87 &  x90 & ~x1 & ~x22 & ~x23 & ~x24 & ~x32 & ~x43 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c17 =  x62;
assign c19 = ~x80;
assign c111 =  x36 &  x56 &  x78 &  x81 & ~x9 & ~x42;
assign c113 =  x3 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x30 &  x31 &  x37 &  x39 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x58 &  x59 &  x60 &  x67 &  x68 &  x70 &  x78 &  x80 &  x86 &  x87 &  x89 &  x90 & ~x1 & ~x22 & ~x24 & ~x25 & ~x34 & ~x35 & ~x42 & ~x43 & ~x45 & ~x52 & ~x55 & ~x62 & ~x63 & ~x64 & ~x72 & ~x73 & ~x75 & ~x85 & ~x93 & ~x95;
assign c115 = ~x80;
assign c117 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x3 & ~x4 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c119 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c121 = ~x31;
assign c123 = ~x80;
assign c125 = ~x80;
assign c127 =  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c129 =  x52;
assign c131 =  x82;
assign c133 =  x62;
assign c135 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c137 = ~x90;
assign c139 =  x3 &  x20 &  x27 &  x28 &  x30 &  x48 &  x49 &  x56 &  x76 &  x87 & ~x4 & ~x23 & ~x34 & ~x35 & ~x64 & ~x83;
assign c141 =  x2 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x39 &  x40 &  x46 &  x48 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x88 &  x89 &  x90 & ~x1 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x35 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x73 & ~x74 & ~x75 & ~x82 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c145 =  x72;
assign c147 =  x18 &  x46 &  x61 &  x68 & ~x24 & ~x33 & ~x41 & ~x45 & ~x84 & ~x95;
assign c149 =  x3 &  x18 &  x20 &  x26 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x88 &  x89 & ~x5 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x63 & ~x64 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x94 & ~x95;
assign c151 = ~x80;
assign c153 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c155 =  x0 &  x6 & ~x95;
assign c157 =  x22;
assign c159 =  x52;
assign c161 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x36 &  x37 &  x38 &  x46 &  x49 &  x50 &  x56 &  x57 &  x66 &  x67 &  x68 &  x78 &  x86 &  x87 &  x88 &  x89 & ~x4 & ~x22 & ~x23 & ~x24 & ~x33 & ~x34 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x65 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c163 =  x16 &  x18 &  x36 &  x37 &  x38 &  x46 &  x47 &  x48 &  x56 &  x57 &  x59 &  x66 &  x67 &  x69 &  x70 &  x76 &  x77 &  x86 &  x87 & ~x23 & ~x25 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x84 & ~x85 & ~x91 & ~x92 & ~x93 & ~x94 & ~x95;
assign c165 = ~x70;
assign c167 =  x22;
assign c169 = ~x51;
assign c173 =  x2 &  x17 &  x18 &  x20 &  x26 &  x27 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x60 &  x67 &  x68 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x88 &  x89 &  x91 & ~x4 & ~x22 & ~x23 & ~x24 & ~x33 & ~x34 & ~x35 & ~x44 & ~x53 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x85 & ~x93 & ~x95;
assign c175 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c177 =  x0 &  x5 & ~x44;
assign c179 =  x22;
assign c181 =  x0 &  x5 &  x27 &  x29 &  x36 &  x66 & ~x44 & ~x55 & ~x65;
assign c183 = ~x80;
assign c185 =  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x49 &  x50 &  x51 &  x59 &  x66 &  x67 &  x68 &  x69 &  x71 &  x79 &  x80 &  x86 &  x87 &  x90 & ~x1 & ~x23 & ~x34 & ~x43 & ~x44 & ~x52 & ~x54 & ~x55 & ~x64 & ~x65 & ~x73 & ~x83 & ~x84 & ~x85 & ~x95;
assign c187 =  x92;
assign c189 = ~x71;
assign c191 = ~x71;
assign c193 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x3 & ~x22 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x52 & ~x53 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c195 =  x2 &  x16 &  x18 &  x19 &  x20 &  x26 &  x27 &  x29 &  x30 &  x36 &  x38 &  x39 &  x46 &  x47 &  x48 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x80 &  x86 &  x87 &  x88 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x92 & ~x94 & ~x95;
assign c197 =  x7 &  x16 &  x36 &  x48 &  x49 &  x59 &  x71 &  x80 &  x81 & ~x54;
assign c199 = ~x51;
assign c1101 =  x77 &  x79 &  x80 &  x81 & ~x45;
assign c1103 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c1105 =  x16 &  x17 &  x18 &  x27 &  x37 &  x38 &  x46 &  x47 &  x48 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x77 &  x86 & ~x21 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x91 & ~x92 & ~x93 & ~x94;
assign c1107 =  x1 &  x19 &  x28 &  x36 &  x67 & ~x5 & ~x35 & ~x74 & ~x75;
assign c1109 =  x1 &  x66 & ~x5 & ~x32;
assign c1111 =  x52;
assign c1113 = ~x51;
assign c1115 =  x92;
assign c1117 =  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c1119 = ~x80;
assign c1121 =  x0 &  x5;
assign c1123 =  x32;
assign c1125 =  x82;
assign c1127 =  x1 &  x17 &  x18 &  x19 &  x27 &  x36 &  x46 &  x48 &  x57 &  x76 &  x77 &  x87 &  x88 & ~x5 & ~x24 & ~x34 & ~x43 & ~x44 & ~x45 & ~x53 & ~x55 & ~x65 & ~x84 & ~x85 & ~x93 & ~x94;
assign c1129 = ~x51;
assign c1131 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x22 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x93 & ~x95;
assign c1133 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c1135 =  x3 &  x16 &  x19 &  x26 &  x38 &  x46 &  x49 &  x58 &  x59 &  x66 &  x67 &  x77 &  x86 & ~x4 & ~x24 & ~x25 & ~x34 & ~x44 & ~x54 & ~x55 & ~x74 & ~x75 & ~x83 & ~x84;
assign c1137 =  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x30 &  x37 &  x38 &  x46 &  x47 &  x48 &  x50 &  x51 &  x58 &  x59 &  x67 &  x70 &  x76 &  x77 &  x79 &  x86 &  x87 &  x89 &  x90 & ~x0 & ~x4 & ~x22 & ~x23 & ~x32 & ~x34 & ~x44 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x85 & ~x92 & ~x93 & ~x95;
assign c1139 = ~x51;
assign c1141 = ~x31;
assign c1143 =  x2 &  x18 &  x19 &  x20 &  x26 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x47 &  x48 &  x50 &  x60 &  x67 &  x68 &  x86 &  x88 & ~x5 & ~x23 & ~x24 & ~x25 & ~x33 & ~x43 & ~x44 & ~x45 & ~x52 & ~x54 & ~x55 & ~x63 & ~x64 & ~x73 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x95;
assign c1145 = ~x31;
assign c1147 =  x92;
assign c1149 =  x3 &  x16 &  x17 &  x18 &  x19 &  x27 &  x28 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x56 &  x57 &  x60 &  x66 &  x67 &  x68 &  x77 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x5 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x84 & ~x85 & ~x95;
assign c1151 = ~x31;
assign c1153 =  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x49 &  x51 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x80 &  x86 &  x87 &  x88 &  x89 & ~x2 & ~x24 & ~x25 & ~x33 & ~x34 & ~x43 & ~x44 & ~x45 & ~x53 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x94 & ~x95;
assign c1155 =  x52;
assign c1157 = ~x60;
assign c1161 =  x3 &  x20 &  x26 &  x27 &  x36 &  x37 &  x48 &  x57 &  x58 &  x76 &  x78 &  x79 &  x88 & ~x4 & ~x22 & ~x25 & ~x34 & ~x35 & ~x53 & ~x55 & ~x65 & ~x74 & ~x83 & ~x85 & ~x92 & ~x93;
assign c1165 = ~x51;
assign c1167 = ~x71;
assign c1169 =  x1 &  x16 &  x17 &  x18 &  x19 &  x26 &  x28 &  x29 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x50 &  x57 &  x59 &  x66 &  x68 &  x70 &  x76 &  x78 &  x80 &  x86 &  x87 &  x88 &  x89 & ~x2 & ~x24 & ~x32 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x63 & ~x65 & ~x75 & ~x81 & ~x83 & ~x84 & ~x92 & ~x93 & ~x94 & ~x95;
assign c1171 =  x1 &  x19 &  x20 &  x37 &  x77 &  x86 & ~x5 & ~x24 & ~x33 & ~x34 & ~x45;
assign c1173 = ~x60;
assign c1175 = ~x30;
assign c1177 =  x16 &  x26 &  x46 &  x57 &  x76 & ~x75 & ~x84 & ~x85 & ~x91;
assign c1179 =  x52;
assign c1181 =  x0 &  x5 &  x26 &  x27 &  x78 & ~x24;
assign c1183 =  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x40 &  x46 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x2 & ~x23 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c1185 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x58 &  x59 &  x60 &  x61 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x88 &  x89 &  x90 &  x91 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c1187 =  x22;
assign c1191 =  x3 &  x17 &  x18 &  x19 &  x20 &  x27 &  x28 &  x37 &  x38 &  x47 &  x48 &  x56 &  x59 &  x69 &  x78 &  x79 &  x90 & ~x4 & ~x23 & ~x24 & ~x35 & ~x44 & ~x65 & ~x74 & ~x75 & ~x85 & ~x93;
assign c1193 =  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x4 & ~x22 & ~x23 & ~x24 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c1195 =  x72;
assign c1197 = ~x71;
assign c1199 =  x32;
assign c1201 =  x42;
assign c1203 =  x2 &  x16 &  x17 &  x19 &  x20 &  x26 &  x27 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x86 &  x88 & ~x3 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c1205 =  x92;
assign c1207 =  x3 &  x16 &  x17 &  x18 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x89 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x53 & ~x54 & ~x55 & ~x63 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x94 & ~x95;
assign c1209 = ~x31;
assign c1211 =  x36 &  x37 &  x38 &  x39 &  x48 &  x57 &  x78 &  x79 &  x81 &  x87 & ~x63;
assign c1213 = ~x51;
assign c1215 =  x36 &  x37 &  x66 &  x67 &  x70 &  x76 &  x77 &  x80 &  x81 &  x87 &  x88 & ~x45 & ~x64;
assign c1217 =  x2 &  x17 &  x56 &  x66 &  x67 &  x69 &  x76 &  x77 &  x79 &  x87 &  x89 & ~x23 & ~x65;
assign c1219 =  x72;
assign c1221 = ~x59;
assign c1223 =  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x22 & ~x23 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c1225 =  x82;
assign c1227 =  x2 &  x16 &  x17 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x68 &  x69 &  x76 &  x79 &  x86 &  x87 &  x88 & ~x5 & ~x23 & ~x24 & ~x25 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x84 & ~x85;
assign c1229 =  x16 &  x28 &  x57 &  x81 & ~x5 & ~x25;
assign c1231 =  x32;
assign c1233 =  x92;
assign c1235 =  x62;
assign c1237 =  x62;
assign c1239 =  x42;
assign c1241 = ~x20;
assign c1243 =  x4 &  x81;
assign c1245 =  x3 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c1247 =  x2 &  x17 &  x19 &  x20 &  x27 &  x28 &  x37 &  x38 &  x39 &  x40 &  x47 &  x48 &  x50 &  x57 &  x60 &  x66 &  x68 &  x69 &  x78 &  x79 &  x80 &  x86 &  x88 &  x89 & ~x5 & ~x23 & ~x25 & ~x35 & ~x45 & ~x54 & ~x73 & ~x75 & ~x82 & ~x83 & ~x95;
assign c1249 =  x0 &  x17 &  x27 &  x38 &  x47 &  x50 &  x59 &  x66 &  x76 &  x78 &  x87 &  x88 & ~x35 & ~x54 & ~x75 & ~x83 & ~x85 & ~x95;
assign c1251 =  x52;
assign c1253 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x40 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c1257 =  x72;
assign c1259 =  x2 &  x19 &  x27 &  x29 &  x37 &  x38 &  x39 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x67 &  x69 &  x70 &  x77 &  x78 &  x79 &  x80 &  x89 &  x90 & ~x1 & ~x23 & ~x25 & ~x32 & ~x33 & ~x35 & ~x44 & ~x52 & ~x53 & ~x55 & ~x63 & ~x72 & ~x73 & ~x75 & ~x83 & ~x93;
assign c1261 =  x3 &  x16 &  x27 &  x36 &  x40 &  x79 &  x88 & ~x4 & ~x24 & ~x25 & ~x42 & ~x83;
assign c1263 =  x0 &  x5 &  x26 &  x28 &  x46 &  x56 &  x66 &  x68 &  x86 & ~x34 & ~x54;
assign c1265 =  x52;
assign c1267 =  x32;
assign c1269 =  x3 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x50 &  x56 &  x57 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x76 &  x78 &  x79 &  x80 &  x86 &  x87 &  x90 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x95;
assign c1271 =  x0 &  x5 &  x27 &  x68 &  x69 & ~x24;
assign c1273 =  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c1275 =  x2 &  x17 &  x18 &  x19 &  x20 &  x26 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x80 &  x86 &  x88 &  x89 & ~x1 & ~x22 & ~x23 & ~x24 & ~x25 & ~x34 & ~x35 & ~x42 & ~x44 & ~x45 & ~x52 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93;
assign c1277 =  x27 &  x36 &  x46 &  x47 &  x49 &  x57 &  x58 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x81 &  x88 & ~x35 & ~x42 & ~x43 & ~x65;
assign c1279 =  x0 &  x6 &  x16 &  x17 &  x57 &  x66 &  x67 &  x76 & ~x35 & ~x64 & ~x65 & ~x75;
assign c1283 = ~x71;
assign c1285 =  x42;
assign c1287 = ~x51;
assign c1289 =  x1 &  x28 &  x56 &  x78 &  x80 &  x86 & ~x5 & ~x35 & ~x43;
assign c1291 =  x62;
assign c1293 =  x42;
assign c1295 =  x46 &  x76 & ~x21 & ~x24 & ~x33 & ~x35 & ~x75 & ~x83 & ~x84 & ~x91 & ~x95;
assign c1297 =  x3 &  x16 &  x17 &  x18 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x22 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x94 & ~x95;
assign c1299 =  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x28 &  x29 &  x36 &  x38 &  x47 &  x48 &  x49 &  x56 &  x57 &  x66 &  x67 &  x68 &  x76 &  x77 &  x86 &  x87 &  x88 &  x89 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x55 & ~x64 & ~x65 & ~x74 & ~x84 & ~x93 & ~x94 & ~x95;
assign c1301 =  x17 &  x26 &  x27 &  x36 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x68 &  x76 &  x87 &  x88 & ~x22 & ~x24 & ~x33 & ~x34 & ~x35 & ~x43 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x75 & ~x83 & ~x84 & ~x85 & ~x91 & ~x93 & ~x95;
assign c1303 =  x42;
assign c1307 = ~x20;
assign c1309 = ~x51;
assign c1311 = ~x80;
assign c1313 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c1315 =  x0 &  x4;
assign c1317 =  x32;
assign c1319 = ~x80;
assign c1321 =  x22;
assign c1323 = ~x71;
assign c1325 = ~x51;
assign c1327 =  x3 &  x17 &  x18 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x39 &  x40 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x89 & ~x2 & ~x22 & ~x23 & ~x24 & ~x34 & ~x35 & ~x43 & ~x45 & ~x52 & ~x53 & ~x55 & ~x62 & ~x63 & ~x64 & ~x73 & ~x75 & ~x82 & ~x83 & ~x84 & ~x92 & ~x94 & ~x95;
assign c1329 =  x32;
assign c1331 =  x72;
assign c1333 =  x92;
assign c1335 =  x1 &  x26 &  x58 &  x77 & ~x5 & ~x32 & ~x95;
assign c1337 =  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94;
assign c1341 =  x0 &  x6 &  x66 & ~x53;
assign c1343 =  x1 &  x27 &  x39 &  x47 &  x49 &  x58 &  x77 & ~x5 & ~x43 & ~x44;
assign c1345 = ~x60;
assign c1347 = ~x51;
assign c1349 =  x82;
assign c1351 = ~x60;
assign c1353 =  x2 &  x19 &  x20 &  x26 &  x27 &  x28 &  x30 &  x36 &  x37 &  x46 &  x49 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x68 &  x69 &  x70 &  x77 &  x78 &  x79 &  x87 &  x88 & ~x1 & ~x23 & ~x24 & ~x33 & ~x34 & ~x43 & ~x44 & ~x52 & ~x53 & ~x63 & ~x64 & ~x65 & ~x73 & ~x75 & ~x83 & ~x84 & ~x85 & ~x94 & ~x95;
assign c1355 =  x0 &  x17 &  x26 &  x28;
assign c1357 =  x92;
assign c1359 =  x3 &  x16 &  x18 &  x19 &  x29 &  x30 &  x31 &  x36 &  x38 &  x39 &  x40 &  x46 &  x48 &  x49 &  x50 &  x56 &  x58 &  x60 &  x66 &  x68 &  x76 &  x77 &  x78 &  x79 &  x80 &  x87 &  x89 &  x90 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x35 & ~x42 & ~x43 & ~x45 & ~x53 & ~x54 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x75 & ~x83 & ~x92 & ~x94 & ~x95;
assign c1361 =  x62;
assign c1363 =  x2 &  x17 &  x18 &  x20 &  x26 &  x27 &  x36 &  x37 &  x38 &  x40 &  x47 &  x48 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x67 &  x68 &  x69 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x22 & ~x23 & ~x24 & ~x34 & ~x35 & ~x45 & ~x52 & ~x53 & ~x54 & ~x62 & ~x63 & ~x64 & ~x72 & ~x83 & ~x84 & ~x92 & ~x93 & ~x94 & ~x95;
assign c1365 = ~x31;
assign c1367 =  x52;
assign c1369 =  x62;
assign c1371 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x36 &  x38 &  x39 &  x40 &  x46 &  x47 &  x49 &  x56 &  x58 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x86 &  x87 &  x89 &  x90 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x54 & ~x55 & ~x64 & ~x65 & ~x75 & ~x82 & ~x83 & ~x85 & ~x94 & ~x95;
assign c1373 =  x1 &  x19 &  x20 &  x26 &  x27 &  x28 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x50 &  x56 &  x58 &  x59 &  x79 &  x80 &  x88 &  x89 & ~x4 & ~x33 & ~x43 & ~x45 & ~x52 & ~x53 & ~x64 & ~x84;
assign c1375 =  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x28 &  x29 &  x37 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x58 &  x60 &  x66 &  x67 &  x69 &  x70 &  x77 &  x79 &  x80 &  x86 &  x89 &  x90 & ~x1 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x45 & ~x52 & ~x53 & ~x54 & ~x62 & ~x63 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c1377 = ~x71;
assign c1379 =  x6 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x48 &  x56 &  x57 &  x59 &  x66 &  x67 &  x69 &  x70 &  x71 &  x76 &  x77 &  x79 &  x87 &  x88 &  x89 &  x90 & ~x4 & ~x5 & ~x24 & ~x25 & ~x33 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c1381 =  x81 & ~x42;
assign c1383 =  x3 & ~x51;
assign c1385 =  x62;
assign c1387 =  x5 &  x16 &  x17 &  x18 &  x26 &  x36 &  x37 &  x56 &  x66 &  x67 &  x76 &  x86 &  x87 & ~x34 & ~x45 & ~x54 & ~x55 & ~x73 & ~x74 & ~x85;
assign c1389 =  x2 &  x16 &  x17 &  x18 &  x20 &  x26 &  x28 &  x30 &  x37 &  x39 &  x40 &  x46 &  x47 &  x48 &  x51 &  x56 &  x59 &  x60 &  x66 &  x67 &  x69 &  x70 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x22 & ~x23 & ~x25 & ~x35 & ~x42 & ~x44 & ~x45 & ~x62 & ~x64 & ~x65 & ~x72 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x94;
assign c1391 =  x0 &  x6 &  x30 &  x37 &  x47 &  x66 &  x86 &  x87 & ~x24;
assign c1393 =  x1 &  x26 &  x46 &  x48 &  x50 &  x57 &  x87 & ~x5 & ~x44 & ~x55;
assign c1395 =  x92;
assign c1397 =  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 & ~x3 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c1399 =  x16 &  x17 &  x18 &  x26 &  x27 &  x36 &  x37 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x68 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 & ~x23 & ~x25 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x91 & ~x92 & ~x93 & ~x94;
assign c1401 = ~x71;
assign c1403 = ~x51;
assign c1405 =  x82;
assign c1407 =  x3 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x56 &  x58 &  x67 &  x68 &  x69 &  x70 &  x76 &  x78 &  x86 &  x87 &  x88 &  x90 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x72 & ~x74 & ~x82 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c1409 = ~x90;
assign c1411 =  x16 &  x36 &  x39 &  x46 &  x66 &  x76 &  x86 & ~x21 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x64 & ~x65 & ~x84 & ~x91 & ~x92 & ~x93 & ~x94 & ~x95;
assign c1413 =  x0 &  x4 &  x26 &  x46 &  x58;
assign c1415 = ~x71;
assign c1417 =  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c1419 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c1421 =  x28 &  x36 &  x46 &  x66 &  x68 &  x79 &  x81 & ~x5 & ~x24 & ~x44 & ~x45;
assign c1425 =  x3 &  x19 &  x26 &  x27 &  x28 &  x29 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x50 &  x51 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x77 &  x80 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x22 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x72 & ~x73 & ~x75 & ~x84 & ~x85 & ~x93 & ~x95;
assign c1427 =  x0 &  x5 &  x27 &  x29 &  x36 &  x46 &  x47 &  x87 & ~x34 & ~x75 & ~x85 & ~x94;
assign c1429 =  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x89 & ~x1 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c1431 = ~x71;
assign c1433 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c1435 = ~x71;
assign c1437 =  x26 &  x27 &  x28 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x57 &  x58 &  x59 &  x66 &  x77 &  x86 &  x87 & ~x21 & ~x24 & ~x25 & ~x34 & ~x43 & ~x45 & ~x55 & ~x64 & ~x65 & ~x74 & ~x75 & ~x84 & ~x91 & ~x94;
assign c1439 =  x2 &  x16 &  x18 &  x19 &  x27 &  x28 &  x36 &  x39 &  x40 &  x46 &  x47 &  x49 &  x50 &  x56 &  x58 &  x59 &  x66 &  x68 &  x69 &  x71 &  x76 &  x78 &  x86 &  x87 &  x88 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x74 & ~x83 & ~x84 & ~x85 & ~x93 & ~x95;
assign c1441 =  x2 &  x16 &  x17 &  x18 &  x27 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x48 &  x49 &  x51 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x70 &  x76 &  x77 &  x78 &  x86 &  x87 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x52 & ~x53 & ~x55 & ~x62 & ~x63 & ~x64 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x95;
assign c1443 = ~x60;
assign c1445 =  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x60 &  x66 &  x67 &  x68 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x72 & ~x73 & ~x75 & ~x82 & ~x83 & ~x85 & ~x93 & ~x94 & ~x95;
assign c1447 = ~x51;
assign c1449 =  x19 &  x27 &  x46 &  x66 &  x68 &  x76 &  x78 &  x81 &  x88 &  x89;
assign c1451 =  x0 &  x4 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x66 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x89 &  x90 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x64 & ~x65 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c1453 =  x32;
assign c1455 =  x0 &  x4;
assign c1457 =  x4 &  x68 &  x81 & ~x42;
assign c1459 = ~x71;
assign c1461 =  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x86 &  x87 &  x88 &  x89 & ~x3 & ~x23 & ~x24 & ~x25 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c1463 = ~x51;
assign c1465 =  x52;
assign c1467 =  x2 &  x16 &  x17 &  x18 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x76 &  x78 &  x80 &  x86 &  x87 &  x88 &  x90 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x85 & ~x93 & ~x95;
assign c1469 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x2 & ~x22 & ~x23 & ~x32 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c1471 =  x3 &  x16 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x38 &  x39 &  x47 &  x49 &  x57 &  x59 &  x60 &  x66 &  x67 &  x76 &  x77 &  x78 &  x79 &  x87 &  x88 & ~x5 & ~x24 & ~x25 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x65 & ~x72 & ~x73 & ~x75 & ~x85 & ~x93 & ~x94;
assign c1473 =  x0 &  x16 &  x17 &  x26 &  x56 &  x69 &  x87 &  x90 & ~x73 & ~x74 & ~x75;
assign c1475 =  x32;
assign c1477 =  x52;
assign c1479 =  x62;
assign c1483 =  x92;
assign c1485 =  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x28 &  x29 &  x30 &  x37 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x60 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x80 &  x87 &  x88 &  x90 & ~x1 & ~x22 & ~x23 & ~x24 & ~x25 & ~x34 & ~x35 & ~x43 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x82 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94;
assign c1487 = ~x51;
assign c1489 =  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c1491 =  x22;
assign c1493 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x88 &  x89 &  x90 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c1495 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 & ~x3 & ~x22 & ~x23 & ~x24 & ~x32 & ~x33 & ~x34 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x81 & ~x82 & ~x83 & ~x84 & ~x92 & ~x93 & ~x94 & ~x95;
assign c1497 =  x2 &  x18 &  x27 &  x28 &  x29 &  x36 &  x38 &  x40 &  x47 &  x48 &  x56 &  x57 &  x58 &  x59 &  x66 &  x68 &  x69 &  x76 &  x86 &  x88 &  x89 & ~x5 & ~x23 & ~x24 & ~x25 & ~x33 & ~x42 & ~x43 & ~x44 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x94 & ~x95;
assign c1499 =  x1 &  x20 &  x26 &  x27 &  x30 &  x37 &  x38 &  x48 &  x49 &  x56 &  x67 &  x76 &  x77 &  x78 & ~x5 & ~x22 & ~x25 & ~x32 & ~x33 & ~x43 & ~x52 & ~x53 & ~x54 & ~x55 & ~x64;
assign c20 =  x45 &  x65 & ~x68;
assign c22 = ~x90;
assign c24 = ~x36;
assign c26 =  x22 &  x61;
assign c28 = ~x37;
assign c210 =  x92;
assign c212 =  x92 & ~x0;
assign c216 =  x53;
assign c220 =  x35;
assign c222 =  x5 &  x16 &  x17 &  x20 &  x26 &  x27 &  x28 &  x36 &  x37 &  x38 &  x46 &  x47 &  x56 &  x66 &  x67 &  x77 &  x89 & ~x1 & ~x2 & ~x25 & ~x35 & ~x43 & ~x44 & ~x51 & ~x53 & ~x54 & ~x62 & ~x63 & ~x73 & ~x74 & ~x84 & ~x93 & ~x94;
assign c224 =  x93;
assign c226 = ~x37;
assign c228 = ~x59;
assign c230 = ~x16;
assign c232 = ~x56;
assign c234 = ~x18;
assign c238 = ~x68;
assign c240 =  x17 &  x18 &  x19 &  x20 &  x26 &  x28 &  x29 &  x30 &  x36 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x2 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x55 & ~x62 & ~x63 & ~x64 & ~x72 & ~x73 & ~x75 & ~x80 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x95;
assign c242 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x2 & ~x21 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x91 & ~x92 & ~x93 & ~x94 & ~x95;
assign c244 =  x0 &  x4 &  x16 &  x17 &  x18 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x2 & ~x3 & ~x21 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x91 & ~x92 & ~x93 & ~x94 & ~x95;
assign c246 =  x35;
assign c248 = ~x78;
assign c250 = ~x76;
assign c252 = ~x56;
assign c254 = ~x26;
assign c256 = ~x76;
assign c258 =  x53;
assign c260 = ~x26 & ~x88;
assign c262 = ~x56 & ~x68;
assign c264 = ~x38;
assign c266 = ~x26;
assign c268 =  x0 &  x4 &  x5 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x46 &  x47 &  x48 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x2 & ~x3 & ~x6 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c270 =  x3 &  x16 &  x17 &  x18 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x38 &  x39 &  x40 &  x41 &  x46 &  x48 &  x49 &  x50 &  x56 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x70 &  x76 &  x77 &  x78 &  x80 &  x81 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x75 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c272 =  x85;
assign c274 = ~x66;
assign c276 =  x8 &  x16 &  x20 &  x31 &  x37 &  x46 &  x47 &  x69 &  x76 &  x90 & ~x1 & ~x2 & ~x24 & ~x25 & ~x42 & ~x45 & ~x51;
assign c278 =  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x30 &  x36 &  x37 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x59 &  x60 &  x61 &  x66 &  x67 &  x68 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x2 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x51 & ~x52 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c282 = ~x27 & ~x77;
assign c284 =  x5 &  x17 &  x30 &  x36 &  x38 &  x39 &  x47 &  x57 &  x59 &  x79 &  x88 &  x89 & ~x1 & ~x2 & ~x42 & ~x43 & ~x44 & ~x51 & ~x52 & ~x54 & ~x64 & ~x65 & ~x73 & ~x75;
assign c286 = ~x27;
assign c288 =  x5 &  x17 &  x49 &  x52 & ~x23 & ~x24 & ~x55 & ~x72 & ~x74 & ~x94;
assign c290 = ~x56;
assign c292 =  x5 & ~x50;
assign c294 = ~x76;
assign c296 =  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x0 & ~x1 & ~x2 & ~x9 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c298 =  x0 &  x4 &  x6 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x2 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2100 =  x45;
assign c2104 = ~x76;
assign c2106 =  x5 &  x19 &  x26 &  x37 &  x47 &  x48 &  x49 &  x50 &  x51 &  x52 &  x60 &  x78 &  x86 &  x87 &  x88 &  x90 & ~x1 & ~x2 & ~x64;
assign c2108 = ~x36 & ~x46;
assign c2110 =  x0 &  x4 &  x16 &  x17 &  x19 &  x26 &  x27 &  x28 &  x30 &  x36 &  x37 &  x46 &  x48 &  x57 &  x66 &  x67 &  x76 &  x86 & ~x3 & ~x23 & ~x32 & ~x33 & ~x45 & ~x53 & ~x74 & ~x82 & ~x83 & ~x84 & ~x91 & ~x95;
assign c2112 =  x5 &  x41 &  x53;
assign c2114 =  x92 & ~x0;
assign c2116 =  x5 &  x17 &  x28 &  x29 &  x31 &  x36 &  x37 &  x38 &  x40 &  x46 &  x47 &  x48 &  x49 &  x59 &  x60 &  x66 &  x67 &  x68 &  x76 &  x78 &  x86 &  x87 &  x88 &  x90 & ~x1 & ~x7 & ~x21 & ~x22 & ~x23 & ~x24 & ~x33 & ~x35 & ~x45 & ~x62 & ~x63 & ~x72 & ~x73 & ~x84 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2118 =  x4 &  x16 &  x17 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x56 &  x57 &  x58 &  x59 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x2 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x51 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x84 & ~x85 & ~x93 & ~x94;
assign c2122 = ~x48 & ~x60;
assign c2124 =  x55;
assign c2126 =  x22;
assign c2128 =  x45;
assign c2130 = ~x67;
assign c2132 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x2 & ~x21 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x91 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2134 = ~x57;
assign c2136 = ~x66;
assign c2138 = ~x56;
assign c2140 = ~x86;
assign c2142 =  x85;
assign c2144 =  x3 &  x5 &  x16 &  x17 &  x18 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x57 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x86 &  x87 &  x88 &  x89 & ~x0 & ~x1 & ~x2 & ~x4 & ~x21 & ~x22 & ~x23 & ~x25 & ~x32 & ~x33 & ~x35 & ~x44 & ~x54 & ~x55 & ~x63 & ~x64 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2146 = ~x68;
assign c2148 = ~x38;
assign c2150 = ~x26;
assign c2152 = ~x58;
assign c2154 = ~x78;
assign c2158 = ~x40;
assign c2160 = ~x38;
assign c2162 =  x3 &  x5 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x2 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c2164 =  x55;
assign c2166 = ~x67;
assign c2168 =  x3 &  x5 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x67 &  x68 &  x69 &  x70 &  x77 &  x78 &  x86 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x2 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x95;
assign c2170 =  x22 &  x61;
assign c2172 =  x84;
assign c2174 = ~x46;
assign c2176 = ~x76;
assign c2178 =  x85 & ~x88;
assign c2180 =  x3 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x2 & ~x21 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2182 =  x35;
assign c2184 =  x67 & ~x0 & ~x35 & ~x45 & ~x62 & ~x80;
assign c2186 = ~x26;
assign c2188 =  x4 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x2 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x51 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2190 = ~x48;
assign c2192 = ~x90;
assign c2194 = ~x79;
assign c2196 = ~x5 & ~x90;
assign c2198 = ~x66;
assign c2200 = ~x48;
assign c2202 =  x22;
assign c2204 =  x3 &  x5 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x2 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c2206 = ~x38;
assign c2208 =  x35;
assign c2210 = ~x19;
assign c2212 =  x54;
assign c2214 =  x16 &  x17 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x36 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x50 &  x56 &  x57 &  x58 &  x60 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x80 &  x86 &  x87 &  x88 &  x90 & ~x1 & ~x2 & ~x22 & ~x24 & ~x32 & ~x33 & ~x42 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x62 & ~x64 & ~x65 & ~x71 & ~x72 & ~x73 & ~x74 & ~x84 & ~x85 & ~x92 & ~x93 & ~x95;
assign c2216 =  x5 &  x17 &  x38 &  x39 &  x47 &  x49 &  x51 &  x52 &  x56 &  x57 &  x59 &  x60 &  x68 &  x70 &  x78 &  x87 & ~x1 & ~x2 & ~x34 & ~x44 & ~x45 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x93;
assign c2218 =  x63;
assign c2220 = ~x86;
assign c2222 = ~x38;
assign c2224 = ~x76;
assign c2226 =  x17 &  x18 &  x27 &  x29 &  x39 &  x48 &  x49 &  x56 &  x57 &  x76 &  x86 &  x89 & ~x0 & ~x2 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x65 & ~x80 & ~x81 & ~x84 & ~x93;
assign c2228 = ~x56;
assign c2230 =  x35;
assign c2232 = ~x76;
assign c2234 =  x7 &  x16 &  x19 &  x20 &  x31 &  x36 &  x38 &  x39 &  x40 &  x41 &  x42 &  x46 &  x47 &  x51 &  x56 &  x58 &  x59 &  x60 &  x66 &  x69 &  x70 &  x87 &  x88 &  x90 & ~x2 & ~x24 & ~x25 & ~x33 & ~x35 & ~x43 & ~x44 & ~x64 & ~x73 & ~x84 & ~x85 & ~x94;
assign c2236 = ~x86;
assign c2238 =  x3 &  x5 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x2 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c2240 =  x35;
assign c2242 = ~x56;
assign c2244 = ~x46;
assign c2246 =  x83;
assign c2248 = ~x78;
assign c2250 =  x55;
assign c2252 =  x52 & ~x21 & ~x54 & ~x95;
assign c2254 =  x82 & ~x0;
assign c2256 =  x0 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x2 & ~x3 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2258 = ~x36 & ~x87;
assign c2260 = ~x66;
assign c2262 =  x55;
assign c2264 = ~x26;
assign c2266 = ~x38;
assign c2268 =  x95;
assign c2270 = ~x36;
assign c2272 =  x45;
assign c2274 = ~x38;
assign c2276 =  x0 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x2 & ~x3 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2278 =  x5 &  x38 &  x52 &  x77 & ~x1 & ~x2 & ~x43 & ~x64;
assign c2280 =  x5 &  x16 &  x17 &  x28 &  x29 &  x37 &  x47 &  x49 &  x50 &  x52 &  x59 &  x60 &  x68 &  x69 &  x70 &  x77 &  x79 &  x88 &  x89 & ~x1 & ~x2 & ~x25 & ~x33 & ~x34 & ~x44 & ~x55 & ~x64 & ~x95;
assign c2282 = ~x70;
assign c2286 =  x3 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x0 & ~x1 & ~x2 & ~x5 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2288 =  x7 &  x20 &  x21 &  x42 &  x70 &  x89 & ~x1 & ~x43 & ~x72;
assign c2290 =  x4 &  x19 &  x29 &  x30 &  x37 &  x46 &  x49 &  x51 & ~x2 & ~x23 & ~x24 & ~x32 & ~x33 & ~x45 & ~x75 & ~x80 & ~x81 & ~x94;
assign c2292 = ~x36;
assign c2294 =  x5 & ~x50;
assign c2296 = ~x66;
assign c2298 = ~x37;
assign c2300 =  x65;
assign c2302 =  x31 &  x41 &  x82 & ~x94;
assign c2304 =  x95;
assign c2306 = ~x27;
assign c2308 = ~x27;
assign c2310 =  x5 &  x16 &  x27 &  x37 &  x48 &  x70 &  x76 &  x90 & ~x1 & ~x24 & ~x51 & ~x54 & ~x62 & ~x63 & ~x85 & ~x95;
assign c2312 =  x4 &  x16 &  x17 &  x18 &  x19 &  x26 &  x29 &  x30 &  x36 &  x37 &  x38 &  x46 &  x47 &  x57 &  x66 &  x67 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x89 &  x90 & ~x2 & ~x23 & ~x25 & ~x32 & ~x33 & ~x42 & ~x43 & ~x44 & ~x45 & ~x51 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x84 & ~x93 & ~x94 & ~x95;
assign c2314 =  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x2 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x80 & ~x82 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c2316 = ~x46;
assign c2318 =  x17 &  x18 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x38 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x67 &  x68 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x35 & ~x44 & ~x45 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x80 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x95;
assign c2320 =  x0 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x2 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x61 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2322 =  x20 &  x26 &  x31 &  x37 &  x47 &  x58 &  x69 & ~x2 & ~x50;
assign c2324 =  x3 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x0 & ~x1 & ~x2 & ~x5 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c2328 = ~x28;
assign c2330 =  x65;
assign c2332 =  x75;
assign c2334 =  x16 &  x17 &  x18 &  x28 &  x30 &  x31 &  x36 &  x37 &  x47 &  x57 &  x58 &  x66 &  x67 &  x70 &  x71 &  x76 &  x78 &  x79 &  x80 & ~x25 & ~x32 & ~x33 & ~x34 & ~x42 & ~x44 & ~x45 & ~x51 & ~x74 & ~x75 & ~x82 & ~x93;
assign c2336 = ~x86;
assign c2338 =  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x80 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2340 =  x5 &  x28 &  x30 &  x31 &  x36 &  x39 &  x47 &  x48 &  x56 &  x58 &  x67 &  x71 &  x79 &  x81 &  x89 & ~x8 & ~x25 & ~x33 & ~x34 & ~x44 & ~x45 & ~x83 & ~x85 & ~x92 & ~x93 & ~x94;
assign c2342 =  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x47 &  x48 &  x49 &  x50 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x77 &  x79 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x0 & ~x9 & ~x23 & ~x25 & ~x35 & ~x43 & ~x44 & ~x52 & ~x53 & ~x54 & ~x63 & ~x64 & ~x73 & ~x75 & ~x83 & ~x84 & ~x93 & ~x94 & ~x95;
assign c2344 = ~x86;
assign c2346 =  x64;
assign c2348 = ~x16;
assign c2350 =  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x79 &  x80 &  x81 &  x87 &  x88 &  x89 & ~x2 & ~x21 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c2352 =  x5 &  x52 &  x68 &  x79 &  x88 & ~x1 & ~x63 & ~x64 & ~x73;
assign c2354 =  x45;
assign c2356 =  x4 &  x17 &  x20 &  x30 &  x31 &  x36 &  x40 &  x41 &  x42 &  x46 &  x47 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x67 &  x68 &  x70 &  x76 &  x77 &  x79 &  x87 &  x88 &  x89 & ~x1 & ~x2 & ~x5 & ~x25 & ~x33 & ~x35 & ~x44 & ~x45 & ~x63 & ~x65 & ~x75 & ~x85 & ~x94 & ~x95;
assign c2358 =  x0 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x2 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x61 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2362 = ~x66;
assign c2364 =  x0 &  x4 &  x16 &  x17 &  x18 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x37 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x2 & ~x3 & ~x11 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x75 & ~x82 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2366 =  x42 &  x71;
assign c2368 = ~x56;
assign c2370 = ~x76;
assign c2372 = ~x90;
assign c2374 =  x35;
assign c2376 =  x0 &  x4 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x2 & ~x3 & ~x21 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x91 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2378 =  x5 &  x18 &  x50 &  x52 &  x59 &  x76 &  x77 &  x78 &  x86 &  x87 &  x89 & ~x1 & ~x44 & ~x63 & ~x65 & ~x85 & ~x93;
assign c2380 = ~x88;
assign c2382 =  x83;
assign c2384 =  x4 &  x19 &  x26 &  x28 &  x29 &  x31 &  x37 &  x39 &  x49 &  x56 &  x57 &  x59 &  x60 &  x66 &  x70 &  x71 &  x76 &  x77 &  x80 &  x86 &  x87 &  x88 & ~x1 & ~x2 & ~x25 & ~x33 & ~x35 & ~x44 & ~x45 & ~x51 & ~x52 & ~x53 & ~x62 & ~x64 & ~x73 & ~x74 & ~x75 & ~x84 & ~x85 & ~x95;
assign c2386 =  x4 &  x17 &  x19 &  x20 &  x21 &  x29 &  x36 &  x37 &  x38 &  x39 &  x49 &  x56 &  x66 &  x67 &  x68 &  x69 &  x70 &  x77 &  x78 &  x87 &  x88 & ~x2 & ~x23 & ~x25 & ~x34 & ~x44 & ~x51 & ~x52 & ~x62 & ~x65 & ~x72 & ~x73 & ~x75 & ~x83 & ~x85 & ~x93 & ~x94;
assign c2388 =  x3 &  x5 &  x16 &  x17 &  x18 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x2 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2390 = ~x56;
assign c2392 =  x41 &  x53;
assign c2394 = ~x57;
assign c2396 = ~x86;
assign c2398 =  x16 &  x18 &  x26 &  x29 &  x46 &  x56 &  x57 &  x58 &  x69 &  x76 &  x77 &  x87 &  x88 &  x89 & ~x1 & ~x24 & ~x25 & ~x33 & ~x35 & ~x42 & ~x43 & ~x51 & ~x52 & ~x54 & ~x62 & ~x63 & ~x64 & ~x75 & ~x82 & ~x85 & ~x91 & ~x92 & ~x93 & ~x95;
assign c2400 =  x3 &  x5 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x2 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2402 = ~x86;
assign c2404 =  x5 &  x39 &  x52 &  x56 &  x57 &  x59 &  x78 & ~x1 & ~x2 & ~x44 & ~x63 & ~x64 & ~x83 & ~x93;
assign c2408 =  x0 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x2 & ~x3 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2410 =  x41 &  x53;
assign c2412 =  x5 &  x53;
assign c2414 =  x75;
assign c2416 =  x5 &  x16 &  x17 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x2 & ~x24 & ~x25 & ~x34 & ~x35 & ~x43 & ~x45 & ~x51 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c2418 = ~x66;
assign c2420 =  x55;
assign c2422 = ~x38;
assign c2424 =  x7 &  x20 &  x21 &  x26 &  x42 &  x70 &  x77 & ~x33;
assign c2426 =  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 & ~x0 & ~x1 & ~x2 & ~x5 & ~x7 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2428 =  x16 &  x17 &  x18 &  x19 &  x27 &  x28 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x50 &  x51 &  x56 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x2 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x74 & ~x75 & ~x80 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c2430 =  x5 &  x16 &  x26 &  x27 &  x28 &  x29 &  x30 &  x38 &  x47 &  x58 &  x60 &  x67 &  x68 &  x70 &  x76 &  x79 &  x89 & ~x1 & ~x2 & ~x34 & ~x35 & ~x51 & ~x52 & ~x53 & ~x55 & ~x62 & ~x64 & ~x65 & ~x73 & ~x83 & ~x93 & ~x95;
assign c2432 = ~x48;
assign c2434 = ~x78;
assign c2436 =  x83;
assign c2438 =  x6 &  x16 &  x17 &  x19 &  x28 &  x30 &  x31 &  x39 &  x40 &  x47 &  x49 &  x50 &  x56 &  x58 &  x59 &  x60 &  x66 &  x68 &  x69 &  x70 &  x76 &  x77 &  x86 &  x88 & ~x2 & ~x8 & ~x10 & ~x23 & ~x24 & ~x32 & ~x33 & ~x34 & ~x35 & ~x54 & ~x55 & ~x64 & ~x65 & ~x73 & ~x74 & ~x92 & ~x93 & ~x95;
assign c2440 = ~x27;
assign c2442 =  x5 &  x39 &  x41 &  x48 &  x50 &  x52 &  x56 &  x57 &  x59 &  x60 &  x68 &  x78 &  x86 &  x87 & ~x1 & ~x2 & ~x35 & ~x44 & ~x45 & ~x64 & ~x75 & ~x93;
assign c2444 =  x3 &  x16 &  x17 &  x19 &  x26 &  x28 &  x36 &  x56 &  x68 &  x69 &  x77 &  x87 &  x88 &  x89 & ~x0 & ~x1 & ~x6 & ~x21 & ~x35 & ~x44 & ~x45 & ~x63 & ~x64 & ~x72 & ~x83 & ~x84 & ~x85 & ~x91 & ~x93;
assign c2446 =  x0 &  x4 &  x17 &  x26 &  x28 &  x30 &  x38 &  x40 &  x46 &  x47 &  x49 &  x56 &  x58 &  x67 &  x69 &  x70 &  x78 &  x89 & ~x1 & ~x2 & ~x3 & ~x24 & ~x32 & ~x33 & ~x35 & ~x41 & ~x43 & ~x52 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x74 & ~x82 & ~x95;
assign c2448 =  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x88 &  x89 & ~x1 & ~x2 & ~x21 & ~x22 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x91 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2450 = ~x66;
assign c2452 =  x0 &  x4 &  x5 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x2 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2456 =  x16 &  x17 &  x18 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x80 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2458 =  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x69 &  x70 &  x76 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x2 & ~x21 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x85 & ~x91 & ~x92 & ~x93 & ~x94;
assign c2462 = ~x77;
assign c2464 =  x35 & ~x47;
assign c2466 = ~x38;
assign c2468 =  x3 &  x10 &  x16 &  x19 &  x20 &  x28 &  x36 &  x37 &  x40 &  x46 &  x47 &  x48 &  x58 &  x66 &  x78 &  x86 &  x87 &  x88 &  x90 & ~x0 & ~x1 & ~x2 & ~x9 & ~x22 & ~x23 & ~x24 & ~x25 & ~x35 & ~x42 & ~x44 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x74 & ~x83 & ~x84 & ~x92 & ~x94;
assign c2470 =  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x2 & ~x21 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x91 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2472 =  x55;
assign c2474 =  x3 &  x5 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x2 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c2476 =  x4 &  x10 &  x16 &  x17 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x48 &  x49 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x2 & ~x23 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x41 & ~x42 & ~x43 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2478 = ~x38;
assign c2480 =  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x81 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x2 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c2482 =  x92;
assign c2484 = ~x56;
assign c2486 =  x0 &  x4 &  x15 &  x16 &  x17 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x48 &  x56 &  x57 &  x58 &  x60 &  x66 &  x67 &  x70 &  x76 &  x77 &  x89 &  x90 & ~x2 & ~x3 & ~x22 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x52 & ~x54 & ~x55 & ~x62 & ~x63 & ~x65 & ~x73 & ~x74 & ~x83 & ~x84 & ~x85 & ~x92 & ~x94 & ~x95;
assign c2488 =  x0 &  x4 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x2 & ~x3 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2490 =  x8 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x46 &  x47 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x2 & ~x23 & ~x24 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x51 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x73 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c2492 = ~x28;
assign c2494 =  x4 &  x16 &  x17 &  x27 &  x28 &  x30 &  x59 &  x67 &  x70 &  x71 &  x77 &  x78 &  x80 &  x87 &  x88 &  x90 & ~x1 & ~x2 & ~x23 & ~x24 & ~x32 & ~x33 & ~x43 & ~x44 & ~x45 & ~x51 & ~x52 & ~x53 & ~x54 & ~x55 & ~x65 & ~x73 & ~x74 & ~x75 & ~x93 & ~x95;
assign c2496 =  x3 &  x5 &  x16 &  x26 &  x27 &  x28 &  x29 &  x30 &  x37 &  x39 &  x41 &  x46 &  x47 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x70 &  x76 &  x78 &  x79 &  x86 &  x88 &  x89 & ~x0 & ~x1 & ~x4 & ~x22 & ~x23 & ~x24 & ~x33 & ~x35 & ~x44 & ~x54 & ~x62 & ~x64 & ~x65 & ~x73 & ~x74 & ~x84 & ~x85 & ~x92 & ~x94 & ~x95;
assign c2498 = ~x77;
assign c21 =  x1;
assign c23 =  x2;
assign c25 =  x44;
assign c27 =  x1;
assign c29 =  x0 &  x3 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 & ~x1 & ~x24 & ~x25 & ~x34 & ~x35 & ~x43 & ~x44 & ~x53 & ~x54 & ~x55 & ~x62 & ~x64 & ~x65 & ~x73 & ~x75 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c211 =  x2;
assign c213 =  x1;
assign c215 =  x0 &  x3 &  x16 &  x17 &  x19 &  x26 &  x28 &  x29 &  x36 &  x37 &  x38 &  x40 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x78 &  x79 &  x86 &  x87 &  x88 & ~x1 & ~x2 & ~x24 & ~x25 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x55 & ~x62 & ~x63 & ~x64 & ~x72 & ~x73 & ~x75 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c217 =  x4 &  x5 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x0 & ~x1 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c219 = ~x89;
assign c221 =  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x0 & ~x1 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c223 =  x63;
assign c225 =  x33;
assign c227 =  x1;
assign c229 = ~x30;
assign c233 =  x62;
assign c235 = ~x18;
assign c237 = ~x69;
assign c239 =  x9 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x29 &  x30 &  x36 &  x38 &  x39 &  x40 &  x41 &  x46 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x67 &  x69 &  x78 &  x80 &  x86 &  x87 &  x88 &  x89 &  x91 & ~x1 & ~x2 & ~x22 & ~x23 & ~x25 & ~x32 & ~x33 & ~x35 & ~x43 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x82 & ~x92 & ~x93 & ~x94 & ~x95;
assign c241 =  x18 &  x19 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x59 &  x66 &  x67 &  x68 &  x76 &  x79 &  x88 &  x89 &  x90 & ~x2 & ~x3 & ~x4 & ~x24 & ~x25 & ~x32 & ~x33 & ~x35 & ~x42 & ~x44 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c243 =  x62;
assign c245 =  x24;
assign c247 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x70 &  x71 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x1 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c249 = ~x89;
assign c251 =  x2;
assign c253 =  x18 &  x20 &  x26 &  x28 &  x30 &  x31 &  x46 &  x47 &  x48 &  x49 &  x51 &  x56 &  x57 &  x58 &  x60 &  x67 &  x68 &  x79 &  x87 &  x90 & ~x0 & ~x3 & ~x22 & ~x23 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x53 & ~x55 & ~x62 & ~x63 & ~x73 & ~x74 & ~x75 & ~x82 & ~x84 & ~x95;
assign c255 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x1 & ~x2 & ~x10 & ~x22 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c257 =  x4 &  x5 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c259 =  x3 &  x4 &  x7 &  x16 &  x17 &  x18 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x47 &  x48 &  x58 &  x60 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x22 & ~x25 & ~x33 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x62 & ~x64 & ~x65 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94;
assign c261 =  x16 &  x18 &  x19 &  x26 &  x27 &  x28 &  x30 &  x36 &  x37 &  x39 &  x40 &  x48 &  x49 &  x56 &  x57 &  x58 &  x67 &  x68 &  x70 &  x78 &  x80 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x4 & ~x5 & ~x24 & ~x25 & ~x34 & ~x43 & ~x44 & ~x55 & ~x63 & ~x64 & ~x74 & ~x85 & ~x92 & ~x93 & ~x95;
assign c263 =  x16 &  x17 &  x19 &  x20 &  x26 &  x27 &  x28 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x77 &  x78 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x2 & ~x3 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x54 & ~x55 & ~x62 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c265 =  x93;
assign c267 =  x17 &  x26 &  x27 &  x29 &  x36 &  x38 &  x47 &  x48 &  x60 &  x66 &  x68 &  x70 &  x71 &  x77 &  x80 &  x86 &  x89 & ~x0 & ~x1 & ~x3 & ~x22 & ~x23 & ~x24 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x45 & ~x55 & ~x62 & ~x64 & ~x72 & ~x74 & ~x75 & ~x83 & ~x93;
assign c269 =  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x37 &  x38 &  x46 &  x47 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x69 &  x70 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x90 & ~x2 & ~x3 & ~x4 & ~x22 & ~x23 & ~x24 & ~x32 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c271 =  x1;
assign c273 = ~x89;
assign c275 =  x1;
assign c277 =  x17 &  x20 &  x27 &  x28 &  x30 &  x36 &  x39 &  x46 &  x47 &  x49 &  x56 &  x58 &  x67 &  x68 &  x70 &  x71 &  x76 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x52 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x82 & ~x92 & ~x93 & ~x95;
assign c279 =  x2;
assign c281 =  x1;
assign c283 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x48 &  x49 &  x50 &  x56 &  x58 &  x59 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x3 & ~x4 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x94 & ~x95;
assign c285 =  x0 &  x3 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x30 &  x36 &  x37 &  x38 &  x46 &  x47 &  x48 &  x50 &  x56 &  x57 &  x58 &  x60 &  x66 &  x67 &  x68 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x2 & ~x23 & ~x24 & ~x25 & ~x35 & ~x43 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x93 & ~x95;
assign c287 = ~x89;
assign c289 =  x32;
assign c291 =  x1;
assign c293 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c295 =  x62;
assign c297 =  x0 &  x17 &  x27 &  x29 &  x30 &  x37 &  x48 &  x57 &  x60 &  x66 &  x67 &  x68 &  x69 &  x77 &  x80 & ~x1 & ~x2 & ~x4 & ~x25 & ~x34 & ~x35 & ~x44 & ~x45 & ~x63 & ~x65 & ~x73 & ~x74 & ~x75 & ~x84 & ~x85 & ~x94 & ~x95;
assign c2101 =  x3 &  x32;
assign c2103 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x36 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x59 &  x67 &  x68 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x2 & ~x3 & ~x4 & ~x24 & ~x33 & ~x34 & ~x35 & ~x45 & ~x55 & ~x65 & ~x73 & ~x74 & ~x75 & ~x84 & ~x95;
assign c2105 =  x2;
assign c2107 =  x1;
assign c2109 =  x0 &  x3 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x36 &  x37 &  x38 &  x39 &  x40 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x60 &  x66 &  x67 &  x68 &  x70 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x2 & ~x24 & ~x25 & ~x34 & ~x35 & ~x43 & ~x44 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x85 & ~x94 & ~x95;
assign c2111 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x1 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2113 =  x0 &  x3 &  x16 &  x17 &  x26 &  x27 &  x28 &  x29 &  x36 &  x37 &  x38 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x86 &  x87 & ~x1 & ~x2 & ~x24 & ~x25 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x84 & ~x85 & ~x95;
assign c2115 =  x2;
assign c2117 =  x17 &  x18 &  x19 &  x20 &  x27 &  x30 &  x36 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x57 &  x58 &  x66 &  x67 &  x69 &  x87 &  x90 & ~x4 & ~x5 & ~x22 & ~x25 & ~x32 & ~x33 & ~x43 & ~x44 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x82 & ~x84 & ~x92 & ~x93 & ~x94;
assign c2119 =  x24;
assign c2121 =  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x68 &  x76 &  x88 &  x89 &  x90 & ~x2 & ~x3 & ~x4 & ~x22 & ~x23 & ~x24 & ~x34 & ~x35 & ~x44 & ~x53 & ~x62 & ~x63 & ~x65 & ~x73 & ~x74 & ~x75 & ~x84 & ~x85 & ~x92 & ~x94 & ~x95;
assign c2123 =  x2;
assign c2125 =  x0 &  x3 &  x16 &  x17 &  x18 &  x19 &  x27 &  x30 &  x38 &  x39 &  x40 &  x46 &  x49 &  x50 &  x51 &  x57 &  x58 &  x59 &  x67 &  x68 &  x69 &  x76 &  x86 & ~x1 & ~x2 & ~x24 & ~x35 & ~x53 & ~x55 & ~x64 & ~x65 & ~x75 & ~x84 & ~x85 & ~x93 & ~x95;
assign c2127 = ~x69;
assign c2129 = ~x89;
assign c2131 = ~x89;
assign c2133 =  x25;
assign c2135 =  x2;
assign c2137 =  x54;
assign c2139 =  x24;
assign c2141 =  x4 &  x7 &  x26 &  x27 &  x28 &  x29 &  x30 &  x39 &  x46 &  x47 &  x48 &  x50 &  x51 &  x59 &  x60 &  x68 &  x69 &  x77 &  x78 &  x79 &  x80 &  x88 & ~x0 & ~x25 & ~x34 & ~x35 & ~x42 & ~x43 & ~x54 & ~x63 & ~x74 & ~x82 & ~x92;
assign c2143 = ~x89;
assign c2145 = ~x89;
assign c2147 =  x0 &  x16 &  x17 &  x19 &  x26 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x46 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x76 &  x78 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x4 & ~x24 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x63 & ~x65 & ~x73 & ~x75 & ~x83 & ~x84 & ~x93 & ~x94 & ~x95;
assign c2149 =  x17 &  x18 &  x26 &  x27 &  x30 &  x36 &  x46 &  x47 &  x48 &  x50 &  x56 &  x57 &  x58 &  x59 &  x68 &  x76 &  x86 &  x87 &  x90 &  x91 & ~x2 & ~x3 & ~x4 & ~x24 & ~x34 & ~x53 & ~x55 & ~x63 & ~x64 & ~x73 & ~x75 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c2151 =  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x68 &  x69 &  x76 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x4 & ~x5 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x44 & ~x54 & ~x55 & ~x62 & ~x65 & ~x72 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2153 =  x7 &  x17 &  x18 &  x19 &  x26 &  x28 &  x29 &  x30 &  x31 &  x36 &  x38 &  x40 &  x46 &  x48 &  x49 &  x50 &  x51 &  x57 &  x58 &  x60 &  x66 &  x69 &  x76 &  x77 &  x78 &  x79 &  x80 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x35 & ~x42 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x64 & ~x72 & ~x73 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c2155 =  x93;
assign c2157 =  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x2 & ~x4 & ~x5 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2159 = ~x69;
assign c2161 =  x16 &  x19 &  x26 &  x27 &  x28 &  x29 &  x36 &  x38 &  x39 &  x47 &  x51 &  x56 &  x57 &  x58 &  x60 &  x68 &  x71 &  x78 &  x79 &  x80 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x2 & ~x8 & ~x33 & ~x35 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x72 & ~x73 & ~x74 & ~x81 & ~x82 & ~x92 & ~x94;
assign c2163 = ~x18;
assign c2165 =  x62;
assign c2167 = ~x18;
assign c2169 =  x1;
assign c2171 =  x1;
assign c2173 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x2 & ~x4 & ~x5 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2175 =  x33;
assign c2177 =  x24;
assign c2179 =  x54;
assign c2181 = ~x30;
assign c2183 =  x62;
assign c2185 =  x1;
assign c2187 =  x93;
assign c2189 =  x2;
assign c2191 =  x0 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x46 &  x47 &  x48 &  x56 &  x58 &  x59 &  x66 &  x67 &  x68 &  x76 &  x77 &  x86 &  x87 &  x89 & ~x1 & ~x4 & ~x23 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c2193 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x1 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2195 =  x2;
assign c2197 = ~x69;
assign c2199 =  x93;
assign c2201 =  x1;
assign c2203 =  x2;
assign c2205 =  x1;
assign c2207 =  x44;
assign c2209 = ~x29;
assign c2211 = ~x30;
assign c2213 =  x2;
assign c2215 =  x16 &  x17 &  x18 &  x20 &  x26 &  x27 &  x29 &  x36 &  x38 &  x39 &  x46 &  x49 &  x58 &  x59 &  x68 &  x76 &  x77 &  x78 &  x80 &  x86 &  x89 &  x90 & ~x0 & ~x15 & ~x25 & ~x33 & ~x34 & ~x35 & ~x44 & ~x52 & ~x54 & ~x55 & ~x62 & ~x64 & ~x65 & ~x72 & ~x73 & ~x75 & ~x81 & ~x83 & ~x85 & ~x92 & ~x94 & ~x95;
assign c2217 =  x0 &  x3 &  x16 &  x26 &  x27 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x57 &  x66 &  x67 &  x69 &  x77 &  x79 &  x86 &  x87 &  x88 & ~x2 & ~x24 & ~x54 & ~x55 & ~x62 & ~x64 & ~x65 & ~x72 & ~x75 & ~x92 & ~x93 & ~x94;
assign c2219 =  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x30 &  x36 &  x37 &  x38 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x80 &  x86 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x2 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2221 =  x1;
assign c2223 = ~x89;
assign c2225 =  x0 &  x3 &  x26 &  x27 &  x28 &  x36 &  x37 &  x38 &  x46 &  x47 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x70 &  x76 &  x77 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x44 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x84 & ~x85 & ~x94;
assign c2227 = ~x30;
assign c2231 =  x2;
assign c2233 =  x16 &  x19 &  x20 &  x27 &  x28 &  x31 &  x36 &  x37 &  x39 &  x40 &  x46 &  x48 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2235 =  x33;
assign c2237 =  x0 &  x3 &  x16 &  x27 &  x29 &  x36 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x86 &  x87 &  x89 & ~x1 & ~x2 & ~x24 & ~x25 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x63 & ~x64 & ~x65 & ~x75 & ~x83 & ~x84 & ~x85 & ~x95;
assign c2239 =  x44;
assign c2241 =  x27 &  x56 &  x66 &  x78 &  x80 & ~x4 & ~x5 & ~x24 & ~x25 & ~x33 & ~x34 & ~x45 & ~x52 & ~x64 & ~x82 & ~x84 & ~x94;
assign c2243 =  x0 &  x3 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x46 &  x47 &  x48 &  x56 &  x58 &  x59 &  x60 &  x66 &  x67 &  x69 &  x76 &  x77 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x2 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x54 & ~x55 & ~x63 & ~x64 & ~x73 & ~x75 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c2245 = ~x30;
assign c2247 =  x0 &  x3 &  x16 &  x17 &  x19 &  x26 &  x29 &  x36 &  x38 &  x39 &  x46 &  x47 &  x48 &  x51 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x69 &  x76 &  x77 &  x78 &  x88 & ~x1 & ~x35 & ~x43 & ~x44 & ~x54 & ~x55 & ~x63 & ~x65 & ~x75 & ~x83 & ~x85 & ~x93 & ~x95;
assign c2249 =  x1;
assign c2251 =  x2;
assign c2253 =  x24;
assign c2255 =  x54;
assign c2261 =  x0 &  x17 &  x18 &  x19 &  x28 &  x30 &  x38 &  x47 &  x48 &  x59 &  x60 &  x67 &  x68 &  x69 &  x70 &  x76 &  x88 & ~x1 & ~x4 & ~x24 & ~x32 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x55 & ~x64 & ~x65 & ~x73 & ~x85 & ~x95;
assign c2265 =  x0 &  x3 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 & ~x2 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x94 & ~x95;
assign c2267 =  x93;
assign c2269 =  x62;
assign c2271 =  x62;
assign c2273 = ~x59;
assign c2275 =  x1;
assign c2277 =  x43;
assign c2279 =  x25;
assign c2281 = ~x17;
assign c2283 =  x26 &  x29 &  x49 &  x50 &  x58 &  x68 &  x80 &  x86 &  x87 &  x91 & ~x21 & ~x22 & ~x45 & ~x72 & ~x81 & ~x83;
assign c2285 =  x43;
assign c2287 = ~x18;
assign c2289 =  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2291 =  x2;
assign c2293 =  x1;
assign c2295 =  x16 &  x19 &  x26 &  x27 &  x31 &  x36 &  x37 &  x38 &  x46 &  x47 &  x49 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x90 & ~x0 & ~x1 & ~x2 & ~x3 & ~x22 & ~x23 & ~x25 & ~x33 & ~x34 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x64 & ~x72 & ~x73 & ~x74 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x95;
assign c2297 =  x33;
assign c2299 = ~x18;
assign c2301 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x2 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2303 =  x2;
assign c2305 =  x1;
assign c2307 = ~x89;
assign c2309 =  x1;
assign c2311 =  x1;
assign c2313 =  x33;
assign c2315 =  x1;
assign c2317 =  x93;
assign c2319 =  x7 &  x88 &  x91 & ~x5 & ~x8 & ~x22 & ~x32 & ~x92;
assign c2321 =  x54;
assign c2323 =  x1;
assign c2325 =  x16 &  x18 &  x19 &  x26 &  x28 &  x29 &  x30 &  x36 &  x37 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x58 &  x59 &  x66 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x89 &  x90 & ~x2 & ~x4 & ~x23 & ~x24 & ~x32 & ~x33 & ~x35 & ~x44 & ~x45 & ~x53 & ~x55 & ~x62 & ~x63 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x95;
assign c2327 =  x16 &  x17 &  x18 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x2 & ~x22 & ~x23 & ~x24 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x64 & ~x65 & ~x72 & ~x73 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x95;
assign c2329 =  x0 &  x3 &  x16 &  x17 &  x26 &  x27 &  x36 &  x37 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x58 &  x59 &  x67 &  x69 &  x70 &  x76 &  x77 &  x87 &  x88 & ~x1 & ~x2 & ~x24 & ~x25 & ~x35 & ~x43 & ~x45 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x84 & ~x85 & ~x95;
assign c2331 =  x0 &  x3 &  x17 &  x18 &  x19 &  x27 &  x28 &  x37 &  x38 &  x39 &  x46 &  x48 &  x49 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x70 &  x76 &  x77 &  x79 &  x86 &  x87 &  x88 & ~x1 & ~x24 & ~x25 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x83 & ~x84 & ~x85 & ~x95;
assign c2333 =  x93;
assign c2335 =  x0 &  x3 &  x16 &  x18 &  x19 &  x27 &  x28 &  x36 &  x38 &  x39 &  x46 &  x47 &  x48 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x2 & ~x23 & ~x24 & ~x25 & ~x34 & ~x35 & ~x43 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x74 & ~x75 & ~x84 & ~x85;
assign c2337 =  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x37 &  x38 &  x39 &  x46 &  x56 &  x57 &  x59 &  x60 &  x66 &  x67 &  x68 &  x76 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x2 & ~x4 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x45 & ~x54 & ~x55 & ~x62 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2339 =  x43;
assign c2341 =  x2;
assign c2343 =  x1;
assign c2345 =  x2;
assign c2347 =  x0 &  x18 &  x26 &  x29 &  x30 &  x37 &  x38 &  x47 &  x48 &  x50 &  x56 &  x57 &  x59 &  x66 &  x67 &  x78 &  x86 &  x88 &  x90 & ~x2 & ~x4 & ~x25 & ~x32 & ~x34 & ~x35 & ~x44 & ~x55 & ~x65 & ~x74 & ~x75 & ~x82 & ~x85 & ~x92 & ~x94 & ~x95;
assign c2349 =  x33;
assign c2351 =  x1;
assign c2353 =  x2;
assign c2355 =  x2;
assign c2357 =  x1;
assign c2359 =  x2;
assign c2361 = ~x68;
assign c2363 =  x1;
assign c2365 = ~x30;
assign c2367 =  x94;
assign c2369 =  x1;
assign c2371 =  x1;
assign c2373 =  x0 &  x16 &  x17 &  x19 &  x26 &  x28 &  x29 &  x30 &  x36 &  x37 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x2 & ~x4 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x73 & ~x75 & ~x84 & ~x85 & ~x93 & ~x95;
assign c2375 =  x1;
assign c2377 =  x23;
assign c2379 =  x0 &  x16 &  x18 &  x19 &  x30 &  x37 &  x40 &  x46 &  x50 &  x59 &  x66 &  x77 &  x78 &  x87 & ~x1 & ~x4 & ~x25 & ~x33 & ~x35 & ~x45 & ~x64 & ~x75 & ~x92;
assign c2381 = ~x69;
assign c2385 =  x2;
assign c2387 =  x1;
assign c2389 =  x16 &  x17 &  x26 &  x28 &  x29 &  x30 &  x31 &  x36 &  x38 &  x40 &  x41 &  x48 &  x50 &  x51 &  x56 &  x58 &  x66 &  x67 &  x68 &  x69 &  x77 &  x78 &  x86 &  x90 & ~x0 & ~x2 & ~x7 & ~x22 & ~x23 & ~x24 & ~x43 & ~x44 & ~x52 & ~x53 & ~x62 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x83 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2391 =  x33;
assign c2393 =  x2;
assign c2397 =  x24;
assign c2399 = ~x31;
assign c2401 =  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x36 &  x40 &  x46 &  x47 &  x48 &  x49 &  x51 &  x57 &  x58 &  x59 &  x60 &  x67 &  x68 &  x76 &  x79 &  x86 &  x87 & ~x0 & ~x3 & ~x24 & ~x35 & ~x45 & ~x52 & ~x54 & ~x74 & ~x75 & ~x84 & ~x93 & ~x94;
assign c2403 =  x1;
assign c2405 = ~x60;
assign c2407 =  x1;
assign c2409 =  x0 &  x3 &  x16 &  x17 &  x18 &  x19 &  x27 &  x30 &  x36 &  x38 &  x39 &  x46 &  x47 &  x48 &  x57 &  x59 &  x60 &  x66 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x89 &  x90 & ~x24 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x63 & ~x64 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x95;
assign c2411 = ~x30;
assign c2413 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x1 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x54 & ~x55 & ~x62 & ~x63 & ~x65 & ~x72 & ~x73 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2415 =  x2;
assign c2417 = ~x89;
assign c2419 =  x2;
assign c2421 = ~x90;
assign c2423 = ~x89;
assign c2425 =  x24;
assign c2427 =  x1;
assign c2429 =  x2;
assign c2431 =  x4 &  x6 &  x8 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2433 =  x72;
assign c2435 =  x17 &  x20 &  x28 &  x30 &  x36 &  x57 &  x60 &  x66 &  x69 &  x71 &  x78 &  x80 &  x86 &  x87 & ~x0 & ~x3 & ~x32 & ~x33 & ~x43 & ~x44 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x73 & ~x74 & ~x84 & ~x92 & ~x93 & ~x95;
assign c2437 =  x93;
assign c2439 =  x2;
assign c2441 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x2 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2443 =  x24;
assign c2445 = ~x17;
assign c2447 = ~x59;
assign c2449 =  x4 &  x5 &  x16 &  x17 &  x18 &  x19 &  x26 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x60 &  x66 &  x69 &  x77 &  x78 &  x80 &  x86 &  x88 &  x89 &  x91 & ~x0 & ~x1 & ~x2 & ~x22 & ~x23 & ~x24 & ~x32 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x92 & ~x93 & ~x94;
assign c2451 =  x21 &  x43;
assign c2455 =  x93;
assign c2457 =  x62;
assign c2459 =  x2;
assign c2461 =  x1;
assign c2463 =  x1;
assign c2465 =  x2;
assign c2467 =  x2;
assign c2469 =  x34;
assign c2471 =  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c2473 =  x16 &  x17 &  x26 &  x29 &  x30 &  x36 &  x37 &  x38 &  x40 &  x46 &  x48 &  x49 &  x50 &  x51 &  x56 &  x58 &  x60 &  x66 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x14 & ~x22 & ~x23 & ~x25 & ~x33 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x84 & ~x92 & ~x93;
assign c2475 =  x1;
assign c2477 = ~x89;
assign c2479 =  x0 &  x17 &  x18 &  x26 &  x37 &  x46 &  x56 &  x67 &  x68 &  x87 & ~x1 & ~x3 & ~x4 & ~x24 & ~x25 & ~x34 & ~x55 & ~x93;
assign c2481 =  x73;
assign c2483 =  x0 &  x3 &  x16 &  x30 &  x36 &  x48 &  x56 &  x57 &  x59 &  x60 &  x68 &  x69 &  x70 &  x77 & ~x2 & ~x25 & ~x33 & ~x43 & ~x44 & ~x45 & ~x65 & ~x74 & ~x75 & ~x82 & ~x83 & ~x95;
assign c2485 =  x62;
assign c2487 =  x2;
assign c2489 = ~x18;
assign c2493 =  x73;
assign c2495 =  x93;
assign c2497 =  x2;
assign c2499 = ~x30;
assign c30 = ~x76;
assign c32 =  x0 &  x16 &  x17 &  x19 &  x20 &  x29 &  x38 &  x39 &  x40 &  x60 &  x68 &  x92 & ~x23 & ~x32 & ~x35 & ~x54 & ~x65 & ~x72 & ~x75;
assign c34 =  x0 &  x2 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 & ~x1 & ~x3 & ~x4 & ~x5 & ~x23 & ~x24 & ~x25 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c36 =  x75;
assign c38 = ~x37;
assign c310 =  x0 &  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x3 & ~x4 & ~x5 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x83 & ~x84 & ~x85 & ~x94 & ~x95;
assign c312 = ~x16;
assign c314 = ~x76;
assign c316 =  x2 &  x17 &  x18 &  x19 &  x26 &  x27 &  x29 &  x30 &  x39 &  x40 &  x46 &  x47 &  x48 &  x57 &  x59 &  x60 &  x67 &  x69 & ~x1 & ~x4 & ~x6 & ~x7 & ~x25 & ~x35 & ~x42 & ~x44 & ~x45 & ~x54 & ~x65 & ~x72 & ~x74 & ~x82 & ~x84 & ~x85 & ~x93;
assign c318 =  x0 &  x8 &  x16 &  x17 &  x18 &  x27 &  x28 &  x36 &  x37 &  x40 &  x41 &  x46 &  x47 &  x48 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x67 &  x68 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 & ~x23 & ~x24 & ~x25 & ~x35 & ~x42 & ~x44 & ~x52 & ~x53 & ~x54 & ~x55 & ~x61 & ~x62 & ~x63 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85;
assign c320 =  x5 & ~x30;
assign c322 = ~x27;
assign c324 =  x4 &  x21 &  x27 &  x28 &  x37 &  x41 &  x46 &  x50 &  x56 &  x67 &  x70 &  x79 &  x88 & ~x23 & ~x34 & ~x42 & ~x43 & ~x52 & ~x53 & ~x82 & ~x83 & ~x85 & ~x94;
assign c326 =  x35;
assign c328 = ~x46;
assign c330 =  x4 &  x5 &  x16 &  x17 &  x18 &  x26 &  x27 &  x36 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x68 &  x69 &  x70 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x23 & ~x24 & ~x25 & ~x31 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x95;
assign c332 = ~x76;
assign c334 =  x0 &  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x3 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c336 = ~x26;
assign c338 =  x2 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 & ~x1 & ~x4 & ~x5 & ~x6 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c340 =  x75;
assign c342 = ~x90;
assign c344 =  x2 &  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x4 & ~x5 & ~x6 & ~x23 & ~x24 & ~x25 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c346 =  x55;
assign c348 =  x2 &  x18 &  x20 &  x26 &  x27 &  x36 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x87 & ~x1 & ~x4 & ~x5 & ~x23 & ~x34 & ~x35 & ~x42 & ~x44 & ~x53 & ~x63 & ~x64 & ~x74 & ~x82 & ~x84 & ~x85 & ~x91;
assign c350 =  x0 &  x16 &  x17 &  x20 &  x26 &  x27 &  x28 &  x36 &  x38 &  x39 &  x40 &  x46 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x60 &  x67 &  x69 &  x70 &  x76 &  x77 &  x78 &  x87 &  x90 &  x91 &  x92 & ~x1 & ~x24 & ~x25 & ~x32 & ~x35 & ~x43 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x72 & ~x73 & ~x74 & ~x75 & ~x84 & ~x85 & ~x94 & ~x95;
assign c352 =  x2 &  x5 &  x16 &  x17 &  x18 &  x26 &  x27 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x31 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c354 =  x2 &  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x4 & ~x5 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c356 =  x4 &  x16 &  x18 &  x19 &  x20 &  x28 &  x31 &  x32 &  x36 &  x39 &  x40 &  x41 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x86 &  x87 &  x89 & ~x24 & ~x34 & ~x35 & ~x42 & ~x45 & ~x52 & ~x53 & ~x54 & ~x65 & ~x74 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x94 & ~x95;
assign c358 = ~x57;
assign c360 = ~x46;
assign c362 = ~x56;
assign c364 =  x4 &  x5 &  x16 &  x17 &  x18 &  x19 &  x20 &  x21 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x32 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x25 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x95;
assign c366 =  x2 &  x3 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x36 &  x37 &  x38 &  x40 &  x46 &  x48 &  x49 &  x56 &  x57 &  x58 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x79 &  x80 &  x86 &  x88 &  x89 &  x90 & ~x1 & ~x4 & ~x5 & ~x6 & ~x23 & ~x24 & ~x25 & ~x34 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x65 & ~x72 & ~x73 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c368 = ~x47;
assign c370 =  x2 &  x16 &  x17 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x38 &  x40 &  x46 &  x47 &  x48 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x4 & ~x5 & ~x9 & ~x24 & ~x25 & ~x34 & ~x35 & ~x44 & ~x45 & ~x53 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x75 & ~x84 & ~x85 & ~x94 & ~x95;
assign c372 =  x16 &  x17 &  x18 &  x19 &  x20 &  x21 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x32 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x23 & ~x24 & ~x25 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c374 =  x0 &  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x40 &  x41 &  x46 &  x47 &  x48 &  x50 &  x56 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x71 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x89 &  x90 & ~x3 & ~x4 & ~x22 & ~x23 & ~x25 & ~x32 & ~x33 & ~x35 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x94 & ~x95;
assign c376 = ~x56;
assign c378 =  x33;
assign c380 = ~x67;
assign c384 = ~x67;
assign c386 = ~x37;
assign c388 =  x4 &  x5 &  x9 &  x10 &  x16 &  x17 &  x18 &  x26 &  x36 &  x38 &  x39 &  x40 &  x48 &  x49 &  x50 &  x51 &  x56 &  x58 &  x59 &  x60 &  x66 &  x67 &  x69 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x90 & ~x1 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x64 & ~x73 & ~x83 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c390 =  x2 &  x4 &  x5 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x3 & ~x9 & ~x23 & ~x24 & ~x25 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x75 & ~x83 & ~x84 & ~x85 & ~x94 & ~x95;
assign c392 =  x2 &  x33 &  x86 &  x87 & ~x62 & ~x82 & ~x95;
assign c394 = ~x68;
assign c396 =  x19 &  x20 &  x29 &  x41 &  x49 &  x76 &  x78 &  x92 & ~x24 & ~x63 & ~x83 & ~x95;
assign c398 = ~x76;
assign c3100 =  x2 &  x4 &  x5 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c3102 =  x0 &  x2 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x3 & ~x4 & ~x6 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c3104 =  x85;
assign c3106 =  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x4 & ~x6 & ~x12 & ~x23 & ~x24 & ~x25 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c3108 = ~x89;
assign c3110 =  x55 &  x95;
assign c3112 =  x5 & ~x30;
assign c3114 = ~x16;
assign c3116 =  x2 &  x5 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x3 & ~x6 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c3118 = ~x28;
assign c3120 = ~x76;
assign c3122 = ~x36;
assign c3124 =  x4 &  x16 &  x17 &  x18 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x32 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x67 &  x68 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x87 & ~x23 & ~x25 & ~x35 & ~x42 & ~x45 & ~x53 & ~x55 & ~x63 & ~x73 & ~x74 & ~x82 & ~x92 & ~x93 & ~x94;
assign c3126 =  x20 &  x30 &  x92 & ~x71;
assign c3128 =  x20 &  x92 & ~x71;
assign c3130 =  x5 &  x32 &  x66 &  x67 & ~x1 & ~x34 & ~x42 & ~x45;
assign c3132 =  x85;
assign c3134 = ~x86;
assign c3136 =  x33 & ~x4;
assign c3138 =  x18 &  x27 &  x79 & ~x20 & ~x21 & ~x22 & ~x44 & ~x52 & ~x53 & ~x83 & ~x92 & ~x94;
assign c3140 = ~x56;
assign c3142 = ~x76;
assign c3144 = ~x56;
assign c3146 =  x2 &  x16 &  x17 &  x18 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x48 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x87 &  x89 & ~x1 & ~x3 & ~x23 & ~x24 & ~x25 & ~x33 & ~x35 & ~x43 & ~x52 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x71 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x95;
assign c3148 =  x4 &  x5 &  x18 &  x79 & ~x3 & ~x31 & ~x55 & ~x83;
assign c3150 =  x4 &  x5 &  x16 &  x18 &  x26 &  x27 &  x37 &  x38 &  x39 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x89 &  x90 & ~x1 & ~x23 & ~x24 & ~x25 & ~x31 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x94 & ~x95;
assign c3152 =  x0 &  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x3 & ~x4 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x94 & ~x95;
assign c3154 = ~x76;
assign c3156 =  x4 &  x5 &  x6 &  x7 &  x9 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x59 &  x60 &  x66 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x23 & ~x24 & ~x25 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c3158 =  x64;
assign c3160 = ~x67;
assign c3162 =  x0 &  x2 &  x16 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x36 &  x37 &  x38 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 & ~x1 & ~x3 & ~x4 & ~x5 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x95;
assign c3164 = ~x36;
assign c3166 =  x0 &  x20 &  x92 & ~x23 & ~x73 & ~x84 & ~x94 & ~x95;
assign c3168 = ~x66;
assign c3170 = ~x28;
assign c3172 =  x0 &  x16 &  x18 &  x19 &  x20 &  x29 &  x36 &  x38 &  x39 &  x40 &  x47 &  x49 &  x66 &  x68 &  x69 &  x70 &  x88 &  x92 & ~x1 & ~x23 & ~x24 & ~x32 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x72 & ~x75 & ~x84 & ~x95;
assign c3174 =  x84 & ~x16;
assign c3176 =  x0 &  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x37 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x3 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x73 & ~x74 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c3178 = ~x39;
assign c3180 =  x5 &  x33 & ~x43;
assign c3182 =  x2 &  x16 &  x17 &  x18 &  x26 &  x27 &  x28 &  x29 &  x36 &  x38 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x60 &  x66 &  x68 &  x76 &  x78 &  x79 &  x80 &  x81 &  x86 &  x89 & ~x1 & ~x9 & ~x21 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x65 & ~x75 & ~x84 & ~x85 & ~x94;
assign c3184 =  x33 & ~x7 & ~x83;
assign c3186 =  x2 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x81 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x3 & ~x21 & ~x22 & ~x23 & ~x24 & ~x25 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c3188 =  x2 &  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x4 & ~x5 & ~x6 & ~x23 & ~x24 & ~x25 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c3190 = ~x86;
assign c3192 =  x84;
assign c3194 = ~x16;
assign c3196 = ~x19;
assign c3198 =  x2 &  x16 &  x17 &  x26 &  x27 &  x28 &  x36 &  x37 &  x38 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x67 &  x68 &  x70 &  x76 &  x86 &  x88 & ~x1 & ~x6 & ~x22 & ~x23 & ~x25 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x62 & ~x63 & ~x64 & ~x73 & ~x75 & ~x84 & ~x85 & ~x91 & ~x92 & ~x93 & ~x94 & ~x95;
assign c3200 =  x72;
assign c3202 = ~x37;
assign c3204 =  x2 &  x17 &  x18 &  x27 &  x28 &  x29 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x57 &  x58 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x81 &  x86 &  x87 &  x90 & ~x1 & ~x7 & ~x22 & ~x24 & ~x32 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x94 & ~x95;
assign c3206 =  x4 &  x5 &  x16 &  x17 &  x18 &  x19 &  x21 &  x26 &  x27 &  x28 &  x29 &  x30 &  x32 &  x36 &  x37 &  x39 &  x41 &  x46 &  x48 &  x56 &  x58 &  x59 &  x66 &  x67 &  x69 &  x70 &  x76 &  x77 &  x87 & ~x1 & ~x25 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x94 & ~x95;
assign c3208 = ~x76;
assign c3210 = ~x90;
assign c3212 =  x0 &  x2 &  x17 &  x18 &  x26 &  x27 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x67 &  x68 &  x70 &  x76 &  x78 &  x79 &  x80 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x4 & ~x6 & ~x23 & ~x24 & ~x25 & ~x34 & ~x35 & ~x42 & ~x44 & ~x45 & ~x52 & ~x53 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x74 & ~x75 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c3214 =  x0 &  x20 &  x26 &  x27 &  x37 &  x39 &  x48 &  x49 &  x56 &  x57 &  x58 &  x60 &  x66 &  x77 &  x87 &  x88 &  x90 &  x92 & ~x1 & ~x23 & ~x32 & ~x33 & ~x45 & ~x54 & ~x62 & ~x72 & ~x75 & ~x95;
assign c3216 = ~x66;
assign c3218 =  x55;
assign c3220 =  x84;
assign c3222 =  x2 &  x21 &  x22 &  x38 &  x48 &  x51 &  x77 & ~x44 & ~x72 & ~x83 & ~x85 & ~x95;
assign c3224 =  x2 &  x3 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 & ~x1 & ~x4 & ~x5 & ~x6 & ~x23 & ~x24 & ~x25 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x61 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c3226 =  x0 &  x2 &  x17 &  x18 &  x19 &  x20 &  x27 &  x28 &  x29 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x49 &  x50 &  x57 &  x58 &  x59 &  x67 &  x68 &  x70 &  x76 &  x77 &  x87 &  x88 &  x89 & ~x1 & ~x4 & ~x5 & ~x23 & ~x24 & ~x25 & ~x33 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x55 & ~x62 & ~x72 & ~x83 & ~x84 & ~x93 & ~x94 & ~x95;
assign c3228 = ~x38;
assign c3230 =  x2 &  x4 &  x5 &  x16 &  x17 &  x18 &  x19 &  x20 &  x27 &  x28 &  x29 &  x36 &  x37 &  x38 &  x48 &  x49 &  x50 &  x56 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x78 &  x79 &  x86 &  x87 &  x88 &  x90 & ~x0 & ~x1 & ~x3 & ~x22 & ~x23 & ~x25 & ~x32 & ~x34 & ~x35 & ~x42 & ~x44 & ~x45 & ~x52 & ~x53 & ~x55 & ~x62 & ~x64 & ~x65 & ~x72 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x93 & ~x95;
assign c3232 =  x0 &  x20 &  x48 &  x67 &  x79 &  x92 & ~x23 & ~x32 & ~x64 & ~x73 & ~x84 & ~x95;
assign c3234 = ~x67;
assign c3236 = ~x66;
assign c3238 =  x4 &  x5 &  x6 &  x16 &  x17 &  x18 &  x19 &  x20 &  x21 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x86 &  x87 &  x89 &  x90 & ~x1 & ~x23 & ~x24 & ~x25 & ~x34 & ~x35 & ~x42 & ~x43 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x92 & ~x93 & ~x94;
assign c3240 =  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x21 &  x27 &  x28 &  x29 &  x38 &  x41 &  x48 &  x49 &  x50 &  x51 &  x57 &  x66 &  x68 &  x69 &  x77 &  x78 &  x89 & ~x1 & ~x3 & ~x23 & ~x25 & ~x35 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x65 & ~x71 & ~x73 & ~x75 & ~x82 & ~x84;
assign c3242 = ~x56;
assign c3244 =  x44;
assign c3246 =  x0 &  x2 &  x16 &  x17 &  x18 &  x26 &  x27 &  x28 &  x29 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x67 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x90 & ~x1 & ~x3 & ~x4 & ~x5 & ~x23 & ~x24 & ~x25 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x94 & ~x95;
assign c3248 =  x2 &  x17 &  x20 &  x21 &  x27 &  x28 &  x37 &  x41 &  x47 &  x48 &  x49 &  x51 &  x57 &  x58 &  x59 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 & ~x1 & ~x3 & ~x23 & ~x24 & ~x25 & ~x35 & ~x43 & ~x44 & ~x54 & ~x55 & ~x62 & ~x65 & ~x73 & ~x74 & ~x82 & ~x84 & ~x85 & ~x91 & ~x92 & ~x95;
assign c3250 = ~x37;
assign c3252 =  x0 &  x2 &  x16 &  x17 &  x18 &  x26 &  x36 &  x37 &  x38 &  x40 &  x46 &  x47 &  x48 &  x49 &  x56 &  x58 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x3 & ~x4 & ~x6 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x94 & ~x95;
assign c3254 = ~x16;
assign c3256 =  x0 &  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x4 & ~x6 & ~x24 & ~x25 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c3258 =  x84;
assign c3260 =  x4 &  x5 &  x6 &  x9 &  x16 &  x17 &  x18 &  x19 &  x20 &  x21 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x23 & ~x24 & ~x25 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c3262 =  x44;
assign c3264 =  x45;
assign c3266 = ~x46;
assign c3268 =  x54;
assign c3270 =  x0 &  x7 &  x8 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x1 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c3272 =  x18 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x51 &  x56 &  x67 &  x76 &  x77 &  x79 &  x87 & ~x31 & ~x32 & ~x35 & ~x44 & ~x45 & ~x52 & ~x54 & ~x61 & ~x73 & ~x85 & ~x94;
assign c3274 = ~x16;
assign c3276 =  x0 &  x2 &  x17 &  x18 &  x26 &  x27 &  x28 &  x29 &  x37 &  x38 &  x40 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x87 &  x88 &  x89 & ~x4 & ~x6 & ~x24 & ~x34 & ~x35 & ~x45 & ~x52 & ~x54 & ~x55 & ~x62 & ~x63 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x85 & ~x95;
assign c3278 =  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x61 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x81 &  x86 &  x87 &  x88 & ~x1 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c3282 = ~x16;
assign c3284 = ~x90;
assign c3286 =  x93;
assign c3288 =  x25;
assign c3290 = ~x38;
assign c3292 =  x2 &  x5 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x3 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c3294 = ~x67;
assign c3296 =  x35;
assign c3298 =  x2 &  x5 &  x17 &  x18 &  x27 &  x36 &  x47 &  x49 &  x50 &  x57 &  x60 &  x66 &  x67 &  x68 &  x69 &  x76 &  x78 &  x79 &  x87 &  x88 & ~x3 & ~x22 & ~x23 & ~x31 & ~x32 & ~x53 & ~x55 & ~x63 & ~x64 & ~x65 & ~x74 & ~x83 & ~x84 & ~x92 & ~x94 & ~x95;
assign c3300 = ~x56;
assign c3302 = ~x36;
assign c3304 =  x2 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x4 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x31 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c3306 =  x0 &  x2 &  x16 &  x17 &  x18 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x3 & ~x4 & ~x6 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x75 & ~x83 & ~x84 & ~x85 & ~x95;
assign c3308 = ~x16;
assign c3310 = ~x66;
assign c3312 =  x2 &  x4 &  x18 &  x28 &  x29 &  x30 &  x36 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x58 &  x59 &  x60 &  x66 &  x70 &  x76 &  x77 &  x79 &  x81 &  x88 & ~x0 & ~x22 & ~x23 & ~x24 & ~x35 & ~x43 & ~x45 & ~x52 & ~x53 & ~x54 & ~x62 & ~x63 & ~x65 & ~x72 & ~x73 & ~x75 & ~x92 & ~x93 & ~x94 & ~x95;
assign c3314 =  x85;
assign c3316 = ~x47;
assign c3320 = ~x37;
assign c3322 = ~x56;
assign c3324 =  x85;
assign c3326 = ~x76;
assign c3328 = ~x76;
assign c3330 =  x0 &  x2 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 & ~x1 & ~x3 & ~x4 & ~x5 & ~x23 & ~x24 & ~x25 & ~x34 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x94 & ~x95;
assign c3332 = ~x17;
assign c3334 =  x32;
assign c3336 = ~x46;
assign c3338 =  x2 &  x4 &  x5 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x3 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c3340 =  x35;
assign c3342 = ~x58;
assign c3344 = ~x37;
assign c3346 =  x2 &  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x4 & ~x5 & ~x6 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c3348 =  x71 &  x88 & ~x20;
assign c3350 =  x2 &  x29 &  x50 &  x81 &  x87 &  x90 & ~x0 & ~x61 & ~x82 & ~x83;
assign c3352 =  x5 & ~x30;
assign c3354 = ~x76;
assign c3356 =  x2 &  x18 &  x19 &  x28 &  x37 &  x39 &  x40 &  x46 &  x47 &  x49 &  x50 &  x56 &  x57 &  x58 &  x60 &  x66 &  x67 &  x70 &  x76 &  x77 &  x78 &  x88 &  x89 & ~x1 & ~x3 & ~x7 & ~x24 & ~x25 & ~x35 & ~x43 & ~x45 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x75 & ~x82 & ~x85 & ~x91 & ~x92 & ~x93 & ~x95;
assign c3358 = ~x66;
assign c3360 = ~x16;
assign c3362 = ~x37 & ~x76;
assign c3364 =  x2 &  x16 &  x17 &  x18 &  x26 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 & ~x1 & ~x4 & ~x5 & ~x6 & ~x8 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x95;
assign c3366 =  x2 &  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x4 & ~x5 & ~x6 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c3368 =  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x81 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x21 & ~x22 & ~x23 & ~x24 & ~x25 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c3370 =  x0 &  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x29 &  x30 &  x36 &  x38 &  x39 &  x40 &  x46 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x60 &  x66 &  x67 &  x68 &  x70 &  x77 &  x78 &  x79 &  x80 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x3 & ~x4 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x44 & ~x45 & ~x52 & ~x53 & ~x55 & ~x62 & ~x63 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x94 & ~x95;
assign c3372 = ~x46;
assign c3374 =  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x4 & ~x5 & ~x9 & ~x23 & ~x24 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x64 & ~x72 & ~x74 & ~x75 & ~x82 & ~x83 & ~x85 & ~x93 & ~x95;
assign c3376 =  x2 &  x5 & ~x30;
assign c3378 = ~x57;
assign c3382 =  x0 &  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x4 & ~x6 & ~x24 & ~x25 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x94 & ~x95;
assign c3384 = ~x66;
assign c3386 =  x19 &  x20 &  x29 &  x38 &  x39 &  x41 &  x47 &  x49 &  x50 &  x59 &  x60 &  x67 &  x70 &  x77 &  x79 &  x86 &  x88 &  x89 &  x90 & ~x23 & ~x24 & ~x25 & ~x31 & ~x34 & ~x42 & ~x43 & ~x44 & ~x45 & ~x62 & ~x65 & ~x75 & ~x83 & ~x84 & ~x85 & ~x94;
assign c3388 = ~x37;
assign c3390 =  x16 &  x17 &  x19 &  x20 &  x27 &  x28 &  x29 &  x36 &  x38 &  x39 &  x40 &  x41 &  x47 &  x48 &  x49 &  x51 &  x56 &  x57 &  x58 &  x60 &  x67 &  x68 &  x70 &  x78 &  x86 &  x88 &  x89 & ~x1 & ~x3 & ~x23 & ~x24 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x55 & ~x63 & ~x64 & ~x71 & ~x72 & ~x73 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x95;
assign c3394 =  x2 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x77 &  x78 &  x86 &  x87 & ~x1 & ~x4 & ~x6 & ~x23 & ~x24 & ~x25 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x91 & ~x92 & ~x93 & ~x94 & ~x95;
assign c3398 = ~x86;
assign c3400 =  x33 & ~x42 & ~x82 & ~x95;
assign c3402 =  x0 &  x7 &  x8 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x1 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x94 & ~x95;
assign c3404 =  x19 &  x82 & ~x21;
assign c3406 = ~x26;
assign c3408 =  x85;
assign c3412 =  x0 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x39 &  x40 &  x47 &  x48 &  x49 &  x57 &  x58 &  x59 &  x67 &  x70 &  x77 &  x78 &  x79 &  x87 &  x88 &  x89 &  x92 & ~x1 & ~x23 & ~x24 & ~x35 & ~x44 & ~x45 & ~x53 & ~x54 & ~x64 & ~x83 & ~x85 & ~x94 & ~x95;
assign c3414 =  x16 &  x17 &  x26 &  x28 &  x36 &  x39 &  x40 &  x41 &  x47 &  x49 &  x51 &  x56 &  x60 &  x66 &  x68 &  x70 &  x76 &  x87 &  x88 & ~x1 & ~x3 & ~x23 & ~x32 & ~x33 & ~x45 & ~x55 & ~x65 & ~x74 & ~x75 & ~x82 & ~x85 & ~x91 & ~x92 & ~x93;
assign c3416 =  x2 &  x3 &  x18 &  x27 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x49 &  x51 &  x56 &  x57 &  x59 &  x60 &  x66 &  x76 &  x78 &  x79 &  x90 & ~x1 & ~x4 & ~x5 & ~x6 & ~x25 & ~x33 & ~x34 & ~x44 & ~x45 & ~x52 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x85 & ~x95;
assign c3418 =  x79 & ~x30;
assign c3420 =  x2 &  x26 &  x27 &  x36 &  x38 &  x48 &  x49 &  x51 &  x58 &  x59 &  x66 &  x67 &  x77 &  x78 &  x79 &  x88 & ~x1 & ~x6 & ~x23 & ~x25 & ~x32 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x62 & ~x63 & ~x74 & ~x75 & ~x85 & ~x91 & ~x92 & ~x95;
assign c3422 = ~x16;
assign c3424 =  x0 &  x2 &  x10 &  x16 &  x17 &  x18 &  x26 &  x27 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x3 & ~x4 & ~x23 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c3426 = ~x30 & ~x91;
assign c3428 =  x2 &  x17 &  x19 &  x27 &  x32 &  x36 &  x48 &  x49 &  x50 &  x51 &  x56 &  x60 &  x67 &  x68 &  x69 &  x70 &  x77 &  x78 &  x88 &  x89 & ~x0 & ~x1 & ~x3 & ~x25 & ~x43 & ~x44 & ~x53 & ~x54 & ~x62 & ~x64 & ~x74 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c3430 =  x8 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x32 &  x39 &  x48 &  x66 &  x69 &  x70 &  x76 &  x77 &  x80 &  x87 &  x88 &  x89 &  x90 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x75 & ~x92 & ~x93 & ~x94;
assign c3432 =  x18 &  x71 & ~x20;
assign c3434 = ~x26;
assign c3436 =  x4 &  x27 &  x32 &  x39 &  x40 &  x41 &  x46 &  x50 &  x56 &  x59 &  x60 &  x68 &  x78 &  x79 & ~x23 & ~x25 & ~x34 & ~x42 & ~x64;
assign c3438 = ~x27;
assign c3440 = ~x67;
assign c3442 =  x2 &  x4 &  x5 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c3444 =  x32 &  x33 & ~x43 & ~x82 & ~x94 & ~x95;
assign c3446 = ~x89;
assign c3448 =  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x3 & ~x23 & ~x24 & ~x25 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x71 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c3450 =  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x21 &  x26 &  x28 &  x29 &  x30 &  x32 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x69 &  x70 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x23 & ~x24 & ~x25 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x92 & ~x93 & ~x94 & ~x95;
assign c3452 = ~x61 & ~x80;
assign c3454 =  x45;
assign c3458 = ~x38;
assign c3460 =  x33 & ~x45 & ~x82 & ~x94;
assign c3462 =  x93;
assign c3464 = ~x76;
assign c3466 =  x2 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x36 &  x40 &  x48 &  x49 &  x57 &  x58 &  x60 &  x66 &  x69 &  x76 &  x78 &  x79 &  x87 & ~x1 & ~x6 & ~x7 & ~x24 & ~x63 & ~x72 & ~x74 & ~x94 & ~x95;
assign c3468 =  x2 &  x16 &  x17 &  x26 &  x27 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 & ~x6 & ~x24 & ~x25 & ~x31 & ~x35 & ~x44 & ~x45 & ~x53 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94;
assign c3470 = ~x56;
assign c3472 =  x93;
assign c3474 =  x64 & ~x57;
assign c3476 =  x2 &  x4 &  x5 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x0 & ~x1 & ~x3 & ~x24 & ~x25 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x85 & ~x92 & ~x93 & ~x95;
assign c3478 =  x85;
assign c3480 =  x0 &  x2 &  x16 &  x17 &  x18 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x3 & ~x4 & ~x6 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x95;
assign c3482 =  x0 &  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x3 & ~x4 & ~x23 & ~x24 & ~x25 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c3484 =  x0 &  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x3 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c3486 =  x2 &  x22 &  x70 &  x90 & ~x82;
assign c3488 =  x0 &  x2 &  x17 &  x19 &  x26 &  x36 &  x37 &  x38 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 & ~x4 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x34 & ~x35 & ~x43 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x72 & ~x73 & ~x74 & ~x75 & ~x84 & ~x85 & ~x92 & ~x94 & ~x95;
assign c3490 =  x84;
assign c3492 = ~x56;
assign c3494 =  x32 &  x33 & ~x43 & ~x82;
assign c3496 =  x4 &  x5 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x31 &  x32 &  x36 &  x37 &  x41 &  x46 &  x47 &  x50 &  x56 &  x57 &  x58 &  x60 &  x66 &  x69 &  x70 &  x76 &  x77 &  x87 & ~x1 & ~x25 & ~x43 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x65 & ~x72 & ~x74 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94;
assign c3498 =  x2 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 & ~x1 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x31 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c31 =  x3 &  x42;
assign c33 = ~x36;
assign c35 =  x13 &  x18 &  x19 &  x20 &  x26 &  x27 &  x30 &  x36 &  x37 &  x38 &  x56 &  x57 &  x58 &  x60 &  x67 &  x69 &  x80 &  x88 & ~x7 & ~x22 & ~x25 & ~x33 & ~x34 & ~x42 & ~x43 & ~x44 & ~x53 & ~x55 & ~x65 & ~x73 & ~x81;
assign c37 =  x52;
assign c39 =  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x71 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x0 & ~x3 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x52 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c311 = ~x39;
assign c313 =  x6 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x36 &  x37 &  x38 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x71 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 & ~x1 & ~x7 & ~x22 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c315 =  x4 &  x16 &  x17 &  x18 &  x36 &  x37 &  x39 &  x46 &  x47 &  x49 &  x50 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x69 &  x76 &  x77 &  x78 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x5 & ~x23 & ~x24 & ~x25 & ~x44 & ~x45 & ~x52 & ~x54 & ~x55 & ~x64 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x95;
assign c317 =  x91;
assign c319 =  x3 &  x4;
assign c323 =  x5 &  x6 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c325 = ~x70;
assign c327 =  x2 &  x3 &  x6 &  x16 &  x17 &  x19 &  x28 &  x30 &  x36 &  x37 &  x38 &  x46 &  x67 &  x77 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x22 & ~x23 & ~x24 & ~x25 & ~x34 & ~x35 & ~x44 & ~x85 & ~x95;
assign c329 =  x25;
assign c331 =  x0 &  x2 &  x4 &  x16 &  x17 &  x19 &  x26 &  x29 &  x36 &  x49 &  x56 &  x58 &  x66 &  x76 &  x79 &  x80 &  x86 & ~x22 & ~x25 & ~x33 & ~x35 & ~x65 & ~x82 & ~x85 & ~x92;
assign c333 =  x1;
assign c335 =  x6 &  x46 &  x47 &  x51 & ~x41 & ~x52 & ~x92;
assign c339 =  x16 &  x17 &  x18 &  x20 &  x26 &  x28 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x61 &  x66 &  x67 &  x69 &  x70 &  x71 &  x76 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x1 & ~x22 & ~x23 & ~x24 & ~x33 & ~x34 & ~x43 & ~x44 & ~x53 & ~x55 & ~x62 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x85 & ~x92 & ~x94 & ~x95;
assign c341 = ~x2;
assign c343 =  x4 &  x18 &  x19 &  x20 &  x27 &  x30 &  x36 &  x38 &  x39 &  x48 &  x50 &  x51 &  x56 &  x57 &  x59 &  x67 &  x68 &  x70 &  x76 &  x87 &  x90 & ~x5 & ~x23 & ~x24 & ~x25 & ~x45 & ~x52 & ~x62 & ~x74 & ~x84 & ~x93 & ~x94;
assign c345 =  x42;
assign c347 =  x1;
assign c349 =  x1;
assign c351 = ~x60;
assign c353 =  x0 & ~x51;
assign c355 =  x4 &  x16 &  x17 &  x26 &  x38 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x86 & ~x1 & ~x5 & ~x23 & ~x24 & ~x25 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x62 & ~x64 & ~x65 & ~x75 & ~x81 & ~x83 & ~x84 & ~x85;
assign c357 = ~x60;
assign c359 =  x3 &  x5 & ~x7;
assign c361 = ~x7;
assign c365 =  x4 &  x16 &  x26 &  x36 &  x37 &  x38 &  x46 &  x47 &  x49 &  x56 &  x57 &  x58 &  x60 &  x66 &  x67 &  x68 &  x69 &  x76 &  x86 & ~x5 & ~x21 & ~x23 & ~x24 & ~x44 & ~x52 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x84 & ~x85 & ~x93 & ~x94;
assign c367 =  x28 &  x29 &  x31 & ~x21 & ~x61 & ~x81 & ~x95;
assign c369 =  x6 & ~x7;
assign c371 =  x52;
assign c373 =  x3 &  x8 &  x61 & ~x92;
assign c375 =  x63;
assign c377 = ~x4;
assign c379 = ~x70;
assign c381 = ~x88;
assign c383 =  x16 &  x20 &  x37 &  x38 &  x39 &  x58 &  x70 &  x76 &  x78 &  x86 &  x88 & ~x2 & ~x32 & ~x43 & ~x52 & ~x92;
assign c385 =  x2 &  x17 &  x19 &  x26 &  x27 &  x29 &  x37 &  x38 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x58 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x78 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x0 & ~x1 & ~x4 & ~x22 & ~x23 & ~x25 & ~x33 & ~x34 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x93 & ~x94;
assign c387 =  x1;
assign c389 =  x62;
assign c391 =  x0 &  x3 & ~x51;
assign c393 =  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x21 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x1 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c395 = ~x70;
assign c397 =  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x4 & ~x22 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c399 = ~x2 & ~x6;
assign c3101 = ~x60;
assign c3103 =  x52;
assign c3105 = ~x60;
assign c3107 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x61 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c3109 =  x6 &  x16 &  x17 &  x20 &  x28 &  x36 &  x37 &  x40 &  x46 &  x48 &  x49 &  x50 &  x57 &  x58 &  x59 &  x67 &  x68 &  x70 &  x76 &  x77 &  x78 &  x80 &  x86 &  x88 &  x89 &  x90 & ~x1 & ~x9 & ~x22 & ~x23 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x52 & ~x62 & ~x64 & ~x65 & ~x73 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x94 & ~x95;
assign c3111 =  x64;
assign c3113 =  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x0 & ~x1 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c3115 =  x73;
assign c3117 = ~x60;
assign c3119 =  x94;
assign c3121 =  x1;
assign c3123 =  x5 &  x18 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x39 &  x46 &  x47 &  x49 &  x57 &  x58 &  x59 &  x66 &  x68 &  x69 &  x76 &  x77 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 & ~x0 & ~x1 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x35 & ~x43 & ~x45 & ~x52 & ~x53 & ~x54 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x84 & ~x85 & ~x93 & ~x95;
assign c3125 =  x52;
assign c3127 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c3129 =  x1;
assign c3131 = ~x2 & ~x7;
assign c3133 =  x4 &  x16 &  x26 &  x27 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x57 &  x58 &  x59 &  x60 &  x66 &  x68 &  x69 &  x76 &  x77 &  x86 & ~x1 & ~x5 & ~x22 & ~x23 & ~x25 & ~x34 & ~x35 & ~x42 & ~x44 & ~x45 & ~x53 & ~x54 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84;
assign c3135 =  x4 &  x17 &  x18 &  x20 &  x26 &  x28 &  x36 &  x38 &  x39 &  x40 &  x46 &  x48 &  x49 &  x50 &  x56 &  x58 &  x60 &  x66 &  x68 &  x69 &  x76 &  x77 &  x79 &  x86 &  x87 &  x89 & ~x5 & ~x23 & ~x24 & ~x35 & ~x52 & ~x53 & ~x54 & ~x65 & ~x75 & ~x94 & ~x95;
assign c3137 =  x4 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x59 &  x66 &  x68 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x89 &  x90 & ~x1 & ~x5 & ~x24 & ~x25 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x63 & ~x65 & ~x72 & ~x73 & ~x75 & ~x85 & ~x94;
assign c3141 =  x52;
assign c3143 =  x1;
assign c3145 =  x4 &  x16 &  x36 &  x37 &  x46 &  x48 &  x56 &  x58 &  x66 &  x67 &  x68 &  x71 &  x77 &  x86 &  x87 &  x88 & ~x5 & ~x23 & ~x24 & ~x33 & ~x35 & ~x43 & ~x62 & ~x63 & ~x73 & ~x85 & ~x94;
assign c3147 =  x0 &  x2 &  x4 &  x16 &  x17 &  x18 &  x20 &  x28 &  x30 &  x38 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x60 &  x66 &  x67 &  x69 &  x77 &  x79 &  x86 &  x87 &  x89 & ~x1 & ~x22 & ~x23 & ~x24 & ~x33 & ~x34 & ~x44 & ~x52 & ~x53 & ~x55 & ~x64 & ~x65 & ~x75 & ~x83 & ~x85 & ~x92 & ~x94 & ~x95;
assign c3149 =  x16 &  x36 &  x48 &  x56 & ~x2 & ~x32 & ~x44 & ~x92;
assign c3151 = ~x0 & ~x2;
assign c3153 =  x4 &  x56 &  x57 & ~x5 & ~x10 & ~x55;
assign c3155 =  x16 &  x27 &  x28 &  x29 &  x30 &  x37 &  x38 &  x48 &  x49 &  x50 &  x56 &  x67 &  x76 & ~x21 & ~x22 & ~x41 & ~x43 & ~x45 & ~x52 & ~x53 & ~x81 & ~x84 & ~x92 & ~x93;
assign c3157 =  x1;
assign c3159 =  x16 &  x27 &  x56 &  x86 &  x87 & ~x2 & ~x24 & ~x25 & ~x32 & ~x44 & ~x75;
assign c3161 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x0 & ~x1 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c3163 = ~x6;
assign c3165 =  x1;
assign c3167 = ~x50;
assign c3169 = ~x41;
assign c3171 = ~x2;
assign c3173 =  x2 &  x16 &  x17 &  x19 &  x20 &  x26 &  x28 &  x29 &  x30 &  x31 &  x36 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x70 &  x71 &  x76 &  x79 &  x80 &  x86 &  x87 &  x89 &  x90 &  x91 & ~x22 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x65 & ~x72 & ~x73 & ~x74 & ~x81 & ~x82 & ~x84 & ~x95;
assign c3175 =  x1;
assign c3177 = ~x2 & ~x3;
assign c3179 =  x0 &  x3 & ~x8;
assign c3181 =  x3 &  x18 &  x20 &  x28 &  x36 &  x57 & ~x1 & ~x24 & ~x52 & ~x55 & ~x65 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x91 & ~x93;
assign c3183 = ~x70;
assign c3185 =  x3 &  x72;
assign c3187 = ~x2 & ~x6;
assign c3189 =  x2 &  x5 &  x16 &  x18 &  x20 &  x21 &  x26 &  x27 &  x28 &  x29 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c3191 =  x19 &  x28 &  x37 &  x39 &  x57 &  x58 &  x66 &  x67 &  x69 &  x70 &  x76 &  x91 & ~x7 & ~x32 & ~x33 & ~x42 & ~x43 & ~x52 & ~x63 & ~x74 & ~x81 & ~x82 & ~x83 & ~x92 & ~x93;
assign c3193 =  x63;
assign c3195 =  x52;
assign c3197 = ~x60;
assign c3199 = ~x78;
assign c3201 = ~x50;
assign c3203 =  x5 &  x6 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x1 & ~x4 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x95;
assign c3205 = ~x58;
assign c3209 = ~x88;
assign c3211 =  x2 &  x3 &  x5 &  x56;
assign c3213 =  x52;
assign c3215 =  x1;
assign c3217 =  x1;
assign c3219 =  x36 &  x50 &  x59 &  x67 &  x77 &  x87 & ~x2 & ~x32 & ~x33 & ~x44 & ~x54 & ~x62 & ~x92;
assign c3221 =  x1;
assign c3223 = ~x2;
assign c3225 =  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x30 &  x36 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 & ~x0 & ~x1 & ~x3 & ~x5 & ~x24 & ~x25 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c3227 = ~x70;
assign c3229 =  x61 & ~x41 & ~x92;
assign c3231 =  x19 &  x21 &  x27 &  x30 &  x31 &  x37 &  x39 &  x40 &  x51 &  x57 &  x58 &  x59 &  x68 &  x69 &  x70 &  x71 &  x76 &  x78 &  x80 &  x86 &  x88 & ~x0 & ~x1 & ~x22 & ~x23 & ~x32 & ~x44 & ~x53 & ~x54 & ~x63 & ~x65 & ~x73 & ~x82 & ~x83 & ~x84;
assign c3233 = ~x60;
assign c3235 =  x1;
assign c3237 =  x5 &  x6 &  x16 &  x17 &  x18 &  x20 &  x26 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x60 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x87 &  x89 & ~x1 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x54 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x95;
assign c3239 =  x1;
assign c3241 = ~x2 & ~x6;
assign c3243 = ~x51;
assign c3245 =  x19 &  x46 &  x47 &  x48 &  x51 &  x58 &  x60 &  x66 &  x67 &  x68 &  x70 &  x77 &  x78 & ~x0 & ~x3 & ~x5 & ~x22 & ~x32 & ~x33 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x54 & ~x55 & ~x75 & ~x82 & ~x85 & ~x92 & ~x95;
assign c3247 = ~x69;
assign c3249 =  x4 &  x16 &  x17 &  x18 &  x26 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x5 & ~x23 & ~x24 & ~x25 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c3251 =  x52;
assign c3253 = ~x50;
assign c3255 = ~x2 & ~x6;
assign c3257 =  x16 &  x19 &  x21 &  x26 &  x27 &  x28 &  x30 &  x31 &  x37 &  x39 &  x46 &  x48 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x68 &  x69 &  x70 &  x71 &  x76 &  x78 &  x80 &  x88 &  x89 &  x90 &  x91 & ~x1 & ~x3 & ~x23 & ~x24 & ~x32 & ~x42 & ~x44 & ~x52 & ~x53 & ~x54 & ~x62 & ~x63 & ~x64 & ~x72 & ~x73 & ~x74 & ~x82 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c3259 = ~x50;
assign c3261 =  x4 &  x17 &  x26 &  x37 &  x39 &  x47 &  x48 &  x57 &  x67 &  x69 &  x86 &  x88 & ~x1 & ~x5 & ~x23 & ~x33 & ~x35 & ~x42 & ~x43 & ~x45 & ~x52 & ~x54 & ~x62 & ~x63 & ~x64 & ~x73 & ~x75 & ~x84 & ~x92 & ~x93 & ~x94 & ~x95;
assign c3265 =  x75;
assign c3267 =  x2 &  x17 &  x18 &  x19 &  x20 &  x21 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x48 &  x51 &  x56 &  x58 &  x59 &  x60 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x80 &  x86 &  x87 &  x89 &  x90 & ~x0 & ~x1 & ~x22 & ~x23 & ~x24 & ~x25 & ~x35 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x73 & ~x74 & ~x75 & ~x82 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94;
assign c3269 =  x16 &  x17 &  x19 &  x20 &  x26 &  x28 &  x29 &  x31 &  x36 &  x37 &  x38 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x60 &  x66 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x91 & ~x1 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x52 & ~x62 & ~x63 & ~x64 & ~x73 & ~x74 & ~x81 & ~x83 & ~x84 & ~x92 & ~x95;
assign c3273 =  x0 &  x2 &  x4 &  x16 &  x20 &  x26 &  x27 &  x29 &  x30 &  x37 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x60 &  x70 &  x78 &  x79 &  x88 &  x89 &  x90 & ~x23 & ~x24 & ~x25 & ~x34 & ~x35 & ~x43 & ~x45 & ~x55 & ~x63 & ~x64 & ~x74 & ~x75 & ~x82;
assign c3275 =  x83;
assign c3277 =  x1;
assign c3279 =  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x1 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c3281 =  x3 &  x56 & ~x22 & ~x71;
assign c3283 =  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x3 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c3285 =  x2 &  x4 &  x16 &  x26 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x69 &  x76 &  x77 &  x86 &  x88 &  x89 & ~x0 & ~x1 & ~x5 & ~x25 & ~x42 & ~x43 & ~x45 & ~x52 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x72 & ~x74 & ~x83 & ~x85 & ~x94 & ~x95;
assign c3287 =  x2 &  x3 &  x5;
assign c3289 =  x4 &  x16 &  x17 &  x19 &  x26 &  x28 &  x30 &  x36 &  x38 &  x39 &  x46 &  x47 &  x50 &  x56 &  x60 &  x66 &  x67 & ~x6 & ~x24 & ~x25 & ~x32 & ~x35 & ~x43 & ~x45 & ~x53 & ~x54 & ~x63 & ~x64 & ~x65 & ~x85;
assign c3291 = ~x2;
assign c3293 =  x1;
assign c3295 =  x95;
assign c3297 =  x63;
assign c3299 =  x1;
assign c3301 = ~x0 & ~x2;
assign c3303 =  x53;
assign c3305 =  x21 &  x92;
assign c3307 =  x62;
assign c3309 =  x52;
assign c3311 = ~x60;
assign c3313 =  x3 &  x6 &  x37 &  x40 &  x48 &  x57 &  x67 &  x79 & ~x9 & ~x44 & ~x45 & ~x65 & ~x72 & ~x75 & ~x85 & ~x92;
assign c3315 =  x16 &  x17 &  x18 &  x20 &  x26 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x1 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x61 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c3317 =  x4 &  x16 &  x19 &  x20 &  x26 &  x27 &  x28 &  x36 &  x38 &  x40 &  x46 &  x47 &  x50 &  x56 &  x68 &  x69 &  x70 &  x76 &  x77 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x5 & ~x23 & ~x24 & ~x25 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x65 & ~x72 & ~x73 & ~x83 & ~x85 & ~x94;
assign c3319 =  x3;
assign c3323 =  x3 &  x72;
assign c3325 = ~x2;
assign c3327 = ~x2;
assign c3329 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c3331 =  x2 &  x6 &  x16 &  x77 & ~x43 & ~x84;
assign c3333 = ~x2 & ~x7;
assign c3335 =  x31 &  x58 & ~x2 & ~x32 & ~x62;
assign c3337 =  x0 &  x2 &  x4 &  x26 &  x46 &  x59 &  x67 &  x77 &  x78 &  x79 &  x80 &  x86 &  x88 & ~x24 & ~x43 & ~x54 & ~x62 & ~x64 & ~x73 & ~x75 & ~x92;
assign c3339 =  x4 &  x16 &  x18 &  x26 &  x39 &  x47 &  x48 &  x56 &  x57 &  x68 &  x69 &  x70 &  x78 & ~x32 & ~x35 & ~x45 & ~x62 & ~x63 & ~x64 & ~x82 & ~x84 & ~x85 & ~x93;
assign c3343 = ~x70;
assign c3345 =  x74;
assign c3347 =  x1;
assign c3349 =  x0 &  x2 &  x4 &  x16 &  x19 &  x26 &  x27 &  x28 &  x36 &  x39 &  x46 &  x48 &  x56 &  x57 &  x59 &  x66 &  x76 &  x86 & ~x23 & ~x25 & ~x33 & ~x34 & ~x43 & ~x45 & ~x72 & ~x73 & ~x74 & ~x82 & ~x83 & ~x93 & ~x94;
assign c3351 =  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x48 &  x56 &  x57 &  x66 &  x67 &  x69 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x5 & ~x23 & ~x24 & ~x44 & ~x45 & ~x52 & ~x53 & ~x55 & ~x62 & ~x65 & ~x72 & ~x83 & ~x84 & ~x85 & ~x94 & ~x95;
assign c3353 =  x1;
assign c3355 =  x1;
assign c3357 = ~x2 & ~x6;
assign c3359 =  x0 &  x4 &  x16 &  x47 &  x68 &  x86 & ~x6 & ~x24 & ~x65 & ~x75 & ~x82 & ~x94;
assign c3361 = ~x70;
assign c3363 = ~x6;
assign c3365 =  x2 &  x3;
assign c3367 =  x43;
assign c3369 =  x52;
assign c3371 =  x73;
assign c3375 = ~x60;
assign c3377 =  x6 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c3379 =  x84;
assign c3381 =  x83;
assign c3387 =  x52;
assign c3389 =  x1;
assign c3391 =  x0 &  x4 &  x16 &  x17 &  x26 &  x28 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x60 &  x67 &  x78 & ~x6 & ~x45 & ~x55 & ~x65 & ~x73 & ~x85 & ~x94;
assign c3393 = ~x60;
assign c3395 =  x2 &  x3 &  x5 &  x77;
assign c3397 =  x73;
assign c3399 = ~x2 & ~x4;
assign c3401 =  x6 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x1 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c3403 =  x43;
assign c3405 = ~x50;
assign c3407 =  x16 &  x18 &  x20 &  x26 &  x27 &  x28 &  x29 &  x31 &  x36 &  x38 &  x39 &  x40 &  x41 &  x48 &  x49 &  x56 &  x57 &  x59 &  x60 &  x66 &  x67 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x87 &  x89 &  x90 & ~x0 & ~x22 & ~x24 & ~x25 & ~x33 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x64 & ~x65 & ~x72 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c3409 =  x1;
assign c3411 =  x42;
assign c3413 =  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x91 & ~x1 & ~x8 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c3415 = ~x18;
assign c3417 =  x1;
assign c3419 =  x52;
assign c3421 = ~x40;
assign c3423 = ~x39;
assign c3425 =  x0 &  x2 &  x4 &  x17 &  x20 &  x26 &  x28 &  x29 &  x30 &  x37 &  x38 &  x46 &  x47 &  x48 &  x49 &  x57 &  x58 &  x60 &  x66 &  x69 &  x76 &  x79 &  x86 &  x87 &  x88 &  x90 & ~x1 & ~x22 & ~x23 & ~x33 & ~x34 & ~x35 & ~x55 & ~x62 & ~x65 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c3427 = ~x2 & ~x4;
assign c3429 =  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x1 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c3431 =  x3 &  x6 &  x17 &  x46 &  x76 & ~x5 & ~x35 & ~x75;
assign c3433 =  x52;
assign c3435 = ~x88;
assign c3437 = ~x60;
assign c3439 = ~x7;
assign c3441 =  x53;
assign c3443 = ~x3;
assign c3445 = ~x2 & ~x5;
assign c3447 =  x74;
assign c3449 = ~x2;
assign c3451 =  x0 &  x2 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x47 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x86 &  x88 &  x89 & ~x1 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x92 & ~x93 & ~x94 & ~x95;
assign c3453 = ~x2 & ~x92;
assign c3455 =  x64;
assign c3457 =  x2 &  x3 &  x6;
assign c3459 =  x9 &  x20 &  x26 &  x30 &  x31 &  x36 &  x37 &  x39 &  x40 &  x57 &  x61 &  x68 &  x70 &  x76 &  x90 & ~x22 & ~x64 & ~x72 & ~x83 & ~x94;
assign c3461 = ~x68;
assign c3463 =  x1;
assign c3465 = ~x2;
assign c3467 =  x1;
assign c3469 =  x91;
assign c3471 = ~x50;
assign c3473 = ~x70;
assign c3475 =  x2 &  x16 &  x18 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x90 & ~x1 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c3477 =  x6 &  x42 &  x90 &  x91;
assign c3479 =  x52;
assign c3481 =  x1;
assign c3483 =  x1;
assign c3485 = ~x79;
assign c3487 =  x0 &  x4 & ~x7 & ~x45;
assign c3489 =  x72;
assign c3491 =  x2 &  x3 &  x5;
assign c3493 =  x2 &  x3 &  x5;
assign c3495 =  x2 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x70 &  x71 &  x77 &  x78 &  x86 &  x87 &  x89 &  x90 &  x91 & ~x1 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x65 & ~x72 & ~x74 & ~x75 & ~x81 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c3497 = ~x60;
assign c3499 =  x6 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x7 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x52 & ~x53 & ~x54 & ~x63 & ~x64 & ~x72 & ~x73 & ~x74 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c40 = ~x36;
assign c42 =  x0 &  x2 &  x3 &  x19 &  x21 &  x28 &  x31 &  x39 &  x47 &  x76 &  x80 &  x86 &  x91 & ~x1 & ~x7 & ~x22 & ~x24 & ~x35 & ~x54 & ~x84;
assign c44 = ~x46;
assign c46 = ~x26;
assign c48 =  x67 &  x91 & ~x71;
assign c410 =  x0 &  x2 &  x3 &  x4 &  x16 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x52 & ~x55 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c412 =  x20 &  x26 &  x27 &  x29 &  x30 &  x37 &  x38 &  x39 &  x40 &  x59 &  x61 &  x62 &  x66 &  x67 &  x68 &  x69 &  x76 &  x78 &  x79 &  x88 &  x89 & ~x8 & ~x22 & ~x32 & ~x35 & ~x42 & ~x43 & ~x53 & ~x55 & ~x74 & ~x75 & ~x83 & ~x92 & ~x93 & ~x95;
assign c414 =  x5 &  x59 & ~x4 & ~x6 & ~x21 & ~x81 & ~x91;
assign c416 =  x24;
assign c418 =  x5 &  x17 &  x19 &  x20 &  x21 &  x26 &  x28 &  x29 &  x30 &  x31 &  x37 &  x40 &  x47 &  x56 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x81 &  x86 &  x87 &  x89 &  x90 &  x91 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x45 & ~x54 & ~x55 & ~x63 & ~x64 & ~x84 & ~x92 & ~x94 & ~x95;
assign c420 =  x21 &  x31 &  x42 &  x48 &  x91 & ~x43 & ~x83;
assign c422 = ~x17;
assign c424 =  x31 &  x47 & ~x58;
assign c426 = ~x58;
assign c428 = ~x17;
assign c430 =  x92;
assign c432 = ~x86;
assign c434 =  x50 &  x56 &  x59 &  x62 &  x63 & ~x32 & ~x42 & ~x54;
assign c436 = ~x28;
assign c438 =  x16 &  x21 &  x31 &  x38 &  x40 &  x50 &  x70 &  x71 &  x76 &  x77 &  x80 &  x91 & ~x4 & ~x10 & ~x35 & ~x75 & ~x84;
assign c440 = ~x77;
assign c442 =  x16 &  x20 &  x26 &  x27 &  x28 &  x30 &  x39 &  x46 &  x47 &  x48 &  x49 &  x66 &  x67 &  x68 &  x76 &  x77 &  x86 &  x88 &  x90 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x60 & ~x63 & ~x65 & ~x82 & ~x92 & ~x95;
assign c444 =  x48 &  x68 &  x69 &  x89 &  x90 & ~x4 & ~x33 & ~x44 & ~x52 & ~x60 & ~x83 & ~x95;
assign c446 =  x1 &  x17 &  x19 &  x20 &  x26 &  x29 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x59 &  x66 &  x67 &  x69 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x3 & ~x4 & ~x14 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x74 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c448 =  x82;
assign c450 =  x5 & ~x4 & ~x69;
assign c452 = ~x76;
assign c454 = ~x36;
assign c456 =  x0 &  x2 &  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x57 &  x58 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x1 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x42 & ~x43 & ~x44 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x95;
assign c458 =  x82;
assign c462 = ~x66;
assign c464 =  x16 &  x17 &  x20 &  x26 &  x27 &  x29 &  x30 &  x31 &  x36 &  x46 &  x47 &  x52 &  x67 &  x77 &  x86 &  x88 &  x90 & ~x0 & ~x2 & ~x3 & ~x4 & ~x22 & ~x23 & ~x25 & ~x32 & ~x33 & ~x35 & ~x44 & ~x45 & ~x65 & ~x74 & ~x84 & ~x92 & ~x94 & ~x95;
assign c466 = ~x19;
assign c468 =  x1 &  x7 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x3 & ~x4 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c470 =  x18 &  x19 &  x36 &  x38 &  x46 &  x59 &  x67 &  x78 & ~x22 & ~x33 & ~x41 & ~x45 & ~x54 & ~x70 & ~x71 & ~x72 & ~x73 & ~x82 & ~x84 & ~x85 & ~x94 & ~x95;
assign c472 =  x10 &  x63 & ~x54;
assign c474 = ~x86;
assign c476 = ~x27;
assign c478 =  x75 & ~x36;
assign c480 = ~x66;
assign c482 =  x0 &  x2 &  x3 &  x5 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x31 &  x36 &  x37 &  x39 &  x46 &  x56 &  x66 &  x67 &  x68 &  x76 &  x77 &  x78 &  x79 &  x80 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x44 & ~x45 & ~x55 & ~x65 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c484 = ~x87;
assign c486 = ~x86;
assign c488 =  x32 &  x82;
assign c490 =  x29 &  x47 &  x67 &  x77 &  x86 &  x87 &  x89 & ~x24 & ~x32 & ~x33 & ~x41 & ~x43 & ~x70 & ~x74 & ~x81 & ~x82 & ~x92 & ~x94;
assign c492 = ~x17;
assign c494 =  x45;
assign c496 =  x23;
assign c498 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x3 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4100 =  x0 &  x2 &  x3 &  x5 &  x16 &  x17 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x36 &  x37 &  x38 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x55 & ~x65 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x95;
assign c4102 = ~x48;
assign c4104 =  x1 &  x5 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x56 &  x57 &  x66 &  x67 &  x68 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x3 & ~x4 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4106 = ~x76;
assign c4108 =  x0 &  x2 &  x3 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x57 &  x58 &  x59 &  x66 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x6 & ~x23 & ~x24 & ~x32 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x71 & ~x73 & ~x82 & ~x83 & ~x84 & ~x92 & ~x95;
assign c4110 =  x55;
assign c4112 = ~x17;
assign c4116 =  x5 & ~x70;
assign c4118 = ~x40;
assign c4120 = ~x48;
assign c4122 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x29 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x57 &  x59 &  x60 &  x61 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x23 & ~x24 & ~x25 & ~x32 & ~x43 & ~x44 & ~x63 & ~x65 & ~x71 & ~x72 & ~x73 & ~x74 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x95;
assign c4124 =  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x50 &  x51 &  x57 &  x58 &  x66 &  x67 &  x77 &  x78 &  x88 &  x90 & ~x6 & ~x22 & ~x24 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x54 & ~x55 & ~x64 & ~x65 & ~x71 & ~x72 & ~x82 & ~x83 & ~x85 & ~x92 & ~x93;
assign c4126 =  x0 &  x2 &  x3 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x46 &  x47 &  x48 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x62 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x80 &  x86 &  x87 &  x88 &  x90 & ~x1 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x95;
assign c4128 = ~x76;
assign c4130 = ~x76;
assign c4132 =  x0 &  x2 &  x3 &  x5 &  x16 &  x17 &  x19 &  x20 &  x27 &  x29 &  x30 &  x38 &  x48 &  x76 &  x77 &  x90 & ~x1 & ~x4 & ~x22 & ~x34 & ~x35 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4136 = ~x86;
assign c4138 = ~x69;
assign c4140 = ~x86;
assign c4142 = ~x16;
assign c4144 = ~x88;
assign c4146 =  x0 &  x2 &  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x65 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4148 = ~x46;
assign c4150 =  x31 & ~x58;
assign c4152 =  x0 &  x2 &  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x61 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x54 & ~x55 & ~x65 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4154 = ~x87;
assign c4156 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x3 & ~x4 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4160 =  x50 &  x73 &  x80 &  x91 & ~x54 & ~x83 & ~x84;
assign c4162 =  x25;
assign c4164 =  x73;
assign c4166 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x3 & ~x4 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4168 =  x16 &  x17 &  x26 &  x36 &  x39 &  x49 &  x67 &  x76 &  x77 &  x78 &  x80 &  x86 &  x89 &  x90 & ~x6 & ~x23 & ~x24 & ~x25 & ~x43 & ~x53 & ~x60 & ~x62 & ~x64 & ~x75 & ~x84 & ~x85 & ~x93;
assign c4170 =  x0 &  x2 &  x3 &  x5 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x36 &  x37 &  x38 &  x46 &  x47 &  x56 &  x57 &  x58 &  x66 &  x67 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x64 & ~x65 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x94 & ~x95;
assign c4172 =  x5 & ~x69;
assign c4174 =  x0 &  x2 &  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x7 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4176 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x21 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x3 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4178 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x59 &  x60 &  x61 &  x66 &  x67 &  x68 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x3 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4180 =  x0 &  x2 &  x3 &  x5 &  x16 &  x18 &  x19 &  x20 &  x26 &  x28 &  x29 &  x36 &  x37 &  x38 &  x57 &  x66 &  x77 &  x86 &  x88 &  x90 & ~x1 & ~x4 & ~x22 & ~x23 & ~x24 & ~x32 & ~x33 & ~x35 & ~x42 & ~x44 & ~x45 & ~x55 & ~x64 & ~x83 & ~x84 & ~x85 & ~x95;
assign c4182 =  x34;
assign c4184 = ~x86;
assign c4186 =  x31 & ~x43 & ~x58;
assign c4188 =  x16 &  x18 &  x19 &  x20 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x60 &  x62 &  x66 &  x67 &  x68 &  x69 &  x76 &  x78 &  x79 &  x80 &  x87 &  x89 &  x90 & ~x5 & ~x7 & ~x22 & ~x23 & ~x32 & ~x33 & ~x45 & ~x74 & ~x75 & ~x82 & ~x83 & ~x85 & ~x92 & ~x93 & ~x94;
assign c4190 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x76 &  x77 &  x78 &  x79 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x3 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4192 =  x1 &  x16 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x80 &  x86 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x3 & ~x4 & ~x11 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4194 =  x0 &  x2 &  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x59 &  x66 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x71 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4196 = ~x18;
assign c4198 =  x16 &  x17 &  x19 &  x26 &  x30 &  x38 &  x39 &  x46 &  x48 &  x49 &  x50 &  x56 &  x66 &  x67 &  x69 &  x80 &  x89 & ~x6 & ~x22 & ~x53 & ~x54 & ~x60 & ~x61 & ~x63 & ~x65 & ~x83 & ~x84 & ~x85 & ~x93;
assign c4200 = ~x66;
assign c4202 =  x73 &  x80;
assign c4204 =  x0 &  x2 &  x5 &  x16 &  x18 &  x19 &  x20 &  x26 &  x28 &  x29 &  x36 &  x37 &  x38 &  x39 &  x47 &  x48 &  x49 &  x56 &  x57 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x4 & ~x24 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x53 & ~x54 & ~x65 & ~x74 & ~x75 & ~x83 & ~x85 & ~x93 & ~x94;
assign c4206 =  x0 &  x2 &  x3 &  x5 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x57 &  x66 &  x67 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4210 =  x55;
assign c4212 =  x16 &  x21 &  x38 &  x40 &  x67 &  x69 &  x72 &  x77 &  x90 & ~x6 & ~x23 & ~x25 & ~x55 & ~x65 & ~x84 & ~x85 & ~x93;
assign c4214 =  x18 &  x19 &  x38 &  x46 &  x49 &  x56 &  x57 &  x62 &  x77 &  x78 &  x87 & ~x22 & ~x24 & ~x33 & ~x34 & ~x35 & ~x43 & ~x54 & ~x55 & ~x71 & ~x73 & ~x74 & ~x83 & ~x84 & ~x94;
assign c4216 = ~x27 & ~x76;
assign c4218 =  x19 &  x20 &  x21 &  x27 &  x37 &  x38 &  x39 &  x56 &  x66 &  x69 &  x80 &  x88 & ~x6 & ~x23 & ~x24 & ~x51 & ~x53 & ~x54 & ~x65 & ~x84 & ~x93 & ~x95;
assign c4220 =  x16 &  x17 &  x18 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x6 & ~x21 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x45 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x91 & ~x93 & ~x94;
assign c4222 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x21 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x41 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x91 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4224 = ~x28 & ~x67;
assign c4226 =  x0 &  x2 &  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x46 &  x48 &  x49 &  x56 &  x57 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x11 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x65 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4228 =  x82;
assign c4230 = ~x76;
assign c4232 = ~x0 & ~x2 & ~x4 & ~x70;
assign c4234 =  x0 &  x2 &  x3 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x57 &  x58 &  x59 &  x66 &  x68 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x61 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4236 =  x0 &  x2 &  x3 &  x5 &  x16 &  x18 &  x19 &  x20 &  x29 &  x30 &  x37 &  x56 &  x57 &  x66 &  x67 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x4 & ~x22 & ~x24 & ~x32 & ~x43 & ~x44 & ~x45 & ~x53 & ~x74 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x95;
assign c4238 = ~x56;
assign c4240 =  x16 &  x17 &  x18 &  x20 &  x26 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x47 &  x48 &  x66 &  x67 &  x68 &  x69 &  x71 &  x72 &  x76 &  x78 &  x80 &  x87 &  x90 & ~x0 & ~x2 & ~x3 & ~x4 & ~x22 & ~x23 & ~x24 & ~x34 & ~x35 & ~x45 & ~x55 & ~x65 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c4242 = ~x36;
assign c4244 =  x61 & ~x4 & ~x54 & ~x71;
assign c4246 = ~x56;
assign c4248 = ~x76;
assign c4250 =  x1 &  x16 &  x18 &  x19 &  x20 &  x26 &  x27 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x3 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x34 & ~x35 & ~x41 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x54 & ~x55 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4252 =  x28 &  x31 &  x50 &  x59 &  x73 & ~x92;
assign c4254 =  x2 &  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x40 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x59 &  x66 &  x67 &  x68 &  x76 &  x77 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x9 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x74 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x95;
assign c4256 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x3 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x55 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4258 =  x45;
assign c4262 = ~x58;
assign c4264 = ~x66;
assign c4266 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x3 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4270 =  x20 &  x27 &  x28 &  x30 &  x37 &  x40 &  x47 &  x57 &  x67 &  x68 &  x80 &  x90 &  x91 & ~x6 & ~x22 & ~x23 & ~x33 & ~x34 & ~x44 & ~x45 & ~x82 & ~x83 & ~x84 & ~x92 & ~x93;
assign c4272 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x30 &  x36 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x3 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x35 & ~x41 & ~x42 & ~x43 & ~x52 & ~x54 & ~x55 & ~x63 & ~x64 & ~x73 & ~x74 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4274 =  x63 & ~x42 & ~x54 & ~x92;
assign c4276 = ~x26;
assign c4278 =  x17 &  x30 &  x36 &  x39 &  x41 &  x59 &  x60 &  x62 &  x77 & ~x4 & ~x23 & ~x32 & ~x33 & ~x43 & ~x55 & ~x74 & ~x83 & ~x85 & ~x94;
assign c4280 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x3 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4282 = ~x76;
assign c4284 = ~x56;
assign c4286 = ~x58;
assign c4288 =  x0 &  x2 &  x3 &  x16 &  x29 &  x30 &  x36 &  x37 &  x38 &  x40 &  x46 &  x47 &  x49 &  x50 &  x51 &  x56 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x90 & ~x1 & ~x21 & ~x22 & ~x23 & ~x32 & ~x33 & ~x42 & ~x43 & ~x44 & ~x52 & ~x53 & ~x55 & ~x64 & ~x75 & ~x82 & ~x93 & ~x95;
assign c4290 = ~x76;
assign c4292 = ~x26;
assign c4294 =  x31 &  x47 &  x67 &  x91 & ~x43 & ~x58;
assign c4296 =  x5 & ~x69;
assign c4298 =  x0 &  x2 &  x3 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x40 &  x47 &  x48 &  x56 &  x57 &  x59 &  x66 &  x67 &  x68 &  x76 &  x86 &  x87 &  x88 &  x90 & ~x5 & ~x22 & ~x25 & ~x32 & ~x33 & ~x34 & ~x43 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x94 & ~x95;
assign c4300 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x3 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4302 = ~x43 & ~x58;
assign c4304 = ~x86;
assign c4306 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 & ~x0 & ~x2 & ~x3 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4308 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x61 &  x62 &  x66 &  x68 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x3 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4310 =  x17 &  x18 &  x19 &  x20 &  x28 &  x29 &  x30 &  x46 &  x47 &  x49 &  x50 &  x56 &  x59 &  x60 &  x61 &  x62 &  x67 &  x68 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x90 & ~x4 & ~x23 & ~x24 & ~x32 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x64 & ~x72 & ~x73 & ~x74 & ~x82 & ~x84 & ~x93 & ~x94;
assign c4312 = ~x18;
assign c4314 =  x10 &  x63;
assign c4316 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x0 & ~x2 & ~x3 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4318 =  x0 &  x2 &  x3 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x46 &  x48 &  x49 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x77 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x5 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x65 & ~x74 & ~x75 & ~x82 & ~x83 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4320 = ~x66;
assign c4322 =  x16 &  x17 &  x18 &  x19 &  x20 &  x27 &  x28 &  x36 &  x38 &  x47 &  x48 &  x49 &  x57 &  x58 &  x59 &  x60 &  x66 &  x68 &  x76 &  x77 &  x78 &  x88 &  x89 &  x90 & ~x9 & ~x21 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x42 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x65 & ~x72 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x91 & ~x92 & ~x93 & ~x94;
assign c4324 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x21 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x56 &  x57 &  x58 &  x59 &  x60 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x3 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4328 =  x17 &  x18 &  x19 &  x20 &  x21 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x50 &  x56 &  x59 &  x60 &  x66 &  x67 &  x68 &  x70 &  x71 &  x72 &  x76 &  x77 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x22 & ~x23 & ~x25 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x55 & ~x74 & ~x75 & ~x83 & ~x84 & ~x92 & ~x93 & ~x94;
assign c4330 = ~x76;
assign c4332 =  x62 &  x63 & ~x42 & ~x43 & ~x45 & ~x54;
assign c4334 = ~x26;
assign c4336 = ~x77;
assign c4338 =  x0 &  x2 &  x3 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4340 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x0 & ~x2 & ~x3 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4342 =  x92;
assign c4344 = ~x86;
assign c4346 =  x21 &  x27 &  x72 & ~x6;
assign c4348 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x56 &  x57 &  x70 &  x77 &  x78 &  x79 &  x80 &  x81 &  x86 &  x87 &  x88 &  x90 & ~x0 & ~x2 & ~x3 & ~x4 & ~x24 & ~x25 & ~x33 & ~x35 & ~x44 & ~x45 & ~x55 & ~x65 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4350 = ~x28;
assign c4352 =  x34;
assign c4354 =  x0 &  x2 &  x3 &  x5 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x46 &  x47 &  x57 &  x58 &  x67 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x35 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x65 & ~x75 & ~x82 & ~x83 & ~x84 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4356 =  x64;
assign c4358 =  x91 & ~x59;
assign c4360 =  x16 &  x18 &  x26 &  x27 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x49 &  x67 &  x68 &  x76 &  x78 &  x86 &  x87 &  x88 & ~x6 & ~x24 & ~x32 & ~x34 & ~x35 & ~x43 & ~x45 & ~x60 & ~x64 & ~x65 & ~x75 & ~x82 & ~x93 & ~x94;
assign c4364 =  x75;
assign c4366 =  x0 &  x2 &  x3 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x5 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4368 =  x0 &  x2 &  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x30 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x89 &  x90 & ~x1 & ~x5 & ~x23 & ~x24 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4370 =  x0 &  x2 &  x3 &  x19 &  x20 &  x26 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x60 &  x66 &  x67 &  x68 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x90 & ~x1 & ~x22 & ~x25 & ~x32 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x73 & ~x74 & ~x75 & ~x82 & ~x85 & ~x92 & ~x93 & ~x94;
assign c4372 =  x95;
assign c4374 =  x18 &  x40 &  x48 &  x49 &  x62 &  x67 &  x68 &  x76 &  x80 & ~x3 & ~x4 & ~x35 & ~x45 & ~x53 & ~x54 & ~x75 & ~x82;
assign c4376 =  x2 &  x3 &  x5 &  x17 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x37 &  x38 &  x56 &  x57 &  x66 &  x68 &  x69 &  x70 &  x71 &  x77 &  x78 &  x79 &  x86 & ~x1 & ~x4 & ~x22 & ~x23 & ~x25 & ~x33 & ~x34 & ~x45 & ~x55 & ~x75 & ~x83 & ~x84 & ~x92 & ~x94 & ~x95;
assign c4378 = ~x16;
assign c4380 =  x16 &  x17 &  x18 &  x20 &  x26 &  x27 &  x30 &  x36 &  x37 &  x39 &  x40 &  x47 &  x48 &  x50 &  x57 &  x66 &  x67 &  x69 &  x77 &  x79 &  x87 &  x88 &  x89 & ~x4 & ~x23 & ~x25 & ~x33 & ~x35 & ~x44 & ~x45 & ~x52 & ~x53 & ~x60 & ~x61 & ~x63 & ~x65 & ~x75 & ~x83 & ~x85 & ~x93;
assign c4382 =  x64 & ~x6;
assign c4384 = ~x77;
assign c4386 =  x8 &  x19 &  x28 &  x47 &  x68 &  x76 &  x79 &  x86 &  x88 &  x89 &  x90 & ~x60 & ~x81;
assign c4388 =  x55;
assign c4390 =  x75;
assign c4392 =  x16 &  x17 &  x18 &  x19 &  x20 &  x27 &  x28 &  x29 &  x30 &  x37 &  x38 &  x46 &  x48 &  x57 &  x59 &  x60 &  x61 &  x62 &  x77 &  x78 &  x79 &  x86 &  x89 &  x90 & ~x4 & ~x22 & ~x23 & ~x32 & ~x33 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x74 & ~x82 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4394 =  x0 &  x2 &  x3 &  x5 &  x16 &  x17 &  x18 &  x19 &  x27 &  x36 &  x38 &  x47 &  x57 &  x67 &  x76 &  x86 &  x88 &  x89 &  x90 & ~x4 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x54 & ~x64 & ~x65 & ~x72 & ~x74 & ~x83 & ~x85 & ~x93 & ~x95;
assign c4396 =  x95;
assign c4398 =  x31 &  x47 & ~x58;
assign c4400 =  x32 &  x92;
assign c4402 =  x35;
assign c4404 =  x23 &  x45;
assign c4406 = ~x79;
assign c4408 =  x0 &  x2 &  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4410 = ~x58;
assign c4412 =  x0 &  x2 &  x3 &  x9 &  x16 &  x18 &  x19 &  x26 &  x27 &  x30 &  x31 &  x38 &  x40 &  x41 &  x46 &  x48 &  x50 &  x56 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 & ~x1 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x44 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x75 & ~x83 & ~x85 & ~x92 & ~x93 & ~x95;
assign c4414 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x49 &  x56 &  x66 &  x67 &  x68 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x3 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x64 & ~x65 & ~x71 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4416 = ~x48 & ~x70;
assign c4420 =  x75;
assign c4422 =  x17 &  x21 &  x29 &  x39 &  x41 &  x42 &  x46 &  x48 &  x57 &  x66 &  x68 &  x78 &  x80 &  x86 &  x91 & ~x22 & ~x23 & ~x61 & ~x62 & ~x63 & ~x84 & ~x93 & ~x95;
assign c4424 = ~x17;
assign c4428 =  x47 &  x48 &  x50 &  x59 &  x71 &  x73 &  x80 &  x86 &  x87 & ~x24 & ~x44 & ~x54 & ~x85 & ~x92;
assign c4430 = ~x66;
assign c4432 =  x0 &  x2 &  x3 &  x5 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x36 &  x37 &  x38 &  x46 &  x47 &  x56 &  x66 &  x76 &  x77 &  x78 &  x86 &  x88 &  x89 &  x90 & ~x1 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x45 & ~x54 & ~x55 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4434 =  x32;
assign c4436 = ~x66;
assign c4438 =  x50 &  x72 &  x73 &  x80 &  x91 & ~x54;
assign c4440 =  x7 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4442 =  x52 &  x67 & ~x70;
assign c4444 =  x1 &  x9 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x3 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x72 & ~x73 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c4446 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x21 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x56 &  x57 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x89 &  x90 & ~x0 & ~x2 & ~x3 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x64 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4448 = ~x18;
assign c4450 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x21 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x0 & ~x2 & ~x3 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x55 & ~x65 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c4452 =  x1 &  x16 &  x17 &  x18 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x40 &  x46 &  x47 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x87 &  x88 &  x90 & ~x0 & ~x2 & ~x3 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x43 & ~x44 & ~x53 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4454 = ~x87;
assign c4456 =  x16 &  x17 &  x18 &  x20 &  x21 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x42 &  x46 &  x47 &  x48 &  x56 &  x57 &  x66 &  x67 &  x68 &  x76 &  x77 &  x78 &  x79 &  x80 &  x87 &  x90 &  x91 & ~x22 & ~x23 & ~x25 & ~x33 & ~x34 & ~x35 & ~x44 & ~x54 & ~x61 & ~x62 & ~x63 & ~x64 & ~x65 & ~x84 & ~x85 & ~x93 & ~x94;
assign c4458 =  x62 & ~x4 & ~x43 & ~x71 & ~x83;
assign c4460 = ~x36;
assign c4462 =  x21 &  x52 &  x66 &  x67 & ~x7 & ~x45 & ~x74 & ~x92;
assign c4464 =  x75;
assign c4466 = ~x86;
assign c4470 =  x2 &  x3 &  x19 &  x20 &  x29 &  x31 &  x36 &  x47 &  x48 &  x76 &  x80 &  x90 & ~x25 & ~x60 & ~x63 & ~x94;
assign c4472 =  x1 &  x10 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x3 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4474 = ~x26;
assign c4476 =  x52;
assign c4478 =  x32 &  x82;
assign c4480 =  x0 &  x2 &  x3 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4482 =  x0 &  x2 &  x3 &  x5 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x46 &  x47 &  x66 &  x67 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x1 & ~x4 & ~x22 & ~x23 & ~x24 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94;
assign c4484 =  x10 &  x20 &  x26 &  x61 &  x62 &  x76 &  x78 &  x86 &  x90 & ~x6 & ~x44 & ~x82;
assign c4486 = ~x77;
assign c4488 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x3 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x61 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4490 = ~x16;
assign c4492 =  x31 &  x40 &  x51 & ~x60 & ~x72;
assign c4496 =  x65;
assign c4498 = ~x19;
assign c41 =  x2 & ~x3;
assign c43 =  x4 & ~x0;
assign c45 = ~x90;
assign c47 =  x54;
assign c49 =  x22;
assign c411 =  x4 & ~x3;
assign c413 =  x43;
assign c415 =  x0 &  x1 &  x16 &  x17 &  x26 &  x37 &  x66 &  x67 &  x78 &  x86 &  x89 & ~x23 & ~x25 & ~x32 & ~x44 & ~x54 & ~x85;
assign c417 =  x4 & ~x3;
assign c419 =  x3 &  x19 &  x27 &  x28 &  x29 &  x30 &  x36 &  x38 &  x46 &  x49 &  x50 &  x51 &  x59 &  x66 &  x67 &  x70 &  x79 &  x86 &  x87 & ~x25 & ~x43 & ~x62 & ~x63 & ~x65 & ~x74 & ~x75 & ~x83 & ~x85 & ~x94;
assign c421 = ~x20;
assign c423 =  x2 &  x16 &  x20 &  x26 &  x27 &  x28 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x56 &  x66 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x90 & ~x4 & ~x5 & ~x23 & ~x24 & ~x34 & ~x35 & ~x44 & ~x45 & ~x54 & ~x62 & ~x63 & ~x64 & ~x65 & ~x83 & ~x84 & ~x94 & ~x95;
assign c425 =  x83;
assign c427 =  x16 &  x20 &  x21 &  x36 &  x48 &  x58 &  x68 &  x70 &  x86 &  x89 &  x90 & ~x33 & ~x43 & ~x52 & ~x73 & ~x81 & ~x82 & ~x94;
assign c429 =  x2 &  x19 &  x21 &  x51 & ~x52;
assign c431 =  x4;
assign c433 =  x0 &  x28 &  x30 &  x49 &  x66 &  x78 & ~x3 & ~x43 & ~x84 & ~x92;
assign c435 =  x1 &  x4;
assign c437 = ~x38;
assign c439 =  x3 &  x16 &  x19 &  x26 &  x36 &  x46 &  x47 &  x56 &  x57 &  x66 &  x67 &  x76 & ~x2 & ~x64 & ~x74 & ~x75 & ~x84;
assign c441 =  x4 &  x5 &  x30 &  x88 & ~x55 & ~x83 & ~x84;
assign c443 =  x81 & ~x91;
assign c445 =  x8 &  x16 &  x17 &  x18 &  x20 &  x26 &  x37 &  x39 &  x40 &  x47 &  x51 &  x56 &  x57 &  x59 &  x66 &  x68 &  x69 &  x76 &  x80 &  x86 &  x90 & ~x7 & ~x35 & ~x43 & ~x53 & ~x54 & ~x55 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x93 & ~x95;
assign c447 = ~x2;
assign c449 = ~x39;
assign c451 = ~x20;
assign c455 =  x4 & ~x2;
assign c457 = ~x89;
assign c459 =  x74;
assign c461 = ~x90;
assign c463 =  x93;
assign c465 =  x16 &  x18 &  x20 &  x26 &  x31 &  x36 &  x38 &  x40 &  x46 &  x56 &  x67 &  x70 &  x86 &  x89 &  x90 & ~x6 & ~x7 & ~x22 & ~x24 & ~x62 & ~x63 & ~x73 & ~x75 & ~x84 & ~x93;
assign c467 =  x92;
assign c469 =  x53 & ~x9;
assign c471 =  x17 &  x19 &  x26 &  x27 &  x29 &  x30 &  x31 &  x37 &  x40 &  x59 &  x60 &  x61 &  x67 &  x70 &  x89 & ~x62 & ~x63 & ~x73 & ~x82 & ~x83 & ~x84 & ~x85;
assign c473 = ~x30;
assign c475 =  x4 &  x6 &  x7;
assign c477 =  x3 &  x16 &  x17 &  x18 &  x26 &  x27 &  x28 &  x36 &  x46 &  x47 &  x48 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x69 &  x70 &  x77 &  x78 &  x79 &  x80 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x23 & ~x25 & ~x34 & ~x35 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93;
assign c479 =  x4 & ~x2;
assign c481 =  x19 &  x26 &  x36 &  x39 &  x46 &  x47 &  x59 &  x60 &  x66 &  x67 &  x68 &  x88 & ~x1 & ~x4 & ~x45 & ~x62 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x84;
assign c483 =  x56 & ~x1 & ~x3;
assign c485 =  x5 &  x18 &  x19 &  x20 &  x26 &  x29 &  x30 &  x36 &  x37 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x59 &  x60 &  x67 &  x68 &  x69 &  x76 &  x77 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x74 & ~x75 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c487 = ~x90;
assign c489 =  x6 &  x8 &  x17 &  x19 &  x20 &  x28 &  x30 &  x38 &  x46 &  x57 &  x58 &  x66 &  x69 &  x77 &  x89 &  x91 & ~x32 & ~x42 & ~x44 & ~x54 & ~x74 & ~x75 & ~x85 & ~x92;
assign c491 = ~x29;
assign c493 =  x3 &  x46 &  x56 &  x70 &  x78 &  x89 & ~x2;
assign c495 =  x6 &  x16 &  x18 &  x50 &  x60 &  x67 &  x86 & ~x1 & ~x5 & ~x34;
assign c497 =  x17 &  x18 &  x20 &  x21 &  x27 &  x30 &  x36 &  x37 &  x38 &  x46 &  x47 &  x48 &  x50 &  x58 &  x66 &  x67 &  x68 &  x76 &  x86 &  x87 &  x88 &  x90 & ~x22 & ~x24 & ~x34 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x65 & ~x72 & ~x74 & ~x75 & ~x81 & ~x83 & ~x84 & ~x85;
assign c499 = ~x90;
assign c4101 =  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x56 &  x66 &  x67 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x4 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x64 & ~x65 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4103 =  x0 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x4 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x55 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4105 = ~x90;
assign c4109 =  x84;
assign c4111 =  x3 &  x19 &  x27 &  x28 &  x29 &  x30 &  x46 &  x47 &  x56 &  x57 &  x58 &  x67 &  x68 &  x76 &  x86 &  x87 &  x88 &  x89 & ~x2 & ~x22 & ~x34 & ~x85 & ~x94;
assign c4113 =  x33;
assign c4115 =  x22;
assign c4117 = ~x20;
assign c4119 =  x22;
assign c4121 =  x22;
assign c4123 =  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x36 &  x46 &  x47 &  x56 &  x66 &  x67 &  x68 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x34 & ~x35 & ~x43 & ~x45 & ~x53 & ~x54 & ~x55 & ~x74 & ~x75 & ~x83 & ~x84 & ~x93 & ~x94 & ~x95;
assign c4125 =  x6 &  x7 &  x16 &  x17 &  x18 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x66 &  x76 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x22 & ~x24 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x74 & ~x75 & ~x82 & ~x84 & ~x85 & ~x94 & ~x95;
assign c4127 =  x5 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4129 =  x3 &  x16 &  x17 &  x18 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x46 &  x47 &  x48 &  x56 &  x66 &  x67 &  x68 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x0 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x55 & ~x63 & ~x64 & ~x65 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4131 =  x0 &  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x56 &  x66 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x4 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x65 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4133 =  x4 &  x5 &  x16 &  x17 &  x18 &  x28 &  x29 &  x30 &  x37 &  x46 &  x47 &  x56 &  x76 &  x77 &  x86 &  x89 &  x90 & ~x23 & ~x33 & ~x34 & ~x85;
assign c4135 =  x83;
assign c4137 =  x3 &  x28 &  x58 &  x86 & ~x2 & ~x23 & ~x33 & ~x85;
assign c4139 =  x43;
assign c4141 = ~x39;
assign c4143 = ~x49 & ~x60;
assign c4145 =  x92;
assign c4147 =  x4 & ~x3;
assign c4149 =  x0 &  x17 &  x18 &  x19 &  x27 &  x39 &  x46 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x76 &  x78 &  x87 &  x88 &  x90 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x34 & ~x84 & ~x85 & ~x92 & ~x94 & ~x95;
assign c4151 =  x33;
assign c4153 =  x10 &  x16 &  x19 &  x26 &  x29 &  x36 &  x38 &  x40 &  x41 &  x49 &  x50 &  x51 &  x56 &  x57 &  x59 &  x60 &  x76 &  x78 &  x79 & ~x24 & ~x32 & ~x34 & ~x35 & ~x62 & ~x64 & ~x65 & ~x75;
assign c4155 = ~x3;
assign c4157 =  x1 &  x4;
assign c4159 =  x4 &  x5 &  x17 &  x19 &  x20 &  x26 &  x29 &  x36 &  x37 &  x39 &  x47 &  x56 &  x86 & ~x33 & ~x34 & ~x43 & ~x44 & ~x45 & ~x83 & ~x84 & ~x94;
assign c4161 = ~x20;
assign c4163 =  x3 &  x18 &  x67 &  x68 &  x88 &  x90 & ~x2 & ~x34 & ~x43 & ~x94 & ~x95;
assign c4165 =  x1 &  x2 &  x18 &  x26 &  x37 &  x49 &  x57 &  x66 &  x67 &  x76 & ~x23 & ~x25 & ~x32 & ~x35 & ~x45 & ~x54 & ~x64 & ~x85;
assign c4167 = ~x1 & ~x3;
assign c4169 =  x74;
assign c4171 =  x43;
assign c4173 = ~x8 & ~x40 & ~x82;
assign c4175 = ~x3;
assign c4177 =  x4 &  x5 &  x16 &  x18 &  x19 &  x28 &  x29 &  x37 &  x38 &  x46 &  x47 &  x56 &  x66 &  x79 &  x87 &  x88 &  x90 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x83 & ~x85 & ~x94;
assign c4179 = ~x90;
assign c4181 =  x6 &  x8 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4183 = ~x1 & ~x3;
assign c4185 =  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x56 &  x66 &  x67 &  x76 &  x77 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x64 & ~x65 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4187 = ~x89;
assign c4189 = ~x20;
assign c4191 = ~x20;
assign c4193 =  x94;
assign c4195 =  x5 &  x16 &  x18 &  x19 &  x28 &  x56 &  x67 &  x68 &  x79 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x2 & ~x23 & ~x33 & ~x34 & ~x43 & ~x44 & ~x63 & ~x72 & ~x73 & ~x74 & ~x84 & ~x94;
assign c4197 =  x4 &  x5 &  x17 &  x18 &  x27 &  x28 &  x29 &  x30 &  x37 &  x39 &  x46 &  x66 &  x77 &  x90 & ~x55 & ~x83 & ~x85 & ~x94;
assign c4199 =  x92;
assign c4203 = ~x38;
assign c4205 =  x3 &  x17 &  x26 &  x36 &  x37 &  x39 &  x47 &  x58 &  x59 &  x66 &  x68 &  x79 &  x89 &  x90 & ~x0 & ~x54 & ~x75 & ~x85 & ~x92 & ~x94;
assign c4207 =  x19 &  x36 &  x39 &  x87 &  x88 & ~x0 & ~x1 & ~x95;
assign c4209 =  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x56 &  x66 &  x67 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x4 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x65 & ~x73 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4211 =  x17 &  x18 &  x29 &  x30 &  x36 &  x37 &  x39 &  x40 &  x41 &  x46 &  x47 &  x59 &  x76 &  x77 &  x87 & ~x4 & ~x24 & ~x32 & ~x33 & ~x35 & ~x52 & ~x53 & ~x54 & ~x63 & ~x74 & ~x75 & ~x81 & ~x85 & ~x93 & ~x95;
assign c4213 = ~x67;
assign c4217 =  x5 &  x17 &  x20 &  x27 &  x36 &  x37 &  x38 &  x40 &  x41 &  x46 &  x49 &  x50 &  x56 &  x58 &  x60 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x89 &  x90 & ~x22 & ~x23 & ~x24 & ~x25 & ~x43 & ~x45 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x94;
assign c4219 =  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x46 &  x47 &  x48 &  x56 &  x57 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x45 & ~x55 & ~x65 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4221 = ~x47;
assign c4223 =  x81 & ~x21;
assign c4225 =  x4 & ~x2;
assign c4227 =  x4 & ~x2;
assign c4229 =  x83;
assign c4231 =  x92;
assign c4233 =  x32 & ~x82;
assign c4235 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x61 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4237 = ~x79;
assign c4239 =  x22;
assign c4241 = ~x79;
assign c4243 =  x0 &  x17 &  x18 &  x20 &  x30 &  x37 &  x38 &  x56 &  x66 &  x76 &  x87 &  x90 & ~x2 & ~x33 & ~x44 & ~x53 & ~x55 & ~x83 & ~x94;
assign c4245 = ~x1 & ~x2;
assign c4247 = ~x30;
assign c4249 =  x19 &  x20 &  x27 &  x28 &  x37 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x51 &  x56 &  x57 &  x58 &  x59 &  x61 &  x67 &  x68 &  x69 &  x70 &  x76 &  x78 &  x79 &  x86 &  x88 &  x89 & ~x23 & ~x24 & ~x25 & ~x32 & ~x34 & ~x35 & ~x43 & ~x44 & ~x55 & ~x62 & ~x63 & ~x75 & ~x84 & ~x85 & ~x94 & ~x95;
assign c4251 =  x16 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x30 &  x36 &  x37 &  x38 &  x39 &  x47 &  x48 &  x49 &  x50 &  x56 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x35 & ~x43 & ~x44 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4253 = ~x68;
assign c4255 =  x93;
assign c4257 =  x2 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x58 &  x59 &  x66 &  x67 &  x68 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x90 & ~x0 & ~x22 & ~x23 & ~x25 & ~x34 & ~x35 & ~x44 & ~x45 & ~x53 & ~x54 & ~x84;
assign c4259 =  x22;
assign c4261 = ~x68;
assign c4265 =  x0 &  x5 &  x16 &  x17 &  x19 &  x26 &  x28 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x70 &  x76 &  x77 &  x78 &  x87 &  x89 &  x90 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x35 & ~x45 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93;
assign c4267 =  x16 &  x18 &  x36 &  x47 &  x66 &  x76 &  x88 &  x89 & ~x0 & ~x1 & ~x23 & ~x55 & ~x84;
assign c4269 =  x32;
assign c4271 =  x17 &  x18 &  x19 &  x20 &  x26 &  x28 &  x29 &  x36 &  x39 &  x48 &  x49 &  x50 &  x56 &  x59 &  x60 &  x67 &  x68 &  x69 &  x70 &  x79 &  x80 &  x87 &  x89 &  x90 &  x91 & ~x6 & ~x23 & ~x25 & ~x33 & ~x34 & ~x35 & ~x64 & ~x72 & ~x73 & ~x93 & ~x95;
assign c4273 =  x4 &  x5 &  x17 &  x18 &  x19 &  x27 &  x37 &  x77 &  x89 & ~x23 & ~x24 & ~x34 & ~x43 & ~x55 & ~x85 & ~x92 & ~x93 & ~x95;
assign c4275 =  x92;
assign c4277 =  x54;
assign c4279 =  x2 &  x18 &  x19 &  x27 &  x28 &  x30 &  x37 &  x38 &  x46 &  x57 &  x58 &  x66 &  x67 &  x68 &  x76 &  x77 &  x78 &  x79 &  x87 &  x88 &  x90 & ~x0 & ~x33 & ~x34 & ~x35 & ~x43 & ~x45 & ~x53 & ~x55 & ~x64 & ~x65 & ~x75;
assign c4281 = ~x49 & ~x82;
assign c4283 =  x17 &  x31 &  x39 &  x40 &  x48 &  x56 &  x58 &  x59 &  x60 &  x66 &  x71 &  x76 & ~x24 & ~x25 & ~x34 & ~x52 & ~x54 & ~x75 & ~x81 & ~x92 & ~x94;
assign c4285 =  x1 &  x2 &  x87 & ~x22;
assign c4287 =  x2 & ~x5 & ~x80;
assign c4289 =  x33;
assign c4291 = ~x90;
assign c4293 =  x0 &  x17 &  x18 &  x27 &  x28 &  x30 &  x37 &  x46 &  x56 &  x58 &  x66 &  x67 &  x68 &  x77 &  x79 &  x86 &  x89 &  x90 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x44 & ~x54 & ~x55 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4295 = ~x20;
assign c4297 =  x3 &  x20 &  x29 &  x37 &  x67 &  x76 &  x77 &  x86 & ~x2 & ~x35 & ~x75 & ~x84 & ~x85 & ~x95;
assign c4299 =  x54;
assign c4301 =  x0 &  x19 &  x20 &  x30 &  x58 &  x77 &  x87 &  x89 & ~x2 & ~x25 & ~x33 & ~x34 & ~x43 & ~x44 & ~x74 & ~x93 & ~x94;
assign c4303 =  x0 &  x16 &  x17 &  x18 &  x20 &  x26 &  x28 &  x36 &  x37 &  x39 &  x40 &  x46 &  x47 &  x66 &  x67 &  x76 &  x77 &  x78 &  x79 &  x86 &  x89 &  x90 & ~x3 & ~x22 & ~x24 & ~x25 & ~x33 & ~x44 & ~x55 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94;
assign c4305 =  x0 &  x16 &  x17 &  x18 &  x27 &  x28 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x79 &  x86 &  x88 &  x89 & ~x3 & ~x22 & ~x24 & ~x25 & ~x33 & ~x35 & ~x45 & ~x55 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94;
assign c4307 =  x4 & ~x2;
assign c4309 =  x19 &  x26 &  x69 &  x71 & ~x41 & ~x54 & ~x72 & ~x94;
assign c4311 =  x0 &  x16 &  x18 &  x20 &  x26 &  x27 &  x28 &  x30 &  x37 &  x46 &  x56 &  x66 &  x67 &  x68 &  x69 &  x70 &  x77 &  x78 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x45 & ~x55 & ~x75 & ~x82 & ~x83 & ~x84 & ~x93 & ~x95;
assign c4313 =  x53 & ~x21;
assign c4315 =  x82;
assign c4317 =  x22;
assign c4319 = ~x20;
assign c4321 =  x4 & ~x0;
assign c4323 =  x83;
assign c4325 =  x3 &  x74;
assign c4327 =  x0 &  x16 &  x18 &  x20 &  x29 &  x30 &  x36 &  x37 &  x39 &  x46 &  x48 &  x56 &  x57 &  x58 &  x66 &  x67 &  x70 &  x76 &  x77 &  x90 & ~x3 & ~x22 & ~x23 & ~x25 & ~x33 & ~x35 & ~x55 & ~x74 & ~x75 & ~x83 & ~x84;
assign c4329 = ~x20;
assign c4331 =  x6 &  x7 &  x16 &  x26 &  x29 &  x66 &  x77 & ~x1 & ~x5 & ~x24 & ~x32 & ~x73 & ~x84 & ~x85;
assign c4333 =  x0 &  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x46 &  x56 &  x66 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x4 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x55 & ~x63 & ~x64 & ~x65 & ~x83 & ~x84 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4335 =  x83;
assign c4337 =  x36 &  x46 &  x49 &  x51 &  x56 &  x59 &  x60 &  x66 &  x67 &  x71 &  x76 &  x86 &  x91 & ~x4 & ~x6 & ~x32 & ~x34 & ~x85;
assign c4339 =  x38 &  x39 &  x48 &  x59 &  x60 &  x70 &  x71 &  x77 &  x78 &  x90 & ~x1 & ~x24 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x75 & ~x84;
assign c4341 =  x5 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x53 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4343 = ~x1 & ~x3;
assign c4345 =  x22;
assign c4347 =  x74;
assign c4349 = ~x90;
assign c4351 =  x43;
assign c4355 =  x52;
assign c4357 =  x92;
assign c4361 =  x6 &  x27 &  x30 &  x46 &  x50 &  x56 &  x58 &  x68 & ~x1 & ~x25 & ~x43 & ~x84;
assign c4363 =  x17 &  x18 &  x27 &  x28 &  x29 &  x31 &  x38 &  x39 &  x41 &  x48 &  x49 &  x51 &  x58 &  x59 &  x60 &  x69 &  x76 &  x86 & ~x6 & ~x23 & ~x44 & ~x55 & ~x62 & ~x65 & ~x83;
assign c4365 =  x0 &  x1 &  x18 &  x30 &  x36 &  x46 &  x49 &  x58 &  x59 &  x68 &  x69 &  x86 &  x89;
assign c4367 =  x43;
assign c4369 =  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x46 &  x48 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x55 & ~x65 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4371 =  x0 &  x16 &  x17 &  x18 &  x26 &  x68 & ~x2 & ~x44 & ~x64 & ~x72;
assign c4375 =  x2 &  x17 &  x30 &  x49 &  x58 & ~x3 & ~x34 & ~x45 & ~x64;
assign c4377 =  x3 &  x16 &  x17 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x37 &  x46 &  x47 &  x56 &  x57 &  x66 &  x67 &  x68 &  x76 &  x78 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x23 & ~x24 & ~x25 & ~x35 & ~x45 & ~x55 & ~x64 & ~x65 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4379 = ~x30;
assign c4381 = ~x20;
assign c4383 =  x4 & ~x2;
assign c4385 =  x22;
assign c4387 =  x22;
assign c4389 =  x16 &  x18 &  x38 &  x41 &  x56 &  x69 &  x76 &  x78 &  x79 &  x80 &  x88 &  x89 &  x90 & ~x3 & ~x9 & ~x22 & ~x23 & ~x34 & ~x42 & ~x75 & ~x85;
assign c4391 =  x22;
assign c4393 = ~x57;
assign c4395 =  x4 & ~x0;
assign c4397 = ~x30;
assign c4399 =  x92;
assign c4401 =  x83;
assign c4403 = ~x67;
assign c4405 =  x16 &  x26 &  x27 &  x36 &  x71 &  x79 & ~x4 & ~x5 & ~x7 & ~x32 & ~x35 & ~x44 & ~x75;
assign c4407 =  x0 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x29 &  x30 &  x37 &  x38 &  x46 &  x47 &  x56 &  x66 &  x67 &  x68 &  x69 &  x77 &  x86 &  x87 &  x89 &  x90 & ~x2 & ~x22 & ~x25 & ~x34 & ~x35 & ~x73 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4409 =  x0 &  x38 &  x46 &  x48 &  x88 &  x89 & ~x3 & ~x53 & ~x94;
assign c4411 = ~x90;
assign c4413 =  x46 &  x87 & ~x21 & ~x51 & ~x61;
assign c4415 =  x92;
assign c4417 =  x0 &  x6 &  x7 &  x26 &  x29 &  x36 &  x66 &  x76 &  x78 &  x87 &  x90 & ~x5 & ~x23 & ~x34 & ~x45 & ~x83 & ~x84 & ~x85 & ~x94 & ~x95;
assign c4419 =  x43;
assign c4421 = ~x20;
assign c4423 =  x2 &  x18 &  x19 &  x20 &  x21 &  x37 &  x40 &  x51 &  x60 &  x67 &  x76 &  x77 &  x87 & ~x25 & ~x34 & ~x35 & ~x43 & ~x45 & ~x55 & ~x62 & ~x63 & ~x64 & ~x83 & ~x85;
assign c4425 =  x5 &  x6 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x48 &  x49 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x3 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x55 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4427 =  x54;
assign c4429 =  x0 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x66 &  x67 &  x68 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 & ~x4 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x55 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c4431 =  x5 &  x18 &  x20 &  x26 &  x27 &  x29 &  x30 &  x37 &  x40 &  x41 &  x47 &  x48 &  x49 &  x56 &  x58 &  x69 &  x76 &  x87 & ~x22 & ~x24 & ~x45 & ~x62 & ~x64 & ~x81 & ~x82 & ~x83 & ~x84 & ~x94 & ~x95;
assign c4433 = ~x67;
assign c4435 =  x4 & ~x0;
assign c4437 =  x2 &  x79 & ~x3 & ~x25;
assign c4439 =  x4 &  x5 &  x30 &  x36 &  x39 &  x46 &  x77 &  x88 &  x89 & ~x33 & ~x43 & ~x83;
assign c4441 = ~x90;
assign c4443 = ~x20;
assign c4445 =  x19 &  x20 &  x31 &  x37 &  x38 &  x46 &  x47 &  x49 &  x57 &  x58 &  x59 &  x70 &  x77 &  x78 &  x86 &  x87 & ~x4 & ~x10 & ~x23 & ~x25 & ~x34 & ~x52 & ~x53 & ~x54 & ~x55 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x94 & ~x95;
assign c4447 =  x93;
assign c4449 = ~x67;
assign c4451 =  x16 &  x18 &  x27 &  x28 &  x29 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x59 &  x70 &  x86 &  x87 &  x88 &  x91 & ~x6 & ~x24 & ~x34 & ~x35 & ~x55 & ~x65 & ~x73 & ~x74 & ~x83 & ~x92 & ~x93 & ~x95;
assign c4453 =  x1 &  x3 &  x17 &  x18 &  x37 &  x38 &  x46 &  x57 &  x59 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x86 &  x88 &  x89 & ~x34 & ~x35 & ~x44 & ~x45 & ~x65 & ~x85;
assign c4455 =  x0 &  x16 &  x17 &  x27 &  x29 &  x37 &  x77 &  x86 &  x89 & ~x4 & ~x5 & ~x23 & ~x25 & ~x33 & ~x34 & ~x35 & ~x45 & ~x52 & ~x54 & ~x55 & ~x63 & ~x83 & ~x93 & ~x94 & ~x95;
assign c4457 =  x43;
assign c4459 = ~x57;
assign c4461 =  x3 &  x46 &  x56 &  x57 &  x76 &  x77 &  x78 &  x87 &  x88 &  x90 & ~x2 & ~x23 & ~x33 & ~x34 & ~x45 & ~x65 & ~x74 & ~x84;
assign c4463 =  x16 &  x17 &  x19 &  x20 &  x26 &  x27 &  x29 &  x30 &  x36 &  x38 &  x39 &  x46 &  x47 &  x50 &  x56 &  x58 &  x59 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 &  x91 & ~x23 & ~x24 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x65 & ~x75 & ~x81 & ~x82 & ~x83 & ~x92 & ~x93 & ~x95;
assign c4465 =  x74;
assign c4467 =  x83;
assign c4469 =  x2 &  x17 &  x21 &  x27 &  x28 &  x29 &  x36 &  x37 &  x48 &  x50 &  x57 &  x66 & ~x25 & ~x35 & ~x43 & ~x54 & ~x62 & ~x63 & ~x73 & ~x92;
assign c4471 = ~x39;
assign c4473 =  x89 & ~x0 & ~x1 & ~x24 & ~x45;
assign c4475 =  x2 &  x48 &  x67 & ~x3 & ~x23 & ~x65;
assign c4477 =  x46 & ~x0 & ~x1 & ~x23 & ~x45;
assign c4479 =  x3 &  x16 &  x20 &  x26 &  x30 &  x36 &  x38 &  x56 &  x66 &  x76 &  x77 &  x78 &  x86 &  x88 & ~x0 & ~x24 & ~x44 & ~x62 & ~x63 & ~x65 & ~x75 & ~x85 & ~x94 & ~x95;
assign c4481 =  x81 & ~x41 & ~x60;
assign c4483 =  x2 &  x6 &  x7 &  x19 &  x20 &  x28 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x47 &  x56 &  x66 &  x68 &  x76 &  x80 &  x86 &  x87 &  x89 &  x90 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x54 & ~x55 & ~x63 & ~x65 & ~x75 & ~x82 & ~x94;
assign c4485 = ~x90;
assign c4487 =  x5 &  x70 & ~x2 & ~x51 & ~x72 & ~x73 & ~x92;
assign c4489 = ~x67;
assign c4491 =  x3 &  x17 &  x18 &  x19 &  x26 &  x29 &  x30 &  x36 &  x46 &  x56 &  x57 &  x66 &  x67 &  x76 &  x77 &  x78 &  x86 &  x88 &  x90 & ~x4 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x35 & ~x43 & ~x44 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x83 & ~x85 & ~x93 & ~x95;
assign c4493 =  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x56 &  x57 &  x58 &  x66 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x65 & ~x84 & ~x93 & ~x94 & ~x95;
assign c4495 = ~x30;
assign c4497 = ~x39;
assign c4499 =  x93;
assign c54 = ~x38;
assign c56 =  x1 &  x3 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c58 =  x1 &  x3 &  x4 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x37 &  x38 &  x46 &  x47 &  x48 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x90 & ~x2 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x74 & ~x82 & ~x83 & ~x84 & ~x85 & ~x93 & ~x95;
assign c510 =  x1 &  x5 &  x6 &  x7 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x61 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c512 =  x19 &  x38 &  x42 &  x52 & ~x22 & ~x54 & ~x83;
assign c514 =  x0 &  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x40 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x89 &  x90 & ~x2 & ~x3 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c516 =  x1 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c518 =  x0 &  x1 &  x4 &  x16 &  x26 &  x27 &  x28 &  x36 &  x39 &  x40 &  x56 &  x68 &  x70 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x90 & ~x3 & ~x5 & ~x25 & ~x33 & ~x34 & ~x44 & ~x73 & ~x74 & ~x75 & ~x85 & ~x92;
assign c520 =  x1 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x6 & ~x7 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c522 =  x0 &  x1 &  x4 &  x16 &  x29 &  x30 &  x37 &  x38 &  x57 &  x68 &  x78 &  x79 &  x87 &  x88 &  x90 & ~x2 & ~x5 & ~x22 & ~x24 & ~x25 & ~x43 & ~x45 & ~x54 & ~x65 & ~x72 & ~x74 & ~x81 & ~x95;
assign c524 =  x33;
assign c526 =  x85;
assign c528 =  x1 &  x3 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x47 &  x48 &  x49 &  x50 &  x57 &  x58 &  x59 &  x66 &  x68 &  x69 &  x70 &  x77 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x0 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x71 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x95;
assign c530 =  x0 &  x1 &  x4 &  x18 &  x29 &  x30 &  x31 &  x38 &  x39 &  x40 &  x47 &  x48 &  x50 &  x57 &  x58 &  x59 &  x60 &  x67 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x89 &  x90 & ~x2 & ~x3 & ~x8 & ~x25 & ~x32 & ~x45 & ~x63 & ~x65 & ~x72 & ~x73 & ~x83 & ~x85 & ~x92 & ~x93;
assign c532 =  x1 &  x3 &  x16 &  x17 &  x19 &  x20 &  x26 &  x27 &  x28 &  x30 &  x31 &  x38 &  x39 &  x46 &  x47 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x61 &  x62 &  x68 &  x69 &  x70 &  x77 &  x79 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x22 & ~x23 & ~x24 & ~x25 & ~x54 & ~x65 & ~x75 & ~x82 & ~x83 & ~x84 & ~x92 & ~x93;
assign c536 = ~x77;
assign c538 =  x93;
assign c540 =  x21 &  x26 &  x28 &  x31 &  x38 &  x46 &  x50 &  x51 &  x61 &  x62 &  x71 &  x79 & ~x22 & ~x45;
assign c542 =  x1 &  x4 &  x16 &  x17 &  x18 &  x19 &  x28 &  x29 &  x38 &  x46 &  x47 &  x70 &  x76 &  x87 &  x88 &  x89 & ~x6 & ~x22 & ~x23 & ~x24 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x54 & ~x55 & ~x60 & ~x61 & ~x62 & ~x63 & ~x65 & ~x72 & ~x75 & ~x82 & ~x83 & ~x85 & ~x92 & ~x93 & ~x95;
assign c544 =  x24;
assign c546 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x61 &  x62 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x45 & ~x54 & ~x55 & ~x64 & ~x65 & ~x73 & ~x74 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c548 =  x5 &  x17 &  x18 &  x27 &  x29 &  x37 &  x38 &  x42 &  x46 &  x50 &  x67 &  x70 &  x71 &  x78 &  x80 &  x87 &  x90 &  x91 & ~x4 & ~x22 & ~x24 & ~x25 & ~x35 & ~x45 & ~x55;
assign c552 = ~x27;
assign c554 = ~x78;
assign c556 =  x1 &  x4 &  x13 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x38 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x89 &  x90 & ~x2 & ~x6 & ~x7 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c558 =  x0 &  x4 & ~x50;
assign c560 =  x1 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x41 & ~x42 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94;
assign c562 =  x0 &  x1 &  x4 &  x16 &  x17 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x37 &  x39 &  x46 &  x47 &  x48 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x79 &  x87 &  x89 & ~x2 & ~x5 & ~x24 & ~x25 & ~x32 & ~x33 & ~x35 & ~x43 & ~x54 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x84 & ~x92 & ~x94 & ~x95;
assign c564 =  x8 &  x18 &  x58 & ~x45 & ~x60;
assign c566 =  x0 &  x1 &  x10 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c568 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x61 &  x62 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x44 & ~x45 & ~x54 & ~x55 & ~x64 & ~x65 & ~x72 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c570 =  x0 &  x1 &  x4 &  x16 &  x18 &  x19 &  x28 &  x29 &  x30 &  x37 &  x38 &  x39 &  x46 &  x48 &  x49 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x76 &  x78 &  x86 &  x87 &  x88 &  x90 & ~x3 & ~x6 & ~x22 & ~x24 & ~x25 & ~x32 & ~x35 & ~x43 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x65 & ~x73 & ~x74 & ~x82 & ~x83 & ~x84 & ~x93;
assign c572 =  x0 &  x1 &  x16 &  x19 &  x20 &  x26 &  x27 &  x28 &  x30 &  x36 &  x37 &  x48 &  x56 &  x57 &  x66 &  x68 &  x69 &  x79 &  x80 &  x89 &  x90 & ~x2 & ~x25 & ~x33 & ~x34 & ~x42 & ~x43 & ~x51 & ~x53 & ~x54 & ~x61 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x93 & ~x95;
assign c574 =  x85;
assign c576 =  x1 &  x16 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x31 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x51 &  x56 &  x57 &  x58 &  x59 &  x61 &  x62 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x79 &  x80 &  x86 &  x87 &  x88 &  x90 &  x91 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x55 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x93;
assign c578 =  x1 &  x16 &  x17 &  x18 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x37 &  x38 &  x46 &  x47 &  x49 &  x56 &  x58 &  x59 &  x60 &  x66 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x6 & ~x9 & ~x22 & ~x23 & ~x24 & ~x33 & ~x34 & ~x35 & ~x44 & ~x52 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c580 = ~x39;
assign c582 =  x0 &  x1 &  x4 &  x17 &  x18 &  x19 &  x37 &  x39 &  x48 &  x56 &  x57 &  x67 &  x80 &  x88 &  x90 & ~x3 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x45 & ~x54 & ~x82 & ~x84 & ~x93;
assign c584 = ~x59;
assign c586 =  x1 &  x4 &  x5 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x6 & ~x7 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c588 =  x1 &  x5 &  x16 &  x17 &  x18 &  x19 &  x20 &  x27 &  x28 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x57 &  x58 &  x60 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x45 & ~x51 & ~x52 & ~x53 & ~x55 & ~x62 & ~x63 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x92 & ~x93 & ~x94 & ~x95;
assign c590 =  x94;
assign c592 =  x84;
assign c594 =  x0 &  x1 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c596 =  x1 &  x3 &  x4 &  x16 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c598 = ~x59;
assign c5100 =  x0 &  x4 & ~x50;
assign c5102 = ~x89;
assign c5104 =  x1 &  x3 &  x6 &  x16 &  x17 &  x19 &  x20 &  x26 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x46 &  x47 &  x49 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x78 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x0 & ~x2 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5106 =  x43;
assign c5108 =  x55;
assign c5110 =  x1 &  x8 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x61 &  x62 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x45 & ~x54 & ~x55 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5112 =  x4 &  x17 &  x20 &  x30 &  x37 &  x40 &  x52 &  x56 &  x77 & ~x2 & ~x7 & ~x23 & ~x45 & ~x72 & ~x83 & ~x94;
assign c5114 =  x0 &  x1 &  x4 &  x16 &  x19 &  x20 &  x27 &  x28 &  x30 &  x37 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x66 &  x67 &  x69 &  x70 &  x76 &  x77 &  x79 &  x80 &  x86 &  x88 &  x89 & ~x2 & ~x3 & ~x6 & ~x23 & ~x24 & ~x25 & ~x35 & ~x44 & ~x52 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x72 & ~x73 & ~x85 & ~x93 & ~x95;
assign c5116 =  x43;
assign c5118 =  x85;
assign c5120 =  x0 &  x1 &  x4 &  x16 &  x18 &  x20 &  x26 &  x27 &  x28 &  x29 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x78 &  x79 &  x80 &  x86 &  x87 &  x89 &  x90 & ~x2 & ~x3 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x44 & ~x54 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94;
assign c5122 = ~x77;
assign c5124 =  x1 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x61 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5126 =  x35;
assign c5128 =  x0 &  x1 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5130 =  x0 &  x1 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x3 & ~x6 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5132 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x52 &  x56 &  x57 &  x58 &  x59 &  x60 &  x61 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x54 & ~x55 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5134 =  x1 &  x3 &  x5 &  x6 &  x9 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5138 =  x1 &  x3 &  x8 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x61 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5140 =  x1 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x38 &  x39 &  x40 &  x42 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x80 &  x86 &  x88 &  x90 & ~x2 & ~x7 & ~x22 & ~x23 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x54 & ~x55 & ~x65 & ~x74 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x95;
assign c5142 =  x1 &  x3 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5144 =  x0 &  x1 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x38 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x22 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x51 & ~x52 & ~x53 & ~x54 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5146 =  x3 &  x4 &  x16 &  x17 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x36 &  x37 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x67 &  x68 &  x70 &  x76 &  x77 &  x78 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5148 =  x1 &  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x0 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x61 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5150 =  x3 &  x63;
assign c5152 =  x1 &  x16 &  x20 &  x26 &  x27 &  x28 &  x30 &  x31 &  x36 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x58 &  x59 &  x60 &  x62 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x63 & ~x65 & ~x72 & ~x73 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x95;
assign c5154 =  x30 &  x62 &  x70 &  x71 &  x79 &  x81 &  x86 & ~x2 & ~x22 & ~x65 & ~x73 & ~x82;
assign c5156 =  x43;
assign c5158 =  x1 &  x4 &  x16 &  x26 &  x29 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x58 &  x59 &  x66 &  x67 &  x69 &  x70 &  x77 &  x80 &  x89 &  x90 & ~x2 & ~x3 & ~x23 & ~x24 & ~x34 & ~x35 & ~x43 & ~x52 & ~x53 & ~x55 & ~x63 & ~x65 & ~x72 & ~x75 & ~x84 & ~x85 & ~x93;
assign c5160 =  x74;
assign c5162 = ~x18;
assign c5164 =  x0 &  x4 & ~x3 & ~x6;
assign c5166 =  x75;
assign c5168 =  x0 &  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x63 & ~x65 & ~x71 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5170 = ~x59;
assign c5172 =  x0 &  x4 &  x18 &  x19 &  x20 &  x26 &  x28 &  x46 &  x48 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x69 &  x70 &  x76 &  x77 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 & ~x2 & ~x3 & ~x5 & ~x22 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x44 & ~x55 & ~x64 & ~x65 & ~x72 & ~x73 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x93 & ~x95;
assign c5174 =  x35;
assign c5176 =  x1 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x52 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x54 & ~x64 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5178 = ~x57;
assign c5180 =  x35;
assign c5182 =  x1 &  x4 &  x5 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x6 & ~x14 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5186 =  x35;
assign c5188 =  x1 &  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x2 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x51 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5190 =  x43;
assign c5192 =  x1 &  x4 &  x26 &  x47 &  x52 &  x60 &  x76 &  x78 & ~x7 & ~x32 & ~x54 & ~x74 & ~x81 & ~x84;
assign c5194 =  x39 &  x40 & ~x60;
assign c5196 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x42 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x7 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5198 =  x1 &  x3 &  x14 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x79 &  x80 &  x86 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5200 =  x1 &  x8 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x56 &  x57 &  x66 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x91 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x54 & ~x55 & ~x60 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5202 =  x0 &  x1 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5204 =  x1 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x6 & ~x13 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x94 & ~x95;
assign c5206 =  x95;
assign c5208 =  x55;
assign c5210 =  x55;
assign c5212 =  x1 &  x3 &  x16 &  x17 &  x18 &  x20 &  x21 &  x27 &  x28 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x42 &  x46 &  x48 &  x50 &  x56 &  x57 &  x58 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x80 &  x87 &  x88 &  x90 & ~x0 & ~x2 & ~x22 & ~x24 & ~x34 & ~x44 & ~x45 & ~x54 & ~x55 & ~x65 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x92 & ~x93;
assign c5214 = ~x46;
assign c5216 = ~x69;
assign c5218 = ~x77;
assign c5220 =  x1 &  x3 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x54 & ~x55 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5222 =  x34;
assign c5224 =  x1 &  x5 &  x6 &  x8 &  x9 &  x17 &  x18 &  x19 &  x20 &  x21 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x59 &  x66 &  x68 &  x70 &  x79 &  x80 &  x89 &  x90 &  x91 & ~x2 & ~x4 & ~x22 & ~x23 & ~x25 & ~x33 & ~x34 & ~x35 & ~x44 & ~x53 & ~x55 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x92 & ~x93 & ~x94;
assign c5226 = ~x26;
assign c5228 =  x18 &  x19 &  x21 &  x29 &  x38 &  x40 &  x41 &  x42 &  x46 &  x47 &  x56 &  x71 &  x80 &  x89 & ~x4 & ~x25 & ~x45 & ~x65 & ~x73 & ~x74 & ~x82 & ~x92 & ~x93 & ~x94;
assign c5230 =  x43;
assign c5232 =  x55;
assign c5234 =  x83 &  x95;
assign c5236 =  x1 &  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x29 &  x30 &  x36 &  x37 &  x38 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x68 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x87 &  x88 &  x90 &  x91 & ~x0 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x44 & ~x51 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5238 = ~x39;
assign c5240 =  x1 &  x3 &  x5 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x0 & ~x2 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x61 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5242 =  x55;
assign c5244 =  x33;
assign c5246 = ~x27;
assign c5248 =  x33;
assign c5250 =  x1 &  x3 &  x5 &  x6 &  x9 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5252 = ~x76;
assign c5254 =  x0 &  x1 &  x4 &  x16 &  x17 &  x26 &  x27 &  x29 &  x31 &  x36 &  x38 &  x40 &  x41 &  x46 &  x47 &  x49 &  x56 &  x59 &  x60 &  x68 &  x70 &  x78 &  x80 &  x86 &  x87 &  x88 &  x90 & ~x3 & ~x22 & ~x24 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x53 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x74 & ~x75 & ~x82 & ~x83 & ~x85 & ~x92 & ~x93 & ~x95;
assign c5256 =  x0 &  x1 &  x4 &  x17 &  x18 &  x20 &  x26 &  x27 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x47 &  x48 &  x56 &  x57 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5258 =  x34;
assign c5260 =  x16 &  x20 &  x27 &  x36 &  x37 &  x48 &  x49 &  x50 &  x56 &  x59 &  x61 &  x62 &  x66 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x90 & ~x9 & ~x23 & ~x34 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x64 & ~x75 & ~x82 & ~x83 & ~x92 & ~x94 & ~x95;
assign c5262 =  x1 &  x4 &  x16 &  x17 &  x26 &  x28 &  x36 &  x48 &  x49 &  x58 &  x59 &  x70 &  x76 &  x86 &  x87 & ~x2 & ~x5 & ~x15 & ~x24 & ~x33 & ~x35 & ~x44 & ~x45 & ~x54 & ~x65 & ~x74 & ~x75 & ~x84 & ~x92 & ~x94;
assign c5264 =  x43;
assign c5266 =  x1 &  x3 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x36 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x5 & ~x22 & ~x24 & ~x25 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x55 & ~x65 & ~x73 & ~x74 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5268 =  x1 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5270 = ~x48;
assign c5272 =  x55;
assign c5274 =  x1 &  x3 &  x4 &  x16 &  x17 &  x19 &  x27 &  x28 &  x29 &  x30 &  x37 &  x38 &  x46 &  x48 &  x59 &  x66 &  x67 &  x68 &  x69 &  x77 &  x80 &  x86 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x35 & ~x42 & ~x43 & ~x44 & ~x53 & ~x54 & ~x55 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x85 & ~x92 & ~x93 & ~x95;
assign c5276 = ~x38;
assign c5278 =  x55;
assign c5280 =  x0 &  x1 &  x4 &  x16 &  x20 &  x26 &  x27 &  x28 &  x30 &  x38 &  x46 &  x47 &  x56 &  x66 &  x67 &  x69 &  x70 &  x76 &  x77 &  x78 &  x80 & ~x3 & ~x5 & ~x22 & ~x23 & ~x25 & ~x34 & ~x44 & ~x53 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x92 & ~x94 & ~x95;
assign c5282 =  x1 &  x18 &  x28 &  x31 &  x46 &  x50 &  x62 &  x77 &  x78 &  x80 & ~x45 & ~x55 & ~x65 & ~x73 & ~x74 & ~x82;
assign c5284 =  x1 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x61 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5286 =  x1 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x61 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5290 =  x55;
assign c5292 =  x0 &  x1 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x3 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5294 =  x1 &  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x21 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x0 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5296 =  x1 &  x16 &  x17 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x49 &  x50 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x69 &  x70 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x60 & ~x61 & ~x63 & ~x64 & ~x65 & ~x72 & ~x74 & ~x75 & ~x82 & ~x83 & ~x85 & ~x92 & ~x93 & ~x94;
assign c5298 =  x1 &  x3 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x36 &  x38 &  x47 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x90 & ~x0 & ~x2 & ~x5 & ~x23 & ~x24 & ~x25 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x64 & ~x65 & ~x74 & ~x75 & ~x82 & ~x84 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5300 =  x8 & ~x59;
assign c5302 =  x4 &  x16 &  x19 &  x20 &  x26 &  x27 &  x28 &  x30 &  x36 &  x37 &  x46 &  x47 &  x48 &  x49 &  x66 &  x69 &  x70 &  x76 &  x78 &  x80 &  x87 & ~x6 & ~x7 & ~x35 & ~x43 & ~x45 & ~x72 & ~x74 & ~x75 & ~x82 & ~x84 & ~x92;
assign c5304 =  x1 &  x7 &  x16 &  x17 &  x18 &  x20 &  x26 &  x27 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x56 &  x57 &  x66 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x89 &  x90 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x41 & ~x42 & ~x43 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x65 & ~x71 & ~x72 & ~x73 & ~x74 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94;
assign c5306 = ~x38;
assign c5308 =  x1 &  x4 &  x13 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x36 &  x37 &  x38 &  x47 &  x48 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x70 &  x76 &  x77 &  x78 &  x80 &  x89 & ~x2 & ~x5 & ~x23 & ~x25 & ~x34 & ~x35 & ~x45 & ~x53 & ~x55 & ~x63 & ~x73 & ~x74 & ~x82 & ~x83 & ~x84 & ~x92 & ~x95;
assign c5310 =  x83;
assign c5312 =  x1 &  x3 &  x4 &  x18 &  x20 &  x26 &  x30 &  x38 &  x46 &  x48 &  x49 &  x50 &  x58 &  x67 &  x68 &  x69 &  x70 &  x77 &  x80 &  x90 & ~x0 & ~x2 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x44 & ~x45 & ~x54 & ~x55 & ~x63 & ~x84 & ~x92 & ~x93 & ~x95;
assign c5314 =  x0 &  x1 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x27 &  x29 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x57 &  x67 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x88 &  x89 &  x91 & ~x6 & ~x22 & ~x24 & ~x25 & ~x34 & ~x35 & ~x64 & ~x65 & ~x73 & ~x82 & ~x83 & ~x84 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5316 =  x1 &  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x8 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5318 = ~x17;
assign c5320 =  x1 &  x3 &  x4 &  x16 &  x17 &  x18 &  x20 &  x26 &  x29 &  x30 &  x36 &  x37 &  x38 &  x47 &  x48 &  x49 &  x56 &  x57 &  x59 &  x66 &  x67 &  x69 &  x76 &  x78 &  x79 &  x80 &  x87 &  x89 &  x90 & ~x2 & ~x5 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x55 & ~x63 & ~x73 & ~x74 & ~x82 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94;
assign c5322 =  x1 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x60 &  x61 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x5 & ~x22 & ~x23 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x72 & ~x74 & ~x75 & ~x82 & ~x83 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5324 =  x35;
assign c5326 =  x43;
assign c5328 =  x35;
assign c5330 = ~x56;
assign c5332 =  x1 &  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x21 &  x26 &  x28 &  x29 &  x31 &  x36 &  x37 &  x38 &  x39 &  x41 &  x46 &  x48 &  x49 &  x50 &  x51 &  x56 &  x58 &  x59 &  x60 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x8 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x81 & ~x83 & ~x85 & ~x92 & ~x93 & ~x94;
assign c5334 =  x0 &  x1 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x3 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5336 =  x0 &  x1 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5338 =  x0 &  x1 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x61 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x54 & ~x55 & ~x63 & ~x64 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5340 =  x1 &  x3 &  x4 &  x16 &  x19 &  x20 &  x26 &  x27 &  x28 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x54 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x95;
assign c5342 =  x4 &  x68 &  x70 & ~x5 & ~x25 & ~x51 & ~x74;
assign c5344 =  x65;
assign c5348 = ~x77;
assign c5350 =  x0 &  x1 &  x4 &  x17 &  x20 &  x29 &  x30 &  x36 &  x40 &  x46 &  x47 &  x48 &  x57 &  x59 &  x69 &  x70 &  x71 &  x86 & ~x3 & ~x8 & ~x22 & ~x25 & ~x33 & ~x44 & ~x65 & ~x73 & ~x93 & ~x94;
assign c5352 =  x63;
assign c5354 =  x1 &  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x0 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x51 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5356 =  x53;
assign c5358 =  x65;
assign c5360 =  x0 &  x1 &  x4 &  x11 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x60 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x3 & ~x22 & ~x23 & ~x24 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5364 = ~x27;
assign c5366 = ~x36;
assign c5368 = ~x56;
assign c5370 = ~x66;
assign c5374 =  x8 &  x16 &  x29 &  x37 &  x38 &  x46 &  x48 &  x67 &  x68 &  x70 &  x88 &  x91 & ~x22 & ~x23 & ~x25 & ~x34 & ~x44 & ~x60 & ~x62 & ~x63 & ~x74 & ~x82 & ~x84 & ~x94;
assign c5376 = ~x27;
assign c5378 =  x62;
assign c5380 =  x1 &  x4 &  x17 &  x18 &  x20 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x66 &  x67 &  x69 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x5 & ~x22 & ~x24 & ~x25 & ~x32 & ~x34 & ~x35 & ~x42 & ~x43 & ~x45 & ~x55 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5382 = ~x27;
assign c5384 =  x1 &  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x58 &  x59 &  x60 &  x66 &  x67 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x11 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5386 =  x1 &  x5 &  x6 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x40 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x61 &  x62 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x54 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5388 =  x43;
assign c5390 = ~x17;
assign c5392 =  x16 &  x17 &  x27 &  x30 &  x36 &  x40 &  x46 &  x48 &  x49 &  x50 &  x58 &  x59 &  x62 &  x69 &  x77 &  x78 &  x79 &  x80 &  x81 &  x86 &  x87 &  x90 & ~x2 & ~x22 & ~x25 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x74 & ~x82 & ~x83;
assign c5394 =  x3 &  x27 &  x28 &  x46 &  x59 &  x69 &  x70 &  x80 &  x86 &  x88 &  x90 & ~x2 & ~x32 & ~x33 & ~x35 & ~x41 & ~x42 & ~x44 & ~x51 & ~x52 & ~x54 & ~x73 & ~x75 & ~x84;
assign c5396 =  x3 &  x17 &  x20 &  x29 &  x30 &  x37 &  x47 &  x49 &  x50 &  x56 &  x57 &  x59 &  x60 &  x66 &  x67 &  x70 &  x78 &  x80 &  x86 &  x88 &  x90 & ~x2 & ~x23 & ~x24 & ~x33 & ~x51 & ~x52 & ~x62 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x94 & ~x95;
assign c5398 =  x1 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x5 & ~x8 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5400 =  x1 &  x3 &  x5 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x42 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5402 =  x1 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x6 & ~x21 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x41 & ~x42 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5404 = ~x78;
assign c5406 = ~x16;
assign c5408 =  x1 &  x3 &  x16 &  x17 &  x18 &  x20 &  x26 &  x27 &  x28 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x42 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x66 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x44 & ~x45 & ~x54 & ~x55 & ~x61 & ~x63 & ~x64 & ~x73 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x94 & ~x95;
assign c5410 = ~x59 & ~x81;
assign c5412 =  x3 &  x16 &  x18 &  x19 &  x20 &  x21 &  x26 &  x27 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x42 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x58 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x89 &  x90 & ~x0 & ~x22 & ~x23 & ~x24 & ~x33 & ~x34 & ~x35 & ~x45 & ~x54 & ~x55 & ~x65 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x95;
assign c5414 =  x1 &  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x0 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x51 & ~x52 & ~x53 & ~x54 & ~x55 & ~x61 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5416 = ~x37;
assign c5418 =  x1 &  x3 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5420 = ~x26;
assign c5422 =  x34;
assign c5424 =  x74;
assign c5426 = ~x17;
assign c5428 =  x1 &  x3 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5430 =  x1 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x21 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5432 = ~x26;
assign c5434 =  x8 &  x20 &  x26 &  x36 &  x38 &  x39 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x70 &  x76 &  x77 &  x78 &  x86 &  x87 &  x90 & ~x10 & ~x21 & ~x23 & ~x24 & ~x25 & ~x33 & ~x35 & ~x64 & ~x65 & ~x72 & ~x74 & ~x84 & ~x85 & ~x92 & ~x93;
assign c5436 =  x1 &  x3 &  x16 &  x17 &  x18 &  x27 &  x28 &  x29 &  x37 &  x38 &  x39 &  x46 &  x48 &  x49 &  x52 &  x56 &  x57 &  x66 &  x68 &  x69 &  x70 &  x77 &  x78 &  x79 &  x80 &  x86 &  x88 &  x89 & ~x0 & ~x2 & ~x22 & ~x24 & ~x25 & ~x34 & ~x35 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x65 & ~x73 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94;
assign c5438 =  x35;
assign c5440 = ~x88;
assign c5442 =  x0 &  x1 &  x4 &  x26 &  x28 &  x29 &  x30 &  x36 &  x38 &  x39 &  x47 &  x48 &  x50 &  x57 &  x58 &  x59 &  x60 &  x68 &  x77 &  x78 &  x80 &  x87 &  x90 & ~x2 & ~x3 & ~x23 & ~x32 & ~x35 & ~x44 & ~x52 & ~x64 & ~x65 & ~x72 & ~x74 & ~x75 & ~x85 & ~x92;
assign c5444 =  x1 &  x3 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5446 =  x0 &  x1 &  x4 &  x16 &  x18 &  x19 &  x20 &  x27 &  x28 &  x30 &  x37 &  x38 &  x46 &  x47 &  x48 &  x56 &  x70 &  x78 &  x79 &  x80 &  x86 &  x87 &  x89 &  x90 & ~x2 & ~x5 & ~x23 & ~x34 & ~x44 & ~x45 & ~x52 & ~x63 & ~x73 & ~x74 & ~x82 & ~x85 & ~x92 & ~x93;
assign c5448 = ~x38;
assign c5452 =  x0 &  x1 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x78 &  x79 &  x80 &  x86 &  x87 &  x90 & ~x2 & ~x3 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x35 & ~x44 & ~x45 & ~x54 & ~x55 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c5454 =  x1 &  x3 &  x4 &  x17 &  x18 &  x20 &  x27 &  x28 &  x29 &  x30 &  x37 &  x39 &  x46 &  x48 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x5 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5456 = ~x28;
assign c5458 =  x55;
assign c5460 =  x33;
assign c5464 =  x55;
assign c5466 =  x1 &  x4 &  x14 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x36 &  x37 &  x38 &  x39 &  x46 &  x57 &  x58 &  x67 &  x68 &  x70 &  x77 &  x78 &  x79 &  x80 &  x88 & ~x2 & ~x23 & ~x24 & ~x32 & ~x33 & ~x34 & ~x35 & ~x45 & ~x53 & ~x62 & ~x64 & ~x72 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x95;
assign c5468 =  x34;
assign c5470 =  x43;
assign c5472 = ~x36;
assign c5474 =  x0 &  x1 &  x8 &  x16 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c5476 =  x0 &  x1 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x48 &  x49 &  x56 &  x57 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x2 & ~x3 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5478 =  x43;
assign c5480 =  x75;
assign c5482 =  x1 &  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x8 & ~x9 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5486 =  x0 &  x1 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x56 &  x57 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x3 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5488 = ~x49;
assign c5490 =  x62;
assign c5494 =  x0 &  x1 &  x4 &  x52 & ~x72;
assign c5496 =  x0 &  x1 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x29 &  x30 &  x36 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x57 &  x66 &  x68 &  x69 &  x70 &  x76 &  x78 &  x79 &  x80 &  x86 &  x87 &  x90 & ~x2 & ~x3 & ~x11 & ~x22 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5498 =  x1 &  x3 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c51 =  x2;
assign c53 =  x1 &  x16 &  x17 &  x19 &  x20 &  x27 &  x28 &  x29 &  x37 &  x38 &  x46 &  x48 &  x49 &  x56 &  x57 &  x66 &  x68 &  x70 &  x77 &  x78 &  x80 &  x86 &  x87 &  x89 & ~x4 & ~x7 & ~x22 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x64 & ~x75 & ~x82 & ~x84 & ~x85 & ~x92 & ~x93 & ~x95;
assign c55 = ~x80;
assign c57 =  x44;
assign c59 = ~x1;
assign c511 =  x2;
assign c513 = ~x58;
assign c515 =  x2;
assign c517 =  x82;
assign c519 =  x0 &  x27 &  x67 & ~x4 & ~x35 & ~x45 & ~x62 & ~x93 & ~x95;
assign c521 = ~x80;
assign c523 = ~x20;
assign c525 = ~x70;
assign c527 = ~x70;
assign c529 = ~x80;
assign c531 = ~x3 & ~x4;
assign c533 =  x82;
assign c535 =  x73;
assign c537 =  x82;
assign c539 = ~x49;
assign c541 = ~x68;
assign c545 =  x93;
assign c547 =  x36 &  x67 & ~x3 & ~x4 & ~x8 & ~x23 & ~x95;
assign c549 = ~x4 & ~x5;
assign c551 =  x1 &  x17 &  x18 &  x20 &  x26 &  x28 &  x30 &  x37 &  x38 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x89 &  x90 & ~x4 & ~x7 & ~x22 & ~x23 & ~x24 & ~x33 & ~x34 & ~x35 & ~x45 & ~x72 & ~x73 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x95;
assign c553 = ~x4 & ~x5;
assign c555 =  x1 &  x4 &  x5 &  x6 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c557 = ~x1;
assign c559 = ~x4 & ~x5;
assign c561 = ~x1;
assign c563 =  x82;
assign c565 = ~x1;
assign c567 =  x18 & ~x4 & ~x6 & ~x22;
assign c569 =  x29 &  x56 & ~x4 & ~x6;
assign c571 =  x54;
assign c573 = ~x1;
assign c575 = ~x90;
assign c577 = ~x4 & ~x6 & ~x55;
assign c579 =  x82;
assign c581 = ~x70;
assign c583 = ~x90;
assign c585 = ~x1;
assign c587 =  x22;
assign c589 =  x16 &  x69 & ~x4 & ~x6 & ~x73;
assign c591 =  x92;
assign c593 =  x16 &  x17 &  x19 &  x20 &  x26 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x66 &  x68 &  x69 &  x70 &  x77 &  x78 &  x79 &  x80 &  x86 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x3 & ~x22 & ~x24 & ~x25 & ~x33 & ~x34 & ~x42 & ~x43 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c595 =  x2;
assign c597 =  x1 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x39 &  x46 &  x47 &  x48 &  x56 &  x57 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x4 & ~x7 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x64 & ~x65 & ~x73 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x94;
assign c599 = ~x70;
assign c5101 = ~x4 & ~x5;
assign c5103 = ~x80;
assign c5105 = ~x4 & ~x5;
assign c5107 =  x1 &  x4 &  x5 &  x6 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5109 =  x27 &  x28 &  x41 &  x48 &  x51 &  x58 &  x59 &  x60 &  x70 &  x76 &  x80 &  x90 & ~x0 & ~x3 & ~x24 & ~x25 & ~x35 & ~x54 & ~x64 & ~x65 & ~x85 & ~x95;
assign c5111 =  x92;
assign c5113 =  x2;
assign c5115 = ~x1;
assign c5117 =  x2;
assign c5119 =  x22;
assign c5121 = ~x80;
assign c5123 =  x2;
assign c5125 = ~x1;
assign c5127 = ~x80;
assign c5129 = ~x1;
assign c5131 = ~x70;
assign c5133 =  x72;
assign c5135 =  x44;
assign c5137 = ~x70;
assign c5139 =  x92;
assign c5141 = ~x1;
assign c5143 = ~x20;
assign c5145 = ~x4 & ~x5;
assign c5147 = ~x1;
assign c5149 =  x1 &  x4 &  x5 &  x6 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5151 = ~x70;
assign c5153 =  x92;
assign c5155 =  x16 &  x18 &  x20 &  x26 &  x28 &  x29 &  x31 &  x36 &  x37 &  x39 &  x46 &  x50 &  x51 &  x56 &  x58 &  x60 &  x66 &  x67 &  x71 &  x77 &  x78 &  x80 &  x87 &  x88 &  x89 & ~x0 & ~x3 & ~x23 & ~x25 & ~x33 & ~x34 & ~x44 & ~x45 & ~x53 & ~x65 & ~x74 & ~x75 & ~x82 & ~x84 & ~x85 & ~x93 & ~x94;
assign c5157 =  x16 &  x19 &  x26 &  x28 &  x30 &  x36 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x60 &  x66 &  x67 &  x68 &  x69 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 & ~x0 & ~x2 & ~x3 & ~x23 & ~x24 & ~x25 & ~x32 & ~x45 & ~x52 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x74 & ~x82 & ~x85 & ~x93;
assign c5159 =  x22;
assign c5161 = ~x4 & ~x5;
assign c5163 =  x22;
assign c5165 =  x45;
assign c5167 = ~x1;
assign c5169 = ~x20;
assign c5171 = ~x90;
assign c5173 =  x82;
assign c5175 = ~x78;
assign c5177 =  x2;
assign c5179 =  x44;
assign c5181 = ~x4 & ~x6;
assign c5183 =  x69 & ~x4 & ~x6 & ~x83;
assign c5185 =  x1 &  x4 &  x5 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5187 =  x73;
assign c5189 =  x16 &  x17 &  x18 &  x27 &  x37 &  x48 &  x56 &  x66 &  x67 &  x68 &  x69 &  x77 &  x79 &  x87 &  x88 &  x89 & ~x4 & ~x7 & ~x22 & ~x23 & ~x24 & ~x33 & ~x34 & ~x54 & ~x55 & ~x64 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5193 = ~x20;
assign c5195 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x3 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5197 =  x73;
assign c5199 = ~x4 & ~x5;
assign c5201 = ~x4 & ~x5;
assign c5205 = ~x3 & ~x4 & ~x8;
assign c5207 = ~x20;
assign c5209 =  x2;
assign c5211 = ~x20;
assign c5213 =  x92;
assign c5215 =  x72;
assign c5217 = ~x1;
assign c5221 =  x24;
assign c5223 =  x1 &  x4 &  x16 &  x17 &  x19 &  x26 &  x30 &  x37 &  x38 &  x39 &  x47 &  x49 &  x50 &  x58 &  x59 &  x60 &  x69 &  x76 &  x78 &  x79 &  x86 &  x87 &  x88 & ~x0 & ~x3 & ~x22 & ~x23 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x44 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94;
assign c5225 =  x2;
assign c5227 =  x1 &  x16 &  x17 &  x18 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x68 &  x69 &  x76 &  x77 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x0 & ~x2 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x95;
assign c5229 =  x2;
assign c5231 =  x1 &  x16 &  x17 &  x18 &  x20 &  x26 &  x27 &  x29 &  x30 &  x36 &  x37 &  x38 &  x46 &  x47 &  x48 &  x56 &  x57 &  x66 &  x67 &  x68 &  x70 &  x76 &  x77 &  x78 &  x80 &  x90 & ~x2 & ~x4 & ~x7 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x55 & ~x72 & ~x73 & ~x74 & ~x82 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5233 =  x82;
assign c5235 =  x1 &  x16 &  x17 &  x18 &  x19 &  x28 &  x29 &  x30 &  x36 &  x38 &  x39 &  x46 &  x47 &  x56 &  x57 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x79 &  x80 &  x86 &  x87 & ~x2 & ~x4 & ~x7 & ~x23 & ~x25 & ~x33 & ~x35 & ~x55 & ~x65 & ~x74 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c5237 =  x73;
assign c5239 =  x92;
assign c5241 =  x22;
assign c5243 =  x2;
assign c5245 =  x0 &  x71 &  x86 & ~x4 & ~x62 & ~x73;
assign c5247 = ~x70;
assign c5249 = ~x4 & ~x5;
assign c5251 =  x2;
assign c5253 =  x23;
assign c5255 = ~x1;
assign c5257 =  x2;
assign c5259 = ~x70;
assign c5261 = ~x90;
assign c5263 = ~x3 & ~x4 & ~x8;
assign c5265 = ~x1;
assign c5267 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x30 &  x37 &  x38 &  x39 &  x46 &  x47 &  x49 &  x50 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x0 & ~x2 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x62 & ~x63 & ~x64 & ~x73 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5269 =  x92;
assign c5273 =  x2;
assign c5275 = ~x20;
assign c5277 = ~x80;
assign c5279 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x47 &  x56 &  x57 &  x66 &  x68 &  x69 &  x76 &  x78 &  x79 &  x86 &  x87 &  x89 &  x90 & ~x2 & ~x4 & ~x7 & ~x22 & ~x23 & ~x24 & ~x33 & ~x34 & ~x35 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x94 & ~x95;
assign c5281 =  x82;
assign c5283 =  x72;
assign c5285 =  x7 &  x19 &  x29 &  x49 & ~x0 & ~x2 & ~x3 & ~x23 & ~x25 & ~x55 & ~x65 & ~x83 & ~x92;
assign c5287 =  x2;
assign c5289 =  x93;
assign c5291 =  x92;
assign c5293 =  x0 &  x1 &  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x2 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c5295 =  x2;
assign c5297 = ~x80;
assign c5299 = ~x69;
assign c5301 = ~x70;
assign c5303 =  x2;
assign c5305 = ~x1;
assign c5307 = ~x70;
assign c5309 = ~x70;
assign c5311 = ~x20;
assign c5313 = ~x4 & ~x5;
assign c5315 =  x0 & ~x4 & ~x8;
assign c5317 = ~x4 & ~x6 & ~x25;
assign c5319 =  x1 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x39 &  x40 &  x46 &  x47 &  x48 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5321 = ~x4 & ~x31;
assign c5323 =  x2;
assign c5327 = ~x20;
assign c5329 =  x1 &  x16 &  x17 &  x18 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5331 = ~x90;
assign c5333 = ~x80;
assign c5335 = ~x20;
assign c5337 = ~x20;
assign c5339 = ~x1;
assign c5341 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x3 & ~x22 & ~x23 & ~x24 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x62 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x94 & ~x95;
assign c5343 = ~x4 & ~x5;
assign c5345 =  x0 &  x51 &  x60 &  x87 & ~x4 & ~x32 & ~x43 & ~x74;
assign c5347 = ~x70;
assign c5351 =  x26 & ~x4 & ~x6 & ~x85;
assign c5353 =  x18 & ~x3 & ~x4 & ~x8 & ~x84;
assign c5355 =  x1 &  x16 &  x18 &  x19 &  x20 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x66 &  x68 &  x69 &  x76 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x4 & ~x7 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x45 & ~x64 & ~x65 & ~x73 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x94;
assign c5357 = ~x1;
assign c5359 =  x73;
assign c5363 = ~x70;
assign c5365 =  x1 &  x16 &  x17 &  x20 &  x26 &  x27 &  x29 &  x30 &  x31 &  x36 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x80 &  x87 &  x89 & ~x0 & ~x2 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x82 & ~x83 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5367 =  x16 &  x19 &  x20 &  x21 &  x26 &  x27 &  x28 &  x29 &  x36 &  x37 &  x38 &  x40 &  x41 &  x46 &  x47 &  x50 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x70 &  x71 &  x76 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x22 & ~x23 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x95;
assign c5369 = ~x57;
assign c5371 =  x54;
assign c5373 =  x1 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x49 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x80 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x55 & ~x62 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94;
assign c5375 =  x2;
assign c5377 =  x2;
assign c5379 = ~x37;
assign c5381 =  x1 &  x16 &  x20 &  x30 &  x36 &  x37 &  x47 &  x48 &  x50 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x76 &  x77 &  x80 &  x87 &  x89 &  x90 & ~x0 & ~x3 & ~x22 & ~x24 & ~x25 & ~x33 & ~x34 & ~x43 & ~x44 & ~x55 & ~x65 & ~x73 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5383 = ~x80;
assign c5385 = ~x4 & ~x21 & ~x91;
assign c5387 =  x1 &  x4 &  x5 &  x6 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5389 =  x2;
assign c5391 =  x2;
assign c5393 = ~x1;
assign c5395 = ~x80;
assign c5397 =  x2;
assign c5399 = ~x1;
assign c5401 =  x1 &  x17 &  x19 &  x69 &  x88 &  x90 & ~x4 & ~x6 & ~x33 & ~x84 & ~x95;
assign c5403 = ~x1;
assign c5405 =  x22;
assign c5407 =  x72;
assign c5409 =  x2;
assign c5411 =  x92;
assign c5413 =  x53 & ~x4;
assign c5415 = ~x70;
assign c5417 =  x0 & ~x4 & ~x55 & ~x62 & ~x65 & ~x94;
assign c5421 =  x28 & ~x4 & ~x6 & ~x83;
assign c5423 = ~x90;
assign c5425 =  x6 &  x16 &  x17 &  x18 &  x19 &  x21 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5427 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x27 &  x28 &  x29 &  x30 &  x40 &  x46 &  x48 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x79 &  x80 &  x88 &  x89 &  x90 &  x91 & ~x0 & ~x2 & ~x3 & ~x22 & ~x24 & ~x25 & ~x34 & ~x35 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c5429 =  x16 &  x17 &  x20 &  x27 &  x29 &  x30 &  x36 &  x37 &  x40 &  x50 &  x56 &  x57 &  x58 &  x60 &  x67 &  x68 &  x70 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x0 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x45 & ~x64 & ~x65 & ~x72 & ~x73 & ~x82 & ~x83 & ~x95;
assign c5431 = ~x1;
assign c5433 = ~x1;
assign c5435 = ~x1;
assign c5437 =  x73;
assign c5439 = ~x30;
assign c5441 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5443 =  x16 &  x46 &  x70 &  x79 & ~x2 & ~x4 & ~x6 & ~x33 & ~x34 & ~x35 & ~x93 & ~x95;
assign c5445 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x48 &  x49 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x3 & ~x22 & ~x23 & ~x24 & ~x34 & ~x35 & ~x43 & ~x45 & ~x52 & ~x53 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5447 =  x73;
assign c5449 = ~x70;
assign c5451 = ~x20;
assign c5453 = ~x80;
assign c5455 =  x1 &  x4 &  x5 &  x6 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5457 =  x2;
assign c5459 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x27 &  x28 &  x30 &  x36 &  x37 &  x40 &  x46 &  x47 &  x50 &  x56 &  x58 &  x66 &  x67 &  x69 &  x71 &  x76 &  x78 &  x79 &  x80 &  x87 &  x88 & ~x0 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x34 & ~x44 & ~x45 & ~x54 & ~x55 & ~x63 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x95;
assign c5461 =  x72;
assign c5465 = ~x70;
assign c5467 = ~x1;
assign c5469 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x2 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c5471 =  x29 &  x37 &  x79 & ~x4;
assign c5473 =  x83;
assign c5475 =  x92;
assign c5477 =  x92;
assign c5479 = ~x20;
assign c5481 =  x19 &  x26 &  x69 &  x79 & ~x4 & ~x6 & ~x34 & ~x85;
assign c5485 = ~x1;
assign c5487 =  x76 & ~x2 & ~x3 & ~x4 & ~x8;
assign c5489 =  x2;
assign c5491 = ~x47;
assign c5493 = ~x1;
assign c5495 =  x82;
assign c5497 = ~x88;
assign c5499 = ~x80;
assign c60 =  x1 &  x16 &  x19 &  x26 &  x27 &  x28 &  x30 &  x38 &  x46 &  x48 &  x49 &  x50 &  x56 &  x58 &  x66 &  x68 &  x69 &  x70 &  x76 &  x87 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x52 & ~x54 & ~x55 & ~x62 & ~x64 & ~x65 & ~x74 & ~x75 & ~x84 & ~x90 & ~x91 & ~x92 & ~x93 & ~x94 & ~x95;
assign c62 =  x0 &  x1 &  x3 &  x4 &  x5 &  x16 &  x18 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x50 &  x51 &  x59 &  x66 &  x67 &  x77 &  x78 &  x79 &  x86 &  x88 &  x89 & ~x33 & ~x34 & ~x43 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x94 & ~x95;
assign c64 =  x1 &  x19 &  x27 &  x37 &  x39 &  x40 &  x46 &  x56 &  x57 &  x58 &  x60 &  x66 &  x70 & ~x6 & ~x21 & ~x22 & ~x23 & ~x25 & ~x35 & ~x42 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x65 & ~x83 & ~x85 & ~x91 & ~x94 & ~x95;
assign c66 =  x1 &  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 & ~x4 & ~x5 & ~x6 & ~x8 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c68 =  x10 &  x73 & ~x6;
assign c610 =  x43;
assign c612 =  x0 & ~x20;
assign c614 =  x0 &  x32 &  x51 &  x89 & ~x63;
assign c616 = ~x27;
assign c620 =  x1 &  x2 &  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x4 & ~x5 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x95;
assign c622 =  x0 &  x1 &  x3 &  x4 &  x5 &  x18 &  x26 &  x27 &  x29 &  x36 &  x37 &  x39 &  x40 &  x47 &  x49 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x77 &  x79 &  x89 & ~x2 & ~x33 & ~x35 & ~x45 & ~x52 & ~x54 & ~x55 & ~x63 & ~x64 & ~x75 & ~x84 & ~x94;
assign c624 =  x1 &  x2 &  x4 &  x16 &  x17 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x39 &  x46 &  x47 &  x50 &  x56 &  x57 &  x58 &  x66 &  x67 &  x76 &  x77 &  x86 &  x87 & ~x0 & ~x3 & ~x23 & ~x33 & ~x35 & ~x42 & ~x43 & ~x53 & ~x55 & ~x62 & ~x64 & ~x65 & ~x71 & ~x72 & ~x75 & ~x82 & ~x83 & ~x85 & ~x93 & ~x94 & ~x95;
assign c626 =  x1 &  x4 &  x5 &  x16 &  x17 &  x18 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x57 &  x58 &  x59 &  x67 &  x76 &  x77 &  x78 &  x79 &  x88 &  x89 &  x90 & ~x23 & ~x24 & ~x25 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x84 & ~x85;
assign c628 =  x1 &  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x4 & ~x5 & ~x7 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c630 =  x2 &  x62 &  x80 & ~x42 & ~x74;
assign c632 =  x9 &  x16 &  x17 &  x28 &  x37 &  x38 &  x40 &  x57 &  x58 &  x59 &  x78 &  x81 &  x86 &  x87 &  x88 &  x89 &  x91 & ~x5 & ~x22 & ~x24 & ~x34 & ~x53 & ~x55 & ~x65 & ~x73 & ~x83 & ~x92 & ~x93 & ~x94 & ~x95;
assign c634 =  x1 &  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 &  x92 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x75;
assign c636 =  x1 &  x2 &  x11 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 & ~x4 & ~x5 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c638 = ~x39;
assign c640 = ~x27;
assign c642 =  x0 &  x39 &  x78 &  x88 & ~x31 & ~x43 & ~x72 & ~x73 & ~x84;
assign c644 =  x1 &  x4 &  x5 &  x6 &  x16 &  x17 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x38 &  x39 &  x40 &  x46 &  x47 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x86 &  x87 &  x88 & ~x23 & ~x25 & ~x32 & ~x33 & ~x34 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x63 & ~x64 & ~x65 & ~x75 & ~x85 & ~x95;
assign c646 =  x1 &  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x81 &  x86 &  x87 &  x88 & ~x4 & ~x5 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x95;
assign c648 =  x2 &  x39 &  x72 &  x78 & ~x3 & ~x9 & ~x32 & ~x52;
assign c650 =  x1 &  x4 &  x5 &  x16 &  x20 &  x26 &  x27 &  x29 &  x37 &  x38 &  x40 &  x41 &  x46 &  x48 &  x49 &  x51 &  x58 &  x60 &  x66 &  x67 &  x70 &  x76 &  x78 &  x79 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x55 & ~x63 & ~x64 & ~x75 & ~x84;
assign c652 =  x1 &  x2 &  x4 &  x16 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x37 &  x38 &  x40 &  x46 &  x56 &  x57 &  x67 &  x68 &  x76 &  x77 &  x86 &  x87 & ~x0 & ~x3 & ~x14 & ~x24 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x53 & ~x54 & ~x64 & ~x84 & ~x93 & ~x94;
assign c654 =  x0 &  x1 &  x10 &  x19 &  x28 &  x29 &  x38 &  x40 &  x41 &  x46 &  x48 &  x49 &  x50 &  x51 &  x56 &  x59 &  x60 &  x66 &  x68 &  x77 &  x86 &  x90 & ~x24 & ~x32 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x55 & ~x63 & ~x65 & ~x73 & ~x75 & ~x84 & ~x85 & ~x94;
assign c656 =  x2 &  x17 &  x19 &  x26 &  x31 &  x46 &  x47 &  x67 & ~x22 & ~x32 & ~x33 & ~x74 & ~x89;
assign c658 = ~x10;
assign c660 =  x1 &  x2 &  x4 &  x5 &  x16 &  x27 &  x36 &  x38 &  x46 &  x49 &  x50 &  x56 &  x57 &  x58 &  x68 &  x76 &  x87 & ~x3 & ~x33 & ~x42 & ~x43 & ~x52 & ~x55 & ~x64 & ~x65;
assign c662 =  x0 &  x1 &  x16 &  x17 &  x18 &  x19 &  x27 &  x30 &  x37 &  x40 &  x46 &  x47 &  x49 &  x50 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x78 &  x86 &  x87 & ~x5 & ~x23 & ~x24 & ~x25 & ~x34 & ~x43 & ~x45 & ~x52 & ~x55 & ~x62 & ~x64 & ~x75 & ~x83 & ~x85 & ~x94 & ~x95;
assign c666 = ~x77;
assign c668 =  x0 &  x30 & ~x10 & ~x69;
assign c670 =  x2 &  x4 &  x5 &  x19 &  x26 &  x27 &  x28 &  x29 &  x37 &  x39 &  x50 &  x57 &  x59 &  x67 &  x76 &  x86 &  x87 & ~x0 & ~x3 & ~x24 & ~x33 & ~x44 & ~x54 & ~x64 & ~x65 & ~x84 & ~x95;
assign c672 = ~x66;
assign c674 = ~x48;
assign c678 =  x1 &  x4 &  x5 &  x16 &  x17 &  x18 &  x19 &  x21 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x84 & ~x85 & ~x94 & ~x95;
assign c680 =  x1 &  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 & ~x4 & ~x5 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c682 = ~x59;
assign c684 =  x22 &  x41;
assign c686 = ~x77;
assign c688 =  x0 &  x3 &  x4 &  x5 &  x7 &  x17 &  x28 &  x30 &  x37 &  x39 &  x40 &  x47 &  x48 &  x49 &  x58 &  x86 &  x87 &  x88 & ~x34 & ~x43 & ~x44 & ~x53 & ~x74 & ~x75 & ~x95;
assign c690 =  x41 &  x62 & ~x74;
assign c692 = ~x26;
assign c694 =  x0 &  x1 &  x2 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x86 &  x87 &  x88 & ~x4 & ~x5 & ~x7 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x63 & ~x64 & ~x65 & ~x75 & ~x83 & ~x84 & ~x85 & ~x94 & ~x95;
assign c696 =  x0 &  x1 &  x2 &  x16 &  x17 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x38 &  x39 &  x40 &  x48 &  x49 &  x51 &  x57 &  x59 &  x86 & ~x7 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x45 & ~x52 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x84 & ~x94 & ~x95;
assign c698 =  x0 &  x9 &  x10 &  x26 &  x27 &  x28 &  x38 &  x49 &  x50 &  x58 &  x60 &  x71 &  x76 &  x78 &  x79 &  x88 &  x89 & ~x33 & ~x42 & ~x63;
assign c6100 =  x1 &  x2 &  x4 &  x5 &  x17 &  x18 &  x19 &  x27 &  x28 &  x30 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x56 &  x67 &  x86 &  x87 & ~x3 & ~x25 & ~x33 & ~x35 & ~x43 & ~x45 & ~x53 & ~x54 & ~x63 & ~x65 & ~x75 & ~x84 & ~x85 & ~x94;
assign c6102 =  x0 &  x16 &  x82 & ~x74;
assign c6104 =  x2 &  x31 & ~x89 & ~x90;
assign c6106 = ~x89;
assign c6110 =  x1 &  x4 &  x6 &  x17 &  x18 &  x20 &  x26 &  x28 &  x29 &  x30 &  x36 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x77 &  x78 &  x79 &  x80 &  x81 &  x87 &  x88 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x74 & ~x75 & ~x84 & ~x85;
assign c6114 =  x0 &  x2;
assign c6116 =  x1 &  x2 &  x17 &  x18 &  x19 &  x28 &  x30 &  x37 &  x40 &  x47 &  x48 &  x56 &  x57 &  x67 &  x68 &  x69 &  x70 &  x77 &  x78 &  x86 &  x88 &  x89 &  x92 & ~x3 & ~x23 & ~x25 & ~x34 & ~x35 & ~x43 & ~x52 & ~x62 & ~x63 & ~x64 & ~x75;
assign c6118 =  x1 &  x4 &  x5 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x84 & ~x85;
assign c6120 =  x54;
assign c6122 =  x1 &  x4 &  x5 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x84 & ~x85;
assign c6124 =  x1 &  x2 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 & ~x0 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c6126 =  x1 &  x4 &  x5 &  x6 &  x17 &  x27 &  x28 &  x37 &  x40 &  x46 &  x47 &  x48 &  x50 &  x58 &  x86 &  x88 & ~x22 & ~x23 & ~x25 & ~x33 & ~x34 & ~x42 & ~x43 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x74 & ~x85;
assign c6128 =  x50 & ~x20 & ~x85;
assign c6130 =  x16 &  x19 &  x29 &  x30 &  x38 &  x48 &  x49 &  x60 &  x66 &  x76 &  x86 & ~x6 & ~x23 & ~x24 & ~x34 & ~x35 & ~x45 & ~x75 & ~x82 & ~x90 & ~x91 & ~x93;
assign c6132 =  x0 &  x39 & ~x45 & ~x63;
assign c6134 =  x0 &  x3 &  x4 &  x5 &  x7 &  x16 &  x27 &  x37 &  x38 &  x47 &  x48 &  x50 &  x51 &  x86 &  x87 & ~x23 & ~x25 & ~x33 & ~x42 & ~x43 & ~x52 & ~x54 & ~x85;
assign c6136 =  x10 &  x73;
assign c6138 =  x61 &  x73;
assign c6140 =  x1 &  x4 &  x5 &  x17 &  x18 &  x20 &  x26 &  x27 &  x28 &  x31 &  x40 &  x47 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x87 &  x88 & ~x8 & ~x24 & ~x32 & ~x34 & ~x35 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x74 & ~x95;
assign c6144 =  x1 &  x2 &  x16 &  x19 &  x29 &  x30 &  x37 &  x39 &  x40 &  x46 &  x48 &  x49 &  x51 &  x59 &  x68 &  x76 &  x78 & ~x4 & ~x5 & ~x6 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x42 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x74 & ~x75 & ~x81 & ~x84 & ~x93 & ~x94 & ~x95;
assign c6146 =  x31 & ~x89;
assign c6148 =  x0 &  x22;
assign c6150 =  x1 &  x12 &  x17 &  x19 &  x26 &  x29 &  x36 &  x40 &  x49 &  x50 &  x57 &  x58 &  x60 &  x66 &  x67 &  x68 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 & ~x7 & ~x25 & ~x32 & ~x35 & ~x42 & ~x45 & ~x53 & ~x63 & ~x65 & ~x73 & ~x74 & ~x84 & ~x85 & ~x92 & ~x93;
assign c6152 =  x1 &  x4 &  x10 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x30 &  x36 &  x39 &  x48 &  x50 &  x56 &  x57 &  x58 &  x59 &  x69 &  x86 &  x87 & ~x24 & ~x32 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x55 & ~x62 & ~x64 & ~x65 & ~x75 & ~x84 & ~x85 & ~x91 & ~x92;
assign c6154 =  x2 &  x16 &  x18 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x39 &  x40 &  x46 &  x47 &  x48 &  x57 &  x58 &  x59 &  x66 &  x69 &  x70 &  x72 &  x76 &  x79 &  x87 &  x89 & ~x22 & ~x32 & ~x33 & ~x34 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x64 & ~x75 & ~x83 & ~x94;
assign c6156 =  x1 &  x10 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x36 &  x39 &  x40 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x86 &  x87 & ~x34 & ~x35 & ~x42 & ~x44 & ~x55 & ~x62 & ~x65 & ~x75 & ~x80 & ~x81 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c6160 =  x44;
assign c6162 = ~x28;
assign c6164 =  x0 &  x1 &  x3 &  x4 &  x5 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x29 &  x36 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x66 &  x68 &  x69 &  x77 &  x78 &  x88 & ~x2 & ~x42 & ~x43 & ~x45 & ~x54 & ~x62 & ~x63 & ~x75 & ~x85;
assign c6166 =  x2 &  x18 &  x28 &  x36 &  x46 &  x47 &  x57 &  x66 &  x69 &  x79 &  x80 &  x81 &  x82 &  x88 & ~x3 & ~x33 & ~x34 & ~x35 & ~x44 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x65;
assign c6168 =  x0 &  x3 &  x4 &  x16 &  x18 &  x27 &  x29 &  x30 &  x46 &  x47 &  x49 &  x50 &  x57 &  x68 &  x69 &  x77 &  x78 &  x79 &  x87 &  x89 & ~x45 & ~x55 & ~x83 & ~x84 & ~x92;
assign c6170 =  x0 &  x1 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c6172 =  x1 &  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x5 & ~x8 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c6174 =  x55;
assign c6176 =  x1 &  x4 &  x6 &  x10 &  x16 &  x17 &  x18 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x74 & ~x75 & ~x84 & ~x85;
assign c6178 =  x61 &  x72 &  x73 & ~x75;
assign c6180 =  x2 &  x16 &  x17 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x31 &  x36 &  x38 &  x39 &  x46 &  x47 &  x48 &  x49 &  x50 &  x57 &  x58 &  x66 &  x67 &  x68 &  x72 &  x77 &  x78 &  x80 &  x87 &  x89 &  x90 & ~x5 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x65 & ~x75 & ~x83 & ~x84 & ~x85 & ~x95;
assign c6182 =  x2 &  x4 &  x5 &  x16 &  x17 &  x18 &  x20 &  x26 &  x27 &  x31 &  x36 &  x37 &  x39 &  x40 &  x46 &  x49 &  x50 &  x56 &  x58 &  x59 &  x66 &  x69 &  x76 &  x77 &  x86 &  x87 & ~x0 & ~x3 & ~x24 & ~x25 & ~x33 & ~x34 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x64 & ~x65 & ~x75;
assign c6184 =  x0 &  x1 &  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x21 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x3 & ~x4 & ~x5 & ~x23 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75;
assign c6186 = ~x66;
assign c6188 =  x1 &  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 & ~x4 & ~x5 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c6190 =  x19 &  x60 &  x82 & ~x93;
assign c6192 =  x0 &  x1 &  x3 &  x4 &  x5 &  x16 &  x17 &  x18 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x47 &  x48 &  x49 &  x50 &  x56 &  x66 &  x67 &  x76 &  x77 &  x78 &  x79 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x34 & ~x35 & ~x44 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x73 & ~x75 & ~x84 & ~x85 & ~x94;
assign c6194 =  x25 &  x64;
assign c6196 =  x0 &  x1 &  x3 &  x4 &  x5 &  x7 &  x17 &  x18 &  x26 &  x29 &  x36 &  x37 &  x38 &  x39 &  x47 &  x48 &  x49 &  x50 &  x57 &  x66 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x87 & ~x33 & ~x34 & ~x35 & ~x43 & ~x45 & ~x52 & ~x53 & ~x54 & ~x63 & ~x64 & ~x65 & ~x75 & ~x84 & ~x85 & ~x94;
assign c6200 = ~x36;
assign c6202 =  x1 &  x4 &  x5 &  x16 &  x17 &  x26 &  x27 &  x28 &  x29 &  x30 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x57 &  x59 &  x66 &  x68 &  x77 &  x78 &  x79 &  x80 &  x81 &  x88 &  x89 & ~x24 & ~x25 & ~x43 & ~x44 & ~x53 & ~x54 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x84 & ~x85;
assign c6204 =  x25 &  x44;
assign c6206 =  x1 &  x16 &  x17 &  x19 &  x21 &  x26 &  x27 &  x28 &  x29 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x57 &  x58 &  x59 &  x67 &  x70 &  x71 &  x77 &  x78 &  x87 &  x88 &  x90 &  x91 &  x92 & ~x24 & ~x25 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x65 & ~x74 & ~x75;
assign c6208 =  x83;
assign c6210 = ~x27;
assign c6212 =  x1 &  x16 &  x19 &  x27 &  x30 &  x37 &  x48 &  x57 &  x67 &  x69 & ~x22 & ~x23 & ~x24 & ~x42 & ~x43 & ~x44 & ~x55 & ~x62 & ~x65 & ~x72 & ~x80 & ~x81 & ~x84 & ~x93 & ~x94 & ~x95;
assign c6214 = ~x59;
assign c6216 =  x46 &  x58 &  x77 &  x80 &  x81 &  x82 & ~x55 & ~x62;
assign c6218 =  x0 &  x1 &  x2 &  x8 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x39 &  x40 &  x46 &  x47 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 & ~x3 & ~x5 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x55 & ~x64 & ~x65 & ~x75;
assign c6220 =  x1 &  x16 &  x17 &  x18 &  x26 &  x27 &  x28 &  x31 &  x37 &  x48 &  x50 &  x51 &  x57 &  x66 &  x68 &  x69 &  x76 &  x78 &  x86 &  x87 & ~x33 & ~x34 & ~x35 & ~x42 & ~x44 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x72 & ~x73 & ~x74 & ~x75 & ~x80 & ~x83 & ~x85 & ~x93 & ~x95;
assign c6222 =  x1 &  x2 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x76 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x4 & ~x5 & ~x7 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x95;
assign c6224 =  x0 &  x1 &  x2 &  x16 &  x17 &  x19 &  x30 &  x36 &  x38 &  x40 &  x41 &  x47 &  x48 &  x50 &  x51 &  x56 &  x57 &  x67 &  x69 &  x76 &  x86 & ~x3 & ~x5 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x44 & ~x52 & ~x53 & ~x55 & ~x62 & ~x63 & ~x64 & ~x75 & ~x82 & ~x84 & ~x93 & ~x95;
assign c6226 =  x2 & ~x21 & ~x89;
assign c6228 =  x1 &  x4 &  x5 &  x16 &  x17 &  x18 &  x19 &  x28 &  x29 &  x30 &  x31 &  x36 &  x38 &  x40 &  x41 &  x46 &  x48 &  x49 &  x50 &  x51 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x84 & ~x85;
assign c6230 =  x1 &  x4 &  x5 &  x16 &  x17 &  x18 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x70 &  x76 &  x77 &  x78 &  x79 &  x87 &  x88 &  x89 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x53 & ~x54 & ~x55 & ~x63 & ~x73 & ~x74 & ~x75 & ~x84 & ~x85;
assign c6232 = ~x20;
assign c6234 =  x1 &  x2 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x58 &  x59 &  x67 &  x68 &  x69 &  x76 &  x86 &  x87 & ~x3 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x61 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x91 & ~x92 & ~x93 & ~x94 & ~x95;
assign c6236 =  x0 &  x1 &  x3 &  x5 &  x8 & ~x24 & ~x25 & ~x52 & ~x95;
assign c6238 =  x0 &  x1 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x37 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x59 &  x66 &  x67 &  x68 &  x76 &  x77 &  x78 &  x80 &  x81 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x75 & ~x85 & ~x94 & ~x95;
assign c6240 =  x1 &  x16 &  x17 &  x18 &  x19 &  x26 &  x28 &  x29 &  x30 &  x31 &  x36 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x86 &  x87 &  x88 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x80 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94;
assign c6248 =  x1 &  x2 &  x4 &  x5 &  x17 &  x18 &  x27 &  x36 &  x37 &  x39 &  x46 &  x56 &  x58 &  x67 &  x68 &  x77 & ~x0 & ~x3 & ~x23 & ~x24 & ~x25 & ~x45 & ~x75 & ~x85 & ~x95;
assign c6250 =  x5 &  x82;
assign c6252 =  x1 &  x2 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x39 &  x46 &  x47 &  x56 &  x59 &  x67 &  x68 &  x69 &  x76 &  x77 &  x86 & ~x3 & ~x21 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x44 & ~x53 & ~x64 & ~x74 & ~x75 & ~x83 & ~x91 & ~x93 & ~x94;
assign c6256 =  x0 & ~x20;
assign c6260 =  x2 &  x19 &  x46 & ~x34 & ~x74 & ~x89;
assign c6262 =  x54;
assign c6264 =  x1 &  x16 &  x17 &  x19 &  x27 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x51 &  x56 &  x57 &  x58 &  x60 &  x66 &  x68 &  x76 &  x77 &  x78 &  x86 &  x87 &  x89 & ~x4 & ~x5 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x55 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x83 & ~x84 & ~x92 & ~x94 & ~x95;
assign c6266 =  x1 &  x4 &  x5 &  x16 &  x17 &  x18 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x67 &  x76 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x64 & ~x65 & ~x71 & ~x72 & ~x73 & ~x75 & ~x84 & ~x85 & ~x94;
assign c6268 =  x1 &  x4 &  x5 &  x7 &  x16 &  x17 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x59 &  x66 &  x76 &  x87 &  x88 &  x89 & ~x23 & ~x24 & ~x25 & ~x32 & ~x35 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x85 & ~x95;
assign c6270 = ~x69;
assign c6272 =  x16 &  x17 &  x20 &  x31 &  x37 &  x40 &  x46 &  x50 &  x57 &  x68 &  x78 &  x80 & ~x4 & ~x6 & ~x45 & ~x74 & ~x95;
assign c6274 =  x4 &  x5 &  x17 &  x27 &  x29 &  x38 &  x40 &  x48 &  x50 &  x56 &  x57 &  x66 &  x67 &  x68 &  x76 &  x86 & ~x23 & ~x24 & ~x25 & ~x32 & ~x35 & ~x42 & ~x54 & ~x55 & ~x65 & ~x73 & ~x74 & ~x85 & ~x91 & ~x92 & ~x94 & ~x95;
assign c6276 =  x22;
assign c6278 =  x1 &  x17 &  x26 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x76 &  x78 &  x80 &  x81 &  x87 &  x88 & ~x11 & ~x22 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x53 & ~x55 & ~x73 & ~x74 & ~x75 & ~x84 & ~x85 & ~x92 & ~x93 & ~x95;
assign c6280 =  x2 &  x19 &  x21 &  x26 &  x30 &  x31 &  x37 &  x38 &  x39 &  x41 &  x47 &  x49 &  x50 &  x51 &  x59 &  x66 &  x67 &  x76 &  x78 &  x79 &  x81 &  x87 &  x88 &  x89 &  x90 & ~x10 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x54 & ~x55 & ~x62 & ~x63 & ~x65 & ~x75 & ~x85 & ~x94 & ~x95;
assign c6282 = ~x3 & ~x88;
assign c6284 =  x35;
assign c6286 =  x1 &  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x4 & ~x5 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c6288 =  x1 &  x4 &  x5 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x84 & ~x85 & ~x94 & ~x95;
assign c6290 =  x0 &  x1 &  x3 &  x4 &  x5 &  x16 &  x17 &  x18 &  x26 &  x27 &  x28 &  x30 &  x36 &  x37 &  x38 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x76 &  x77 &  x86 &  x87 &  x88 &  x89 & ~x2 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x75 & ~x84 & ~x85 & ~x94 & ~x95;
assign c6292 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x70 &  x71 &  x72 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x75 & ~x84 & ~x85 & ~x94 & ~x95;
assign c6294 = ~x77;
assign c6296 =  x93;
assign c6298 =  x65;
assign c6300 =  x17 &  x19 &  x21 &  x26 &  x27 &  x30 &  x37 &  x38 &  x39 &  x40 &  x47 &  x49 &  x58 &  x59 &  x60 &  x66 &  x68 &  x71 &  x77 &  x78 &  x88 &  x90 &  x91 &  x92 & ~x23 & ~x24 & ~x34 & ~x35 & ~x44 & ~x45 & ~x52 & ~x54 & ~x62 & ~x63 & ~x64 & ~x65;
assign c6302 =  x0 &  x49 &  x56 &  x86 & ~x5 & ~x7 & ~x52 & ~x81;
assign c6304 =  x4 &  x5 &  x31 &  x37 &  x39 &  x40 &  x41 &  x50 &  x56 &  x66 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x24 & ~x33 & ~x34 & ~x35 & ~x53 & ~x75 & ~x83 & ~x85;
assign c6306 =  x1 &  x2 &  x3 &  x17 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x59 &  x60 &  x66 &  x67 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x4 & ~x5 & ~x6 & ~x7 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x34 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x63 & ~x64 & ~x74 & ~x75 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c6308 = ~x87;
assign c6310 =  x0 &  x3 &  x4 &  x5 &  x6 &  x18 &  x26 &  x47 &  x57 &  x66 & ~x34;
assign c6312 =  x55;
assign c6314 =  x2 &  x13 &  x30 &  x48 &  x50 &  x57 &  x69 &  x77 &  x90 & ~x4 & ~x5 & ~x6 & ~x43 & ~x52 & ~x53 & ~x63 & ~x64 & ~x74 & ~x75 & ~x83 & ~x84 & ~x93;
assign c6316 =  x4 &  x5 &  x26 &  x59 &  x67 &  x68 &  x80 &  x88 &  x92 & ~x34 & ~x45 & ~x55;
assign c6318 = ~x77;
assign c6320 = ~x26;
assign c6322 =  x1 &  x4 &  x6 &  x7 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x94 & ~x95;
assign c6324 =  x1 &  x2 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x4 & ~x5 & ~x7 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x94 & ~x95;
assign c6326 =  x85 &  x94;
assign c6328 =  x1 &  x2 &  x4 &  x6 &  x7 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 & ~x0 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x84 & ~x85 & ~x95;
assign c6330 =  x73 & ~x9;
assign c6332 = ~x39;
assign c6334 =  x1 &  x2 &  x3 &  x10 &  x27 &  x30 &  x31 &  x58 &  x66 &  x67 &  x78 &  x86 & ~x4 & ~x5 & ~x6 & ~x25 & ~x42 & ~x44 & ~x45 & ~x53 & ~x55 & ~x64 & ~x75 & ~x83 & ~x84 & ~x85;
assign c6336 =  x4 &  x5 & ~x41;
assign c6338 =  x63;
assign c6340 =  x35;
assign c6342 =  x1 &  x31 &  x40 &  x49 &  x56 &  x58 &  x60 &  x67 &  x70 &  x87 & ~x6 & ~x9 & ~x21 & ~x25 & ~x32 & ~x43 & ~x44 & ~x84 & ~x91;
assign c6344 =  x0 &  x1 &  x3 &  x4 &  x5 &  x16 &  x27 &  x28 &  x29 &  x36 &  x38 &  x39 &  x46 &  x47 &  x49 &  x57 &  x59 &  x60 &  x68 &  x77 &  x78 &  x87 & ~x24 & ~x34 & ~x43 & ~x52 & ~x53 & ~x55 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x85 & ~x95;
assign c6346 =  x1 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x86 &  x87 &  x88 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x64 & ~x65 & ~x75 & ~x80 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c6348 =  x1 &  x2 &  x3 &  x16 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x4 & ~x5 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c6350 =  x1 &  x2 &  x16 &  x17 &  x19 &  x27 &  x28 &  x30 &  x38 &  x40 &  x49 &  x50 &  x56 &  x57 &  x58 &  x60 &  x68 &  x71 &  x76 &  x77 &  x86 &  x89 &  x90 &  x92 & ~x3 & ~x23 & ~x24 & ~x25 & ~x32 & ~x35 & ~x54 & ~x55 & ~x62 & ~x65;
assign c6352 = ~x76;
assign c6354 = ~x66;
assign c6356 = ~x48;
assign c6358 =  x1 &  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x4 & ~x5 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c6360 = ~x46;
assign c6362 =  x22 &  x79;
assign c6364 =  x1 &  x16 &  x17 &  x18 &  x19 &  x27 &  x29 &  x30 &  x38 &  x39 &  x40 &  x50 &  x57 &  x59 &  x68 &  x76 &  x78 &  x79 &  x80 &  x82 &  x86 &  x88 & ~x24 & ~x25 & ~x33 & ~x34 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x84;
assign c6366 =  x1 &  x2 &  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x4 & ~x5 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c6368 =  x0 &  x1 &  x27 &  x37 &  x39 &  x51 &  x66 &  x88 & ~x42 & ~x53 & ~x64 & ~x65 & ~x80 & ~x84 & ~x93 & ~x95;
assign c6370 =  x1 &  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x4 & ~x5 & ~x7 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c6372 = ~x77;
assign c6374 =  x4 &  x5 &  x17 &  x28 &  x30 &  x37 &  x39 &  x48 &  x50 &  x56 &  x57 &  x58 & ~x21 & ~x32 & ~x34 & ~x54 & ~x91 & ~x94;
assign c6376 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x68 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x81 &  x82 &  x86 &  x87 &  x88 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x75;
assign c6378 =  x0 &  x1 &  x17 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x66 &  x76 &  x87 &  x88 & ~x24 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x52 & ~x53 & ~x55 & ~x63 & ~x65 & ~x72 & ~x73 & ~x74 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c6380 =  x1 &  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x76 &  x77 &  x78 &  x79 &  x80 &  x81 &  x86 &  x88 &  x90 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x44 & ~x54 & ~x55 & ~x64 & ~x65 & ~x73 & ~x74 & ~x83 & ~x84 & ~x85 & ~x92 & ~x94 & ~x95;
assign c6382 =  x1 &  x4 &  x5 &  x16 &  x37 &  x48 &  x51 &  x56 & ~x33 & ~x43 & ~x44 & ~x65 & ~x73 & ~x74 & ~x91 & ~x93;
assign c6384 =  x1 &  x2 &  x3 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x4 & ~x5 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c6386 = ~x66;
assign c6388 =  x1 &  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x21 &  x26 &  x27 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x48 &  x51 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x76 &  x77 &  x78 &  x79 &  x80 &  x81 &  x86 &  x87 &  x88 &  x89 &  x90 &  x91 & ~x3 & ~x5 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75;
assign c6390 = ~x60;
assign c6392 =  x1 &  x4 &  x6 &  x7 &  x16 &  x17 &  x18 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x50 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x87 &  x88 & ~x10 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x75 & ~x83 & ~x84 & ~x85 & ~x94;
assign c6394 =  x0 &  x1 &  x16 &  x17 &  x26 &  x27 &  x30 &  x37 &  x41 &  x46 &  x48 &  x50 &  x56 &  x57 &  x67 &  x70 &  x87 &  x88 & ~x33 & ~x42 & ~x43 & ~x44 & ~x45 & ~x55 & ~x62 & ~x65 & ~x72 & ~x74 & ~x75 & ~x84 & ~x85 & ~x94 & ~x95;
assign c6396 =  x1 &  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 & ~x4 & ~x5 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c6398 =  x0 &  x19 &  x30 &  x38 &  x51 &  x59 & ~x33 & ~x53 & ~x55 & ~x80 & ~x85 & ~x94;
assign c6400 =  x1 &  x4 &  x6 &  x16 &  x18 &  x28 &  x36 &  x37 &  x38 &  x48 &  x49 &  x50 &  x57 &  x58 &  x59 &  x60 &  x61 &  x66 &  x67 &  x68 &  x70 &  x76 &  x87 &  x88 &  x89 &  x90 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x62 & ~x63 & ~x64 & ~x75;
assign c6402 =  x65;
assign c6404 =  x1 &  x7 &  x16 &  x19 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x58 &  x59 &  x66 &  x67 &  x69 &  x76 &  x77 &  x78 &  x87 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x75 & ~x80 & ~x81 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94;
assign c6406 =  x1 &  x4 &  x5 &  x16 &  x17 &  x18 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x66 &  x67 &  x76 &  x77 &  x78 &  x86 &  x87 &  x90 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x54 & ~x55 & ~x62 & ~x64 & ~x65 & ~x71 & ~x72 & ~x74 & ~x75 & ~x84 & ~x85 & ~x94 & ~x95;
assign c6408 =  x0 &  x1 &  x3 &  x4 &  x5 &  x17 &  x18 &  x27 &  x29 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x58 &  x67 &  x68 &  x77 &  x78 &  x79 &  x86 &  x89 & ~x23 & ~x24 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x53 & ~x54 & ~x63 & ~x64 & ~x73 & ~x95;
assign c6410 =  x2 &  x4 &  x6 &  x16 &  x17 &  x20 &  x27 &  x29 &  x30 &  x39 &  x48 &  x49 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 & ~x3 & ~x33 & ~x43 & ~x55 & ~x61 & ~x72 & ~x74 & ~x85 & ~x94 & ~x95;
assign c6412 =  x22;
assign c6414 =  x44;
assign c6418 =  x1 &  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x80 &  x81 &  x86 &  x87 &  x88 &  x89 & ~x4 & ~x5 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x94 & ~x95;
assign c6420 =  x1 &  x2 &  x16 &  x17 &  x26 &  x28 &  x38 &  x46 &  x47 &  x48 &  x49 &  x50 &  x58 &  x59 &  x60 &  x68 &  x69 &  x71 &  x72 &  x76 &  x78 & ~x9 & ~x22 & ~x23 & ~x24 & ~x32 & ~x33 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x75;
assign c6422 = ~x76;
assign c6424 =  x1 &  x8 &  x17 &  x19 &  x27 &  x30 &  x40 &  x50 &  x60 &  x67 &  x88 & ~x23 & ~x34 & ~x42 & ~x44 & ~x64 & ~x74 & ~x75 & ~x84 & ~x90 & ~x93;
assign c6428 =  x1 &  x2 &  x7 &  x16 &  x17 &  x18 &  x19 &  x27 &  x29 &  x30 &  x36 &  x37 &  x38 &  x46 &  x47 &  x50 &  x57 &  x58 &  x69 &  x77 &  x78 &  x79 &  x86 &  x87 & ~x0 & ~x23 & ~x24 & ~x25 & ~x33 & ~x42 & ~x43 & ~x52 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x71 & ~x72 & ~x73 & ~x75 & ~x85 & ~x93 & ~x95;
assign c6430 =  x1 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x31 &  x36 &  x38 &  x39 &  x46 &  x50 &  x56 &  x67 &  x76 &  x78 &  x79 &  x86 &  x87 &  x89 &  x91 &  x92 & ~x3 & ~x23 & ~x34 & ~x43 & ~x44 & ~x45 & ~x53 & ~x55 & ~x63 & ~x64 & ~x72;
assign c6432 =  x2 &  x4 &  x5 &  x19 &  x38 &  x50 &  x60 &  x68 &  x87 & ~x3 & ~x23 & ~x32 & ~x35 & ~x44 & ~x45 & ~x63;
assign c6434 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x7 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x91 & ~x92 & ~x93 & ~x94 & ~x95;
assign c6436 =  x1 &  x4 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x39 &  x40 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x59 &  x60 &  x66 &  x68 &  x69 &  x70 &  x87 &  x88 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x52 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x91 & ~x94 & ~x95;
assign c6438 =  x2 &  x16 &  x17 &  x19 &  x20 &  x26 &  x27 &  x29 &  x30 &  x36 &  x38 &  x39 &  x46 &  x48 &  x49 &  x50 &  x51 &  x57 &  x58 &  x66 &  x67 &  x68 &  x76 &  x77 &  x78 &  x86 &  x88 &  x91 & ~x10 & ~x23 & ~x25 & ~x32 & ~x33 & ~x34 & ~x42 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x65 & ~x73 & ~x74 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c6440 =  x4 &  x5 &  x19 &  x29 &  x30 &  x36 &  x39 &  x46 &  x50 &  x58 &  x76 &  x87 &  x89 & ~x23 & ~x25 & ~x32 & ~x42 & ~x61 & ~x64 & ~x73 & ~x74 & ~x75;
assign c6442 = ~x67;
assign c6444 =  x85;
assign c6446 =  x7 & ~x60 & ~x71;
assign c6448 =  x44;
assign c6450 =  x1 &  x2 &  x4 &  x6 &  x16 &  x17 &  x18 &  x19 &  x20 &  x27 &  x28 &  x29 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x0 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x75 & ~x83 & ~x84 & ~x85 & ~x94 & ~x95;
assign c6452 = ~x36;
assign c6454 =  x0 &  x3 &  x4 &  x5 &  x28 &  x39 &  x46 &  x47 &  x49 &  x88 & ~x24 & ~x32 & ~x33 & ~x35 & ~x42 & ~x43 & ~x44 & ~x54 & ~x55 & ~x72 & ~x73 & ~x83 & ~x85;
assign c6456 =  x22;
assign c6458 =  x1 &  x4 &  x5 &  x16 &  x17 &  x26 &  x28 &  x29 &  x30 &  x38 &  x46 &  x47 &  x50 &  x56 &  x57 &  x58 &  x66 &  x67 &  x76 &  x86 & ~x21 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x52 & ~x53 & ~x55 & ~x64 & ~x65 & ~x75 & ~x85 & ~x91 & ~x94 & ~x95;
assign c6460 =  x54;
assign c6462 =  x0 &  x3 &  x4 &  x5 &  x16 &  x17 &  x26 &  x30 &  x37 &  x39 &  x40 &  x46 &  x47 &  x50 &  x56 &  x57 &  x88 & ~x2 & ~x43 & ~x44 & ~x53;
assign c6464 =  x1 &  x4 &  x16 &  x17 &  x18 &  x26 &  x28 &  x29 &  x36 &  x38 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x57 &  x58 &  x59 &  x66 &  x77 &  x78 &  x79 &  x87 &  x88 &  x89 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x71 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c6466 =  x1 &  x2 &  x4 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x3 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c6468 = ~x36;
assign c6470 =  x65;
assign c6472 =  x64;
assign c6474 =  x2 & ~x89;
assign c6476 =  x22 &  x41 &  x79 & ~x83;
assign c6478 = ~x56;
assign c6480 =  x1 &  x4 &  x5 &  x16 &  x17 &  x19 &  x26 &  x27 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x49 &  x56 &  x58 &  x66 &  x67 &  x69 &  x76 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x24 & ~x32 & ~x42 & ~x43 & ~x45 & ~x54 & ~x62 & ~x64 & ~x65 & ~x75 & ~x84 & ~x85 & ~x91 & ~x94;
assign c6482 =  x17 &  x18 &  x28 &  x29 &  x36 &  x37 &  x38 &  x40 &  x46 &  x47 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x77 &  x79 &  x81 &  x86 &  x87 &  x89 &  x90 & ~x5 & ~x7 & ~x22 & ~x25 & ~x33 & ~x34 & ~x42 & ~x43 & ~x44 & ~x52 & ~x55 & ~x63 & ~x73 & ~x75 & ~x85 & ~x94;
assign c6484 =  x1 &  x4 &  x6 &  x16 &  x17 &  x18 &  x19 &  x21 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x69 &  x70 &  x76 &  x77 &  x86 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x85 & ~x93 & ~x94 & ~x95;
assign c6486 =  x56 &  x92 & ~x52 & ~x61;
assign c6488 =  x22 &  x41;
assign c6490 = ~x7 & ~x31;
assign c6492 = ~x59;
assign c6494 =  x65;
assign c6496 =  x16 &  x17 &  x26 &  x28 &  x30 &  x36 &  x37 &  x56 &  x59 &  x60 &  x61 &  x68 &  x69 &  x76 &  x77 &  x80 &  x81 &  x86 &  x87 &  x88 & ~x7 & ~x23 & ~x24 & ~x32 & ~x33 & ~x34 & ~x35 & ~x44 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x75 & ~x85 & ~x95;
assign c6498 =  x0 &  x82;
assign c61 =  x43;
assign c63 =  x1 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x37 &  x38 &  x39 &  x40 &  x41 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c65 = ~x1;
assign c67 =  x95;
assign c69 = ~x2;
assign c611 = ~x1;
assign c613 =  x1 &  x17 &  x18 &  x27 &  x28 &  x30 &  x36 &  x37 &  x38 &  x40 &  x46 &  x47 &  x49 &  x56 &  x57 &  x66 &  x68 &  x69 &  x70 &  x71 &  x76 &  x80 &  x86 &  x88 &  x89 & ~x0 & ~x22 & ~x23 & ~x32 & ~x35 & ~x43 & ~x53 & ~x62 & ~x64 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x92 & ~x93 & ~x94 & ~x95;
assign c615 = ~x50;
assign c617 = ~x1;
assign c619 =  x5 &  x18 &  x19 &  x26 &  x27 &  x28 &  x30 &  x36 &  x37 &  x38 &  x46 &  x56 &  x58 &  x59 &  x66 &  x68 &  x76 &  x77 &  x86 &  x87 & ~x4 & ~x25 & ~x34 & ~x44 & ~x54 & ~x64 & ~x75 & ~x84 & ~x85;
assign c621 =  x54;
assign c623 =  x24;
assign c625 =  x18 &  x19 &  x20 &  x27 &  x29 &  x30 &  x37 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x68 &  x69 &  x70 &  x76 &  x80 &  x86 &  x88 &  x89 &  x90 & ~x2 & ~x22 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x83 & ~x84;
assign c627 = ~x1;
assign c629 = ~x1;
assign c631 =  x17 &  x20 &  x21 &  x28 &  x37 &  x40 &  x46 &  x47 &  x48 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x71 &  x76 &  x77 &  x79 &  x86 &  x87 &  x89 &  x90 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x53 & ~x54 & ~x55 & ~x62 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x85 & ~x92 & ~x93 & ~x95;
assign c633 =  x31 & ~x2 & ~x6 & ~x7;
assign c635 = ~x1;
assign c637 =  x16 &  x17 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x37 &  x49 &  x50 &  x56 &  x57 &  x58 &  x66 &  x67 &  x68 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x2 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x55 & ~x63 & ~x64 & ~x65 & ~x75 & ~x82 & ~x83 & ~x84;
assign c639 =  x1 &  x3 &  x6 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x0 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x94 & ~x95;
assign c641 = ~x2 & ~x3;
assign c643 =  x1 &  x16 &  x19 &  x28 &  x30 &  x31 &  x39 &  x46 &  x47 &  x49 &  x56 &  x58 &  x60 &  x66 &  x70 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x90 &  x91 & ~x23 & ~x24 & ~x25 & ~x32 & ~x34 & ~x35 & ~x42 & ~x45 & ~x52 & ~x54 & ~x61 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x95;
assign c645 = ~x1;
assign c647 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x86 &  x87 &  x88 &  x89 & ~x0 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c649 =  x8 &  x20 &  x29 &  x31 &  x59 &  x60 &  x76 &  x79 &  x90 & ~x3 & ~x22 & ~x23 & ~x24 & ~x44 & ~x45 & ~x55 & ~x73 & ~x85 & ~x92;
assign c651 =  x1 &  x2 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x87 &  x88 &  x89 &  x90 & ~x22 & ~x24 & ~x25 & ~x32 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x85 & ~x92 & ~x93 & ~x95;
assign c653 =  x53;
assign c655 =  x24;
assign c657 = ~x2 & ~x5;
assign c659 = ~x86;
assign c661 =  x1 &  x19 &  x68 &  x69 &  x77 & ~x2 & ~x25 & ~x93;
assign c663 = ~x2 & ~x5;
assign c665 =  x67 & ~x2 & ~x5;
assign c667 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x72 & ~x73 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c669 = ~x58;
assign c671 =  x1 &  x4 &  x16 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x50 &  x56 &  x58 &  x59 &  x76 &  x78 &  x86 &  x87 &  x88 &  x89 & ~x5 & ~x7 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x53 & ~x54 & ~x62 & ~x64 & ~x65 & ~x94 & ~x95;
assign c673 = ~x0 & ~x2;
assign c675 =  x16 &  x19 &  x20 &  x27 &  x28 &  x29 &  x31 &  x40 &  x47 &  x49 &  x50 &  x66 &  x68 &  x69 &  x71 &  x76 &  x78 &  x80 &  x87 &  x89 &  x91 & ~x22 & ~x23 & ~x24 & ~x32 & ~x35 & ~x53 & ~x54 & ~x55 & ~x62 & ~x65 & ~x72 & ~x73 & ~x75 & ~x92 & ~x95;
assign c677 =  x62;
assign c679 =  x1 &  x2 &  x6 &  x7 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x89 & ~x4 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x64 & ~x65 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x94;
assign c681 = ~x50;
assign c683 = ~x1;
assign c685 =  x1 &  x2 &  x6 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x78 &  x79 &  x86 &  x87 &  x88 & ~x0 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x34 & ~x45 & ~x52 & ~x53 & ~x55 & ~x63 & ~x64 & ~x65 & ~x75 & ~x84 & ~x85 & ~x94 & ~x95;
assign c687 = ~x2 & ~x3;
assign c689 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x9 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c691 =  x3 &  x4 & ~x0 & ~x74;
assign c693 =  x16 &  x17 &  x37 &  x38 &  x39 &  x47 &  x50 &  x51 &  x60 &  x67 &  x68 &  x71 &  x77 &  x79 &  x80 &  x89 & ~x0 & ~x10 & ~x23 & ~x25 & ~x35 & ~x43 & ~x54 & ~x62 & ~x73 & ~x84;
assign c695 =  x33;
assign c699 = ~x1;
assign c6101 =  x2 &  x16 &  x17 &  x19 &  x20 &  x28 &  x29 &  x36 &  x47 &  x49 &  x51 &  x58 &  x59 &  x76 &  x80 &  x88 &  x89 & ~x22 & ~x25 & ~x32 & ~x33 & ~x43 & ~x45 & ~x52 & ~x65 & ~x72 & ~x73 & ~x82 & ~x92 & ~x93;
assign c6103 =  x33;
assign c6105 =  x19 &  x31 & ~x2 & ~x6 & ~x7;
assign c6107 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x61 & ~x63 & ~x65 & ~x72 & ~x73 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x94 & ~x95;
assign c6109 =  x16 &  x18 &  x20 &  x27 &  x29 &  x40 &  x47 &  x48 &  x49 &  x50 &  x66 &  x70 &  x76 &  x77 &  x87 &  x88 &  x90 & ~x2 & ~x22 & ~x25 & ~x33 & ~x35 & ~x44 & ~x45 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x82 & ~x83 & ~x85 & ~x93 & ~x94;
assign c6111 =  x17 &  x20 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x58 &  x59 &  x66 &  x67 &  x69 &  x70 &  x71 &  x76 &  x78 &  x79 &  x86 &  x88 &  x89 &  x90 & ~x0 & ~x22 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x94;
assign c6113 =  x33;
assign c6115 =  x21 &  x40 &  x67 &  x69 &  x71 &  x79 &  x89 &  x90 & ~x0 & ~x32 & ~x35 & ~x72 & ~x92;
assign c6117 =  x5 &  x26 &  x28 &  x56 &  x76 &  x77 &  x86 &  x87 &  x88 & ~x4 & ~x24 & ~x43 & ~x84;
assign c6119 =  x20 &  x27 &  x29 &  x38 &  x39 &  x40 &  x41 &  x50 &  x51 &  x56 &  x58 &  x69 &  x77 &  x80 &  x86 &  x91 & ~x0 & ~x22 & ~x24 & ~x33 & ~x34 & ~x35 & ~x52 & ~x53 & ~x54 & ~x62 & ~x65 & ~x72 & ~x75 & ~x82 & ~x83 & ~x84 & ~x95;
assign c6121 = ~x2 & ~x5;
assign c6123 =  x55;
assign c6125 =  x1 &  x2 &  x6 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x4 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c6127 =  x19 & ~x2;
assign c6129 =  x74;
assign c6131 =  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x30 &  x37 &  x38 &  x46 &  x56 &  x57 &  x66 &  x68 &  x76 &  x78 &  x87 &  x90 & ~x2 & ~x32 & ~x34 & ~x35 & ~x42 & ~x44 & ~x45 & ~x52 & ~x63 & ~x73 & ~x74 & ~x75 & ~x82 & ~x84 & ~x85;
assign c6133 = ~x1;
assign c6135 =  x9 &  x26 &  x29 &  x31 &  x36 &  x39 &  x46 &  x47 &  x50 &  x56 &  x68 &  x70 &  x71 &  x77 &  x86 &  x87 &  x89 &  x90 & ~x22 & ~x24 & ~x34 & ~x35 & ~x42 & ~x44 & ~x45 & ~x55 & ~x63 & ~x75 & ~x81 & ~x82 & ~x83 & ~x92 & ~x94 & ~x95;
assign c6137 = ~x39;
assign c6139 = ~x1;
assign c6141 = ~x1;
assign c6143 =  x54;
assign c6145 =  x11 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x29 &  x30 &  x31 &  x39 &  x40 &  x46 &  x47 &  x49 &  x50 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x69 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x89 &  x90 &  x91 & ~x0 & ~x22 & ~x24 & ~x42 & ~x45 & ~x52 & ~x54 & ~x62 & ~x65 & ~x73 & ~x74 & ~x84 & ~x85 & ~x94 & ~x95;
assign c6147 =  x1 &  x2 &  x6 &  x7 &  x16 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x4 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x85;
assign c6149 = ~x1;
assign c6151 = ~x2 & ~x6 & ~x7;
assign c6153 =  x1 &  x5 &  x26 &  x36 &  x46 &  x67 &  x68 &  x76 &  x78 &  x79 &  x88 &  x89 &  x90 & ~x4 & ~x33 & ~x44 & ~x45 & ~x55 & ~x75;
assign c6157 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x71 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x44 & ~x45 & ~x53 & ~x54 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c6159 = ~x50;
assign c6161 = ~x86;
assign c6163 = ~x31;
assign c6165 =  x33;
assign c6167 = ~x2 & ~x5;
assign c6169 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x31 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x89 &  x91 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c6171 = ~x90;
assign c6173 = ~x40;
assign c6175 =  x52;
assign c6177 = ~x47;
assign c6181 = ~x2 & ~x6 & ~x7;
assign c6183 =  x3 & ~x51;
assign c6185 = ~x1;
assign c6187 = ~x2;
assign c6189 = ~x2;
assign c6191 =  x6 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x46 &  x47 &  x48 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 & ~x0 & ~x4 & ~x22 & ~x23 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x95;
assign c6193 =  x19 &  x20 &  x21 &  x28 &  x31 &  x36 &  x38 &  x40 &  x47 &  x49 &  x67 &  x68 &  x71 &  x79 &  x80 &  x89 & ~x22 & ~x23 & ~x24 & ~x32 & ~x33 & ~x34 & ~x45 & ~x72 & ~x81 & ~x84 & ~x85 & ~x92 & ~x94;
assign c6195 =  x52;
assign c6197 =  x1 &  x2 &  x16 &  x18 &  x20 &  x26 &  x28 &  x30 &  x36 &  x38 &  x39 &  x41 &  x46 &  x47 &  x48 &  x49 &  x51 &  x57 &  x58 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x79 &  x80 &  x88 &  x89 & ~x22 & ~x23 & ~x24 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x52 & ~x53 & ~x55 & ~x62 & ~x63 & ~x75 & ~x81 & ~x83 & ~x92 & ~x94 & ~x95;
assign c6199 = ~x1;
assign c6201 = ~x1;
assign c6203 = ~x40;
assign c6205 = ~x30;
assign c6207 = ~x4;
assign c6209 = ~x58;
assign c6211 =  x1 &  x4 &  x16 &  x17 &  x18 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x76 &  x77 &  x86 &  x87 &  x88 & ~x5 & ~x6 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x84 & ~x85 & ~x94 & ~x95;
assign c6213 = ~x88;
assign c6215 =  x1 &  x2 &  x16 &  x17 &  x18 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x76 &  x77 &  x86 &  x87 & ~x0 & ~x3 & ~x5 & ~x7 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x71 & ~x72 & ~x73 & ~x74 & ~x75 & ~x94 & ~x95;
assign c6217 = ~x2;
assign c6219 = ~x1;
assign c6221 = ~x2 & ~x3;
assign c6223 = ~x1;
assign c6225 =  x24;
assign c6227 = ~x4;
assign c6229 =  x53;
assign c6231 = ~x86;
assign c6233 = ~x50;
assign c6235 =  x5 &  x17 &  x18 &  x29 &  x30 &  x46 &  x47 &  x48 &  x66 &  x77 &  x86 &  x88 & ~x24 & ~x35 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x63 & ~x65 & ~x84 & ~x85 & ~x93 & ~x95;
assign c6237 =  x84;
assign c6239 = ~x48;
assign c6243 =  x1 &  x5 &  x20 &  x26 &  x46 &  x49 &  x51 &  x59 &  x66 &  x69 &  x71 &  x78 &  x87 &  x91 & ~x22 & ~x34 & ~x53 & ~x63 & ~x72 & ~x93;
assign c6245 = ~x2 & ~x3;
assign c6247 = ~x1;
assign c6249 =  x16 &  x17 &  x18 &  x20 &  x26 &  x27 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x47 &  x48 &  x56 &  x58 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x79 &  x80 &  x88 &  x90 & ~x0 & ~x22 & ~x25 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x81 & ~x83 & ~x92 & ~x93;
assign c6251 =  x24;
assign c6253 = ~x30;
assign c6255 =  x42;
assign c6257 = ~x2 & ~x6 & ~x7;
assign c6259 = ~x2 & ~x5;
assign c6261 = ~x38;
assign c6263 =  x69 &  x76 &  x80 &  x89 &  x91 & ~x0 & ~x22 & ~x32 & ~x43 & ~x55 & ~x72 & ~x92;
assign c6265 =  x18 &  x26 &  x27 &  x28 &  x30 &  x36 &  x40 &  x46 &  x48 &  x49 &  x56 &  x60 &  x66 &  x68 &  x70 &  x71 &  x76 &  x79 &  x80 &  x86 &  x87 &  x90 & ~x0 & ~x22 & ~x23 & ~x25 & ~x33 & ~x35 & ~x53 & ~x54 & ~x55 & ~x64 & ~x72 & ~x74 & ~x75 & ~x82 & ~x83 & ~x92 & ~x93 & ~x94;
assign c6267 =  x16 &  x17 &  x18 &  x26 &  x27 &  x28 &  x29 &  x36 &  x38 &  x39 &  x40 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x22 & ~x24 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x65 & ~x73 & ~x74 & ~x75 & ~x81 & ~x82 & ~x83 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c6269 = ~x50;
assign c6271 =  x5 &  x28 &  x40 &  x48 &  x49 &  x58 &  x59 &  x88 &  x89 & ~x4 & ~x24 & ~x32 & ~x63 & ~x75;
assign c6273 =  x75;
assign c6275 =  x1 &  x19 &  x38 &  x56 &  x78 & ~x2 & ~x21 & ~x25 & ~x32 & ~x34 & ~x44 & ~x54 & ~x73;
assign c6277 =  x1 &  x16 &  x18 &  x19 &  x20 &  x29 &  x30 &  x39 &  x46 &  x48 &  x50 &  x58 &  x68 &  x70 &  x77 &  x80 &  x86 &  x89 &  x90 & ~x2 & ~x22 & ~x25 & ~x34 & ~x44 & ~x53 & ~x65 & ~x83 & ~x93;
assign c6279 = ~x30;
assign c6281 = ~x2;
assign c6283 =  x42 & ~x0 & ~x81;
assign c6285 = ~x1;
assign c6287 =  x4 & ~x2 & ~x6 & ~x7 & ~x33;
assign c6289 = ~x2 & ~x3;
assign c6291 = ~x1;
assign c6293 =  x1 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x29 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x78 &  x79 &  x80 &  x86 &  x87 &  x89 &  x90 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x53 & ~x61 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c6295 =  x1 &  x5 &  x17 &  x19 &  x20 &  x26 &  x28 &  x37 &  x39 &  x40 &  x46 &  x47 &  x48 &  x56 &  x59 &  x67 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 & ~x4 & ~x24 & ~x34 & ~x35 & ~x44 & ~x45 & ~x54 & ~x65 & ~x75 & ~x85;
assign c6297 =  x52;
assign c6299 =  x5 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x37 &  x38 &  x47 &  x57 &  x58 &  x66 &  x78 &  x86 &  x87 & ~x4 & ~x34 & ~x35 & ~x43 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64;
assign c6301 = ~x2 & ~x88;
assign c6303 = ~x2 & ~x5;
assign c6305 =  x75;
assign c6307 =  x31 & ~x2 & ~x7;
assign c6309 =  x71 &  x91 & ~x10 & ~x11 & ~x42;
assign c6311 = ~x2 & ~x5;
assign c6313 = ~x2 & ~x3;
assign c6315 =  x1 &  x5 &  x16 &  x18 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x47 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x67 &  x68 &  x76 &  x87 &  x89 & ~x4 & ~x35 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x65 & ~x75 & ~x84 & ~x85;
assign c6317 =  x1 &  x5 &  x17 &  x18 &  x29 &  x38 &  x48 &  x49 &  x57 &  x59 &  x67 &  x68 &  x76 &  x78 & ~x4 & ~x25 & ~x33 & ~x34 & ~x35 & ~x43 & ~x54 & ~x65 & ~x84;
assign c6319 = ~x40;
assign c6321 = ~x0 & ~x9;
assign c6323 =  x16 &  x19 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x47 &  x48 &  x50 &  x56 &  x58 &  x66 &  x76 &  x77 &  x86 &  x87 & ~x2 & ~x22 & ~x23 & ~x25 & ~x33 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x64 & ~x72 & ~x74 & ~x82 & ~x83 & ~x85 & ~x93 & ~x94 & ~x95;
assign c6327 = ~x40;
assign c6329 = ~x2;
assign c6331 =  x1 &  x16 &  x17 &  x19 &  x20 &  x26 &  x28 &  x29 &  x30 &  x36 &  x37 &  x39 &  x40 &  x46 &  x47 &  x56 &  x57 &  x58 &  x60 &  x66 &  x67 &  x68 &  x69 &  x76 &  x78 &  x80 &  x86 &  x88 &  x89 &  x90 &  x91 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x61 & ~x63 & ~x64 & ~x73 & ~x74 & ~x82 & ~x83 & ~x84 & ~x92 & ~x93 & ~x95;
assign c6333 = ~x38;
assign c6335 = ~x76;
assign c6337 = ~x2;
assign c6339 =  x53;
assign c6341 =  x52;
assign c6343 =  x33;
assign c6345 =  x20 &  x59 &  x88 &  x91 & ~x21 & ~x35 & ~x73;
assign c6347 = ~x1;
assign c6349 =  x4 &  x16 &  x17 &  x19 &  x20 &  x27 &  x58 & ~x5 & ~x7 & ~x53 & ~x54 & ~x75 & ~x84;
assign c6351 = ~x18;
assign c6353 =  x1 &  x3 &  x6 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 & ~x0 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x94 & ~x95;
assign c6355 =  x52;
assign c6357 = ~x1;
assign c6359 = ~x2;
assign c6361 = ~x1;
assign c6363 =  x1 &  x6 &  x7 &  x16 &  x17 &  x19 &  x20 &  x27 &  x28 &  x29 &  x36 &  x37 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x58 &  x59 &  x60 &  x66 &  x67 &  x69 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x4 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x44 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x84 & ~x85 & ~x94 & ~x95;
assign c6367 = ~x1;
assign c6369 =  x1 &  x2 &  x6 &  x7 &  x16 &  x17 &  x18 &  x19 &  x26 &  x27 &  x28 &  x29 &  x30 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x76 &  x77 &  x78 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x4 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x85 & ~x93 & ~x94 & ~x95;
assign c6371 =  x6 &  x7 &  x16 &  x19 &  x21 &  x29 &  x36 &  x37 &  x59 &  x76 &  x77 &  x78 & ~x4 & ~x24 & ~x34 & ~x35 & ~x43 & ~x45 & ~x55 & ~x64;
assign c6373 =  x65;
assign c6375 = ~x31;
assign c6379 =  x3 &  x5 &  x80 & ~x0;
assign c6381 = ~x1;
assign c6383 =  x10 & ~x70;
assign c6385 = ~x2 & ~x3;
assign c6387 =  x2 &  x17 &  x18 &  x19 &  x26 &  x27 &  x29 &  x30 &  x36 &  x37 &  x39 &  x40 &  x46 &  x47 &  x48 &  x50 &  x60 &  x66 &  x67 &  x69 &  x70 &  x71 &  x78 &  x80 &  x89 & ~x24 & ~x25 & ~x33 & ~x34 & ~x35 & ~x42 & ~x53 & ~x54 & ~x55 & ~x62 & ~x64 & ~x65 & ~x73 & ~x74 & ~x81 & ~x82 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c6389 =  x16 &  x17 &  x18 &  x20 &  x27 &  x29 &  x31 &  x37 &  x38 &  x40 &  x48 &  x49 &  x51 &  x56 &  x57 &  x59 &  x60 &  x68 &  x69 &  x70 &  x77 &  x78 &  x80 &  x86 &  x88 &  x89 & ~x0 & ~x22 & ~x23 & ~x24 & ~x25 & ~x33 & ~x34 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x62 & ~x63 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x84 & ~x92 & ~x94 & ~x95;
assign c6391 =  x3 &  x4 & ~x0;
assign c6393 = ~x2 & ~x5;
assign c6395 =  x84;
assign c6397 = ~x1;
assign c6399 = ~x2 & ~x5;
assign c6401 = ~x2;
assign c6403 = ~x40;
assign c6405 =  x20 &  x29 &  x30 &  x36 &  x37 &  x39 &  x40 &  x46 &  x50 &  x51 &  x57 &  x58 &  x59 &  x67 &  x68 &  x71 &  x78 &  x79 &  x80 & ~x0 & ~x22 & ~x24 & ~x35 & ~x44 & ~x45 & ~x52 & ~x63 & ~x81 & ~x83 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c6407 =  x10 & ~x69;
assign c6409 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x28 &  x29 &  x30 &  x31 &  x36 &  x38 &  x39 &  x40 &  x41 &  x47 &  x48 &  x49 &  x50 &  x56 &  x59 &  x66 &  x67 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x0 & ~x22 & ~x24 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x62 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c6411 =  x1 &  x7 &  x20 &  x26 &  x27 &  x29 &  x30 &  x37 &  x46 &  x48 &  x51 &  x57 &  x59 &  x70 &  x78 &  x79 &  x80 &  x89 & ~x24 & ~x25 & ~x52 & ~x53 & ~x54 & ~x62 & ~x63 & ~x65 & ~x74 & ~x81 & ~x83 & ~x84 & ~x85 & ~x93;
assign c6413 =  x19 &  x26 &  x28 &  x30 &  x31 &  x49 &  x58 &  x68 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 & ~x2 & ~x22 & ~x24 & ~x32 & ~x34 & ~x45 & ~x83 & ~x85;
assign c6415 =  x84 & ~x2;
assign c6417 = ~x1;
assign c6419 = ~x40;
assign c6421 = ~x56;
assign c6423 =  x1 &  x16 &  x19 &  x27 &  x28 &  x30 &  x31 &  x36 &  x38 &  x39 &  x48 &  x49 &  x56 &  x58 &  x59 &  x66 &  x68 &  x71 &  x77 &  x78 &  x79 &  x80 &  x88 &  x89 &  x91 & ~x22 & ~x23 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x42 & ~x43 & ~x45 & ~x53 & ~x54 & ~x55 & ~x64 & ~x65 & ~x72 & ~x73 & ~x83 & ~x85 & ~x92 & ~x93 & ~x95;
assign c6425 =  x3 &  x10 &  x79 &  x91 & ~x0 & ~x72;
assign c6427 =  x1 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x50 &  x56 &  x57 &  x58 &  x59 &  x60 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x33 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x61 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c6429 = ~x1;
assign c6431 = ~x2 & ~x3;
assign c6433 = ~x5;
assign c6435 =  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x41 &  x46 &  x47 &  x48 &  x49 &  x51 &  x56 &  x57 &  x59 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x78 &  x79 &  x80 &  x86 &  x87 &  x89 &  x90 &  x91 & ~x22 & ~x23 & ~x24 & ~x25 & ~x32 & ~x34 & ~x35 & ~x43 & ~x44 & ~x45 & ~x52 & ~x53 & ~x54 & ~x55 & ~x62 & ~x63 & ~x64 & ~x65 & ~x72 & ~x73 & ~x74 & ~x83 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94 & ~x95;
assign c6437 = ~x50;
assign c6439 = ~x1;
assign c6441 = ~x79;
assign c6443 = ~x1;
assign c6445 =  x42;
assign c6447 =  x42 & ~x81;
assign c6449 =  x93 & ~x0 & ~x5;
assign c6451 = ~x2 & ~x5;
assign c6455 =  x33;
assign c6457 =  x3 &  x6 &  x16 &  x20 &  x30 &  x31 &  x38 &  x40 &  x48 &  x51 &  x56 &  x58 &  x59 &  x69 &  x76 &  x77 &  x78 &  x79 &  x87 & ~x0 & ~x23 & ~x24 & ~x25 & ~x33 & ~x43 & ~x44 & ~x52 & ~x54 & ~x55 & ~x64 & ~x73 & ~x74 & ~x84 & ~x94 & ~x95;
assign c6459 = ~x7;
assign c6461 = ~x1;
assign c6463 =  x5 &  x16 &  x17 &  x18 &  x26 &  x27 &  x36 &  x37 &  x39 &  x46 &  x56 &  x76 &  x77 &  x78 &  x89 &  x90 & ~x4 & ~x23 & ~x24 & ~x25 & ~x34 & ~x35 & ~x43 & ~x64 & ~x65 & ~x75;
assign c6465 =  x33;
assign c6467 = ~x50;
assign c6469 =  x84;
assign c6471 = ~x1;
assign c6473 = ~x40;
assign c6475 =  x25;
assign c6477 = ~x1;
assign c6479 =  x49 & ~x2 & ~x6 & ~x7;
assign c6481 = ~x1;
assign c6483 = ~x50;
assign c6485 =  x1 &  x6 &  x17 &  x18 &  x19 &  x26 &  x29 &  x30 &  x36 &  x38 &  x39 &  x46 &  x48 &  x50 &  x56 &  x66 &  x67 &  x68 &  x76 &  x86 & ~x0 & ~x4 & ~x22 & ~x24 & ~x32 & ~x33 & ~x34 & ~x43 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x75 & ~x82 & ~x85 & ~x94 & ~x95;
assign c6487 =  x1 &  x17 &  x19 &  x20 &  x29 &  x37 &  x38 &  x40 &  x41 &  x46 &  x49 &  x50 &  x56 &  x57 &  x66 &  x67 &  x68 &  x69 &  x70 &  x76 &  x77 &  x80 &  x86 &  x87 &  x88 &  x89 &  x90 & ~x22 & ~x25 & ~x33 & ~x34 & ~x35 & ~x44 & ~x54 & ~x61 & ~x62 & ~x74 & ~x75 & ~x84 & ~x85 & ~x92 & ~x93 & ~x94;
assign c6489 =  x52;
assign c6491 =  x1 &  x2 &  x6 &  x7 &  x16 &  x17 &  x18 &  x19 &  x20 &  x26 &  x27 &  x28 &  x29 &  x30 &  x31 &  x36 &  x37 &  x38 &  x39 &  x40 &  x46 &  x47 &  x48 &  x49 &  x50 &  x51 &  x56 &  x57 &  x58 &  x59 &  x66 &  x67 &  x68 &  x76 &  x77 &  x79 &  x86 &  x87 &  x88 &  x89 & ~x4 & ~x23 & ~x24 & ~x25 & ~x32 & ~x34 & ~x35 & ~x42 & ~x43 & ~x44 & ~x45 & ~x53 & ~x54 & ~x55 & ~x63 & ~x64 & ~x65 & ~x75 & ~x83 & ~x85 & ~x94 & ~x95;
assign c6493 = ~x2 & ~x3;
assign c6495 = ~x2 & ~x4;
assign c6497 = ~x2;
assign c6499 =  x42;

endmodule