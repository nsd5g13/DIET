module tm( x0,x1,x2,x3,x4,x5,x6,x7,x8,x9,x10,x11,x12,x13,x14,x15,x16,x17,x18,x19,x20,x21,x22,x23,x24,x25,x26,x27,x28,x29,x30,x31,x32,x33,x34,x35,x36,x37,x38,x39,x40,x41,x42,x43,x44,x45,x46,x47,x48,x49,x50,x51,x52,x53,x54,x55,x56,x57,x58,x59,x60,x61,x62,x63,x64,x65,x66,x67,x68,x69,x70,x71,x72,x73,x74,x75,x76,x77,x78,x79,x80,x81,x82,x83,x84,x85,x86,x87,x88,x89,x90,x91,x92,x93,x94,x95,x96,x97,x98,x99,x100,x101,x102,x103,x104,x105,x106,x107,x108,x109,x110,x111,x112,x113,x114,x115,x116,x117,x118,x119,x120,x121,x122,x123,x124,x125,x126,x127,x128,x129,x130,x131,x132,x133,x134,x135,x136,x137,x138,x139,x140,x141,x142,x143,x144,x145,x146,x147,x148,x149,x150,x151,x152,x153,x154,x155,x156,x157,x158,x159,x160,x161,x162,x163,x164,x165,x166,x167,x168,x169,x170,x171,x172,x173,x174,x175,x176,x177,x178,x179,x180,x181,x182,x183,x184,x185,x186,x187,x188,x189,x190,x191,x192,x193,x194,x195,x196,x197,x198,x199,x200,x201,x202,x203,x204,x205,x206,x207,x208,x209,x210,x211,x212,x213,x214,x215,x216,x217,x218,x219,x220,x221,x222,x223,x224,x225,x226,x227,x228,x229,x230,x231,x232,x233,x234,x235,x236,x237,x238,x239,x240,x241,x242,x243,x244,x245,x246,x247,x248,x249,x250,x251,x252,x253,x254,x255,x256,x257,x258,x259,x260,x261,x262,x263,x264,x265,x266,x267,x268,x269,x270,x271,x272,x273,x274,x275,x276,x277,x278,x279,x280,x281,x282,x283,x284,x285,x286,x287,x288,x289,x290,x291,x292,x293,x294,x295,x296,x297,x298,x299,x300,x301,x302,x303,x304,x305,x306,x307,x308,x309,x310,x311,x312,x313,x314,x315,x316,x317,x318,x319,x320,x321,x322,x323,x324,x325,x326,x327,x328,x329,x330,x331,x332,x333,x334,x335,x336,x337,x338,x339,x340,x341,x342,x343,x344,x345,x346,x347,x348,x349,x350,x351,x352,x353,x354,x355,x356,x357,x358,x359,x360,x361,x362,x363,x364,x365,x366,x367,x368,x369,x370,x371,x372,x373,x374,x375,x376,x377,x378,x379,x380,x381,x382,x383,x384,x385,x386,x387,x388,x389,x390,x391,x392,x393,x394,x395,x396,x397,x398,x399,x400,x401,x402,x403,x404,x405,x406,x407,x408,x409,x410,x411,x412,x413,x414,x415,x416,x417,x418,x419,x420,x421,x422,x423,x424,x425,x426,x427,x428,x429,x430,x431,x432,x433,x434,x435,x436,x437,x438,x439,x440,x441,x442,x443,x444,x445,x446,x447,x448,x449,x450,x451,x452,x453,x454,x455,x456,x457,x458,x459,x460,x461,x462,x463,x464,x465,x466,x467,x468,x469,x470,x471,x472,x473,x474,x475,x476,x477,x478,x479,x480,x481,x482,x483,x484,x485,x486,x487,x488,x489,x490,x491,x492,x493,x494,x495,x496,x497,x498,x499,x500,x501,x502,x503,x504,x505,x506,x507,x508,x509,x510,x511,x512,x513,x514,x515,x516,x517,x518,x519,x520,x521,x522,x523,x524,x525,x526,x527,x528,x529,x530,x531,x532,x533,x534,x535,x536,x537,x538,x539,x540,x541,x542,x543,x544,x545,x546,x547,x548,x549,x550,x551,x552,x553,x554,x555,x556,x557,x558,x559,x560,x561,x562,x563,x564,x565,x566,x567,x568,x569,x570,x571,x572,x573,x574,x575,x576,x577,x578,x579,x580,x581,x582,x583,x584,x585,x586,x587,x588,x589,x590,x591,x592,x593,x594,x595,x596,x597,x598,x599,x600,x601,x602,x603,x604,x605,x606,x607,x608,x609,x610,x611,x612,x613,x614,x615,x616,x617,x618,x619,x620,x621,x622,x623,x624,x625,x626,x627,x628,x629,x630,x631,x632,x633,x634,x635,x636,x637,x638,x639,x640,x641,x642,x643,x644,x645,x646,x647,x648,x649,x650,x651,x652,x653,x654,x655,x656,x657,x658,x659,x660,x661,x662,x663,x664,x665,x666,x667,x668,x669,x670,x671,x672,x673,x674,x675,x676,x677,x678,x679,x680,x681,x682,x683,x684,x685,x686,x687,x688,x689,x690,x691,x692,x693,x694,x695,x696,x697,x698,x699,x700,x701,x702,x703,x704,x705,x706,x707,x708,x709,x710,x711,x712,x713,x714,x715,x716,x717,x718,x719,x720,x721,x722,x723,x724,x725,x726,x727,x728,x729,x730,x731,x732,x733,x734,x735,x736,x737,x738,x739,x740,x741,x742,x743,x744,x745,x746,x747,x748,x749,x750,x751,x752,x753,x754,x755,x756,x757,x758,x759,x760,x761,x762,x763,x764,x765,x766,x767,x768,x769,x770,x771,x772,x773,x774,x775,x776,x777,x778,x779,x780,x781,x782,x783,c8238,c7311,c2224,c3391,c0356,c0309,c8324,c1433,c447,c594,c1176,c6238,c5458,c1360,c4293,c6236,c3480,c5353,c4243,c1154,c090,c0280,c7271,c625,c4371,c5488,c7259,c3355,c4200,c1355,c898,c5429,c7243,c2112,c2430,c8216,c155,c4435,c2171,c882,c5365,c5424,c661,c4483,c6335,c2218,c2358,c7372,c3298,c1349,c8370,c2275,c151,c2370,c7153,c6306,c1292,c7401,c872,c5284,c252,c813,c921,c3135,c6135,c2272,c4185,c6466,c5478,c0131,c5371,c672,c11,c3130,c0460,c6499,c5173,c643,c6221,c248,c4460,c2292,c6256,c4201,c7220,c4120,c6284,c1114,c3468,c958,c1243,c4378,c3166,c7232,c4142,c674,c1208,c9363,c7430,c4158,c111,c8414,c3487,c7446,c050,c6384,c1256,c2242,c33,c054,c0298,c5491,c878,c438,c56,c6333,c982,c7161,c17,c1417,c8108,c837,c2300,c9456,c174,c3435,c8346,c526,c152,c0193,c6259,c4324,c9264,c3296,c0187,c7280,c8301,c6383,c9432,c1340,c5402,c4487,c3206,c9339,c310,c2201,c4242,c6242,c5431,c7484,c8356,c6409,c02,c9202,c2193,c9197,c2438,c8343,c9468,c8368,c5418,c8189,c8469,c3280,c0117,c4325,c5169,c5280,c074,c1211,c4181,c0304,c4427,c436,c191,c8265,c9379,c6397,c1363,c4348,c4179,c845,c2197,c9480,c5253,c9109,c1437,c6245,c3100,c942,c824,c6125,c8194,c8450,c8338,c1139,c8418,c38,c4245,c947,c541,c158,c265,c2221,c8197,c082,c2226,c3378,c8458,c4277,c0328,c6477,c2348,c4123,c4394,c3445,c3372,c1315,c6427,c4192,c9252,c9326,c6181,c8135,c7276,c5413,c9453,c2154,c0282,c3241,c6295,c6382,c2410,c4270,c0237,c232,c2465,c4381,c127,c150,c7371,c4233,c855,c1431,c3218,c1248,c2375,c1117,c6280,c8495,c573,c3396,c2158,c172,c0105,c4311,c2334,c2160,c678,c010,c8272,c6195,c2376,c8396,c5468,c67,c4391,c1104,c0299,c6344,c0224,c8127,c2346,c715,c660,c0429,c721,c2170,c9274,c312,c9455,c5140,c7149,c1423,c3427,c3335,c3244,c3348,c6141,c8257,c2283,c7469,c3159,c0386,c7164,c7320,c4109,c3179,c0235,c767,c5144,c6334,c4498,c0301,c2212,c9140,c544,c3326,c348,c7154,c474,c475,c2187,c341,c7369,c1409,c6229,c6170,c82,c5354,c9411,c365,c5302,c9142,c2259,c812,c3327,c5441,c3395,c463,c945,c2342,c2174,c0365,c5374,c94,c9174,c0389,c9131,c6365,c2281,c7303,c6289,c273,c9106,c1199,c7270,c8274,c4269,c7112,c3461,c6278,c1322,c0121,c7464,c673,c0170,c5333,c3421,c2387,c026,c4218,c5480,c230,c546,c584,c913,c7162,c6310,c1257,c3137,c6401,c3369,c9180,c3278,c0422,c6122,c1399,c0234,c2449,c6426,c6343,c2109,c6468,c6193,c169,c1412,c3132,c7101,c944,c9436,c1185,c520,c5124,c2326,c0379,c9290,c640,c3172,c8134,c765,c8440,c1454,c7425,c3129,c7116,c554,c598,c8276,c8145,c7221,c373,c4207,c5182,c3410,c1387,c4261,c123,c124,c2111,c069,c292,c1375,c677,c4300,c5330,c7485,c2217,c3307,c7419,c1283,c5394,c4428,c5219,c4422,c578,c3371,c4276,c4376,c1175,c3367,c6451,c828,c0362,c1233,c1195,c4164,c5421,c750,c5249,c9428,c926,c9417,c3401,c5203,c9120,c2405,c8120,c453,c6173,c4363,c0452,c8220,c5324,c8410,c6430,c8123,c0263,c1366,c5148,c2440,c8192,c9145,c0394,c3323,c4336,c1448,c0339,c5289,c2454,c2310,c8153,c1462,c6434,c5412,c7121,c2118,c148,c1141,c494,c5447,c3476,c0238,c0122,c973,c8404,c2391,c9205,c4190,c9403,c9254,c1266,c8481,c9158,c9136,c857,c3162,c8201,c5114,c1328,c9380,c166,c4256,c8491,c994,c6108,c330,c4306,c0127,c0376,c6304,c5137,c636,c3169,c6227,c7340,c7314,c55,c6348,c2386,c2280,c8184,c5361,c071,c2403,c6439,c4331,c2196,c5296,c189,c2361,c2415,c6157,c8371,c9209,c4284,c161,c2455,c0189,c4301,c371,c1100,c798,c7454,c8333,c8222,c889,c255,c9165,c4113,c4401,c6201,c1472,c9222,c5464,c0442,c4267,c7102,c6241,c1142,c626,c5310,c0164,c560,c0323,c0271,c6407,c449,c0307,c632,c1113,c2336,c5244,c7200,c9152,c2175,c088,c0229,c2211,c5428,c2227,c326,c5107,c962,c2228,c1353,c3418,c7412,c4161,c2324,c99,c8116,c760,c9425,c2425,c2417,c76,c42,c3309,c5462,c9128,c4356,c156,c496,c9334,c8330,c5479,c1204,c0286,c0120,c7323,c911,c8292,c3158,c0216,c2492,c5454,c421,c2349,c3358,c4407,c9323,c6474,c8415,c3328,c545,c4316,c0126,c9465,c028,c1258,c1157,c6375,c417,c1441,c9329,c1183,c491,c0269,c7302,c6381,c6161,c1140,c5298,c0469,c793,c740,c359,c610,c492,c5294,c290,c5326,c7351,c826,c286,c8428,c6286,c4477,c9198,c9275,c5134,c9451,c2433,c8334,c1476,c3313,c1226,c3190,c7130,c3469,c2318,c185,c2265,c2305,c3282,c8471,c5383,c6362,c1498,c5443,c8214,c8365,c6312,c5337,c1249,c1273,c1300,c5452,c4388,c2467,c680,c1488,c4297,c32,c9315,c411,c7228,c7409,c4280,c1302,c7189,c1336,c3250,c0268,c8489,c5279,c7181,c4247,c1390,c8305,c0487,c194,c3446,c0156,c1389,c8420,c4328,c1215,c3433,c7240,c747,c8316,c4167,c3155,c1136,c1445,c7146,c5494,c774,c8455,c4104,c2289,c1484,c8223,c5293,c8164,c953,c9195,c2140,c0161,c7295,c1324,c8209,c6494,c7173,c3204,c3214,c4106,c8364,c8466,c1430,c241,c7207,c1259,c055,c0132,c5196,c693,c3340,c5271,c0311,c2252,c3268,c3473,c5256,c2115,c6366,c815,c7444,c3160,c7234,c0142,c7266,c3294,c2341,c9291,c8255,c8213,c6103,c7174,c1466,c1343,c8297,c3163,c9235,c6274,c3337,c8394,c051,c7157,c3411,c6352,c8230,c5269,c9313,c6449,c1331,c1110,c6353,c458,c0145,c716,c7187,c818,c1285,c1339,c5103,c451,c454,c8319,c8434,c2328,c5372,c3212,c97,c0230,c4423,c7134,c8186,c1486,c2119,c6483,c2452,c8403,c6452,c6443,c2245,c8101,c434,c823,c5328,c2393,c685,c6249,c0239,c6124,c3108,c9104,c8487,c3393,c6296,c7337,c6140,c0212,c0147,c66,c9385,c8438,c3128,c7279,c038,c4220,c7452,c7145,c9317,c8448,c9439,c791,c4319,c5387,c072,c1229,c1293,c0139,c5455,c861,c9194,c0439,c90,c4229,c3414,c5235,c5432,c1106,c7325,c6217,c162,c3426,c3439,c323,c4114,c5175,c937,c4495,c9355,c8485,c8332,c5396,c1213,c4272,c8309,c6291,c3248,c9210,c8149,c2389,c441,c4490,c6169,c4160,c0138,c382,c2472,c4406,c6264,c6413,c5282,c1179,c1133,c2478,c8401,c05,c7290,c5180,c0162,c7439,c3114,c7109,c4469,c0134,c999,c426,c7343,c2277,c9207,c7250,c7477,c5277,c2264,c6402,c7427,c240,c5135,c836,c029,c1449,c3432,c7410,c8185,c0283,c8442,c8203,c0450,c0399,c4443,c9191,c1305,c6301,c5187,c9306,c6408,c4399,c043,c3290,c650,c1290,c4408,c8315,c4214,c4492,c5236,c1304,c7471,c9259,c4365,c954,c6204,c2404,c5286,c2262,c779,c5313,c274,c4188,c1414,c3255,c1210,c2434,c5498,c2241,c4400,c2480,c2458,c4126,c3381,c3403,c1319,c8241,c135,c8114,c5314,c1272,c5445,c874,c7291,c9437,c2457,c5217,c6471,c777,c4159,c497,c4395,c023,c4102,c1307,c9260,c079,c5362,c4380,c8329,c61,c9310,c6487,c631,c7176,c036,c7330,c1144,c3201,c138,c4402,c9107,c9249,c8247,c2355,c1357,c5411,c8175,c5426,c2339,c2491,c299,c280,c555,c0419,c2340,c048,c629,c0418,c532,c357,c6233,c8493,c0318,c6438,c3161,c0409,c015,c4144,c676,c134,c3232,c0295,c2219,c0293,c0314,c5246,c1458,c1201,c1291,c9175,c0378,c4398,c1347,c9253,c1244,c3270,c618,c4235,c3247,c5204,c7432,c0326,c80,c7208,c3123,c4491,c7193,c0416,c1497,c4292,c4128,c9188,c9467,c0359,c785,c0233,c912,c662,c0231,c8100,c0471,c7496,c5482,c3291,c3287,c0173,c4252,c7365,c6196,c7479,c098,c9176,c8179,c4372,c9123,c9256,c8398,c2347,c8360,c8113,c26,c792,c4318,c8441,c5391,c2151,c0372,c9189,c7195,c8181,c4479,c2448,c1162,c219,c1489,c078,c7177,c0265,c8421,c2150,c192,c0168,c3302,c7186,c3279,c3138,c8300,c6254,c360,c1469,c7169,c6493,c3380,c9459,c784,c2205,c3219,c259,c8278,c968,c7206,c3322,c6360,c485,c0243,c8363,c9200,c7499,c963,c0259,c440,c5177,c4411,c659,c1228,c7281,c227,c2304,c7442,c0249,c5146,c1187,c5250,c4101,c5473,c887,c5202,c62,c159,c1327,c1483,c4335,c9489,c695,c4121,c2311,c3120,c095,c3240,c649,c4143,c461,c375,c1317,c334,c745,c8411,c4458,c2279,c1169,c3472,c3168,c1391,c910,c6320,c628,c424,c2251,c2314,c2141,c0346,c69,c3448,c3254,c413,c2236,c1278,c267,c4386,c9354,c6479,c1194,c9134,c0488,c2412,c6226,c8166,c5106,c9150,c140,c4278,c8497,c420,c032,c667,c0458,c2294,c3239,c3178,c07,c6482,c559,c9450,c0186,c2497,c1383,c0101,c9217,c7133,c2401,c2416,c1107,c627,c1218,c0375,c0447,c3273,c825,c4141,c0445,c1212,c780,c8242,c7141,c92,c8124,c9257,c9345,c764,c4184,c918,c9416,c2315,c2223,c5306,c5380,c167,c4354,c429,c5435,c2469,c60,c6172,c7418,c9356,c3467,c543,c5194,c247,c6458,c343,c6210,c4414,c24,c7236,c5168,c8349,c7472,c6441,c5232,c49,c9105,c1186,c0251,c6191,c2129,c4263,c9283,c2490,c1372,c3269,c2424,c1270,c5496,c0264,c6142,c534,c8159,c3375,c040,c1282,c2200,c8492,c45,c0400,c5319,c665,c5228,c3289,c3419,c8144,c9204,c0148,c6123,c3127,c1122,c362,c2384,c099,c5410,c28,c9299,c216,c1173,c40,c067,c3231,c790,c0114,c5405,c5419,c0197,c950,c0440,c9314,c077,c8252,c6368,c3141,c6455,c36,c8399,c0177,c6246,c8187,c4118,c0451,c1224,c446,c085,c2488,c638,c3385,c585,c8169,c177,c09,c8382,c0130,c4177,c0167,c498,c1150,c094,c2456,c7213,c9384,c372,c768,c34,c024,c25,c2186,c9117,c4205,c7408,c7455,c1180,c875,c5312,c0402,c0437,c48,c8167,c1214,c7275,c8240,c9401,c2317,c564,c0158,c853,c8425,c8476,c4339,c2431,c8224,c3305,c0383,c8484,c646,c457,c4239,c8172,c9348,c0462,c52,c7483,c712,c849,c766,c7128,c514,c2216,c021,c3466,c8110,c3402,c7445,c8443,c0414,c260,c851,c635,c246,c0492,c1358,c4396,c6341,c2266,c2498,c7197,c8325,c3321,c3453,c838,c3424,c7284,c2409,c841,c8464,c1312,c896,c3482,c0496,c8161,c1130,c093,c3389,c985,c7470,c7350,c9155,c3237,c0215,c4285,c0102,c6418,c562,c9161,c0473,c5185,c9182,c2466,c940,c23,c7241,c9292,c31,c7367,c178,c5170,c4148,c734,c0455,c6116,c4127,c9132,c7272,c7406,c1111,c5363,c9469,c483,c4367,c2192,c3374,c9273,c4384,c2437,c5297,c675,c288,c9172,c4456,c7482,c990,c9479,c9298,c7185,c535,c9476,c8447,c4397,c381,c2330,c9496,c0223,c6118,c2214,c4204,c3324,c5122,c0332,c9387,c3494,c9272,c4221,c6194,c276,c8477,c9393,c4232,c5255,c0334,c0116,c3242,c523,c060,c21,c1475,c9395,c6361,c1216,c3266,c5497,c669,c0103,c7288,c5440,c8251,c5223,c8452,c9446,c5199,c1286,c4466,c0274,c2156,c7215,c8208,c7385,c0354,c8146,c1368,c744,c1235,c2177,c746,c2207,c5492,c691,c756,c7120,c9143,c380,c8367,c3346,c9285,c0465,c199,c3471,c053,c5207,c9466,c2383,c5477,c8467,c0349,c8171,c1261,c2208,c262,c8381,c8277,c186,c1496,c0371,c9386,c2378,c7322,c4299,c738,c915,c7138,c6156,c336,c6429,c9399,c0241,c5300,c4186,c955,c6190,c5210,c88,c9370,c3102,c8296,c6475,c3257,c637,c6228,c6112,c515,c3397,c271,c4281,c4410,c1251,c6216,c0136,c5112,c353,c8429,c8388,c4360,c4382,c0482,c3265,c7125,c6447,c5247,c6182,c4482,c7268,c7392,c4488,c9477,c4494,c6391,c4115,c658,c9376,c7405,c684,c786,c0443,c1168,c1170,c0316,c931,c810,c4165,c936,c2209,c547,c8253,c9497,c925,c6215,c5357,c5470,c6389,c7478,c850,c3205,c283,c1188,c1492,c1275,c634,c112,c338,c6442,c58,c1129,c862,c2320,c8160,c3303,c4283,c264,c741,c195,c5299,c176,c1231,c93,c5367,c6218,c8341,c3183,c8227,c2256,c1356,c0163,c4219,c6110,c894,c1246,c6314,c7301,c596,c340,c3113,c7166,c4462,c6386,c5358,c1178,c1264,c8170,c0470,c7399,c1354,c4441,c8210,c6244,c8221,c017,c9138,c775,c2327,c549,c3315,c6425,c114,c9447,c5157,c9358,c8298,c444,c927,c9367,c6199,c6349,c460,c081,c8314,c9365,c9471,c1333,c4343,c1351,c5476,c2253,c7370,c0110,c2360,c416,c7165,c7489,c8486,c835,c1297,c1435,c0258,c1344,c9223,c0250,c1374,c8111,c8354,c039,c225,c5215,c2357,c725,c6114,c7473,c414,c686,c4369,c966,c6354,c9427,c6260,c510,c020,c3134,c8342,c258,c1242,c6219,c7474,c9119,c6130,c9375,c7435,c6356,c2247,c7143,c834,c9475,c6345,c047,c3308,c4342,c250,c8313,c4340,c315,c9337,c8498,c754,c5123,c063,c9216,c0444,c428,c6145,c8431,c8427,c2153,c987,c012,c3230,c8359,c6105,c7468,c1236,c5150,c6371,c867,c3208,c3470,c1223,c2445,c228,c9281,c9301,c9335,c2374,c1125,c4146,c6357,c0474,c7306,c4442,c5189,c29,c184,c6410,c3437,c8225,c5152,c9141,c6177,c9248,c7317,c0353,c3460,c4217,c2225,c394,c175,c9343,c8475,c844,c1143,c8307,c1370,c0310,c415,c193,c5285,c5101,c9168,c0252,c5274,c1237,c3122,c8361,c0185,c3259,c3185,c5242,c7364,c8358,c5119,c3330,c1401,c5188,c9265,c8182,c7231,c6168,c848,c1380,c9359,c164,c452,c7310,c369,c2390,c1485,c1181,c6347,c7417,c7475,c989,c7115,c6326,c1329,c7424,c928,c4129,c1296,c7493,c43,c3317,c3142,c9196,c7449,c9118,c1207,c7394,c2359,c5343,c619,c3184,c8336,c5212,c7386,c04,c8340,c3124,c1422,c0279,c9173,c057,c5471,c1220,c8384,c8306,c014,c8280,c1478,c883,c187,c8321,c2285,c2267,c7168,c2400,c4172,c9346,c1316,c2477,c548,c5305,c0253,c8337,c8419,c4350,c7278,c3188,c9234,c1442,c5335,c8417,c5417,c8432,c731,c450,c8383,c718,c84,c0137,c0245,c671,c3415,c8142,c4417,c933,c1398,c6432,c294,c2476,c0192,c3118,c6331,c8357,c7247,c4438,c9405,c4211,c68,c4162,c688,c5238,c443,c351,c0497,c1203,c6462,c3398,c2139,c7457,c4418,c4264,c9231,c7368,c6406,c3136,c4287,c7363,c287,c4275,c3293,c1450,c0355,c2483,c9181,c9151,c7338,c4334,c6139,c2142,c0342,c7431,c412,c5376,c3262,c1385,c486,c235,c7196,c6265,c2260,c1135,c0499,c6120,c422,c822,c5422,c50,c7205,c8268,c8335,c4375,c1166,c8289,c737,c8320,c9352,c6251,c9311,c3119,c3148,c6363,c6399,c4213,c7248,c3246,c27,c5149,c089,c456,c0387,c183,c4454,c2333,c2319,c1205,c3377,c3339,c7321,c1280,c0266,c6109,c6269,c367,c445,c2407,c3392,c552,c7172,c4116,c0361,c4450,c6138,c751,c6213,c7108,c3111,c7264,c2351,c2474,c8317,c6160,c8283,c7210,c1474,c980,c4244,c0303,c3474,c6311,c513,c2296,c8456,c9250,c1455,c5213,c0438,c9464,c4323,c8390,c871,c2271,c0300,c331,c4327,c3353,c7150,c3365,c425,c5266,c6396,c4176,c4366,c0370,c6250,c6131,c034,c2429,c2379,c0369,c8294,c4266,c2338,c5290,c7233,c6174,c6492,c3479,c2427,c0149,c654,c2234,c663,c20,c9430,c9139,c6137,c877,c6450,c8465,c4447,c9486,c2100,c9338,c7495,c8326,c4326,c4183,c5377,c8318,c8129,c530,c6297,c895,c6186,c0169,c2274,c5221,c6121,c6283,c096,c7267,c08,c879,c0219,c1134,c0113,c384,c78,c814,c4344,c042,c5193,c5252,c9201,c5258,c3215,c1119,c3101,c4282,c7345,c1245,c0154,c2248,c4199,c1338,c5220,c0407,c1174,c1345,c0475,c1403,c0420,c1428,c1427,c8291,c4403,c8380,c3288,c215,c153,c9396,c2366,c2273,c5104,c314,c0174,c8496,c6431,c5161,c6411,c4431,c0207,c1121,c7467,c2309,c4302,c8408,c8323,c9438,c0125,c8200,c7298,c0351,c666,c6147,c8459,c77,c119,c2484,c5110,c6373,c4445,c253,c390,c0277,c7124,c8204,c3150,c3370,c3361,c7342,c9327,c3192,c3457,c876,c5154,c9242,c4476,c1424,c266,c9241,c3404,c86,c970,c795,c6469,c1318,c218,c7334,c3182,c1323,c2302,c5311,c2372,c1313,c3139,c4246,c87,c527,c0182,c9321,c1240,c8375,c770,c2134,c6200,c9316,c6393,c682,c473,c773,c4472,c0213,c3364,c3486,c070,c4426,c1400,c9460,c6307,c3228,c5147,c278,c8446,c6134,c771,c648,c679,c2436,c1127,c6448,c5483,c0175,c5321,c1196,c7198,c8302,c4209,c3116,c237,c692,c9244,c739,c4404,c5218,c1429,c3490,c7421,c6294,c6424,c0373,c586,c4250,c1418,c431,c7201,c3416,c6211,c2444,c7211,c8219,c3344,c5272,c2116,c952,c2329,c9280,c7309,c3144,c616,c2499,c0480,c5457,c1101,c9440,c5227,c0287,c2308,c346,c0153,c137,c1163,c5257,c9478,c5115,c1155,c317,c8295,c0448,c0199,c4208,c6158,c1147,c8479,c3236,c068,c6351,c1308,c978,c8232,c9149,c16,c495,c2133,c6370,c296,c387,c4153,c4187,c2269,c7428,c9286,c2443,c8198,c484,c9233,c0296,c8474,c5270,c6467,c1432,c3264,c1394,c5225,c4265,c9353,c6277,c7359,c2147,c8122,c9276,c493,c6390,c7255,c1276,c6299,c419,c7178,c881,c244,c8173,c524,c917,c0432,c0415,c0247,c220,c7413,c1447,c8254,c7104,c1238,c7438,c4174,c2268,c946,c2291,c8444,c3197,c956,c3352,c3151,c755,c3388,c132,c5465,c5109,c2202,c395,c4119,c7118,c6364,c9277,c061,c4499,c1348,c827,c4421,c2120,c7107,c243,c0226,c2249,c295,c6367,c8439,c5407,c0367,c551,c5323,c019,c2408,c3356,c5197,c0227,c1277,c2354,c0313,c4178,c7105,c9390,c0324,c7123,c9407,c3422,c988,c2493,c5261,c2222,c977,c8387,c5320,c1255,c9404,c9351,c9360,c6346,c9144,c7258,c291,c0248,c1112,c2419,c1410,c6253,c0463,c9307,c9262,c542,c914,c7341,c749,c8269,c7110,c110,c131,c5348,c689,c7216,c3112,c0320,c3354,c5327,c2420,c4258,c4170,c4346,c591,c7466,c3440,c3405,c9113,c4355,c5341,c762,c763,c0278,c7152,c8183,c6179,c2344,c939,c2352,c9295,c6209,c7393,c9178,c1151,c9340,c1197,c7307,c1115,c269,c8157,c6257,c8118,c6394,c9369,c0204,c376,c142,c5172,c6497,c2363,c056,c0391,c5133,c668,c4295,c2421,c4175,c3430,c3225,c9238,c6222,c7226,c5239,c4212,c2494,c9383,c9322,c2121,c9499,c2106,c8190,c4189,c6267,c0178,c455,c1408,c5448,c4459,c9485,c7456,c0179,c5102,c9214,c0201,c2369,c7277,c7103,c6446,c1330,c0352,c8426,c5325,c5308,c0423,c9330,c3253,c5459,c7122,c5142,c8275,c0111,c15,c4455,c0327,c3299,c0106,c0200,c2399,c899,c091,c6164,c9108,c196,c1198,c9402,c0411,c478,c8121,c9372,c2371,c397,c6152,c9415,c4107,c9336,c9341,c2392,c433,c1120,c4374,c8457,c058,c4312,c960,c5100,c459,c6379,c9392,c2331,c7353,c1191,c3284,c251,c761,c2235,c6206,c7335,c2243,c0461,c6263,c2337,c2124,c9493,c4210,c3386,c0100,c472,c8193,c8156,c9484,c9229,c1108,c7265,c2233,c2276,c224,c0467,c858,c683,c9170,c4485,c1473,c7415,c182,c572,c7443,c711,c839,c890,c8199,c9371,c7261,c0424,c6266,c5171,c5381,c1468,c0218,c1379,c7182,c6205,c8109,c96,c2191,c7378,c699,c3496,c4385,c4486,c234,c8155,c2380,c2210,c4286,c0336,c556,c5206,c313,c3351,c6273,c2231,c3481,c9167,c2220,c736,c4349,c4481,c2215,c6243,c4110,c8206,c6208,c0466,c0403,c7390,c8151,c8286,c0398,c611,c2462,c4132,c8264,c568,c3311,c9187,c986,c5434,c8141,c8271,c3384,c4420,c9333,c0128,c5439,c5444,c2442,c9266,c9474,c480,c8461,c0214,c7142,c4238,c3394,c794,c6176,c4268,c3462,c769,c8311,c641,c0344,c690,c329,c8245,c0484,c254,c5400,c389,c7373,c6490,c8366,c168,c1219,c6330,c2131,c9350,c4405,c075,c7362,c0436,c9458,c2377,c1311,c5174,c6106,c272,c18,c0343,c7488,c2244,c080,c4383,c8212,c9121,c1482,c0210,c471,c432,c6189,c8445,c748,c6167,c4122,c0146,c3252,c8215,c1463,c9190,c5451,c0453,c5141,c181,c7179,c3319,c8158,c9452,c8119,c4130,c3193,c7188,c0498,c2485,c5121,c9166,c5359,c866,c9137,c9101,c8228,c0392,c1262,c7331,c1131,c0388,c3316,c6392,c7225,c670,c3332,c6317,c561,c5222,c840,c920,c035,c7230,c5385,c1126,c3233,c8136,c4138,c64,c0291,c7254,c022,c7273,c6332,c2135,c5181,c5347,c6175,c30,c4288,c8233,c870,c2254,c0180,c4453,c5481,c2288,c9193,c342,c6358,c4193,c9377,c971,c6470,c7358,c1303,c393,c3441,c9441,c3436,c7333,c7462,c1301,c533,c7416,c512,c9126,c3464,c5248,c0184,c4262,c279,c3217,c115,c5234,c984,c5364,c8130,c8102,c1386,c8262,c1165,c3131,c1415,c117,c4437,c1470,c213,c6154,c967,c9294,c4223,c2213,c5420,c5155,c319,c2381,c727,c0255,c820,c2323,c3210,c229,c5344,c5138,c2278,c7313,c7147,c5336,c930,c7274,c339,c3413,c7167,c5129,c592,c7384,c8372,c7404,c5389,c6188,c81,c2188,c5404,c8322,c318,c8327,c7119,c8202,c7171,c8347,c10,c6350,c0292,c0254,c2411,c6465,c0363,c22,c355,c1487,c423,c9304,c789,c3407,c0408,c4182,c7304,c0202,c717,c787,c7346,c0425,c9433,c5153,c5368,c2418,c3149,c8259,c6329,c5263,c3181,c180,c1420,c4361,c2203,c4155,c466,c7366,c3207,c7360,c6324,c1160,c1269,c3498,c0493,c7319,c819,c4329,c9413,c65,c165,c3412,c1459,c577,c146,c1289,c1287,c9240,c8237,c4253,c3484,c1309,c9203,c856,c6318,c6119,c0350,c4206,c0208,c0489,c719,c0133,c7249,c4171,c5397,c0155,c9237,c7286,c4463,c464,c8231,c3459,c6444,c7235,c1471,c4173,c8273,c3107,c5351,c7411,c4303,c5423,c4226,c3199,c8462,c0322,c1271,c0195,c2195,c4216,c0435,c1247,c2107,c5105,c5265,c7429,c5456,c7227,c9279,c8405,c7170,c9462,c3209,c2143,c3211,c959,c231,c5216,c5179,c3454,c1260,c8226,c6419,c7465,c0330,c811,c4124,c0368,c1426,c2435,c1225,c9444,c932,c7199,c1299,c4475,c6498,c6247,c2179,c3295,c5406,c569,c681,c0123,c3452,c51,c5446,c1407,c2335,c8140,c0104,c0348,c880,c1377,c5430,c3229,c297,c1402,c6275,c5489,c9129,c0481,c5190,c9381,c9324,c817,c2166,c9463,c4440,c5264,c579,c1172,c4433,c470,c5467,c0141,c1161,c7318,c9435,c972,c6339,c6202,c8117,c3115,c612,c8378,c614,c2145,c4345,c1265,c4135,c5111,c1153,c4314,c5229,c1267,c8243,c47,c6261,c7344,c582,c3312,c8385,c4133,c7183,c4478,c0377,c758,c6378,c860,c5268,c4191,c4112,c5403,c6136,c7214,c116,c521,c9208,c7180,c6454,c6453,c1326,c8331,c8132,c489,c01,c320,c5237,c3373,c2137,c9445,c9368,c0430,c7159,c2402,c6385,c2128,c3285,c3379,c282,c796,c5388,c8104,c2185,c6268,c8133,c275,c6237,c7263,c1137,c3235,c5292,c6197,c122,c488,c8126,c1217,c332,c9227,c8470,c157,c4294,c0196,c0211,c7184,c0236,c4168,c529,c5484,c4430,c8345,c9331,c5233,c467,c6486,c7299,c8377,c5356,c6148,c3145,c0194,c8162,c7151,c9408,c540,c0427,c4353,c54,c7194,c7292,c0205,c9409,c3431,c8180,c558,c39,c7100,c537,c975,c9115,c8391,c3491,c490,c0225,c5490,c6403,c2101,c7402,c8362,c6184,c8246,c5463,c2198,c9258,c086,c7379,c7339,c2345,c0319,c2306,c8191,c5415,c656,c5145,c3350,c593,c4315,c9389,c4444,c5267,c1200,c5201,c0109,c6484,c7217,c713,c4468,c8433,c95,c9179,c4241,c149,c72,c9461,c3334,c9245,c4497,c1452,c8499,c2446,c3292,c782,c8355,c6308,c620,c141,c1352,c3297,c5382,c696,c0382,c2159,c6457,c0118,c4222,c7476,c783,c9224,c9378,c256,c630,c1193,c730,c1388,c9470,c333,c1491,c349,c5209,c1495,c3195,c335,c8234,c2257,c2103,c1461,c4260,c3304,c979,c57,c3447,c6372,c1425,c9400,c9454,c2172,c3475,c6328,c6285,c2343,c4140,c4496,c7487,c5165,c5200,c8400,c7111,c4251,c7224,c8249,c1189,c3360,c2388,c2258,c2316,c3198,c2413,c0308,c4150,c4228,c5143,c4389,c9164,c0405,c6155,c664,c7458,c1298,c729,c5332,c5241,c1465,c0290,c5425,c6101,c7283,c4464,c2453,c6104,c9362,c5198,c3425,c949,c4364,c344,c5486,c5370,c1421,c622,c5116,c6305,c4248,c0267,c3226,c6478,c7414,c9112,c7131,c6460,c3170,c1192,c2136,c0464,c4413,c1281,c9297,c0347,c2146,c0209,c0410,c0261,c388,c6340,c6293,c7440,c724,c7289,c7296,c2475,c3423,c9220,c8454,c410,c639,c4432,c7348,c1397,c7396,c8392,c4105,c6395,c4446,c5108,c9391,c7352,c214,c7222,c4197,c3463,c687,c0395,c2204,c2149,c1320,c9221,c0390,c733,c1477,c5113,c356,c2183,c4240,c5342,c6338,c268,c7246,c6298,c8165,c4259,c8250,c6281,c2468,c6319,c6111,c2394,c468,c8256,c8115,c016,c5450,c7380,c528,c8150,c7374,c8267,c3171,c6359,c2181,c0406,c5287,c6230,c7287,c753,c2303,c0244,c12,c3442,c7420,c5375,c788,c1232,c7355,c4321,c525,c3359,c5386,c5315,c580,c893,c7349,c3383,c2397,c6485,c938,c5346,c9157,c13,c3104,c9122,c9219,c041,c4393,c0479,c210,c3200,c1378,c4154,c6271,c9344,c5466,c8293,c9102,c6239,c0494,c7426,c062,c923,c3275,c8413,c1376,c35,c2487,c0404,c3443,c1230,c366,c816,c6127,c821,c0401,c2482,c0431,c113,c1493,c7175,c261,c3133,c2450,c0374,c9397,c7354,c3121,c8374,c8416,c9398,c2157,c8284,c0143,c4379,c4134,c9426,c7437,c9442,c065,c2261,c3449,c5366,c590,c7316,c133,c4493,c5414,c9491,c7129,c221,c2148,c0472,c3165,c8287,c8351,c934,c0302,c6214,c1480,c9268,c7461,c1384,c0454,c8236,c553,c6488,c6435,c14,c2123,c8244,c2463,c0285,c6472,c8423,c2127,c0338,c4157,c211,c345,c8217,c0176,c0364,c3382,c8389,c0129,c5369,c7450,c5438,c052,c8229,c233,c481,c0441,c2144,c3263,c170,c2297,c9282,c757,c4338,c5350,c3143,c8107,c4111,c4358,c7135,c9328,c5214,c2287,c073,c1373,c8148,c1274,c0151,c479,c969,c595,c9162,c1263,c3409,c385,c8131,c3429,c1190,c9492,c6422,c9421,c4231,c7490,c6400,c8348,c37,c8473,c7252,c6463,c3301,c8353,c8482,c0335,c863,c4257,c7253,c6322,c891,c645,c8103,c9199,c3387,c5276,c4332,c6415,c3333,c2496,c7257,c2104,c4255,c3234,c045,c4236,c5309,c7262,c3286,c5399,c723,c6380,c2229,c742,c4362,c171,c3261,c743,c1295,c7282,c1364,c469,c6337,c5136,c797,c8177,c19,c9239,c2432,c7144,c599,c378,c076,c7223,c9267,c623,c8478,c8235,c2182,c013,c9289,c2290,c9364,c4254,c1221,c1145,c6287,c139,c9319,c3390,c4234,c0222,c9156,c430,c2365,c2307,c6224,c3428,c5158,c6151,c143,c239,c2423,c9308,c7155,c5262,c9284,c9406,c5259,c3362,c570,c7486,c0357,c1411,c576,c1337,c3177,c6262,c4434,c3493,c9116,c7156,c9296,c1306,c8424,c3488,c3408,c6437,c5163,c8196,c2238,c4320,c71,c0159,c8409,c2460,c1234,c6456,c538,c991,c4412,c0217,c859,c044,c418,c8163,c8290,c0228,c4274,c8147,c3103,c4117,c1350,c7256,c4196,c1438,c263,c3174,c9135,c2286,c9130,c027,c2298,c830,c0140,c5162,c1456,c1167,c6398,c3478,c8239,c8369,c5487,c121,c477,c1321,c7329,c2199,c7327,c4461,c892,c2132,c8379,c7497,c0183,c3345,c4230,c1132,c9287,c2255,c352,c4357,c6166,c7336,c4368,c7136,c5251,c9100,c8422,c4298,c4480,c567,c4237,c3406,c6220,c3277,c7114,c5184,c6232,c4290,c9183,c9251,c2184,c6428,c9488,c3483,c1227,c7381,c8407,c1164,c9361,c651,c6480,c1443,c5164,c011,c3223,c031,c9171,c759,c5340,c5166,c9424,c2396,c025,c3310,c2189,c7139,c4198,c2206,c924,c8328,c482,c9347,c7347,c8168,c0190,c1253,c8174,c6459,c9481,c277,c5409,c6192,c7491,c0397,c732,c3434,c6445,c4436,c6327,c965,c1382,c3271,c5245,c0240,c4392,c4180,c4457,c217,c633,c321,c3202,c3106,c4448,c5191,c7453,c2165,c4308,c951,c4194,c6323,c3417,c4341,c6421,c4305,c53,c1209,c1252,c8112,c961,c3196,c698,c3274,c0284,c997,c8207,c6276,c163,c0172,c5449,c3458,c396,c8261,c884,c2250,c7460,c9110,c565,c5240,c8105,c778,c0220,c9247,c2163,c4352,c4489,c852,c587,c5301,c1171,c8143,c531,c0380,c1118,c5273,c922,c9448,c1419,c993,c772,c0107,c5195,c9410,c722,c9394,c8397,c8188,c03,c5393,c4296,c9305,c197,c7163,c3318,c0483,c519,c4152,c2470,c842,c3276,c7382,c9288,c6321,c7209,c0203,c4273,c4333,c6117,c8125,c7300,c7397,c144,c0242,c6423,c3451,c8178,c6240,c4202,c7212,c4452,c7422,c8137,c9270,c9225,c5416,c4195,c1393,c3126,c1334,c3368,c0345,c6481,c9230,c2322,c1182,c8303,c4373,c5295,c5151,c4100,c7245,c9483,c9163,c9212,c1413,c5131,c059,c1381,c9320,c710,c0385,c3485,c3497,c5392,c1453,c3349,c1361,c75,c6376,c995,c7459,c7494,c160,c285,c4147,c6107,c720,c3456,c198,c73,c0381,c6144,c128,c9498,c4227,c7242,c5224,c6316,c1206,c0341,c3221,c8263,c6252,c8460,c0456,c642,c3157,c0449,c427,c3331,c5192,c9318,c2176,c5378,c1494,c311,c8299,c1310,c2362,c0433,c6128,c63,c0446,c8154,c6290,c1367,c1103,c9269,c3189,c5433,c3167,c2293,c5156,c7383,c4224,c5130,c8310,c0257,c3376,c4203,c226,c4347,c2459,c9211,c91,c6355,c7357,c222,c2464,c363,c6436,c652,c0232,c0384,c5345,c2155,c6153,c087,c4289,c5176,c6146,c4359,c1177,c2178,c442,c4439,c864,c41,c6198,c6143,c1467,c4390,c289,c2108,c4387,c6185,c2138,c8288,c7202,c0144,c1268,c8128,c589,c4225,c5401,c3194,c083,c0275,c1284,c8350,c1128,c3243,c7315,c781,c2152,c462,c1314,c644,c0340,c9342,c3249,c2117,c6309,c0476,c752,c0198,c0317,c6300,c2364,c2169,c6149,c9263,c2105,c6417,c5288,c6387,c0171,c9243,c6113,c1444,c8490,c8449,c8393,c0181,c2190,c0272,c3455,c539,c2168,c7387,c4139,c0417,c3227,c1116,c6404,c8195,c347,c6223,c981,c3153,c4467,c4474,c6315,c7158,c9309,c2489,c4415,c9357,c4310,c4249,c0221,c5307,c8248,c0413,c566,c3125,c976,c6433,c3110,c5495,c6496,c0108,c1395,c0412,c2422,c9159,c868,c5329,c435,c943,c7294,c5339,c6369,c8406,c0333,c7391,c0434,c4151,c581,c9226,c5278,c9302,c337,c7192,c2102,c370,c8430,c499,c7436,c5205,c8211,c398,c364,c3272,c257,c4377,c0276,c6414,c0294,c7229,c1346,c2332,c5291,c9431,c0428,c6491,c5281,c0288,c3283,c4337,c238,c3154,c574,c3146,c5352,c897,c7376,c647,c1105,c4429,c1332,c6292,c465,c8480,c136,c2382,c033,c5126,c0270,c6313,c9382,c0206,c776,c0366,c399,c0289,c1250,c518,c6412,c7190,c5132,c2180,c2110,c7498,c8373,c8218,c9422,c3220,c829,c3117,c0393,c4419,c8463,c0321,c5186,c3338,c223,c374,c3222,c974,c613,c2428,c126,c0246,c0468,c3342,c8152,c212,c929,c5338,c9255,c98,c1392,c7148,c0119,c5159,c3314,c324,c5355,c2350,c4425,c5349,c4103,c6258,c1479,c4317,c4156,c9111,c517,c0115,c6183,c4313,c1457,c293,c9373,c9418,c7356,c888,c3329,c7239,c46,c358,c7237,c9412,c7375,c6248,c6207,c1335,c377,c3156,c6303,c4163,c657,c714,c190,c2284,c9125,c7395,c3191,c7117,c9494,c7447,c2130,c0457,c147,c8412,c3152,c9332,c7285,c3489,c7312,c2439,c1124,c847,c0306,c7492,c0421,c8483,c0477,c7324,c3213,c1288,c2495,c7137,c037,c694,c7308,c3224,c4484,c5211,c6150,c7269,c9423,c0360,c487,c4351,c049,c1254,c6374,c5316,c7407,c5398,c511,c1451,c89,c2299,c1342,c0124,c5128,c575,c1436,c9228,c386,c8386,c1439,c2367,c2473,c188,c3109,c550,c1159,c2451,c3306,c120,c2270,c1148,c154,c5117,c2481,c2368,c3238,c5461,c6377,c9449,c3477,c0315,c9127,c3267,c242,c7451,c8472,c0396,c7361,c2414,c281,c4169,c5120,c1434,c0491,c4125,c1362,c8205,c2325,c6180,c7481,c6163,c064,c3180,c4149,c3420,c4471,c8402,c3399,c8339,c018,c6270,c9177,c885,c536,c476,c173,c06,c2122,c992,c7328,c8453,c5436,c615,c7191,c0166,c4307,c916,c869,c4271,c236,c1406,c2194,c9215,c8282,c6171,c1365,c843,c9206,c5474,c2125,c5460,c1146,c6461,c0490,c5493,c5125,c3444,c249,c9490,c328,c2395,c7332,c9300,c9293,c3343,c5390,c6100,c7132,c5472,c9184,c0135,c8376,c9325,c44,c4304,c5230,c2406,c728,c1222,c1123,c284,c6178,c9414,c2164,c2353,c0329,c3341,c3175,c655,c0160,c2426,c1149,c9114,c0281,c437,c5442,c7126,c6129,c2161,c092,c9472,c1371,c350,c3105,c8344,c6440,c1241,c9487,c6255,c0337,c4322,c2312,c0358,c2321,c5260,c179,c7434,c4470,c9271,c8494,c4473,c0305,c4131,c9261,c3499,c7244,c1279,c6159,c957,c270,c0459,c1138,c983,c9303,c3260,c4166,c9482,c3495,c9374,c799,c130,c125,c7204,c6302,c8308,c6416,c7293,c3176,c854,c4108,c9192,c7326,c9473,c3258,c8281,c8139,c5499,c9236,c516,c5183,c6231,c4330,c0165,c448,c4424,c1404,c6282,c361,c379,c9218,c0260,c8266,c83,c865,c6495,c9153,c2461,c4291,c1158,c7480,c2232,c5322,c2301,c4137,c3450,c6336,c391,c964,c392,c030,c522,c5384,c6132,c2113,c8260,c3203,c74,c1341,c621,c0312,c2486,c2167,c7441,c5127,c5118,c7433,c6288,c1490,c327,c0152,c5475,c3336,c588,c6133,c9148,c6272,c6476,c0426,c9246,c7127,c0485,c066,c6279,c5178,c5379,c5160,c5254,c097,c4449,c6388,c5437,c0478,c3320,c6212,c8304,c563,c9457,c1405,c0191,c3186,c5334,c383,c322,c8395,c9124,c084,c846,c0273,c948,c1440,c8106,c996,c0157,c2447,c8437,c9169,c439,c245,c8436,c8270,c7398,c79,c2230,c8258,c5139,c6115,c8138,c3256,c0150,c5395,c8352,c5304,c941,c2398,c7448,c2246,c9495,c583,c6225,c1202,c3173,c118,c2313,c3347,c7203,c7305,c3245,c7251,c2114,c735,c9213,c2239,c9154,c3147,c046,c6235,c5243,c3251,c873,c9232,c1152,c7297,c59,c6126,c7160,c0325,c1102,c571,c3300,c7463,c1359,c2126,c6162,c3140,c8488,c5317,c1446,c833,c129,c0495,c2373,c7106,c5331,c9349,c4465,c4145,c9429,c5303,c7389,c831,c9185,c6342,c4279,c3438,c4416,c9420,c2479,c832,c3465,c70,c1294,c2356,c8279,c7377,c6405,c2240,c4215,c0486,c5208,c2471,c1416,c3363,c3187,c7113,c6489,c325,c5453,c597,c5408,c5427,c5373,c1156,c2295,c1369,c8435,c8176,c5318,c2282,c3281,c3216,c6464,c4409,c9388,c1109,c1239,c624,c4309,c9443,c3164,c354,c85,c8451,c2162,c145,c9366,c9133,c5360,c6325,c935,c557,c9160,c7260,c6473,c6203,c697,c919,c2237,c8285,c3366,c3492,c4136,c6102,c6234,c9103,c726,c7140,c7388,c1499,c00,c0256,c5226,c0297,c5485,c7423,c9186,c7219,c5167,c8468,c298,c6165,c7238,c1464,c0112,c5283,c5275,c1184,c3400,c2441,c998,c2263,c617,c886,c4451,c368,c0331,c2173,c0262,c1325,c6187,c7403,c653,c9312,c1396,c9147,c5469,c316,c2385,c9278,c7400,c3325,c1481,c0188,c9434,c3357,c7218,c1460,c5231,c9419,c4370,c8312,c6420,c9146 );

input x0;
input x1;
input x2;
input x3;
input x4;
input x5;
input x6;
input x7;
input x8;
input x9;
input x10;
input x11;
input x12;
input x13;
input x14;
input x15;
input x16;
input x17;
input x18;
input x19;
input x20;
input x21;
input x22;
input x23;
input x24;
input x25;
input x26;
input x27;
input x28;
input x29;
input x30;
input x31;
input x32;
input x33;
input x34;
input x35;
input x36;
input x37;
input x38;
input x39;
input x40;
input x41;
input x42;
input x43;
input x44;
input x45;
input x46;
input x47;
input x48;
input x49;
input x50;
input x51;
input x52;
input x53;
input x54;
input x55;
input x56;
input x57;
input x58;
input x59;
input x60;
input x61;
input x62;
input x63;
input x64;
input x65;
input x66;
input x67;
input x68;
input x69;
input x70;
input x71;
input x72;
input x73;
input x74;
input x75;
input x76;
input x77;
input x78;
input x79;
input x80;
input x81;
input x82;
input x83;
input x84;
input x85;
input x86;
input x87;
input x88;
input x89;
input x90;
input x91;
input x92;
input x93;
input x94;
input x95;
input x96;
input x97;
input x98;
input x99;
input x100;
input x101;
input x102;
input x103;
input x104;
input x105;
input x106;
input x107;
input x108;
input x109;
input x110;
input x111;
input x112;
input x113;
input x114;
input x115;
input x116;
input x117;
input x118;
input x119;
input x120;
input x121;
input x122;
input x123;
input x124;
input x125;
input x126;
input x127;
input x128;
input x129;
input x130;
input x131;
input x132;
input x133;
input x134;
input x135;
input x136;
input x137;
input x138;
input x139;
input x140;
input x141;
input x142;
input x143;
input x144;
input x145;
input x146;
input x147;
input x148;
input x149;
input x150;
input x151;
input x152;
input x153;
input x154;
input x155;
input x156;
input x157;
input x158;
input x159;
input x160;
input x161;
input x162;
input x163;
input x164;
input x165;
input x166;
input x167;
input x168;
input x169;
input x170;
input x171;
input x172;
input x173;
input x174;
input x175;
input x176;
input x177;
input x178;
input x179;
input x180;
input x181;
input x182;
input x183;
input x184;
input x185;
input x186;
input x187;
input x188;
input x189;
input x190;
input x191;
input x192;
input x193;
input x194;
input x195;
input x196;
input x197;
input x198;
input x199;
input x200;
input x201;
input x202;
input x203;
input x204;
input x205;
input x206;
input x207;
input x208;
input x209;
input x210;
input x211;
input x212;
input x213;
input x214;
input x215;
input x216;
input x217;
input x218;
input x219;
input x220;
input x221;
input x222;
input x223;
input x224;
input x225;
input x226;
input x227;
input x228;
input x229;
input x230;
input x231;
input x232;
input x233;
input x234;
input x235;
input x236;
input x237;
input x238;
input x239;
input x240;
input x241;
input x242;
input x243;
input x244;
input x245;
input x246;
input x247;
input x248;
input x249;
input x250;
input x251;
input x252;
input x253;
input x254;
input x255;
input x256;
input x257;
input x258;
input x259;
input x260;
input x261;
input x262;
input x263;
input x264;
input x265;
input x266;
input x267;
input x268;
input x269;
input x270;
input x271;
input x272;
input x273;
input x274;
input x275;
input x276;
input x277;
input x278;
input x279;
input x280;
input x281;
input x282;
input x283;
input x284;
input x285;
input x286;
input x287;
input x288;
input x289;
input x290;
input x291;
input x292;
input x293;
input x294;
input x295;
input x296;
input x297;
input x298;
input x299;
input x300;
input x301;
input x302;
input x303;
input x304;
input x305;
input x306;
input x307;
input x308;
input x309;
input x310;
input x311;
input x312;
input x313;
input x314;
input x315;
input x316;
input x317;
input x318;
input x319;
input x320;
input x321;
input x322;
input x323;
input x324;
input x325;
input x326;
input x327;
input x328;
input x329;
input x330;
input x331;
input x332;
input x333;
input x334;
input x335;
input x336;
input x337;
input x338;
input x339;
input x340;
input x341;
input x342;
input x343;
input x344;
input x345;
input x346;
input x347;
input x348;
input x349;
input x350;
input x351;
input x352;
input x353;
input x354;
input x355;
input x356;
input x357;
input x358;
input x359;
input x360;
input x361;
input x362;
input x363;
input x364;
input x365;
input x366;
input x367;
input x368;
input x369;
input x370;
input x371;
input x372;
input x373;
input x374;
input x375;
input x376;
input x377;
input x378;
input x379;
input x380;
input x381;
input x382;
input x383;
input x384;
input x385;
input x386;
input x387;
input x388;
input x389;
input x390;
input x391;
input x392;
input x393;
input x394;
input x395;
input x396;
input x397;
input x398;
input x399;
input x400;
input x401;
input x402;
input x403;
input x404;
input x405;
input x406;
input x407;
input x408;
input x409;
input x410;
input x411;
input x412;
input x413;
input x414;
input x415;
input x416;
input x417;
input x418;
input x419;
input x420;
input x421;
input x422;
input x423;
input x424;
input x425;
input x426;
input x427;
input x428;
input x429;
input x430;
input x431;
input x432;
input x433;
input x434;
input x435;
input x436;
input x437;
input x438;
input x439;
input x440;
input x441;
input x442;
input x443;
input x444;
input x445;
input x446;
input x447;
input x448;
input x449;
input x450;
input x451;
input x452;
input x453;
input x454;
input x455;
input x456;
input x457;
input x458;
input x459;
input x460;
input x461;
input x462;
input x463;
input x464;
input x465;
input x466;
input x467;
input x468;
input x469;
input x470;
input x471;
input x472;
input x473;
input x474;
input x475;
input x476;
input x477;
input x478;
input x479;
input x480;
input x481;
input x482;
input x483;
input x484;
input x485;
input x486;
input x487;
input x488;
input x489;
input x490;
input x491;
input x492;
input x493;
input x494;
input x495;
input x496;
input x497;
input x498;
input x499;
input x500;
input x501;
input x502;
input x503;
input x504;
input x505;
input x506;
input x507;
input x508;
input x509;
input x510;
input x511;
input x512;
input x513;
input x514;
input x515;
input x516;
input x517;
input x518;
input x519;
input x520;
input x521;
input x522;
input x523;
input x524;
input x525;
input x526;
input x527;
input x528;
input x529;
input x530;
input x531;
input x532;
input x533;
input x534;
input x535;
input x536;
input x537;
input x538;
input x539;
input x540;
input x541;
input x542;
input x543;
input x544;
input x545;
input x546;
input x547;
input x548;
input x549;
input x550;
input x551;
input x552;
input x553;
input x554;
input x555;
input x556;
input x557;
input x558;
input x559;
input x560;
input x561;
input x562;
input x563;
input x564;
input x565;
input x566;
input x567;
input x568;
input x569;
input x570;
input x571;
input x572;
input x573;
input x574;
input x575;
input x576;
input x577;
input x578;
input x579;
input x580;
input x581;
input x582;
input x583;
input x584;
input x585;
input x586;
input x587;
input x588;
input x589;
input x590;
input x591;
input x592;
input x593;
input x594;
input x595;
input x596;
input x597;
input x598;
input x599;
input x600;
input x601;
input x602;
input x603;
input x604;
input x605;
input x606;
input x607;
input x608;
input x609;
input x610;
input x611;
input x612;
input x613;
input x614;
input x615;
input x616;
input x617;
input x618;
input x619;
input x620;
input x621;
input x622;
input x623;
input x624;
input x625;
input x626;
input x627;
input x628;
input x629;
input x630;
input x631;
input x632;
input x633;
input x634;
input x635;
input x636;
input x637;
input x638;
input x639;
input x640;
input x641;
input x642;
input x643;
input x644;
input x645;
input x646;
input x647;
input x648;
input x649;
input x650;
input x651;
input x652;
input x653;
input x654;
input x655;
input x656;
input x657;
input x658;
input x659;
input x660;
input x661;
input x662;
input x663;
input x664;
input x665;
input x666;
input x667;
input x668;
input x669;
input x670;
input x671;
input x672;
input x673;
input x674;
input x675;
input x676;
input x677;
input x678;
input x679;
input x680;
input x681;
input x682;
input x683;
input x684;
input x685;
input x686;
input x687;
input x688;
input x689;
input x690;
input x691;
input x692;
input x693;
input x694;
input x695;
input x696;
input x697;
input x698;
input x699;
input x700;
input x701;
input x702;
input x703;
input x704;
input x705;
input x706;
input x707;
input x708;
input x709;
input x710;
input x711;
input x712;
input x713;
input x714;
input x715;
input x716;
input x717;
input x718;
input x719;
input x720;
input x721;
input x722;
input x723;
input x724;
input x725;
input x726;
input x727;
input x728;
input x729;
input x730;
input x731;
input x732;
input x733;
input x734;
input x735;
input x736;
input x737;
input x738;
input x739;
input x740;
input x741;
input x742;
input x743;
input x744;
input x745;
input x746;
input x747;
input x748;
input x749;
input x750;
input x751;
input x752;
input x753;
input x754;
input x755;
input x756;
input x757;
input x758;
input x759;
input x760;
input x761;
input x762;
input x763;
input x764;
input x765;
input x766;
input x767;
input x768;
input x769;
input x770;
input x771;
input x772;
input x773;
input x774;
input x775;
input x776;
input x777;
input x778;
input x779;
input x780;
input x781;
input x782;
input x783;
output c8238;
output c7311;
output c2224;
output c3391;
output c0356;
output c0309;
output c8324;
output c1433;
output c447;
output c594;
output c1176;
output c6238;
output c5458;
output c1360;
output c4293;
output c6236;
output c3480;
output c5353;
output c4243;
output c1154;
output c090;
output c0280;
output c7271;
output c625;
output c4371;
output c5488;
output c7259;
output c3355;
output c4200;
output c1355;
output c898;
output c5429;
output c7243;
output c2112;
output c2430;
output c8216;
output c155;
output c4435;
output c2171;
output c882;
output c5365;
output c5424;
output c661;
output c4483;
output c6335;
output c2218;
output c2358;
output c7372;
output c3298;
output c1349;
output c8370;
output c2275;
output c151;
output c2370;
output c7153;
output c6306;
output c1292;
output c7401;
output c872;
output c5284;
output c252;
output c813;
output c921;
output c3135;
output c6135;
output c2272;
output c4185;
output c6466;
output c5478;
output c0131;
output c5371;
output c672;
output c11;
output c3130;
output c0460;
output c6499;
output c5173;
output c643;
output c6221;
output c248;
output c4460;
output c2292;
output c6256;
output c4201;
output c7220;
output c4120;
output c6284;
output c1114;
output c3468;
output c958;
output c1243;
output c4378;
output c3166;
output c7232;
output c4142;
output c674;
output c1208;
output c9363;
output c7430;
output c4158;
output c111;
output c8414;
output c3487;
output c7446;
output c050;
output c6384;
output c1256;
output c2242;
output c33;
output c054;
output c0298;
output c5491;
output c878;
output c438;
output c56;
output c6333;
output c982;
output c7161;
output c17;
output c1417;
output c8108;
output c837;
output c2300;
output c9456;
output c174;
output c3435;
output c8346;
output c526;
output c152;
output c0193;
output c6259;
output c4324;
output c9264;
output c3296;
output c0187;
output c7280;
output c8301;
output c6383;
output c9432;
output c1340;
output c5402;
output c4487;
output c3206;
output c9339;
output c310;
output c2201;
output c4242;
output c6242;
output c5431;
output c7484;
output c8356;
output c6409;
output c02;
output c9202;
output c2193;
output c9197;
output c2438;
output c8343;
output c9468;
output c8368;
output c5418;
output c8189;
output c8469;
output c3280;
output c0117;
output c4325;
output c5169;
output c5280;
output c074;
output c1211;
output c4181;
output c0304;
output c4427;
output c436;
output c191;
output c8265;
output c9379;
output c6397;
output c1363;
output c4348;
output c4179;
output c845;
output c2197;
output c9480;
output c5253;
output c9109;
output c1437;
output c6245;
output c3100;
output c942;
output c824;
output c6125;
output c8194;
output c8450;
output c8338;
output c1139;
output c8418;
output c38;
output c4245;
output c947;
output c541;
output c158;
output c265;
output c2221;
output c8197;
output c082;
output c2226;
output c3378;
output c8458;
output c4277;
output c0328;
output c6477;
output c2348;
output c4123;
output c4394;
output c3445;
output c3372;
output c1315;
output c6427;
output c4192;
output c9252;
output c9326;
output c6181;
output c8135;
output c7276;
output c5413;
output c9453;
output c2154;
output c0282;
output c3241;
output c6295;
output c6382;
output c2410;
output c4270;
output c0237;
output c232;
output c2465;
output c4381;
output c127;
output c150;
output c7371;
output c4233;
output c855;
output c1431;
output c3218;
output c1248;
output c2375;
output c1117;
output c6280;
output c8495;
output c573;
output c3396;
output c2158;
output c172;
output c0105;
output c4311;
output c2334;
output c2160;
output c678;
output c010;
output c8272;
output c6195;
output c2376;
output c8396;
output c5468;
output c67;
output c4391;
output c1104;
output c0299;
output c6344;
output c0224;
output c8127;
output c2346;
output c715;
output c660;
output c0429;
output c721;
output c2170;
output c9274;
output c312;
output c9455;
output c5140;
output c7149;
output c1423;
output c3427;
output c3335;
output c3244;
output c3348;
output c6141;
output c8257;
output c2283;
output c7469;
output c3159;
output c0386;
output c7164;
output c7320;
output c4109;
output c3179;
output c0235;
output c767;
output c5144;
output c6334;
output c4498;
output c0301;
output c2212;
output c9140;
output c544;
output c3326;
output c348;
output c7154;
output c474;
output c475;
output c2187;
output c341;
output c7369;
output c1409;
output c6229;
output c6170;
output c82;
output c5354;
output c9411;
output c365;
output c5302;
output c9142;
output c2259;
output c812;
output c3327;
output c5441;
output c3395;
output c463;
output c945;
output c2342;
output c2174;
output c0365;
output c5374;
output c94;
output c9174;
output c0389;
output c9131;
output c6365;
output c2281;
output c7303;
output c6289;
output c273;
output c9106;
output c1199;
output c7270;
output c8274;
output c4269;
output c7112;
output c3461;
output c6278;
output c1322;
output c0121;
output c7464;
output c673;
output c0170;
output c5333;
output c3421;
output c2387;
output c026;
output c4218;
output c5480;
output c230;
output c546;
output c584;
output c913;
output c7162;
output c6310;
output c1257;
output c3137;
output c6401;
output c3369;
output c9180;
output c3278;
output c0422;
output c6122;
output c1399;
output c0234;
output c2449;
output c6426;
output c6343;
output c2109;
output c6468;
output c6193;
output c169;
output c1412;
output c3132;
output c7101;
output c944;
output c9436;
output c1185;
output c520;
output c5124;
output c2326;
output c0379;
output c9290;
output c640;
output c3172;
output c8134;
output c765;
output c8440;
output c1454;
output c7425;
output c3129;
output c7116;
output c554;
output c598;
output c8276;
output c8145;
output c7221;
output c373;
output c4207;
output c5182;
output c3410;
output c1387;
output c4261;
output c123;
output c124;
output c2111;
output c069;
output c292;
output c1375;
output c677;
output c4300;
output c5330;
output c7485;
output c2217;
output c3307;
output c7419;
output c1283;
output c5394;
output c4428;
output c5219;
output c4422;
output c578;
output c3371;
output c4276;
output c4376;
output c1175;
output c3367;
output c6451;
output c828;
output c0362;
output c1233;
output c1195;
output c4164;
output c5421;
output c750;
output c5249;
output c9428;
output c926;
output c9417;
output c3401;
output c5203;
output c9120;
output c2405;
output c8120;
output c453;
output c6173;
output c4363;
output c0452;
output c8220;
output c5324;
output c8410;
output c6430;
output c8123;
output c0263;
output c1366;
output c5148;
output c2440;
output c8192;
output c9145;
output c0394;
output c3323;
output c4336;
output c1448;
output c0339;
output c5289;
output c2454;
output c2310;
output c8153;
output c1462;
output c6434;
output c5412;
output c7121;
output c2118;
output c148;
output c1141;
output c494;
output c5447;
output c3476;
output c0238;
output c0122;
output c973;
output c8404;
output c2391;
output c9205;
output c4190;
output c9403;
output c9254;
output c1266;
output c8481;
output c9158;
output c9136;
output c857;
output c3162;
output c8201;
output c5114;
output c1328;
output c9380;
output c166;
output c4256;
output c8491;
output c994;
output c6108;
output c330;
output c4306;
output c0127;
output c0376;
output c6304;
output c5137;
output c636;
output c3169;
output c6227;
output c7340;
output c7314;
output c55;
output c6348;
output c2386;
output c2280;
output c8184;
output c5361;
output c071;
output c2403;
output c6439;
output c4331;
output c2196;
output c5296;
output c189;
output c2361;
output c2415;
output c6157;
output c8371;
output c9209;
output c4284;
output c161;
output c2455;
output c0189;
output c4301;
output c371;
output c1100;
output c798;
output c7454;
output c8333;
output c8222;
output c889;
output c255;
output c9165;
output c4113;
output c4401;
output c6201;
output c1472;
output c9222;
output c5464;
output c0442;
output c4267;
output c7102;
output c6241;
output c1142;
output c626;
output c5310;
output c0164;
output c560;
output c0323;
output c0271;
output c6407;
output c449;
output c0307;
output c632;
output c1113;
output c2336;
output c5244;
output c7200;
output c9152;
output c2175;
output c088;
output c0229;
output c2211;
output c5428;
output c2227;
output c326;
output c5107;
output c962;
output c2228;
output c1353;
output c3418;
output c7412;
output c4161;
output c2324;
output c99;
output c8116;
output c760;
output c9425;
output c2425;
output c2417;
output c76;
output c42;
output c3309;
output c5462;
output c9128;
output c4356;
output c156;
output c496;
output c9334;
output c8330;
output c5479;
output c1204;
output c0286;
output c0120;
output c7323;
output c911;
output c8292;
output c3158;
output c0216;
output c2492;
output c5454;
output c421;
output c2349;
output c3358;
output c4407;
output c9323;
output c6474;
output c8415;
output c3328;
output c545;
output c4316;
output c0126;
output c9465;
output c028;
output c1258;
output c1157;
output c6375;
output c417;
output c1441;
output c9329;
output c1183;
output c491;
output c0269;
output c7302;
output c6381;
output c6161;
output c1140;
output c5298;
output c0469;
output c793;
output c740;
output c359;
output c610;
output c492;
output c5294;
output c290;
output c5326;
output c7351;
output c826;
output c286;
output c8428;
output c6286;
output c4477;
output c9198;
output c9275;
output c5134;
output c9451;
output c2433;
output c8334;
output c1476;
output c3313;
output c1226;
output c3190;
output c7130;
output c3469;
output c2318;
output c185;
output c2265;
output c2305;
output c3282;
output c8471;
output c5383;
output c6362;
output c1498;
output c5443;
output c8214;
output c8365;
output c6312;
output c5337;
output c1249;
output c1273;
output c1300;
output c5452;
output c4388;
output c2467;
output c680;
output c1488;
output c4297;
output c32;
output c9315;
output c411;
output c7228;
output c7409;
output c4280;
output c1302;
output c7189;
output c1336;
output c3250;
output c0268;
output c8489;
output c5279;
output c7181;
output c4247;
output c1390;
output c8305;
output c0487;
output c194;
output c3446;
output c0156;
output c1389;
output c8420;
output c4328;
output c1215;
output c3433;
output c7240;
output c747;
output c8316;
output c4167;
output c3155;
output c1136;
output c1445;
output c7146;
output c5494;
output c774;
output c8455;
output c4104;
output c2289;
output c1484;
output c8223;
output c5293;
output c8164;
output c953;
output c9195;
output c2140;
output c0161;
output c7295;
output c1324;
output c8209;
output c6494;
output c7173;
output c3204;
output c3214;
output c4106;
output c8364;
output c8466;
output c1430;
output c241;
output c7207;
output c1259;
output c055;
output c0132;
output c5196;
output c693;
output c3340;
output c5271;
output c0311;
output c2252;
output c3268;
output c3473;
output c5256;
output c2115;
output c6366;
output c815;
output c7444;
output c3160;
output c7234;
output c0142;
output c7266;
output c3294;
output c2341;
output c9291;
output c8255;
output c8213;
output c6103;
output c7174;
output c1466;
output c1343;
output c8297;
output c3163;
output c9235;
output c6274;
output c3337;
output c8394;
output c051;
output c7157;
output c3411;
output c6352;
output c8230;
output c5269;
output c9313;
output c6449;
output c1331;
output c1110;
output c6353;
output c458;
output c0145;
output c716;
output c7187;
output c818;
output c1285;
output c1339;
output c5103;
output c451;
output c454;
output c8319;
output c8434;
output c2328;
output c5372;
output c3212;
output c97;
output c0230;
output c4423;
output c7134;
output c8186;
output c1486;
output c2119;
output c6483;
output c2452;
output c8403;
output c6452;
output c6443;
output c2245;
output c8101;
output c434;
output c823;
output c5328;
output c2393;
output c685;
output c6249;
output c0239;
output c6124;
output c3108;
output c9104;
output c8487;
output c3393;
output c6296;
output c7337;
output c6140;
output c0212;
output c0147;
output c66;
output c9385;
output c8438;
output c3128;
output c7279;
output c038;
output c4220;
output c7452;
output c7145;
output c9317;
output c8448;
output c9439;
output c791;
output c4319;
output c5387;
output c072;
output c1229;
output c1293;
output c0139;
output c5455;
output c861;
output c9194;
output c0439;
output c90;
output c4229;
output c3414;
output c5235;
output c5432;
output c1106;
output c7325;
output c6217;
output c162;
output c3426;
output c3439;
output c323;
output c4114;
output c5175;
output c937;
output c4495;
output c9355;
output c8485;
output c8332;
output c5396;
output c1213;
output c4272;
output c8309;
output c6291;
output c3248;
output c9210;
output c8149;
output c2389;
output c441;
output c4490;
output c6169;
output c4160;
output c0138;
output c382;
output c2472;
output c4406;
output c6264;
output c6413;
output c5282;
output c1179;
output c1133;
output c2478;
output c8401;
output c05;
output c7290;
output c5180;
output c0162;
output c7439;
output c3114;
output c7109;
output c4469;
output c0134;
output c999;
output c426;
output c7343;
output c2277;
output c9207;
output c7250;
output c7477;
output c5277;
output c2264;
output c6402;
output c7427;
output c240;
output c5135;
output c836;
output c029;
output c1449;
output c3432;
output c7410;
output c8185;
output c0283;
output c8442;
output c8203;
output c0450;
output c0399;
output c4443;
output c9191;
output c1305;
output c6301;
output c5187;
output c9306;
output c6408;
output c4399;
output c043;
output c3290;
output c650;
output c1290;
output c4408;
output c8315;
output c4214;
output c4492;
output c5236;
output c1304;
output c7471;
output c9259;
output c4365;
output c954;
output c6204;
output c2404;
output c5286;
output c2262;
output c779;
output c5313;
output c274;
output c4188;
output c1414;
output c3255;
output c1210;
output c2434;
output c5498;
output c2241;
output c4400;
output c2480;
output c2458;
output c4126;
output c3381;
output c3403;
output c1319;
output c8241;
output c135;
output c8114;
output c5314;
output c1272;
output c5445;
output c874;
output c7291;
output c9437;
output c2457;
output c5217;
output c6471;
output c777;
output c4159;
output c497;
output c4395;
output c023;
output c4102;
output c1307;
output c9260;
output c079;
output c5362;
output c4380;
output c8329;
output c61;
output c9310;
output c6487;
output c631;
output c7176;
output c036;
output c7330;
output c1144;
output c3201;
output c138;
output c4402;
output c9107;
output c9249;
output c8247;
output c2355;
output c1357;
output c5411;
output c8175;
output c5426;
output c2339;
output c2491;
output c299;
output c280;
output c555;
output c0419;
output c2340;
output c048;
output c629;
output c0418;
output c532;
output c357;
output c6233;
output c8493;
output c0318;
output c6438;
output c3161;
output c0409;
output c015;
output c4144;
output c676;
output c134;
output c3232;
output c0295;
output c2219;
output c0293;
output c0314;
output c5246;
output c1458;
output c1201;
output c1291;
output c9175;
output c0378;
output c4398;
output c1347;
output c9253;
output c1244;
output c3270;
output c618;
output c4235;
output c3247;
output c5204;
output c7432;
output c0326;
output c80;
output c7208;
output c3123;
output c4491;
output c7193;
output c0416;
output c1497;
output c4292;
output c4128;
output c9188;
output c9467;
output c0359;
output c785;
output c0233;
output c912;
output c662;
output c0231;
output c8100;
output c0471;
output c7496;
output c5482;
output c3291;
output c3287;
output c0173;
output c4252;
output c7365;
output c6196;
output c7479;
output c098;
output c9176;
output c8179;
output c4372;
output c9123;
output c9256;
output c8398;
output c2347;
output c8360;
output c8113;
output c26;
output c792;
output c4318;
output c8441;
output c5391;
output c2151;
output c0372;
output c9189;
output c7195;
output c8181;
output c4479;
output c2448;
output c1162;
output c219;
output c1489;
output c078;
output c7177;
output c0265;
output c8421;
output c2150;
output c192;
output c0168;
output c3302;
output c7186;
output c3279;
output c3138;
output c8300;
output c6254;
output c360;
output c1469;
output c7169;
output c6493;
output c3380;
output c9459;
output c784;
output c2205;
output c3219;
output c259;
output c8278;
output c968;
output c7206;
output c3322;
output c6360;
output c485;
output c0243;
output c8363;
output c9200;
output c7499;
output c963;
output c0259;
output c440;
output c5177;
output c4411;
output c659;
output c1228;
output c7281;
output c227;
output c2304;
output c7442;
output c0249;
output c5146;
output c1187;
output c5250;
output c4101;
output c5473;
output c887;
output c5202;
output c62;
output c159;
output c1327;
output c1483;
output c4335;
output c9489;
output c695;
output c4121;
output c2311;
output c3120;
output c095;
output c3240;
output c649;
output c4143;
output c461;
output c375;
output c1317;
output c334;
output c745;
output c8411;
output c4458;
output c2279;
output c1169;
output c3472;
output c3168;
output c1391;
output c910;
output c6320;
output c628;
output c424;
output c2251;
output c2314;
output c2141;
output c0346;
output c69;
output c3448;
output c3254;
output c413;
output c2236;
output c1278;
output c267;
output c4386;
output c9354;
output c6479;
output c1194;
output c9134;
output c0488;
output c2412;
output c6226;
output c8166;
output c5106;
output c9150;
output c140;
output c4278;
output c8497;
output c420;
output c032;
output c667;
output c0458;
output c2294;
output c3239;
output c3178;
output c07;
output c6482;
output c559;
output c9450;
output c0186;
output c2497;
output c1383;
output c0101;
output c9217;
output c7133;
output c2401;
output c2416;
output c1107;
output c627;
output c1218;
output c0375;
output c0447;
output c3273;
output c825;
output c4141;
output c0445;
output c1212;
output c780;
output c8242;
output c7141;
output c92;
output c8124;
output c9257;
output c9345;
output c764;
output c4184;
output c918;
output c9416;
output c2315;
output c2223;
output c5306;
output c5380;
output c167;
output c4354;
output c429;
output c5435;
output c2469;
output c60;
output c6172;
output c7418;
output c9356;
output c3467;
output c543;
output c5194;
output c247;
output c6458;
output c343;
output c6210;
output c4414;
output c24;
output c7236;
output c5168;
output c8349;
output c7472;
output c6441;
output c5232;
output c49;
output c9105;
output c1186;
output c0251;
output c6191;
output c2129;
output c4263;
output c9283;
output c2490;
output c1372;
output c3269;
output c2424;
output c1270;
output c5496;
output c0264;
output c6142;
output c534;
output c8159;
output c3375;
output c040;
output c1282;
output c2200;
output c8492;
output c45;
output c0400;
output c5319;
output c665;
output c5228;
output c3289;
output c3419;
output c8144;
output c9204;
output c0148;
output c6123;
output c3127;
output c1122;
output c362;
output c2384;
output c099;
output c5410;
output c28;
output c9299;
output c216;
output c1173;
output c40;
output c067;
output c3231;
output c790;
output c0114;
output c5405;
output c5419;
output c0197;
output c950;
output c0440;
output c9314;
output c077;
output c8252;
output c6368;
output c3141;
output c6455;
output c36;
output c8399;
output c0177;
output c6246;
output c8187;
output c4118;
output c0451;
output c1224;
output c446;
output c085;
output c2488;
output c638;
output c3385;
output c585;
output c8169;
output c177;
output c09;
output c8382;
output c0130;
output c4177;
output c0167;
output c498;
output c1150;
output c094;
output c2456;
output c7213;
output c9384;
output c372;
output c768;
output c34;
output c024;
output c25;
output c2186;
output c9117;
output c4205;
output c7408;
output c7455;
output c1180;
output c875;
output c5312;
output c0402;
output c0437;
output c48;
output c8167;
output c1214;
output c7275;
output c8240;
output c9401;
output c2317;
output c564;
output c0158;
output c853;
output c8425;
output c8476;
output c4339;
output c2431;
output c8224;
output c3305;
output c0383;
output c8484;
output c646;
output c457;
output c4239;
output c8172;
output c9348;
output c0462;
output c52;
output c7483;
output c712;
output c849;
output c766;
output c7128;
output c514;
output c2216;
output c021;
output c3466;
output c8110;
output c3402;
output c7445;
output c8443;
output c0414;
output c260;
output c851;
output c635;
output c246;
output c0492;
output c1358;
output c4396;
output c6341;
output c2266;
output c2498;
output c7197;
output c8325;
output c3321;
output c3453;
output c838;
output c3424;
output c7284;
output c2409;
output c841;
output c8464;
output c1312;
output c896;
output c3482;
output c0496;
output c8161;
output c1130;
output c093;
output c3389;
output c985;
output c7470;
output c7350;
output c9155;
output c3237;
output c0215;
output c4285;
output c0102;
output c6418;
output c562;
output c9161;
output c0473;
output c5185;
output c9182;
output c2466;
output c940;
output c23;
output c7241;
output c9292;
output c31;
output c7367;
output c178;
output c5170;
output c4148;
output c734;
output c0455;
output c6116;
output c4127;
output c9132;
output c7272;
output c7406;
output c1111;
output c5363;
output c9469;
output c483;
output c4367;
output c2192;
output c3374;
output c9273;
output c4384;
output c2437;
output c5297;
output c675;
output c288;
output c9172;
output c4456;
output c7482;
output c990;
output c9479;
output c9298;
output c7185;
output c535;
output c9476;
output c8447;
output c4397;
output c381;
output c2330;
output c9496;
output c0223;
output c6118;
output c2214;
output c4204;
output c3324;
output c5122;
output c0332;
output c9387;
output c3494;
output c9272;
output c4221;
output c6194;
output c276;
output c8477;
output c9393;
output c4232;
output c5255;
output c0334;
output c0116;
output c3242;
output c523;
output c060;
output c21;
output c1475;
output c9395;
output c6361;
output c1216;
output c3266;
output c5497;
output c669;
output c0103;
output c7288;
output c5440;
output c8251;
output c5223;
output c8452;
output c9446;
output c5199;
output c1286;
output c4466;
output c0274;
output c2156;
output c7215;
output c8208;
output c7385;
output c0354;
output c8146;
output c1368;
output c744;
output c1235;
output c2177;
output c746;
output c2207;
output c5492;
output c691;
output c756;
output c7120;
output c9143;
output c380;
output c8367;
output c3346;
output c9285;
output c0465;
output c199;
output c3471;
output c053;
output c5207;
output c9466;
output c2383;
output c5477;
output c8467;
output c0349;
output c8171;
output c1261;
output c2208;
output c262;
output c8381;
output c8277;
output c186;
output c1496;
output c0371;
output c9386;
output c2378;
output c7322;
output c4299;
output c738;
output c915;
output c7138;
output c6156;
output c336;
output c6429;
output c9399;
output c0241;
output c5300;
output c4186;
output c955;
output c6190;
output c5210;
output c88;
output c9370;
output c3102;
output c8296;
output c6475;
output c3257;
output c637;
output c6228;
output c6112;
output c515;
output c3397;
output c271;
output c4281;
output c4410;
output c1251;
output c6216;
output c0136;
output c5112;
output c353;
output c8429;
output c8388;
output c4360;
output c4382;
output c0482;
output c3265;
output c7125;
output c6447;
output c5247;
output c6182;
output c4482;
output c7268;
output c7392;
output c4488;
output c9477;
output c4494;
output c6391;
output c4115;
output c658;
output c9376;
output c7405;
output c684;
output c786;
output c0443;
output c1168;
output c1170;
output c0316;
output c931;
output c810;
output c4165;
output c936;
output c2209;
output c547;
output c8253;
output c9497;
output c925;
output c6215;
output c5357;
output c5470;
output c6389;
output c7478;
output c850;
output c3205;
output c283;
output c1188;
output c1492;
output c1275;
output c634;
output c112;
output c338;
output c6442;
output c58;
output c1129;
output c862;
output c2320;
output c8160;
output c3303;
output c4283;
output c264;
output c741;
output c195;
output c5299;
output c176;
output c1231;
output c93;
output c5367;
output c6218;
output c8341;
output c3183;
output c8227;
output c2256;
output c1356;
output c0163;
output c4219;
output c6110;
output c894;
output c1246;
output c6314;
output c7301;
output c596;
output c340;
output c3113;
output c7166;
output c4462;
output c6386;
output c5358;
output c1178;
output c1264;
output c8170;
output c0470;
output c7399;
output c1354;
output c4441;
output c8210;
output c6244;
output c8221;
output c017;
output c9138;
output c775;
output c2327;
output c549;
output c3315;
output c6425;
output c114;
output c9447;
output c5157;
output c9358;
output c8298;
output c444;
output c927;
output c9367;
output c6199;
output c6349;
output c460;
output c081;
output c8314;
output c9365;
output c9471;
output c1333;
output c4343;
output c1351;
output c5476;
output c2253;
output c7370;
output c0110;
output c2360;
output c416;
output c7165;
output c7489;
output c8486;
output c835;
output c1297;
output c1435;
output c0258;
output c1344;
output c9223;
output c0250;
output c1374;
output c8111;
output c8354;
output c039;
output c225;
output c5215;
output c2357;
output c725;
output c6114;
output c7473;
output c414;
output c686;
output c4369;
output c966;
output c6354;
output c9427;
output c6260;
output c510;
output c020;
output c3134;
output c8342;
output c258;
output c1242;
output c6219;
output c7474;
output c9119;
output c6130;
output c9375;
output c7435;
output c6356;
output c2247;
output c7143;
output c834;
output c9475;
output c6345;
output c047;
output c3308;
output c4342;
output c250;
output c8313;
output c4340;
output c315;
output c9337;
output c8498;
output c754;
output c5123;
output c063;
output c9216;
output c0444;
output c428;
output c6145;
output c8431;
output c8427;
output c2153;
output c987;
output c012;
output c3230;
output c8359;
output c6105;
output c7468;
output c1236;
output c5150;
output c6371;
output c867;
output c3208;
output c3470;
output c1223;
output c2445;
output c228;
output c9281;
output c9301;
output c9335;
output c2374;
output c1125;
output c4146;
output c6357;
output c0474;
output c7306;
output c4442;
output c5189;
output c29;
output c184;
output c6410;
output c3437;
output c8225;
output c5152;
output c9141;
output c6177;
output c9248;
output c7317;
output c0353;
output c3460;
output c4217;
output c2225;
output c394;
output c175;
output c9343;
output c8475;
output c844;
output c1143;
output c8307;
output c1370;
output c0310;
output c415;
output c193;
output c5285;
output c5101;
output c9168;
output c0252;
output c5274;
output c1237;
output c3122;
output c8361;
output c0185;
output c3259;
output c3185;
output c5242;
output c7364;
output c8358;
output c5119;
output c3330;
output c1401;
output c5188;
output c9265;
output c8182;
output c7231;
output c6168;
output c848;
output c1380;
output c9359;
output c164;
output c452;
output c7310;
output c369;
output c2390;
output c1485;
output c1181;
output c6347;
output c7417;
output c7475;
output c989;
output c7115;
output c6326;
output c1329;
output c7424;
output c928;
output c4129;
output c1296;
output c7493;
output c43;
output c3317;
output c3142;
output c9196;
output c7449;
output c9118;
output c1207;
output c7394;
output c2359;
output c5343;
output c619;
output c3184;
output c8336;
output c5212;
output c7386;
output c04;
output c8340;
output c3124;
output c1422;
output c0279;
output c9173;
output c057;
output c5471;
output c1220;
output c8384;
output c8306;
output c014;
output c8280;
output c1478;
output c883;
output c187;
output c8321;
output c2285;
output c2267;
output c7168;
output c2400;
output c4172;
output c9346;
output c1316;
output c2477;
output c548;
output c5305;
output c0253;
output c8337;
output c8419;
output c4350;
output c7278;
output c3188;
output c9234;
output c1442;
output c5335;
output c8417;
output c5417;
output c8432;
output c731;
output c450;
output c8383;
output c718;
output c84;
output c0137;
output c0245;
output c671;
output c3415;
output c8142;
output c4417;
output c933;
output c1398;
output c6432;
output c294;
output c2476;
output c0192;
output c3118;
output c6331;
output c8357;
output c7247;
output c4438;
output c9405;
output c4211;
output c68;
output c4162;
output c688;
output c5238;
output c443;
output c351;
output c0497;
output c1203;
output c6462;
output c3398;
output c2139;
output c7457;
output c4418;
output c4264;
output c9231;
output c7368;
output c6406;
output c3136;
output c4287;
output c7363;
output c287;
output c4275;
output c3293;
output c1450;
output c0355;
output c2483;
output c9181;
output c9151;
output c7338;
output c4334;
output c6139;
output c2142;
output c0342;
output c7431;
output c412;
output c5376;
output c3262;
output c1385;
output c486;
output c235;
output c7196;
output c6265;
output c2260;
output c1135;
output c0499;
output c6120;
output c422;
output c822;
output c5422;
output c50;
output c7205;
output c8268;
output c8335;
output c4375;
output c1166;
output c8289;
output c737;
output c8320;
output c9352;
output c6251;
output c9311;
output c3119;
output c3148;
output c6363;
output c6399;
output c4213;
output c7248;
output c3246;
output c27;
output c5149;
output c089;
output c456;
output c0387;
output c183;
output c4454;
output c2333;
output c2319;
output c1205;
output c3377;
output c3339;
output c7321;
output c1280;
output c0266;
output c6109;
output c6269;
output c367;
output c445;
output c2407;
output c3392;
output c552;
output c7172;
output c4116;
output c0361;
output c4450;
output c6138;
output c751;
output c6213;
output c7108;
output c3111;
output c7264;
output c2351;
output c2474;
output c8317;
output c6160;
output c8283;
output c7210;
output c1474;
output c980;
output c4244;
output c0303;
output c3474;
output c6311;
output c513;
output c2296;
output c8456;
output c9250;
output c1455;
output c5213;
output c0438;
output c9464;
output c4323;
output c8390;
output c871;
output c2271;
output c0300;
output c331;
output c4327;
output c3353;
output c7150;
output c3365;
output c425;
output c5266;
output c6396;
output c4176;
output c4366;
output c0370;
output c6250;
output c6131;
output c034;
output c2429;
output c2379;
output c0369;
output c8294;
output c4266;
output c2338;
output c5290;
output c7233;
output c6174;
output c6492;
output c3479;
output c2427;
output c0149;
output c654;
output c2234;
output c663;
output c20;
output c9430;
output c9139;
output c6137;
output c877;
output c6450;
output c8465;
output c4447;
output c9486;
output c2100;
output c9338;
output c7495;
output c8326;
output c4326;
output c4183;
output c5377;
output c8318;
output c8129;
output c530;
output c6297;
output c895;
output c6186;
output c0169;
output c2274;
output c5221;
output c6121;
output c6283;
output c096;
output c7267;
output c08;
output c879;
output c0219;
output c1134;
output c0113;
output c384;
output c78;
output c814;
output c4344;
output c042;
output c5193;
output c5252;
output c9201;
output c5258;
output c3215;
output c1119;
output c3101;
output c4282;
output c7345;
output c1245;
output c0154;
output c2248;
output c4199;
output c1338;
output c5220;
output c0407;
output c1174;
output c1345;
output c0475;
output c1403;
output c0420;
output c1428;
output c1427;
output c8291;
output c4403;
output c8380;
output c3288;
output c215;
output c153;
output c9396;
output c2366;
output c2273;
output c5104;
output c314;
output c0174;
output c8496;
output c6431;
output c5161;
output c6411;
output c4431;
output c0207;
output c1121;
output c7467;
output c2309;
output c4302;
output c8408;
output c8323;
output c9438;
output c0125;
output c8200;
output c7298;
output c0351;
output c666;
output c6147;
output c8459;
output c77;
output c119;
output c2484;
output c5110;
output c6373;
output c4445;
output c253;
output c390;
output c0277;
output c7124;
output c8204;
output c3150;
output c3370;
output c3361;
output c7342;
output c9327;
output c3192;
output c3457;
output c876;
output c5154;
output c9242;
output c4476;
output c1424;
output c266;
output c9241;
output c3404;
output c86;
output c970;
output c795;
output c6469;
output c1318;
output c218;
output c7334;
output c3182;
output c1323;
output c2302;
output c5311;
output c2372;
output c1313;
output c3139;
output c4246;
output c87;
output c527;
output c0182;
output c9321;
output c1240;
output c8375;
output c770;
output c2134;
output c6200;
output c9316;
output c6393;
output c682;
output c473;
output c773;
output c4472;
output c0213;
output c3364;
output c3486;
output c070;
output c4426;
output c1400;
output c9460;
output c6307;
output c3228;
output c5147;
output c278;
output c8446;
output c6134;
output c771;
output c648;
output c679;
output c2436;
output c1127;
output c6448;
output c5483;
output c0175;
output c5321;
output c1196;
output c7198;
output c8302;
output c4209;
output c3116;
output c237;
output c692;
output c9244;
output c739;
output c4404;
output c5218;
output c1429;
output c3490;
output c7421;
output c6294;
output c6424;
output c0373;
output c586;
output c4250;
output c1418;
output c431;
output c7201;
output c3416;
output c6211;
output c2444;
output c7211;
output c8219;
output c3344;
output c5272;
output c2116;
output c952;
output c2329;
output c9280;
output c7309;
output c3144;
output c616;
output c2499;
output c0480;
output c5457;
output c1101;
output c9440;
output c5227;
output c0287;
output c2308;
output c346;
output c0153;
output c137;
output c1163;
output c5257;
output c9478;
output c5115;
output c1155;
output c317;
output c8295;
output c0448;
output c0199;
output c4208;
output c6158;
output c1147;
output c8479;
output c3236;
output c068;
output c6351;
output c1308;
output c978;
output c8232;
output c9149;
output c16;
output c495;
output c2133;
output c6370;
output c296;
output c387;
output c4153;
output c4187;
output c2269;
output c7428;
output c9286;
output c2443;
output c8198;
output c484;
output c9233;
output c0296;
output c8474;
output c5270;
output c6467;
output c1432;
output c3264;
output c1394;
output c5225;
output c4265;
output c9353;
output c6277;
output c7359;
output c2147;
output c8122;
output c9276;
output c493;
output c6390;
output c7255;
output c1276;
output c6299;
output c419;
output c7178;
output c881;
output c244;
output c8173;
output c524;
output c917;
output c0432;
output c0415;
output c0247;
output c220;
output c7413;
output c1447;
output c8254;
output c7104;
output c1238;
output c7438;
output c4174;
output c2268;
output c946;
output c2291;
output c8444;
output c3197;
output c956;
output c3352;
output c3151;
output c755;
output c3388;
output c132;
output c5465;
output c5109;
output c2202;
output c395;
output c4119;
output c7118;
output c6364;
output c9277;
output c061;
output c4499;
output c1348;
output c827;
output c4421;
output c2120;
output c7107;
output c243;
output c0226;
output c2249;
output c295;
output c6367;
output c8439;
output c5407;
output c0367;
output c551;
output c5323;
output c019;
output c2408;
output c3356;
output c5197;
output c0227;
output c1277;
output c2354;
output c0313;
output c4178;
output c7105;
output c9390;
output c0324;
output c7123;
output c9407;
output c3422;
output c988;
output c2493;
output c5261;
output c2222;
output c977;
output c8387;
output c5320;
output c1255;
output c9404;
output c9351;
output c9360;
output c6346;
output c9144;
output c7258;
output c291;
output c0248;
output c1112;
output c2419;
output c1410;
output c6253;
output c0463;
output c9307;
output c9262;
output c542;
output c914;
output c7341;
output c749;
output c8269;
output c7110;
output c110;
output c131;
output c5348;
output c689;
output c7216;
output c3112;
output c0320;
output c3354;
output c5327;
output c2420;
output c4258;
output c4170;
output c4346;
output c591;
output c7466;
output c3440;
output c3405;
output c9113;
output c4355;
output c5341;
output c762;
output c763;
output c0278;
output c7152;
output c8183;
output c6179;
output c2344;
output c939;
output c2352;
output c9295;
output c6209;
output c7393;
output c9178;
output c1151;
output c9340;
output c1197;
output c7307;
output c1115;
output c269;
output c8157;
output c6257;
output c8118;
output c6394;
output c9369;
output c0204;
output c376;
output c142;
output c5172;
output c6497;
output c2363;
output c056;
output c0391;
output c5133;
output c668;
output c4295;
output c2421;
output c4175;
output c3430;
output c3225;
output c9238;
output c6222;
output c7226;
output c5239;
output c4212;
output c2494;
output c9383;
output c9322;
output c2121;
output c9499;
output c2106;
output c8190;
output c4189;
output c6267;
output c0178;
output c455;
output c1408;
output c5448;
output c4459;
output c9485;
output c7456;
output c0179;
output c5102;
output c9214;
output c0201;
output c2369;
output c7277;
output c7103;
output c6446;
output c1330;
output c0352;
output c8426;
output c5325;
output c5308;
output c0423;
output c9330;
output c3253;
output c5459;
output c7122;
output c5142;
output c8275;
output c0111;
output c15;
output c4455;
output c0327;
output c3299;
output c0106;
output c0200;
output c2399;
output c899;
output c091;
output c6164;
output c9108;
output c196;
output c1198;
output c9402;
output c0411;
output c478;
output c8121;
output c9372;
output c2371;
output c397;
output c6152;
output c9415;
output c4107;
output c9336;
output c9341;
output c2392;
output c433;
output c1120;
output c4374;
output c8457;
output c058;
output c4312;
output c960;
output c5100;
output c459;
output c6379;
output c9392;
output c2331;
output c7353;
output c1191;
output c3284;
output c251;
output c761;
output c2235;
output c6206;
output c7335;
output c2243;
output c0461;
output c6263;
output c2337;
output c2124;
output c9493;
output c4210;
output c3386;
output c0100;
output c472;
output c8193;
output c8156;
output c9484;
output c9229;
output c1108;
output c7265;
output c2233;
output c2276;
output c224;
output c0467;
output c858;
output c683;
output c9170;
output c4485;
output c1473;
output c7415;
output c182;
output c572;
output c7443;
output c711;
output c839;
output c890;
output c8199;
output c9371;
output c7261;
output c0424;
output c6266;
output c5171;
output c5381;
output c1468;
output c0218;
output c1379;
output c7182;
output c6205;
output c8109;
output c96;
output c2191;
output c7378;
output c699;
output c3496;
output c4385;
output c4486;
output c234;
output c8155;
output c2380;
output c2210;
output c4286;
output c0336;
output c556;
output c5206;
output c313;
output c3351;
output c6273;
output c2231;
output c3481;
output c9167;
output c2220;
output c736;
output c4349;
output c4481;
output c2215;
output c6243;
output c4110;
output c8206;
output c6208;
output c0466;
output c0403;
output c7390;
output c8151;
output c8286;
output c0398;
output c611;
output c2462;
output c4132;
output c8264;
output c568;
output c3311;
output c9187;
output c986;
output c5434;
output c8141;
output c8271;
output c3384;
output c4420;
output c9333;
output c0128;
output c5439;
output c5444;
output c2442;
output c9266;
output c9474;
output c480;
output c8461;
output c0214;
output c7142;
output c4238;
output c3394;
output c794;
output c6176;
output c4268;
output c3462;
output c769;
output c8311;
output c641;
output c0344;
output c690;
output c329;
output c8245;
output c0484;
output c254;
output c5400;
output c389;
output c7373;
output c6490;
output c8366;
output c168;
output c1219;
output c6330;
output c2131;
output c9350;
output c4405;
output c075;
output c7362;
output c0436;
output c9458;
output c2377;
output c1311;
output c5174;
output c6106;
output c272;
output c18;
output c0343;
output c7488;
output c2244;
output c080;
output c4383;
output c8212;
output c9121;
output c1482;
output c0210;
output c471;
output c432;
output c6189;
output c8445;
output c748;
output c6167;
output c4122;
output c0146;
output c3252;
output c8215;
output c1463;
output c9190;
output c5451;
output c0453;
output c5141;
output c181;
output c7179;
output c3319;
output c8158;
output c9452;
output c8119;
output c4130;
output c3193;
output c7188;
output c0498;
output c2485;
output c5121;
output c9166;
output c5359;
output c866;
output c9137;
output c9101;
output c8228;
output c0392;
output c1262;
output c7331;
output c1131;
output c0388;
output c3316;
output c6392;
output c7225;
output c670;
output c3332;
output c6317;
output c561;
output c5222;
output c840;
output c920;
output c035;
output c7230;
output c5385;
output c1126;
output c3233;
output c8136;
output c4138;
output c64;
output c0291;
output c7254;
output c022;
output c7273;
output c6332;
output c2135;
output c5181;
output c5347;
output c6175;
output c30;
output c4288;
output c8233;
output c870;
output c2254;
output c0180;
output c4453;
output c5481;
output c2288;
output c9193;
output c342;
output c6358;
output c4193;
output c9377;
output c971;
output c6470;
output c7358;
output c1303;
output c393;
output c3441;
output c9441;
output c3436;
output c7333;
output c7462;
output c1301;
output c533;
output c7416;
output c512;
output c9126;
output c3464;
output c5248;
output c0184;
output c4262;
output c279;
output c3217;
output c115;
output c5234;
output c984;
output c5364;
output c8130;
output c8102;
output c1386;
output c8262;
output c1165;
output c3131;
output c1415;
output c117;
output c4437;
output c1470;
output c213;
output c6154;
output c967;
output c9294;
output c4223;
output c2213;
output c5420;
output c5155;
output c319;
output c2381;
output c727;
output c0255;
output c820;
output c2323;
output c3210;
output c229;
output c5344;
output c5138;
output c2278;
output c7313;
output c7147;
output c5336;
output c930;
output c7274;
output c339;
output c3413;
output c7167;
output c5129;
output c592;
output c7384;
output c8372;
output c7404;
output c5389;
output c6188;
output c81;
output c2188;
output c5404;
output c8322;
output c318;
output c8327;
output c7119;
output c8202;
output c7171;
output c8347;
output c10;
output c6350;
output c0292;
output c0254;
output c2411;
output c6465;
output c0363;
output c22;
output c355;
output c1487;
output c423;
output c9304;
output c789;
output c3407;
output c0408;
output c4182;
output c7304;
output c0202;
output c717;
output c787;
output c7346;
output c0425;
output c9433;
output c5153;
output c5368;
output c2418;
output c3149;
output c8259;
output c6329;
output c5263;
output c3181;
output c180;
output c1420;
output c4361;
output c2203;
output c4155;
output c466;
output c7366;
output c3207;
output c7360;
output c6324;
output c1160;
output c1269;
output c3498;
output c0493;
output c7319;
output c819;
output c4329;
output c9413;
output c65;
output c165;
output c3412;
output c1459;
output c577;
output c146;
output c1289;
output c1287;
output c9240;
output c8237;
output c4253;
output c3484;
output c1309;
output c9203;
output c856;
output c6318;
output c6119;
output c0350;
output c4206;
output c0208;
output c0489;
output c719;
output c0133;
output c7249;
output c4171;
output c5397;
output c0155;
output c9237;
output c7286;
output c4463;
output c464;
output c8231;
output c3459;
output c6444;
output c7235;
output c1471;
output c4173;
output c8273;
output c3107;
output c5351;
output c7411;
output c4303;
output c5423;
output c4226;
output c3199;
output c8462;
output c0322;
output c1271;
output c0195;
output c2195;
output c4216;
output c0435;
output c1247;
output c2107;
output c5105;
output c5265;
output c7429;
output c5456;
output c7227;
output c9279;
output c8405;
output c7170;
output c9462;
output c3209;
output c2143;
output c3211;
output c959;
output c231;
output c5216;
output c5179;
output c3454;
output c1260;
output c8226;
output c6419;
output c7465;
output c0330;
output c811;
output c4124;
output c0368;
output c1426;
output c2435;
output c1225;
output c9444;
output c932;
output c7199;
output c1299;
output c4475;
output c6498;
output c6247;
output c2179;
output c3295;
output c5406;
output c569;
output c681;
output c0123;
output c3452;
output c51;
output c5446;
output c1407;
output c2335;
output c8140;
output c0104;
output c0348;
output c880;
output c1377;
output c5430;
output c3229;
output c297;
output c1402;
output c6275;
output c5489;
output c9129;
output c0481;
output c5190;
output c9381;
output c9324;
output c817;
output c2166;
output c9463;
output c4440;
output c5264;
output c579;
output c1172;
output c4433;
output c470;
output c5467;
output c0141;
output c1161;
output c7318;
output c9435;
output c972;
output c6339;
output c6202;
output c8117;
output c3115;
output c612;
output c8378;
output c614;
output c2145;
output c4345;
output c1265;
output c4135;
output c5111;
output c1153;
output c4314;
output c5229;
output c1267;
output c8243;
output c47;
output c6261;
output c7344;
output c582;
output c3312;
output c8385;
output c4133;
output c7183;
output c4478;
output c0377;
output c758;
output c6378;
output c860;
output c5268;
output c4191;
output c4112;
output c5403;
output c6136;
output c7214;
output c116;
output c521;
output c9208;
output c7180;
output c6454;
output c6453;
output c1326;
output c8331;
output c8132;
output c489;
output c01;
output c320;
output c5237;
output c3373;
output c2137;
output c9445;
output c9368;
output c0430;
output c7159;
output c2402;
output c6385;
output c2128;
output c3285;
output c3379;
output c282;
output c796;
output c5388;
output c8104;
output c2185;
output c6268;
output c8133;
output c275;
output c6237;
output c7263;
output c1137;
output c3235;
output c5292;
output c6197;
output c122;
output c488;
output c8126;
output c1217;
output c332;
output c9227;
output c8470;
output c157;
output c4294;
output c0196;
output c0211;
output c7184;
output c0236;
output c4168;
output c529;
output c5484;
output c4430;
output c8345;
output c9331;
output c5233;
output c467;
output c6486;
output c7299;
output c8377;
output c5356;
output c6148;
output c3145;
output c0194;
output c8162;
output c7151;
output c9408;
output c540;
output c0427;
output c4353;
output c54;
output c7194;
output c7292;
output c0205;
output c9409;
output c3431;
output c8180;
output c558;
output c39;
output c7100;
output c537;
output c975;
output c9115;
output c8391;
output c3491;
output c490;
output c0225;
output c5490;
output c6403;
output c2101;
output c7402;
output c8362;
output c6184;
output c8246;
output c5463;
output c2198;
output c9258;
output c086;
output c7379;
output c7339;
output c2345;
output c0319;
output c2306;
output c8191;
output c5415;
output c656;
output c5145;
output c3350;
output c593;
output c4315;
output c9389;
output c4444;
output c5267;
output c1200;
output c5201;
output c0109;
output c6484;
output c7217;
output c713;
output c4468;
output c8433;
output c95;
output c9179;
output c4241;
output c149;
output c72;
output c9461;
output c3334;
output c9245;
output c4497;
output c1452;
output c8499;
output c2446;
output c3292;
output c782;
output c8355;
output c6308;
output c620;
output c141;
output c1352;
output c3297;
output c5382;
output c696;
output c0382;
output c2159;
output c6457;
output c0118;
output c4222;
output c7476;
output c783;
output c9224;
output c9378;
output c256;
output c630;
output c1193;
output c730;
output c1388;
output c9470;
output c333;
output c1491;
output c349;
output c5209;
output c1495;
output c3195;
output c335;
output c8234;
output c2257;
output c2103;
output c1461;
output c4260;
output c3304;
output c979;
output c57;
output c3447;
output c6372;
output c1425;
output c9400;
output c9454;
output c2172;
output c3475;
output c6328;
output c6285;
output c2343;
output c4140;
output c4496;
output c7487;
output c5165;
output c5200;
output c8400;
output c7111;
output c4251;
output c7224;
output c8249;
output c1189;
output c3360;
output c2388;
output c2258;
output c2316;
output c3198;
output c2413;
output c0308;
output c4150;
output c4228;
output c5143;
output c4389;
output c9164;
output c0405;
output c6155;
output c664;
output c7458;
output c1298;
output c729;
output c5332;
output c5241;
output c1465;
output c0290;
output c5425;
output c6101;
output c7283;
output c4464;
output c2453;
output c6104;
output c9362;
output c5198;
output c3425;
output c949;
output c4364;
output c344;
output c5486;
output c5370;
output c1421;
output c622;
output c5116;
output c6305;
output c4248;
output c0267;
output c3226;
output c6478;
output c7414;
output c9112;
output c7131;
output c6460;
output c3170;
output c1192;
output c2136;
output c0464;
output c4413;
output c1281;
output c9297;
output c0347;
output c2146;
output c0209;
output c0410;
output c0261;
output c388;
output c6340;
output c6293;
output c7440;
output c724;
output c7289;
output c7296;
output c2475;
output c3423;
output c9220;
output c8454;
output c410;
output c639;
output c4432;
output c7348;
output c1397;
output c7396;
output c8392;
output c4105;
output c6395;
output c4446;
output c5108;
output c9391;
output c7352;
output c214;
output c7222;
output c4197;
output c3463;
output c687;
output c0395;
output c2204;
output c2149;
output c1320;
output c9221;
output c0390;
output c733;
output c1477;
output c5113;
output c356;
output c2183;
output c4240;
output c5342;
output c6338;
output c268;
output c7246;
output c6298;
output c8165;
output c4259;
output c8250;
output c6281;
output c2468;
output c6319;
output c6111;
output c2394;
output c468;
output c8256;
output c8115;
output c016;
output c5450;
output c7380;
output c528;
output c8150;
output c7374;
output c8267;
output c3171;
output c6359;
output c2181;
output c0406;
output c5287;
output c6230;
output c7287;
output c753;
output c2303;
output c0244;
output c12;
output c3442;
output c7420;
output c5375;
output c788;
output c1232;
output c7355;
output c4321;
output c525;
output c3359;
output c5386;
output c5315;
output c580;
output c893;
output c7349;
output c3383;
output c2397;
output c6485;
output c938;
output c5346;
output c9157;
output c13;
output c3104;
output c9122;
output c9219;
output c041;
output c4393;
output c0479;
output c210;
output c3200;
output c1378;
output c4154;
output c6271;
output c9344;
output c5466;
output c8293;
output c9102;
output c6239;
output c0494;
output c7426;
output c062;
output c923;
output c3275;
output c8413;
output c1376;
output c35;
output c2487;
output c0404;
output c3443;
output c1230;
output c366;
output c816;
output c6127;
output c821;
output c0401;
output c2482;
output c0431;
output c113;
output c1493;
output c7175;
output c261;
output c3133;
output c2450;
output c0374;
output c9397;
output c7354;
output c3121;
output c8374;
output c8416;
output c9398;
output c2157;
output c8284;
output c0143;
output c4379;
output c4134;
output c9426;
output c7437;
output c9442;
output c065;
output c2261;
output c3449;
output c5366;
output c590;
output c7316;
output c133;
output c4493;
output c5414;
output c9491;
output c7129;
output c221;
output c2148;
output c0472;
output c3165;
output c8287;
output c8351;
output c934;
output c0302;
output c6214;
output c1480;
output c9268;
output c7461;
output c1384;
output c0454;
output c8236;
output c553;
output c6488;
output c6435;
output c14;
output c2123;
output c8244;
output c2463;
output c0285;
output c6472;
output c8423;
output c2127;
output c0338;
output c4157;
output c211;
output c345;
output c8217;
output c0176;
output c0364;
output c3382;
output c8389;
output c0129;
output c5369;
output c7450;
output c5438;
output c052;
output c8229;
output c233;
output c481;
output c0441;
output c2144;
output c3263;
output c170;
output c2297;
output c9282;
output c757;
output c4338;
output c5350;
output c3143;
output c8107;
output c4111;
output c4358;
output c7135;
output c9328;
output c5214;
output c2287;
output c073;
output c1373;
output c8148;
output c1274;
output c0151;
output c479;
output c969;
output c595;
output c9162;
output c1263;
output c3409;
output c385;
output c8131;
output c3429;
output c1190;
output c9492;
output c6422;
output c9421;
output c4231;
output c7490;
output c6400;
output c8348;
output c37;
output c8473;
output c7252;
output c6463;
output c3301;
output c8353;
output c8482;
output c0335;
output c863;
output c4257;
output c7253;
output c6322;
output c891;
output c645;
output c8103;
output c9199;
output c3387;
output c5276;
output c4332;
output c6415;
output c3333;
output c2496;
output c7257;
output c2104;
output c4255;
output c3234;
output c045;
output c4236;
output c5309;
output c7262;
output c3286;
output c5399;
output c723;
output c6380;
output c2229;
output c742;
output c4362;
output c171;
output c3261;
output c743;
output c1295;
output c7282;
output c1364;
output c469;
output c6337;
output c5136;
output c797;
output c8177;
output c19;
output c9239;
output c2432;
output c7144;
output c599;
output c378;
output c076;
output c7223;
output c9267;
output c623;
output c8478;
output c8235;
output c2182;
output c013;
output c9289;
output c2290;
output c9364;
output c4254;
output c1221;
output c1145;
output c6287;
output c139;
output c9319;
output c3390;
output c4234;
output c0222;
output c9156;
output c430;
output c2365;
output c2307;
output c6224;
output c3428;
output c5158;
output c6151;
output c143;
output c239;
output c2423;
output c9308;
output c7155;
output c5262;
output c9284;
output c9406;
output c5259;
output c3362;
output c570;
output c7486;
output c0357;
output c1411;
output c576;
output c1337;
output c3177;
output c6262;
output c4434;
output c3493;
output c9116;
output c7156;
output c9296;
output c1306;
output c8424;
output c3488;
output c3408;
output c6437;
output c5163;
output c8196;
output c2238;
output c4320;
output c71;
output c0159;
output c8409;
output c2460;
output c1234;
output c6456;
output c538;
output c991;
output c4412;
output c0217;
output c859;
output c044;
output c418;
output c8163;
output c8290;
output c0228;
output c4274;
output c8147;
output c3103;
output c4117;
output c1350;
output c7256;
output c4196;
output c1438;
output c263;
output c3174;
output c9135;
output c2286;
output c9130;
output c027;
output c2298;
output c830;
output c0140;
output c5162;
output c1456;
output c1167;
output c6398;
output c3478;
output c8239;
output c8369;
output c5487;
output c121;
output c477;
output c1321;
output c7329;
output c2199;
output c7327;
output c4461;
output c892;
output c2132;
output c8379;
output c7497;
output c0183;
output c3345;
output c4230;
output c1132;
output c9287;
output c2255;
output c352;
output c4357;
output c6166;
output c7336;
output c4368;
output c7136;
output c5251;
output c9100;
output c8422;
output c4298;
output c4480;
output c567;
output c4237;
output c3406;
output c6220;
output c3277;
output c7114;
output c5184;
output c6232;
output c4290;
output c9183;
output c9251;
output c2184;
output c6428;
output c9488;
output c3483;
output c1227;
output c7381;
output c8407;
output c1164;
output c9361;
output c651;
output c6480;
output c1443;
output c5164;
output c011;
output c3223;
output c031;
output c9171;
output c759;
output c5340;
output c5166;
output c9424;
output c2396;
output c025;
output c3310;
output c2189;
output c7139;
output c4198;
output c2206;
output c924;
output c8328;
output c482;
output c9347;
output c7347;
output c8168;
output c0190;
output c1253;
output c8174;
output c6459;
output c9481;
output c277;
output c5409;
output c6192;
output c7491;
output c0397;
output c732;
output c3434;
output c6445;
output c4436;
output c6327;
output c965;
output c1382;
output c3271;
output c5245;
output c0240;
output c4392;
output c4180;
output c4457;
output c217;
output c633;
output c321;
output c3202;
output c3106;
output c4448;
output c5191;
output c7453;
output c2165;
output c4308;
output c951;
output c4194;
output c6323;
output c3417;
output c4341;
output c6421;
output c4305;
output c53;
output c1209;
output c1252;
output c8112;
output c961;
output c3196;
output c698;
output c3274;
output c0284;
output c997;
output c8207;
output c6276;
output c163;
output c0172;
output c5449;
output c3458;
output c396;
output c8261;
output c884;
output c2250;
output c7460;
output c9110;
output c565;
output c5240;
output c8105;
output c778;
output c0220;
output c9247;
output c2163;
output c4352;
output c4489;
output c852;
output c587;
output c5301;
output c1171;
output c8143;
output c531;
output c0380;
output c1118;
output c5273;
output c922;
output c9448;
output c1419;
output c993;
output c772;
output c0107;
output c5195;
output c9410;
output c722;
output c9394;
output c8397;
output c8188;
output c03;
output c5393;
output c4296;
output c9305;
output c197;
output c7163;
output c3318;
output c0483;
output c519;
output c4152;
output c2470;
output c842;
output c3276;
output c7382;
output c9288;
output c6321;
output c7209;
output c0203;
output c4273;
output c4333;
output c6117;
output c8125;
output c7300;
output c7397;
output c144;
output c0242;
output c6423;
output c3451;
output c8178;
output c6240;
output c4202;
output c7212;
output c4452;
output c7422;
output c8137;
output c9270;
output c9225;
output c5416;
output c4195;
output c1393;
output c3126;
output c1334;
output c3368;
output c0345;
output c6481;
output c9230;
output c2322;
output c1182;
output c8303;
output c4373;
output c5295;
output c5151;
output c4100;
output c7245;
output c9483;
output c9163;
output c9212;
output c1413;
output c5131;
output c059;
output c1381;
output c9320;
output c710;
output c0385;
output c3485;
output c3497;
output c5392;
output c1453;
output c3349;
output c1361;
output c75;
output c6376;
output c995;
output c7459;
output c7494;
output c160;
output c285;
output c4147;
output c6107;
output c720;
output c3456;
output c198;
output c73;
output c0381;
output c6144;
output c128;
output c9498;
output c4227;
output c7242;
output c5224;
output c6316;
output c1206;
output c0341;
output c3221;
output c8263;
output c6252;
output c8460;
output c0456;
output c642;
output c3157;
output c0449;
output c427;
output c3331;
output c5192;
output c9318;
output c2176;
output c5378;
output c1494;
output c311;
output c8299;
output c1310;
output c2362;
output c0433;
output c6128;
output c63;
output c0446;
output c8154;
output c6290;
output c1367;
output c1103;
output c9269;
output c3189;
output c5433;
output c3167;
output c2293;
output c5156;
output c7383;
output c4224;
output c5130;
output c8310;
output c0257;
output c3376;
output c4203;
output c226;
output c4347;
output c2459;
output c9211;
output c91;
output c6355;
output c7357;
output c222;
output c2464;
output c363;
output c6436;
output c652;
output c0232;
output c0384;
output c5345;
output c2155;
output c6153;
output c087;
output c4289;
output c5176;
output c6146;
output c4359;
output c1177;
output c2178;
output c442;
output c4439;
output c864;
output c41;
output c6198;
output c6143;
output c1467;
output c4390;
output c289;
output c2108;
output c4387;
output c6185;
output c2138;
output c8288;
output c7202;
output c0144;
output c1268;
output c8128;
output c589;
output c4225;
output c5401;
output c3194;
output c083;
output c0275;
output c1284;
output c8350;
output c1128;
output c3243;
output c7315;
output c781;
output c2152;
output c462;
output c1314;
output c644;
output c0340;
output c9342;
output c3249;
output c2117;
output c6309;
output c0476;
output c752;
output c0198;
output c0317;
output c6300;
output c2364;
output c2169;
output c6149;
output c9263;
output c2105;
output c6417;
output c5288;
output c6387;
output c0171;
output c9243;
output c6113;
output c1444;
output c8490;
output c8449;
output c8393;
output c0181;
output c2190;
output c0272;
output c3455;
output c539;
output c2168;
output c7387;
output c4139;
output c0417;
output c3227;
output c1116;
output c6404;
output c8195;
output c347;
output c6223;
output c981;
output c3153;
output c4467;
output c4474;
output c6315;
output c7158;
output c9309;
output c2489;
output c4415;
output c9357;
output c4310;
output c4249;
output c0221;
output c5307;
output c8248;
output c0413;
output c566;
output c3125;
output c976;
output c6433;
output c3110;
output c5495;
output c6496;
output c0108;
output c1395;
output c0412;
output c2422;
output c9159;
output c868;
output c5329;
output c435;
output c943;
output c7294;
output c5339;
output c6369;
output c8406;
output c0333;
output c7391;
output c0434;
output c4151;
output c581;
output c9226;
output c5278;
output c9302;
output c337;
output c7192;
output c2102;
output c370;
output c8430;
output c499;
output c7436;
output c5205;
output c8211;
output c398;
output c364;
output c3272;
output c257;
output c4377;
output c0276;
output c6414;
output c0294;
output c7229;
output c1346;
output c2332;
output c5291;
output c9431;
output c0428;
output c6491;
output c5281;
output c0288;
output c3283;
output c4337;
output c238;
output c3154;
output c574;
output c3146;
output c5352;
output c897;
output c7376;
output c647;
output c1105;
output c4429;
output c1332;
output c6292;
output c465;
output c8480;
output c136;
output c2382;
output c033;
output c5126;
output c0270;
output c6313;
output c9382;
output c0206;
output c776;
output c0366;
output c399;
output c0289;
output c1250;
output c518;
output c6412;
output c7190;
output c5132;
output c2180;
output c2110;
output c7498;
output c8373;
output c8218;
output c9422;
output c3220;
output c829;
output c3117;
output c0393;
output c4419;
output c8463;
output c0321;
output c5186;
output c3338;
output c223;
output c374;
output c3222;
output c974;
output c613;
output c2428;
output c126;
output c0246;
output c0468;
output c3342;
output c8152;
output c212;
output c929;
output c5338;
output c9255;
output c98;
output c1392;
output c7148;
output c0119;
output c5159;
output c3314;
output c324;
output c5355;
output c2350;
output c4425;
output c5349;
output c4103;
output c6258;
output c1479;
output c4317;
output c4156;
output c9111;
output c517;
output c0115;
output c6183;
output c4313;
output c1457;
output c293;
output c9373;
output c9418;
output c7356;
output c888;
output c3329;
output c7239;
output c46;
output c358;
output c7237;
output c9412;
output c7375;
output c6248;
output c6207;
output c1335;
output c377;
output c3156;
output c6303;
output c4163;
output c657;
output c714;
output c190;
output c2284;
output c9125;
output c7395;
output c3191;
output c7117;
output c9494;
output c7447;
output c2130;
output c0457;
output c147;
output c8412;
output c3152;
output c9332;
output c7285;
output c3489;
output c7312;
output c2439;
output c1124;
output c847;
output c0306;
output c7492;
output c0421;
output c8483;
output c0477;
output c7324;
output c3213;
output c1288;
output c2495;
output c7137;
output c037;
output c694;
output c7308;
output c3224;
output c4484;
output c5211;
output c6150;
output c7269;
output c9423;
output c0360;
output c487;
output c4351;
output c049;
output c1254;
output c6374;
output c5316;
output c7407;
output c5398;
output c511;
output c1451;
output c89;
output c2299;
output c1342;
output c0124;
output c5128;
output c575;
output c1436;
output c9228;
output c386;
output c8386;
output c1439;
output c2367;
output c2473;
output c188;
output c3109;
output c550;
output c1159;
output c2451;
output c3306;
output c120;
output c2270;
output c1148;
output c154;
output c5117;
output c2481;
output c2368;
output c3238;
output c5461;
output c6377;
output c9449;
output c3477;
output c0315;
output c9127;
output c3267;
output c242;
output c7451;
output c8472;
output c0396;
output c7361;
output c2414;
output c281;
output c4169;
output c5120;
output c1434;
output c0491;
output c4125;
output c1362;
output c8205;
output c2325;
output c6180;
output c7481;
output c6163;
output c064;
output c3180;
output c4149;
output c3420;
output c4471;
output c8402;
output c3399;
output c8339;
output c018;
output c6270;
output c9177;
output c885;
output c536;
output c476;
output c173;
output c06;
output c2122;
output c992;
output c7328;
output c8453;
output c5436;
output c615;
output c7191;
output c0166;
output c4307;
output c916;
output c869;
output c4271;
output c236;
output c1406;
output c2194;
output c9215;
output c8282;
output c6171;
output c1365;
output c843;
output c9206;
output c5474;
output c2125;
output c5460;
output c1146;
output c6461;
output c0490;
output c5493;
output c5125;
output c3444;
output c249;
output c9490;
output c328;
output c2395;
output c7332;
output c9300;
output c9293;
output c3343;
output c5390;
output c6100;
output c7132;
output c5472;
output c9184;
output c0135;
output c8376;
output c9325;
output c44;
output c4304;
output c5230;
output c2406;
output c728;
output c1222;
output c1123;
output c284;
output c6178;
output c9414;
output c2164;
output c2353;
output c0329;
output c3341;
output c3175;
output c655;
output c0160;
output c2426;
output c1149;
output c9114;
output c0281;
output c437;
output c5442;
output c7126;
output c6129;
output c2161;
output c092;
output c9472;
output c1371;
output c350;
output c3105;
output c8344;
output c6440;
output c1241;
output c9487;
output c6255;
output c0337;
output c4322;
output c2312;
output c0358;
output c2321;
output c5260;
output c179;
output c7434;
output c4470;
output c9271;
output c8494;
output c4473;
output c0305;
output c4131;
output c9261;
output c3499;
output c7244;
output c1279;
output c6159;
output c957;
output c270;
output c0459;
output c1138;
output c983;
output c9303;
output c3260;
output c4166;
output c9482;
output c3495;
output c9374;
output c799;
output c130;
output c125;
output c7204;
output c6302;
output c8308;
output c6416;
output c7293;
output c3176;
output c854;
output c4108;
output c9192;
output c7326;
output c9473;
output c3258;
output c8281;
output c8139;
output c5499;
output c9236;
output c516;
output c5183;
output c6231;
output c4330;
output c0165;
output c448;
output c4424;
output c1404;
output c6282;
output c361;
output c379;
output c9218;
output c0260;
output c8266;
output c83;
output c865;
output c6495;
output c9153;
output c2461;
output c4291;
output c1158;
output c7480;
output c2232;
output c5322;
output c2301;
output c4137;
output c3450;
output c6336;
output c391;
output c964;
output c392;
output c030;
output c522;
output c5384;
output c6132;
output c2113;
output c8260;
output c3203;
output c74;
output c1341;
output c621;
output c0312;
output c2486;
output c2167;
output c7441;
output c5127;
output c5118;
output c7433;
output c6288;
output c1490;
output c327;
output c0152;
output c5475;
output c3336;
output c588;
output c6133;
output c9148;
output c6272;
output c6476;
output c0426;
output c9246;
output c7127;
output c0485;
output c066;
output c6279;
output c5178;
output c5379;
output c5160;
output c5254;
output c097;
output c4449;
output c6388;
output c5437;
output c0478;
output c3320;
output c6212;
output c8304;
output c563;
output c9457;
output c1405;
output c0191;
output c3186;
output c5334;
output c383;
output c322;
output c8395;
output c9124;
output c084;
output c846;
output c0273;
output c948;
output c1440;
output c8106;
output c996;
output c0157;
output c2447;
output c8437;
output c9169;
output c439;
output c245;
output c8436;
output c8270;
output c7398;
output c79;
output c2230;
output c8258;
output c5139;
output c6115;
output c8138;
output c3256;
output c0150;
output c5395;
output c8352;
output c5304;
output c941;
output c2398;
output c7448;
output c2246;
output c9495;
output c583;
output c6225;
output c1202;
output c3173;
output c118;
output c2313;
output c3347;
output c7203;
output c7305;
output c3245;
output c7251;
output c2114;
output c735;
output c9213;
output c2239;
output c9154;
output c3147;
output c046;
output c6235;
output c5243;
output c3251;
output c873;
output c9232;
output c1152;
output c7297;
output c59;
output c6126;
output c7160;
output c0325;
output c1102;
output c571;
output c3300;
output c7463;
output c1359;
output c2126;
output c6162;
output c3140;
output c8488;
output c5317;
output c1446;
output c833;
output c129;
output c0495;
output c2373;
output c7106;
output c5331;
output c9349;
output c4465;
output c4145;
output c9429;
output c5303;
output c7389;
output c831;
output c9185;
output c6342;
output c4279;
output c3438;
output c4416;
output c9420;
output c2479;
output c832;
output c3465;
output c70;
output c1294;
output c2356;
output c8279;
output c7377;
output c6405;
output c2240;
output c4215;
output c0486;
output c5208;
output c2471;
output c1416;
output c3363;
output c3187;
output c7113;
output c6489;
output c325;
output c5453;
output c597;
output c5408;
output c5427;
output c5373;
output c1156;
output c2295;
output c1369;
output c8435;
output c8176;
output c5318;
output c2282;
output c3281;
output c3216;
output c6464;
output c4409;
output c9388;
output c1109;
output c1239;
output c624;
output c4309;
output c9443;
output c3164;
output c354;
output c85;
output c8451;
output c2162;
output c145;
output c9366;
output c9133;
output c5360;
output c6325;
output c935;
output c557;
output c9160;
output c7260;
output c6473;
output c6203;
output c697;
output c919;
output c2237;
output c8285;
output c3366;
output c3492;
output c4136;
output c6102;
output c6234;
output c9103;
output c726;
output c7140;
output c7388;
output c1499;
output c00;
output c0256;
output c5226;
output c0297;
output c5485;
output c7423;
output c9186;
output c7219;
output c5167;
output c8468;
output c298;
output c6165;
output c7238;
output c1464;
output c0112;
output c5283;
output c5275;
output c1184;
output c3400;
output c2441;
output c998;
output c2263;
output c617;
output c886;
output c4451;
output c368;
output c0331;
output c2173;
output c0262;
output c1325;
output c6187;
output c7403;
output c653;
output c9312;
output c1396;
output c9147;
output c5469;
output c316;
output c2385;
output c9278;
output c7400;
output c3325;
output c1481;
output c0188;
output c9434;
output c3357;
output c7218;
output c1460;
output c5231;
output c9419;
output c4370;
output c8312;
output c6420;
output c9146;

assign c00 =  x231 &  x534 & ~x123 & ~x414 & ~x637;
assign c02 =  x408 &  x436 & ~x38 & ~x149 & ~x291 & ~x579 & ~x666 & ~x744;
assign c04 =  x431 &  x549 &  x603 & ~x420 & ~x545;
assign c06 =  x93 &  x149 &  x206 &  x262 &  x346 &  x402;
assign c08 =  x167;
assign c010 =  x594 & ~x9 & ~x43 & ~x241 & ~x379 & ~x380 & ~x428 & ~x431 & ~x436 & ~x641;
assign c012 =  x205 &  x261 & ~x183 & ~x356 & ~x395 & ~x438 & ~x720;
assign c014 =  x634 & ~x240 & ~x664;
assign c016 =  x261 &  x288 &  x316 &  x456 & ~x152 & ~x187 & ~x449 & ~x617;
assign c018 =  x26 &  x53;
assign c020 =  x312 &  x484 &  x509 & ~x13 & ~x66 & ~x93 & ~x293 & ~x714 & ~x726;
assign c022 =  x783;
assign c024 =  x332 &  x419;
assign c026 =  x231 &  x232 &  x315 &  x316 &  x480 & ~x588;
assign c028 =  x204 &  x232 & ~x125 & ~x198 & ~x293 & ~x328 & ~x348 & ~x435 & ~x751;
assign c030 =  x521 & ~x2 & ~x48 & ~x61 & ~x77 & ~x108 & ~x139 & ~x155 & ~x392 & ~x395 & ~x476 & ~x478 & ~x705 & ~x722;
assign c032 =  x544 &  x545 &  x594;
assign c034 =  x26;
assign c036 =  x177 &  x552 & ~x99 & ~x239 & ~x356;
assign c038 = ~x39 & ~x53 & ~x80 & ~x98 & ~x111 & ~x209 & ~x210 & ~x240 & ~x246 & ~x266 & ~x353 & ~x505 & ~x720 & ~x745;
assign c040 =  x289 &  x317 &  x456 &  x484 &  x485 & ~x14 & ~x108 & ~x140 & ~x394 & ~x421 & ~x504 & ~x697 & ~x703 & ~x721 & ~x746 & ~x753 & ~x757 & ~x779;
assign c042 =  x509 &  x512 &  x536;
assign c044 =  x371 & ~x180 & ~x243 & ~x269 & ~x364 & ~x475 & ~x607 & ~x619 & ~x645 & ~x647 & ~x687 & ~x719;
assign c046 =  x167;
assign c048 =  x146 &  x232 & ~x65 & ~x157 & ~x324;
assign c050 =  x65 &  x93 &  x261 &  x373;
assign c052 = ~x121 & ~x181 & ~x218 & ~x243 & ~x411 & ~x551 & ~x576 & ~x579 & ~x580 & ~x650 & ~x709 & ~x776;
assign c054 =  x498 & ~x1 & ~x184 & ~x337 & ~x356 & ~x602 & ~x709;
assign c056 =  x460 &  x577 & ~x148;
assign c058 =  x177 & ~x80 & ~x266 & ~x356 & ~x414 & ~x467;
assign c060 =  x122 &  x289 & ~x68 & ~x74 & ~x153 & ~x336 & ~x672 & ~x776;
assign c062 =  x173 &  x258 &  x397 &  x480 & ~x11 & ~x65 & ~x150 & ~x239;
assign c064 =  x26;
assign c066 =  x65 &  x93 &  x149 &  x177 & ~x213 & ~x605;
assign c068 =  x232 &  x260 &  x427 & ~x311 & ~x659 & ~x757;
assign c070 =  x27 &  x699;
assign c072 =  x543 &  x569 &  x595 & ~x176 & ~x379;
assign c074 =  x167 &  x223;
assign c076 =  x0;
assign c078 =  x439 &  x493 &  x494 &  x521 & ~x38 & ~x59 & ~x66 & ~x96 & ~x123 & ~x744;
assign c080 =  x511 & ~x38 & ~x328 & ~x345 & ~x709;
assign c082 = ~x71 & ~x129 & ~x138 & ~x213 & ~x243 & ~x269 & ~x270 & ~x272 & ~x328 & ~x356 & ~x474 & ~x517 & ~x680 & ~x706 & ~x713 & ~x775;
assign c084 =  x515 &  x577 & ~x36 & ~x367 & ~x393 & ~x395 & ~x422 & ~x764;
assign c086 =  x285 &  x433 &  x456 & ~x123;
assign c088 =  x65 &  x94 &  x260 &  x372 & ~x740;
assign c092 =  x203 & ~x11 & ~x39 & ~x53 & ~x156 & ~x302 & ~x317 & ~x347 & ~x356 & ~x358 & ~x449 & ~x520 & ~x547;
assign c094 =  x174 &  x204 & ~x38 & ~x74 & ~x208 & ~x237 & ~x606;
assign c096 =  x140;
assign c098 =  x204 &  x484 & ~x185 & ~x266 & ~x492 & ~x671 & ~x705 & ~x745;
assign c0100 =  x517 &  x542 &  x567 & ~x14 & ~x750;
assign c0102 =  x261 &  x262 &  x289 &  x317 &  x512 & ~x29 & ~x85 & ~x86 & ~x505 & ~x641;
assign c0104 =  x559 &  x573;
assign c0106 =  x517 & ~x48 & ~x320 & ~x354;
assign c0108 =  x55;
assign c0110 =  x172 &  x173 &  x174 & ~x123 & ~x619 & ~x665 & ~x750 & ~x767;
assign c0114 =  x473 &  x484 &  x547 & ~x11 & ~x71 & ~x779;
assign c0116 = ~x42 & ~x94 & ~x108 & ~x161 & ~x187 & ~x271 & ~x647 & ~x653 & ~x692;
assign c0118 =  x204 &  x232 &  x483 &  x536 & ~x38 & ~x125 & ~x182 & ~x686 & ~x712;
assign c0120 =  x261 &  x262 &  x288 &  x345 &  x540 & ~x14 & ~x322 & ~x326;
assign c0122 = ~x22 & ~x25 & ~x41 & ~x52 & ~x102 & ~x123 & ~x267 & ~x320 & ~x327 & ~x410 & ~x449 & ~x531 & ~x665 & ~x668 & ~x712 & ~x716;
assign c0124 =  x91 &  x204 &  x260 &  x316 & ~x599;
assign c0126 =  x120 & ~x69 & ~x266 & ~x271 & ~x436 & ~x502 & ~x515 & ~x692;
assign c0128 =  x200 &  x506 & ~x726;
assign c0130 =  x83;
assign c0132 =  x83;
assign c0134 =  x463 &  x484 &  x536 & ~x11;
assign c0136 =  x27;
assign c0138 =  x167;
assign c0140 =  x456 &  x484 &  x509 & ~x395;
assign c0142 =  x150 &  x261 &  x289 & ~x106 & ~x269 & ~x306 & ~x605;
assign c0144 =  x281 &  x481;
assign c0146 =  x83;
assign c0148 =  x599 &  x623 & ~x10 & ~x86 & ~x106 & ~x449;
assign c0150 =  x205 &  x261 & ~x60 & ~x223 & ~x324 & ~x395 & ~x616 & ~x752 & ~x772;
assign c0154 =  x147 &  x231 & ~x10 & ~x22 & ~x151 & ~x327 & ~x384 & ~x731;
assign c0156 =  x388 &  x484 &  x547 & ~x298 & ~x336;
assign c0158 =  x261 &  x343 &  x511 & ~x366 & ~x410 & ~x627;
assign c0160 =  x494 &  x521 &  x549 & ~x39 & ~x68 & ~x124 & ~x641 & ~x705;
assign c0162 =  x461 &  x503 &  x511 & ~x424;
assign c0164 =  x232 &  x427 &  x567 & ~x263 & ~x410 & ~x520;
assign c0166 =  x368 & ~x30 & ~x269 & ~x320 & ~x561 & ~x686 & ~x693 & ~x697;
assign c0170 = ~x30 & ~x124 & ~x187 & ~x212 & ~x215 & ~x321 & ~x328 & ~x351 & ~x379 & ~x572 & ~x641;
assign c0172 =  x111;
assign c0174 =  x459 & ~x272 & ~x404 & ~x687;
assign c0176 =  x599 &  x620 & ~x326 & ~x395;
assign c0178 =  x457 & ~x44 & ~x73 & ~x212 & ~x269 & ~x270 & ~x299 & ~x356 & ~x357 & ~x702 & ~x726 & ~x776 & ~x782;
assign c0180 =  x199 &  x478;
assign c0182 =  x408 & ~x289 & ~x582 & ~x583 & ~x675;
assign c0184 = ~x125 & ~x187 & ~x302 & ~x318 & ~x446;
assign c0186 =  x231 &  x232 &  x371 & ~x328 & ~x547 & ~x602 & ~x721;
assign c0188 =  x783;
assign c0190 =  x147 &  x258 & ~x11 & ~x39 & ~x318 & ~x378 & ~x434;
assign c0192 =  x85;
assign c0194 =  x452 & ~x11 & ~x27 & ~x32 & ~x49 & ~x78 & ~x102 & ~x110 & ~x134 & ~x150 & ~x161 & ~x327 & ~x602 & ~x696 & ~x751;
assign c0196 =  x226;
assign c0198 =  x378 &  x453 & ~x210;
assign c0200 =  x550 & ~x638 & ~x664;
assign c0202 =  x479;
assign c0204 =  x518 &  x592 & ~x34 & ~x101 & ~x186 & ~x422;
assign c0206 =  x24;
assign c0208 =  x316 &  x317 &  x318 &  x486 &  x512 & ~x46 & ~x718;
assign c0210 =  x510 &  x518 & ~x496;
assign c0212 =  x173 & ~x22 & ~x196 & ~x465 & ~x550 & ~x579 & ~x586 & ~x694;
assign c0214 = ~x105 & ~x184 & ~x213 & ~x223 & ~x240 & ~x246 & ~x350 & ~x380 & ~x410 & ~x414 & ~x492 & ~x551 & ~x578 & ~x671;
assign c0216 =  x756;
assign c0218 =  x83;
assign c0220 =  x261 &  x262 &  x317 &  x345 &  x513 & ~x395;
assign c0222 =  x544 &  x622;
assign c0224 =  x379 & ~x183 & ~x271 & ~x272 & ~x673;
assign c0226 =  x27;
assign c0228 =  x111;
assign c0230 =  x489 &  x516 &  x539 &  x566 & ~x395 & ~x713 & ~x774;
assign c0232 =  x227 &  x534 & ~x318;
assign c0234 =  x0;
assign c0236 =  x534 & ~x318 & ~x344 & ~x638;
assign c0238 =  x141;
assign c0240 =  x401 & ~x160 & ~x318 & ~x337 & ~x604 & ~x645 & ~x646 & ~x697 & ~x713 & ~x760;
assign c0242 = ~x14 & ~x145 & ~x158 & ~x242 & ~x328 & ~x410 & ~x413 & ~x414 & ~x711 & ~x770;
assign c0244 =  x480 & ~x275 & ~x330;
assign c0246 =  x55;
assign c0248 =  x147 & ~x15 & ~x155 & ~x196 & ~x296 & ~x308 & ~x354 & ~x574 & ~x616 & ~x640 & ~x672;
assign c0250 =  x389 & ~x155 & ~x216 & ~x236 & ~x289 & ~x318 & ~x551 & ~x705 & ~x730;
assign c0252 =  x544 &  x570 & ~x132 & ~x382 & ~x414 & ~x450;
assign c0254 =  x317 &  x567 &  x652 & ~x159;
assign c0256 =  x728;
assign c0258 =  x757;
assign c0260 =  x381 &  x409 &  x441 &  x464;
assign c0262 =  x261 &  x262 &  x345 &  x484 & ~x55 & ~x82 & ~x130 & ~x254 & ~x424 & ~x749;
assign c0264 =  x289 &  x540 &  x563 &  x568;
assign c0266 =  x783;
assign c0268 =  x550 &  x577 & ~x11 & ~x41 & ~x45 & ~x183 & ~x308 & ~x422 & ~x450 & ~x546 & ~x668 & ~x754;
assign c0270 =  x140;
assign c0272 =  x502 &  x530 &  x542;
assign c0274 =  x206 &  x318 &  x402 & ~x134 & ~x161 & ~x192 & ~x479 & ~x732 & ~x777;
assign c0276 =  x120 &  x148 &  x204 & ~x11 & ~x213 & ~x328 & ~x366 & ~x632;
assign c0278 =  x261 &  x262 &  x287 &  x512 &  x539 & ~x277 & ~x745;
assign c0280 =  x26;
assign c0282 =  x25;
assign c0284 =  x261 &  x289 & ~x13 & ~x99 & ~x153 & ~x215 & ~x243 & ~x421 & ~x423 & ~x687 & ~x776;
assign c0286 =  x503 &  x505;
assign c0288 =  x408 &  x438 &  x563 & ~x294;
assign c0290 =  x484 &  x547 & ~x515;
assign c0294 =  x167;
assign c0296 =  x226 & ~x18 & ~x143 & ~x319;
assign c0298 =  x120 &  x148 &  x176 & ~x74 & ~x240 & ~x576 & ~x704;
assign c0302 =  x559;
assign c0306 =  x206 &  x556 & ~x158 & ~x367 & ~x708;
assign c0308 =  x27;
assign c0310 =  x458 & ~x15 & ~x78 & ~x327 & ~x356 & ~x377 & ~x385 & ~x558 & ~x559 & ~x670 & ~x691 & ~x720 & ~x722 & ~x745;
assign c0312 =  x378 &  x436 & ~x150 & ~x488 & ~x638 & ~x662;
assign c0314 =  x459 &  x550 &  x577 & ~x10 & ~x16 & ~x33 & ~x43 & ~x103 & ~x449 & ~x643 & ~x690 & ~x722 & ~x735 & ~x775;
assign c0316 =  x522 &  x549 &  x577 &  x604 & ~x421;
assign c0318 =  x172 &  x201 &  x451 & ~x6 & ~x46 & ~x328 & ~x613 & ~x673 & ~x712 & ~x717 & ~x743;
assign c0320 =  x83;
assign c0322 = ~x11 & ~x75 & ~x88 & ~x155 & ~x187 & ~x212 & ~x327 & ~x465 & ~x680 & ~x686;
assign c0324 =  x230 &  x436 &  x510 &  x536 & ~x94 & ~x123 & ~x150 & ~x675;
assign c0326 =  x479 & ~x94 & ~x150 & ~x243 & ~x289;
assign c0328 =  x55;
assign c0330 =  x121 &  x291 &  x318 &  x402 & ~x242 & ~x325;
assign c0332 =  x333 &  x401 &  x426 &  x480 & ~x319 & ~x586;
assign c0334 =  x597 &  x622 &  x624 & ~x9;
assign c0336 =  x401 &  x480 & ~x42 & ~x217 & ~x551 & ~x580;
assign c0338 =  x510 &  x518 & ~x421;
assign c0340 =  x483 & ~x190 & ~x225 & ~x270 & ~x299 & ~x380 & ~x384 & ~x411;
assign c0342 =  x261 &  x318 &  x345 &  x457 & ~x33 & ~x44 & ~x113 & ~x125 & ~x135 & ~x183;
assign c0344 = ~x13 & ~x32 & ~x39 & ~x54 & ~x94 & ~x122 & ~x129 & ~x271 & ~x500 & ~x519 & ~x551 & ~x557 & ~x579 & ~x607 & ~x620 & ~x624 & ~x638 & ~x646 & ~x672 & ~x719 & ~x763 & ~x768;
assign c0346 = ~x39 & ~x192 & ~x240 & ~x275 & ~x328 & ~x352 & ~x356 & ~x474 & ~x560 & ~x717 & ~x740 & ~x752;
assign c0348 = ~x17 & ~x35 & ~x71 & ~x72 & ~x77 & ~x97 & ~x105 & ~x132 & ~x137 & ~x212 & ~x298 & ~x327 & ~x328 & ~x330 & ~x336 & ~x379 & ~x383 & ~x435 & ~x611 & ~x617 & ~x693 & ~x731 & ~x779;
assign c0350 =  x556 &  x610 & ~x12 & ~x303 & ~x697;
assign c0352 =  x28;
assign c0354 =  x544 &  x570 & ~x37 & ~x53 & ~x78 & ~x102 & ~x111 & ~x130 & ~x356 & ~x736;
assign c0356 =  x594 & ~x39 & ~x270 & ~x298 & ~x363 & ~x414 & ~x457 & ~x682;
assign c0358 =  x278 &  x377;
assign c0360 =  x118 &  x147 &  x172 &  x480 & ~x708;
assign c0362 = ~x153 & ~x187 & ~x206 & ~x243 & ~x266 & ~x318 & ~x357 & ~x601 & ~x671 & ~x683 & ~x705 & ~x779;
assign c0364 =  x232 &  x260 &  x427 & ~x375 & ~x576;
assign c0366 =  x783;
assign c0368 =  x332 &  x441 & ~x181;
assign c0370 =  x144 &  x174 &  x425 & ~x338;
assign c0372 =  x459 &  x519 &  x599;
assign c0374 =  x232 &  x427 &  x483 &  x595 &  x623 & ~x1 & ~x319 & ~x731;
assign c0376 =  x26;
assign c0378 =  x106;
assign c0380 =  x113 &  x341 &  x480;
assign c0382 =  x204 &  x457 & ~x10 & ~x69 & ~x152 & ~x236 & ~x269 & ~x640 & ~x642 & ~x719;
assign c0384 =  x234 &  x262 &  x595 & ~x101 & ~x699 & ~x773;
assign c0386 =  x544 &  x596 & ~x4 & ~x11 & ~x105 & ~x134;
assign c0388 =  x617;
assign c0390 =  x480 &  x567 & ~x153 & ~x212 & ~x614;
assign c0392 =  x540 & ~x265 & ~x266 & ~x327 & ~x351 & ~x664 & ~x686;
assign c0394 =  x489 & ~x106 & ~x130 & ~x144 & ~x356 & ~x379 & ~x560;
assign c0398 =  x83;
assign c0400 =  x147 &  x231 &  x506 & ~x125 & ~x694;
assign c0402 =  x261 &  x289 &  x317 &  x345 &  x513 & ~x155 & ~x395 & ~x719;
assign c0404 =  x379 &  x389 & ~x714 & ~x740;
assign c0406 =  x446 &  x510 &  x512 & ~x125 & ~x337 & ~x717;
assign c0408 =  x84;
assign c0410 =  x252;
assign c0412 =  x230 &  x480 &  x508 & ~x240 & ~x320 & ~x330 & ~x390;
assign c0414 =  x118 &  x119 &  x147 &  x174 &  x231 &  x370 & ~x598 & ~x703;
assign c0416 =  x540 & ~x189 & ~x408 & ~x548;
assign c0418 =  x147 &  x452 & ~x269 & ~x440;
assign c0420 =  x756;
assign c0422 =  x258 &  x313 &  x456 &  x507 &  x509 & ~x374 & ~x639 & ~x640 & ~x719 & ~x773;
assign c0426 =  x227 &  x479 & ~x159 & ~x366 & ~x580 & ~x692 & ~x775;
assign c0428 =  x32;
assign c0430 =  x204 &  x260 &  x316 &  x344 &  x484 &  x679;
assign c0432 = ~x16 & ~x38 & ~x57 & ~x101 & ~x267 & ~x269 & ~x270 & ~x318 & ~x328 & ~x332 & ~x334 & ~x420 & ~x434 & ~x660 & ~x666 & ~x710 & ~x719 & ~x722 & ~x737 & ~x773 & ~x777;
assign c0434 =  x34 &  x232 &  x372;
assign c0436 =  x54;
assign c0438 =  x261 &  x289 &  x317 & ~x47 & ~x55 & ~x240 & ~x269 & ~x367 & ~x395 & ~x492 & ~x643 & ~x775;
assign c0440 =  x232 &  x508 &  x510 & ~x181 & ~x318 & ~x691 & ~x745 & ~x781;
assign c0442 =  x480 & ~x20 & ~x47 & ~x56 & ~x65 & ~x93 & ~x98 & ~x184 & ~x266 & ~x290 & ~x298 & ~x328 & ~x393 & ~x688 & ~x754 & ~x759;
assign c0444 =  x23 &  x763;
assign c0446 =  x672;
assign c0448 =  x387 &  x548 & ~x394 & ~x420;
assign c0450 =  x397 &  x480 & ~x47 & ~x67 & ~x237 & ~x641;
assign c0454 =  x203 & ~x213 & ~x303 & ~x318 & ~x385 & ~x559 & ~x724;
assign c0456 =  x84;
assign c0458 =  x486 & ~x61 & ~x101 & ~x139 & ~x155 & ~x193 & ~x211 & ~x271 & ~x410 & ~x693;
assign c0460 =  x517 & ~x18 & ~x192 & ~x493;
assign c0462 =  x65 &  x93 &  x121 &  x205 &  x261 &  x344 & ~x575;
assign c0464 =  x399 & ~x11 & ~x187 & ~x318 & ~x320 & ~x421 & ~x557 & ~x638 & ~x689 & ~x710;
assign c0466 =  x204 &  x623 & ~x348 & ~x377 & ~x520;
assign c0468 =  x597 & ~x29 & ~x42 & ~x46 & ~x63 & ~x86 & ~x100 & ~x102 & ~x129 & ~x134 & ~x155 & ~x196 & ~x221 & ~x377 & ~x379 & ~x641 & ~x669 & ~x740 & ~x759 & ~x772;
assign c0470 =  x617 &  x620 &  x654;
assign c0472 =  x461 &  x475;
assign c0474 = ~x10 & ~x95 & ~x221 & ~x318 & ~x650;
assign c0476 =  x167;
assign c0478 =  x457 &  x547 & ~x328 & ~x466;
assign c0480 =  x521 &  x549 & ~x128 & ~x267 & ~x704;
assign c0482 =  x3;
assign c0484 =  x53;
assign c0486 =  x225 &  x285 &  x509;
assign c0488 =  x446 &  x457 &  x463 &  x537 & ~x424;
assign c0490 = ~x36 & ~x39 & ~x40 & ~x136 & ~x160 & ~x183 & ~x212 & ~x240 & ~x452 & ~x613 & ~x616 & ~x658 & ~x726 & ~x733 & ~x740 & ~x779;
assign c0492 =  x426 & ~x89 & ~x121 & ~x144 & ~x187 & ~x217 & ~x271 & ~x272 & ~x290 & ~x579 & ~x654 & ~x718;
assign c0494 =  x112;
assign c0496 =  x55;
assign c0498 =  x509 & ~x39 & ~x129 & ~x289 & ~x294 & ~x324 & ~x356 & ~x450;
assign c01 =  x358 &  x359 &  x415 & ~x28 & ~x32 & ~x60 & ~x83 & ~x115 & ~x731 & ~x764;
assign c03 =  x276 &  x304 & ~x95 & ~x354 & ~x630;
assign c05 =  x675 & ~x418 & ~x543 & ~x657;
assign c07 = ~x12 & ~x23 & ~x29 & ~x369 & ~x418 & ~x425 & ~x445 & ~x498 & ~x507 & ~x536 & ~x558 & ~x563 & ~x617 & ~x701;
assign c09 = ~x54 & ~x209 & ~x332 & ~x335 & ~x339 & ~x418 & ~x441 & ~x499 & ~x528 & ~x534 & ~x611 & ~x640 & ~x735;
assign c011 =  x501 & ~x7 & ~x21 & ~x145 & ~x378 & ~x431 & ~x458 & ~x459 & ~x542 & ~x543 & ~x700;
assign c013 =  x228 &  x256 &  x311 &  x338;
assign c015 =  x181 &  x208 &  x235 &  x314;
assign c017 =  x534 & ~x0 & ~x57 & ~x133 & ~x142 & ~x432 & ~x435 & ~x543 & ~x783;
assign c019 =  x357 &  x385 &  x412 &  x413 &  x414 & ~x30;
assign c021 =  x619 &  x647 & ~x53 & ~x57 & ~x85 & ~x392 & ~x419 & ~x710 & ~x711 & ~x755;
assign c023 =  x407 &  x601 &  x628 &  x629 & ~x29 & ~x87 & ~x129 & ~x166 & ~x726 & ~x727;
assign c025 = ~x21 & ~x22 & ~x30 & ~x152 & ~x198 & ~x304 & ~x305 & ~x361 & ~x362 & ~x389 & ~x418 & ~x419 & ~x433 & ~x445 & ~x488 & ~x542 & ~x559 & ~x781;
assign c027 =  x661 &  x662 & ~x55 & ~x112 & ~x497 & ~x498 & ~x559 & ~x616 & ~x783;
assign c029 =  x649 &  x676 &  x677 & ~x23 & ~x253 & ~x448 & ~x531 & ~x684 & ~x685;
assign c031 =  x153 &  x154 &  x180 &  x181 &  x208;
assign c033 =  x182 &  x183 &  x209 & ~x58 & ~x765;
assign c035 =  x331 &  x359 & ~x461 & ~x518;
assign c037 = ~x4 & ~x5 & ~x35 & ~x107 & ~x112 & ~x113 & ~x322 & ~x351 & ~x409 & ~x433 & ~x459 & ~x486 & ~x543 & ~x598 & ~x635 & ~x683;
assign c039 = ~x90 & ~x402 & ~x431 & ~x438 & ~x459 & ~x594 & ~x710;
assign c041 = ~x83 & ~x92 & ~x96 & ~x121 & ~x137 & ~x160 & ~x174 & ~x201 & ~x202 & ~x228 & ~x229 & ~x283 & ~x284 & ~x626 & ~x759;
assign c043 =  x273 &  x302 &  x330 & ~x281 & ~x657;
assign c045 =  x245 &  x273 &  x301 & ~x82 & ~x83 & ~x109 & ~x466 & ~x756 & ~x763;
assign c047 = ~x21 & ~x31 & ~x64 & ~x86 & ~x117 & ~x138 & ~x141 & ~x172 & ~x174 & ~x202 & ~x228 & ~x229 & ~x257 & ~x284 & ~x311 & ~x339 & ~x605 & ~x615 & ~x711 & ~x726 & ~x727 & ~x763 & ~x767 & ~x782;
assign c049 =  x708 &  x709 & ~x455;
assign c051 = ~x83 & ~x343 & ~x370 & ~x371 & ~x549 & ~x608 & ~x644 & ~x783;
assign c053 =  x69 &  x97 &  x124 & ~x475 & ~x532 & ~x783;
assign c055 = ~x21 & ~x91 & ~x115 & ~x145 & ~x229 & ~x459 & ~x517 & ~x691;
assign c057 =  x369 & ~x90 & ~x105 & ~x143 & ~x171 & ~x402 & ~x459 & ~x770 & ~x783;
assign c059 =  x90 &  x650 & ~x51 & ~x81 & ~x480;
assign c061 = ~x140 & ~x171 & ~x204 & ~x232 & ~x259 & ~x260 & ~x433 & ~x616 & ~x630;
assign c063 = ~x96 & ~x343 & ~x370 & ~x371 & ~x425 & ~x498 & ~x507 & ~x526 & ~x702;
assign c065 =  x266 &  x267 &  x268 & ~x51 & ~x447 & ~x751;
assign c067 =  x619 &  x647 & ~x28 & ~x336 & ~x391 & ~x543 & ~x710 & ~x775;
assign c069 =  x659 & ~x362 & ~x445 & ~x472 & ~x529 & ~x698;
assign c071 =  x219 &  x248 &  x249 & ~x112 & ~x494 & ~x710;
assign c073 =  x295 &  x322 &  x323 &  x403;
assign c075 =  x181 &  x208 &  x209 &  x236 & ~x34 & ~x62 & ~x168 & ~x224 & ~x559 & ~x587 & ~x675 & ~x703 & ~x761;
assign c077 = ~x238 & ~x399 & ~x400 & ~x402 & ~x427 & ~x455 & ~x456 & ~x482 & ~x503 & ~x510 & ~x511 & ~x538 & ~x539 & ~x559;
assign c079 = ~x239 & ~x361 & ~x389 & ~x441 & ~x444 & ~x445 & ~x480 & ~x497 & ~x536 & ~x733 & ~x783;
assign c081 = ~x368 & ~x395 & ~x453 & ~x480 & ~x481 & ~x507 & ~x509 & ~x534 & ~x536 & ~x537 & ~x563 & ~x564 & ~x581 & ~x593 & ~x649 & ~x706 & ~x763;
assign c083 = ~x22 & ~x75 & ~x181 & ~x333 & ~x339 & ~x360 & ~x362 & ~x393 & ~x420 & ~x445 & ~x447 & ~x536 & ~x564 & ~x584 & ~x783;
assign c085 = ~x50 & ~x60 & ~x79 & ~x103 & ~x220 & ~x247 & ~x305 & ~x418 & ~x445 & ~x447 & ~x573 & ~x584;
assign c087 =  x657 &  x658 & ~x72 & ~x498 & ~x524 & ~x530 & ~x549 & ~x587 & ~x670 & ~x727 & ~x753;
assign c089 = ~x24 & ~x48 & ~x86 & ~x117 & ~x408 & ~x459 & ~x460 & ~x462 & ~x596 & ~x655 & ~x681 & ~x716;
assign c091 =  x267 &  x294 & ~x331;
assign c093 =  x238 &  x265 &  x292 & ~x3 & ~x4 & ~x5 & ~x599 & ~x734;
assign c095 =  x297 & ~x17 & ~x29 & ~x279 & ~x314 & ~x504 & ~x531 & ~x733 & ~x762 & ~x763 & ~x766;
assign c097 = ~x62 & ~x349 & ~x406 & ~x459 & ~x489 & ~x568 & ~x596 & ~x599 & ~x601 & ~x630 & ~x706 & ~x783;
assign c099 = ~x202 & ~x203 & ~x230 & ~x257 & ~x259 & ~x286 & ~x313 & ~x314;
assign c0101 = ~x50 & ~x147 & ~x223 & ~x295 & ~x337 & ~x433 & ~x459 & ~x514 & ~x771;
assign c0103 =  x157 &  x158 & ~x25 & ~x58 & ~x112 & ~x142 & ~x143 & ~x196 & ~x197 & ~x491 & ~x710 & ~x748 & ~x755 & ~x765;
assign c0105 = ~x21 & ~x79 & ~x193 & ~x201 & ~x202 & ~x229 & ~x433 & ~x459;
assign c0107 = ~x19 & ~x54 & ~x287 & ~x288 & ~x314 & ~x342 & ~x343 & ~x370 & ~x616 & ~x772 & ~x775;
assign c0109 =  x157 &  x158 & ~x21 & ~x59 & ~x61 & ~x68 & ~x281;
assign c0111 = ~x21 & ~x53 & ~x201 & ~x229 & ~x257 & ~x284 & ~x307 & ~x332 & ~x333 & ~x418 & ~x529 & ~x587;
assign c0113 =  x236 &  x240 &  x268 & ~x40;
assign c0115 =  x580 &  x581 & ~x509 & ~x537;
assign c0117 =  x659 &  x687 &  x688 &  x689 & ~x57 & ~x531;
assign c0119 =  x274 &  x358 & ~x407 & ~x574;
assign c0121 =  x708 &  x711 &  x739;
assign c0123 = ~x336 & ~x371 & ~x399 & ~x401 & ~x402 & ~x455 & ~x531 & ~x537 & ~x727 & ~x783;
assign c0125 =  x67 &  x68 & ~x23 & ~x51 & ~x445 & ~x528;
assign c0127 =  x428 & ~x90 & ~x174 & ~x201 & ~x202 & ~x229 & ~x257 & ~x258 & ~x285 & ~x313;
assign c0129 =  x268 &  x269 &  x295 &  x296 &  x430;
assign c0131 =  x682 &  x683 & ~x0 & ~x2 & ~x55 & ~x83 & ~x109 & ~x167 & ~x221 & ~x245 & ~x418 & ~x478 & ~x531 & ~x534 & ~x586 & ~x588 & ~x617 & ~x646 & ~x701 & ~x759;
assign c0133 =  x276 &  x304 &  x445 &  x501;
assign c0135 = ~x0 & ~x21 & ~x22 & ~x103 & ~x208 & ~x223 & ~x226 & ~x276 & ~x305 & ~x332 & ~x335 & ~x362 & ~x418 & ~x445 & ~x526 & ~x664;
assign c0137 =  x238 & ~x360 & ~x445 & ~x459;
assign c0139 =  x695 & ~x196 & ~x419 & ~x503 & ~x783;
assign c0141 =  x360 & ~x92 & ~x171 & ~x173 & ~x201 & ~x202 & ~x225 & ~x284 & ~x308;
assign c0143 =  x211 &  x239 & ~x27 & ~x260 & ~x335 & ~x710 & ~x783;
assign c0145 = ~x91 & ~x92 & ~x142 & ~x280 & ~x408 & ~x512 & ~x513 & ~x599 & ~x634 & ~x652 & ~x732;
assign c0147 = ~x24 & ~x60 & ~x169 & ~x336 & ~x353 & ~x374 & ~x402 & ~x429 & ~x431 & ~x456 & ~x458 & ~x484 & ~x511 & ~x703 & ~x729 & ~x779;
assign c0149 = ~x2 & ~x14 & ~x17 & ~x53 & ~x167 & ~x169 & ~x170 & ~x248 & ~x273 & ~x279 & ~x280 & ~x302 & ~x305 & ~x360 & ~x362 & ~x389 & ~x418 & ~x445 & ~x474 & ~x498 & ~x503 & ~x531 & ~x589 & ~x748;
assign c0151 =  x212 &  x213 &  x240 &  x241 & ~x28 & ~x225 & ~x710;
assign c0153 =  x180 &  x423 & ~x763;
assign c0155 =  x738 &  x739;
assign c0157 =  x407 & ~x86 & ~x399 & ~x455 & ~x482 & ~x510;
assign c0159 = ~x50 & ~x180 & ~x343 & ~x370 & ~x371 & ~x372 & ~x399 & ~x503 & ~x765;
assign c0161 =  x405 &  x406 & ~x280 & ~x361 & ~x418 & ~x534 & ~x644 & ~x697;
assign c0163 =  x244 &  x329 & ~x418;
assign c0165 =  x659 &  x687 &  x688 &  x689 & ~x23 & ~x56 & ~x281 & ~x447 & ~x559;
assign c0167 =  x269 &  x295 & ~x767;
assign c0169 = ~x180 & ~x232 & ~x278 & ~x307 & ~x332 & ~x445 & ~x472 & ~x505 & ~x561;
assign c0171 =  x208 &  x209 &  x342;
assign c0173 =  x124 &  x125 &  x151 &  x179 & ~x3 & ~x60 & ~x280 & ~x781 & ~x783;
assign c0175 =  x453 & ~x18 & ~x93 & ~x267 & ~x383 & ~x458 & ~x543 & ~x652 & ~x688 & ~x709 & ~x733;
assign c0177 =  x334 & ~x57 & ~x350 & ~x484 & ~x538 & ~x540 & ~x710;
assign c0179 =  x648 &  x675 &  x703 & ~x96 & ~x140 & ~x167 & ~x168 & ~x738;
assign c0181 = ~x90 & ~x92 & ~x174 & ~x201 & ~x202 & ~x225 & ~x229 & ~x230 & ~x257 & ~x285 & ~x311 & ~x312 & ~x727;
assign c0183 = ~x33 & ~x83 & ~x122 & ~x151 & ~x349 & ~x378 & ~x404 & ~x410 & ~x460 & ~x514 & ~x568 & ~x599 & ~x659 & ~x710;
assign c0185 =  x209 &  x210 & ~x55 & ~x169 & ~x503 & ~x671;
assign c0187 =  x435 & ~x40 & ~x129 & ~x454 & ~x504 & ~x509 & ~x536 & ~x537 & ~x620 & ~x754 & ~x781;
assign c0189 = ~x0 & ~x63 & ~x135 & ~x168 & ~x174 & ~x351 & ~x402 & ~x459 & ~x625 & ~x628 & ~x674 & ~x680 & ~x762;
assign c0191 =  x276 &  x417 & ~x353 & ~x459;
assign c0193 =  x416 & ~x33 & ~x187 & ~x455 & ~x482 & ~x484 & ~x511 & ~x537 & ~x594 & ~x700 & ~x783;
assign c0195 = ~x19 & ~x425 & ~x453 & ~x454 & ~x455 & ~x481 & ~x482 & ~x509 & ~x510 & ~x536 & ~x537 & ~x621 & ~x635 & ~x747 & ~x774;
assign c0197 =  x405 &  x490 & ~x0 & ~x418 & ~x445;
assign c0199 = ~x201 & ~x458 & ~x486 & ~x518 & ~x573 & ~x596 & ~x783;
assign c0201 =  x125 &  x152 & ~x30 & ~x112 & ~x308 & ~x692 & ~x775 & ~x777;
assign c0203 =  x710 &  x711 &  x712 & ~x418;
assign c0205 =  x185 &  x212 & ~x22 & ~x57 & ~x202;
assign c0207 =  x428 &  x510 &  x590 & ~x406 & ~x433;
assign c0209 =  x209 &  x236 & ~x57 & ~x165 & ~x197 & ~x224 & ~x652;
assign c0211 = ~x43 & ~x131 & ~x332 & ~x333 & ~x402 & ~x503 & ~x540 & ~x587;
assign c0213 =  x554 &  x583 & ~x445;
assign c0215 =  x240 & ~x445;
assign c0217 = ~x99 & ~x103 & ~x158 & ~x425 & ~x453 & ~x507 & ~x509 & ~x534 & ~x536 & ~x537 & ~x538 & ~x565 & ~x594 & ~x638 & ~x646 & ~x754;
assign c0219 =  x90 & ~x342 & ~x343;
assign c0221 = ~x237 & ~x263 & ~x369 & ~x453 & ~x480 & ~x509 & ~x536 & ~x537;
assign c0223 =  x304 & ~x13 & ~x88 & ~x147 & ~x597 & ~x627 & ~x657 & ~x709 & ~x734 & ~x754 & ~x756 & ~x757 & ~x762 & ~x764;
assign c0225 = ~x57 & ~x79 & ~x117 & ~x133 & ~x191 & ~x200 & ~x201 & ~x229 & ~x282 & ~x305 & ~x361 & ~x363 & ~x418 & ~x419 & ~x445 & ~x559;
assign c0227 = ~x30 & ~x166 & ~x254 & ~x282 & ~x305 & ~x332 & ~x418 & ~x445 & ~x450 & ~x479 & ~x499 & ~x531 & ~x563 & ~x669 & ~x700 & ~x729 & ~x775;
assign c0229 =  x212 &  x239 &  x240 &  x267 & ~x782;
assign c0231 = ~x43 & ~x183 & ~x396 & ~x453 & ~x454 & ~x480 & ~x481 & ~x507 & ~x508 & ~x509 & ~x510 & ~x532 & ~x535 & ~x537 & ~x559 & ~x565 & ~x612 & ~x642 & ~x644 & ~x722 & ~x728 & ~x731 & ~x775;
assign c0233 =  x748;
assign c0235 =  x647 &  x675 & ~x21 & ~x57 & ~x97 & ~x197 & ~x632 & ~x683;
assign c0237 = ~x21 & ~x86 & ~x114 & ~x142 & ~x226 & ~x402 & ~x429 & ~x431 & ~x456 & ~x484 & ~x511;
assign c0239 =  x181 &  x182 &  x208 & ~x504;
assign c0241 =  x303 & ~x204 & ~x599 & ~x656;
assign c0243 =  x405 & ~x3 & ~x26 & ~x30 & ~x103 & ~x498 & ~x499 & ~x504 & ~x506 & ~x529 & ~x536 & ~x759;
assign c0245 =  x183 &  x184 &  x210 &  x428;
assign c0247 =  x298 &  x326 &  x354 & ~x83 & ~x361 & ~x418 & ~x419 & ~x443 & ~x445;
assign c0249 =  x209 &  x210 &  x211 & ~x144 & ~x652;
assign c0251 =  x619 &  x646 &  x647 &  x674 & ~x710;
assign c0253 =  x208 &  x366;
assign c0255 =  x465 & ~x134 & ~x218 & ~x332 & ~x335 & ~x359 & ~x418 & ~x459 & ~x499;
assign c0257 = ~x24 & ~x83 & ~x90 & ~x257 & ~x285 & ~x553 & ~x573 & ~x749;
assign c0259 =  x342 & ~x16 & ~x31 & ~x45 & ~x108 & ~x115 & ~x142 & ~x143 & ~x170 & ~x197 & ~x227 & ~x276 & ~x305 & ~x337 & ~x418 & ~x445 & ~x562 & ~x726 & ~x728;
assign c0261 =  x97 &  x124 &  x125 &  x179 & ~x196;
assign c0263 =  x283 &  x310 &  x338 &  x366;
assign c0265 = ~x53 & ~x399 & ~x400 & ~x426 & ~x454 & ~x455 & ~x456 & ~x509 & ~x511 & ~x537 & ~x621 & ~x777;
assign c0267 =  x255 &  x311 &  x338 &  x339;
assign c0269 = ~x24 & ~x40 & ~x83 & ~x147 & ~x402 & ~x408 & ~x431 & ~x459 & ~x541 & ~x707 & ~x757;
assign c0271 =  x437 & ~x28 & ~x87 & ~x167 & ~x222 & ~x248 & ~x251 & ~x306 & ~x308 & ~x418 & ~x469 & ~x497 & ~x504 & ~x558 & ~x586;
assign c0273 =  x265 &  x266 &  x292 & ~x625 & ~x682;
assign c0275 =  x245 &  x273 & ~x44 & ~x59 & ~x434 & ~x476 & ~x494 & ~x725 & ~x783;
assign c0277 =  x407 & ~x251 & ~x253 & ~x279 & ~x282 & ~x305 & ~x310 & ~x332 & ~x361 & ~x362 & ~x418 & ~x445 & ~x533 & ~x586;
assign c0279 =  x299 &  x326 &  x327 &  x429 & ~x475;
assign c0281 = ~x28 & ~x55 & ~x62 & ~x72 & ~x87 & ~x92 & ~x114 & ~x174 & ~x196 & ~x201 & ~x202 & ~x229 & ~x251 & ~x257 & ~x284 & ~x339 & ~x684;
assign c0283 = ~x2 & ~x83 & ~x234 & ~x369 & ~x398 & ~x399 & ~x479 & ~x480 & ~x532;
assign c0285 =  x294 &  x295 &  x322 &  x323 & ~x3 & ~x28 & ~x165 & ~x170 & ~x197 & ~x503 & ~x559 & ~x759;
assign c0287 =  x268 &  x269 & ~x23 & ~x146 & ~x201;
assign c0289 =  x342 & ~x21 & ~x112 & ~x305 & ~x307 & ~x332 & ~x339 & ~x366 & ~x418 & ~x445 & ~x503 & ~x528 & ~x771;
assign c0291 =  x627 &  x683 & ~x81 & ~x418 & ~x557;
assign c0293 =  x187 & ~x1 & ~x7 & ~x435 & ~x521 & ~x598 & ~x754 & ~x757 & ~x766;
assign c0295 =  x124 &  x125 &  x151 &  x152 & ~x56 & ~x82 & ~x475 & ~x530 & ~x556 & ~x652;
assign c0297 = ~x167 & ~x192 & ~x201 & ~x228 & ~x385 & ~x418 & ~x445 & ~x524;
assign c0299 = ~x52 & ~x96 & ~x117 & ~x137 & ~x138 & ~x145 & ~x147 & ~x170 & ~x195 & ~x284 & ~x339 & ~x410 & ~x669 & ~x739 & ~x752 & ~x757 & ~x782;
assign c0301 =  x301 &  x329 &  x593 & ~x489;
assign c0303 = ~x2 & ~x20 & ~x23 & ~x57 & ~x59 & ~x60 & ~x150 & ~x249 & ~x252 & ~x279 & ~x335 & ~x391 & ~x419 & ~x459 & ~x514 & ~x597 & ~x652 & ~x762 & ~x763;
assign c0305 = ~x5 & ~x8 & ~x19 & ~x26 & ~x55 & ~x82 & ~x253 & ~x333 & ~x358 & ~x387 & ~x418 & ~x445 & ~x447 & ~x507 & ~x524 & ~x529 & ~x535 & ~x753 & ~x783;
assign c0307 =  x229 & ~x98 & ~x112 & ~x426 & ~x453 & ~x509 & ~x510 & ~x565;
assign c0309 =  x324 & ~x4 & ~x98 & ~x305 & ~x336 & ~x361 & ~x391 & ~x418 & ~x445 & ~x474;
assign c0311 =  x744 &  x745 &  x746 & ~x280 & ~x672;
assign c0313 =  x564 & ~x109 & ~x139 & ~x196 & ~x222 & ~x324 & ~x404 & ~x459 & ~x514 & ~x627 & ~x659 & ~x710;
assign c0315 = ~x95 & ~x98 & ~x150 & ~x178 & ~x204 & ~x232 & ~x432 & ~x433 & ~x543 & ~x573 & ~x599 & ~x629 & ~x687 & ~x710 & ~x712 & ~x736 & ~x759;
assign c0317 =  x239 &  x266 & ~x251 & ~x362 & ~x391 & ~x503;
assign c0319 = ~x23 & ~x180 & ~x398 & ~x418 & ~x445 & ~x506 & ~x528 & ~x533 & ~x534 & ~x557;
assign c0321 = ~x57 & ~x285 & ~x286 & ~x287 & ~x313 & ~x314 & ~x342 & ~x343 & ~x370;
assign c0323 = ~x177 & ~x258 & ~x285 & ~x286 & ~x314 & ~x341;
assign c0325 = ~x369 & ~x453 & ~x454 & ~x482 & ~x507 & ~x509 & ~x510 & ~x536 & ~x537 & ~x767;
assign c0327 =  x399 & ~x23 & ~x202 & ~x229 & ~x257 & ~x284 & ~x782;
assign c0329 =  x360 &  x500 & ~x30 & ~x33 & ~x83 & ~x174 & ~x504;
assign c0331 = ~x237 & ~x343 & ~x371 & ~x399 & ~x454 & ~x510;
assign c0333 =  x247 & ~x148 & ~x524 & ~x783;
assign c0335 = ~x0 & ~x2 & ~x300 & ~x354 & ~x402 & ~x486 & ~x568 & ~x593 & ~x597;
assign c0337 =  x40 &  x94 & ~x23 & ~x26 & ~x249 & ~x476;
assign c0339 =  x210 &  x211 &  x236 &  x237 &  x369 & ~x196;
assign c0341 =  x487 & ~x453 & ~x481 & ~x509 & ~x536 & ~x537 & ~x580 & ~x593;
assign c0343 = ~x0 & ~x25 & ~x28 & ~x53 & ~x181 & ~x196 & ~x280 & ~x314 & ~x341 & ~x342 & ~x368 & ~x369 & ~x452 & ~x587 & ~x670 & ~x763 & ~x777;
assign c0345 =  x294 & ~x28 & ~x30 & ~x54 & ~x280 & ~x305 & ~x330 & ~x360 & ~x389 & ~x418 & ~x446 & ~x475 & ~x529;
assign c0347 = ~x6 & ~x12 & ~x55 & ~x107 & ~x112 & ~x431 & ~x438 & ~x571 & ~x595 & ~x631 & ~x732;
assign c0349 =  x370 &  x507 & ~x18 & ~x64 & ~x78 & ~x81 & ~x114 & ~x459 & ~x515 & ~x627 & ~x702 & ~x754;
assign c0351 = ~x148 & ~x201 & ~x202 & ~x203 & ~x229 & ~x258 & ~x311 & ~x681;
assign c0353 =  x658 &  x659 &  x687 & ~x53 & ~x445 & ~x447 & ~x473 & ~x502 & ~x530 & ~x646 & ~x702 & ~x732;
assign c0355 =  x249 &  x334 & ~x408 & ~x711 & ~x762;
assign c0357 =  x462 & ~x26 & ~x53 & ~x160 & ~x210 & ~x419 & ~x481 & ~x507 & ~x509 & ~x620;
assign c0359 =  x228 & ~x398 & ~x425 & ~x452 & ~x454 & ~x508;
assign c0361 = ~x300 & ~x373 & ~x402 & ~x459 & ~x484 & ~x511 & ~x538;
assign c0363 = ~x24 & ~x346 & ~x454 & ~x481 & ~x482 & ~x509 & ~x510 & ~x537 & ~x635;
assign c0365 = ~x18 & ~x19 & ~x21 & ~x22 & ~x79 & ~x83 & ~x89 & ~x91 & ~x118 & ~x145 & ~x147 & ~x202 & ~x224 & ~x228 & ~x229 & ~x596 & ~x615 & ~x682 & ~x700 & ~x705;
assign c0367 =  x228 &  x255 &  x311 & ~x27 & ~x111 & ~x139 & ~x729;
assign c0369 = ~x51 & ~x57 & ~x108 & ~x197 & ~x220 & ~x221 & ~x305 & ~x329 & ~x332 & ~x335 & ~x362 & ~x418 & ~x477 & ~x498 & ~x529 & ~x587;
assign c0371 =  x245 &  x273 & ~x22 & ~x445;
assign c0373 =  x297 & ~x24 & ~x305 & ~x332 & ~x387 & ~x418 & ~x445 & ~x472 & ~x503 & ~x690 & ~x755 & ~x782;
assign c0375 =  x41 & ~x105 & ~x143 & ~x778;
assign c0377 =  x301 &  x329 &  x330 & ~x84 & ~x174 & ~x710 & ~x756;
assign c0379 =  x127 &  x154 & ~x59 & ~x82 & ~x141 & ~x642;
assign c0381 =  x264 &  x265 &  x292 &  x425 & ~x193;
assign c0383 =  x334 &  x417 &  x418 & ~x10 & ~x84 & ~x88 & ~x174 & ~x196 & ~x201 & ~x655 & ~x678 & ~x706 & ~x708 & ~x733;
assign c0385 =  x240 &  x241;
assign c0387 = ~x5 & ~x98 & ~x247 & ~x305 & ~x311 & ~x332 & ~x335 & ~x339 & ~x362 & ~x498 & ~x506 & ~x530 & ~x589 & ~x641 & ~x783;
assign c0389 = ~x55 & ~x72 & ~x85 & ~x139 & ~x220 & ~x339 & ~x361 & ~x418 & ~x445 & ~x471 & ~x495 & ~x506 & ~x562 & ~x702;
assign c0391 =  x302 &  x330 & ~x60 & ~x310 & ~x543;
assign c0393 = ~x16 & ~x19 & ~x41 & ~x114 & ~x319 & ~x454 & ~x455 & ~x477 & ~x482 & ~x507 & ~x509 & ~x510 & ~x536 & ~x537 & ~x538 & ~x561 & ~x564 & ~x565 & ~x593 & ~x639 & ~x644 & ~x750 & ~x770;
assign c0395 =  x407 & ~x2 & ~x26 & ~x28 & ~x167 & ~x250 & ~x418 & ~x445 & ~x475 & ~x614 & ~x616 & ~x694;
assign c0397 = ~x13 & ~x23 & ~x263 & ~x280 & ~x370 & ~x399 & ~x421 & ~x452 & ~x453 & ~x756 & ~x782;
assign c0399 =  x714 & ~x83 & ~x280 & ~x473 & ~x524 & ~x534 & ~x587 & ~x589 & ~x728;
assign c0401 =  x237 &  x240;
assign c0403 =  x314 & ~x7 & ~x9 & ~x35 & ~x59 & ~x105 & ~x459 & ~x464 & ~x486 & ~x541 & ~x568 & ~x571 & ~x597 & ~x601 & ~x667;
assign c0405 =  x434 & ~x79 & ~x453 & ~x455 & ~x482 & ~x509 & ~x537 & ~x538 & ~x593 & ~x620 & ~x741;
assign c0407 =  x668 & ~x531;
assign c0409 = ~x40 & ~x169 & ~x171 & ~x364 & ~x401 & ~x402 & ~x431 & ~x456 & ~x484 & ~x511 & ~x538 & ~x676 & ~x749;
assign c0411 =  x331 &  x359 &  x528 & ~x167;
assign c0413 =  x434 & ~x399 & ~x454 & ~x455 & ~x481;
assign c0415 = ~x5 & ~x6 & ~x33 & ~x86 & ~x102 & ~x107 & ~x173 & ~x308 & ~x322 & ~x431 & ~x459 & ~x571 & ~x627 & ~x655 & ~x708 & ~x727 & ~x761 & ~x783;
assign c0417 =  x240 &  x242 &  x267 & ~x35;
assign c0419 =  x266 &  x293 &  x294 & ~x655 & ~x656;
assign c0421 =  x380 & ~x251 & ~x331 & ~x332 & ~x334 & ~x418 & ~x445 & ~x497;
assign c0423 =  x338 &  x366 &  x393 &  x394 & ~x19 & ~x33;
assign c0425 =  x369 &  x423 & ~x79 & ~x86 & ~x107 & ~x197 & ~x201 & ~x228 & ~x587;
assign c0427 = ~x79 & ~x197 & ~x418 & ~x422 & ~x445 & ~x475 & ~x496 & ~x498 & ~x532 & ~x534 & ~x554 & ~x587 & ~x617 & ~x759 & ~x777 & ~x783;
assign c0429 = ~x20 & ~x23 & ~x57 & ~x111 & ~x426 & ~x453 & ~x480 & ~x481 & ~x507 & ~x508 & ~x509 & ~x536 & ~x557 & ~x562 & ~x580 & ~x642 & ~x727 & ~x771;
assign c0431 =  x329 & ~x3 & ~x6 & ~x17 & ~x60 & ~x207 & ~x280 & ~x462 & ~x476 & ~x549 & ~x751 & ~x783;
assign c0433 =  x268 &  x295 & ~x230;
assign c0435 =  x154 &  x180 &  x181 &  x207 &  x208 & ~x108;
assign c0437 =  x238 &  x265 &  x292 &  x293 & ~x625 & ~x681 & ~x742;
assign c0439 =  x369 & ~x18 & ~x21 & ~x51 & ~x57 & ~x85 & ~x138 & ~x144 & ~x198 & ~x200 & ~x223 & ~x249 & ~x276 & ~x280 & ~x305 & ~x336 & ~x362 & ~x416 & ~x417 & ~x418 & ~x587 & ~x615 & ~x756;
assign c0441 = ~x8 & ~x61 & ~x120 & ~x133 & ~x139 & ~x381 & ~x432 & ~x459 & ~x462 & ~x541 & ~x568 & ~x573 & ~x597 & ~x630 & ~x706 & ~x735;
assign c0443 =  x722 & ~x527;
assign c0445 = ~x218 & ~x370 & ~x398 & ~x399 & ~x454 & ~x536 & ~x549;
assign c0447 = ~x2 & ~x28 & ~x201 & ~x202 & ~x257 & ~x284 & ~x285 & ~x313 & ~x339 & ~x475 & ~x549;
assign c0449 = ~x131 & ~x237 & ~x399 & ~x455 & ~x509 & ~x510 & ~x511 & ~x537 & ~x538;
assign c0451 = ~x79 & ~x177 & ~x179 & ~x204 & ~x232 & ~x279 & ~x338 & ~x433 & ~x736;
assign c0453 = ~x15 & ~x18 & ~x33 & ~x51 & ~x54 & ~x81 & ~x83 & ~x108 & ~x132 & ~x193 & ~x221 & ~x226 & ~x227 & ~x248 & ~x253 & ~x339 & ~x363 & ~x418 & ~x420 & ~x421 & ~x445 & ~x447 & ~x585 & ~x764 & ~x782;
assign c0455 =  x97 &  x98 &  x124 &  x125;
assign c0457 =  x334 & ~x15 & ~x511 & ~x537 & ~x538 & ~x597;
assign c0459 =  x310 & ~x507 & ~x536;
assign c0461 =  x323 & ~x83 & ~x96 & ~x153 & ~x279 & ~x305 & ~x332 & ~x362 & ~x418 & ~x587 & ~x726 & ~x770 & ~x776;
assign c0463 =  x154 &  x155 &  x181 &  x182 &  x208 & ~x167;
assign c0465 =  x256 &  x311 & ~x83 & ~x84 & ~x195 & ~x481 & ~x509 & ~x537 & ~x589 & ~x615 & ~x616 & ~x766;
assign c0467 =  x213 &  x214 & ~x335 & ~x418 & ~x445;
assign c0469 =  x13;
assign c0471 =  x286 &  x314 & ~x51 & ~x171 & ~x193 & ~x196 & ~x222 & ~x227 & ~x251 & ~x304 & ~x305 & ~x335 & ~x362 & ~x418 & ~x419 & ~x445 & ~x472 & ~x475 & ~x529 & ~x534;
assign c0473 =  x219 &  x275 & ~x461 & ~x543;
assign c0475 =  x238 &  x239 &  x266 &  x267 & ~x172 & ~x223 & ~x530;
assign c0477 =  x264 &  x268 & ~x691;
assign c0479 =  x299 &  x300 &  x325 & ~x21 & ~x43 & ~x74;
assign c0481 =  x311 &  x338 &  x365 &  x366;
assign c0483 =  x658 &  x659 &  x661 & ~x13 & ~x281 & ~x756;
assign c0485 =  x129 &  x156 &  x183 & ~x53 & ~x224 & ~x280;
assign c0487 =  x564 & ~x247 & ~x391 & ~x418 & ~x445 & ~x531 & ~x542 & ~x543 & ~x597 & ~x627;
assign c0489 =  x302 &  x330 &  x331 &  x358 & ~x22 & ~x32 & ~x109 & ~x767;
assign c0491 =  x187 &  x212;
assign c0493 =  x304 & ~x51 & ~x174 & ~x201 & ~x594 & ~x783;
assign c0495 = ~x6 & ~x81 & ~x114 & ~x143 & ~x402 & ~x411 & ~x430 & ~x431 & ~x441 & ~x459 & ~x469 & ~x513 & ~x540 & ~x699 & ~x732 & ~x764;
assign c0497 =  x12 &  x39;
assign c0499 = ~x53 & ~x86 & ~x196 & ~x203 & ~x230 & ~x409 & ~x412 & ~x632 & ~x688;
assign c10 =  x378 & ~x0 & ~x73 & ~x143 & ~x173 & ~x175 & ~x186 & ~x197 & ~x203 & ~x216 & ~x220 & ~x221 & ~x226 & ~x242 & ~x243 & ~x244 & ~x258 & ~x284 & ~x355 & ~x368 & ~x370 & ~x381 & ~x420 & ~x452 & ~x453 & ~x505 & ~x509 & ~x538 & ~x585 & ~x638 & ~x667 & ~x696 & ~x761 & ~x777 & ~x782;
assign c12 =  x322 &  x408 & ~x87 & ~x104 & ~x119 & ~x146 & ~x149 & ~x175 & ~x194 & ~x203 & ~x258 & ~x278 & ~x304 & ~x387 & ~x538 & ~x693 & ~x696 & ~x727;
assign c14 =  x626 &  x655 &  x684 & ~x371 & ~x600;
assign c16 =  x146 &  x646;
assign c18 =  x97 &  x211 &  x325 &  x353 & ~x87 & ~x257 & ~x338 & ~x342 & ~x722;
assign c110 = ~x73 & ~x188 & ~x248 & ~x249 & ~x258 & ~x260 & ~x370 & ~x402 & ~x404 & ~x473 & ~x498 & ~x636 & ~x699 & ~x704;
assign c112 = ~x7 & ~x24 & ~x86 & ~x104 & ~x111 & ~x120 & ~x138 & ~x144 & ~x146 & ~x148 & ~x170 & ~x173 & ~x176 & ~x188 & ~x202 & ~x203 & ~x204 & ~x224 & ~x230 & ~x232 & ~x233 & ~x249 & ~x260 & ~x261 & ~x287 & ~x288 & ~x304 & ~x315 & ~x317 & ~x332 & ~x333 & ~x337 & ~x367 & ~x373 & ~x396 & ~x397 & ~x401 & ~x453 & ~x454 & ~x500 & ~x512 & ~x557 & ~x587 & ~x618 & ~x672 & ~x718 & ~x728;
assign c114 =  x640;
assign c116 =  x37 &  x151 &  x294 & ~x397;
assign c118 =  x124 &  x322 & ~x121 & ~x538;
assign c120 =  x295 &  x324 &  x409 & ~x74 & ~x78 & ~x119 & ~x192 & ~x220 & ~x231 & ~x329 & ~x398 & ~x400 & ~x423 & ~x506 & ~x592 & ~x648 & ~x649 & ~x670 & ~x779;
assign c122 =  x580 &  x581 &  x585;
assign c124 =  x98 &  x241 &  x269 &  x298 & ~x394 & ~x406;
assign c126 =  x269 &  x384 &  x411 &  x743;
assign c128 = ~x82 & ~x176 & ~x204 & ~x229 & ~x288 & ~x375 & ~x402 & ~x406 & ~x604 & ~x676;
assign c130 =  x63 &  x675 & ~x97;
assign c132 =  x176 &  x233 &  x705;
assign c134 =  x411 & ~x76 & ~x82 & ~x115 & ~x141 & ~x258 & ~x395 & ~x434 & ~x454 & ~x637 & ~x723 & ~x724;
assign c136 =  x677 & ~x153 & ~x434 & ~x454;
assign c138 =  x663 & ~x578 & ~x771;
assign c140 = ~x95 & ~x97 & ~x126 & ~x155 & ~x290 & ~x388 & ~x736;
assign c142 =  x701;
assign c144 =  x634 & ~x73 & ~x658 & ~x744;
assign c146 =  x711 & ~x53 & ~x256 & ~x288 & ~x485 & ~x584 & ~x628 & ~x775;
assign c148 =  x405 &  x406 & ~x91 & ~x116 & ~x215 & ~x231 & ~x268 & ~x270 & ~x315 & ~x371 & ~x389 & ~x691;
assign c150 =  x608 &  x609 & ~x688 & ~x722;
assign c152 =  x241 &  x469 & ~x107 & ~x222 & ~x278 & ~x476 & ~x640 & ~x646 & ~x666 & ~x724;
assign c154 =  x551 & ~x54 & ~x58 & ~x79 & ~x110 & ~x187 & ~x314 & ~x388 & ~x453 & ~x504 & ~x531 & ~x661 & ~x666 & ~x692 & ~x697 & ~x750 & ~x782;
assign c156 =  x243 &  x483 & ~x306;
assign c158 =  x146 &  x483 & ~x467 & ~x624;
assign c160 =  x380 &  x408 &  x465 & ~x91 & ~x136 & ~x195 & ~x217 & ~x258 & ~x286 & ~x309 & ~x442 & ~x647 & ~x677 & ~x718 & ~x719 & ~x724;
assign c162 =  x0;
assign c164 =  x626 &  x655 &  x684 & ~x88 & ~x140 & ~x165 & ~x199 & ~x248 & ~x273 & ~x724 & ~x778;
assign c166 =  x325 & ~x73 & ~x120 & ~x261 & ~x406;
assign c168 = ~x4 & ~x27 & ~x31 & ~x72 & ~x88 & ~x108 & ~x134 & ~x162 & ~x168 & ~x175 & ~x222 & ~x228 & ~x232 & ~x272 & ~x273 & ~x286 & ~x344 & ~x399 & ~x419 & ~x473 & ~x505 & ~x526 & ~x553 & ~x574 & ~x647 & ~x665 & ~x666 & ~x675 & ~x692 & ~x695 & ~x696 & ~x722 & ~x725 & ~x730 & ~x748 & ~x754;
assign c170 =  x679 &  x706 & ~x480 & ~x584 & ~x629;
assign c172 =  x5 &  x6;
assign c174 =  x662 &  x664 & ~x773;
assign c176 =  x739 & ~x340 & ~x426 & ~x687 & ~x744 & ~x765;
assign c178 =  x731 & ~x322 & ~x516;
assign c180 =  x711 & ~x196 & ~x204 & ~x314 & ~x716;
assign c182 =  x325 &  x439 & ~x199 & ~x286 & ~x397 & ~x463 & ~x639 & ~x666 & ~x725;
assign c184 =  x231 &  x429 & ~x153 & ~x515;
assign c186 =  x636 &  x641;
assign c188 =  x435 &  x577 & ~x121 & ~x299;
assign c190 =  x324 & ~x7 & ~x92 & ~x106 & ~x142 & ~x143 & ~x193 & ~x260 & ~x278 & ~x375 & ~x661 & ~x692 & ~x720;
assign c192 =  x378 &  x436 &  x464 & ~x62 & ~x119 & ~x166 & ~x184 & ~x201 & ~x212 & ~x229 & ~x286 & ~x315 & ~x384 & ~x705;
assign c194 =  x455 & ~x150 & ~x296 & ~x377;
assign c196 =  x644;
assign c198 =  x655 & ~x121 & ~x212 & ~x341 & ~x372 & ~x398 & ~x412 & ~x424 & ~x667 & ~x691 & ~x722;
assign c1100 = ~x73 & ~x81 & ~x344 & ~x361 & ~x377 & ~x402 & ~x406 & ~x482 & ~x546;
assign c1102 =  x676 & ~x325 & ~x434;
assign c1104 = ~x47 & ~x51 & ~x112 & ~x116 & ~x133 & ~x149 & ~x173 & ~x176 & ~x199 & ~x244 & ~x253 & ~x258 & ~x259 & ~x275 & ~x288 & ~x304 & ~x331 & ~x361 & ~x367 & ~x370 & ~x402 & ~x418 & ~x475 & ~x556 & ~x584 & ~x619 & ~x662 & ~x677 & ~x703 & ~x706 & ~x718 & ~x722 & ~x733 & ~x757;
assign c1106 =  x351 &  x549 &  x655 & ~x258 & ~x691;
assign c1108 =  x605 & ~x83 & ~x159 & ~x164 & ~x229 & ~x242 & ~x251 & ~x270 & ~x282 & ~x297 & ~x306 & ~x315 & ~x382 & ~x422 & ~x453 & ~x471 & ~x496 & ~x675 & ~x691;
assign c1110 =  x119 &  x674;
assign c1112 = ~x3 & ~x49 & ~x63 & ~x115 & ~x140 & ~x196 & ~x197 & ~x203 & ~x231 & ~x260 & ~x304 & ~x317 & ~x334 & ~x364 & ~x399 & ~x427 & ~x429 & ~x430 & ~x447 & ~x473 & ~x501 & ~x584 & ~x605 & ~x691 & ~x692 & ~x693 & ~x719 & ~x780;
assign c1114 =  x324 &  x409 & ~x19 & ~x53 & ~x55 & ~x82 & ~x106 & ~x108 & ~x114 & ~x115 & ~x118 & ~x120 & ~x122 & ~x139 & ~x168 & ~x172 & ~x219 & ~x227 & ~x275 & ~x281 & ~x306 & ~x308 & ~x335 & ~x336 & ~x358 & ~x360 & ~x363 & ~x365 & ~x366 & ~x367 & ~x369 & ~x424 & ~x480 & ~x482 & ~x502 & ~x503 & ~x504 & ~x508 & ~x509 & ~x530 & ~x535 & ~x562 & ~x565 & ~x583 & ~x620 & ~x637 & ~x638 & ~x640 & ~x646 & ~x647 & ~x650 & ~x691 & ~x695 & ~x696 & ~x724 & ~x760;
assign c1116 =  x174 &  x674 & ~x241;
assign c1118 =  x623 &  x651 & ~x73 & ~x118 & ~x139 & ~x145 & ~x284 & ~x393 & ~x472 & ~x475 & ~x481 & ~x509 & ~x510 & ~x527 & ~x529 & ~x538 & ~x560 & ~x667 & ~x669 & ~x693 & ~x724 & ~x725 & ~x727 & ~x758;
assign c1120 = ~x34 & ~x60 & ~x141 & ~x147 & ~x156 & ~x188 & ~x210 & ~x220 & ~x229 & ~x242 & ~x259 & ~x304 & ~x325 & ~x329 & ~x383 & ~x415 & ~x482 & ~x722;
assign c1122 = ~x2 & ~x26 & ~x92 & ~x181 & ~x183 & ~x258 & ~x383 & ~x512 & ~x526 & ~x589 & ~x591 & ~x617 & ~x690 & ~x694 & ~x753;
assign c1124 =  x35 &  x648;
assign c1126 =  x326 &  x469 & ~x143 & ~x310 & ~x313 & ~x341 & ~x393 & ~x446 & ~x504;
assign c1128 =  x68 &  x96 &  x322 &  x379 & ~x31 & ~x51 & ~x90 & ~x197 & ~x198 & ~x229 & ~x482 & ~x779;
assign c1130 =  x577 & ~x6 & ~x98 & ~x184 & ~x191 & ~x192 & ~x241 & ~x304 & ~x506 & ~x510;
assign c1132 =  x551 & ~x82 & ~x119 & ~x173 & ~x188 & ~x203 & ~x282 & ~x427 & ~x460 & ~x505 & ~x559 & ~x732;
assign c1134 =  x322 &  x351 & ~x1 & ~x74 & ~x78 & ~x84 & ~x106 & ~x120 & ~x143 & ~x148 & ~x225 & ~x258 & ~x311 & ~x357 & ~x388 & ~x415 & ~x416 & ~x455 & ~x478 & ~x481 & ~x507 & ~x510 & ~x537 & ~x539 & ~x555 & ~x557 & ~x621 & ~x666 & ~x699 & ~x701 & ~x724 & ~x728 & ~x735 & ~x736 & ~x780;
assign c1136 =  x678 &  x705 & ~x73 & ~x265;
assign c1138 =  x9 &  x401 & ~x198;
assign c1140 =  x217 &  x647;
assign c1142 =  x372;
assign c1144 =  x330 &  x667 & ~x742;
assign c1146 =  x647 & ~x39 & ~x152;
assign c1148 = ~x47 & ~x73 & ~x102 & ~x121 & ~x164 & ~x167 & ~x171 & ~x199 & ~x202 & ~x229 & ~x231 & ~x232 & ~x260 & ~x271 & ~x279 & ~x285 & ~x287 & ~x330 & ~x339 & ~x357 & ~x373 & ~x415 & ~x423 & ~x428 & ~x429 & ~x447 & ~x455 & ~x478 & ~x536 & ~x555 & ~x567 & ~x722 & ~x738 & ~x752 & ~x758;
assign c1150 =  x700;
assign c1152 =  x41 &  x296 & ~x8 & ~x202 & ~x230 & ~x371 & ~x373 & ~x424 & ~x547 & ~x748;
assign c1154 =  x579 &  x710 & ~x220 & ~x312 & ~x657 & ~x693;
assign c1156 =  x202 &  x371 &  x548;
assign c1158 =  x39 &  x295 &  x542;
assign c1160 = ~x47 & ~x59 & ~x81 & ~x88 & ~x112 & ~x160 & ~x174 & ~x200 & ~x246 & ~x259 & ~x273 & ~x307 & ~x314 & ~x329 & ~x338 & ~x386 & ~x399 & ~x402 & ~x406 & ~x429 & ~x449 & ~x499 & ~x505 & ~x555 & ~x582 & ~x609 & ~x637 & ~x644 & ~x667 & ~x668 & ~x695 & ~x696 & ~x698 & ~x699 & ~x720 & ~x723 & ~x725 & ~x759 & ~x783;
assign c1162 =  x379 &  x435 & ~x203 & ~x240 & ~x258 & ~x298 & ~x355 & ~x367 & ~x672 & ~x696 & ~x719 & ~x724;
assign c1164 = ~x93 & ~x94 & ~x149 & ~x150 & ~x177 & ~x178 & ~x232 & ~x259 & ~x288 & ~x294 & ~x303 & ~x314 & ~x396 & ~x442 & ~x481 & ~x526 & ~x564 & ~x693 & ~x705;
assign c1166 =  x69 &  x296 &  x409 &  x466 & ~x133 & ~x134 & ~x555 & ~x695 & ~x696 & ~x728;
assign c1168 =  x324 & ~x73 & ~x87 & ~x371 & ~x377 & ~x606;
assign c1170 =  x492 & ~x149 & ~x333 & ~x386 & ~x410 & ~x514;
assign c1172 =  x485 &  x540 &  x595 &  x677 & ~x155 & ~x475 & ~x618;
assign c1174 =  x322 &  x492 & ~x297 & ~x383 & ~x466;
assign c1176 =  x435 & ~x43 & ~x77 & ~x195 & ~x196 & ~x212 & ~x223 & ~x229 & ~x255 & ~x270 & ~x286 & ~x298 & ~x315 & ~x384 & ~x390 & ~x396 & ~x421 & ~x423 & ~x505 & ~x538 & ~x691;
assign c1178 =  x540 &  x704 & ~x182 & ~x236;
assign c1180 =  x647 & ~x95 & ~x97 & ~x335 & ~x624;
assign c1182 =  x695 & ~x552;
assign c1184 =  x739 & ~x91 & ~x170 & ~x202 & ~x314 & ~x454 & ~x598 & ~x673 & ~x717;
assign c1186 =  x39 &  x68 &  x97 & ~x74 & ~x94 & ~x120 & ~x133 & ~x360 & ~x503 & ~x504 & ~x612 & ~x733 & ~x777;
assign c1188 =  x370 &  x484 & ~x153;
assign c1190 =  x703;
assign c1192 =  x672;
assign c1194 =  x374 &  x380 &  x550 & ~x666;
assign c1196 =  x241 &  x299 &  x327 &  x356 & ~x81 & ~x199;
assign c1198 =  x741 &  x742 &  x770 & ~x106 & ~x117 & ~x146 & ~x198 & ~x612 & ~x690 & ~x694 & ~x722 & ~x745;
assign c1200 =  x677 & ~x44 & ~x169 & ~x223 & ~x367 & ~x452 & ~x518 & ~x645 & ~x670 & ~x685 & ~x725 & ~x729 & ~x756;
assign c1202 =  x634 & ~x325 & ~x552 & ~x715;
assign c1204 =  x311;
assign c1206 =  x380 &  x551 &  x710 & ~x505;
assign c1208 =  x656 & ~x120 & ~x196 & ~x260 & ~x288 & ~x402 & ~x612 & ~x645 & ~x690 & ~x693;
assign c1210 =  x651 & ~x73 & ~x196 & ~x197 & ~x200 & ~x290 & ~x309 & ~x444 & ~x587 & ~x702 & ~x725;
assign c1212 =  x354 & ~x33 & ~x95 & ~x259 & ~x427 & ~x638 & ~x692 & ~x697;
assign c1214 = ~x19 & ~x106 & ~x115 & ~x196 & ~x231 & ~x286 & ~x311 & ~x341 & ~x371 & ~x374 & ~x377 & ~x394 & ~x453 & ~x546 & ~x635 & ~x693;
assign c1216 =  x211 & ~x32 & ~x89 & ~x103 & ~x137 & ~x173 & ~x388 & ~x424 & ~x431 & ~x450 & ~x454 & ~x633 & ~x661 & ~x693 & ~x730 & ~x750 & ~x766 & ~x779;
assign c1218 =  x124 &  x294 &  x322 & ~x120;
assign c1220 =  x244 &  x619;
assign c1222 =  x174 &  x483;
assign c1224 =  x324 &  x552 &  x771 & ~x60 & ~x669;
assign c1226 =  x90;
assign c1228 =  x551 &  x744 & ~x368 & ~x662 & ~x692;
assign c1230 =  x68 &  x378 &  x379 &  x403 & ~x537;
assign c1232 =  x757;
assign c1234 =  x70 &  x155 &  x298 &  x496 & ~x258;
assign c1236 =  x757;
assign c1238 =  x218;
assign c1240 =  x68 &  x266 &  x351 &  x408 & ~x388 & ~x498 & ~x620;
assign c1242 =  x520 &  x605 & ~x298 & ~x594;
assign c1244 =  x300 &  x380 & ~x322;
assign c1246 =  x297 &  x439 & ~x2 & ~x52 & ~x106 & ~x193 & ~x219 & ~x229 & ~x248 & ~x250 & ~x340 & ~x369 & ~x429 & ~x501 & ~x507 & ~x531 & ~x556;
assign c1248 =  x90 &  x483 & ~x179;
assign c1250 =  x327 &  x441 & ~x201 & ~x258 & ~x332 & ~x477 & ~x781;
assign c1252 =  x219;
assign c1254 = ~x59 & ~x144 & ~x183 & ~x184 & ~x192 & ~x196 & ~x285 & ~x304 & ~x325 & ~x330 & ~x342 & ~x365 & ~x384 & ~x418 & ~x426 & ~x438 & ~x446 & ~x472 & ~x498 & ~x589 & ~x637 & ~x639 & ~x669 & ~x727 & ~x750 & ~x761;
assign c1256 =  x246 &  x647 & ~x241 & ~x269;
assign c1258 =  x704 & ~x127 & ~x155 & ~x209 & ~x236;
assign c1260 =  x295 &  x324 & ~x84 & ~x142 & ~x229 & ~x341 & ~x342 & ~x395 & ~x402 & ~x414 & ~x577 & ~x668;
assign c1262 =  x607 &  x609 &  x612 & ~x690;
assign c1264 =  x296 &  x324 & ~x1 & ~x21 & ~x53 & ~x59 & ~x88 & ~x331 & ~x360 & ~x368 & ~x429 & ~x430 & ~x453 & ~x454 & ~x456 & ~x560 & ~x575 & ~x591 & ~x610 & ~x693 & ~x700 & ~x727 & ~x749 & ~x763;
assign c1266 =  x273 &  x353 &  x483;
assign c1268 =  x124 &  x379 & ~x3 & ~x59 & ~x73 & ~x134 & ~x159 & ~x242 & ~x285 & ~x286 & ~x298 & ~x301 & ~x311 & ~x331 & ~x359 & ~x382 & ~x561 & ~x566 & ~x757 & ~x758;
assign c1270 =  x175 & ~x40 & ~x45 & ~x69 & ~x97 & ~x254 & ~x296 & ~x468 & ~x629 & ~x736;
assign c1272 =  x273 & ~x406;
assign c1274 =  x353 &  x551 &  x710;
assign c1276 =  x274 & ~x352 & ~x444 & ~x742;
assign c1278 = ~x98 & ~x118 & ~x126 & ~x221 & ~x283 & ~x298 & ~x307 & ~x318 & ~x320 & ~x423 & ~x454 & ~x479 & ~x600 & ~x674;
assign c1280 =  x520 & ~x150 & ~x325 & ~x326 & ~x438 & ~x442 & ~x467;
assign c1282 =  x152 &  x153 &  x324 & ~x16 & ~x691;
assign c1284 =  x556;
assign c1286 =  x298 &  x441 & ~x78 & ~x133 & ~x258 & ~x340 & ~x614 & ~x726;
assign c1288 =  x229 &  x427;
assign c1290 =  x540 &  x705 & ~x153 & ~x601;
assign c1292 = ~x127 & ~x130 & ~x148 & ~x157 & ~x162 & ~x184 & ~x221 & ~x225 & ~x258 & ~x268 & ~x276 & ~x298 & ~x302 & ~x314 & ~x324 & ~x325 & ~x398 & ~x410 & ~x420 & ~x451 & ~x468 & ~x478 & ~x623;
assign c1294 =  x758;
assign c1296 =  x324 &  x325 &  x741 &  x743 &  x744 & ~x663 & ~x694;
assign c1298 =  x378 &  x520 & ~x312 & ~x325 & ~x454 & ~x481 & ~x615 & ~x721;
assign c1300 =  x552 &  x555 & ~x152 & ~x476;
assign c1302 =  x268 &  x382 & ~x399 & ~x406 & ~x435 & ~x696;
assign c1304 =  x6;
assign c1306 =  x585;
assign c1308 =  x757;
assign c1310 =  x70 &  x325 & ~x18 & ~x107 & ~x117 & ~x314 & ~x334 & ~x393 & ~x430 & ~x454 & ~x642;
assign c1312 =  x297 & ~x312 & ~x406 & ~x429 & ~x661;
assign c1314 =  x579 & ~x80 & ~x443 & ~x492 & ~x514 & ~x667;
assign c1316 =  x655 & ~x217 & ~x233 & ~x288 & ~x314 & ~x574 & ~x602;
assign c1318 =  x68 &  x266 &  x323 &  x408 & ~x442;
assign c1320 =  x520 & ~x159 & ~x201 & ~x213 & ~x219 & ~x240 & ~x242 & ~x275 & ~x298 & ~x355 & ~x450 & ~x454 & ~x455 & ~x649;
assign c1322 =  x380 &  x550 & ~x269 & ~x298;
assign c1324 =  x241 &  x469 & ~x283 & ~x361 & ~x395 & ~x639;
assign c1326 =  x520 & ~x43 & ~x60 & ~x88 & ~x134 & ~x172 & ~x195 & ~x197 & ~x251 & ~x269 & ~x270 & ~x337 & ~x442 & ~x531 & ~x534 & ~x553 & ~x696 & ~x779;
assign c1328 = ~x78 & ~x98 & ~x127 & ~x130 & ~x163 & ~x168 & ~x193 & ~x254 & ~x261 & ~x270 & ~x361 & ~x478 & ~x487 & ~x516 & ~x653;
assign c1330 =  x662 &  x693;
assign c1332 = ~x0 & ~x63 & ~x78 & ~x79 & ~x136 & ~x202 & ~x204 & ~x205 & ~x342 & ~x344 & ~x398 & ~x403 & ~x418 & ~x482 & ~x548 & ~x642 & ~x674 & ~x777 & ~x778 & ~x780;
assign c1334 =  x97 &  x267 & ~x73 & ~x251 & ~x314 & ~x398;
assign c1336 =  x241 &  x354 & ~x229;
assign c1338 =  x173 &  x455;
assign c1340 =  x124 & ~x33 & ~x100 & ~x103 & ~x116 & ~x164 & ~x241 & ~x268 & ~x275 & ~x298 & ~x312 & ~x335 & ~x355 & ~x364 & ~x385 & ~x397 & ~x455 & ~x471 & ~x724;
assign c1342 =  x324 & ~x28 & ~x73 & ~x91 & ~x116 & ~x146 & ~x172 & ~x173 & ~x174 & ~x188 & ~x258 & ~x281 & ~x313 & ~x314 & ~x372 & ~x452 & ~x633 & ~x689 & ~x690 & ~x705;
assign c1344 =  x427 &  x720;
assign c1346 =  x677 & ~x211 & ~x422 & ~x481;
assign c1348 = ~x6 & ~x27 & ~x43 & ~x197 & ~x270 & ~x286 & ~x328 & ~x357 & ~x384 & ~x454 & ~x482 & ~x544 & ~x586 & ~x645 & ~x666 & ~x693 & ~x716 & ~x754;
assign c1350 =  x295 &  x380 &  x409 &  x437 & ~x20 & ~x24 & ~x77 & ~x340 & ~x511 & ~x520 & ~x723 & ~x750;
assign c1352 =  x552 &  x555;
assign c1354 =  x39 &  x68 &  x96 &  x296 & ~x200 & ~x639 & ~x695;
assign c1356 =  x664 &  x667;
assign c1358 = ~x21 & ~x28 & ~x51 & ~x52 & ~x73 & ~x80 & ~x85 & ~x93 & ~x103 & ~x109 & ~x141 & ~x145 & ~x156 & ~x162 & ~x167 & ~x176 & ~x192 & ~x203 & ~x228 & ~x232 & ~x249 & ~x255 & ~x260 & ~x272 & ~x275 & ~x282 & ~x288 & ~x301 & ~x304 & ~x316 & ~x342 & ~x361 & ~x365 & ~x389 & ~x413 & ~x414 & ~x415 & ~x417 & ~x421 & ~x423 & ~x447 & ~x449 & ~x452 & ~x455 & ~x470 & ~x528 & ~x560 & ~x581 & ~x617 & ~x699 & ~x719 & ~x720 & ~x722 & ~x730 & ~x746 & ~x749 & ~x756 & ~x763 & ~x776;
assign c1360 =  x726;
assign c1362 =  x239 &  x268 &  x409 & ~x73 & ~x451 & ~x464;
assign c1364 =  x684 & ~x249 & ~x259 & ~x438 & ~x439 & ~x580 & ~x767;
assign c1366 =  x662 & ~x714;
assign c1368 =  x41 & ~x134 & ~x146 & ~x167 & ~x197 & ~x203 & ~x341 & ~x362 & ~x377 & ~x393 & ~x402 & ~x700;
assign c1370 =  x70 &  x269 &  x440 & ~x314 & ~x725 & ~x753;
assign c1372 =  x406 & ~x91 & ~x119 & ~x184 & ~x204 & ~x260 & ~x315 & ~x326 & ~x353 & ~x384 & ~x538 & ~x621;
assign c1374 =  x190;
assign c1376 =  x98 &  x184 &  x269 &  x297 &  x326 & ~x781;
assign c1378 =  x353 & ~x146 & ~x190 & ~x230 & ~x249 & ~x260 & ~x284 & ~x331 & ~x373 & ~x427 & ~x430 & ~x666 & ~x668 & ~x719;
assign c1380 =  x578 &  x579 &  x580 & ~x387 & ~x532 & ~x665 & ~x692;
assign c1382 =  x655 &  x685 &  x742 &  x743 & ~x193 & ~x303 & ~x591 & ~x615 & ~x695 & ~x738;
assign c1384 =  x701;
assign c1386 =  x520 & ~x119 & ~x127 & ~x138 & ~x184 & ~x298 & ~x417 & ~x510;
assign c1388 =  x156 &  x297 &  x326 & ~x20 & ~x106 & ~x170 & ~x393 & ~x425 & ~x633 & ~x666;
assign c1390 =  x727;
assign c1392 =  x428 &  x731;
assign c1394 =  x98 &  x268 &  x297 & ~x399 & ~x548 & ~x669 & ~x704 & ~x751;
assign c1396 =  x567 &  x676 & ~x98 & ~x680;
assign c1398 =  x380 &  x550 & ~x90 & ~x117 & ~x229 & ~x257 & ~x269 & ~x314 & ~x539;
assign c1400 =  x760;
assign c1402 =  x523 &  x743 &  x773 & ~x115;
assign c1404 = ~x29 & ~x77 & ~x106 & ~x173 & ~x202 & ~x204 & ~x288 & ~x317 & ~x369 & ~x373 & ~x406 & ~x481 & ~x508 & ~x690 & ~x749;
assign c1406 =  x641;
assign c1408 =  x325 & ~x385 & ~x401 & ~x605 & ~x618 & ~x636 & ~x693;
assign c1410 =  x127 &  x184 &  x297 &  x382 & ~x103 & ~x453 & ~x535;
assign c1412 =  x411 &  x667;
assign c1414 =  x272 &  x353;
assign c1416 =  x608 &  x612;
assign c1418 =  x297 &  x685 &  x743 & ~x201 & ~x750;
assign c1420 =  x8 & ~x56 & ~x83 & ~x117 & ~x199 & ~x309 & ~x368 & ~x506 & ~x536 & ~x591 & ~x670;
assign c1422 =  x297 &  x439 & ~x341 & ~x366 & ~x401 & ~x638 & ~x676;
assign c1424 = ~x98 & ~x121 & ~x145 & ~x187 & ~x240 & ~x258 & ~x260 & ~x371 & ~x586;
assign c1426 =  x413;
assign c1428 =  x465 &  x539 &  x648;
assign c1430 =  x229 &  x371;
assign c1432 =  x742 & ~x406 & ~x608 & ~x649;
assign c1434 =  x40 &  x69 &  x268 &  x297 & ~x766;
assign c1436 =  x294 &  x409 &  x570 & ~x395 & ~x450;
assign c1438 =  x579 &  x580 &  x581 & ~x81 & ~x251 & ~x388 & ~x478 & ~x666 & ~x691 & ~x724 & ~x756;
assign c1440 =  x274 &  x647;
assign c1442 = ~x24 & ~x29 & ~x82 & ~x147 & ~x165 & ~x172 & ~x203 & ~x204 & ~x221 & ~x229 & ~x285 & ~x303 & ~x334 & ~x373 & ~x377 & ~x395 & ~x402 & ~x417 & ~x502 & ~x691 & ~x706 & ~x722;
assign c1444 = ~x91 & ~x127 & ~x198 & ~x244 & ~x248 & ~x272 & ~x288 & ~x298 & ~x362 & ~x425 & ~x516 & ~x529 & ~x545 & ~x554;
assign c1446 =  x580 &  x585;
assign c1448 =  x428 & ~x290 & ~x389;
assign c1450 =  x124 &  x152 & ~x147 & ~x314 & ~x326 & ~x342 & ~x353 & ~x393 & ~x423 & ~x510;
assign c1452 =  x484 &  x511 & ~x95 & ~x96 & ~x99 & ~x126 & ~x180;
assign c1454 =  x577 &  x771 & ~x437 & ~x468;
assign c1456 =  x153 &  x294 &  x295 & ~x430 & ~x431 & ~x510 & ~x533 & ~x573 & ~x733;
assign c1458 =  x759 & ~x384;
assign c1460 =  x70 &  x156 &  x184 & ~x277;
assign c1462 =  x359;
assign c1464 =  x677 & ~x142 & ~x153 & ~x452 & ~x592 & ~x681 & ~x682;
assign c1466 =  x272 &  x325 & ~x88 & ~x110 & ~x195 & ~x198 & ~x199 & ~x220 & ~x221 & ~x225 & ~x226 & ~x331;
assign c1468 =  x68 &  x153 &  x324 &  x351 &  x380 & ~x143 & ~x366 & ~x702;
assign c1470 =  x37 &  x268 &  x717;
assign c1472 =  x294 & ~x138 & ~x148 & ~x184 & ~x222 & ~x230 & ~x298 & ~x315 & ~x326 & ~x382 & ~x447 & ~x511 & ~x512 & ~x566 & ~x723;
assign c1474 =  x297 &  x326 & ~x259 & ~x311 & ~x333 & ~x435 & ~x674 & ~x694 & ~x781;
assign c1476 =  x684 & ~x138 & ~x171 & ~x175 & ~x251 & ~x270 & ~x286 & ~x288 & ~x297 & ~x298 & ~x421 & ~x527 & ~x529 & ~x539 & ~x725;
assign c1478 =  x322 &  x465 &  x522 & ~x190 & ~x229 & ~x230 & ~x330 & ~x421 & ~x427 & ~x619 & ~x675 & ~x724 & ~x763;
assign c1480 = ~x18 & ~x31 & ~x45 & ~x49 & ~x51 & ~x56 & ~x58 & ~x73 & ~x83 & ~x131 & ~x145 & ~x172 & ~x173 & ~x219 & ~x242 & ~x244 & ~x255 & ~x260 & ~x276 & ~x286 & ~x288 & ~x298 & ~x308 & ~x316 & ~x331 & ~x357 & ~x368 & ~x390 & ~x398 & ~x454 & ~x473 & ~x509 & ~x526 & ~x557 & ~x562 & ~x568 & ~x616 & ~x622 & ~x623 & ~x691 & ~x693 & ~x755 & ~x763 & ~x765 & ~x777;
assign c1482 =  x654 &  x655 &  x743 & ~x202 & ~x315 & ~x534;
assign c1484 = ~x98 & ~x236 & ~x253 & ~x325 & ~x326 & ~x406 & ~x443 & ~x496 & ~x504 & ~x528 & ~x600 & ~x710;
assign c1486 =  x577 &  x578 &  x579 &  x580 & ~x168 & ~x194 & ~x281 & ~x366 & ~x692;
assign c1488 =  x579 &  x609 & ~x571 & ~x659;
assign c1490 =  x374 &  x376 & ~x212 & ~x220 & ~x304 & ~x694 & ~x728;
assign c1492 = ~x53 & ~x87 & ~x91 & ~x104 & ~x142 & ~x149 & ~x184 & ~x185 & ~x197 & ~x259 & ~x260 & ~x285 & ~x327 & ~x329 & ~x384 & ~x401 & ~x442 & ~x449 & ~x450 & ~x479 & ~x504 & ~x621 & ~x692 & ~x693 & ~x732 & ~x760;
assign c1494 =  x98 &  x268 &  x269 & ~x140 & ~x219 & ~x258 & ~x305 & ~x314 & ~x333 & ~x402 & ~x670 & ~x676;
assign c1496 =  x40 &  x297 & ~x94;
assign c1498 =  x324 & ~x20 & ~x220 & ~x401 & ~x406 & ~x429 & ~x583 & ~x634 & ~x693 & ~x704 & ~x753;
assign c11 =  x516 &  x544 & ~x272 & ~x299 & ~x659;
assign c13 =  x95 & ~x140 & ~x195 & ~x238 & ~x266 & ~x416 & ~x530 & ~x536 & ~x590 & ~x595;
assign c15 =  x533;
assign c17 =  x462 &  x488 &  x516 & ~x160 & ~x213 & ~x245 & ~x271;
assign c19 =  x490 &  x518 & ~x521 & ~x548 & ~x619;
assign c111 =  x487 &  x515 &  x543 & ~x85 & ~x140 & ~x141 & ~x189 & ~x242 & ~x249 & ~x256 & ~x280 & ~x447 & ~x528 & ~x563 & ~x756;
assign c113 =  x317 & ~x72 & ~x82 & ~x204 & ~x630;
assign c115 = ~x10 & ~x12 & ~x13 & ~x65 & ~x87 & ~x362 & ~x429 & ~x455 & ~x458 & ~x482 & ~x501 & ~x568 & ~x623 & ~x644 & ~x672 & ~x674 & ~x729;
assign c117 =  x194;
assign c119 =  x166;
assign c121 =  x333 & ~x669;
assign c123 =  x535 & ~x306 & ~x517;
assign c125 =  x712 &  x713 & ~x25 & ~x106 & ~x111 & ~x521 & ~x578 & ~x592 & ~x605 & ~x617;
assign c127 =  x517 &  x518 &  x545 &  x571 & ~x109;
assign c129 =  x206 &  x286 & ~x376;
assign c131 =  x395;
assign c133 = ~x113 & ~x140 & ~x319 & ~x372 & ~x423 & ~x513 & ~x589 & ~x590 & ~x653 & ~x708 & ~x711 & ~x756;
assign c135 = ~x33 & ~x56 & ~x195 & ~x223 & ~x226 & ~x263 & ~x348 & ~x461 & ~x487 & ~x542 & ~x768;
assign c137 =  x207 &  x235 &  x262 &  x290 &  x318 & ~x379 & ~x672;
assign c139 =  x43 &  x491 & ~x783;
assign c141 =  x454 & ~x169 & ~x188 & ~x215 & ~x227;
assign c143 =  x394;
assign c145 =  x519 &  x546 &  x573 &  x601;
assign c147 =  x575 &  x630 &  x657 & ~x29 & ~x54 & ~x196 & ~x476 & ~x501 & ~x588;
assign c149 =  x261 &  x288 & ~x1 & ~x10 & ~x39 & ~x72;
assign c151 =  x423 & ~x114 & ~x699 & ~x780;
assign c153 = ~x195 & ~x354 & ~x380 & ~x408 & ~x462 & ~x465 & ~x492 & ~x493 & ~x521 & ~x522 & ~x548 & ~x643;
assign c155 =  x660 &  x688 & ~x513 & ~x668;
assign c157 =  x313 &  x495 & ~x701 & ~x775;
assign c159 = ~x15 & ~x32 & ~x110 & ~x137 & ~x219 & ~x266 & ~x295 & ~x339 & ~x366 & ~x392 & ~x417 & ~x420 & ~x424 & ~x501 & ~x581 & ~x615 & ~x625 & ~x669 & ~x678 & ~x701 & ~x760;
assign c161 =  x377 & ~x22 & ~x28 & ~x130 & ~x466 & ~x467 & ~x494 & ~x521 & ~x522 & ~x549 & ~x760;
assign c163 = ~x25 & ~x51 & ~x58 & ~x89 & ~x101 & ~x113 & ~x137 & ~x140 & ~x160 & ~x187 & ~x197 & ~x214 & ~x251 & ~x310 & ~x361 & ~x493 & ~x494 & ~x505 & ~x521 & ~x548 & ~x644 & ~x699 & ~x703 & ~x730 & ~x756 & ~x761;
assign c165 =  x463 &  x491 &  x519 &  x546 & ~x224 & ~x284 & ~x338 & ~x356 & ~x475 & ~x588;
assign c167 =  x100 &  x183 & ~x87 & ~x414 & ~x469 & ~x582 & ~x584 & ~x753;
assign c169 =  x201 &  x228;
assign c171 = ~x182 & ~x238 & ~x266 & ~x321 & ~x406 & ~x443 & ~x533 & ~x538 & ~x613 & ~x680 & ~x765;
assign c173 =  x533;
assign c175 =  x95 &  x122 &  x149 &  x150 &  x177 &  x206;
assign c177 =  x507 &  x535 & ~x87 & ~x473 & ~x520 & ~x576;
assign c179 = ~x23 & ~x24 & ~x30 & ~x88 & ~x90 & ~x108 & ~x163 & ~x220 & ~x251 & ~x276 & ~x280 & ~x303 & ~x458 & ~x476 & ~x515 & ~x683 & ~x687 & ~x711 & ~x713 & ~x735 & ~x737 & ~x762;
assign c181 =  x249;
assign c183 =  x513 &  x541 &  x569 &  x653;
assign c185 =  x285 & ~x32 & ~x53 & ~x87 & ~x142 & ~x372 & ~x529 & ~x562 & ~x586 & ~x729 & ~x765;
assign c187 =  x525 & ~x306 & ~x319 & ~x711 & ~x768;
assign c189 =  x417;
assign c191 =  x490 &  x517 &  x518 &  x545 & ~x51 & ~x86 & ~x108 & ~x110 & ~x116 & ~x280 & ~x356 & ~x478 & ~x563 & ~x729 & ~x759;
assign c193 =  x508 & ~x30 & ~x463 & ~x576 & ~x602 & ~x730;
assign c195 =  x431 &  x459 &  x487 &  x515 & ~x137 & ~x167 & ~x187 & ~x388;
assign c197 =  x214 &  x494 & ~x302 & ~x658;
assign c199 =  x206 &  x262 &  x464 &  x519 & ~x3;
assign c1101 =  x462 &  x490 &  x517 & ~x132 & ~x251 & ~x273 & ~x370 & ~x498 & ~x657;
assign c1103 =  x348 &  x430 & ~x8 & ~x80 & ~x284 & ~x420 & ~x451 & ~x502 & ~x507 & ~x550 & ~x781;
assign c1105 =  x565 &  x621 & ~x30 & ~x329 & ~x711 & ~x712 & ~x741 & ~x770;
assign c1107 =  x42 &  x462 &  x490 & ~x85 & ~x110 & ~x416 & ~x699;
assign c1109 =  x95 &  x315 &  x342;
assign c1111 =  x486 &  x513 & ~x10 & ~x38 & ~x109 & ~x176 & ~x760;
assign c1113 =  x495 &  x524 & ~x170 & ~x445 & ~x477 & ~x711 & ~x727 & ~x740 & ~x741;
assign c1115 = ~x12 & ~x39 & ~x85 & ~x86 & ~x263 & ~x264 & ~x276 & ~x309 & ~x375 & ~x487 & ~x558 & ~x584 & ~x589 & ~x732 & ~x760;
assign c1117 =  x631 &  x659 &  x660 &  x713 & ~x673;
assign c1119 =  x396 &  x467 & ~x247 & ~x305;
assign c1121 =  x660 &  x687 &  x688 &  x713 & ~x112 & ~x251;
assign c1123 =  x459 &  x487 & ~x81 & ~x521 & ~x522 & ~x549 & ~x578 & ~x613 & ~x783;
assign c1125 =  x462 &  x463 &  x490 &  x518 & ~x1 & ~x3 & ~x5 & ~x54 & ~x392 & ~x418 & ~x419 & ~x423 & ~x523;
assign c1127 =  x547 &  x573 &  x574 &  x601 &  x629 & ~x0 & ~x308;
assign c1129 =  x576 &  x603 &  x631 & ~x30 & ~x54 & ~x141 & ~x168 & ~x309 & ~x310 & ~x314 & ~x475 & ~x560 & ~x596 & ~x779 & ~x782;
assign c1131 =  x226;
assign c1133 =  x226;
assign c1135 =  x513 &  x541 & ~x8 & ~x10 & ~x191 & ~x669 & ~x688 & ~x775;
assign c1137 =  x405 &  x460 & ~x113 & ~x414 & ~x554 & ~x601 & ~x700;
assign c1139 = ~x15 & ~x168 & ~x264 & ~x319 & ~x499 & ~x540 & ~x557 & ~x642 & ~x693 & ~x711 & ~x757 & ~x764;
assign c1141 =  x633 &  x660 &  x688 & ~x85 & ~x137 & ~x250 & ~x567 & ~x595 & ~x706 & ~x707 & ~x729;
assign c1143 =  x72 &  x211 & ~x568;
assign c1145 = ~x89 & ~x107 & ~x111 & ~x113 & ~x392 & ~x413 & ~x494 & ~x521 & ~x536 & ~x548 & ~x568 & ~x605 & ~x649 & ~x760;
assign c1147 =  x519 &  x546 &  x573 &  x600 & ~x32 & ~x53 & ~x55 & ~x280 & ~x420;
assign c1149 =  x207 &  x547 &  x574 &  x601;
assign c1151 =  x369 &  x494 & ~x170 & ~x218 & ~x224 & ~x770;
assign c1153 =  x72 &  x128 &  x212 & ~x331 & ~x412 & ~x530;
assign c1155 =  x507 &  x535 & ~x547;
assign c1157 =  x99 & ~x684;
assign c1159 =  x433 & ~x1 & ~x87 & ~x185 & ~x420 & ~x521 & ~x522 & ~x548;
assign c1161 = ~x238 & ~x266 & ~x377 & ~x405 & ~x474 & ~x592 & ~x644 & ~x680 & ~x697;
assign c1163 =  x444 &  x527;
assign c1165 =  x489 &  x516 &  x517 &  x544;
assign c1167 =  x481 &  x509 &  x621 & ~x1 & ~x339;
assign c1169 =  x320 &  x321 &  x348 &  x432 & ~x10 & ~x56 & ~x83 & ~x475 & ~x586;
assign c1171 =  x439 & ~x234 & ~x596 & ~x597 & ~x707 & ~x711;
assign c1173 =  x568 &  x736 & ~x628;
assign c1175 =  x278;
assign c1177 =  x339 & ~x219 & ~x779;
assign c1179 =  x154 &  x209 &  x237 &  x265 &  x321 & ~x190;
assign c1181 = ~x5 & ~x25 & ~x26 & ~x30 & ~x51 & ~x201 & ~x394 & ~x420 & ~x470 & ~x486 & ~x498 & ~x502 & ~x514 & ~x530 & ~x563 & ~x568 & ~x569 & ~x580 & ~x582 & ~x585 & ~x597 & ~x618 & ~x621 & ~x623 & ~x678 & ~x699 & ~x727 & ~x781;
assign c1183 =  x659 & ~x17 & ~x85 & ~x398 & ~x513 & ~x514 & ~x566 & ~x567 & ~x649 & ~x675 & ~x697 & ~x707;
assign c1185 =  x130 &  x158 &  x214 & ~x84;
assign c1187 =  x43 &  x323 & ~x441 & ~x568;
assign c1189 =  x390;
assign c1191 =  x332 & ~x524 & ~x609 & ~x667;
assign c1193 =  x334 & ~x775;
assign c1195 =  x631 &  x659 &  x686 & ~x596 & ~x702;
assign c1197 =  x508 & ~x115 & ~x335 & ~x476 & ~x504 & ~x656 & ~x657 & ~x661 & ~x683 & ~x728;
assign c1199 =  x534 & ~x376;
assign c1201 =  x164 &  x491;
assign c1203 =  x459 &  x486 &  x487 & ~x20 & ~x140 & ~x158 & ~x159 & ~x186 & ~x360 & ~x365 & ~x414 & ~x560 & ~x671 & ~x754;
assign c1205 =  x533;
assign c1207 =  x289 &  x317 &  x345 & ~x184 & ~x210 & ~x310 & ~x671;
assign c1209 =  x582 &  x668;
assign c1211 =  x459 &  x543 & ~x9 & ~x56 & ~x478;
assign c1213 =  x461 &  x488 &  x715 &  x716 & ~x21 & ~x58 & ~x85 & ~x163 & ~x335 & ~x416 & ~x589 & ~x760;
assign c1215 =  x129 & ~x55 & ~x318 & ~x597 & ~x684;
assign c1217 = ~x25 & ~x79 & ~x220 & ~x276 & ~x380 & ~x409 & ~x460 & ~x517 & ~x521 & ~x548 & ~x577 & ~x603 & ~x684 & ~x711;
assign c1219 = ~x108 & ~x120 & ~x409 & ~x521 & ~x572 & ~x577 & ~x602 & ~x711;
assign c1221 =  x109;
assign c1223 =  x488 &  x513 & ~x10;
assign c1225 = ~x38 & ~x111 & ~x113 & ~x148 & ~x229 & ~x342 & ~x597 & ~x599 & ~x637 & ~x711 & ~x765;
assign c1227 =  x463 &  x490 &  x518 &  x546 & ~x1 & ~x3 & ~x20 & ~x32 & ~x338 & ~x561 & ~x760;
assign c1229 = ~x1 & ~x3 & ~x36 & ~x54 & ~x84 & ~x164 & ~x220 & ~x249 & ~x408 & ~x464 & ~x476 & ~x491 & ~x493 & ~x519 & ~x521 & ~x548 & ~x560 & ~x574 & ~x578 & ~x588 & ~x712 & ~x782;
assign c1231 =  x72 &  x100 &  x128 &  x212 &  x240 & ~x3 & ~x84 & ~x358 & ~x588 & ~x727;
assign c1233 = ~x8 & ~x58 & ~x85 & ~x215 & ~x225 & ~x251 & ~x330 & ~x332 & ~x420 & ~x464 & ~x467 & ~x492 & ~x493 & ~x494 & ~x521 & ~x522 & ~x580 & ~x583 & ~x673 & ~x725 & ~x781;
assign c1235 = ~x192 & ~x263 & ~x304 & ~x659 & ~x662 & ~x684 & ~x711 & ~x745 & ~x769;
assign c1237 =  x181 &  x265 &  x321 & ~x84;
assign c1239 =  x633 &  x659 &  x660 &  x686 &  x687 & ~x4 & ~x108 & ~x483;
assign c1241 =  x339;
assign c1243 =  x396 & ~x198 & ~x364 & ~x427;
assign c1245 =  x490 &  x518 &  x545 & ~x22 & ~x61 & ~x118 & ~x141 & ~x190 & ~x218 & ~x226 & ~x272 & ~x302 & ~x388 & ~x420 & ~x443 & ~x445 & ~x479 & ~x564 & ~x672 & ~x697 & ~x731;
assign c1247 =  x347 & ~x8 & ~x224 & ~x521 & ~x530 & ~x603 & ~x619 & ~x731 & ~x783;
assign c1249 =  x562 & ~x223;
assign c1251 =  x165 &  x323 & ~x530;
assign c1253 =  x562 & ~x272 & ~x274;
assign c1255 =  x341 &  x369 &  x397 & ~x113 & ~x114 & ~x165 & ~x222 & ~x227 & ~x310 & ~x337 & ~x562 & ~x617 & ~x672 & ~x754;
assign c1257 =  x389;
assign c1259 = ~x1 & ~x13 & ~x65 & ~x471 & ~x521 & ~x568 & ~x570 & ~x577 & ~x696 & ~x730;
assign c1261 =  x541 &  x596 &  x624 &  x652 &  x708;
assign c1263 =  x404 &  x431 &  x459 &  x486 & ~x419 & ~x612;
assign c1265 =  x262 &  x290 &  x291 & ~x3 & ~x238 & ~x420 & ~x613 & ~x699 & ~x759 & ~x760;
assign c1267 =  x490 &  x517 &  x545 &  x572 & ~x58 & ~x307 & ~x531 & ~x782;
assign c1269 =  x748 & ~x578;
assign c1271 =  x474;
assign c1273 =  x306;
assign c1275 =  x433 &  x461 &  x489 &  x517;
assign c1277 =  x519 &  x547 &  x574 & ~x140 & ~x458 & ~x540;
assign c1279 =  x487 &  x543 &  x571 & ~x26 & ~x54 & ~x55 & ~x84 & ~x391 & ~x532 & ~x696 & ~x763;
assign c1281 =  x576 & ~x530 & ~x557 & ~x597 & ~x626 & ~x675;
assign c1283 =  x691 &  x692 &  x719 & ~x29 & ~x251 & ~x362 & ~x367 & ~x632 & ~x729;
assign c1285 =  x342 & ~x5 & ~x20 & ~x132 & ~x134 & ~x144 & ~x215;
assign c1287 =  x632 &  x659 &  x660 &  x687 &  x713 & ~x28 & ~x111;
assign c1289 =  x342 &  x343 & ~x6 & ~x47 & ~x59 & ~x79 & ~x86 & ~x217 & ~x366 & ~x458 & ~x689;
assign c1291 =  x73 &  x129 & ~x330 & ~x358 & ~x444 & ~x474;
assign c1293 =  x519 &  x574 & ~x51 & ~x54 & ~x84 & ~x111 & ~x195 & ~x363 & ~x513 & ~x756 & ~x759;
assign c1295 =  x388;
assign c1297 =  x93 &  x95 &  x122 &  x150 &  x177;
assign c1299 =  x433 &  x461 &  x488 & ~x340 & ~x589;
assign c1303 =  x232 & ~x348 & ~x597;
assign c1305 =  x743 & ~x28 & ~x32 & ~x238 & ~x266 & ~x521 & ~x522 & ~x534 & ~x700;
assign c1307 =  x417;
assign c1309 =  x362 & ~x40;
assign c1311 =  x262 &  x263 &  x291 &  x319 &  x347 &  x430;
assign c1313 =  x454 &  x482 &  x537 &  x593 &  x621 &  x622 & ~x5 & ~x8;
assign c1315 =  x602 &  x603 &  x629 &  x657 & ~x478;
assign c1317 =  x423;
assign c1319 =  x100 &  x128 & ~x358 & ~x756;
assign c1321 =  x418;
assign c1323 =  x446;
assign c1325 =  x509 &  x593 &  x621 & ~x33 & ~x60 & ~x136 & ~x168 & ~x280 & ~x335 & ~x393 & ~x684;
assign c1327 =  x283 & ~x5 & ~x18 & ~x32 & ~x162 & ~x508 & ~x775;
assign c1329 =  x632 &  x659 &  x686 & ~x565;
assign c1331 =  x575 &  x576 &  x603 &  x630 & ~x4 & ~x24 & ~x50 & ~x51 & ~x54 & ~x223 & ~x506 & ~x507 & ~x530 & ~x588 & ~x753;
assign c1333 =  x517 &  x600 & ~x1 & ~x164 & ~x216 & ~x253;
assign c1335 =  x576 &  x603 &  x631 &  x658 & ~x1 & ~x84 & ~x363 & ~x392 & ~x423 & ~x451 & ~x501 & ~x532 & ~x558 & ~x588 & ~x617 & ~x673 & ~x755;
assign c1337 =  x349 &  x460 & ~x606;
assign c1339 =  x459 &  x487 & ~x215 & ~x307 & ~x578;
assign c1341 =  x630 &  x657 &  x683 & ~x112 & ~x140 & ~x169 & ~x729;
assign c1343 =  x450;
assign c1345 = ~x87 & ~x136 & ~x169 & ~x408 & ~x462 & ~x464 & ~x521 & ~x522 & ~x549 & ~x578 & ~x587 & ~x708 & ~x762;
assign c1347 = ~x38 & ~x160 & ~x286 & ~x522 & ~x570 & ~x578 & ~x606 & ~x621 & ~x622 & ~x636;
assign c1349 =  x367 & ~x56 & ~x60 & ~x83 & ~x85 & ~x142 & ~x699 & ~x748 & ~x783;
assign c1351 =  x554;
assign c1353 =  x431 &  x459 &  x516 & ~x1 & ~x141 & ~x471;
assign c1355 =  x100 &  x128 & ~x187;
assign c1357 =  x72 & ~x0 & ~x524 & ~x610;
assign c1359 =  x563 &  x591 & ~x278 & ~x408;
assign c1361 =  x317 & ~x6 & ~x10 & ~x186 & ~x364 & ~x522 & ~x549 & ~x750;
assign c1363 =  x80;
assign c1365 =  x397 &  x425 &  x453 & ~x33 & ~x113 & ~x116 & ~x168 & ~x197;
assign c1367 =  x461 & ~x264;
assign c1369 = ~x63 & ~x169 & ~x250 & ~x368 & ~x392 & ~x421 & ~x446 & ~x453 & ~x457 & ~x486 & ~x500 & ~x501 & ~x514 & ~x539 & ~x540 & ~x542 & ~x560 & ~x568 & ~x597 & ~x646 & ~x654 & ~x666 & ~x676 & ~x703 & ~x710 & ~x723 & ~x726 & ~x735 & ~x737;
assign c1371 =  x43 &  x235 & ~x440 & ~x467;
assign c1373 =  x181 &  x209 & ~x46 & ~x223 & ~x380;
assign c1375 =  x415 &  x443 & ~x775;
assign c1377 =  x347 &  x430 & ~x35 & ~x109 & ~x190 & ~x578 & ~x657 & ~x730;
assign c1379 = ~x71 & ~x379 & ~x380 & ~x409 & ~x465 & ~x491 & ~x494 & ~x522 & ~x606 & ~x630;
assign c1381 =  x137 & ~x248 & ~x274 & ~x276;
assign c1383 =  x509 &  x537 & ~x117 & ~x196 & ~x366 & ~x577 & ~x604 & ~x605 & ~x766;
assign c1385 =  x508 &  x621 & ~x1 & ~x61;
assign c1387 =  x108 & ~x501 & ~x558;
assign c1389 = ~x10 & ~x64 & ~x313 & ~x392 & ~x420 & ~x508 & ~x534 & ~x535 & ~x536 & ~x584 & ~x670 & ~x686 & ~x711 & ~x714 & ~x729 & ~x740 & ~x756;
assign c1391 =  x129 & ~x8 & ~x84 & ~x339 & ~x388 & ~x597 & ~x626;
assign c1393 =  x221;
assign c1395 =  x490 &  x517 &  x545 & ~x58 & ~x77 & ~x109 & ~x160 & ~x169 & ~x256 & ~x307 & ~x310 & ~x330 & ~x336 & ~x364 & ~x416;
assign c1397 = ~x1 & ~x4 & ~x12 & ~x14 & ~x39 & ~x40 & ~x94 & ~x224 & ~x475 & ~x543 & ~x620 & ~x646 & ~x647 & ~x672 & ~x685 & ~x711 & ~x712 & ~x731 & ~x736 & ~x737 & ~x760 & ~x765;
assign c1399 =  x397 &  x425 & ~x57 & ~x87 & ~x117 & ~x169 & ~x170 & ~x249 & ~x251 & ~x277 & ~x419 & ~x445 & ~x472 & ~x473 & ~x588 & ~x674 & ~x700 & ~x727 & ~x730;
assign c1401 =  x582 &  x610 & ~x251 & ~x418 & ~x475 & ~x741 & ~x756;
assign c1403 =  x547 &  x574 &  x575 &  x601 &  x629 & ~x473 & ~x728;
assign c1405 =  x194 & ~x42 & ~x388 & ~x523 & ~x558 & ~x587 & ~x778;
assign c1407 =  x461 &  x489 & ~x1 & ~x3 & ~x105 & ~x130 & ~x214 & ~x253 & ~x577 & ~x606 & ~x640;
assign c1409 =  x310;
assign c1411 =  x573 &  x600 & ~x319 & ~x737 & ~x775;
assign c1413 = ~x45 & ~x47 & ~x356 & ~x436 & ~x437 & ~x440 & ~x521 & ~x549 & ~x577 & ~x608 & ~x611 & ~x676 & ~x728 & ~x753 & ~x759;
assign c1415 =  x244 & ~x165 & ~x408 & ~x488 & ~x659 & ~x711 & ~x713;
assign c1417 =  x602 &  x657 &  x683 & ~x451;
assign c1419 =  x462 &  x490 &  x516 &  x543 & ~x187 & ~x188;
assign c1421 = ~x31 & ~x47 & ~x84 & ~x111 & ~x112 & ~x117 & ~x141 & ~x158 & ~x228 & ~x252 & ~x387 & ~x416 & ~x420 & ~x421 & ~x424 & ~x467 & ~x475 & ~x494 & ~x501 & ~x521 & ~x522 & ~x549 & ~x580 & ~x611 & ~x646 & ~x696 & ~x728;
assign c1423 =  x488 &  x516 &  x543 & ~x27 & ~x135 & ~x280 & ~x358 & ~x420 & ~x443 & ~x531 & ~x734 & ~x778;
assign c1425 =  x631 &  x659 &  x686 &  x712;
assign c1427 =  x603 &  x630 &  x631 &  x657 & ~x507 & ~x618;
assign c1429 =  x564 & ~x144 & ~x251 & ~x684;
assign c1431 = ~x5 & ~x56 & ~x59 & ~x186 & ~x493 & ~x521 & ~x522 & ~x524 & ~x533 & ~x548 & ~x568 & ~x578 & ~x707 & ~x722 & ~x765 & ~x781;
assign c1433 =  x497 &  x582 & ~x279 & ~x769;
assign c1435 =  x181 &  x208 &  x236 &  x264 &  x292 & ~x273;
assign c1437 = ~x8 & ~x10 & ~x23 & ~x28 & ~x52 & ~x114 & ~x432 & ~x486 & ~x513 & ~x534 & ~x568 & ~x656 & ~x711 & ~x737 & ~x762 & ~x765;
assign c1439 =  x406 & ~x12 & ~x18 & ~x42 & ~x52 & ~x67 & ~x110 & ~x111 & ~x252 & ~x264 & ~x451 & ~x612 & ~x641;
assign c1441 =  x719 & ~x36 & ~x166 & ~x218 & ~x273 & ~x361 & ~x427 & ~x501 & ~x502 & ~x640 & ~x781;
assign c1443 =  x519 &  x546 &  x572 &  x573;
assign c1445 =  x631 &  x659 &  x686 &  x712 & ~x420 & ~x536;
assign c1447 = ~x4 & ~x12 & ~x33 & ~x40 & ~x55 & ~x80 & ~x424 & ~x504 & ~x529 & ~x568 & ~x586 & ~x592 & ~x619 & ~x644 & ~x646 & ~x649 & ~x650 & ~x668 & ~x675 & ~x676 & ~x730 & ~x760 & ~x769 & ~x770 & ~x780;
assign c1449 =  x534;
assign c1451 =  x391;
assign c1453 = ~x80 & ~x82 & ~x251 & ~x304 & ~x351 & ~x360 & ~x380 & ~x390 & ~x406 & ~x408 & ~x437 & ~x446 & ~x474 & ~x643 & ~x683 & ~x684 & ~x711 & ~x712 & ~x740;
assign c1455 =  x660 &  x687 & ~x27 & ~x34 & ~x50 & ~x166 & ~x335 & ~x389 & ~x445 & ~x560 & ~x568 & ~x589 & ~x649 & ~x697 & ~x707 & ~x729 & ~x782;
assign c1457 = ~x13 & ~x37 & ~x237 & ~x416 & ~x619 & ~x699 & ~x711 & ~x737 & ~x741 & ~x769 & ~x780;
assign c1459 = ~x26 & ~x85 & ~x264 & ~x282 & ~x291 & ~x319 & ~x347 & ~x403 & ~x458 & ~x461 & ~x513 & ~x655 & ~x708 & ~x711 & ~x755 & ~x758;
assign c1461 =  x200 & ~x264 & ~x586;
assign c1463 =  x519 &  x546 &  x573;
assign c1465 =  x568 &  x624 &  x652 &  x708;
assign c1467 =  x575 &  x602 &  x603 &  x630 &  x657 & ~x775;
assign c1469 =  x424 &  x452 & ~x194 & ~x255 & ~x282 & ~x641 & ~x642 & ~x776;
assign c1471 =  x418;
assign c1473 = ~x1 & ~x12 & ~x13 & ~x164 & ~x311 & ~x562 & ~x568 & ~x578 & ~x589 & ~x611 & ~x645 & ~x646 & ~x737 & ~x763;
assign c1475 =  x236 &  x458 &  x513 & ~x22 & ~x588;
assign c1477 =  x603 &  x630 &  x631 &  x657 &  x658;
assign c1479 =  x150 &  x177 & ~x5 & ~x7 & ~x20 & ~x32 & ~x81 & ~x111 & ~x252 & ~x391 & ~x514 & ~x560 & ~x588 & ~x766;
assign c1481 =  x604 &  x631 &  x659 & ~x25 & ~x32 & ~x83 & ~x676 & ~x678 & ~x704 & ~x730 & ~x748;
assign c1483 =  x513 & ~x5 & ~x8 & ~x9 & ~x34 & ~x112 & ~x121 & ~x220 & ~x449 & ~x758;
assign c1485 =  x288 & ~x13 & ~x293 & ~x294 & ~x321 & ~x422 & ~x643 & ~x699 & ~x705 & ~x731 & ~x732 & ~x778;
assign c1487 =  x349 &  x433 &  x461 & ~x65 & ~x80 & ~x110 & ~x371 & ~x414 & ~x445 & ~x703 & ~x729;
assign c1489 =  x261 &  x316 &  x344 & ~x58 & ~x302 & ~x522 & ~x587;
assign c1491 =  x214 &  x242 & ~x318 & ~x514 & ~x741;
assign c1493 =  x763 &  x764;
assign c1495 =  x347 & ~x20 & ~x133 & ~x252 & ~x305 & ~x469 & ~x503;
assign c1497 =  x610 & ~x30 & ~x31 & ~x359 & ~x389 & ~x444 & ~x531 & ~x770;
assign c1499 =  x547 &  x575 &  x602 &  x629 & ~x12 & ~x25 & ~x250;
assign c20 =  x238 &  x490 &  x601 & ~x60 & ~x626;
assign c22 =  x155 &  x157 &  x184 & ~x82 & ~x112 & ~x243 & ~x270 & ~x276 & ~x289 & ~x366 & ~x778;
assign c24 =  x100 &  x128 & ~x214 & ~x271 & ~x272 & ~x298 & ~x299 & ~x308 & ~x392 & ~x395 & ~x478 & ~x496 & ~x533 & ~x553 & ~x616 & ~x618 & ~x634 & ~x637 & ~x651 & ~x664 & ~x668 & ~x676 & ~x693 & ~x721 & ~x732;
assign c26 =  x72 & ~x29 & ~x86 & ~x196 & ~x197 & ~x281 & ~x328 & ~x331 & ~x392 & ~x471 & ~x503 & ~x551 & ~x553 & ~x569 & ~x579 & ~x587 & ~x596 & ~x597 & ~x606 & ~x609 & ~x611 & ~x612 & ~x625 & ~x634 & ~x651 & ~x669 & ~x680 & ~x696 & ~x702 & ~x720 & ~x758;
assign c28 =  x369 &  x513 & ~x519;
assign c210 =  x102 &  x103 & ~x57 & ~x290 & ~x346 & ~x638;
assign c212 =  x493 & ~x269 & ~x352 & ~x353 & ~x406 & ~x473 & ~x578 & ~x579 & ~x604 & ~x608 & ~x633;
assign c214 =  x733 & ~x518;
assign c216 =  x349 & ~x3 & ~x20 & ~x21 & ~x32 & ~x50 & ~x59 & ~x63 & ~x81 & ~x86 & ~x106 & ~x110 & ~x137 & ~x157 & ~x166 & ~x187 & ~x201 & ~x218 & ~x256 & ~x276 & ~x278 & ~x279 & ~x280 & ~x303 & ~x304 & ~x308 & ~x310 & ~x335 & ~x360 & ~x361 & ~x362 & ~x391 & ~x436 & ~x502 & ~x553 & ~x563 & ~x606 & ~x620 & ~x670 & ~x693 & ~x696 & ~x701 & ~x708 & ~x735 & ~x750 & ~x760;
assign c218 =  x101 &  x102 & ~x31 & ~x216 & ~x272 & ~x335 & ~x386 & ~x503 & ~x693 & ~x731 & ~x752 & ~x763;
assign c220 =  x519 &  x546 & ~x61 & ~x299 & ~x326 & ~x577 & ~x581 & ~x605 & ~x631 & ~x632 & ~x734 & ~x750 & ~x752 & ~x755;
assign c222 =  x187 & ~x151 & ~x362 & ~x619 & ~x671;
assign c224 =  x12 & ~x445 & ~x518 & ~x546 & ~x603;
assign c226 =  x542 &  x597 & ~x30 & ~x170 & ~x248 & ~x282 & ~x501 & ~x519 & ~x520 & ~x546 & ~x547 & ~x603 & ~x629;
assign c228 =  x154 &  x155 &  x267 & ~x0 & ~x58 & ~x189 & ~x242 & ~x264 & ~x355 & ~x533 & ~x553 & ~x555 & ~x764 & ~x783;
assign c230 =  x467 &  x774 & ~x763;
assign c232 =  x326 & ~x80 & ~x158 & ~x168 & ~x212 & ~x240 & ~x251 & ~x255 & ~x443 & ~x465 & ~x475 & ~x518 & ~x546 & ~x586 & ~x613;
assign c234 =  x267 &  x574 & ~x208 & ~x442 & ~x570 & ~x578 & ~x599 & ~x649;
assign c236 =  x184 &  x185 &  x212 & ~x136 & ~x300 & ~x302 & ~x341 & ~x356 & ~x385 & ~x386 & ~x411 & ~x418 & ~x422 & ~x476 & ~x507 & ~x525 & ~x553 & ~x560 & ~x561 & ~x608 & ~x641 & ~x649 & ~x666 & ~x675 & ~x678 & ~x722 & ~x726 & ~x733 & ~x734 & ~x752;
assign c238 = ~x29 & ~x106 & ~x129 & ~x170 & ~x172 & ~x201 & ~x212 & ~x240 & ~x241 & ~x295 & ~x363 & ~x418 & ~x482 & ~x549 & ~x554 & ~x597 & ~x608 & ~x651 & ~x669 & ~x672 & ~x693;
assign c240 =  x466 &  x518 & ~x228 & ~x260 & ~x380;
assign c242 =  x181 &  x237 & ~x110 & ~x115 & ~x192 & ~x241 & ~x352 & ~x559 & ~x603 & ~x604 & ~x631;
assign c244 =  x184 &  x212 & ~x291 & ~x318 & ~x357 & ~x382 & ~x524 & ~x612 & ~x613 & ~x677 & ~x752 & ~x781;
assign c246 = ~x181 & ~x452 & ~x453 & ~x485 & ~x502 & ~x515 & ~x623 & ~x651 & ~x680 & ~x685 & ~x706 & ~x726;
assign c248 =  x381 &  x435 & ~x199 & ~x214 & ~x224 & ~x268 & ~x548 & ~x550 & ~x578 & ~x668 & ~x697;
assign c250 = ~x5 & ~x36 & ~x53 & ~x157 & ~x165 & ~x167 & ~x185 & ~x213 & ~x224 & ~x225 & ~x228 & ~x240 & ~x247 & ~x268 & ~x270 & ~x451 & ~x522 & ~x549 & ~x583 & ~x586 & ~x621 & ~x649 & ~x668 & ~x694 & ~x733 & ~x751 & ~x763 & ~x777;
assign c252 =  x384 & ~x152 & ~x261 & ~x454 & ~x490 & ~x573;
assign c254 =  x632 & ~x38 & ~x198 & ~x503 & ~x535 & ~x569 & ~x570 & ~x625 & ~x656 & ~x696;
assign c256 =  x459 & ~x21 & ~x79 & ~x135 & ~x168 & ~x189 & ~x197 & ~x201 & ~x220 & ~x222 & ~x226 & ~x227 & ~x240 & ~x308 & ~x338 & ~x439 & ~x447 & ~x502 & ~x553 & ~x577 & ~x578 & ~x606 & ~x644 & ~x651 & ~x753;
assign c258 =  x339 & ~x152 & ~x472;
assign c260 =  x466 &  x544 & ~x352;
assign c262 =  x630 & ~x117 & ~x307 & ~x356 & ~x386 & ~x450 & ~x451 & ~x495 & ~x578 & ~x579 & ~x587 & ~x592 & ~x621 & ~x647 & ~x745 & ~x750 & ~x771;
assign c264 = ~x139 & ~x291 & ~x398 & ~x442 & ~x443 & ~x566 & ~x570 & ~x596 & ~x600 & ~x629 & ~x656;
assign c266 =  x97 &  x237 &  x293 & ~x29 & ~x50 & ~x76 & ~x83 & ~x164 & ~x167 & ~x334 & ~x419 & ~x449 & ~x552 & ~x556 & ~x578 & ~x579 & ~x580 & ~x603 & ~x604 & ~x606 & ~x637 & ~x640 & ~x669 & ~x735 & ~x753;
assign c268 =  x589;
assign c270 =  x533;
assign c272 =  x440 & ~x491 & ~x602 & ~x629 & ~x739;
assign c274 =  x104 & ~x123;
assign c276 =  x459 &  x541 & ~x491 & ~x545 & ~x600 & ~x629;
assign c278 =  x188 &  x213 & ~x318 & ~x399 & ~x445 & ~x503 & ~x647;
assign c280 =  x69 &  x96 &  x432;
assign c282 =  x96 &  x381 &  x460 & ~x212 & ~x546;
assign c284 =  x104 & ~x518;
assign c286 =  x571 &  x627 &  x744 & ~x113 & ~x118 & ~x219 & ~x226 & ~x281 & ~x283 & ~x392 & ~x449 & ~x603 & ~x604 & ~x607;
assign c288 =  x310;
assign c290 =  x213 &  x214 &  x215 &  x216 & ~x329 & ~x362 & ~x389 & ~x415 & ~x779;
assign c292 =  x95 &  x297;
assign c294 =  x185 &  x492 &  x520 &  x547 & ~x8 & ~x86 & ~x446 & ~x509 & ~x530 & ~x553 & ~x558 & ~x698 & ~x732;
assign c296 = ~x203 & ~x363 & ~x412 & ~x495 & ~x550 & ~x553 & ~x569 & ~x580 & ~x596 & ~x598 & ~x626 & ~x628 & ~x690 & ~x696;
assign c298 =  x98 &  x238 & ~x133 & ~x240 & ~x251 & ~x616 & ~x680 & ~x695 & ~x759;
assign c2100 =  x485 &  x570 &  x684 & ~x579 & ~x608 & ~x621 & ~x640;
assign c2102 =  x533 &  x618;
assign c2104 = ~x1 & ~x196 & ~x302 & ~x400 & ~x468 & ~x485 & ~x486 & ~x522 & ~x578 & ~x628 & ~x710 & ~x725;
assign c2106 = ~x3 & ~x8 & ~x90 & ~x112 & ~x223 & ~x247 & ~x252 & ~x334 & ~x363 & ~x471 & ~x538 & ~x543 & ~x558 & ~x561 & ~x572 & ~x625 & ~x628 & ~x629 & ~x649 & ~x656 & ~x673 & ~x680 & ~x733 & ~x738 & ~x739 & ~x753 & ~x775 & ~x781;
assign c2108 =  x98 &  x126 &  x238 & ~x34 & ~x117 & ~x147 & ~x193 & ~x223 & ~x240 & ~x241 & ~x298 & ~x419 & ~x451 & ~x531 & ~x558 & ~x581 & ~x587 & ~x588 & ~x609 & ~x637 & ~x643 & ~x668 & ~x692 & ~x724 & ~x751;
assign c2110 =  x72 & ~x214 & ~x264 & ~x580 & ~x720;
assign c2112 =  x188 &  x216 & ~x150 & ~x151 & ~x755 & ~x761 & ~x774;
assign c2114 =  x69 &  x124 &  x571 & ~x49 & ~x106 & ~x110 & ~x112 & ~x115 & ~x222 & ~x223 & ~x278 & ~x310 & ~x362 & ~x364 & ~x502 & ~x505 & ~x525 & ~x528 & ~x530 & ~x531 & ~x581 & ~x609 & ~x638 & ~x639 & ~x695 & ~x729 & ~x755 & ~x757;
assign c2116 = ~x53 & ~x263 & ~x274 & ~x281 & ~x490 & ~x518 & ~x545 & ~x600 & ~x602 & ~x627 & ~x628 & ~x630 & ~x726 & ~x730;
assign c2118 =  x159 &  x160 & ~x291 & ~x566 & ~x780;
assign c2120 =  x381 & ~x22 & ~x57 & ~x80 & ~x88 & ~x166 & ~x169 & ~x212 & ~x213 & ~x214 & ~x220 & ~x240 & ~x268 & ~x275 & ~x295 & ~x365 & ~x474 & ~x476 & ~x556 & ~x582 & ~x701 & ~x731;
assign c2122 =  x97 &  x125 &  x181 &  x209 &  x237 & ~x18 & ~x24 & ~x29 & ~x51 & ~x56 & ~x74 & ~x82 & ~x108 & ~x114 & ~x136 & ~x143 & ~x163 & ~x168 & ~x171 & ~x199 & ~x200 & ~x214 & ~x222 & ~x223 & ~x240 & ~x241 & ~x244 & ~x251 & ~x275 & ~x276 & ~x333 & ~x392 & ~x477 & ~x531 & ~x553 & ~x558 & ~x559 & ~x560 & ~x580 & ~x614 & ~x618 & ~x669 & ~x698 & ~x701 & ~x759 & ~x761 & ~x764 & ~x780 & ~x783;
assign c2124 = ~x45 & ~x112 & ~x158 & ~x202 & ~x212 & ~x228 & ~x282 & ~x359 & ~x500 & ~x528 & ~x578 & ~x597 & ~x604 & ~x611 & ~x612 & ~x624 & ~x625 & ~x635 & ~x651 & ~x663 & ~x671 & ~x676 & ~x753 & ~x779;
assign c2126 =  x40 &  x68 & ~x30 & ~x199 & ~x238 & ~x360 & ~x387 & ~x469 & ~x530 & ~x550 & ~x674;
assign c2128 = ~x11 & ~x73 & ~x113 & ~x147 & ~x214 & ~x240 & ~x295 & ~x549;
assign c2130 =  x45 &  x576 & ~x625;
assign c2132 =  x290 & ~x83 & ~x85 & ~x186 & ~x212 & ~x239 & ~x306 & ~x496 & ~x553 & ~x578 & ~x644 & ~x699 & ~x720 & ~x781;
assign c2134 =  x367 & ~x490;
assign c2136 =  x477;
assign c2138 =  x132 &  x158 & ~x222 & ~x373;
assign c2140 = ~x262 & ~x434 & ~x461 & ~x490 & ~x518 & ~x519 & ~x544 & ~x545 & ~x546 & ~x629 & ~x656 & ~x658;
assign c2142 = ~x577 & ~x633;
assign c2144 = ~x3 & ~x263 & ~x264 & ~x360 & ~x398 & ~x450 & ~x526 & ~x533 & ~x562 & ~x600 & ~x622 & ~x628 & ~x651 & ~x683 & ~x700 & ~x702 & ~x710 & ~x723 & ~x729;
assign c2146 =  x382 &  x409 &  x435 &  x436 &  x489 & ~x25 & ~x84 & ~x214 & ~x251 & ~x308 & ~x610 & ~x613 & ~x614;
assign c2148 =  x421 &  x449 &  x589;
assign c2150 =  x40 & ~x6 & ~x73 & ~x102 & ~x129 & ~x138 & ~x159 & ~x170 & ~x173 & ~x492 & ~x530 & ~x551 & ~x579 & ~x622 & ~x755;
assign c2152 =  x570 &  x773 & ~x262 & ~x763;
assign c2154 =  x326 & ~x32 & ~x183 & ~x266 & ~x389 & ~x518 & ~x547 & ~x629;
assign c2156 =  x411 &  x542 & ~x51 & ~x54 & ~x82 & ~x111 & ~x165 & ~x169 & ~x194 & ~x195 & ~x219 & ~x224 & ~x241 & ~x277 & ~x279 & ~x296 & ~x308 & ~x471 & ~x525 & ~x612;
assign c2158 =  x618 &  x675;
assign c2160 =  x216 & ~x7 & ~x96 & ~x150 & ~x514 & ~x612 & ~x653;
assign c2162 =  x184 &  x185 &  x212 & ~x58 & ~x152 & ~x279 & ~x310 & ~x319 & ~x388 & ~x418 & ~x647;
assign c2164 =  x125 &  x490 & ~x74 & ~x103 & ~x114 & ~x132 & ~x219 & ~x240 & ~x241 & ~x254 & ~x500 & ~x550 & ~x603 & ~x609 & ~x702 & ~x733;
assign c2166 =  x130 &  x131 &  x132 & ~x273 & ~x291;
assign c2168 =  x464 &  x490 &  x517 & ~x28 & ~x33 & ~x58 & ~x143 & ~x166 & ~x171 & ~x173 & ~x193 & ~x194 & ~x197 & ~x221 & ~x222 & ~x282 & ~x285 & ~x298 & ~x301 & ~x304 & ~x306 & ~x313 & ~x338 & ~x341 & ~x393 & ~x395 & ~x446 & ~x524 & ~x527 & ~x577 & ~x583 & ~x607 & ~x619 & ~x640 & ~x648 & ~x675 & ~x681 & ~x731 & ~x735 & ~x737 & ~x762;
assign c2170 =  x184 &  x521 & ~x33 & ~x291 & ~x328 & ~x394 & ~x675;
assign c2172 =  x181 &  x467 & ~x272 & ~x638;
assign c2174 =  x104 & ~x97 & ~x359 & ~x669;
assign c2176 =  x155 &  x574 & ~x52 & ~x263 & ~x264 & ~x308 & ~x583 & ~x587 & ~x671;
assign c2178 =  x129 &  x155 &  x156 & ~x52 & ~x82 & ~x84 & ~x218 & ~x220 & ~x226 & ~x235 & ~x236 & ~x263 & ~x308 & ~x336 & ~x473 & ~x588 & ~x615 & ~x675 & ~x700 & ~x759 & ~x783;
assign c2180 =  x155 & ~x141 & ~x214 & ~x222 & ~x226 & ~x242 & ~x251 & ~x263 & ~x264 & ~x365 & ~x392 & ~x419 & ~x527 & ~x563 & ~x651 & ~x677 & ~x680 & ~x731 & ~x755 & ~x778;
assign c2182 =  x77;
assign c2184 =  x435 & ~x213 & ~x241 & ~x310 & ~x378 & ~x698 & ~x750 & ~x760;
assign c2186 =  x542 &  x597 & ~x30 & ~x54 & ~x246 & ~x281 & ~x419 & ~x500 & ~x520 & ~x546 & ~x573 & ~x631 & ~x756;
assign c2188 =  x296 &  x602 & ~x423 & ~x477 & ~x510 & ~x598 & ~x771 & ~x772 & ~x783;
assign c2190 =  x412 & ~x217 & ~x242 & ~x270 & ~x297 & ~x394 & ~x446 & ~x504 & ~x579 & ~x668 & ~x669 & ~x730 & ~x761 & ~x765;
assign c2192 =  x158 &  x184 &  x185 & ~x243 & ~x338 & ~x558;
assign c2194 =  x372 & ~x77 & ~x84 & ~x85 & ~x112 & ~x136 & ~x137 & ~x140 & ~x146 & ~x190 & ~x199 & ~x224 & ~x277 & ~x282 & ~x305 & ~x308 & ~x388 & ~x393 & ~x447 & ~x448 & ~x526 & ~x552 & ~x556 & ~x581 & ~x604 & ~x664 & ~x673 & ~x674 & ~x680 & ~x700 & ~x707;
assign c2196 =  x703 & ~x490;
assign c2198 =  x214 &  x241 & ~x0 & ~x181 & ~x434 & ~x462 & ~x490;
assign c2200 =  x155 &  x349 & ~x24 & ~x52 & ~x87 & ~x167 & ~x219 & ~x241 & ~x249 & ~x273 & ~x297 & ~x302 & ~x305 & ~x327 & ~x333 & ~x418 & ~x587 & ~x588 & ~x609 & ~x633 & ~x662 & ~x705 & ~x720 & ~x752 & ~x759;
assign c2202 =  x187 &  x189 & ~x151 & ~x399;
assign c2204 =  x125 &  x435 &  x461 & ~x22 & ~x78 & ~x109 & ~x114 & ~x135 & ~x166 & ~x200 & ~x214 & ~x241 & ~x281 & ~x304 & ~x308 & ~x338 & ~x414 & ~x418 & ~x503 & ~x524 & ~x534 & ~x549 & ~x551 & ~x609 & ~x617 & ~x622 & ~x637 & ~x638 & ~x673 & ~x679 & ~x706 & ~x728;
assign c2206 =  x95 &  x377 & ~x437 & ~x518 & ~x668;
assign c2208 =  x460 &  x515 & ~x33 & ~x50 & ~x59 & ~x108 & ~x224 & ~x248 & ~x360 & ~x471 & ~x476 & ~x490 & ~x518 & ~x560 & ~x731;
assign c2210 = ~x31 & ~x261 & ~x302 & ~x490 & ~x518 & ~x529 & ~x544 & ~x545 & ~x547 & ~x602 & ~x603 & ~x629 & ~x630 & ~x658 & ~x685 & ~x746;
assign c2212 =  x366 & ~x152;
assign c2214 =  x270 &  x271 &  x297 & ~x138 & ~x212 & ~x518;
assign c2216 =  x381 &  x632 & ~x5 & ~x412 & ~x597 & ~x611 & ~x656 & ~x669;
assign c2218 = ~x35 & ~x83 & ~x133 & ~x156 & ~x157 & ~x213 & ~x214 & ~x239 & ~x240 & ~x241 & ~x266 & ~x279 & ~x295 & ~x312 & ~x445 & ~x549 & ~x550 & ~x556 & ~x558 & ~x578 & ~x579 & ~x618 & ~x679 & ~x732;
assign c2220 =  x384 & ~x379 & ~x434 & ~x629 & ~x738;
assign c2222 =  x96 &  x406 & ~x27 & ~x45 & ~x141 & ~x198 & ~x240 & ~x309 & ~x394 & ~x493 & ~x518 & ~x520 & ~x672;
assign c2224 =  x267 &  x517 & ~x21 & ~x64 & ~x81 & ~x85 & ~x173 & ~x560 & ~x586 & ~x590 & ~x593 & ~x625 & ~x627 & ~x645 & ~x702 & ~x720 & ~x751 & ~x755;
assign c2226 =  x490 & ~x60 & ~x114 & ~x240 & ~x549 & ~x604 & ~x679 & ~x766;
assign c2228 =  x103 &  x130 & ~x245 & ~x274 & ~x545 & ~x665;
assign c2230 =  x466 & ~x0 & ~x30 & ~x51 & ~x58 & ~x60 & ~x75 & ~x78 & ~x84 & ~x111 & ~x137 & ~x171 & ~x190 & ~x200 & ~x228 & ~x247 & ~x253 & ~x269 & ~x270 & ~x272 & ~x301 & ~x326 & ~x327 & ~x366 & ~x392 & ~x553 & ~x562 & ~x586 & ~x611 & ~x641 & ~x671 & ~x672 & ~x697 & ~x732 & ~x756 & ~x763;
assign c2232 = ~x25 & ~x29 & ~x57 & ~x58 & ~x85 & ~x114 & ~x141 & ~x152 & ~x167 & ~x248 & ~x250 & ~x278 & ~x335 & ~x344 & ~x416 & ~x419 & ~x435 & ~x518 & ~x531 & ~x545 & ~x572 & ~x601 & ~x756;
assign c2234 =  x438 & ~x0 & ~x27 & ~x57 & ~x134 & ~x196 & ~x200 & ~x226 & ~x254 & ~x353 & ~x361 & ~x366 & ~x418 & ~x422 & ~x477 & ~x527 & ~x531 & ~x532 & ~x550 & ~x551 & ~x560 & ~x561 & ~x584 & ~x613 & ~x647 & ~x665 & ~x667 & ~x696 & ~x701 & ~x724 & ~x729 & ~x756 & ~x761 & ~x782;
assign c2236 =  x464 & ~x268 & ~x270 & ~x352 & ~x406 & ~x577;
assign c2238 =  x406 &  x433 & ~x56 & ~x109 & ~x167 & ~x212 & ~x214 & ~x225 & ~x227 & ~x254 & ~x256 & ~x296 & ~x309 & ~x366 & ~x393 & ~x394 & ~x444 & ~x446 & ~x465 & ~x467 & ~x471 & ~x492 & ~x503 & ~x525 & ~x531 & ~x551 & ~x585 & ~x586 & ~x620 & ~x649 & ~x674;
assign c2240 =  x67 &  x95 & ~x24 & ~x26 & ~x191 & ~x211 & ~x224 & ~x239 & ~x248 & ~x308 & ~x413 & ~x446 & ~x473 & ~x519 & ~x521 & ~x531 & ~x579 & ~x581 & ~x725 & ~x758;
assign c2242 =  x161 & ~x276 & ~x318 & ~x622 & ~x726;
assign c2244 = ~x1 & ~x33 & ~x76 & ~x90 & ~x113 & ~x118 & ~x149 & ~x170 & ~x178 & ~x208 & ~x229 & ~x417 & ~x455 & ~x485 & ~x501 & ~x529 & ~x556 & ~x568 & ~x569 & ~x581 & ~x583 & ~x592 & ~x599 & ~x623 & ~x626 & ~x627 & ~x638 & ~x650 & ~x693 & ~x704 & ~x705 & ~x710 & ~x720 & ~x750;
assign c2246 =  x533 & ~x426 & ~x491;
assign c2248 =  x186 &  x213 &  x548 & ~x356 & ~x596 & ~x680;
assign c2250 =  x456 &  x513 & ~x25 & ~x50 & ~x58 & ~x131 & ~x132 & ~x165 & ~x192 & ~x198 & ~x219 & ~x242 & ~x307 & ~x338 & ~x364 & ~x474 & ~x553 & ~x556 & ~x561 & ~x577 & ~x582 & ~x642 & ~x668 & ~x696 & ~x705;
assign c2252 =  x492 & ~x5 & ~x30 & ~x48 & ~x201 & ~x230 & ~x249 & ~x325 & ~x380 & ~x391 & ~x407 & ~x434 & ~x696;
assign c2254 = ~x51 & ~x84 & ~x159 & ~x203 & ~x214 & ~x219 & ~x242 & ~x256 & ~x295 & ~x305 & ~x336 & ~x633 & ~x646 & ~x722;
assign c2256 =  x518 & ~x192 & ~x324 & ~x575 & ~x603 & ~x604 & ~x609 & ~x630 & ~x634;
assign c2258 =  x70 &  x98 &  x125 &  x127 &  x266 & ~x185 & ~x190 & ~x213 & ~x701;
assign c2260 =  x534;
assign c2262 =  x490 & ~x25 & ~x63 & ~x111 & ~x161 & ~x255 & ~x269 & ~x270 & ~x285 & ~x303 & ~x406 & ~x552 & ~x636 & ~x638 & ~x731 & ~x762;
assign c2264 =  x381 & ~x88 & ~x194 & ~x213 & ~x218 & ~x242 & ~x243 & ~x296 & ~x364 & ~x449 & ~x493 & ~x521 & ~x550 & ~x578 & ~x581;
assign c2266 =  x215 &  x216 &  x238 & ~x151 & ~x566;
assign c2268 = ~x98 & ~x135 & ~x490 & ~x502 & ~x518 & ~x547 & ~x601 & ~x628 & ~x629 & ~x630 & ~x658 & ~x718 & ~x745 & ~x774;
assign c2270 =  x95 & ~x1 & ~x6 & ~x21 & ~x55 & ~x63 & ~x102 & ~x103 & ~x144 & ~x145 & ~x161 & ~x162 & ~x183 & ~x278 & ~x363 & ~x443 & ~x478 & ~x503 & ~x532 & ~x549 & ~x563 & ~x577 & ~x578 & ~x590 & ~x606 & ~x609 & ~x641 & ~x676 & ~x679 & ~x703 & ~x723 & ~x733 & ~x759;
assign c2272 =  x11 & ~x113 & ~x190 & ~x200 & ~x224 & ~x338 & ~x490 & ~x547 & ~x728;
assign c2274 =  x76 &  x104 & ~x247 & ~x400;
assign c2276 =  x297 & ~x5 & ~x21 & ~x35 & ~x142 & ~x170 & ~x306 & ~x358 & ~x364 & ~x436 & ~x491 & ~x492 & ~x518 & ~x729;
assign c2278 =  x96 &  x433 &  x460 & ~x546;
assign c2280 =  x212 &  x240 &  x491 &  x574 & ~x608;
assign c2282 =  x158 &  x185 & ~x263 & ~x357 & ~x448 & ~x731;
assign c2284 =  x130 &  x131 & ~x67 & ~x398 & ~x610 & ~x646 & ~x774;
assign c2286 =  x153 &  x237 &  x321 &  x544 & ~x242;
assign c2288 =  x189 & ~x123 & ~x124 & ~x510;
assign c2290 =  x216 & ~x125 & ~x347 & ~x362 & ~x455 & ~x612 & ~x648 & ~x702 & ~x759;
assign c2292 =  x96 &  x124 &  x152 &  x180 & ~x17 & ~x28 & ~x30 & ~x34 & ~x84 & ~x145 & ~x161 & ~x162 & ~x163 & ~x173 & ~x184 & ~x201 & ~x240 & ~x253 & ~x443 & ~x475 & ~x496 & ~x497 & ~x528 & ~x548 & ~x549 & ~x550 & ~x560 & ~x606 & ~x608 & ~x610 & ~x645 & ~x648 & ~x667 & ~x672 & ~x701 & ~x726 & ~x735;
assign c2294 = ~x5 & ~x78 & ~x168 & ~x251 & ~x326 & ~x367 & ~x385 & ~x443 & ~x536 & ~x541 & ~x552 & ~x569 & ~x579 & ~x592 & ~x626 & ~x639 & ~x662 & ~x690 & ~x691 & ~x704 & ~x743 & ~x770 & ~x771;
assign c2296 =  x486 &  x713 &  x714 & ~x141 & ~x240 & ~x250 & ~x607;
assign c2298 =  x412 & ~x0 & ~x17 & ~x113 & ~x519 & ~x547 & ~x558 & ~x600 & ~x601 & ~x603 & ~x628 & ~x629 & ~x631 & ~x657 & ~x658;
assign c2300 =  x185 &  x241 &  x521 & ~x440 & ~x618 & ~x729;
assign c2302 =  x213 &  x521 & ~x35 & ~x55 & ~x151;
assign c2304 =  x181 &  x571 & ~x57 & ~x90 & ~x137 & ~x221 & ~x242 & ~x249 & ~x254 & ~x268 & ~x270 & ~x276 & ~x311 & ~x586 & ~x638 & ~x670 & ~x700;
assign c2306 =  x159 &  x160 & ~x69 & ~x371;
assign c2308 =  x705 & ~x547 & ~x738 & ~x768;
assign c2310 =  x130 &  x131 & ~x29 & ~x54 & ~x58 & ~x85 & ~x167 & ~x302 & ~x348 & ~x371 & ~x420 & ~x428 & ~x478 & ~x479 & ~x500 & ~x527 & ~x531 & ~x534 & ~x535 & ~x562 & ~x566 & ~x591 & ~x621 & ~x649 & ~x696 & ~x723 & ~x729 & ~x758 & ~x783;
assign c2312 = ~x29 & ~x143 & ~x218 & ~x264 & ~x424 & ~x442 & ~x448 & ~x484 & ~x506 & ~x510 & ~x544 & ~x627 & ~x649 & ~x669 & ~x681 & ~x704 & ~x757;
assign c2314 = ~x23 & ~x61 & ~x73 & ~x85 & ~x172 & ~x176 & ~x190 & ~x240 & ~x241 & ~x244 & ~x258 & ~x300 & ~x389 & ~x499 & ~x551 & ~x578 & ~x612 & ~x623 & ~x634 & ~x643 & ~x651 & ~x662 & ~x677 & ~x678 & ~x680 & ~x691 & ~x693 & ~x705 & ~x738 & ~x755;
assign c2316 =  x214 &  x217 &  x239 & ~x596;
assign c2318 =  x466 &  x519 & ~x172 & ~x353 & ~x582 & ~x583 & ~x764;
assign c2320 =  x213 &  x217 & ~x652 & ~x680;
assign c2322 = ~x2 & ~x5 & ~x7 & ~x25 & ~x53 & ~x76 & ~x88 & ~x89 & ~x104 & ~x117 & ~x128 & ~x131 & ~x132 & ~x163 & ~x164 & ~x194 & ~x212 & ~x213 & ~x223 & ~x286 & ~x308 & ~x330 & ~x384 & ~x447 & ~x473 & ~x474 & ~x495 & ~x559 & ~x560 & ~x612 & ~x614 & ~x673 & ~x679 & ~x705 & ~x721 & ~x733 & ~x734 & ~x754 & ~x778 & ~x781;
assign c2324 =  x158 &  x466;
assign c2326 =  x187 &  x189 & ~x152 & ~x400 & ~x454;
assign c2328 =  x589;
assign c2332 =  x243 &  x440 &  x468 & ~x685;
assign c2334 =  x490 &  x516 & ~x0 & ~x6 & ~x58 & ~x117 & ~x171 & ~x199 & ~x222 & ~x226 & ~x241 & ~x254 & ~x275 & ~x284 & ~x335 & ~x363 & ~x364 & ~x498 & ~x521 & ~x549 & ~x550 & ~x555 & ~x558 & ~x575 & ~x603 & ~x604 & ~x633 & ~x694 & ~x703;
assign c2336 =  x601 & ~x5 & ~x34 & ~x36 & ~x53 & ~x106 & ~x166 & ~x223 & ~x360 & ~x512 & ~x525 & ~x554 & ~x598 & ~x615 & ~x623 & ~x625 & ~x712 & ~x731;
assign c2338 =  x677 & ~x295;
assign c2340 =  x328 &  x358 & ~x519 & ~x547;
assign c2342 =  x75 &  x76 & ~x219 & ~x427;
assign c2344 =  x602 & ~x141 & ~x189 & ~x551 & ~x570 & ~x578 & ~x579 & ~x625 & ~x626 & ~x676 & ~x683 & ~x693 & ~x720;
assign c2346 =  x188 & ~x87 & ~x123 & ~x151 & ~x152 & ~x390 & ~x537;
assign c2348 = ~x60 & ~x214 & ~x244 & ~x269 & ~x275 & ~x297 & ~x303 & ~x335 & ~x359 & ~x386 & ~x394 & ~x415 & ~x476 & ~x526 & ~x530 & ~x561 & ~x578 & ~x605 & ~x612 & ~x617 & ~x647 & ~x661 & ~x663 & ~x666 & ~x707 & ~x739 & ~x748 & ~x759 & ~x762;
assign c2350 =  x69 &  x544 & ~x1 & ~x7 & ~x27 & ~x53 & ~x90 & ~x106 & ~x131 & ~x140 & ~x187 & ~x192 & ~x196 & ~x198 & ~x216 & ~x217 & ~x251 & ~x280 & ~x281 & ~x364 & ~x393 & ~x421 & ~x474 & ~x530 & ~x551 & ~x558 & ~x578 & ~x580 & ~x611 & ~x640 & ~x643 & ~x669 & ~x702 & ~x730 & ~x754 & ~x755 & ~x757;
assign c2352 = ~x3 & ~x32 & ~x81 & ~x114 & ~x248 & ~x308 & ~x385 & ~x395 & ~x429 & ~x470 & ~x480 & ~x503 & ~x541 & ~x565 & ~x570 & ~x581 & ~x597 & ~x600 & ~x622 & ~x627 & ~x628 & ~x648 & ~x649 & ~x669 & ~x676 & ~x678 & ~x683 & ~x708 & ~x755;
assign c2354 = ~x54 & ~x63 & ~x82 & ~x83 & ~x101 & ~x212 & ~x214 & ~x240 & ~x241 & ~x243 & ~x248 & ~x273 & ~x313 & ~x418 & ~x419 & ~x445 & ~x447 & ~x470 & ~x475 & ~x497 & ~x549 & ~x556 & ~x587 & ~x623 & ~x639 & ~x675 & ~x680 & ~x703 & ~x720 & ~x782;
assign c2356 = ~x86 & ~x162 & ~x168 & ~x253 & ~x274 & ~x357 & ~x362 & ~x440 & ~x441 & ~x468 & ~x469 & ~x479 & ~x492 & ~x495 & ~x549 & ~x578 & ~x620 & ~x634 & ~x695 & ~x779;
assign c2358 =  x478;
assign c2360 =  x155 &  x183 & ~x219 & ~x240 & ~x352 & ~x420 & ~x637 & ~x755;
assign c2362 =  x412 &  x413 &  x439 & ~x577 & ~x603 & ~x605 & ~x630;
assign c2364 =  x98 &  x266 &  x290 & ~x35 & ~x331 & ~x441 & ~x554 & ~x569 & ~x625;
assign c2366 =  x765 & ~x467 & ~x469 & ~x720;
assign c2368 =  x70 &  x98 &  x406 &  x432 & ~x20 & ~x28 & ~x35 & ~x112 & ~x140 & ~x225 & ~x226 & ~x550 & ~x579 & ~x581 & ~x610 & ~x614 & ~x642 & ~x664 & ~x755;
assign c2370 =  x618;
assign c2372 =  x124 &  x406 & ~x22 & ~x77 & ~x106 & ~x135 & ~x137 & ~x144 & ~x158 & ~x169 & ~x193 & ~x198 & ~x200 & ~x226 & ~x229 & ~x240 & ~x251 & ~x278 & ~x303 & ~x307 & ~x309 & ~x334 & ~x442 & ~x467 & ~x470 & ~x502 & ~x519 & ~x520 & ~x526 & ~x555 & ~x580 & ~x583 & ~x673 & ~x676;
assign c2374 =  x459 & ~x44 & ~x87 & ~x168 & ~x282 & ~x305 & ~x306 & ~x337 & ~x463 & ~x491 & ~x518 & ~x545 & ~x573 & ~x586;
assign c2376 =  x214 &  x241 &  x269 & ~x113 & ~x137 & ~x181 & ~x385 & ~x450 & ~x477 & ~x501 & ~x510 & ~x561 & ~x752;
assign c2378 =  x438 &  x464 & ~x88 & ~x172 & ~x173 & ~x216 & ~x226 & ~x243 & ~x255 & ~x258 & ~x352 & ~x557 & ~x578 & ~x603 & ~x608 & ~x609 & ~x639 & ~x752 & ~x759;
assign c2380 =  x299 &  x367;
assign c2382 =  x67 &  x377 &  x402 & ~x393 & ~x550 & ~x579 & ~x702;
assign c2384 =  x158 &  x185 & ~x290 & ~x291 & ~x337 & ~x356 & ~x359 & ~x692 & ~x752;
assign c2386 =  x212 &  x576 & ~x496 & ~x530 & ~x534 & ~x626 & ~x677 & ~x731;
assign c2388 =  x508 &  x625;
assign c2390 =  x161 & ~x123 & ~x755;
assign c2392 =  x184 &  x212 & ~x26 & ~x33 & ~x48 & ~x57 & ~x151 & ~x153 & ~x362 & ~x391 & ~x412 & ~x420 & ~x503 & ~x505 & ~x532 & ~x533 & ~x584 & ~x612 & ~x681 & ~x682 & ~x700 & ~x704 & ~x707 & ~x752 & ~x780;
assign c2394 =  x124 &  x152 & ~x56 & ~x75 & ~x78 & ~x84 & ~x89 & ~x104 & ~x157 & ~x164 & ~x182 & ~x195 & ~x212 & ~x238 & ~x240 & ~x245 & ~x249 & ~x275 & ~x279 & ~x281 & ~x283 & ~x335 & ~x361 & ~x365 & ~x445 & ~x474 & ~x478 & ~x522 & ~x523 & ~x531 & ~x534 & ~x550 & ~x556 & ~x560 & ~x588 & ~x640 & ~x646 & ~x667 & ~x694 & ~x724 & ~x752;
assign c2396 =  x39 & ~x3 & ~x89 & ~x142 & ~x164 & ~x238 & ~x282 & ~x416 & ~x447 & ~x491 & ~x518 & ~x555 & ~x587 & ~x641 & ~x668 & ~x677;
assign c2398 =  x75 & ~x393 & ~x590 & ~x594 & ~x622 & ~x706;
assign c2400 =  x519 &  x545 & ~x1 & ~x9 & ~x58 & ~x113 & ~x142 & ~x168 & ~x327 & ~x357 & ~x381 & ~x475 & ~x577 & ~x579 & ~x591 & ~x632 & ~x638 & ~x646 & ~x670 & ~x680 & ~x698 & ~x700 & ~x734;
assign c2402 =  x180 & ~x62 & ~x143 & ~x193 & ~x238 & ~x240 & ~x254 & ~x255 & ~x305 & ~x338 & ~x391 & ~x392 & ~x531 & ~x582 & ~x602 & ~x777;
assign c2404 =  x155 &  x184 &  x212 & ~x57 & ~x61 & ~x87 & ~x139 & ~x298 & ~x299 & ~x336 & ~x444 & ~x534 & ~x606 & ~x634 & ~x635 & ~x668 & ~x692 & ~x733 & ~x734 & ~x750 & ~x752 & ~x781;
assign c2406 =  x437 &  x490 & ~x3 & ~x87 & ~x136 & ~x165 & ~x191 & ~x200 & ~x298 & ~x338 & ~x351 & ~x444 & ~x469 & ~x523 & ~x552 & ~x588 & ~x617 & ~x645 & ~x646 & ~x647 & ~x668 & ~x678 & ~x698 & ~x701 & ~x730 & ~x754;
assign c2408 =  x439 &  x773 & ~x325;
assign c2410 =  x396 &  x541;
assign c2412 =  x75 &  x76 &  x104;
assign c2414 =  x381 &  x382 & ~x59 & ~x79 & ~x83 & ~x142 & ~x167 & ~x307 & ~x331 & ~x419 & ~x447 & ~x529 & ~x545 & ~x546 & ~x561 & ~x587 & ~x629 & ~x630 & ~x671 & ~x731;
assign c2416 =  x95 &  x263 & ~x30 & ~x82 & ~x84 & ~x135 & ~x156 & ~x170 & ~x171 & ~x184 & ~x200 & ~x226 & ~x228 & ~x279 & ~x305 & ~x308 & ~x309 & ~x336 & ~x337 & ~x395 & ~x447 & ~x448 & ~x557 & ~x588 & ~x607 & ~x608 & ~x616 & ~x619 & ~x638 & ~x648 & ~x756;
assign c2418 =  x69 &  x70 &  x97 &  x237 & ~x2 & ~x29 & ~x85 & ~x121 & ~x422 & ~x623;
assign c2420 =  x602 & ~x481 & ~x570 & ~x578 & ~x627 & ~x633 & ~x679 & ~x680 & ~x771 & ~x776;
assign c2422 = ~x43 & ~x98 & ~x235 & ~x407 & ~x472 & ~x490 & ~x519 & ~x547 & ~x600 & ~x629 & ~x739;
assign c2424 =  x459 &  x515 & ~x1 & ~x137 & ~x219 & ~x228 & ~x285 & ~x451 & ~x525 & ~x552 & ~x597 & ~x649 & ~x680;
assign c2426 =  x213 &  x214 &  x241 &  x242 & ~x376 & ~x536 & ~x648 & ~x673;
assign c2428 =  x483 &  x511 & ~x22 & ~x46 & ~x55 & ~x85 & ~x112 & ~x171 & ~x198 & ~x222 & ~x223 & ~x226 & ~x228 & ~x248 & ~x270 & ~x283 & ~x297 & ~x334 & ~x364 & ~x421 & ~x450 & ~x581 & ~x614 & ~x639 & ~x665 & ~x694 & ~x723 & ~x729 & ~x734 & ~x735;
assign c2430 =  x158 &  x159 &  x184 &  x185 & ~x302 & ~x306 & ~x364 & ~x695 & ~x730;
assign c2432 =  x241 &  x242 &  x243 & ~x80 & ~x83 & ~x181 & ~x640 & ~x643 & ~x648;
assign c2434 =  x369 &  x625;
assign c2436 =  x397 &  x542 & ~x32 & ~x56 & ~x59 & ~x112 & ~x191 & ~x277 & ~x309 & ~x474 & ~x504 & ~x528 & ~x549 & ~x574 & ~x576 & ~x701 & ~x757;
assign c2438 =  x181 &  x411 & ~x268 & ~x504 & ~x604;
assign c2440 =  x682 & ~x24 & ~x87 & ~x111 & ~x115 & ~x143 & ~x191 & ~x222 & ~x240 & ~x256 & ~x268 & ~x339 & ~x360 & ~x421 & ~x447 & ~x528 & ~x602 & ~x629;
assign c2442 =  x405 & ~x25 & ~x59 & ~x81 & ~x86 & ~x88 & ~x104 & ~x109 & ~x112 & ~x156 & ~x161 & ~x186 & ~x188 & ~x198 & ~x213 & ~x249 & ~x252 & ~x306 & ~x310 & ~x336 & ~x358 & ~x364 & ~x437 & ~x440 & ~x444 & ~x472 & ~x475 & ~x492 & ~x503 & ~x521 & ~x524 & ~x549 & ~x550 & ~x579 & ~x583 & ~x584 & ~x639 & ~x649 & ~x693 & ~x702 & ~x734 & ~x755 & ~x759 & ~x781 & ~x782;
assign c2444 =  x183 &  x184 &  x212 & ~x20 & ~x50 & ~x75 & ~x79 & ~x87 & ~x151 & ~x152 & ~x252 & ~x327 & ~x364 & ~x411 & ~x524 & ~x615 & ~x644 & ~x724 & ~x755;
assign c2446 =  x421;
assign c2448 =  x186 &  x438 &  x466 &  x521 & ~x456;
assign c2450 =  x69 &  x97 &  x181 &  x209 &  x237 & ~x57 & ~x84 & ~x162 & ~x213 & ~x281 & ~x283 & ~x391 & ~x532 & ~x578 & ~x580 & ~x644 & ~x645 & ~x647 & ~x705 & ~x734 & ~x752 & ~x761;
assign c2452 =  x603 & ~x221 & ~x391 & ~x394 & ~x439 & ~x457 & ~x495 & ~x580 & ~x600 & ~x643 & ~x649 & ~x680 & ~x761;
assign c2454 =  x483 & ~x105 & ~x162 & ~x163 & ~x173 & ~x186 & ~x214 & ~x216 & ~x227 & ~x256 & ~x393 & ~x417 & ~x420 & ~x421 & ~x445 & ~x446 & ~x474 & ~x476 & ~x527 & ~x552 & ~x557 & ~x558 & ~x579 & ~x581 & ~x589 & ~x590 & ~x612 & ~x613 & ~x614 & ~x636 & ~x666 & ~x667 & ~x703 & ~x763 & ~x783;
assign c2456 =  x67 &  x95 & ~x49 & ~x163 & ~x183 & ~x218 & ~x442 & ~x518 & ~x548 & ~x550 & ~x616;
assign c2458 =  x372 &  x377 & ~x81 & ~x108 & ~x113 & ~x133 & ~x142 & ~x190 & ~x198 & ~x200 & ~x282 & ~x420 & ~x527 & ~x551 & ~x577 & ~x579 & ~x580 & ~x583 & ~x606 & ~x610 & ~x668 & ~x698 & ~x732 & ~x735 & ~x781;
assign c2460 =  x377 & ~x6 & ~x186 & ~x248 & ~x466 & ~x598 & ~x770;
assign c2462 =  x98 &  x354 &  x381 & ~x252 & ~x268 & ~x554 & ~x669 & ~x707;
assign c2464 = ~x26 & ~x29 & ~x58 & ~x118 & ~x181 & ~x198 & ~x225 & ~x306 & ~x360 & ~x390 & ~x456 & ~x483 & ~x498 & ~x500 & ~x566 & ~x589 & ~x594 & ~x598 & ~x625 & ~x626 & ~x651 & ~x656 & ~x752;
assign c2466 =  x184 &  x464 &  x491 & ~x87 & ~x291 & ~x300 & ~x319 & ~x553 & ~x587;
assign c2468 =  x366;
assign c2470 =  x648 & ~x462 & ~x491 & ~x546 & ~x628;
assign c2472 =  x74 & ~x263 & ~x598;
assign c2474 =  x155 &  x492 & ~x1 & ~x32 & ~x113 & ~x144 & ~x221 & ~x248 & ~x270 & ~x272 & ~x282 & ~x300 & ~x326 & ~x391 & ~x417 & ~x500 & ~x504 & ~x507 & ~x533 & ~x550 & ~x578 & ~x581 & ~x588 & ~x667 & ~x673 & ~x676 & ~x678 & ~x694 & ~x702 & ~x704 & ~x751 & ~x780;
assign c2476 =  x412 &  x746 & ~x679 & ~x727;
assign c2478 =  x674;
assign c2480 =  x372 &  x570 & ~x107 & ~x143 & ~x166 & ~x198 & ~x256 & ~x547 & ~x583 & ~x586;
assign c2482 = ~x263 & ~x264 & ~x275 & ~x280 & ~x359 & ~x369 & ~x414 & ~x442 & ~x450 & ~x500 & ~x501 & ~x505 & ~x539 & ~x544 & ~x612 & ~x616 & ~x622 & ~x629 & ~x646 & ~x656 & ~x657 & ~x675 & ~x702 & ~x704 & ~x759;
assign c2484 = ~x151 & ~x351 & ~x490 & ~x518 & ~x544 & ~x600 & ~x628 & ~x685 & ~x743 & ~x756;
assign c2486 =  x427 &  x455 &  x570 & ~x309 & ~x585;
assign c2488 = ~x98 & ~x151 & ~x350 & ~x488 & ~x489 & ~x490 & ~x491 & ~x544 & ~x628 & ~x710;
assign c2490 =  x733 & ~x518;
assign c2492 = ~x304 & ~x319 & ~x389 & ~x414 & ~x452 & ~x485 & ~x488 & ~x511 & ~x515 & ~x544 & ~x588 & ~x600 & ~x621 & ~x629 & ~x656 & ~x755;
assign c2494 =  x394 & ~x206 & ~x434;
assign c2496 =  x95 &  x433 &  x460 & ~x111 & ~x117 & ~x145 & ~x197 & ~x337 & ~x389 & ~x519 & ~x529 & ~x549 & ~x611 & ~x675;
assign c2498 =  x714 & ~x2 & ~x50 & ~x57 & ~x74 & ~x89 & ~x91 & ~x113 & ~x116 & ~x159 & ~x170 & ~x200 & ~x214 & ~x218 & ~x242 & ~x296 & ~x330 & ~x395 & ~x422 & ~x500 & ~x534 & ~x535 & ~x560 & ~x577 & ~x587 & ~x589 & ~x604 & ~x605 & ~x608 & ~x615 & ~x631 & ~x639 & ~x645 & ~x667 & ~x672 & ~x673 & ~x694 & ~x733 & ~x735 & ~x755 & ~x765 & ~x783;
assign c21 =  x316 & ~x293 & ~x460 & ~x464;
assign c23 =  x389;
assign c25 =  x447;
assign c27 = ~x64 & ~x78 & ~x199 & ~x203 & ~x232 & ~x249 & ~x287 & ~x340 & ~x343 & ~x395 & ~x402 & ~x428 & ~x430 & ~x457 & ~x459 & ~x483 & ~x504 & ~x530 & ~x618 & ~x671 & ~x674 & ~x733 & ~x761 & ~x767;
assign c29 =  x473;
assign c211 = ~x20 & ~x21 & ~x44 & ~x71 & ~x75 & ~x85 & ~x100 & ~x127 & ~x641 & ~x705 & ~x713 & ~x742 & ~x770;
assign c213 =  x703;
assign c215 =  x362;
assign c217 =  x348 & ~x7 & ~x10 & ~x33 & ~x61 & ~x64 & ~x82 & ~x86 & ~x136 & ~x177 & ~x204 & ~x258 & ~x260 & ~x278 & ~x283 & ~x314 & ~x359 & ~x366 & ~x369 & ~x392 & ~x421 & ~x621 & ~x648 & ~x704 & ~x733 & ~x751;
assign c219 =  x323 &  x409 &  x771 & ~x25 & ~x82 & ~x87 & ~x89 & ~x163 & ~x229 & ~x246 & ~x248 & ~x306 & ~x341 & ~x366 & ~x389 & ~x392 & ~x454 & ~x497 & ~x531 & ~x699;
assign c221 =  x205 & ~x270 & ~x350 & ~x769;
assign c223 =  x118 &  x147 & ~x476;
assign c225 =  x112;
assign c227 =  x323 & ~x6 & ~x24 & ~x28 & ~x51 & ~x58 & ~x59 & ~x105 & ~x111 & ~x112 & ~x139 & ~x140 & ~x163 & ~x167 & ~x188 & ~x193 & ~x201 & ~x202 & ~x203 & ~x247 & ~x249 & ~x255 & ~x273 & ~x277 & ~x285 & ~x286 & ~x288 & ~x303 & ~x311 & ~x312 & ~x333 & ~x387 & ~x413 & ~x416 & ~x427 & ~x429 & ~x452 & ~x457 & ~x470 & ~x477 & ~x484 & ~x498 & ~x502 & ~x504 & ~x507 & ~x539 & ~x558 & ~x614 & ~x694 & ~x696 & ~x720 & ~x729 & ~x754 & ~x762 & ~x764;
assign c229 =  x221;
assign c231 =  x333;
assign c233 =  x177 &  x232 & ~x43 & ~x431;
assign c235 =  x306;
assign c237 =  x426 &  x507;
assign c239 = ~x8 & ~x19 & ~x30 & ~x51 & ~x53 & ~x60 & ~x63 & ~x133 & ~x203 & ~x204 & ~x216 & ~x227 & ~x250 & ~x257 & ~x277 & ~x282 & ~x285 & ~x316 & ~x329 & ~x335 & ~x337 & ~x341 & ~x396 & ~x402 & ~x403 & ~x417 & ~x430 & ~x440 & ~x454 & ~x478 & ~x496 & ~x512 & ~x528 & ~x559 & ~x565 & ~x589 & ~x607 & ~x634 & ~x648 & ~x704 & ~x721 & ~x729 & ~x731 & ~x737 & ~x759 & ~x764 & ~x776 & ~x777;
assign c243 =  x66 &  x177;
assign c245 =  x348 &  x376 & ~x107 & ~x160 & ~x177 & ~x226 & ~x232 & ~x310 & ~x338 & ~x370 & ~x424 & ~x439 & ~x452;
assign c247 =  x472;
assign c249 =  x117 &  x378;
assign c251 =  x700;
assign c253 =  x718 & ~x202 & ~x280 & ~x287 & ~x398 & ~x419 & ~x444 & ~x450 & ~x510 & ~x534 & ~x549;
assign c255 =  x387 & ~x99;
assign c257 =  x445;
assign c259 =  x112;
assign c261 =  x194;
assign c263 =  x389;
assign c265 =  x655 &  x656 &  x657 & ~x400 & ~x767;
assign c267 = ~x43 & ~x53 & ~x64 & ~x119 & ~x350 & ~x682 & ~x687 & ~x715 & ~x721 & ~x722 & ~x732 & ~x744 & ~x756 & ~x769;
assign c269 =  x363;
assign c271 =  x472;
assign c273 = ~x8 & ~x20 & ~x75 & ~x81 & ~x119 & ~x141 & ~x148 & ~x205 & ~x255 & ~x260 & ~x277 & ~x288 & ~x339 & ~x345 & ~x347 & ~x387 & ~x449 & ~x455 & ~x496 & ~x506 & ~x672 & ~x704 & ~x732 & ~x774;
assign c275 =  x465 & ~x103 & ~x219 & ~x230 & ~x286 & ~x312 & ~x445 & ~x456 & ~x538 & ~x723;
assign c277 =  x739 & ~x176 & ~x204 & ~x455 & ~x592;
assign c279 =  x454 & ~x459;
assign c281 =  x391;
assign c283 =  x739 &  x769 & ~x177;
assign c285 =  x251;
assign c287 =  x277;
assign c289 =  x207 & ~x106 & ~x191 & ~x200 & ~x227 & ~x229 & ~x255 & ~x283 & ~x404 & ~x456 & ~x458 & ~x459 & ~x536 & ~x564 & ~x666 & ~x733;
assign c291 =  x207 & ~x3 & ~x84 & ~x88 & ~x106 & ~x145 & ~x249 & ~x284 & ~x311 & ~x312 & ~x366 & ~x395 & ~x430 & ~x431 & ~x453 & ~x456 & ~x459 & ~x672 & ~x704;
assign c293 =  x594;
assign c295 =  x343 & ~x294;
assign c297 =  x302 & ~x292 & ~x689;
assign c299 =  x690 & ~x82 & ~x287 & ~x311 & ~x343 & ~x384 & ~x728;
assign c2101 =  x173 &  x202 & ~x292;
assign c2103 =  x501;
assign c2105 =  x700;
assign c2107 =  x334;
assign c2109 =  x509 & ~x154 & ~x403;
assign c2111 =  x147 & ~x13 & ~x40 & ~x154 & ~x280 & ~x336 & ~x392 & ~x727;
assign c2113 =  x426 & ~x433 & ~x742 & ~x744;
assign c2115 =  x140;
assign c2117 =  x454 &  x592;
assign c2119 =  x525 & ~x146;
assign c2121 =  x203 &  x247;
assign c2123 =  x742 &  x743 &  x770 & ~x117 & ~x167 & ~x343 & ~x345 & ~x368 & ~x428 & ~x767 & ~x775;
assign c2125 =  x681 & ~x455 & ~x470 & ~x764 & ~x778;
assign c2127 =  x711 &  x740 & ~x85 & ~x170 & ~x285 & ~x371 & ~x452 & ~x453 & ~x476;
assign c2129 =  x391;
assign c2131 =  x203 & ~x17 & ~x100;
assign c2133 =  x681 &  x711 & ~x429;
assign c2135 =  x653 & ~x191 & ~x226 & ~x227 & ~x366 & ~x397 & ~x427 & ~x444 & ~x480 & ~x592 & ~x728 & ~x762 & ~x763;
assign c2137 =  x174 & ~x293;
assign c2141 =  x397 &  x481 & ~x599 & ~x654 & ~x680;
assign c2143 =  x582 & ~x308 & ~x365 & ~x532 & ~x643 & ~x762;
assign c2145 =  x717 &  x738 &  x740;
assign c2147 =  x581 & ~x8 & ~x367 & ~x392 & ~x733;
assign c2149 = ~x2 & ~x77 & ~x88 & ~x94 & ~x195 & ~x276 & ~x333 & ~x343 & ~x384 & ~x430 & ~x431 & ~x442 & ~x455 & ~x459 & ~x466 & ~x482 & ~x485 & ~x541 & ~x565 & ~x694 & ~x774;
assign c2151 =  x291 &  x320 & ~x83 & ~x287 & ~x317;
assign c2153 =  x191 &  x203;
assign c2155 =  x319 &  x718 & ~x343 & ~x356;
assign c2157 =  x390;
assign c2159 = ~x22 & ~x27 & ~x48 & ~x55 & ~x56 & ~x57 & ~x58 & ~x75 & ~x83 & ~x86 & ~x160 & ~x174 & ~x177 & ~x229 & ~x245 & ~x250 & ~x256 & ~x274 & ~x276 & ~x286 & ~x345 & ~x346 & ~x364 & ~x392 & ~x415 & ~x416 & ~x420 & ~x423 & ~x428 & ~x457 & ~x480 & ~x560 & ~x565 & ~x580 & ~x584 & ~x589 & ~x612 & ~x623 & ~x669 & ~x689 & ~x698 & ~x702 & ~x724 & ~x733 & ~x737 & ~x754;
assign c2161 =  x672;
assign c2163 =  x359;
assign c2165 =  x655 & ~x92 & ~x120 & ~x177 & ~x341 & ~x372 & ~x427 & ~x594 & ~x779;
assign c2167 =  x739 &  x743 & ~x682;
assign c2169 =  x771 & ~x102 & ~x229 & ~x257 & ~x287 & ~x288 & ~x314 & ~x316 & ~x399 & ~x441 & ~x444 & ~x450 & ~x501 & ~x506 & ~x535;
assign c2171 =  x740 &  x742 & ~x130 & ~x230 & ~x252 & ~x401 & ~x428 & ~x509 & ~x777;
assign c2173 =  x386 & ~x77 & ~x135 & ~x509 & ~x564 & ~x565 & ~x620 & ~x645 & ~x692;
assign c2175 =  x482 &  x535;
assign c2177 =  x359 & ~x41;
assign c2179 =  x424 &  x426;
assign c2181 =  x178 &  x205 &  x233 & ~x198 & ~x432 & ~x447 & ~x664 & ~x723;
assign c2183 =  x418;
assign c2185 =  x178 &  x206 &  x207 & ~x430;
assign c2187 =  x343 & ~x71 & ~x381 & ~x433;
assign c2189 =  x231 & ~x13 & ~x42 & ~x44 & ~x71 & ~x99 & ~x269;
assign c2191 =  x207 &  x295 &  x715 & ~x77 & ~x339 & ~x459 & ~x567;
assign c2195 =  x361;
assign c2197 =  x507 & ~x349 & ~x376;
assign c2199 =  x331;
assign c2203 =  x267 &  x742 &  x769 & ~x77 & ~x166 & ~x204 & ~x232 & ~x286 & ~x367 & ~x426 & ~x470 & ~x610 & ~x752;
assign c2205 =  x202 & ~x207 & ~x292 & ~x625 & ~x654;
assign c2207 =  x457;
assign c2209 =  x330 & ~x265 & ~x292 & ~x293 & ~x436 & ~x719 & ~x745;
assign c2211 =  x391;
assign c2213 =  x737 &  x739 & ~x509;
assign c2215 =  x110;
assign c2217 =  x389;
assign c2219 =  x582 & ~x385 & ~x413;
assign c2221 =  x136;
assign c2223 =  x178 &  x233 &  x234 &  x261;
assign c2225 = ~x11 & ~x40 & ~x420 & ~x458 & ~x689 & ~x700 & ~x744 & ~x756 & ~x769 & ~x779;
assign c2227 =  x507 & ~x41 & ~x515;
assign c2229 =  x550 & ~x708;
assign c2231 =  x293 & ~x202 & ~x287 & ~x372 & ~x411 & ~x458 & ~x459 & ~x471 & ~x497 & ~x501 & ~x560 & ~x689;
assign c2233 =  x566 & ~x209 & ~x477 & ~x543 & ~x630;
assign c2235 =  x352 &  x743 & ~x3 & ~x221 & ~x230 & ~x259 & ~x332 & ~x426 & ~x457 & ~x702;
assign c2237 =  x246 &  x429 &  x430;
assign c2239 =  x169;
assign c2241 = ~x55 & ~x79 & ~x89 & ~x121 & ~x122 & ~x201 & ~x202 & ~x230 & ~x247 & ~x257 & ~x260 & ~x278 & ~x290 & ~x313 & ~x451 & ~x458 & ~x528 & ~x563 & ~x621 & ~x636 & ~x671 & ~x688 & ~x696 & ~x703 & ~x707 & ~x736 & ~x753 & ~x757;
assign c2243 =  x203 & ~x209 & ~x322 & ~x459;
assign c2245 =  x334;
assign c2247 =  x425 & ~x69 & ~x431 & ~x486 & ~x654;
assign c2249 =  x500;
assign c2251 =  x626 & ~x312 & ~x397 & ~x426 & ~x455 & ~x458 & ~x484 & ~x621 & ~x670;
assign c2253 =  x292 & ~x77 & ~x95 & ~x140 & ~x176 & ~x202 & ~x227 & ~x231 & ~x246 & ~x259 & ~x339 & ~x438 & ~x475 & ~x501 & ~x553 & ~x567 & ~x650;
assign c2255 =  x294 & ~x21 & ~x29 & ~x76 & ~x78 & ~x91 & ~x110 & ~x113 & ~x163 & ~x223 & ~x232 & ~x258 & ~x310 & ~x342 & ~x358 & ~x373 & ~x391 & ~x392 & ~x399 & ~x402 & ~x403 & ~x416 & ~x424 & ~x431 & ~x476 & ~x480 & ~x482 & ~x483 & ~x620 & ~x672 & ~x694 & ~x699 & ~x775;
assign c2257 =  x608 & ~x188;
assign c2259 =  x637 & ~x77 & ~x340;
assign c2261 =  x757;
assign c2263 =  x151 &  x516 & ~x202 & ~x429 & ~x502;
assign c2265 =  x207 &  x716 & ~x202 & ~x260 & ~x284 & ~x368 & ~x423 & ~x445 & ~x469 & ~x496;
assign c2267 =  x114;
assign c2269 =  x573 & ~x28 & ~x140 & ~x311 & ~x339 & ~x394 & ~x422 & ~x426 & ~x433 & ~x458 & ~x459;
assign c2271 =  x262 &  x350 &  x435 & ~x44;
assign c2273 =  x127 & ~x18 & ~x107 & ~x174 & ~x435 & ~x445 & ~x464 & ~x520 & ~x673 & ~x764 & ~x767;
assign c2275 =  x700;
assign c2277 =  x201 & ~x10 & ~x236 & ~x265;
assign c2279 =  x728;
assign c2281 =  x291 &  x346 &  x633;
assign c2283 =  x347 &  x430 &  x457 & ~x91 & ~x450;
assign c2285 =  x414;
assign c2287 =  x315 & ~x420 & ~x541 & ~x654 & ~x775;
assign c2289 =  x236 & ~x39 & ~x66 & ~x219 & ~x225 & ~x289 & ~x316 & ~x359 & ~x371 & ~x395 & ~x396 & ~x479 & ~x481 & ~x639 & ~x679 & ~x767;
assign c2291 =  x361;
assign c2293 =  x71 & ~x23 & ~x299 & ~x312 & ~x400 & ~x432 & ~x459 & ~x512 & ~x717;
assign c2295 = ~x46 & ~x104 & ~x127 & ~x212 & ~x587 & ~x767 & ~x769 & ~x774 & ~x776;
assign c2297 =  x736;
assign c2299 =  x719 & ~x11 & ~x202 & ~x471;
assign c2301 =  x739 &  x740 & ~x94 & ~x120 & ~x147 & ~x148 & ~x189 & ~x192 & ~x230 & ~x416 & ~x509 & ~x556 & ~x672;
assign c2303 =  x582 & ~x119 & ~x501;
assign c2305 =  x334;
assign c2307 =  x718 &  x719 & ~x256;
assign c2309 =  x391;
assign c2311 =  x375 &  x718 & ~x372 & ~x411;
assign c2313 =  x296 & ~x60 & ~x62 & ~x75 & ~x83 & ~x89 & ~x148 & ~x149 & ~x160 & ~x166 & ~x168 & ~x177 & ~x203 & ~x226 & ~x246 & ~x282 & ~x311 & ~x312 & ~x316 & ~x343 & ~x375 & ~x414 & ~x530 & ~x587 & ~x611 & ~x635 & ~x639 & ~x669 & ~x674 & ~x726 & ~x753;
assign c2315 =  x136 &  x193;
assign c2317 =  x178 &  x262 & ~x48 & ~x114 & ~x167 & ~x423 & ~x425 & ~x534 & ~x562 & ~x673 & ~x700 & ~x761;
assign c2319 =  x656 & ~x432 & ~x540 & ~x668;
assign c2321 =  x122 &  x123 &  x178 &  x205;
assign c2323 =  x716 &  x742 & ~x48 & ~x289 & ~x341 & ~x343 & ~x401 & ~x422 & ~x505 & ~x558 & ~x565;
assign c2325 =  x740 & ~x176 & ~x311 & ~x401 & ~x428 & ~x429 & ~x475 & ~x529;
assign c2327 =  x207 &  x319 & ~x67 & ~x342;
assign c2329 =  x435 &  x626 & ~x485 & ~x594;
assign c2331 =  x391;
assign c2333 =  x663 & ~x2 & ~x28 & ~x106 & ~x218 & ~x252 & ~x307 & ~x312 & ~x387 & ~x422 & ~x482 & ~x559;
assign c2335 = ~x6 & ~x73 & ~x286 & ~x301 & ~x330 & ~x360 & ~x370 & ~x432 & ~x433 & ~x458 & ~x459 & ~x505 & ~x513 & ~x719;
assign c2337 =  x250;
assign c2339 =  x289 &  x344;
assign c2341 =  x410 &  x554;
assign c2343 =  x573 & ~x29 & ~x133 & ~x203 & ~x230 & ~x232 & ~x274 & ~x287 & ~x370 & ~x372 & ~x393 & ~x401 & ~x420 & ~x426 & ~x431 & ~x459 & ~x482 & ~x509 & ~x568 & ~x640 & ~x644 & ~x663 & ~x678 & ~x689 & ~x706 & ~x755 & ~x762 & ~x773 & ~x776;
assign c2345 =  x86;
assign c2347 =  x553 &  x594 & ~x612;
assign c2349 =  x234 &  x262 &  x345 &  x346;
assign c2351 =  x203 &  x259 & ~x42 & ~x765 & ~x769;
assign c2353 =  x418;
assign c2355 =  x5 &  x729;
assign c2357 =  x592;
assign c2359 =  x446;
assign c2361 =  x653 & ~x166 & ~x219 & ~x286 & ~x372;
assign c2363 =  x207 &  x234 &  x262 & ~x52 & ~x195 & ~x219 & ~x251 & ~x252 & ~x588 & ~x592 & ~x643 & ~x751;
assign c2365 =  x540 & ~x230 & ~x312 & ~x393 & ~x585;
assign c2367 =  x295 & ~x119 & ~x204 & ~x232 & ~x261 & ~x283 & ~x310 & ~x347 & ~x374 & ~x427 & ~x561 & ~x565 & ~x650;
assign c2369 =  x178 &  x206 &  x234 &  x261 & ~x54 & ~x83 & ~x479 & ~x564;
assign c2371 =  x718 &  x719 & ~x312 & ~x355 & ~x466;
assign c2373 =  x220 & ~x297 & ~x464;
assign c2375 =  x430 & ~x350 & ~x413 & ~x426 & ~x463;
assign c2377 =  x430 &  x512;
assign c2379 =  x681 & ~x91 & ~x310 & ~x483 & ~x707 & ~x779;
assign c2381 =  x149 &  x262;
assign c2383 =  x398 & ~x348;
assign c2385 = ~x27 & ~x52 & ~x81 & ~x112 & ~x119 & ~x120 & ~x134 & ~x145 & ~x225 & ~x288 & ~x339 & ~x404 & ~x425 & ~x430 & ~x432 & ~x450 & ~x458 & ~x459 & ~x513 & ~x539 & ~x556 & ~x564 & ~x651 & ~x678 & ~x699 & ~x724 & ~x733;
assign c2387 =  x537 & ~x42 & ~x208 & ~x459 & ~x460;
assign c2389 =  x581 & ~x194 & ~x394 & ~x753;
assign c2391 =  x697;
assign c2393 =  x390;
assign c2395 =  x151 &  x234 & ~x455;
assign c2397 =  x174 & ~x293;
assign c2399 =  x718 & ~x77 & ~x107 & ~x133 & ~x140 & ~x256 & ~x372 & ~x399 & ~x415 & ~x453 & ~x564 & ~x753;
assign c2401 =  x222;
assign c2403 =  x621 & ~x265 & ~x422;
assign c2405 =  x205 &  x356 & ~x48 & ~x480 & ~x666 & ~x694;
assign c2407 =  x595 & ~x145 & ~x146 & ~x282 & ~x370 & ~x590 & ~x762;
assign c2409 =  x390;
assign c2411 =  x419;
assign c2413 =  x628 &  x631 & ~x313 & ~x458 & ~x459;
assign c2415 =  x389;
assign c2417 =  x121 &  x122 &  x233 & ~x110 & ~x450 & ~x643 & ~x696 & ~x759;
assign c2419 =  x769 & ~x48 & ~x230 & ~x331 & ~x430 & ~x458 & ~x744;
assign c2421 =  x236 & ~x109 & ~x119 & ~x121 & ~x148 & ~x189 & ~x199 & ~x234 & ~x422 & ~x590 & ~x767;
assign c2423 = ~x24 & ~x47 & ~x48 & ~x108 & ~x167 & ~x218 & ~x278 & ~x287 & ~x360 & ~x405 & ~x427 & ~x430 & ~x458 & ~x459 & ~x500 & ~x538 & ~x588 & ~x670 & ~x696 & ~x737 & ~x752;
assign c2425 =  x149;
assign c2427 =  x378 &  x771 & ~x43 & ~x458;
assign c2429 =  x359;
assign c2431 =  x276;
assign c2433 =  x302 &  x329;
assign c2435 =  x375 &  x718 & ~x175;
assign c2437 =  x173 & ~x293;
assign c2439 =  x333;
assign c2441 =  x71 &  x348 & ~x204 & ~x329;
assign c2443 =  x512 &  x566 & ~x279 & ~x360 & ~x480 & ~x532;
assign c2445 = ~x293 & ~x769;
assign c2447 =  x430 &  x457 &  x484 & ~x227 & ~x369 & ~x452;
assign c2449 =  x201 &  x230 & ~x40;
assign c2451 =  x403 &  x458 &  x718 & ~x399;
assign c2453 =  x672;
assign c2455 =  x500;
assign c2457 =  x681 & ~x104 & ~x283 & ~x456 & ~x511 & ~x766 & ~x777;
assign c2459 =  x291 &  x319 &  x347 &  x348 & ~x122 & ~x767;
assign c2463 =  x424 &  x425 &  x426;
assign c2465 =  x454 &  x591 & ~x569;
assign c2467 =  x315 &  x594 & ~x653;
assign c2469 =  x193;
assign c2471 =  x526 &  x594 & ~x476;
assign c2473 =  x389;
assign c2475 =  x737 &  x746;
assign c2477 =  x176 &  x428 & ~x488;
assign c2479 =  x636 & ~x220 & ~x223 & ~x254 & ~x285 & ~x304 & ~x364 & ~x778;
assign c2481 =  x430 &  x718 & ~x356;
assign c2483 =  x502;
assign c2485 =  x503;
assign c2487 =  x418;
assign c2489 =  x528;
assign c2491 =  x414 & ~x105 & ~x566;
assign c2493 =  x191;
assign c2495 =  x512 &  x539 &  x594 & ~x424 & ~x476 & ~x479;
assign c2497 =  x320 & ~x26 & ~x48 & ~x177 & ~x194 & ~x204 & ~x261 & ~x276 & ~x300 & ~x303 & ~x368 & ~x413 & ~x533 & ~x585 & ~x589 & ~x615 & ~x667 & ~x678;
assign c2499 =  x739 &  x742 & ~x219 & ~x425 & ~x500 & ~x513;
assign c30 =  x610 & ~x18 & ~x35 & ~x84 & ~x170 & ~x199 & ~x412 & ~x466 & ~x589 & ~x602 & ~x631 & ~x640 & ~x641 & ~x669 & ~x672;
assign c32 =  x250 &  x418;
assign c34 =  x46 &  x245;
assign c36 =  x556 & ~x245 & ~x470 & ~x523;
assign c38 =  x399 & ~x23 & ~x28 & ~x32 & ~x134 & ~x136 & ~x191 & ~x192 & ~x200 & ~x247 & ~x255 & ~x257 & ~x283 & ~x331 & ~x340 & ~x359 & ~x418 & ~x452 & ~x517 & ~x584 & ~x589 & ~x590 & ~x591 & ~x619 & ~x620 & ~x643 & ~x671 & ~x673 & ~x695 & ~x702 & ~x763 & ~x778 & ~x781 & ~x783;
assign c310 =  x721 & ~x327 & ~x577;
assign c312 =  x499 & ~x54 & ~x328 & ~x411 & ~x440 & ~x467 & ~x494 & ~x495 & ~x496 & ~x517 & ~x522 & ~x588 & ~x705 & ~x726;
assign c314 =  x218 &  x498 &  x499 & ~x561 & ~x585;
assign c316 =  x334 & ~x465 & ~x570;
assign c318 = ~x146 & ~x227 & ~x465 & ~x467 & ~x472 & ~x515 & ~x518 & ~x570;
assign c320 =  x526 &  x554 & ~x384 & ~x477 & ~x551 & ~x568;
assign c322 = ~x11 & ~x60 & ~x256 & ~x261 & ~x278 & ~x309 & ~x376 & ~x555 & ~x574;
assign c324 =  x363 & ~x304 & ~x486;
assign c326 =  x608 & ~x6 & ~x51 & ~x134 & ~x146 & ~x460 & ~x466 & ~x492 & ~x677 & ~x705;
assign c328 =  x775 & ~x150 & ~x194 & ~x519;
assign c330 =  x445 & ~x454 & ~x465 & ~x495;
assign c332 =  x635 & ~x190 & ~x334 & ~x470 & ~x627 & ~x675;
assign c334 =  x722 & ~x573 & ~x580 & ~x603 & ~x688;
assign c336 =  x190 &  x218 &  x526;
assign c338 =  x136 &  x305;
assign c340 =  x356 &  x636 & ~x110 & ~x113 & ~x135 & ~x194 & ~x220 & ~x223 & ~x278 & ~x305 & ~x616 & ~x629;
assign c342 =  x356 &  x408 & ~x50 & ~x54 & ~x80 & ~x136 & ~x279 & ~x545 & ~x600 & ~x603 & ~x713;
assign c344 = ~x8 & ~x24 & ~x25 & ~x26 & ~x51 & ~x55 & ~x61 & ~x82 & ~x83 & ~x92 & ~x106 & ~x109 & ~x113 & ~x171 & ~x190 & ~x191 & ~x222 & ~x224 & ~x249 & ~x278 & ~x336 & ~x466 & ~x571 & ~x574 & ~x577 & ~x604 & ~x624 & ~x626 & ~x656 & ~x712 & ~x763 & ~x783;
assign c346 =  x386 &  x537 &  x638 & ~x521;
assign c348 =  x243 & ~x384 & ~x502 & ~x628 & ~x711;
assign c350 =  x650 & ~x30 & ~x154 & ~x166 & ~x233 & ~x260 & ~x337 & ~x421 & ~x476 & ~x571 & ~x587 & ~x728;
assign c352 =  x306 &  x334 &  x418 & ~x543;
assign c354 =  x326 &  x328 &  x378;
assign c356 =  x221 & ~x294 & ~x430;
assign c358 =  x356 &  x384 & ~x166 & ~x470 & ~x544 & ~x702;
assign c360 =  x763;
assign c362 =  x498 &  x526 &  x666 & ~x384 & ~x705;
assign c364 =  x296 &  x327 &  x609;
assign c366 =  x73 &  x101 &  x129 & ~x114 & ~x234 & ~x375 & ~x475;
assign c368 =  x375 &  x424 & ~x545;
assign c370 =  x747 & ~x60 & ~x65 & ~x322 & ~x419 & ~x445 & ~x476 & ~x544 & ~x546 & ~x627 & ~x659;
assign c372 =  x466 &  x494 & ~x289 & ~x348 & ~x405;
assign c374 =  x262 & ~x58 & ~x224 & ~x225 & ~x412 & ~x438 & ~x457 & ~x650 & ~x709;
assign c376 =  x501;
assign c378 =  x45 &  x71 &  x72;
assign c380 =  x129 &  x678;
assign c382 =  x310 & ~x95 & ~x244;
assign c384 =  x749 & ~x278 & ~x551 & ~x654 & ~x687;
assign c386 =  x385 &  x693 & ~x109;
assign c388 =  x232 & ~x90 & ~x164 & ~x261 & ~x359 & ~x640;
assign c390 =  x192 & ~x45 & ~x61 & ~x328 & ~x586 & ~x645 & ~x719;
assign c392 =  x355 &  x408 & ~x38 & ~x51 & ~x166 & ~x192 & ~x278 & ~x306 & ~x543 & ~x657 & ~x671;
assign c394 =  x363 & ~x440;
assign c396 =  x73 & ~x104 & ~x168 & ~x472 & ~x504;
assign c398 =  x129 &  x212 & ~x164 & ~x208 & ~x249 & ~x278 & ~x334 & ~x391 & ~x555;
assign c3100 =  x160 &  x216 &  x356 &  x384 & ~x350 & ~x529;
assign c3102 =  x503 & ~x466;
assign c3104 =  x638 & ~x440 & ~x523 & ~x576 & ~x607 & ~x631;
assign c3106 =  x423 & ~x328 & ~x467 & ~x469 & ~x494 & ~x521 & ~x545 & ~x575;
assign c3108 =  x394 &  x422 &  x450 & ~x470 & ~x489 & ~x626;
assign c3110 =  x241 &  x394 &  x422 &  x450;
assign c3112 =  x387 &  x414 &  x496 &  x524 & ~x0 & ~x26 & ~x348 & ~x505 & ~x588 & ~x617 & ~x647 & ~x697 & ~x700 & ~x702;
assign c3114 =  x239 & ~x352 & ~x467 & ~x561 & ~x593 & ~x618 & ~x677;
assign c3116 =  x241 &  x267 & ~x384 & ~x440 & ~x600 & ~x627 & ~x693;
assign c3118 =  x611 & ~x467 & ~x496 & ~x522;
assign c3120 =  x44 & ~x178 & ~x306 & ~x403 & ~x543;
assign c3122 = ~x60 & ~x298 & ~x374 & ~x379 & ~x380 & ~x402 & ~x431 & ~x450 & ~x479 & ~x507 & ~x538 & ~x563 & ~x564 & ~x570 & ~x612 & ~x664 & ~x726 & ~x745 & ~x749 & ~x755 & ~x779;
assign c3124 =  x585 & ~x580;
assign c3126 =  x306 &  x334 & ~x411 & ~x413 & ~x489;
assign c3128 =  x47 &  x413 & ~x349 & ~x419;
assign c3130 =  x383 &  x635 &  x691 & ~x51 & ~x65 & ~x673 & ~x757;
assign c3132 =  x216 &  x267 & ~x8 & ~x34 & ~x385 & ~x546;
assign c3134 =  x734 & ~x363 & ~x373 & ~x400 & ~x728;
assign c3136 = ~x34 & ~x60 & ~x88 & ~x111 & ~x113 & ~x144 & ~x167 & ~x170 & ~x180 & ~x190 & ~x218 & ~x219 & ~x220 & ~x225 & ~x249 & ~x282 & ~x306 & ~x334 & ~x366 & ~x368 & ~x422 & ~x451 & ~x476 & ~x499 & ~x531 & ~x555 & ~x583 & ~x617 & ~x642 & ~x653 & ~x704 & ~x707 & ~x710;
assign c3138 =  x238 &  x239 & ~x251 & ~x327 & ~x384 & ~x461 & ~x466 & ~x521;
assign c3140 =  x584 & ~x469 & ~x580 & ~x624;
assign c3142 =  x107 &  x332;
assign c3144 =  x45 & ~x80 & ~x306 & ~x334 & ~x587 & ~x737;
assign c3146 =  x294 & ~x159 & ~x278 & ~x329 & ~x405 & ~x520 & ~x599;
assign c3148 =  x145 & ~x14 & ~x52 & ~x120 & ~x279 & ~x288 & ~x318 & ~x518 & ~x584 & ~x782;
assign c3150 =  x443 &  x470 &  x498 & ~x59 & ~x87 & ~x384 & ~x458 & ~x518 & ~x557;
assign c3152 =  x291 &  x525 & ~x88 & ~x439 & ~x466 & ~x490 & ~x668 & ~x703;
assign c3154 =  x551 & ~x109 & ~x493 & ~x507 & ~x539 & ~x549 & ~x682;
assign c3156 =  x245 &  x494 & ~x178 & ~x306 & ~x614 & ~x639;
assign c3158 =  x156 & ~x34 & ~x52 & ~x86 & ~x269 & ~x378 & ~x476 & ~x486 & ~x532 & ~x542 & ~x571 & ~x585 & ~x641 & ~x645;
assign c3160 =  x247 & ~x7 & ~x168 & ~x254 & ~x306 & ~x353 & ~x433 & ~x572 & ~x757;
assign c3162 =  x579 & ~x5 & ~x173 & ~x249 & ~x306 & ~x508 & ~x532 & ~x542 & ~x544 & ~x587 & ~x601;
assign c3164 =  x220 & ~x167 & ~x385;
assign c3166 =  x267 &  x268 &  x294 & ~x58 & ~x380 & ~x414 & ~x489 & ~x542 & ~x574;
assign c3168 =  x442 &  x524 &  x551 & ~x78 & ~x196 & ~x640 & ~x664;
assign c3170 =  x385 &  x509 &  x637 & ~x392;
assign c3172 =  x157 &  x539 & ~x25 & ~x124 & ~x141 & ~x533 & ~x559 & ~x639;
assign c3174 =  x444 &  x501 &  x668 & ~x118;
assign c3176 =  x696 & ~x496;
assign c3178 = ~x124 & ~x130 & ~x402 & ~x469 & ~x470 & ~x605 & ~x628 & ~x739;
assign c3180 = ~x9 & ~x94 & ~x163 & ~x167 & ~x193 & ~x219 & ~x242 & ~x249 & ~x303 & ~x341 & ~x548 & ~x549 & ~x699 & ~x711 & ~x749;
assign c3182 =  x552 &  x580 &  x608 & ~x306 & ~x466 & ~x535 & ~x669 & ~x710;
assign c3184 = ~x5 & ~x60 & ~x191 & ~x301 & ~x414 & ~x441 & ~x465 & ~x467 & ~x470 & ~x496 & ~x521 & ~x622 & ~x623 & ~x731;
assign c3186 =  x128 &  x156 &  x524 & ~x542 & ~x598 & ~x729;
assign c3188 =  x74 & ~x113 & ~x166 & ~x167 & ~x181 & ~x320 & ~x560;
assign c3190 =  x494 & ~x194 & ~x261 & ~x431;
assign c3192 =  x102 &  x129 & ~x7 & ~x225 & ~x226 & ~x432 & ~x560 & ~x585;
assign c3194 =  x497 &  x524 & ~x2 & ~x59 & ~x75 & ~x163 & ~x422 & ~x598 & ~x703;
assign c3196 =  x444 & ~x199;
assign c3198 =  x24;
assign c3200 =  x585 & ~x493 & ~x498;
assign c3202 =  x770 & ~x249 & ~x488 & ~x517 & ~x629 & ~x682 & ~x710;
assign c3204 =  x233 & ~x34 & ~x90 & ~x174 & ~x198 & ~x227 & ~x306 & ~x363 & ~x465 & ~x545 & ~x546 & ~x622 & ~x643 & ~x680 & ~x751;
assign c3206 =  x239 &  x240 & ~x412 & ~x440 & ~x464 & ~x469 & ~x691 & ~x739;
assign c3208 =  x385 &  x721 & ~x1 & ~x114 & ~x222 & ~x350;
assign c3210 =  x193 & ~x139 & ~x299 & ~x328 & ~x352 & ~x354 & ~x376 & ~x380 & ~x382 & ~x403 & ~x404 & ~x431 & ~x448 & ~x481;
assign c3212 =  x366 & ~x355 & ~x467 & ~x521;
assign c3214 =  x359 &  x666;
assign c3216 =  x723 & ~x495;
assign c3218 =  x247 &  x734;
assign c3220 =  x579 &  x607 & ~x143 & ~x197 & ~x227 & ~x228 & ~x255 & ~x275 & ~x282 & ~x304 & ~x306 & ~x701 & ~x705 & ~x706;
assign c3222 =  x218 &  x470 & ~x81 & ~x278 & ~x336 & ~x405 & ~x434 & ~x461 & ~x505 & ~x534 & ~x643 & ~x672 & ~x697 & ~x728;
assign c3224 =  x132 &  x161 &  x385 & ~x166 & ~x588;
assign c3226 =  x73 &  x157 & ~x66 & ~x306 & ~x546;
assign c3228 =  x162 & ~x244 & ~x530 & ~x540;
assign c3230 = ~x8 & ~x56 & ~x89 & ~x130 & ~x133 & ~x229 & ~x255 & ~x382 & ~x405 & ~x432 & ~x434 & ~x465 & ~x505 & ~x535 & ~x546 & ~x570 & ~x670 & ~x700 & ~x701 & ~x727;
assign c3232 =  x186 &  x211 & ~x16 & ~x327;
assign c3234 =  x498 & ~x327 & ~x396 & ~x476 & ~x585 & ~x592 & ~x594 & ~x624 & ~x677 & ~x701 & ~x704 & ~x772 & ~x774;
assign c3236 =  x334 & ~x274 & ~x431 & ~x588 & ~x715;
assign c3238 =  x748 & ~x57 & ~x599;
assign c3240 =  x214 &  x706 & ~x1 & ~x376 & ~x431 & ~x487;
assign c3242 =  x205 &  x316 & ~x34 & ~x52 & ~x139 & ~x166 & ~x546 & ~x556 & ~x588 & ~x672 & ~x704 & ~x758;
assign c3244 = ~x92 & ~x106 & ~x134 & ~x135 & ~x174 & ~x467 & ~x518 & ~x521 & ~x561 & ~x563 & ~x598 & ~x672 & ~x725 & ~x762;
assign c3246 = ~x36 & ~x71 & ~x193 & ~x263 & ~x308 & ~x363 & ~x368 & ~x395 & ~x422 & ~x466 & ~x503 & ~x507 & ~x545 & ~x546 & ~x547 & ~x598 & ~x602 & ~x678 & ~x709;
assign c3248 =  x528 & ~x440 & ~x498 & ~x521 & ~x580;
assign c3250 =  x556 & ~x226 & ~x358 & ~x440 & ~x465 & ~x467;
assign c3252 =  x129 &  x635 & ~x37 & ~x113 & ~x168 & ~x226 & ~x505 & ~x561 & ~x618 & ~x703;
assign c3254 =  x277 & ~x1 & ~x45 & ~x196 & ~x357 & ~x384 & ~x434 & ~x513 & ~x514 & ~x515 & ~x588 & ~x692 & ~x693;
assign c3256 = ~x28 & ~x29 & ~x321 & ~x326 & ~x344 & ~x374 & ~x407 & ~x422 & ~x424 & ~x426 & ~x431 & ~x457 & ~x482 & ~x560 & ~x716 & ~x717 & ~x750;
assign c3258 =  x320 &  x501 & ~x570;
assign c3260 =  x498 & ~x253 & ~x412 & ~x466 & ~x495 & ~x674;
assign c3262 =  x218;
assign c3264 =  x268 & ~x1 & ~x19 & ~x95 & ~x191 & ~x249 & ~x253 & ~x255 & ~x278 & ~x309 & ~x470 & ~x503 & ~x570;
assign c3266 =  x324 & ~x92 & ~x166 & ~x459 & ~x519 & ~x573 & ~x576 & ~x656 & ~x739;
assign c3268 = ~x311 & ~x405 & ~x416 & ~x459 & ~x460 & ~x503 & ~x526 & ~x534 & ~x562 & ~x583 & ~x608;
assign c3270 =  x529 & ~x33 & ~x440 & ~x466 & ~x541 & ~x571;
assign c3272 =  x77 &  x219;
assign c3274 =  x323 & ~x155 & ~x216 & ~x657;
assign c3276 =  x384 &  x411 &  x465 &  x466 & ~x66 & ~x392 & ~x433;
assign c3278 =  x501 &  x590;
assign c3280 =  x584 &  x612 & ~x200 & ~x467 & ~x496;
assign c3282 =  x411 &  x635 &  x663 & ~x153 & ~x227 & ~x307 & ~x639 & ~x657;
assign c3284 =  x580 &  x608 & ~x89 & ~x113 & ~x117 & ~x165 & ~x168 & ~x255 & ~x437 & ~x546 & ~x561 & ~x699 & ~x708 & ~x723 & ~x760;
assign c3286 =  x501 & ~x384 & ~x387 & ~x467 & ~x496;
assign c3288 =  x334 & ~x303 & ~x327 & ~x350 & ~x403;
assign c3290 =  x192 &  x276 & ~x354 & ~x427 & ~x449;
assign c3292 =  x526 & ~x85 & ~x89 & ~x167 & ~x327 & ~x383 & ~x406 & ~x436 & ~x506 & ~x532 & ~x585 & ~x587 & ~x620 & ~x641 & ~x645 & ~x648 & ~x729;
assign c3294 =  x243 &  x423 & ~x490 & ~x546 & ~x598 & ~x700 & ~x727;
assign c3296 =  x294 & ~x50 & ~x75 & ~x170 & ~x280 & ~x281 & ~x384 & ~x431 & ~x457 & ~x671 & ~x683;
assign c3298 =  x678 & ~x95 & ~x178 & ~x261 & ~x475 & ~x500 & ~x561 & ~x669 & ~x696 & ~x711;
assign c3300 =  x233 &  x316 & ~x63 & ~x82 & ~x86 & ~x137 & ~x190 & ~x199 & ~x250 & ~x365 & ~x476 & ~x571 & ~x734 & ~x782;
assign c3302 =  x326 &  x606 &  x662 & ~x545 & ~x574;
assign c3304 =  x221 &  x445 & ~x486;
assign c3306 =  x697;
assign c3308 =  x267 &  x579 & ~x135 & ~x375 & ~x376 & ~x460 & ~x616;
assign c3310 =  x299 &  x635 & ~x106 & ~x194 & ~x665;
assign c3312 =  x438 &  x678 & ~x376 & ~x527;
assign c3314 =  x328 &  x637 & ~x5 & ~x278 & ~x306 & ~x363 & ~x572 & ~x642 & ~x734;
assign c3316 =  x129 &  x156 & ~x14 & ~x53 & ~x110 & ~x242 & ~x319 & ~x475 & ~x488 & ~x491 & ~x517 & ~x670 & ~x698;
assign c3318 =  x326 &  x327 &  x378 & ~x250;
assign c3320 =  x44 & ~x264 & ~x570 & ~x774;
assign c3322 =  x356 &  x357 &  x383 &  x384 &  x411 & ~x498 & ~x754;
assign c3324 =  x288 &  x316 & ~x175 & ~x611 & ~x629 & ~x735;
assign c3326 = ~x110 & ~x243 & ~x354 & ~x376 & ~x426 & ~x505 & ~x512 & ~x513 & ~x515 & ~x531 & ~x570 & ~x594 & ~x646 & ~x690 & ~x692 & ~x746 & ~x774;
assign c3328 =  x583 &  x611 & ~x61 & ~x141 & ~x199 & ~x440 & ~x608;
assign c3330 =  x391 & ~x440;
assign c3332 =  x537 & ~x212 & ~x466 & ~x467 & ~x521 & ~x523 & ~x549 & ~x571 & ~x680;
assign c3334 =  x638 & ~x466 & ~x467 & ~x522 & ~x580 & ~x607 & ~x674;
assign c3336 =  x764;
assign c3338 = ~x25 & ~x60 & ~x291 & ~x327 & ~x354 & ~x380 & ~x400 & ~x408 & ~x423 & ~x427 & ~x478 & ~x596 & ~x615 & ~x674 & ~x721 & ~x726 & ~x748 & ~x754;
assign c3340 =  x501 & ~x469 & ~x470 & ~x523;
assign c3342 =  x103 &  x158 & ~x141 & ~x278 & ~x306 & ~x504 & ~x587 & ~x646 & ~x739;
assign c3344 =  x771 & ~x68 & ~x95;
assign c3346 =  x706 & ~x10 & ~x92 & ~x404 & ~x587;
assign c3348 =  x211 & ~x97 & ~x114 & ~x348 & ~x375 & ~x519 & ~x556 & ~x585 & ~x612 & ~x617 & ~x682;
assign c3350 =  x278 &  x306 &  x334 & ~x116 & ~x330 & ~x377 & ~x439 & ~x486 & ~x541;
assign c3352 =  x585 & ~x86 & ~x470 & ~x522;
assign c3354 =  x317 & ~x119 & ~x176 & ~x284 & ~x465 & ~x466 & ~x510 & ~x543 & ~x629 & ~x661;
assign c3356 =  x418 & ~x143 & ~x467 & ~x509 & ~x515 & ~x535;
assign c3358 =  x499 & ~x327 & ~x328 & ~x406 & ~x496;
assign c3360 =  x498 & ~x113 & ~x380 & ~x384 & ~x410 & ~x466 & ~x467 & ~x520 & ~x529 & ~x546 & ~x548 & ~x562;
assign c3362 =  x528 & ~x273 & ~x327 & ~x466;
assign c3364 = ~x3 & ~x168 & ~x216 & ~x273 & ~x353 & ~x383 & ~x435 & ~x465 & ~x484 & ~x485 & ~x486 & ~x535 & ~x537 & ~x587 & ~x642 & ~x670 & ~x772;
assign c3366 =  x527 & ~x492 & ~x521 & ~x534;
assign c3368 = ~x57 & ~x130 & ~x141 & ~x170 & ~x172 & ~x256 & ~x273 & ~x436 & ~x467 & ~x470 & ~x519 & ~x523 & ~x560 & ~x598 & ~x652 & ~x680 & ~x741 & ~x756;
assign c3370 =  x441 & ~x167 & ~x376 & ~x507 & ~x517 & ~x543 & ~x560 & ~x585 & ~x610 & ~x772;
assign c3372 =  x278 & ~x377 & ~x384 & ~x431 & ~x508;
assign c3374 =  x331 &  x499 & ~x466 & ~x589;
assign c3376 =  x160 &  x357 &  x384 &  x412 &  x440 & ~x586;
assign c3378 =  x721 & ~x306 & ~x607 & ~x716;
assign c3380 =  x157 &  x158 &  x650 & ~x95 & ~x668;
assign c3382 =  x762;
assign c3384 =  x241 &  x313 &  x368 & ~x227 & ~x252 & ~x356 & ~x398 & ~x559;
assign c3386 =  x386 &  x414 &  x666 & ~x199 & ~x337 & ~x574 & ~x780 & ~x781;
assign c3388 =  x584 & ~x577 & ~x580;
assign c3390 =  x246 &  x765;
assign c3392 = ~x75 & ~x142 & ~x199 & ~x226 & ~x356 & ~x357 & ~x384 & ~x412 & ~x466 & ~x488 & ~x521 & ~x591 & ~x622 & ~x624 & ~x706 & ~x745 & ~x774;
assign c3394 =  x131 &  x285 & ~x43 & ~x140 & ~x460 & ~x561 & ~x616 & ~x675;
assign c3396 =  x352 &  x439 &  x691;
assign c3398 =  x165 &  x334 & ~x328;
assign c3400 =  x735 & ~x66 & ~x82 & ~x585;
assign c3402 = ~x45 & ~x114 & ~x141 & ~x299 & ~x300 & ~x357 & ~x405 & ~x412 & ~x466 & ~x467 & ~x505 & ~x532 & ~x561 & ~x672 & ~x761;
assign c3404 =  x320 &  x528 & ~x156 & ~x493;
assign c3406 =  x366 & ~x384 & ~x412 & ~x467;
assign c3408 =  x499 &  x526 &  x553 & ~x412 & ~x493 & ~x570 & ~x645;
assign c3410 =  x296 &  x664 & ~x249;
assign c3412 =  x771 & ~x61 & ~x78 & ~x616 & ~x629 & ~x674 & ~x740;
assign c3414 =  x73 &  x101 &  x129 & ~x28 & ~x84 & ~x136 & ~x226 & ~x306 & ~x435 & ~x445 & ~x616 & ~x644 & ~x660 & ~x700 & ~x756;
assign c3416 =  x46 &  x245;
assign c3418 =  x474 & ~x102 & ~x112 & ~x226 & ~x467 & ~x469 & ~x522 & ~x623 & ~x681 & ~x711 & ~x737;
assign c3420 =  x327 &  x662 & ~x181;
assign c3422 =  x499 &  x527 & ~x6 & ~x328 & ~x385 & ~x522 & ~x523 & ~x576 & ~x586 & ~x747;
assign c3424 =  x441 & ~x368 & ~x402 & ~x580 & ~x592;
assign c3426 = ~x203 & ~x402 & ~x541;
assign c3428 =  x320 &  x418 & ~x31;
assign c3430 =  x324 &  x356 & ~x278 & ~x306 & ~x685 & ~x739;
assign c3432 =  x411 &  x466 & ~x137 & ~x305 & ~x319 & ~x432 & ~x612 & ~x637 & ~x668 & ~x729;
assign c3434 =  x250 &  x334 & ~x427;
assign c3436 = ~x36 & ~x60 & ~x63 & ~x168 & ~x198 & ~x229 & ~x276 & ~x338 & ~x422 & ~x424 & ~x450 & ~x478 & ~x518 & ~x528 & ~x545 & ~x573 & ~x575 & ~x588 & ~x601 & ~x669 & ~x681 & ~x701;
assign c3438 =  x501 & ~x141;
assign c3440 =  x357 &  x385 &  x412 &  x466 & ~x641;
assign c3442 =  x636 & ~x78 & ~x242 & ~x306 & ~x307 & ~x310 & ~x656 & ~x725;
assign c3444 =  x317 &  x502 & ~x469 & ~x544;
assign c3446 =  x719 &  x746 & ~x124 & ~x557;
assign c3448 =  x147 &  x158 &  x203 & ~x9 & ~x41 & ~x96 & ~x251 & ~x529 & ~x585 & ~x618;
assign c3450 =  x582 & ~x467 & ~x580 & ~x669;
assign c3452 =  x414 &  x442 &  x443 &  x470 & ~x137 & ~x512 & ~x543 & ~x625 & ~x669 & ~x720;
assign c3454 =  x339 &  x367 &  x705 & ~x1 & ~x470;
assign c3456 =  x556 & ~x196 & ~x468 & ~x470 & ~x496 & ~x522 & ~x576;
assign c3458 =  x73 &  x101 &  x128 & ~x515 & ~x543;
assign c3460 =  x411 &  x412 &  x494 & ~x78;
assign c3462 =  x73 &  x129 &  x328;
assign c3464 =  x414 &  x470 & ~x54 & ~x112 & ~x243 & ~x465 & ~x505 & ~x618 & ~x775;
assign c3466 =  x636 & ~x69 & ~x278 & ~x362 & ~x492 & ~x574 & ~x577 & ~x605 & ~x669 & ~x708 & ~x709;
assign c3468 =  x161 &  x357 &  x385 & ~x308 & ~x309 & ~x555 & ~x556 & ~x672;
assign c3470 =  x470 &  x524 &  x551 & ~x465 & ~x513 & ~x515 & ~x537 & ~x561 & ~x643 & ~x726;
assign c3472 = ~x195 & ~x327 & ~x356 & ~x402 & ~x424 & ~x508 & ~x585 & ~x646;
assign c3474 =  x706 & ~x178;
assign c3476 = ~x7 & ~x217 & ~x412 & ~x433 & ~x458 & ~x467 & ~x513 & ~x519 & ~x626 & ~x657 & ~x669;
assign c3478 =  x350 & ~x132 & ~x159 & ~x184 & ~x212 & ~x215 & ~x466 & ~x489 & ~x492 & ~x709;
assign c3480 =  x276 & ~x327 & ~x371 & ~x434 & ~x487 & ~x517 & ~x559;
assign c3482 =  x691;
assign c3484 =  x305 &  x501 & ~x495 & ~x515 & ~x719;
assign c3486 =  x356 &  x408 & ~x221 & ~x279;
assign c3488 =  x44 & ~x207 & ~x292 & ~x320 & ~x515 & ~x729 & ~x743;
assign c3490 =  x395 &  x423 & ~x157 & ~x384 & ~x386 & ~x463 & ~x467;
assign c3492 =  x191 &  x219 &  x247 & ~x308 & ~x344 & ~x580;
assign c3494 =  x443 &  x470 & ~x243 & ~x356 & ~x451 & ~x611;
assign c3496 =  x73 &  x128 & ~x376 & ~x672 & ~x680;
assign c3498 =  x353 & ~x84 & ~x237 & ~x278 & ~x293 & ~x470 & ~x472 & ~x516 & ~x571 & ~x670 & ~x682 & ~x776;
assign c31 =  x150 &  x151 &  x179 & ~x1 & ~x169 & ~x303 & ~x445;
assign c33 =  x269 & ~x82 & ~x110 & ~x201 & ~x285 & ~x342 & ~x361 & ~x702 & ~x725 & ~x747;
assign c35 =  x269 &  x409 & ~x482 & ~x537 & ~x719 & ~x766;
assign c37 =  x659 &  x660 &  x687 & ~x87 & ~x307 & ~x363 & ~x760 & ~x764 & ~x768;
assign c39 =  x598 &  x599;
assign c311 =  x301 &  x330 &  x472 & ~x635;
assign c313 =  x425 &  x534 & ~x70 & ~x459 & ~x660 & ~x684 & ~x700 & ~x720 & ~x736 & ~x740 & ~x753;
assign c315 =  x200 &  x509;
assign c317 = ~x126 & ~x180 & ~x235 & ~x325 & ~x466 & ~x613 & ~x630 & ~x642 & ~x722 & ~x759 & ~x769;
assign c319 = ~x27 & ~x143 & ~x145 & ~x247 & ~x258 & ~x278 & ~x286 & ~x287 & ~x315 & ~x316 & ~x386 & ~x392 & ~x396 & ~x397 & ~x444 & ~x505 & ~x586 & ~x614 & ~x618 & ~x669;
assign c321 = ~x46 & ~x93 & ~x173 & ~x258 & ~x259 & ~x285 & ~x368 & ~x393 & ~x396 & ~x416 & ~x425 & ~x470 & ~x480 & ~x534 & ~x556 & ~x777;
assign c323 =  x404 & ~x55 & ~x481 & ~x672;
assign c325 =  x124 &  x153 &  x689 &  x716;
assign c327 =  x547 & ~x0 & ~x60 & ~x137 & ~x190 & ~x192 & ~x221 & ~x475 & ~x622 & ~x705;
assign c329 =  x433 & ~x310 & ~x588;
assign c331 =  x343 &  x400 & ~x129;
assign c333 =  x201 &  x231 &  x258 &  x259 & ~x43;
assign c335 =  x543 & ~x48 & ~x75 & ~x136;
assign c337 = ~x34 & ~x173 & ~x286 & ~x341 & ~x365 & ~x399 & ~x481 & ~x483 & ~x509 & ~x732;
assign c339 =  x425 & ~x70 & ~x324 & ~x401 & ~x484;
assign c341 =  x213 &  x547 & ~x622 & ~x731 & ~x736;
assign c343 =  x619 & ~x40 & ~x43 & ~x166 & ~x388 & ~x733;
assign c345 =  x487 & ~x695 & ~x722 & ~x774;
assign c347 =  x544 & ~x103 & ~x195;
assign c349 =  x460 &  x488;
assign c351 =  x490;
assign c353 =  x478 & ~x93 & ~x239 & ~x294;
assign c355 =  x677 & ~x222 & ~x339 & ~x460 & ~x745;
assign c357 =  x627 &  x655 & ~x7 & ~x734;
assign c359 =  x491 &  x519 &  x547;
assign c361 =  x275 & ~x19 & ~x267 & ~x350 & ~x598 & ~x622 & ~x768;
assign c363 = ~x103 & ~x150 & ~x267 & ~x269 & ~x379 & ~x581 & ~x719 & ~x764;
assign c365 =  x312 &  x397 & ~x6 & ~x10 & ~x58 & ~x96 & ~x98 & ~x205 & ~x208 & ~x290 & ~x628 & ~x720 & ~x767;
assign c367 =  x483 &  x566 & ~x73 & ~x97 & ~x181 & ~x490 & ~x716;
assign c369 =  x514 & ~x46;
assign c371 =  x432 & ~x11 & ~x564 & ~x693;
assign c373 =  x171;
assign c375 = ~x51 & ~x169 & ~x226 & ~x250 & ~x272 & ~x358 & ~x397 & ~x444 & ~x528 & ~x559 & ~x591 & ~x618 & ~x690 & ~x703 & ~x730 & ~x754;
assign c377 =  x314 & ~x210 & ~x263 & ~x770;
assign c379 =  x330 & ~x1 & ~x203 & ~x325 & ~x604 & ~x696 & ~x767;
assign c381 =  x343 &  x427 & ~x324 & ~x365 & ~x461 & ~x602;
assign c383 =  x351 & ~x71 & ~x610 & ~x621 & ~x634 & ~x635 & ~x662;
assign c385 =  x491 & ~x26 & ~x75 & ~x700 & ~x767;
assign c387 =  x673 & ~x70 & ~x71;
assign c389 =  x409 & ~x2 & ~x359 & ~x454 & ~x481 & ~x510 & ~x538 & ~x581 & ~x635 & ~x647 & ~x704;
assign c391 =  x533 & ~x108 & ~x295 & ~x434 & ~x722;
assign c393 =  x321 &  x430 &  x484 & ~x224;
assign c395 = ~x16 & ~x36 & ~x43 & ~x44 & ~x57 & ~x75 & ~x84 & ~x113 & ~x114 & ~x126 & ~x180 & ~x265 & ~x392 & ~x486 & ~x487 & ~x575 & ~x624 & ~x658 & ~x659 & ~x662 & ~x716 & ~x717 & ~x725 & ~x777;
assign c397 =  x485 &  x511 &  x648 & ~x360;
assign c399 =  x520 & ~x46 & ~x127 & ~x359 & ~x770;
assign c3101 =  x571 &  x572 & ~x75;
assign c3103 =  x236 &  x382 & ~x565 & ~x760;
assign c3105 =  x427 &  x456 &  x566 & ~x406;
assign c3107 =  x623 & ~x24 & ~x26 & ~x201 & ~x304 & ~x333 & ~x388 & ~x390 & ~x547 & ~x717 & ~x719 & ~x745 & ~x749;
assign c3109 =  x546 & ~x53 & ~x78 & ~x108 & ~x137 & ~x363 & ~x484 & ~x566 & ~x700 & ~x703 & ~x757;
assign c3111 =  x398 &  x425 & ~x178 & ~x207;
assign c3113 =  x269 & ~x170 & ~x313 & ~x334 & ~x342 & ~x359 & ~x391 & ~x397 & ~x421 & ~x424;
assign c3115 =  x459 & ~x534 & ~x636 & ~x722;
assign c3117 =  x564 & ~x43 & ~x70 & ~x351 & ~x358 & ~x379 & ~x773;
assign c3119 =  x148 &  x149 & ~x10 & ~x43;
assign c3121 =  x314 & ~x70 & ~x236 & ~x380 & ~x574 & ~x656 & ~x741 & ~x748 & ~x777;
assign c3123 =  x484 &  x620 & ~x479;
assign c3125 =  x236 &  x263 &  x689 & ~x561 & ~x767;
assign c3127 =  x573 & ~x20 & ~x160 & ~x761;
assign c3129 =  x228 &  x401;
assign c3131 =  x210 &  x492 & ~x160 & ~x752;
assign c3133 =  x321 &  x430 &  x457;
assign c3135 =  x396 & ~x93 & ~x263 & ~x270 & ~x354 & ~x722;
assign c3137 =  x152 &  x488;
assign c3139 =  x304 & ~x19 & ~x48 & ~x82 & ~x184 & ~x319 & ~x326 & ~x548;
assign c3141 =  x154 &  x321 & ~x85 & ~x564;
assign c3143 =  x177 &  x484 & ~x26 & ~x360;
assign c3145 = ~x70 & ~x84 & ~x100 & ~x180 & ~x211 & ~x213 & ~x267 & ~x348 & ~x356 & ~x778;
assign c3147 =  x352 & ~x27 & ~x118 & ~x593 & ~x612 & ~x633 & ~x637 & ~x662;
assign c3149 =  x620 &  x674;
assign c3151 =  x64 & ~x305 & ~x658 & ~x661;
assign c3153 =  x402 &  x431 & ~x481;
assign c3155 = ~x45 & ~x79 & ~x98 & ~x152 & ~x294 & ~x375 & ~x632 & ~x721;
assign c3157 =  x122 &  x150 &  x151 & ~x26 & ~x80 & ~x171 & ~x533;
assign c3159 =  x304 &  x417 & ~x355;
assign c3161 =  x516 &  x517 & ~x46;
assign c3163 =  x483 &  x623 & ~x434;
assign c3165 =  x181 & ~x11 & ~x228 & ~x390 & ~x591;
assign c3167 =  x227 &  x427;
assign c3169 =  x460 & ~x554;
assign c3171 =  x260 &  x428 &  x456 & ~x19 & ~x46 & ~x351 & ~x448;
assign c3173 =  x543 &  x571 &  x572;
assign c3175 =  x430 &  x675;
assign c3177 = ~x23 & ~x397 & ~x399 & ~x446 & ~x481 & ~x591 & ~x717;
assign c3179 =  x548 &  x714;
assign c3181 =  x397 & ~x16 & ~x93 & ~x234 & ~x236 & ~x637 & ~x692 & ~x741;
assign c3183 =  x321 &  x349 & ~x12 & ~x581 & ~x590 & ~x698;
assign c3185 = ~x89 & ~x140 & ~x174 & ~x202 & ~x204 & ~x224 & ~x229 & ~x246 & ~x248 & ~x253 & ~x260 & ~x283 & ~x306 & ~x397 & ~x418 & ~x419 & ~x427 & ~x456 & ~x460 & ~x473 & ~x474 & ~x489 & ~x498 & ~x531 & ~x640 & ~x644 & ~x751 & ~x755 & ~x762;
assign c3187 = ~x91 & ~x140 & ~x193 & ~x254 & ~x284 & ~x286 & ~x317 & ~x339 & ~x343 & ~x360 & ~x368 & ~x540 & ~x561 & ~x587 & ~x671 & ~x673;
assign c3189 =  x149 &  x631 & ~x77 & ~x479;
assign c3191 =  x485 &  x512 &  x621 & ~x777;
assign c3193 = ~x24 & ~x70 & ~x100 & ~x125 & ~x236 & ~x449 & ~x693 & ~x744 & ~x779;
assign c3195 =  x507 & ~x70 & ~x325 & ~x708 & ~x717 & ~x770 & ~x772;
assign c3197 =  x231 &  x400 &  x427 & ~x80;
assign c3199 =  x64 &  x428;
assign c3201 =  x428 &  x674;
assign c3203 =  x681 &  x712 & ~x104;
assign c3205 = ~x48 & ~x75 & ~x97 & ~x100 & ~x192 & ~x359 & ~x388 & ~x559 & ~x687;
assign c3207 =  x69 &  x97 & ~x59 & ~x103 & ~x142 & ~x447 & ~x509;
assign c3209 = ~x19 & ~x46 & ~x73 & ~x236 & ~x239 & ~x267 & ~x382 & ~x431 & ~x570 & ~x601 & ~x721 & ~x724 & ~x768 & ~x770;
assign c3211 =  x520 &  x549 & ~x359 & ~x652 & ~x728 & ~x765 & ~x767;
assign c3213 =  x181 &  x182 &  x210 & ~x51 & ~x174 & ~x502;
assign c3215 =  x625 &  x712;
assign c3217 =  x603 &  x604 &  x631 &  x660 & ~x82 & ~x337 & ~x561 & ~x657 & ~x739;
assign c3219 =  x712;
assign c3221 =  x150 &  x457 & ~x102;
assign c3223 =  x425 & ~x16 & ~x235 & ~x322 & ~x689 & ~x747 & ~x770;
assign c3225 =  x510 &  x564 & ~x268;
assign c3227 =  x321 &  x430 &  x457;
assign c3229 =  x171 &  x257;
assign c3231 =  x274 &  x330 &  x360 & ~x713;
assign c3233 =  x534 & ~x37 & ~x70 & ~x75 & ~x150 & ~x180 & ~x206 & ~x657 & ~x751 & ~x765;
assign c3235 =  x311 &  x564;
assign c3237 =  x346 & ~x426 & ~x452 & ~x502 & ~x554 & ~x581;
assign c3239 =  x436 & ~x421 & ~x482 & ~x534 & ~x564 & ~x708 & ~x736;
assign c3241 =  x653 &  x683;
assign c3243 =  x229 &  x314 & ~x16;
assign c3245 =  x65 &  x93 & ~x17 & ~x60 & ~x250 & ~x301 & ~x471;
assign c3247 =  x370 & ~x103 & ~x345 & ~x351 & ~x630 & ~x776;
assign c3249 =  x453 & ~x103 & ~x125 & ~x160 & ~x405 & ~x433 & ~x572 & ~x660 & ~x706 & ~x736;
assign c3251 =  x463 & ~x20 & ~x80 & ~x142 & ~x415 & ~x427 & ~x476 & ~x566 & ~x721 & ~x729;
assign c3253 =  x432 & ~x309 & ~x535 & ~x767;
assign c3255 =  x69 &  x154 & ~x144;
assign c3257 =  x388 & ~x66 & ~x70 & ~x93 & ~x136 & ~x262 & ~x326 & ~x383 & ~x406 & ~x459 & ~x654;
assign c3259 =  x177 &  x400 &  x565 & ~x110 & ~x138 & ~x489;
assign c3261 =  x397 &  x533;
assign c3263 =  x293 & ~x252 & ~x286 & ~x420 & ~x506;
assign c3265 =  x487 &  x515 & ~x749;
assign c3267 =  x519 & ~x194 & ~x419 & ~x456 & ~x509 & ~x532 & ~x623 & ~x724 & ~x754;
assign c3269 =  x409 & ~x91 & ~x173 & ~x452 & ~x529 & ~x558 & ~x581;
assign c3271 = ~x143 & ~x219 & ~x227 & ~x313 & ~x473 & ~x475 & ~x483 & ~x525 & ~x538 & ~x553 & ~x556 & ~x581 & ~x584 & ~x591 & ~x778;
assign c3273 = ~x145 & ~x172 & ~x233 & ~x258 & ~x286 & ~x313 & ~x337 & ~x359 & ~x444 & ~x455 & ~x583 & ~x695 & ~x696 & ~x731;
assign c3275 =  x599 & ~x75 & ~x115;
assign c3277 =  x458 &  x485 &  x512 &  x567;
assign c3279 =  x209 & ~x3 & ~x32 & ~x64 & ~x88 & ~x414 & ~x473 & ~x538 & ~x563 & ~x617;
assign c3281 =  x304 & ~x178 & ~x236 & ~x291 & ~x294 & ~x325 & ~x706;
assign c3283 =  x66 & ~x24 & ~x217 & ~x359 & ~x360 & ~x393;
assign c3285 =  x400 &  x401 & ~x180 & ~x390 & ~x391;
assign c3287 = ~x6 & ~x27 & ~x29 & ~x43 & ~x103 & ~x105 & ~x120 & ~x126 & ~x194 & ~x323 & ~x336 & ~x364 & ~x381 & ~x392 & ~x461 & ~x466 & ~x549 & ~x630 & ~x700 & ~x750;
assign c3289 =  x66 &  x623 & ~x19 & ~x24 & ~x55 & ~x143 & ~x275 & ~x361 & ~x700;
assign c3291 =  x175 & ~x0 & ~x183 & ~x365 & ~x682 & ~x701 & ~x757;
assign c3293 =  x312 &  x398 & ~x45 & ~x571 & ~x714 & ~x770;
assign c3295 =  x547 & ~x8 & ~x79 & ~x117 & ~x482 & ~x649 & ~x672 & ~x760 & ~x767;
assign c3297 =  x269 &  x492 & ~x25 & ~x30 & ~x559 & ~x595 & ~x598 & ~x736 & ~x764;
assign c3299 = ~x93 & ~x260 & ~x272 & ~x372 & ~x541;
assign c3301 =  x517 & ~x75;
assign c3303 =  x231 &  x427 & ~x40 & ~x726 & ~x767;
assign c3305 =  x509 & ~x42 & ~x46 & ~x180 & ~x325;
assign c3307 =  x314 &  x533;
assign c3309 =  x314 & ~x126 & ~x268 & ~x269 & ~x406 & ~x713 & ~x773;
assign c3311 =  x453 &  x507 & ~x181 & ~x207 & ~x235;
assign c3313 =  x407 & ~x57 & ~x230 & ~x252 & ~x474 & ~x482 & ~x509 & ~x538 & ~x589;
assign c3315 = ~x23 & ~x48 & ~x147 & ~x173 & ~x246 & ~x260 & ~x276 & ~x358 & ~x369 & ~x384 & ~x391 & ~x396 & ~x400 & ~x426 & ~x459 & ~x498 & ~x515 & ~x586;
assign c3317 =  x567 & ~x57 & ~x74 & ~x75 & ~x769;
assign c3319 =  x514 & ~x113 & ~x481 & ~x504;
assign c3321 =  x229 &  x314 & ~x182;
assign c3323 =  x518 & ~x5 & ~x308 & ~x535 & ~x561 & ~x617 & ~x641 & ~x707 & ~x731 & ~x760 & ~x763;
assign c3325 =  x545 & ~x79 & ~x224 & ~x613 & ~x778;
assign c3327 =  x427 &  x428 &  x595 & ~x365;
assign c3329 =  x533 & ~x16 & ~x42 & ~x69 & ~x150 & ~x750 & ~x753 & ~x777;
assign c3331 =  x463 & ~x2 & ~x55 & ~x81 & ~x115 & ~x196 & ~x482 & ~x533 & ~x589 & ~x679 & ~x704 & ~x707 & ~x733 & ~x763;
assign c3333 =  x369 &  x452 & ~x122 & ~x576 & ~x715 & ~x765;
assign c3335 = ~x22 & ~x228 & ~x313 & ~x342 & ~x391 & ~x414 & ~x484 & ~x663 & ~x730;
assign c3337 =  x453 & ~x46 & ~x180 & ~x268 & ~x406;
assign c3339 =  x256 &  x314 & ~x654;
assign c3341 =  x436 & ~x119 & ~x509 & ~x570 & ~x595 & ~x736 & ~x751 & ~x761;
assign c3343 =  x269 & ~x29 & ~x199 & ~x224 & ~x397 & ~x451 & ~x479 & ~x483 & ~x505 & ~x532 & ~x584 & ~x673 & ~x778;
assign c3345 =  x381 & ~x24 & ~x283 & ~x311 & ~x428 & ~x533 & ~x540 & ~x582 & ~x583 & ~x593 & ~x704;
assign c3347 =  x479 & ~x72 & ~x122 & ~x324 & ~x599;
assign c3349 =  x398 & ~x41 & ~x84 & ~x235 & ~x270 & ~x294 & ~x381 & ~x407 & ~x598 & ~x776;
assign c3351 =  x120 & ~x18 & ~x30 & ~x156 & ~x210 & ~x335 & ~x360 & ~x444 & ~x475 & ~x700 & ~x783;
assign c3353 =  x457 &  x485 & ~x480;
assign c3355 =  x314 &  x425 & ~x43 & ~x70 & ~x323 & ~x769;
assign c3357 =  x38 & ~x80 & ~x416;
assign c3359 =  x491 & ~x6 & ~x46 & ~x224 & ~x280 & ~x473 & ~x532 & ~x707 & ~x760;
assign c3361 =  x489 & ~x8 & ~x9 & ~x20 & ~x109 & ~x337 & ~x559 & ~x563 & ~x589 & ~x707;
assign c3363 = ~x24 & ~x46 & ~x75 & ~x197 & ~x285 & ~x286 & ~x312 & ~x330 & ~x334 & ~x344 & ~x417 & ~x426 & ~x446 & ~x642 & ~x700;
assign c3365 =  x680 & ~x118 & ~x142 & ~x203 & ~x222 & ~x417 & ~x476;
assign c3367 =  x153 &  x410;
assign c3369 =  x345 &  x542;
assign c3371 =  x516 &  x543 & ~x78;
assign c3373 = ~x14 & ~x54 & ~x55 & ~x61 & ~x73 & ~x83 & ~x95 & ~x110 & ~x121 & ~x150 & ~x164 & ~x188 & ~x258 & ~x351 & ~x614 & ~x627 & ~x657 & ~x688;
assign c3375 =  x427 &  x509 &  x536 & ~x322;
assign c3377 =  x573 & ~x107 & ~x706 & ~x777;
assign c3379 =  x301 & ~x18 & ~x24 & ~x53 & ~x74 & ~x103 & ~x351 & ~x524 & ~x598 & ~x771;
assign c3381 =  x396 &  x397 & ~x71 & ~x177 & ~x375 & ~x660 & ~x661 & ~x717 & ~x725 & ~x782;
assign c3383 =  x429 &  x430 & ~x397 & ~x423 & ~x559;
assign c3385 =  x738;
assign c3387 =  x461 & ~x103 & ~x336 & ~x454 & ~x565 & ~x751 & ~x752;
assign c3389 =  x512 &  x594 &  x703;
assign c3391 =  x329 &  x360 & ~x208 & ~x550 & ~x770;
assign c3393 =  x535 & ~x44 & ~x126 & ~x406 & ~x459 & ~x669 & ~x683 & ~x721 & ~x767;
assign c3395 =  x627 & ~x161 & ~x277 & ~x279 & ~x282;
assign c3397 =  x275 &  x304 &  x333 & ~x252 & ~x263 & ~x294 & ~x574 & ~x763 & ~x781;
assign c3399 =  x435 & ~x111 & ~x538 & ~x584 & ~x617 & ~x693 & ~x730;
assign c3401 = ~x9 & ~x16 & ~x36 & ~x39 & ~x41 & ~x73 & ~x81 & ~x139 & ~x210 & ~x253 & ~x336 & ~x378 & ~x517 & ~x587 & ~x737 & ~x743 & ~x761 & ~x768;
assign c3403 =  x461;
assign c3405 =  x325 & ~x34 & ~x257 & ~x397 & ~x482 & ~x641 & ~x754;
assign c3407 =  x425 & ~x178 & ~x325 & ~x662;
assign c3409 =  x314 &  x343 & ~x84 & ~x150 & ~x269 & ~x294 & ~x764;
assign c3411 =  x573 &  x601 & ~x103 & ~x586;
assign c3413 =  x456 &  x483 &  x510 &  x566 & ~x180 & ~x405 & ~x633;
assign c3415 =  x201 &  x314 & ~x267;
assign c3417 =  x427 & ~x20 & ~x26 & ~x213 & ~x322 & ~x716 & ~x777;
assign c3419 =  x124 &  x152 & ~x258 & ~x476 & ~x478 & ~x614;
assign c3421 =  x401 &  x402 &  x429 &  x483;
assign c3423 =  x483 &  x566 & ~x153 & ~x180 & ~x235 & ~x535 & ~x718 & ~x742;
assign c3425 =  x343 &  x510 &  x511 & ~x100 & ~x542;
assign c3427 = ~x18 & ~x111 & ~x126 & ~x180 & ~x208 & ~x236 & ~x267 & ~x268 & ~x485 & ~x655 & ~x693 & ~x718;
assign c3429 =  x231 &  x428 &  x456 & ~x396;
assign c3431 =  x325 &  x352 & ~x133 & ~x302;
assign c3433 =  x66 &  x124;
assign c3435 =  x589 & ~x16 & ~x603 & ~x724 & ~x777;
assign c3437 =  x596 & ~x62 & ~x278 & ~x282 & ~x360 & ~x362 & ~x420 & ~x588 & ~x634 & ~x656 & ~x757 & ~x776;
assign c3439 =  x589 & ~x1 & ~x79 & ~x166 & ~x351 & ~x364 & ~x776;
assign c3441 =  x456 &  x565 &  x593 & ~x235;
assign c3443 =  x571 & ~x300 & ~x763 & ~x769;
assign c3445 =  x483 &  x510 &  x648;
assign c3447 =  x490 & ~x75 & ~x85 & ~x222 & ~x441;
assign c3449 =  x66 &  x95 & ~x73;
assign c3451 =  x180 &  x207 & ~x387 & ~x390 & ~x444 & ~x475 & ~x533 & ~x565 & ~x612 & ~x616;
assign c3453 =  x149 &  x428 & ~x81 & ~x391 & ~x408 & ~x416 & ~x419;
assign c3455 =  x263 & ~x18 & ~x85 & ~x446 & ~x482 & ~x536 & ~x539 & ~x581 & ~x613 & ~x616;
assign c3457 =  x403 &  x430 &  x485 &  x512;
assign c3459 =  x427 &  x456 &  x483 &  x511 & ~x448 & ~x660 & ~x741;
assign c3461 =  x293 & ~x89 & ~x111 & ~x165 & ~x280 & ~x482 & ~x534 & ~x584 & ~x672 & ~x761 & ~x767;
assign c3463 =  x540 &  x596 & ~x269;
assign c3465 =  x269 & ~x247 & ~x337 & ~x388 & ~x397 & ~x420 & ~x540 & ~x587;
assign c3467 =  x425 & ~x294 & ~x324;
assign c3469 =  x404 & ~x372 & ~x480 & ~x537 & ~x640 & ~x717;
assign c3471 =  x518 & ~x18 & ~x88 & ~x466 & ~x595 & ~x643;
assign c3473 = ~x37 & ~x77 & ~x229 & ~x279 & ~x280 & ~x341 & ~x358 & ~x365 & ~x370 & ~x401 & ~x427 & ~x450 & ~x535 & ~x557 & ~x646;
assign c3475 =  x120 &  x149 &  x150 & ~x29 & ~x79;
assign c3477 = ~x19 & ~x40 & ~x128 & ~x141 & ~x153 & ~x207 & ~x210 & ~x211 & ~x263 & ~x324 & ~x374 & ~x404 & ~x436 & ~x489 & ~x736 & ~x768;
assign c3479 =  x312 &  x370 &  x564 & ~x777;
assign c3481 =  x229 &  x314 &  x344 & ~x661;
assign c3483 =  x407 & ~x360 & ~x452 & ~x455 & ~x479 & ~x482 & ~x526 & ~x566;
assign c3485 =  x269 & ~x331 & ~x425 & ~x538;
assign c3487 =  x258 &  x259 &  x400 &  x427 & ~x57;
assign c3489 =  x200 &  x314;
assign c3491 =  x417 & ~x70 & ~x147 & ~x148 & ~x149 & ~x553 & ~x664 & ~x693 & ~x724 & ~x741;
assign c3493 =  x390 & ~x150 & ~x179 & ~x214 & ~x642;
assign c3495 =  x182 &  x210 & ~x58 & ~x143 & ~x160 & ~x171 & ~x443 & ~x444;
assign c3497 =  x436 & ~x143 & ~x197 & ~x425 & ~x566 & ~x582 & ~x593 & ~x611 & ~x646;
assign c3499 = ~x17 & ~x75 & ~x178 & ~x199 & ~x213 & ~x350 & ~x581 & ~x661 & ~x696;
assign c40 =  x27;
assign c42 =  x588;
assign c44 =  x122 &  x150 & ~x1 & ~x237 & ~x303 & ~x306 & ~x418 & ~x503 & ~x611 & ~x653 & ~x733 & ~x735 & ~x764;
assign c46 =  x407 &  x491 & ~x60 & ~x171 & ~x221 & ~x225 & ~x227 & ~x266 & ~x450 & ~x503 & ~x662 & ~x663 & ~x708;
assign c48 =  x236 &  x553 &  x581 & ~x144 & ~x620;
assign c410 =  x147 &  x338 &  x624 &  x652;
assign c412 =  x146 &  x393 & ~x69 & ~x154;
assign c414 =  x95 &  x178 &  x179 & ~x105 & ~x143 & ~x345;
assign c416 =  x172 &  x283 & ~x411;
assign c418 =  x574 & ~x0 & ~x155 & ~x437 & ~x439 & ~x465 & ~x468 & ~x475 & ~x503;
assign c420 =  x177 &  x301 &  x357;
assign c422 =  x23;
assign c424 =  x153 &  x519 &  x658;
assign c426 =  x30;
assign c428 =  x549 &  x577 &  x632 & ~x45 & ~x496 & ~x625;
assign c430 =  x264 &  x291 &  x318 &  x345 & ~x86 & ~x109 & ~x199 & ~x225 & ~x246 & ~x275 & ~x303 & ~x405 & ~x700 & ~x701 & ~x728;
assign c432 =  x179 &  x550 & ~x580;
assign c434 =  x257 &  x339 & ~x4 & ~x14 & ~x46 & ~x126 & ~x154 & ~x636 & ~x669;
assign c436 =  x92 &  x122 & ~x14 & ~x26 & ~x44 & ~x70 & ~x166 & ~x587 & ~x588 & ~x669 & ~x706 & ~x732;
assign c438 =  x440 &  x468 &  x579 & ~x106 & ~x508 & ~x677 & ~x725;
assign c440 =  x575 &  x603 &  x630 &  x684 &  x685 & ~x14 & ~x668 & ~x748;
assign c442 =  x549 &  x632 &  x660 & ~x44 & ~x72 & ~x113 & ~x561 & ~x723 & ~x756 & ~x763;
assign c444 =  x550 &  x660 & ~x22 & ~x130 & ~x509 & ~x587;
assign c446 =  x122 &  x491 & ~x111 & ~x237 & ~x763;
assign c448 =  x497 &  x525 & ~x76 & ~x104 & ~x106 & ~x108 & ~x186 & ~x226 & ~x246 & ~x500 & ~x501 & ~x592;
assign c450 =  x228 &  x282 & ~x130 & ~x698;
assign c452 =  x494 &  x633 & ~x14;
assign c454 =  x579 &  x607 &  x689;
assign c456 =  x471 &  x625 & ~x24;
assign c458 =  x28 &  x762;
assign c460 =  x682 & ~x70 & ~x167 & ~x301 & ~x327 & ~x439 & ~x577;
assign c462 =  x105;
assign c464 =  x179 &  x492 &  x520 & ~x1 & ~x87 & ~x100 & ~x534 & ~x675;
assign c466 =  x490 & ~x154 & ~x439 & ~x464 & ~x492 & ~x723 & ~x760;
assign c468 =  x27;
assign c470 =  x264 &  x496 & ~x215 & ~x620;
assign c472 =  x148 &  x625 & ~x70 & ~x491;
assign c474 =  x610 &  x638 & ~x618;
assign c476 =  x499 &  x574;
assign c478 =  x336;
assign c480 =  x284 &  x652 & ~x197 & ~x266 & ~x495 & ~x603;
assign c482 =  x180 &  x497 & ~x396;
assign c484 =  x283 & ~x210 & ~x238 & ~x272 & ~x525 & ~x552 & ~x632;
assign c486 =  x175 &  x284 & ~x399;
assign c488 =  x41 &  x153 &  x181 &  x492;
assign c490 =  x316 &  x371 & ~x209 & ~x210 & ~x237 & ~x279 & ~x321 & ~x330 & ~x332;
assign c492 =  x394 &  x680;
assign c494 =  x523 &  x578 &  x660 & ~x130 & ~x424 & ~x479 & ~x733;
assign c496 =  x181 &  x209 &  x492;
assign c498 =  x492 &  x520 &  x576 &  x631 &  x658 & ~x19 & ~x223 & ~x308 & ~x391 & ~x753;
assign c4100 =  x39 &  x69 &  x497;
assign c4102 =  x632 &  x660 & ~x86 & ~x463 & ~x765;
assign c4104 =  x149 &  x187 &  x243 &  x494;
assign c4106 =  x180 &  x493 & ~x350 & ~x378 & ~x505;
assign c4108 =  x364;
assign c4110 =  x549 &  x632 &  x660 & ~x130 & ~x556 & ~x557 & ~x580 & ~x617 & ~x673;
assign c4112 =  x204 &  x257 & ~x13 & ~x454;
assign c4114 =  x471 & ~x425 & ~x479 & ~x536;
assign c4116 =  x422 & ~x213 & ~x328;
assign c4118 =  x148 & ~x29 & ~x127 & ~x154 & ~x155 & ~x210 & ~x263 & ~x273 & ~x300 & ~x301 & ~x359 & ~x439;
assign c4120 =  x610 & ~x594;
assign c4122 =  x0;
assign c4124 =  x182 &  x209 &  x264 &  x292 &  x319 & ~x28 & ~x87 & ~x170 & ~x218 & ~x275 & ~x359 & ~x448 & ~x503;
assign c4126 =  x490 & ~x72 & ~x143 & ~x248 & ~x275 & ~x309 & ~x410 & ~x478 & ~x479 & ~x533 & ~x548 & ~x555 & ~x556 & ~x563 & ~x584 & ~x588 & ~x610 & ~x614 & ~x645 & ~x670 & ~x694 & ~x728 & ~x747 & ~x761 & ~x776 & ~x778 & ~x781;
assign c4128 =  x123 &  x178 & ~x71 & ~x73 & ~x114 & ~x137 & ~x193 & ~x199 & ~x218 & ~x220 & ~x450 & ~x479 & ~x528 & ~x563 & ~x700 & ~x723;
assign c4132 =  x180 &  x262 & ~x52 & ~x322 & ~x376 & ~x489 & ~x667;
assign c4134 =  x94 &  x188 & ~x168 & ~x197 & ~x237 & ~x617;
assign c4136 =  x208 &  x498 &  x623 & ~x330;
assign c4138 =  x284 &  x338;
assign c4140 =  x39 &  x207 &  x498 & ~x579;
assign c4142 =  x65 & ~x237 & ~x538 & ~x625 & ~x641;
assign c4144 =  x340 &  x651 & ~x663 & ~x664 & ~x748;
assign c4146 =  x1;
assign c4148 =  x628 &  x654 &  x682 & ~x543;
assign c4150 =  x575 &  x603 &  x658 &  x685 & ~x308 & ~x335 & ~x478 & ~x503 & ~x578 & ~x633;
assign c4152 =  x150 &  x178 &  x203 & ~x318;
assign c4154 =  x782;
assign c4156 =  x120 &  x653 &  x654 &  x681;
assign c4158 =  x125 &  x181 & ~x75 & ~x118 & ~x170 & ~x461 & ~x544 & ~x648 & ~x700 & ~x730;
assign c4160 =  x133 &  x148 & ~x154 & ~x156 & ~x249 & ~x385 & ~x413 & ~x468 & ~x554 & ~x695 & ~x722;
assign c4162 =  x65 &  x95 &  x604 & ~x317;
assign c4164 =  x435 & ~x52 & ~x77 & ~x166 & ~x167 & ~x168 & ~x172 & ~x186 & ~x187 & ~x247 & ~x392 & ~x425 & ~x474 & ~x479 & ~x562 & ~x617 & ~x680 & ~x703 & ~x729 & ~x730 & ~x752;
assign c4166 =  x145 & ~x70 & ~x103 & ~x195 & ~x209 & ~x302 & ~x428 & ~x636 & ~x750;
assign c4168 =  x493 &  x521 &  x549 &  x604 &  x631 & ~x74 & ~x158 & ~x528;
assign c4170 =  x26;
assign c4172 =  x523 &  x551 &  x606 &  x661 & ~x501;
assign c4174 =  x627 & ~x170 & ~x494;
assign c4176 =  x347 &  x402 & ~x281 & ~x330 & ~x350 & ~x503 & ~x673 & ~x697;
assign c4178 = ~x29 & ~x266 & ~x293 & ~x301 & ~x328 & ~x329 & ~x349 & ~x376 & ~x415 & ~x431 & ~x440 & ~x441 & ~x473 & ~x498 & ~x527 & ~x557 & ~x581 & ~x720;
assign c4180 =  x153 &  x468;
assign c4182 =  x152 &  x410 &  x605;
assign c4184 =  x120 &  x598 & ~x70 & ~x685;
assign c4186 =  x318 &  x624 & ~x322 & ~x330 & ~x386;
assign c4188 =  x257 &  x652 & ~x13;
assign c4190 =  x662 &  x773 & ~x748;
assign c4192 =  x662 &  x690 &  x773 & ~x433;
assign c4194 =  x153 &  x208 &  x235 & ~x76 & ~x171 & ~x406 & ~x424 & ~x545 & ~x699;
assign c4196 =  x0;
assign c4198 =  x151 &  x179 &  x435 &  x490 & ~x88 & ~x223 & ~x275 & ~x653;
assign c4200 =  x400 & ~x334 & ~x349 & ~x364 & ~x390 & ~x391 & ~x405 & ~x479 & ~x506 & ~x569;
assign c4202 =  x292 &  x581 & ~x214;
assign c4204 =  x346 &  x597 &  x625;
assign c4206 =  x574 & ~x238 & ~x283 & ~x293 & ~x403;
assign c4208 =  x207 &  x292 &  x400 & ~x517;
assign c4210 =  x121 & ~x98 & ~x194 & ~x210 & ~x248 & ~x275 & ~x278 & ~x303 & ~x305 & ~x410 & ~x673 & ~x721 & ~x731;
assign c4212 =  x133 &  x598;
assign c4214 =  x150 & ~x237 & ~x330 & ~x439 & ~x563 & ~x625 & ~x738;
assign c4216 =  x154 &  x181 &  x236 & ~x339 & ~x350 & ~x459;
assign c4218 =  x610 &  x719;
assign c4220 =  x265 &  x578 &  x659 & ~x47;
assign c4222 =  x289 &  x525 & ~x190 & ~x645 & ~x721;
assign c4224 =  x236 &  x469 &  x524;
assign c4226 =  x92 &  x93 &  x94 &  x122 & ~x4 & ~x13 & ~x23 & ~x27 & ~x42 & ~x44 & ~x223 & ~x224 & ~x450 & ~x558 & ~x614;
assign c4228 =  x1 &  x112;
assign c4230 =  x465 &  x493 &  x521 &  x576 &  x603 & ~x23 & ~x52 & ~x130 & ~x478 & ~x563;
assign c4232 =  x97 &  x179 &  x207 & ~x254 & ~x284 & ~x396 & ~x445 & ~x479 & ~x503 & ~x682 & ~x697 & ~x707 & ~x738 & ~x748;
assign c4234 =  x493 &  x521 &  x604 &  x632 &  x659 & ~x225;
assign c4236 =  x498 &  x655;
assign c4238 =  x492 &  x520 &  x576 &  x631 & ~x82 & ~x223 & ~x351 & ~x502 & ~x504 & ~x561 & ~x564 & ~x568 & ~x607 & ~x617 & ~x645 & ~x725 & ~x729;
assign c4240 =  x609 &  x773;
assign c4242 =  x124 &  x243 & ~x44 & ~x423;
assign c4244 =  x95 &  x123 &  x175 &  x631;
assign c4246 =  x205 &  x207 &  x208 &  x438 & ~x75;
assign c4248 =  x345 &  x597 & ~x572 & ~x577;
assign c4250 =  x182 &  x265 &  x292 & ~x31 & ~x202 & ~x246 & ~x406 & ~x433;
assign c4252 =  x55;
assign c4254 =  x318 & ~x59 & ~x70 & ~x271 & ~x280 & ~x328 & ~x330 & ~x335 & ~x359 & ~x614 & ~x670 & ~x741 & ~x764 & ~x770;
assign c4256 =  x27;
assign c4258 =  x365 & ~x184 & ~x210;
assign c4260 =  x654 &  x709 & ~x2 & ~x98 & ~x124 & ~x153 & ~x169 & ~x439;
assign c4262 =  x575 &  x603 &  x630 &  x631 &  x685 & ~x14 & ~x43 & ~x221 & ~x536;
assign c4264 =  x622 &  x656 & ~x715;
assign c4266 =  x602 &  x629 &  x656 & ~x16 & ~x52 & ~x70 & ~x100 & ~x108 & ~x427 & ~x454 & ~x531 & ~x614 & ~x616 & ~x667 & ~x668 & ~x760;
assign c4268 =  x39 &  x69;
assign c4270 =  x286 &  x441 & ~x372 & ~x425;
assign c4272 =  x119 &  x120 &  x653 &  x654 & ~x98;
assign c4274 =  x681 &  x708 &  x709 & ~x70 & ~x459 & ~x745;
assign c4276 =  x179 &  x437 &  x465 &  x521 &  x549 & ~x449;
assign c4278 =  x37 &  x178 & ~x197 & ~x772;
assign c4280 =  x450 & ~x549;
assign c4282 =  x337 &  x625;
assign c4284 =  x207 &  x235 &  x262 & ~x169 & ~x193 & ~x228 & ~x247 & ~x253 & ~x376 & ~x445 & ~x501 & ~x695 & ~x702 & ~x774;
assign c4286 =  x123 &  x151 &  x243 & ~x18 & ~x424 & ~x478 & ~x535;
assign c4288 =  x783;
assign c4290 =  x93 & ~x129 & ~x210 & ~x302 & ~x431 & ~x534;
assign c4292 = ~x113 & ~x141 & ~x247 & ~x276 & ~x308 & ~x320 & ~x321 & ~x393 & ~x418 & ~x501 & ~x589 & ~x615 & ~x619 & ~x645 & ~x651 & ~x702 & ~x725 & ~x730 & ~x774;
assign c4294 =  x622 &  x677 &  x709;
assign c4296 =  x133 &  x150 &  x371 &  x372 & ~x391;
assign c4298 =  x547 &  x575 &  x630 & ~x251 & ~x253 & ~x335 & ~x466 & ~x480 & ~x521 & ~x549 & ~x600 & ~x617 & ~x641 & ~x672 & ~x747 & ~x748;
assign c4300 =  x92 &  x93 &  x120 &  x545 & ~x14 & ~x617 & ~x721;
assign c4302 =  x182 &  x209 &  x236 &  x264 &  x291 &  x292 & ~x17 & ~x19 & ~x20 & ~x249 & ~x308 & ~x405 & ~x503 & ~x588 & ~x671 & ~x782;
assign c4304 =  x124 &  x382;
assign c4306 =  x610;
assign c4308 =  x126 & ~x59 & ~x230 & ~x266 & ~x417 & ~x457 & ~x765 & ~x774;
assign c4310 =  x292 &  x581 &  x654 & ~x274 & ~x311;
assign c4312 =  x606 &  x661 &  x689 & ~x25 & ~x44 & ~x75 & ~x197 & ~x335 & ~x446 & ~x582 & ~x703;
assign c4314 =  x125 &  x318 & ~x257 & ~x456 & ~x717;
assign c4316 =  x66 &  x94 &  x95 & ~x14 & ~x44;
assign c4318 =  x423;
assign c4320 =  x149 &  x332 &  x358;
assign c4322 =  x133 &  x626 &  x627;
assign c4324 =  x491 &  x546 & ~x130 & ~x159 & ~x171 & ~x230 & ~x272 & ~x303 & ~x454 & ~x480 & ~x648 & ~x673 & ~x699 & ~x772;
assign c4326 =  x522 &  x689 & ~x463;
assign c4328 =  x756;
assign c4330 =  x655 & ~x316;
assign c4332 =  x783;
assign c4334 =  x151 &  x179 &  x355 & ~x198 & ~x696 & ~x738;
assign c4336 = ~x15 & ~x30 & ~x44 & ~x55 & ~x70 & ~x72 & ~x195 & ~x210 & ~x214 & ~x236 & ~x237 & ~x330 & ~x410 & ~x438 & ~x548 & ~x660 & ~x716;
assign c4338 =  x574 & ~x185 & ~x281 & ~x293 & ~x305 & ~x387 & ~x432 & ~x472 & ~x571;
assign c4340 =  x493 &  x521 &  x632 &  x659 & ~x1 & ~x18 & ~x171 & ~x697;
assign c4342 =  x449 &  x651 & ~x13;
assign c4344 =  x462 & ~x42 & ~x87 & ~x270 & ~x273 & ~x331 & ~x410 & ~x480 & ~x606;
assign c4346 =  x574 &  x602 &  x629 &  x656 & ~x46 & ~x72 & ~x158 & ~x166 & ~x186 & ~x479 & ~x509 & ~x535 & ~x559 & ~x672 & ~x750 & ~x782;
assign c4348 =  x243 &  x467;
assign c4350 =  x175 &  x654 & ~x13 & ~x210 & ~x273 & ~x638;
assign c4352 =  x603 &  x631 &  x685 & ~x14 & ~x44 & ~x303;
assign c4354 =  x464 &  x492 &  x520 &  x603 &  x658 & ~x14 & ~x44 & ~x719 & ~x721;
assign c4356 =  x96 &  x179 &  x206 &  x207 & ~x321 & ~x725;
assign c4358 =  x247 &  x283;
assign c4360 =  x755;
assign c4362 =  x257 &  x467 & ~x75 & ~x102 & ~x371;
assign c4364 =  x206 &  x262 & ~x4 & ~x169 & ~x255 & ~x293 & ~x303 & ~x330 & ~x376 & ~x392;
assign c4366 =  x524 &  x552 &  x662 & ~x105 & ~x592;
assign c4368 =  x395 &  x709 & ~x70;
assign c4370 =  x471 &  x542 &  x570;
assign c4372 =  x357 &  x442 & ~x25 & ~x160 & ~x532 & ~x646 & ~x647;
assign c4374 =  x146 &  x147 &  x651;
assign c4376 =  x145 & ~x520 & ~x579;
assign c4378 =  x464 &  x575 &  x602 & ~x112 & ~x272 & ~x617 & ~x668 & ~x754 & ~x758;
assign c4380 =  x206 &  x208 &  x412 &  x440;
assign c4382 =  x523 &  x578 &  x605 &  x660 & ~x507;
assign c4384 =  x521 &  x549 &  x632 & ~x24 & ~x30 & ~x44 & ~x83 & ~x525 & ~x592 & ~x608 & ~x671 & ~x722;
assign c4386 =  x180 &  x207 &  x286 &  x467;
assign c4388 =  x421 & ~x137 & ~x266 & ~x439 & ~x689;
assign c4390 =  x413 & ~x345 & ~x425;
assign c4392 =  x553 & ~x450 & ~x703;
assign c4394 =  x69 &  x379 & ~x256 & ~x373 & ~x711;
assign c4396 =  x407 & ~x86 & ~x139 & ~x279 & ~x328 & ~x404 & ~x432 & ~x448 & ~x496 & ~x597 & ~x731;
assign c4398 =  x175 & ~x14 & ~x69 & ~x140 & ~x155 & ~x180 & ~x181 & ~x266 & ~x301 & ~x328 & ~x386 & ~x580;
assign c4400 =  x414 &  x550 & ~x373;
assign c4402 =  x182 &  x237 &  x522;
assign c4404 = ~x44 & ~x72 & ~x209 & ~x210 & ~x235 & ~x236 & ~x301 & ~x409 & ~x410 & ~x526 & ~x644 & ~x688;
assign c4406 =  x147 & ~x154 & ~x235 & ~x272 & ~x328 & ~x410 & ~x439 & ~x526;
assign c4408 =  x174 & ~x55 & ~x56 & ~x195 & ~x209 & ~x223 & ~x237 & ~x271 & ~x328 & ~x471 & ~x551 & ~x641 & ~x662 & ~x720 & ~x756;
assign c4410 = ~x0 & ~x155 & ~x196 & ~x222 & ~x225 & ~x252 & ~x266 & ~x293 & ~x321 & ~x415 & ~x469 & ~x473 & ~x524 & ~x528 & ~x532 & ~x608 & ~x614 & ~x637 & ~x652 & ~x707 & ~x750 & ~x759 & ~x765;
assign c4412 =  x492 &  x520 &  x576 &  x631 & ~x51 & ~x605 & ~x758;
assign c4414 =  x659 &  x687 & ~x240 & ~x249 & ~x367 & ~x445 & ~x516 & ~x532 & ~x568 & ~x624;
assign c4416 =  x256 &  x625 & ~x138 & ~x159;
assign c4418 =  x180 &  x467;
assign c4420 =  x151 &  x179 &  x270 & ~x293 & ~x374;
assign c4422 =  x208 &  x469 &  x497 & ~x245;
assign c4424 =  x94 &  x121 &  x545 & ~x210 & ~x308;
assign c4426 =  x602 &  x685 & ~x430 & ~x702;
assign c4428 =  x96 &  x150 & ~x197 & ~x237 & ~x346;
assign c4430 =  x699;
assign c4432 =  x180 &  x491 &  x519 &  x547 & ~x51 & ~x256 & ~x396 & ~x508 & ~x691;
assign c4434 =  x92 &  x471;
assign c4436 =  x68 &  x574 & ~x266;
assign c4438 =  x119 &  x707 &  x709 & ~x70;
assign c4440 =  x546 &  x600 & ~x29 & ~x57 & ~x166 & ~x193 & ~x221 & ~x359 & ~x612 & ~x614 & ~x689;
assign c4442 =  x781;
assign c4444 =  x655 &  x681 &  x682 &  x709 & ~x154 & ~x755;
assign c4446 =  x151 &  x410 &  x492;
assign c4448 =  x27;
assign c4450 =  x150 &  x179 & ~x2 & ~x155 & ~x388 & ~x625 & ~x680;
assign c4452 =  x92 &  x121 &  x653 &  x681;
assign c4454 =  x602 & ~x293 & ~x410 & ~x411 & ~x418 & ~x419 & ~x431 & ~x449 & ~x499;
assign c4456 =  x123 &  x262 & ~x218 & ~x293 & ~x305 & ~x719;
assign c4458 =  x265 &  x320 &  x492 & ~x433 & ~x619 & ~x673 & ~x675 & ~x697;
assign c4460 =  x683 &  x709 &  x737 & ~x246 & ~x247;
assign c4462 =  x526 &  x609 & ~x396;
assign c4464 =  x365 &  x597;
assign c4466 =  x653 &  x681 & ~x13 & ~x69 & ~x408 & ~x411 & ~x520 & ~x549 & ~x686;
assign c4468 =  x394 & ~x130 & ~x155 & ~x210 & ~x272;
assign c4470 = ~x129 & ~x155 & ~x210 & ~x237 & ~x238 & ~x273 & ~x303 & ~x430 & ~x501 & ~x612 & ~x652 & ~x702;
assign c4472 =  x96 &  x153 & ~x281 & ~x387 & ~x490;
assign c4474 =  x547 &  x574 & ~x86 & ~x115 & ~x183 & ~x226 & ~x247 & ~x256 & ~x285 & ~x313 & ~x388 & ~x445 & ~x505 & ~x533 & ~x673 & ~x698 & ~x725 & ~x764 & ~x773;
assign c4476 =  x680 & ~x436 & ~x692;
assign c4478 =  x123 &  x151 &  x179 &  x204 & ~x13 & ~x30 & ~x197 & ~x316 & ~x421 & ~x728 & ~x736;
assign c4480 =  x28;
assign c4482 =  x26;
assign c4484 =  x65 &  x94 &  x122 &  x576;
assign c4486 =  x783;
assign c4488 =  x496 &  x524 &  x579 &  x607 & ~x21 & ~x528;
assign c4490 = ~x50 & ~x70 & ~x169 & ~x207 & ~x300 & ~x308 & ~x329 & ~x330 & ~x389 & ~x499 & ~x548 & ~x715 & ~x774 & ~x783;
assign c4492 =  x463 & ~x217 & ~x424 & ~x454 & ~x689 & ~x711 & ~x778;
assign c4494 = ~x53 & ~x113 & ~x130 & ~x225 & ~x257 & ~x266 & ~x396 & ~x431 & ~x459 & ~x680 & ~x702 & ~x707;
assign c4496 =  x463 &  x491 &  x519 & ~x0 & ~x52 & ~x156 & ~x167 & ~x186 & ~x196 & ~x197 & ~x245 & ~x273 & ~x364 & ~x365 & ~x392 & ~x454 & ~x534 & ~x692 & ~x725 & ~x759 & ~x774;
assign c41 =  x45 & ~x529;
assign c43 =  x416 & ~x352;
assign c45 = ~x125 & ~x319 & ~x598 & ~x628 & ~x656;
assign c47 =  x417 & ~x32 & ~x37 & ~x64 & ~x66 & ~x722;
assign c49 =  x459 &  x460 &  x461 & ~x25 & ~x34 & ~x48 & ~x51 & ~x55 & ~x104 & ~x112 & ~x584 & ~x677 & ~x733 & ~x734 & ~x757 & ~x758 & ~x783;
assign c411 =  x266 &  x294 &  x351 & ~x36 & ~x83 & ~x440 & ~x447 & ~x585;
assign c413 = ~x96 & ~x114 & ~x320 & ~x582 & ~x598;
assign c415 =  x432 &  x461 & ~x34 & ~x494 & ~x532 & ~x553 & ~x590 & ~x594 & ~x617;
assign c417 =  x361 & ~x594 & ~x598;
assign c419 =  x381 &  x408 & ~x53 & ~x320 & ~x364 & ~x559 & ~x696 & ~x781;
assign c421 = ~x152 & ~x166 & ~x220 & ~x276 & ~x332 & ~x360 & ~x390 & ~x391 & ~x393 & ~x517 & ~x546 & ~x628 & ~x629 & ~x697;
assign c423 =  x487 &  x488 &  x516 & ~x77 & ~x104 & ~x194 & ~x224 & ~x413 & ~x440 & ~x615 & ~x643 & ~x762;
assign c425 =  x428 &  x456 &  x484 &  x488 & ~x53;
assign c427 = ~x1 & ~x18 & ~x67 & ~x74 & ~x77 & ~x85 & ~x96 & ~x295 & ~x615 & ~x640 & ~x676 & ~x693 & ~x694 & ~x707 & ~x737 & ~x745;
assign c429 =  x741 &  x742 & ~x688;
assign c431 =  x322 &  x350 &  x378 &  x714 & ~x106 & ~x139 & ~x191 & ~x481;
assign c433 =  x745 &  x746 & ~x364 & ~x550 & ~x609 & ~x644;
assign c435 =  x742 & ~x187 & ~x299 & ~x603;
assign c437 =  x456 &  x512 &  x620;
assign c439 =  x287 &  x342 &  x509;
assign c441 =  x566 &  x594 & ~x23 & ~x53 & ~x54 & ~x140 & ~x198 & ~x254 & ~x334 & ~x368 & ~x422 & ~x444;
assign c443 = ~x5 & ~x32 & ~x80 & ~x82 & ~x108 & ~x135 & ~x145 & ~x164 & ~x201 & ~x203 & ~x220 & ~x253 & ~x270 & ~x286 & ~x326 & ~x353 & ~x393 & ~x472 & ~x478 & ~x502 & ~x644;
assign c445 =  x287 &  x333 &  x343;
assign c447 =  x185 &  x211 &  x237 & ~x429 & ~x645;
assign c449 =  x405 & ~x77 & ~x82 & ~x309 & ~x340 & ~x368 & ~x424 & ~x445 & ~x453 & ~x471 & ~x496 & ~x504 & ~x522 & ~x553 & ~x557 & ~x565 & ~x583 & ~x756 & ~x763;
assign c451 =  x743 &  x745 & ~x106 & ~x134 & ~x161 & ~x191 & ~x219 & ~x280 & ~x528 & ~x585;
assign c453 =  x710 &  x740 &  x741 & ~x657 & ~x676;
assign c455 =  x741 &  x742 & ~x25 & ~x162 & ~x537 & ~x585 & ~x661;
assign c457 =  x98 &  x239 &  x267 &  x323;
assign c459 = ~x61 & ~x145 & ~x167 & ~x249 & ~x423 & ~x571 & ~x631 & ~x688;
assign c461 =  x259 &  x287 &  x288 &  x316 & ~x29 & ~x324 & ~x522 & ~x739 & ~x744 & ~x765;
assign c463 =  x232 &  x288 &  x333 &  x334 & ~x771;
assign c465 =  x745 & ~x108 & ~x134 & ~x139 & ~x188 & ~x196 & ~x222 & ~x244 & ~x333 & ~x420 & ~x529 & ~x555 & ~x610 & ~x648 & ~x704 & ~x782;
assign c467 =  x288 &  x342 &  x388;
assign c469 =  x75 & ~x398 & ~x484;
assign c471 =  x155 &  x156 &  x183 &  x184 & ~x484 & ~x487;
assign c473 =  x417 &  x446 & ~x14 & ~x32 & ~x55 & ~x142 & ~x358 & ~x722 & ~x723 & ~x763 & ~x766 & ~x778;
assign c475 = ~x289 & ~x336 & ~x544 & ~x601 & ~x627 & ~x742 & ~x743 & ~x770;
assign c477 =  x453 &  x481 &  x509 &  x566;
assign c479 =  x239 &  x267 &  x324 &  x352 &  x380 & ~x106 & ~x144 & ~x483;
assign c481 =  x715 & ~x53 & ~x107 & ~x108 & ~x270 & ~x565 & ~x577 & ~x580 & ~x701;
assign c483 =  x515 &  x516 &  x539 &  x540;
assign c485 =  x75 & ~x54 & ~x371 & ~x503;
assign c487 =  x713 & ~x0 & ~x52 & ~x56 & ~x105 & ~x308 & ~x527 & ~x586 & ~x603 & ~x608 & ~x633 & ~x728;
assign c489 =  x742 &  x743 &  x745 & ~x163;
assign c491 =  x741 & ~x26 & ~x30 & ~x32 & ~x159 & ~x603 & ~x605 & ~x606 & ~x613 & ~x631 & ~x696;
assign c493 =  x485 &  x486 &  x487 &  x515 &  x516;
assign c495 = ~x204 & ~x213 & ~x220 & ~x231 & ~x239 & ~x249 & ~x276 & ~x379 & ~x533 & ~x677;
assign c497 = ~x327 & ~x380 & ~x484 & ~x519 & ~x641 & ~x645 & ~x649 & ~x670;
assign c499 =  x484 &  x487 &  x488 &  x513;
assign c4101 =  x489 &  x517 & ~x4 & ~x106 & ~x242 & ~x283 & ~x296 & ~x471 & ~x525 & ~x527 & ~x558 & ~x644;
assign c4103 =  x324 &  x349 &  x352 & ~x364 & ~x442;
assign c4105 =  x473 &  x500 & ~x68;
assign c4107 =  x305 & ~x594 & ~x721 & ~x744 & ~x771;
assign c4109 =  x455 &  x537 & ~x75 & ~x769;
assign c4111 =  x316 &  x456 &  x457 &  x458;
assign c4113 = ~x33 & ~x49 & ~x74 & ~x87 & ~x106 & ~x109 & ~x130 & ~x134 & ~x160 & ~x185 & ~x212 & ~x214 & ~x245 & ~x246 & ~x272 & ~x286 & ~x296 & ~x324 & ~x365 & ~x368 & ~x394 & ~x526 & ~x579 & ~x584 & ~x585 & ~x609 & ~x612 & ~x617 & ~x669 & ~x723 & ~x783;
assign c4115 =  x459 &  x460 &  x461 & ~x29 & ~x368 & ~x394 & ~x526;
assign c4117 =  x101 & ~x25 & ~x33 & ~x224 & ~x280 & ~x336 & ~x372 & ~x400 & ~x484 & ~x558 & ~x586 & ~x615;
assign c4119 = ~x46 & ~x77 & ~x189 & ~x200 & ~x211 & ~x243 & ~x328 & ~x380 & ~x408 & ~x728;
assign c4121 =  x327 & ~x41 & ~x100 & ~x125 & ~x179;
assign c4123 =  x269 &  x324 & ~x258 & ~x286;
assign c4125 =  x258 & ~x39 & ~x40 & ~x66 & ~x67 & ~x94 & ~x340 & ~x366 & ~x421 & ~x769;
assign c4127 = ~x26 & ~x174 & ~x203 & ~x204 & ~x380 & ~x407 & ~x708;
assign c4129 =  x451 & ~x2 & ~x26 & ~x52 & ~x652 & ~x707;
assign c4131 =  x731 & ~x95;
assign c4133 = ~x179 & ~x288 & ~x289 & ~x420 & ~x517 & ~x629;
assign c4135 =  x740 &  x741 &  x742 & ~x662;
assign c4137 = ~x40 & ~x67 & ~x484 & ~x571 & ~x598 & ~x628;
assign c4139 =  x184 &  x352 & ~x485;
assign c4141 =  x746 &  x747 & ~x579;
assign c4143 = ~x119 & ~x139 & ~x145 & ~x201 & ~x203 & ~x313 & ~x314 & ~x422 & ~x601 & ~x603;
assign c4145 =  x306 & ~x242 & ~x243;
assign c4147 =  x115;
assign c4149 =  x277 & ~x243 & ~x244 & ~x245 & ~x593;
assign c4151 =  x636 & ~x59 & ~x421 & ~x741 & ~x749 & ~x754 & ~x772 & ~x774;
assign c4153 =  x742 &  x744;
assign c4155 =  x259 &  x509 &  x510;
assign c4157 =  x342 &  x370 &  x455 &  x483 &  x484 & ~x615;
assign c4159 =  x432 & ~x52 & ~x211 & ~x340 & ~x418 & ~x536 & ~x552 & ~x648 & ~x765;
assign c4161 =  x274 & ~x38 & ~x65 & ~x106;
assign c4163 =  x269 &  x296 &  x297 &  x323 &  x324 &  x352 & ~x22 & ~x27 & ~x53 & ~x360 & ~x361 & ~x387;
assign c4165 =  x326 &  x352 &  x353 & ~x80 & ~x341 & ~x419 & ~x470 & ~x591 & ~x724;
assign c4167 =  x432 &  x461 & ~x54 & ~x395 & ~x397 & ~x414 & ~x443 & ~x498 & ~x505 & ~x639 & ~x754 & ~x759 & ~x779;
assign c4169 =  x342 &  x370 &  x483 &  x509 &  x510;
assign c4171 =  x160 &  x184 &  x185;
assign c4173 = ~x61 & ~x62 & ~x400 & ~x487 & ~x489 & ~x544 & ~x547;
assign c4175 =  x566 & ~x201 & ~x360 & ~x422;
assign c4177 =  x428 &  x456 &  x457 &  x459 & ~x19 & ~x107;
assign c4179 =  x537 &  x667;
assign c4181 = ~x26 & ~x109 & ~x110 & ~x203 & ~x285 & ~x671 & ~x687 & ~x716;
assign c4183 =  x274 & ~x38 & ~x64 & ~x66;
assign c4185 =  x743 &  x744 &  x745 & ~x196 & ~x219 & ~x305 & ~x530 & ~x604;
assign c4187 =  x287 & ~x64 & ~x108 & ~x323 & ~x379 & ~x493;
assign c4189 =  x214 & ~x204 & ~x233;
assign c4191 =  x457 &  x486 & ~x6 & ~x40 & ~x57 & ~x134 & ~x136 & ~x166 & ~x615 & ~x756 & ~x774;
assign c4193 =  x744 &  x745 & ~x18 & ~x45 & ~x54 & ~x55 & ~x77 & ~x133 & ~x136 & ~x167 & ~x191 & ~x195 & ~x199 & ~x200 & ~x311 & ~x364 & ~x479 & ~x558 & ~x586 & ~x669 & ~x728 & ~x729 & ~x759;
assign c4195 =  x183 &  x211 &  x239 & ~x19 & ~x481 & ~x484 & ~x583 & ~x609 & ~x759;
assign c4197 =  x296 & ~x66 & ~x93 & ~x122 & ~x305;
assign c4199 =  x239 &  x592;
assign c4201 =  x287 &  x333 &  x343;
assign c4203 =  x352 &  x376 &  x379 & ~x340 & ~x499 & ~x673;
assign c4205 =  x185 &  x213 &  x240 &  x241 &  x242;
assign c4207 =  x397 &  x453 &  x481 &  x509 &  x537;
assign c4209 =  x185 &  x212 &  x213 &  x240 &  x242;
assign c4211 =  x306;
assign c4213 =  x156 &  x324 & ~x456;
assign c4215 =  x742 &  x745 & ~x136 & ~x248;
assign c4217 =  x211 &  x239 &  x267 &  x352 & ~x5;
assign c4219 =  x485 &  x486 &  x515 & ~x355 & ~x763 & ~x777;
assign c4221 =  x348 &  x350 &  x376 & ~x338 & ~x414 & ~x559;
assign c4223 =  x333 & ~x563;
assign c4225 = ~x175 & ~x258 & ~x285 & ~x314 & ~x575 & ~x605;
assign c4227 =  x483 &  x538 &  x539 & ~x112 & ~x192 & ~x615 & ~x746 & ~x769;
assign c4229 =  x483 &  x484 &  x509 &  x536 & ~x30 & ~x42;
assign c4231 =  x12 & ~x2 & ~x23 & ~x27 & ~x58 & ~x81 & ~x170 & ~x224 & ~x251 & ~x277 & ~x281 & ~x333 & ~x388 & ~x444 & ~x472 & ~x476 & ~x530 & ~x533 & ~x584 & ~x586 & ~x587 & ~x589 & ~x591 & ~x616 & ~x619 & ~x638 & ~x643 & ~x644 & ~x698 & ~x759 & ~x782;
assign c4233 =  x376 &  x405 & ~x24 & ~x54 & ~x312 & ~x397 & ~x439 & ~x443 & ~x535 & ~x617 & ~x706 & ~x734 & ~x752;
assign c4235 =  x211 &  x239 &  x267 &  x295 & ~x399;
assign c4237 =  x156 &  x296 &  x324 & ~x537;
assign c4239 = ~x96 & ~x370 & ~x419 & ~x457 & ~x483 & ~x541 & ~x544 & ~x643;
assign c4241 = ~x51 & ~x58 & ~x134 & ~x164 & ~x211 & ~x243 & ~x273 & ~x553 & ~x589 & ~x607 & ~x695 & ~x732;
assign c4243 =  x269 &  x295 &  x296 &  x352 &  x380 & ~x644;
assign c4245 =  x131 & ~x540 & ~x627;
assign c4247 = ~x3 & ~x22 & ~x29 & ~x59 & ~x77 & ~x241 & ~x244 & ~x442 & ~x446 & ~x448 & ~x477 & ~x497 & ~x502 & ~x553 & ~x580 & ~x605 & ~x606 & ~x609 & ~x639 & ~x668 & ~x670 & ~x672 & ~x760;
assign c4249 =  x333 & ~x139 & ~x598 & ~x622 & ~x650 & ~x677 & ~x759;
assign c4251 = ~x111 & ~x151 & ~x152 & ~x179 & ~x447 & ~x477 & ~x598 & ~x658 & ~x659;
assign c4253 =  x459 &  x460 &  x461 & ~x24 & ~x57 & ~x336 & ~x609 & ~x766;
assign c4255 =  x540 & ~x137 & ~x220 & ~x253 & ~x259 & ~x314;
assign c4257 =  x263 &  x489 & ~x4 & ~x80 & ~x86 & ~x163 & ~x296 & ~x352 & ~x695 & ~x701 & ~x733 & ~x762;
assign c4259 = ~x203 & ~x289 & ~x314 & ~x319 & ~x347;
assign c4261 =  x202 &  x341 &  x369;
assign c4263 = ~x22 & ~x99 & ~x112 & ~x168 & ~x200 & ~x349 & ~x475 & ~x485 & ~x598 & ~x644 & ~x712 & ~x714;
assign c4265 = ~x257 & ~x287 & ~x408 & ~x602 & ~x603;
assign c4267 = ~x38 & ~x66 & ~x377 & ~x380 & ~x408 & ~x504 & ~x611 & ~x644 & ~x695 & ~x771 & ~x772;
assign c4269 =  x417 & ~x38 & ~x380;
assign c4271 =  x316 &  x372 &  x373 &  x401 &  x430 &  x601;
assign c4273 =  x516 &  x743 &  x744 & ~x106;
assign c4275 =  x740 &  x741 &  x742 & ~x365 & ~x636 & ~x660 & ~x755;
assign c4277 = ~x93 & ~x121 & ~x203 & ~x687 & ~x741 & ~x744;
assign c4279 =  x674 & ~x391;
assign c4281 =  x323 &  x351 & ~x7 & ~x33 & ~x251 & ~x259 & ~x279 & ~x280 & ~x285 & ~x390 & ~x442 & ~x453 & ~x480 & ~x506 & ~x507 & ~x640 & ~x673 & ~x762;
assign c4283 = ~x55 & ~x67 & ~x96 & ~x371 & ~x421 & ~x455 & ~x628 & ~x677 & ~x709 & ~x778 & ~x780;
assign c4285 =  x287 & ~x19 & ~x37 & ~x320 & ~x598 & ~x744;
assign c4287 = ~x206 & ~x233 & ~x288 & ~x315 & ~x490 & ~x517 & ~x644;
assign c4289 =  x401 &  x429 &  x460 & ~x34 & ~x191 & ~x308 & ~x777;
assign c4291 =  x457 &  x486 & ~x134 & ~x138 & ~x140 & ~x162 & ~x191 & ~x215 & ~x758 & ~x759;
assign c4293 =  x741 &  x770 & ~x52 & ~x107 & ~x108 & ~x163 & ~x558 & ~x698;
assign c4295 =  x71 &  x99 &  x351;
assign c4297 =  x488 &  x489 &  x518 & ~x21 & ~x51 & ~x64 & ~x85 & ~x89 & ~x721 & ~x734;
assign c4299 =  x324 &  x352 &  x353 &  x381 & ~x259 & ~x585 & ~x587 & ~x615;
assign c4301 = ~x13 & ~x40 & ~x66 & ~x67 & ~x68 & ~x154 & ~x211 & ~x294 & ~x347 & ~x734 & ~x765;
assign c4303 =  x485 &  x486 &  x487 &  x488 &  x516 & ~x757 & ~x761;
assign c4305 =  x693 &  x694 & ~x366 & ~x421 & ~x530 & ~x776;
assign c4307 =  x452 & ~x62 & ~x73 & ~x90 & ~x310;
assign c4309 =  x326 & ~x27 & ~x67 & ~x93 & ~x122 & ~x150;
assign c4311 =  x460 &  x461 & ~x146 & ~x161 & ~x560 & ~x649 & ~x673 & ~x754;
assign c4313 =  x456 &  x480 &  x481;
assign c4315 = ~x96 & ~x178 & ~x206 & ~x489 & ~x544 & ~x726;
assign c4317 = ~x6 & ~x26 & ~x50 & ~x62 & ~x82 & ~x87 & ~x137 & ~x167 & ~x241 & ~x250 & ~x276 & ~x309 & ~x362 & ~x394 & ~x395 & ~x415 & ~x444 & ~x448 & ~x449 & ~x521 & ~x522 & ~x525 & ~x553 & ~x579 & ~x590 & ~x722 & ~x733 & ~x754 & ~x760;
assign c4319 =  x131 & ~x121 & ~x371;
assign c4321 = ~x28 & ~x58 & ~x82 & ~x89 & ~x188 & ~x212 & ~x308 & ~x310 & ~x313 & ~x363 & ~x366 & ~x393 & ~x453 & ~x475 & ~x479 & ~x495 & ~x499 & ~x565 & ~x567 & ~x580 & ~x593 & ~x594 & ~x609 & ~x615 & ~x623 & ~x673 & ~x732 & ~x733;
assign c4323 =  x696;
assign c4325 =  x102 &  x103 & ~x400;
assign c4327 =  x376 &  x406 & ~x77 & ~x285 & ~x395 & ~x423 & ~x472 & ~x502 & ~x524 & ~x526 & ~x564;
assign c4329 =  x323 &  x324 &  x348 &  x351 & ~x587 & ~x695;
assign c4331 =  x266 &  x294 & ~x52 & ~x63 & ~x113 & ~x201 & ~x282 & ~x557 & ~x639 & ~x729 & ~x752;
assign c4333 =  x389 &  x417 & ~x650 & ~x722;
assign c4335 =  x288 &  x418;
assign c4337 =  x480 &  x507 &  x508 &  x535 & ~x394;
assign c4339 =  x277 & ~x539 & ~x560 & ~x593 & ~x650 & ~x774;
assign c4341 =  x510 &  x511 &  x512 &  x539 & ~x134 & ~x324;
assign c4343 =  x221 & ~x565 & ~x591 & ~x617;
assign c4345 = ~x178 & ~x233 & ~x288 & ~x572;
assign c4347 = ~x62 & ~x220 & ~x365 & ~x408 & ~x571 & ~x655 & ~x656;
assign c4349 =  x323 &  x350 &  x351 & ~x121 & ~x285;
assign c4351 = ~x176 & ~x211 & ~x232 & ~x287 & ~x519;
assign c4353 =  x194;
assign c4355 = ~x127 & ~x306 & ~x391 & ~x598 & ~x628 & ~x629 & ~x712 & ~x756;
assign c4357 =  x466 & ~x1 & ~x215 & ~x269 & ~x553 & ~x662;
assign c4359 =  x98 &  x267 &  x323 &  x351;
assign c4361 =  x13 & ~x85 & ~x109 & ~x253 & ~x504 & ~x574 & ~x730;
assign c4363 =  x535 &  x562 & ~x280 & ~x708 & ~x772;
assign c4365 =  x705 & ~x710;
assign c4367 =  x104 & ~x26 & ~x52 & ~x481 & ~x503 & ~x616;
assign c4369 = ~x181 & ~x234 & ~x598 & ~x627 & ~x628 & ~x629 & ~x653 & ~x656 & ~x671 & ~x683 & ~x777 & ~x782;
assign c4371 =  x156 &  x184 &  x212 & ~x312 & ~x428 & ~x585;
assign c4373 =  x296 &  x323 &  x324 &  x348 & ~x31 & ~x79;
assign c4375 =  x298 &  x324 &  x326 &  x353 & ~x60 & ~x305 & ~x336 & ~x340 & ~x443 & ~x474;
assign c4377 =  x333 & ~x110 & ~x245 & ~x592 & ~x649 & ~x719 & ~x720 & ~x747 & ~x749 & ~x773 & ~x776 & ~x780;
assign c4379 =  x240 &  x266 &  x267 &  x268 & ~x328;
assign c4381 = ~x107 & ~x114 & ~x118 & ~x145 & ~x168 & ~x174 & ~x189 & ~x203 & ~x211 & ~x239 & ~x276 & ~x324 & ~x365 & ~x420 & ~x443 & ~x450 & ~x472 & ~x523 & ~x706 & ~x734;
assign c4383 =  x157 &  x184 & ~x430 & ~x627;
assign c4385 =  x242 &  x267 &  x269 & ~x356;
assign c4387 =  x342 &  x425 &  x426 & ~x31 & ~x49 & ~x51 & ~x83 & ~x106 & ~x113 & ~x138 & ~x394 & ~x724 & ~x736 & ~x756;
assign c4389 =  x267 &  x269 &  x294 &  x297;
assign c4391 =  x380 &  x381 & ~x4 & ~x7 & ~x33 & ~x50 & ~x78 & ~x81 & ~x164 & ~x191 & ~x416 & ~x441 & ~x498 & ~x528 & ~x609;
assign c4393 =  x343 &  x484 &  x540 &  x568;
assign c4395 =  x718 & ~x21 & ~x30 & ~x33 & ~x61 & ~x78 & ~x81 & ~x82 & ~x163 & ~x500 & ~x552 & ~x559 & ~x584 & ~x609;
assign c4397 = ~x67 & ~x94 & ~x122 & ~x294 & ~x320 & ~x640 & ~x641 & ~x677 & ~x706 & ~x729 & ~x747;
assign c4399 =  x268 &  x296 & ~x67 & ~x251 & ~x314;
assign c4401 =  x428 &  x456 &  x483 &  x510 &  x536 & ~x393;
assign c4403 = ~x67 & ~x93 & ~x94 & ~x96 & ~x121 & ~x122 & ~x140 & ~x150 & ~x172;
assign c4405 = ~x33 & ~x289 & ~x400 & ~x408 & ~x575 & ~x601;
assign c4407 =  x445 & ~x78 & ~x380 & ~x408 & ~x641 & ~x644;
assign c4409 =  x183 &  x212 & ~x61 & ~x81 & ~x88 & ~x416 & ~x427 & ~x484 & ~x555 & ~x645;
assign c4411 =  x454 &  x480 &  x481 & ~x768;
assign c4413 =  x156 &  x296 &  x324 & ~x483 & ~x640;
assign c4415 =  x327 & ~x267 & ~x413 & ~x772;
assign c4417 =  x232 & ~x64 & ~x172 & ~x211 & ~x504;
assign c4419 =  x278 & ~x594 & ~x624;
assign c4421 = ~x38 & ~x40 & ~x90 & ~x484 & ~x541 & ~x598 & ~x627 & ~x741;
assign c4423 =  x248 & ~x536 & ~x537 & ~x538 & ~x565 & ~x619;
assign c4425 =  x327 & ~x1 & ~x96 & ~x152 & ~x367;
assign c4427 = ~x15 & ~x130 & ~x162 & ~x189 & ~x211 & ~x268 & ~x351 & ~x352 & ~x394 & ~x471 & ~x529;
assign c4429 =  x277 & ~x566 & ~x593;
assign c4431 = ~x53 & ~x66 & ~x67 & ~x175 & ~x282 & ~x687 & ~x741;
assign c4433 =  x193 & ~x587 & ~x616 & ~x716 & ~x768;
assign c4435 =  x713 & ~x392 & ~x501 & ~x609 & ~x615 & ~x659 & ~x665 & ~x755;
assign c4437 =  x405 & ~x4 & ~x6 & ~x22 & ~x26 & ~x31 & ~x61 & ~x84 & ~x89 & ~x114 & ~x342 & ~x366 & ~x368 & ~x370 & ~x387 & ~x412 & ~x416 & ~x426 & ~x470 & ~x478 & ~x525 & ~x529 & ~x532 & ~x565 & ~x594 & ~x622 & ~x642 & ~x670 & ~x672 & ~x676 & ~x700 & ~x730 & ~x778;
assign c4439 = ~x32 & ~x33 & ~x142 & ~x195 & ~x281 & ~x334 & ~x368 & ~x371 & ~x389 & ~x391 & ~x393 & ~x425 & ~x430 & ~x447 & ~x454 & ~x488 & ~x564 & ~x722 & ~x759 & ~x780;
assign c4441 = ~x282 & ~x289 & ~x489 & ~x603 & ~x628;
assign c4443 = ~x178 & ~x206 & ~x233 & ~x288 & ~x573 & ~x575;
assign c4445 =  x296 & ~x286 & ~x314 & ~x429;
assign c4447 =  x294 &  x321 &  x350 & ~x61 & ~x64 & ~x91 & ~x643 & ~x756;
assign c4449 =  x323 & ~x52 & ~x258 & ~x288 & ~x303 & ~x362 & ~x396 & ~x400 & ~x414 & ~x458 & ~x617 & ~x703 & ~x705 & ~x758;
assign c4451 =  x267 &  x323 & ~x62 & ~x106 & ~x141 & ~x145 & ~x170 & ~x171 & ~x398 & ~x456 & ~x535 & ~x614 & ~x755 & ~x783;
assign c4453 =  x431 &  x460 &  x461 & ~x8 & ~x51 & ~x223 & ~x365 & ~x366 & ~x615 & ~x645 & ~x674 & ~x677 & ~x702 & ~x736 & ~x780;
assign c4455 =  x220 & ~x188 & ~x456;
assign c4457 = ~x6 & ~x29 & ~x55 & ~x90 & ~x172 & ~x174 & ~x285 & ~x314 & ~x395 & ~x519 & ~x658 & ~x671 & ~x687;
assign c4459 =  x620 &  x675 & ~x197;
assign c4461 =  x741 &  x742 & ~x5 & ~x51 & ~x56 & ~x336 & ~x586 & ~x609 & ~x631 & ~x701 & ~x754;
assign c4463 =  x741 &  x742 & ~x27 & ~x32 & ~x80 & ~x164 & ~x364 & ~x426 & ~x453 & ~x480 & ~x529 & ~x562 & ~x564 & ~x584 & ~x611 & ~x642;
assign c4465 =  x385 &  x539 & ~x26 & ~x57 & ~x61 & ~x199 & ~x254 & ~x255 & ~x449 & ~x504;
assign c4467 = ~x61 & ~x233 & ~x254 & ~x443 & ~x472 & ~x487 & ~x489 & ~x531 & ~x644;
assign c4469 =  x518 & ~x107 & ~x137 & ~x252 & ~x399 & ~x400 & ~x429 & ~x442 & ~x468 & ~x486 & ~x527;
assign c4471 = ~x60 & ~x200 & ~x290 & ~x408 & ~x477 & ~x517 & ~x544 & ~x629;
assign c4473 =  x212 &  x240 &  x268 & ~x287;
assign c4475 =  x416 & ~x49 & ~x84 & ~x678 & ~x681;
assign c4477 =  x45 & ~x588;
assign c4479 = ~x6 & ~x88 & ~x298 & ~x510 & ~x598 & ~x616 & ~x627 & ~x666 & ~x667 & ~x727 & ~x729;
assign c4481 =  x460 &  x482 &  x510;
assign c4483 = ~x59 & ~x61 & ~x110 & ~x400 & ~x629 & ~x631 & ~x642 & ~x727 & ~x757 & ~x773;
assign c4485 =  x44 &  x45;
assign c4487 =  x741 & ~x83 & ~x139 & ~x269 & ~x530 & ~x583 & ~x603 & ~x644;
assign c4489 =  x620 & ~x233 & ~x288;
assign c4491 =  x232 &  x277 & ~x243;
assign c4493 =  x479 &  x507 &  x535 & ~x113 & ~x771;
assign c4495 =  x427 &  x483 &  x511 &  x539 & ~x79 & ~x424;
assign c4497 =  x544 &  x742 &  x743 &  x744 & ~x106 & ~x135;
assign c4499 =  x314 & ~x38 & ~x296 & ~x347 & ~x376 & ~x379 & ~x726;
assign c50 =  x485 &  x512 &  x513 &  x540 &  x541 & ~x0 & ~x76 & ~x104 & ~x114 & ~x253 & ~x256 & ~x339 & ~x351 & ~x379 & ~x383 & ~x385 & ~x396;
assign c52 =  x239 &  x295 &  x601;
assign c54 =  x385 &  x443 &  x500;
assign c56 =  x423 & ~x38 & ~x269 & ~x323 & ~x345 & ~x566 & ~x593;
assign c58 =  x688 &  x689 & ~x31 & ~x77 & ~x201 & ~x247 & ~x250 & ~x276 & ~x340 & ~x379 & ~x410 & ~x464 & ~x470 & ~x492 & ~x500 & ~x501 & ~x556 & ~x701;
assign c510 =  x245 &  x304 & ~x235 & ~x688;
assign c512 =  x237 &  x348 &  x376 & ~x79 & ~x104 & ~x218 & ~x246 & ~x301 & ~x330 & ~x331 & ~x340 & ~x369 & ~x371 & ~x398 & ~x527 & ~x595 & ~x596 & ~x625 & ~x675 & ~x710 & ~x765 & ~x780;
assign c514 =  x361 &  x451 & ~x110 & ~x265 & ~x270 & ~x511 & ~x710;
assign c516 =  x375 & ~x3 & ~x5 & ~x7 & ~x18 & ~x32 & ~x48 & ~x61 & ~x92 & ~x108 & ~x115 & ~x119 & ~x134 & ~x137 & ~x146 & ~x162 & ~x166 & ~x173 & ~x174 & ~x188 & ~x196 & ~x198 & ~x200 & ~x217 & ~x219 & ~x225 & ~x230 & ~x254 & ~x255 & ~x271 & ~x275 & ~x277 & ~x286 & ~x303 & ~x311 & ~x313 & ~x314 & ~x327 & ~x331 & ~x333 & ~x340 & ~x363 & ~x369 & ~x370 & ~x384 & ~x386 & ~x389 & ~x397 & ~x412 & ~x413 & ~x419 & ~x421 & ~x424 & ~x453 & ~x473 & ~x505 & ~x506 & ~x527 & ~x536 & ~x557 & ~x567 & ~x584 & ~x594 & ~x596 & ~x598 & ~x614 & ~x619 & ~x624 & ~x638 & ~x641 & ~x644 & ~x652 & ~x667 & ~x673 & ~x674 & ~x675 & ~x676 & ~x708 & ~x723 & ~x729 & ~x731 & ~x732 & ~x782;
assign c518 = ~x123 & ~x150 & ~x209 & ~x347 & ~x349 & ~x409 & ~x487 & ~x566 & ~x593;
assign c520 =  x486 &  x541 &  x685 &  x713 &  x743 & ~x93 & ~x272 & ~x303 & ~x314 & ~x333 & ~x354 & ~x370 & ~x385 & ~x733;
assign c522 =  x397 &  x398 &  x453 & ~x321 & ~x347 & ~x459;
assign c524 =  x385 &  x412 & ~x209 & ~x215;
assign c526 =  x321 &  x460 &  x513 &  x541 &  x714 &  x773 & ~x151 & ~x380;
assign c528 =  x453;
assign c530 =  x659 &  x687 & ~x86 & ~x113 & ~x217 & ~x222 & ~x226 & ~x230 & ~x243 & ~x258 & ~x274 & ~x296 & ~x298 & ~x308 & ~x311 & ~x329 & ~x330 & ~x354 & ~x368 & ~x382 & ~x383 & ~x413 & ~x445 & ~x478 & ~x479 & ~x531 & ~x533 & ~x534 & ~x555 & ~x556 & ~x588 & ~x590 & ~x627 & ~x667 & ~x668 & ~x699 & ~x704 & ~x730 & ~x760;
assign c532 =  x523 &  x579 & ~x150 & ~x246 & ~x305 & ~x586 & ~x709;
assign c534 =  x223 &  x421;
assign c536 =  x453 &  x482 & ~x228 & ~x347 & ~x458;
assign c538 =  x301 &  x387 & ~x154 & ~x744;
assign c540 =  x209 &  x348 &  x576 & ~x413 & ~x451;
assign c542 =  x155 &  x157 & ~x252 & ~x335 & ~x357 & ~x382 & ~x385 & ~x413 & ~x443 & ~x526 & ~x528 & ~x585 & ~x700 & ~x755 & ~x762;
assign c544 =  x426 &  x456 &  x510 & ~x436;
assign c546 =  x689 & ~x1 & ~x8 & ~x22 & ~x26 & ~x28 & ~x46 & ~x50 & ~x54 & ~x55 & ~x77 & ~x79 & ~x81 & ~x83 & ~x84 & ~x110 & ~x137 & ~x141 & ~x164 & ~x190 & ~x194 & ~x195 & ~x220 & ~x247 & ~x255 & ~x256 & ~x274 & ~x282 & ~x284 & ~x307 & ~x308 & ~x312 & ~x330 & ~x332 & ~x337 & ~x339 & ~x340 & ~x352 & ~x360 & ~x361 & ~x365 & ~x386 & ~x391 & ~x393 & ~x394 & ~x406 & ~x422 & ~x423 & ~x435 & ~x446 & ~x474 & ~x475 & ~x506 & ~x531 & ~x560 & ~x590 & ~x614 & ~x615 & ~x643 & ~x698 & ~x727 & ~x757 & ~x782 & ~x783;
assign c548 =  x454 &  x472 &  x536 & ~x235;
assign c550 =  x292 &  x293 &  x350 &  x459 & ~x151 & ~x201 & ~x451 & ~x735 & ~x737;
assign c552 =  x426 &  x509 & ~x125 & ~x348 & ~x358 & ~x430;
assign c554 =  x423 & ~x179 & ~x203 & ~x242 & ~x299 & ~x541 & ~x556;
assign c556 =  x746 &  x747 & ~x5 & ~x75 & ~x162 & ~x220 & ~x331 & ~x340 & ~x342 & ~x383 & ~x413 & ~x435 & ~x468 & ~x494 & ~x522;
assign c558 =  x373 &  x402 &  x456 & ~x465 & ~x466 & ~x768;
assign c560 =  x315 &  x371 &  x398 &  x426 & ~x149 & ~x742;
assign c562 =  x355 &  x413 & ~x212;
assign c564 =  x188 &  x199 &  x503;
assign c566 = ~x123 & ~x293 & ~x295 & ~x319 & ~x347 & ~x349 & ~x373 & ~x377 & ~x379 & ~x392 & ~x430 & ~x445 & ~x473 & ~x486 & ~x559 & ~x643 & ~x712;
assign c568 =  x358 & ~x605;
assign c570 = ~x6 & ~x75 & ~x78 & ~x84 & ~x117 & ~x169 & ~x172 & ~x225 & ~x226 & ~x229 & ~x283 & ~x294 & ~x323 & ~x325 & ~x326 & ~x355 & ~x358 & ~x382 & ~x383 & ~x387 & ~x406 & ~x413 & ~x421 & ~x435 & ~x443 & ~x497 & ~x583 & ~x669 & ~x708 & ~x735 & ~x737 & ~x761 & ~x765;
assign c572 =  x240 &  x543 &  x571 &  x599 & ~x385 & ~x414 & ~x435 & ~x438 & ~x527;
assign c574 = ~x39 & ~x69 & ~x110 & ~x211 & ~x265 & ~x378 & ~x430 & ~x596 & ~x739;
assign c576 =  x340 & ~x213 & ~x236 & ~x317;
assign c578 =  x524 &  x578 & ~x294 & ~x417;
assign c580 =  x662 &  x705;
assign c582 =  x236 &  x264 &  x458 &  x512 &  x684 & ~x370;
assign c584 =  x265 &  x602 &  x742 &  x772;
assign c586 =  x403 &  x487 &  x629 &  x743 &  x744 &  x745;
assign c588 =  x340 & ~x184 & ~x211 & ~x241 & ~x265;
assign c590 =  x659 &  x687 & ~x90 & ~x114 & ~x143 & ~x164 & ~x199 & ~x201 & ~x219 & ~x243 & ~x247 & ~x252 & ~x285 & ~x286 & ~x303 & ~x330 & ~x331 & ~x364 & ~x366 & ~x367 & ~x369 & ~x386 & ~x414 & ~x444 & ~x473 & ~x527 & ~x627 & ~x648 & ~x656 & ~x683;
assign c592 =  x397 & ~x347 & ~x374 & ~x537;
assign c594 =  x346 &  x373 &  x374 &  x401 & ~x183 & ~x188 & ~x211 & ~x216 & ~x286 & ~x314 & ~x365 & ~x702;
assign c596 =  x383 &  x469 &  x471;
assign c598 =  x331 & ~x541;
assign c5100 =  x635 &  x662 & ~x166 & ~x331 & ~x334 & ~x391 & ~x409 & ~x470 & ~x473 & ~x684;
assign c5102 =  x661 &  x693 & ~x302 & ~x443;
assign c5104 =  x355 &  x413 &  x414 &  x471;
assign c5106 =  x413 &  x469;
assign c5108 =  x660;
assign c5110 =  x266 &  x321 &  x433 & ~x67 & ~x144 & ~x286 & ~x380 & ~x425 & ~x454 & ~x681;
assign c5112 =  x419;
assign c5114 =  x552 & ~x375 & ~x409 & ~x499;
assign c5116 =  x236 &  x375 & ~x184 & ~x215 & ~x228 & ~x300 & ~x330 & ~x342 & ~x359 & ~x538 & ~x562 & ~x665 & ~x695;
assign c5118 =  x72 &  x100 & ~x229 & ~x247 & ~x251 & ~x274 & ~x300 & ~x301 & ~x313 & ~x333 & ~x355 & ~x410 & ~x468 & ~x494 & ~x497 & ~x528 & ~x556;
assign c5120 =  x420;
assign c5122 =  x452 & ~x347 & ~x373 & ~x485 & ~x514 & ~x622;
assign c5124 = ~x125 & ~x203 & ~x375 & ~x621;
assign c5126 =  x457 &  x512 &  x539 &  x541 &  x568 & ~x22 & ~x576;
assign c5128 =  x576 & ~x183 & ~x184 & ~x185 & ~x219 & ~x240 & ~x241 & ~x284 & ~x300 & ~x342 & ~x388 & ~x424 & ~x588;
assign c5130 =  x375 &  x403 &  x457 &  x484 & ~x498 & ~x523 & ~x524 & ~x548 & ~x606 & ~x695 & ~x726;
assign c5132 =  x293 &  x404 &  x433 &  x486 &  x687 &  x773 & ~x397;
assign c5134 =  x348 &  x375 & ~x63 & ~x113 & ~x159 & ~x162 & ~x163 & ~x170 & ~x173 & ~x218 & ~x219 & ~x222 & ~x246 & ~x251 & ~x278 & ~x283 & ~x296 & ~x299 & ~x300 & ~x301 & ~x305 & ~x314 & ~x316 & ~x365 & ~x395 & ~x396 & ~x414 & ~x425 & ~x473 & ~x481 & ~x501 & ~x506 & ~x507 & ~x528 & ~x565 & ~x621 & ~x626 & ~x648 & ~x665 & ~x676 & ~x682 & ~x696 & ~x728;
assign c5136 =  x746 &  x775 & ~x93 & ~x121 & ~x330 & ~x358 & ~x380 & ~x381 & ~x471;
assign c5138 =  x426 &  x509 & ~x436 & ~x741;
assign c5140 =  x632 & ~x2 & ~x20 & ~x172 & ~x218 & ~x267 & ~x269 & ~x276 & ~x300 & ~x324 & ~x379 & ~x381 & ~x389 & ~x408 & ~x416 & ~x419 & ~x476 & ~x499 & ~x504 & ~x506 & ~x532 & ~x586 & ~x730;
assign c5142 =  x27;
assign c5144 =  x182 &  x237 &  x264 &  x293 &  x512 &  x746 & ~x342 & ~x388 & ~x418 & ~x705;
assign c5146 =  x543 &  x714 &  x717 & ~x303 & ~x436 & ~x466 & ~x472 & ~x492 & ~x763;
assign c5148 =  x274 &  x275 &  x447 & ~x462;
assign c5150 =  x100 & ~x116 & ~x134 & ~x143 & ~x167 & ~x190 & ~x247 & ~x250 & ~x286 & ~x296 & ~x297 & ~x314 & ~x328 & ~x334 & ~x354 & ~x367 & ~x368 & ~x380 & ~x381 & ~x413 & ~x436 & ~x439 & ~x470 & ~x473 & ~x583 & ~x651 & ~x703;
assign c5152 =  x343 &  x360 & ~x459;
assign c5154 =  x414 &  x471 &  x557;
assign c5156 =  x552 &  x576 &  x578 & ~x30 & ~x142 & ~x333 & ~x352 & ~x403;
assign c5158 =  x687 &  x717 &  x719 & ~x109 & ~x165 & ~x173 & ~x359 & ~x360 & ~x436 & ~x443 & ~x472 & ~x494;
assign c5160 =  x759;
assign c5162 =  x457 &  x512 &  x539 & ~x5 & ~x49 & ~x381 & ~x395 & ~x423 & ~x450 & ~x490 & ~x551;
assign c5164 =  x346 & ~x61 & ~x63 & ~x140 & ~x222 & ~x271 & ~x298 & ~x323 & ~x325 & ~x342 & ~x350 & ~x358 & ~x364 & ~x391 & ~x444 & ~x556 & ~x651 & ~x754;
assign c5166 =  x187 &  x189 &  x510;
assign c5168 =  x426 &  x481 &  x536 & ~x123;
assign c5170 =  x431 &  x485 & ~x138 & ~x162 & ~x167 & ~x191 & ~x287 & ~x299 & ~x301 & ~x316 & ~x339 & ~x342 & ~x370 & ~x453 & ~x619 & ~x637 & ~x641 & ~x669 & ~x710 & ~x726 & ~x734 & ~x738;
assign c5172 =  x180 & ~x55 & ~x215 & ~x218 & ~x254 & ~x299 & ~x369 & ~x370 & ~x450 & ~x629 & ~x740;
assign c5174 =  x746 & ~x24 & ~x36 & ~x86 & ~x88 & ~x143 & ~x144 & ~x161 & ~x169 & ~x191 & ~x201 & ~x219 & ~x221 & ~x252 & ~x274 & ~x287 & ~x299 & ~x313 & ~x353 & ~x356 & ~x358 & ~x380 & ~x383 & ~x384 & ~x386 & ~x417 & ~x466 & ~x468 & ~x472 & ~x473 & ~x478 & ~x674 & ~x726 & ~x731 & ~x764;
assign c5176 =  x303 &  x304 & ~x583;
assign c5178 = ~x65 & ~x264 & ~x270 & ~x293 & ~x319 & ~x347 & ~x375 & ~x402 & ~x430 & ~x591 & ~x614;
assign c5180 =  x374 &  x401 & ~x77 & ~x86 & ~x104 & ~x145 & ~x163 & ~x188 & ~x189 & ~x214 & ~x219 & ~x228 & ~x229 & ~x294 & ~x301 & ~x310 & ~x312 & ~x323 & ~x326 & ~x359 & ~x388 & ~x391 & ~x451 & ~x473 & ~x478 & ~x501 & ~x507 & ~x528 & ~x583 & ~x595 & ~x615 & ~x621 & ~x731 & ~x764;
assign c5182 =  x560;
assign c5184 =  x454 &  x510 &  x538 & ~x38 & ~x462 & ~x466 & ~x514 & ~x694 & ~x740;
assign c5186 =  x487 &  x515 &  x629 &  x744 & ~x65 & ~x328 & ~x361 & ~x387;
assign c5188 =  x487 &  x515 &  x542 &  x714 &  x743 & ~x50 & ~x90 & ~x93 & ~x108 & ~x136 & ~x141 & ~x143 & ~x193 & ~x226 & ~x306 & ~x330 & ~x333 & ~x342 & ~x354 & ~x370 & ~x371 & ~x415 & ~x502 & ~x588 & ~x733 & ~x735 & ~x736 & ~x764 & ~x765;
assign c5190 =  x159 &  x188 & ~x403 & ~x557;
assign c5192 =  x485 &  x512 & ~x5 & ~x8 & ~x23 & ~x79 & ~x80 & ~x106 & ~x286 & ~x326 & ~x358 & ~x381 & ~x385 & ~x397 & ~x413 & ~x450 & ~x479 & ~x492 & ~x696;
assign c5194 =  x188 &  x475 & ~x583;
assign c5196 =  x349 &  x405 &  x433 & ~x64 & ~x89 & ~x93 & ~x177 & ~x358 & ~x389 & ~x481 & ~x538 & ~x563 & ~x566 & ~x665 & ~x693 & ~x766;
assign c5198 =  x302 &  x387 &  x530;
assign c5200 = ~x100 & ~x205 & ~x319 & ~x347 & ~x349 & ~x405 & ~x538;
assign c5202 =  x272 &  x330;
assign c5204 =  x327 & ~x548 & ~x715;
assign c5206 =  x481 &  x509 & ~x149 & ~x378 & ~x403 & ~x569 & ~x771;
assign c5208 =  x387 &  x415 &  x473 & ~x688;
assign c5210 = ~x5 & ~x26 & ~x54 & ~x107 & ~x110 & ~x117 & ~x172 & ~x218 & ~x245 & ~x296 & ~x298 & ~x301 & ~x331 & ~x378 & ~x393 & ~x413 & ~x417 & ~x435 & ~x478 & ~x492 & ~x534 & ~x553 & ~x583 & ~x617 & ~x621 & ~x624 & ~x641 & ~x645 & ~x651 & ~x667 & ~x697 & ~x728;
assign c5212 =  x248 &  x419;
assign c5214 =  x423 & ~x270 & ~x293 & ~x347;
assign c5216 =  x334 & ~x459;
assign c5218 =  x374 & ~x5 & ~x20 & ~x21 & ~x58 & ~x84 & ~x106 & ~x112 & ~x138 & ~x145 & ~x170 & ~x183 & ~x185 & ~x199 & ~x211 & ~x253 & ~x276 & ~x281 & ~x286 & ~x309 & ~x312 & ~x342 & ~x415 & ~x419 & ~x451 & ~x499 & ~x504 & ~x527 & ~x556 & ~x598 & ~x679 & ~x682 & ~x699 & ~x706 & ~x708 & ~x755;
assign c5220 =  x760;
assign c5222 =  x209 &  x236 &  x264 &  x320 &  x376 & ~x257 & ~x313 & ~x327 & ~x328 & ~x385;
assign c5224 =  x552 &  x579 &  x608 & ~x45 & ~x109 & ~x169 & ~x375 & ~x444 & ~x446 & ~x473;
assign c5226 =  x514 &  x600 & ~x200 & ~x357 & ~x383 & ~x415 & ~x417 & ~x435 & ~x439 & ~x443 & ~x736;
assign c5228 = ~x21 & ~x54 & ~x58 & ~x75 & ~x142 & ~x161 & ~x172 & ~x186 & ~x187 & ~x188 & ~x244 & ~x294 & ~x298 & ~x310 & ~x314 & ~x330 & ~x334 & ~x368 & ~x379 & ~x424 & ~x441 & ~x449 & ~x469 & ~x476 & ~x533 & ~x535 & ~x562 & ~x564 & ~x569 & ~x614 & ~x643 & ~x668 & ~x674 & ~x694 & ~x700 & ~x703 & ~x729 & ~x753 & ~x755 & ~x765;
assign c5230 =  x433 &  x576 & ~x172 & ~x299 & ~x303 & ~x323 & ~x498 & ~x572;
assign c5232 =  x509 &  x510 &  x537 & ~x90 & ~x356 & ~x464 & ~x543 & ~x767;
assign c5234 =  x415 &  x502;
assign c5236 =  x125 & ~x7 & ~x29 & ~x31 & ~x59 & ~x76 & ~x84 & ~x110 & ~x113 & ~x135 & ~x136 & ~x143 & ~x146 & ~x161 & ~x174 & ~x186 & ~x215 & ~x218 & ~x219 & ~x223 & ~x224 & ~x226 & ~x246 & ~x297 & ~x299 & ~x304 & ~x307 & ~x314 & ~x324 & ~x325 & ~x327 & ~x328 & ~x331 & ~x333 & ~x334 & ~x338 & ~x354 & ~x355 & ~x357 & ~x385 & ~x391 & ~x396 & ~x413 & ~x417 & ~x418 & ~x421 & ~x423 & ~x424 & ~x445 & ~x446 & ~x451 & ~x467 & ~x473 & ~x479 & ~x502 & ~x503 & ~x532 & ~x535 & ~x538 & ~x554 & ~x561 & ~x569 & ~x583 & ~x617 & ~x618 & ~x620 & ~x644 & ~x646 & ~x653 & ~x680 & ~x695 & ~x698 & ~x729 & ~x732 & ~x734 & ~x756;
assign c5238 =  x348 &  x405 & ~x63 & ~x92 & ~x104 & ~x138 & ~x149 & ~x168 & ~x174 & ~x185 & ~x187 & ~x201 & ~x202 & ~x215 & ~x245 & ~x248 & ~x286 & ~x299 & ~x301 & ~x302 & ~x312 & ~x315 & ~x359 & ~x505 & ~x562 & ~x596 & ~x615 & ~x625 & ~x650 & ~x671 & ~x681 & ~x706;
assign c5240 =  x377 &  x632 & ~x214 & ~x269 & ~x271 & ~x352 & ~x356 & ~x357 & ~x380 & ~x414 & ~x510 & ~x583;
assign c5242 =  x304 &  x453 & ~x292;
assign c5244 =  x293 &  x404 &  x460 &  x743 & ~x66 & ~x372;
assign c5246 =  x745 & ~x3 & ~x5 & ~x18 & ~x32 & ~x33 & ~x47 & ~x49 & ~x55 & ~x57 & ~x60 & ~x77 & ~x86 & ~x105 & ~x190 & ~x201 & ~x218 & ~x224 & ~x281 & ~x298 & ~x302 & ~x307 & ~x329 & ~x330 & ~x342 & ~x355 & ~x361 & ~x394 & ~x397 & ~x398 & ~x410 & ~x423 & ~x441 & ~x444 & ~x450 & ~x451 & ~x467 & ~x500 & ~x527 & ~x529 & ~x530 & ~x532 & ~x555 & ~x558 & ~x585 & ~x614 & ~x675 & ~x680 & ~x726 & ~x732 & ~x735 & ~x766 & ~x781;
assign c5248 =  x353;
assign c5250 =  x373 &  x426 &  x510 & ~x572;
assign c5252 =  x601 &  x761;
assign c5254 =  x245 &  x303 &  x390;
assign c5256 =  x327 &  x443;
assign c5258 =  x212 &  x599 &  x714;
assign c5260 =  x331 &  x503;
assign c5262 =  x216 &  x390;
assign c5264 =  x662 &  x690 &  x691 &  x718 & ~x378;
assign c5266 =  x370 &  x389 & ~x319 & ~x458;
assign c5268 = ~x148 & ~x180 & ~x235 & ~x263 & ~x319 & ~x347 & ~x403 & ~x566 & ~x623;
assign c5270 =  x605 & ~x77 & ~x79 & ~x83 & ~x111 & ~x112 & ~x203 & ~x227 & ~x230 & ~x241 & ~x247 & ~x272 & ~x324 & ~x383 & ~x386 & ~x446 & ~x473 & ~x527 & ~x600 & ~x655 & ~x749;
assign c5272 =  x557;
assign c5274 =  x424 & ~x294 & ~x319;
assign c5276 =  x188 &  x481;
assign c5278 =  x98 &  x749 & ~x381 & ~x411 & ~x435 & ~x763;
assign c5280 =  x266 &  x404 &  x567 &  x568 & ~x548;
assign c5282 =  x283;
assign c5284 =  x376 &  x404 &  x687 & ~x202 & ~x228 & ~x270 & ~x273 & ~x286 & ~x324 & ~x342 & ~x708 & ~x709;
assign c5286 =  x97 & ~x244 & ~x271 & ~x470 & ~x543 & ~x568 & ~x710;
assign c5288 =  x510 & ~x110 & ~x145 & ~x224 & ~x347 & ~x348 & ~x432 & ~x451 & ~x557 & ~x588 & ~x712 & ~x774;
assign c5290 =  x459 &  x686 &  x687 & ~x16 & ~x29 & ~x80 & ~x88 & ~x89 & ~x106 & ~x164 & ~x165 & ~x193 & ~x197 & ~x201 & ~x202 & ~x220 & ~x230 & ~x232 & ~x251 & ~x252 & ~x276 & ~x277 & ~x283 & ~x299 & ~x302 & ~x311 & ~x325 & ~x330 & ~x331 & ~x335 & ~x358 & ~x389 & ~x413 & ~x419 & ~x479 & ~x501 & ~x556 & ~x583 & ~x762;
assign c5292 =  x237 &  x321 &  x377 &  x404 & ~x93 & ~x148 & ~x172 & ~x173 & ~x373 & ~x397 & ~x425 & ~x428 & ~x453 & ~x482 & ~x707;
assign c5294 =  x348 & ~x37 & ~x77 & ~x80 & ~x90 & ~x105 & ~x115 & ~x132 & ~x142 & ~x172 & ~x173 & ~x191 & ~x193 & ~x215 & ~x217 & ~x218 & ~x226 & ~x232 & ~x249 & ~x251 & ~x275 & ~x277 & ~x299 & ~x300 & ~x301 & ~x307 & ~x330 & ~x331 & ~x333 & ~x334 & ~x340 & ~x360 & ~x361 & ~x363 & ~x365 & ~x370 & ~x371 & ~x388 & ~x390 & ~x394 & ~x413 & ~x414 & ~x416 & ~x422 & ~x424 & ~x506 & ~x507 & ~x528 & ~x534 & ~x555 & ~x566 & ~x570 & ~x571 & ~x588 & ~x596 & ~x620 & ~x623 & ~x626 & ~x640 & ~x641 & ~x646 & ~x648 & ~x650 & ~x651 & ~x674 & ~x693 & ~x696 & ~x703 & ~x709 & ~x726 & ~x728 & ~x729 & ~x731 & ~x737 & ~x762 & ~x767 & ~x779 & ~x780 & ~x781 & ~x783;
assign c5296 = ~x38 & ~x93 & ~x150 & ~x180 & ~x235 & ~x265 & ~x320 & ~x403 & ~x457;
assign c5298 =  x424 &  x452 & ~x319;
assign c5300 = ~x209 & ~x263 & ~x291 & ~x347 & ~x351 & ~x514 & ~x540 & ~x676 & ~x743;
assign c5302 =  x319 &  x347 &  x375 & ~x163 & ~x189 & ~x297 & ~x339 & ~x340 & ~x369 & ~x413 & ~x423 & ~x445 & ~x499 & ~x514 & ~x570 & ~x619 & ~x648 & ~x682 & ~x759;
assign c5304 = ~x84 & ~x167 & ~x216 & ~x266 & ~x275 & ~x302 & ~x326 & ~x339 & ~x342 & ~x358 & ~x360 & ~x378 & ~x383 & ~x388 & ~x413 & ~x436 & ~x473 & ~x526 & ~x555 & ~x622 & ~x668 & ~x758;
assign c5306 =  x375 & ~x63 & ~x76 & ~x218 & ~x227 & ~x272 & ~x284 & ~x303 & ~x342 & ~x421 & ~x480 & ~x524 & ~x535 & ~x538 & ~x543 & ~x566 & ~x599 & ~x650 & ~x654 & ~x696 & ~x709 & ~x761 & ~x765;
assign c5308 =  x578 & ~x134 & ~x138 & ~x140 & ~x142 & ~x158 & ~x161 & ~x166 & ~x174 & ~x241 & ~x270 & ~x274 & ~x276 & ~x278 & ~x283 & ~x326 & ~x361 & ~x386 & ~x414 & ~x416 & ~x472 & ~x476 & ~x534 & ~x558 & ~x598 & ~x701 & ~x736;
assign c5310 =  x357 &  x501;
assign c5312 =  x264 &  x431 &  x485 & ~x3 & ~x7 & ~x105 & ~x117 & ~x164 & ~x255 & ~x257 & ~x258 & ~x275 & ~x285 & ~x287 & ~x298 & ~x306 & ~x310 & ~x313 & ~x326 & ~x329 & ~x330 & ~x353 & ~x356 & ~x358 & ~x365 & ~x367 & ~x370 & ~x371 & ~x383 & ~x384 & ~x423 & ~x505 & ~x652 & ~x669 & ~x676 & ~x709 & ~x736 & ~x762;
assign c5314 =  x687 &  x718 & ~x166 & ~x330 & ~x331 & ~x358 & ~x361 & ~x384 & ~x414 & ~x465 & ~x492 & ~x764;
assign c5316 =  x441 & ~x294 & ~x319 & ~x418 & ~x430;
assign c5318 =  x451 & ~x264 & ~x430;
assign c5320 =  x281 &  x615;
assign c5322 =  x606;
assign c5324 =  x315 &  x416 &  x426 & ~x458;
assign c5326 =  x131 &  x426;
assign c5328 =  x415;
assign c5330 =  x541 &  x568 &  x713 &  x742 &  x743 & ~x33 & ~x115 & ~x142 & ~x247 & ~x326 & ~x353 & ~x354 & ~x383 & ~x414 & ~x415 & ~x441 & ~x707 & ~x735 & ~x736;
assign c5332 =  x396 & ~x319;
assign c5334 =  x376 &  x460 & ~x88 & ~x271 & ~x301 & ~x306 & ~x332 & ~x444 & ~x656 & ~x684 & ~x712 & ~x736;
assign c5336 =  x30;
assign c5338 =  x300 &  x358 & ~x656 & ~x771;
assign c5340 =  x320 &  x349 & ~x26 & ~x38 & ~x80 & ~x93 & ~x116 & ~x136 & ~x189 & ~x217 & ~x220 & ~x250 & ~x253 & ~x286 & ~x287 & ~x297 & ~x299 & ~x300 & ~x301 & ~x304 & ~x362 & ~x365 & ~x385 & ~x396 & ~x411 & ~x415 & ~x424 & ~x499 & ~x529 & ~x620 & ~x627 & ~x638 & ~x654 & ~x668 & ~x682 & ~x683 & ~x697 & ~x707 & ~x726 & ~x727 & ~x736 & ~x737 & ~x758 & ~x760;
assign c5342 =  x96 & ~x30 & ~x104 & ~x132 & ~x142 & ~x171 & ~x215 & ~x240 & ~x299 & ~x331 & ~x379 & ~x412 & ~x413 & ~x416 & ~x447 & ~x498 & ~x506 & ~x555 & ~x640 & ~x649 & ~x650 & ~x652 & ~x676 & ~x700 & ~x708 & ~x729 & ~x765;
assign c5344 =  x248 &  x251;
assign c5346 =  x340 & ~x289 & ~x374 & ~x510;
assign c5348 =  x161 &  x198 &  x419;
assign c5350 =  x339 &  x423 & ~x209 & ~x263;
assign c5352 =  x237 &  x348 &  x375 &  x376 & ~x88 & ~x133 & ~x190 & ~x254 & ~x334 & ~x342 & ~x362 & ~x425 & ~x478 & ~x479 & ~x566 & ~x677 & ~x697 & ~x710 & ~x757;
assign c5354 =  x761;
assign c5356 = ~x9 & ~x35 & ~x77 & ~x143 & ~x270 & ~x325 & ~x351 & ~x379 & ~x383 & ~x421 & ~x436 & ~x438 & ~x520 & ~x527 & ~x551 & ~x576 & ~x610 & ~x611 & ~x706 & ~x708;
assign c5358 =  x163 &  x357;
assign c5360 =  x778;
assign c5362 =  x405 &  x687 & ~x57 & ~x115 & ~x116 & ~x147 & ~x170 & ~x189 & ~x191 & ~x194 & ~x204 & ~x222 & ~x229 & ~x246 & ~x247 & ~x258 & ~x286 & ~x287 & ~x327 & ~x328 & ~x329 & ~x358 & ~x361 & ~x362 & ~x368 & ~x372 & ~x373 & ~x389 & ~x416 & ~x427 & ~x454 & ~x529 & ~x534 & ~x535 & ~x707 & ~x779;
assign c5364 =  x605 &  x606 &  x633 & ~x49 & ~x59 & ~x83 & ~x104 & ~x105 & ~x162 & ~x185 & ~x195 & ~x243 & ~x257 & ~x276 & ~x279 & ~x282 & ~x297 & ~x386 & ~x390 & ~x397 & ~x413 & ~x419 & ~x424 & ~x536 & ~x561 & ~x681 & ~x727 & ~x736 & ~x751 & ~x760;
assign c5366 =  x212 &  x213 &  x571 &  x599 & ~x275 & ~x441 & ~x558;
assign c5368 =  x515 &  x543 &  x776 & ~x436 & ~x520;
assign c5370 =  x571 &  x750;
assign c5372 =  x487 &  x601 &  x748;
assign c5374 =  x414 &  x471 & ~x218;
assign c5376 =  x211 &  x293 &  x405 &  x545 &  x687 & ~x370;
assign c5378 =  x460 &  x515 &  x659 &  x745 & ~x218 & ~x248 & ~x358 & ~x361 & ~x366 & ~x384 & ~x393 & ~x413;
assign c5380 =  x235 &  x263 & ~x88 & ~x131 & ~x134 & ~x215 & ~x218 & ~x274 & ~x295 & ~x325 & ~x384 & ~x596 & ~x652 & ~x694 & ~x752 & ~x753;
assign c5382 =  x552 &  x580 &  x635 & ~x137 & ~x306 & ~x358 & ~x757;
assign c5384 =  x329 &  x415 &  x501;
assign c5386 =  x443 &  x471 &  x499 & ~x129 & ~x133 & ~x275 & ~x688;
assign c5388 =  x385 &  x414 &  x472 &  x556 & ~x546;
assign c5390 =  x370 &  x398 &  x453 & ~x347 & ~x430 & ~x485;
assign c5392 =  x315 &  x371 & ~x208 & ~x435 & ~x458;
assign c5394 =  x188 &  x199 &  x302;
assign c5396 =  x373 &  x401 & ~x110 & ~x210 & ~x267 & ~x271 & ~x293 & ~x358 & ~x652;
assign c5398 =  x358 &  x415 & ~x716;
assign c5400 =  x333 &  x390 & ~x98 & ~x208 & ~x235 & ~x459;
assign c5402 =  x215 &  x244 &  x388;
assign c5404 = ~x97 & ~x299 & ~x319 & ~x323 & ~x489 & ~x620;
assign c5406 =  x190 &  x589;
assign c5408 =  x745 &  x746 & ~x135 & ~x219 & ~x220 & ~x246 & ~x284 & ~x302 & ~x342 & ~x355 & ~x385 & ~x407 & ~x468 & ~x492 & ~x494 & ~x522;
assign c5410 =  x441;
assign c5412 =  x360 &  x426 &  x562 & ~x571;
assign c5414 =  x273 &  x388;
assign c5416 =  x284 &  x397 & ~x347;
assign c5418 = ~x138 & ~x165 & ~x188 & ~x211 & ~x215 & ~x217 & ~x219 & ~x239 & ~x247 & ~x254 & ~x257 & ~x270 & ~x271 & ~x287 & ~x294 & ~x325 & ~x326 & ~x355 & ~x358 & ~x361 & ~x369 & ~x383 & ~x388 & ~x417 & ~x419 & ~x423 & ~x499 & ~x508 & ~x560 & ~x584 & ~x587 & ~x597 & ~x643 & ~x645 & ~x651 & ~x705 & ~x732 & ~x736;
assign c5420 =  x24;
assign c5422 =  x239 &  x350 &  x545 &  x773;
assign c5424 =  x209 &  x348 & ~x3 & ~x27 & ~x32 & ~x60 & ~x107 & ~x200 & ~x202 & ~x270 & ~x299 & ~x301 & ~x335 & ~x360 & ~x365 & ~x368 & ~x369 & ~x397 & ~x425 & ~x448 & ~x451 & ~x534 & ~x535 & ~x542 & ~x560 & ~x567 & ~x569 & ~x570 & ~x593 & ~x596 & ~x597 & ~x611 & ~x621 & ~x622 & ~x650 & ~x653 & ~x669 & ~x678 & ~x679 & ~x705 & ~x708 & ~x710 & ~x726 & ~x738 & ~x761 & ~x783;
assign c5426 =  x2;
assign c5428 =  x780;
assign c5430 =  x385 &  x414 &  x443 & ~x185 & ~x712 & ~x713;
assign c5432 =  x746 &  x747 & ~x9 & ~x81 & ~x247 & ~x249 & ~x274 & ~x306 & ~x326 & ~x331 & ~x382 & ~x408 & ~x417 & ~x499 & ~x527 & ~x577 & ~x729;
assign c5434 =  x773 &  x775 & ~x410 & ~x466;
assign c5436 = ~x39 & ~x97 & ~x150 & ~x153 & ~x209 & ~x263 & ~x325 & ~x430 & ~x440 & ~x458 & ~x593 & ~x649;
assign c5438 =  x424 & ~x263;
assign c5440 =  x228 &  x371 &  x388;
assign c5442 =  x747 &  x776 & ~x302 & ~x330 & ~x436 & ~x470 & ~x709;
assign c5444 =  x348 &  x375 &  x376 & ~x25 & ~x54 & ~x65 & ~x103 & ~x106 & ~x163 & ~x170 & ~x219 & ~x271 & ~x272 & ~x274 & ~x284 & ~x301 & ~x303 & ~x304 & ~x343 & ~x357 & ~x358 & ~x360 & ~x367 & ~x370 & ~x388 & ~x419 & ~x425 & ~x445 & ~x449 & ~x450 & ~x471 & ~x479 & ~x533 & ~x534 & ~x570 & ~x594 & ~x619 & ~x622 & ~x624 & ~x626 & ~x641 & ~x647 & ~x676 & ~x678 & ~x704 & ~x705 & ~x734 & ~x736 & ~x764;
assign c5446 =  x644;
assign c5448 =  x189 & ~x321 & ~x530;
assign c5450 =  x376 &  x431 &  x629 &  x743 & ~x91 & ~x359 & ~x470;
assign c5452 =  x760;
assign c5454 =  x431 &  x457 & ~x47 & ~x92 & ~x217 & ~x229 & ~x259 & ~x270 & ~x276 & ~x283 & ~x330 & ~x386 & ~x417 & ~x504 & ~x597 & ~x651 & ~x693 & ~x761 & ~x763;
assign c5456 =  x457 &  x485 &  x512 &  x539 &  x540 &  x567 & ~x547 & ~x552;
assign c5458 =  x438 &  x454;
assign c5460 = ~x21 & ~x23 & ~x59 & ~x76 & ~x80 & ~x104 & ~x135 & ~x140 & ~x162 & ~x165 & ~x174 & ~x201 & ~x202 & ~x222 & ~x244 & ~x247 & ~x249 & ~x259 & ~x272 & ~x285 & ~x296 & ~x297 & ~x298 & ~x306 & ~x309 & ~x312 & ~x314 & ~x324 & ~x338 & ~x379 & ~x383 & ~x385 & ~x396 & ~x397 & ~x408 & ~x410 & ~x412 & ~x413 & ~x441 & ~x452 & ~x469 & ~x500 & ~x583 & ~x585 & ~x592 & ~x594 & ~x611 & ~x627 & ~x666 & ~x672 & ~x680 & ~x703 & ~x709 & ~x725 & ~x736 & ~x759;
assign c5462 = ~x235 & ~x293 & ~x319 & ~x374 & ~x378 & ~x403 & ~x678;
assign c5464 =  x368 & ~x265 & ~x347 & ~x457 & ~x459 & ~x566;
assign c5466 =  x606 & ~x1 & ~x26 & ~x50 & ~x59 & ~x84 & ~x89 & ~x90 & ~x110 & ~x167 & ~x169 & ~x171 & ~x173 & ~x177 & ~x191 & ~x218 & ~x225 & ~x230 & ~x253 & ~x280 & ~x300 & ~x306 & ~x312 & ~x314 & ~x334 & ~x335 & ~x365 & ~x411 & ~x413 & ~x417 & ~x418 & ~x424 & ~x500 & ~x502 & ~x527 & ~x533 & ~x588 & ~x592 & ~x617 & ~x655 & ~x708 & ~x754 & ~x759 & ~x763;
assign c5468 =  x298 &  x356;
assign c5470 =  x377 &  x404 &  x658 & ~x37 & ~x80 & ~x86 & ~x90 & ~x92 & ~x119 & ~x134 & ~x146 & ~x175 & ~x177 & ~x230 & ~x256 & ~x258 & ~x310 & ~x330 & ~x335 & ~x368 & ~x369 & ~x370 & ~x412 & ~x420 & ~x423 & ~x424 & ~x426 & ~x451 & ~x505 & ~x508 & ~x669 & ~x681 & ~x704 & ~x708 & ~x723 & ~x735;
assign c5472 =  x19 &  x192;
assign c5474 =  x474;
assign c5476 =  x293 &  x403 &  x457 & ~x36 & ~x314 & ~x342 & ~x343 & ~x676;
assign c5478 =  x246 &  x503;
assign c5480 =  x543 &  x688 &  x717 & ~x386 & ~x465;
assign c5482 =  x485 & ~x25 & ~x31 & ~x162 & ~x172 & ~x189 & ~x228 & ~x232 & ~x325 & ~x330 & ~x339 & ~x343 & ~x352 & ~x357 & ~x358 & ~x364 & ~x534 & ~x596 & ~x597 & ~x645 & ~x669 & ~x708 & ~x722 & ~x726 & ~x737 & ~x752 & ~x764;
assign c5484 =  x389 &  x534 & ~x235;
assign c5486 =  x304 & ~x98 & ~x293 & ~x430 & ~x541;
assign c5488 =  x71 & ~x53 & ~x60 & ~x107 & ~x108 & ~x109 & ~x110 & ~x140 & ~x163 & ~x200 & ~x201 & ~x219 & ~x221 & ~x224 & ~x229 & ~x239 & ~x246 & ~x272 & ~x276 & ~x282 & ~x299 & ~x301 & ~x314 & ~x327 & ~x328 & ~x332 & ~x334 & ~x359 & ~x383 & ~x387 & ~x417 & ~x421 & ~x445 & ~x446 & ~x452 & ~x502 & ~x527 & ~x534 & ~x536 & ~x560 & ~x562 & ~x599 & ~x619 & ~x668 & ~x674 & ~x683 & ~x697 & ~x710 & ~x735 & ~x755;
assign c5490 =  x301 &  x387 &  x388 &  x502;
assign c5492 =  x172 &  x469;
assign c5494 =  x413 &  x499 & ~x129 & ~x716;
assign c5496 =  x552 &  x635 & ~x319 & ~x416;
assign c5498 =  x240 &  x487 & ~x435 & ~x496;
assign c51 =  x533 &  x593;
assign c53 =  x158 & ~x6 & ~x28 & ~x55 & ~x473 & ~x627 & ~x644 & ~x748 & ~x749 & ~x751 & ~x753;
assign c55 =  x652 & ~x98 & ~x127;
assign c57 =  x381 & ~x79 & ~x82 & ~x261 & ~x725;
assign c59 =  x380 &  x408;
assign c511 =  x278 &  x306 & ~x454 & ~x482 & ~x560 & ~x618 & ~x648 & ~x704 & ~x705;
assign c513 =  x175 & ~x2 & ~x18 & ~x239 & ~x298 & ~x548 & ~x644 & ~x674 & ~x693 & ~x696 & ~x731 & ~x749;
assign c515 =  x184 & ~x460 & ~x481 & ~x484 & ~x591 & ~x748 & ~x751 & ~x765;
assign c517 =  x556 &  x582 &  x583 & ~x31 & ~x469;
assign c519 =  x202 &  x312 &  x535 & ~x95 & ~x364 & ~x672 & ~x760;
assign c521 =  x638 & ~x140 & ~x279 & ~x490 & ~x514 & ~x574 & ~x606;
assign c523 =  x407 & ~x318;
assign c525 =  x483 &  x517;
assign c527 =  x128 &  x409;
assign c529 =  x653 & ~x28 & ~x108 & ~x410 & ~x735 & ~x765;
assign c531 =  x466 &  x494;
assign c533 =  x353 & ~x21 & ~x50 & ~x529;
assign c535 =  x654 & ~x10 & ~x67 & ~x213 & ~x477 & ~x725;
assign c537 =  x80;
assign c539 =  x146 &  x174 &  x201 & ~x15 & ~x24 & ~x317 & ~x503;
assign c541 =  x296 & ~x21 & ~x196 & ~x530 & ~x588 & ~x751 & ~x753 & ~x760;
assign c543 =  x80;
assign c545 =  x123 & ~x33 & ~x463 & ~x485 & ~x572 & ~x751;
assign c547 =  x505 & ~x56 & ~x388 & ~x672;
assign c549 =  x179 &  x180 & ~x399 & ~x403 & ~x482 & ~x509;
assign c551 =  x317 & ~x0 & ~x7 & ~x223 & ~x456 & ~x541 & ~x548 & ~x591 & ~x592 & ~x722 & ~x761;
assign c553 =  x546 & ~x12 & ~x130 & ~x710 & ~x720 & ~x757;
assign c555 =  x682 & ~x767;
assign c557 =  x491 & ~x631 & ~x699;
assign c559 =  x319 &  x422;
assign c561 =  x133 & ~x509 & ~x545;
assign c563 =  x737;
assign c565 =  x572 & ~x41 & ~x78 & ~x83 & ~x84 & ~x636 & ~x753;
assign c567 =  x296 & ~x52 & ~x168 & ~x314 & ~x753;
assign c569 =  x463 &  x491 & ~x2 & ~x102 & ~x586 & ~x755;
assign c571 =  x79;
assign c573 =  x148 & ~x2 & ~x3 & ~x8 & ~x26 & ~x34 & ~x35 & ~x45 & ~x56 & ~x98 & ~x196 & ~x214 & ~x223 & ~x266 & ~x336 & ~x615 & ~x647 & ~x757;
assign c575 =  x175 &  x535 & ~x421 & ~x503 & ~x701 & ~x702 & ~x729 & ~x761;
assign c577 =  x517 & ~x3 & ~x76 & ~x436 & ~x660;
assign c579 =  x516 & ~x0 & ~x7 & ~x21 & ~x36 & ~x47 & ~x52 & ~x59 & ~x60 & ~x83 & ~x110 & ~x111 & ~x169 & ~x381 & ~x411 & ~x607 & ~x611 & ~x664 & ~x685 & ~x692 & ~x702 & ~x713 & ~x748 & ~x750 & ~x751 & ~x762 & ~x764 & ~x768 & ~x773 & ~x778;
assign c581 =  x434 & ~x24 & ~x128 & ~x235;
assign c583 =  x517 &  x566;
assign c585 =  x205 &  x232 &  x286 & ~x91 & ~x174;
assign c587 =  x261 &  x288 & ~x12 & ~x55 & ~x68 & ~x168 & ~x493 & ~x677 & ~x751;
assign c589 =  x572 & ~x7 & ~x49 & ~x86 & ~x110 & ~x183 & ~x609 & ~x666 & ~x690 & ~x719 & ~x730 & ~x751 & ~x775;
assign c591 =  x365 & ~x140 & ~x481 & ~x592;
assign c593 =  x736;
assign c595 =  x679 & ~x703;
assign c597 =  x325 & ~x87 & ~x530 & ~x673 & ~x693 & ~x695 & ~x701 & ~x729 & ~x757;
assign c599 =  x64 &  x91 & ~x16 & ~x54 & ~x503 & ~x761;
assign c5101 =  x149 & ~x168 & ~x224 & ~x619 & ~x629 & ~x703 & ~x730 & ~x757 & ~x775;
assign c5103 =  x465 & ~x6 & ~x52 & ~x261 & ~x755 & ~x761;
assign c5105 =  x381 & ~x363 & ~x666 & ~x778;
assign c5107 =  x352 & ~x545 & ~x641;
assign c5109 =  x353 &  x381 & ~x509;
assign c5111 =  x678 & ~x16 & ~x248 & ~x364 & ~x634;
assign c5113 =  x289 & ~x88 & ~x92 & ~x481 & ~x575;
assign c5115 =  x296 & ~x420 & ~x503 & ~x572 & ~x602 & ~x627;
assign c5117 =  x735;
assign c5119 =  x519 &  x546 & ~x0 & ~x19 & ~x63 & ~x662;
assign c5121 = ~x60 & ~x260 & ~x277 & ~x399 & ~x408 & ~x603 & ~x631 & ~x660 & ~x746 & ~x776;
assign c5123 =  x650 & ~x82 & ~x195 & ~x605 & ~x662;
assign c5125 =  x488 & ~x13 & ~x26 & ~x101 & ~x128 & ~x308 & ~x554 & ~x609 & ~x641 & ~x643 & ~x698 & ~x723 & ~x741;
assign c5127 =  x238 &  x317 & ~x49 & ~x51 & ~x80 & ~x483 & ~x650 & ~x673 & ~x696 & ~x726;
assign c5129 =  x317 & ~x4 & ~x64 & ~x111 & ~x113 & ~x142 & ~x146 & ~x253 & ~x483 & ~x538 & ~x549 & ~x551 & ~x697 & ~x703 & ~x732 & ~x735 & ~x753 & ~x775;
assign c5131 =  x736;
assign c5133 =  x325 & ~x24 & ~x28 & ~x226 & ~x336 & ~x364 & ~x392 & ~x517 & ~x643 & ~x733 & ~x736;
assign c5135 =  x769 & ~x684;
assign c5137 =  x389 &  x631 & ~x35 & ~x52 & ~x364 & ~x743;
assign c5139 =  x464 &  x492 &  x519 &  x547;
assign c5141 =  x262 &  x554;
assign c5143 =  x464 &  x492;
assign c5145 =  x232 & ~x31 & ~x65 & ~x127 & ~x128 & ~x269 & ~x420 & ~x554 & ~x614 & ~x675 & ~x722 & ~x777;
assign c5147 =  x570 & ~x197 & ~x691 & ~x733 & ~x775;
assign c5149 =  x241 &  x269 & ~x26 & ~x91 & ~x171 & ~x172 & ~x308 & ~x485 & ~x597;
assign c5151 =  x322 & ~x254 & ~x279 & ~x492;
assign c5153 =  x175 &  x488 & ~x41 & ~x105 & ~x107 & ~x697;
assign c5155 =  x144 & ~x19 & ~x310;
assign c5157 =  x261 & ~x229 & ~x491 & ~x511 & ~x643 & ~x673 & ~x685 & ~x727 & ~x750 & ~x783;
assign c5159 = ~x56 & ~x127 & ~x234 & ~x346 & ~x366 & ~x443 & ~x473 & ~x691 & ~x744 & ~x755;
assign c5161 =  x278 & ~x2 & ~x83 & ~x275 & ~x303 & ~x672 & ~x759 & ~x761;
assign c5163 =  x262 &  x527;
assign c5165 =  x380 & ~x596 & ~x681 & ~x724;
assign c5167 =  x535 &  x651;
assign c5169 =  x70 &  x266 & ~x82 & ~x376;
assign c5171 =  x259 & ~x16 & ~x46 & ~x79 & ~x240 & ~x279 & ~x294 & ~x647 & ~x666 & ~x674 & ~x699 & ~x723 & ~x765 & ~x780;
assign c5173 =  x260 &  x597 & ~x127;
assign c5175 =  x707 & ~x606;
assign c5177 =  x260 &  x287 & ~x30 & ~x55 & ~x130 & ~x142 & ~x173 & ~x450 & ~x670 & ~x723 & ~x749 & ~x756;
assign c5179 =  x609 &  x610 & ~x307 & ~x335 & ~x488 & ~x629 & ~x681;
assign c5181 =  x257 &  x631 & ~x1 & ~x30 & ~x81 & ~x84 & ~x752;
assign c5183 =  x381 & ~x12 & ~x250;
assign c5185 =  x362 & ~x23 & ~x33 & ~x34 & ~x55 & ~x72 & ~x87 & ~x114 & ~x140 & ~x166 & ~x385 & ~x507 & ~x511 & ~x535 & ~x538 & ~x590 & ~x594 & ~x653 & ~x679 & ~x725 & ~x746 & ~x747 & ~x763 & ~x773 & ~x782;
assign c5187 =  x151 &  x178 &  x205 & ~x484;
assign c5189 =  x36;
assign c5191 =  x103 &  x556;
assign c5193 =  x352 & ~x26 & ~x49 & ~x557 & ~x754 & ~x761;
assign c5195 =  x202 &  x488 & ~x19 & ~x43 & ~x136 & ~x138 & ~x392 & ~x585 & ~x642 & ~x670 & ~x671 & ~x699 & ~x703 & ~x726 & ~x728 & ~x753 & ~x767 & ~x781 & ~x782;
assign c5197 =  x127 &  x437;
assign c5199 =  x233 &  x286 & ~x2 & ~x5 & ~x6 & ~x7 & ~x26 & ~x31 & ~x53 & ~x79 & ~x112 & ~x117 & ~x364 & ~x381 & ~x385 & ~x677 & ~x705 & ~x725 & ~x764 & ~x776;
assign c5201 =  x150 & ~x43 & ~x483 & ~x485 & ~x519 & ~x761 & ~x782;
assign c5203 =  x323 & ~x178 & ~x196 & ~x433;
assign c5205 =  x627 & ~x354 & ~x393 & ~x697 & ~x711 & ~x731 & ~x733;
assign c5207 =  x458 &  x459 & ~x41 & ~x49 & ~x584 & ~x674;
assign c5209 =  x208 &  x555 & ~x82 & ~x226 & ~x494 & ~x629;
assign c5211 =  x68 & ~x456 & ~x629;
assign c5213 =  x324 &  x352 & ~x164 & ~x336;
assign c5215 =  x546 & ~x20 & ~x103 & ~x131 & ~x158 & ~x161 & ~x382 & ~x607 & ~x751;
assign c5217 =  x435 & ~x509 & ~x576;
assign c5219 =  x621 &  x649 & ~x26 & ~x56 & ~x85 & ~x249 & ~x254 & ~x604 & ~x671;
assign c5221 =  x65 & ~x58 & ~x138 & ~x281 & ~x308 & ~x419 & ~x503 & ~x544 & ~x598 & ~x599 & ~x604 & ~x782;
assign c5223 =  x214 &  x554 &  x581 & ~x690;
assign c5225 = ~x317 & ~x539;
assign c5227 =  x306 & ~x481 & ~x551 & ~x591 & ~x593;
assign c5229 =  x666 & ~x23 & ~x194 & ~x225 & ~x574 & ~x629 & ~x660 & ~x672 & ~x683 & ~x711 & ~x756 & ~x780 & ~x781;
assign c5231 =  x611 &  x638 & ~x280 & ~x439;
assign c5233 =  x208 & ~x4 & ~x43 & ~x55 & ~x82 & ~x485 & ~x649 & ~x650 & ~x672 & ~x723 & ~x730 & ~x769 & ~x777 & ~x781;
assign c5235 = ~x0 & ~x2 & ~x3 & ~x30 & ~x56 & ~x111 & ~x224 & ~x399 & ~x427 & ~x449 & ~x463 & ~x481 & ~x487 & ~x515 & ~x521 & ~x532 & ~x547 & ~x562 & ~x599 & ~x672 & ~x676 & ~x703 & ~x731 & ~x732;
assign c5237 =  x267 &  x317;
assign c5239 =  x123 &  x232 & ~x90 & ~x684;
assign c5241 =  x67;
assign c5243 =  x627 & ~x158 & ~x751 & ~x765;
assign c5245 =  x261 &  x660 & ~x7 & ~x20 & ~x28 & ~x637 & ~x666 & ~x676 & ~x698 & ~x722 & ~x723 & ~x724 & ~x749 & ~x757;
assign c5247 = ~x29 & ~x36 & ~x55 & ~x59 & ~x62 & ~x64 & ~x86 & ~x92 & ~x112 & ~x167 & ~x229 & ~x377 & ~x484 & ~x489 & ~x509 & ~x558 & ~x622 & ~x647 & ~x669 & ~x672 & ~x695 & ~x725 & ~x758 & ~x777 & ~x778;
assign c5249 =  x94 & ~x254 & ~x549;
assign c5251 =  x122 & ~x625 & ~x629 & ~x672 & ~x731;
assign c5253 =  x287 & ~x16 & ~x37 & ~x48 & ~x51 & ~x59 & ~x82 & ~x86 & ~x168 & ~x171 & ~x317 & ~x394 & ~x559 & ~x560 & ~x587 & ~x605 & ~x617 & ~x672 & ~x698 & ~x699 & ~x755 & ~x768 & ~x783;
assign c5255 =  x178 &  x179 &  x180 & ~x23 & ~x146 & ~x751;
assign c5257 =  x465 &  x483 & ~x21 & ~x47 & ~x783;
assign c5259 = ~x10 & ~x19 & ~x37 & ~x72 & ~x86 & ~x101 & ~x279 & ~x381 & ~x559 & ~x560 & ~x607 & ~x616 & ~x644 & ~x652 & ~x653 & ~x659 & ~x668 & ~x759 & ~x763 & ~x771;
assign c5261 =  x204 &  x205 & ~x29 & ~x36 & ~x116 & ~x252 & ~x421 & ~x586 & ~x615 & ~x672 & ~x676 & ~x711 & ~x754 & ~x757 & ~x780;
assign c5263 =  x145 &  x146 & ~x95 & ~x134 & ~x154;
assign c5265 =  x154 &  x179 & ~x402 & ~x481;
assign c5267 =  x296 & ~x203 & ~x281 & ~x601 & ~x713 & ~x747;
assign c5269 =  x289 &  x527 & ~x6 & ~x86 & ~x89 & ~x223;
assign c5271 =  x372 &  x546 & ~x7 & ~x746 & ~x782;
assign c5273 =  x533 &  x561 & ~x249 & ~x361 & ~x391;
assign c5275 = ~x22 & ~x34 & ~x220 & ~x290 & ~x345 & ~x437 & ~x463 & ~x470 & ~x662 & ~x687 & ~x774;
assign c5277 =  x434 &  x684;
assign c5279 =  x290 &  x318 & ~x359 & ~x385 & ~x456 & ~x511 & ~x520 & ~x589;
assign c5281 =  x262 &  x445 & ~x4 & ~x12 & ~x23 & ~x142 & ~x760;
assign c5283 =  x465 & ~x2 & ~x23 & ~x26 & ~x58 & ~x163 & ~x165 & ~x250 & ~x261 & ~x554 & ~x560 & ~x586;
assign c5285 =  x707 & ~x633 & ~x757;
assign c5287 =  x709 &  x710;
assign c5289 =  x325 & ~x111 & ~x454 & ~x569 & ~x644;
assign c5291 =  x230 &  x282 & ~x96 & ~x337 & ~x641;
assign c5293 =  x254 & ~x45 & ~x301;
assign c5295 = ~x19 & ~x24 & ~x408 & ~x480 & ~x481 & ~x495 & ~x509 & ~x571 & ~x622 & ~x744 & ~x755 & ~x773;
assign c5297 =  x527 & ~x29 & ~x57 & ~x88 & ~x142 & ~x194 & ~x198 & ~x279 & ~x412 & ~x560;
assign c5299 =  x479 &  x593 & ~x40 & ~x223 & ~x365 & ~x420 & ~x647 & ~x692;
assign c5301 =  x709;
assign c5303 =  x230 &  x604 & ~x7;
assign c5305 =  x638 & ~x196 & ~x335 & ~x517 & ~x548 & ~x629 & ~x653 & ~x728 & ~x780 & ~x781;
assign c5307 =  x206 &  x207 & ~x116 & ~x172 & ~x174 & ~x409 & ~x655 & ~x684 & ~x725 & ~x751 & ~x783;
assign c5309 = ~x0 & ~x8 & ~x9 & ~x261 & ~x308 & ~x463 & ~x503 & ~x604 & ~x742 & ~x748 & ~x778 & ~x779;
assign c5311 =  x435 & ~x513;
assign c5313 =  x740;
assign c5315 =  x79;
assign c5317 =  x458 & ~x10 & ~x39 & ~x106 & ~x136 & ~x555 & ~x558 & ~x617 & ~x637 & ~x672 & ~x691 & ~x692 & ~x761 & ~x770 & ~x775;
assign c5319 =  x262 &  x554;
assign c5321 =  x260 &  x261 &  x262 & ~x8 & ~x12 & ~x22 & ~x58 & ~x64 & ~x130 & ~x198 & ~x674 & ~x722 & ~x754 & ~x757 & ~x759 & ~x780;
assign c5323 =  x232 & ~x75 & ~x102 & ~x154 & ~x317 & ~x610 & ~x767;
assign c5325 =  x290 &  x555 & ~x32;
assign c5327 =  x175 &  x479 & ~x14 & ~x98 & ~x113 & ~x587 & ~x615 & ~x757;
assign c5329 =  x491 &  x712;
assign c5331 =  x217 &  x554 & ~x5 & ~x23 & ~x62 & ~x141 & ~x165 & ~x222 & ~x279 & ~x726;
assign c5333 =  x620 & ~x41 & ~x221 & ~x289 & ~x304 & ~x309 & ~x316 & ~x336;
assign c5335 =  x436 &  x464 & ~x63 & ~x291;
assign c5337 =  x491 &  x628;
assign c5339 =  x435 &  x572;
assign c5341 =  x463 &  x628;
assign c5343 =  x563 &  x595;
assign c5345 =  x525 & ~x0 & ~x22 & ~x33 & ~x51 & ~x52 & ~x55 & ~x58 & ~x252 & ~x279 & ~x448 & ~x607 & ~x662 & ~x691 & ~x717 & ~x775 & ~x776;
assign c5347 =  x479 &  x593 & ~x336 & ~x364 & ~x780;
assign c5349 =  x322 & ~x29 & ~x282 & ~x461 & ~x774;
assign c5351 =  x682 & ~x156;
assign c5353 =  x129 & ~x31 & ~x72 & ~x225 & ~x572 & ~x780;
assign c5355 =  x151 & ~x0 & ~x22 & ~x224 & ~x378 & ~x447 & ~x545 & ~x643;
assign c5357 =  x205 & ~x0 & ~x1 & ~x28 & ~x38 & ~x54 & ~x56 & ~x85 & ~x101 & ~x223 & ~x323 & ~x351 & ~x352 & ~x560 & ~x671 & ~x673 & ~x685 & ~x702 & ~x704 & ~x734;
assign c5359 =  x407 & ~x551;
assign c5361 =  x306 & ~x482 & ~x483 & ~x509 & ~x533 & ~x560 & ~x593;
assign c5363 =  x410 & ~x34 & ~x165 & ~x223 & ~x468 & ~x654;
assign c5365 =  x491 &  x519 &  x547 & ~x8 & ~x26 & ~x35 & ~x777;
assign c5367 =  x230 &  x506 & ~x249;
assign c5369 =  x151 &  x243 & ~x705;
assign c5371 =  x547 &  x631 & ~x748;
assign c5373 =  x296 &  x521;
assign c5375 =  x260 &  x311 & ~x12 & ~x51 & ~x422 & ~x670 & ~x733;
assign c5377 =  x265 &  x395 & ~x42 & ~x700;
assign c5379 =  x410 & ~x378 & ~x467 & ~x645;
assign c5381 =  x553 & ~x639 & ~x663 & ~x746;
assign c5383 =  x178 & ~x8 & ~x29 & ~x51 & ~x56 & ~x280 & ~x348 & ~x350 & ~x629 & ~x643 & ~x655 & ~x704 & ~x729 & ~x753;
assign c5385 =  x175 &  x177 &  x660 & ~x680 & ~x704 & ~x731;
assign c5387 =  x50;
assign c5389 =  x204 &  x205 & ~x30 & ~x128 & ~x268 & ~x337 & ~x695 & ~x705 & ~x726 & ~x733 & ~x759;
assign c5391 =  x592 & ~x31 & ~x55 & ~x244 & ~x715 & ~x732 & ~x769;
assign c5393 =  x260 &  x310 & ~x643;
assign c5395 =  x710 & ~x482;
assign c5397 =  x570 & ~x35 & ~x111 & ~x704 & ~x705 & ~x724 & ~x730 & ~x732 & ~x746 & ~x755;
assign c5399 =  x624 & ~x27 & ~x127 & ~x336 & ~x634 & ~x662 & ~x759 & ~x777;
assign c5401 =  x136 & ~x60 & ~x89 & ~x362;
assign c5403 =  x517 & ~x66 & ~x156 & ~x494;
assign c5405 =  x193 & ~x279 & ~x498 & ~x560 & ~x588;
assign c5407 =  x710;
assign c5409 =  x461 & ~x2 & ~x128 & ~x156 & ~x467 & ~x554;
assign c5411 =  x582 & ~x58 & ~x61 & ~x81 & ~x87 & ~x112 & ~x167 & ~x171 & ~x199 & ~x489 & ~x515 & ~x532 & ~x669;
assign c5413 =  x205 & ~x46 & ~x261 & ~x670 & ~x726;
assign c5415 =  x90 &  x91 & ~x14 & ~x27 & ~x55 & ~x98 & ~x503;
assign c5417 =  x68 &  x69 & ~x485 & ~x486;
assign c5419 =  x261 &  x310;
assign c5421 =  x323 &  x521;
assign c5423 =  x378 & ~x0 & ~x69 & ~x409 & ~x503 & ~x699 & ~x749;
assign c5425 = ~x0 & ~x2 & ~x3 & ~x5 & ~x19 & ~x194 & ~x281 & ~x303 & ~x353 & ~x432 & ~x462 & ~x491 & ~x598 & ~x629 & ~x686;
assign c5427 =  x306 & ~x32 & ~x172 & ~x481 & ~x510 & ~x511 & ~x532 & ~x621;
assign c5429 =  x243 & ~x55 & ~x223 & ~x254 & ~x560 & ~x564 & ~x769;
assign c5431 =  x483 &  x517 & ~x776;
assign c5433 =  x517 & ~x19 & ~x82 & ~x164 & ~x551 & ~x639 & ~x659;
assign c5435 =  x582 & ~x227 & ~x280 & ~x309 & ~x363 & ~x579;
assign c5437 =  x136 & ~x332;
assign c5439 =  x593 & ~x1 & ~x55 & ~x70 & ~x280 & ~x343 & ~x659;
assign c5441 =  x119 &  x147 & ~x28 & ~x70 & ~x154 & ~x223 & ~x691 & ~x752;
assign c5443 =  x533 &  x621;
assign c5445 =  x380 &  x407 & ~x83 & ~x783;
assign c5447 =  x610 &  x611 & ~x4 & ~x5 & ~x22 & ~x111 & ~x112;
assign c5449 =  x422 & ~x1 & ~x31 & ~x84 & ~x138 & ~x172 & ~x196 & ~x198 & ~x281 & ~x358 & ~x672;
assign c5451 =  x498 & ~x133 & ~x165 & ~x554;
assign c5453 =  x137;
assign c5455 =  x626 & ~x85 & ~x99 & ~x101 & ~x732 & ~x735 & ~x740 & ~x754 & ~x764 & ~x774;
assign c5457 =  x352 & ~x0 & ~x757;
assign c5459 =  x158 & ~x6 & ~x288 & ~x491 & ~x573 & ~x600;
assign c5461 =  x407;
assign c5463 =  x462 &  x572 & ~x8 & ~x60 & ~x168 & ~x691 & ~x753;
assign c5465 =  x267 &  x491;
assign c5467 =  x322 & ~x41 & ~x42 & ~x72 & ~x223;
assign c5469 =  x181 &  x345 & ~x34 & ~x420 & ~x550 & ~x551 & ~x749;
assign c5471 =  x305 & ~x0 & ~x1 & ~x481 & ~x484 & ~x504 & ~x532 & ~x535 & ~x616;
assign c5473 =  x435 & ~x107 & ~x112 & ~x476 & ~x668 & ~x671;
assign c5475 =  x654 & ~x722 & ~x778;
assign c5477 =  x186 & ~x34 & ~x197 & ~x484 & ~x588 & ~x622 & ~x681 & ~x732 & ~x739 & ~x765 & ~x777;
assign c5479 =  x619 & ~x2 & ~x56 & ~x58 & ~x123 & ~x419 & ~x447 & ~x660 & ~x688;
assign c5481 =  x241 &  x269 &  x410;
assign c5483 =  x379 & ~x560;
assign c5485 =  x466 & ~x87 & ~x379 & ~x496 & ~x503 & ~x526 & ~x630 & ~x761;
assign c5487 =  x626 &  x627 & ~x770;
assign c5489 =  x175 &  x202 &  x506 & ~x29 & ~x83 & ~x107;
assign c5491 =  x294 &  x322 & ~x26 & ~x82 & ~x101 & ~x198 & ~x224 & ~x279 & ~x755 & ~x775;
assign c5493 =  x69 &  x123;
assign c5495 =  x260 &  x261 &  x286 &  x577 & ~x89 & ~x279 & ~x749;
assign c5497 =  x488 & ~x71 & ~x101 & ~x492 & ~x583 & ~x610 & ~x723;
assign c5499 =  x639 &  x640 &  x666;
assign c60 = ~x25 & ~x34 & ~x60 & ~x66 & ~x135 & ~x204 & ~x229 & ~x232 & ~x249 & ~x259 & ~x315 & ~x354 & ~x446 & ~x468 & ~x478 & ~x480 & ~x584 & ~x597 & ~x625 & ~x636 & ~x652 & ~x721;
assign c62 =  x295 &  x323 &  x379 &  x491 &  x547 &  x575 & ~x45 & ~x90 & ~x495;
assign c64 = ~x8 & ~x104 & ~x135 & ~x143 & ~x202 & ~x232 & ~x305 & ~x307 & ~x318 & ~x330 & ~x342 & ~x359 & ~x419 & ~x442 & ~x445 & ~x451 & ~x497 & ~x534 & ~x540 & ~x552 & ~x556 & ~x562 & ~x610 & ~x618 & ~x638 & ~x649 & ~x703 & ~x726 & ~x730 & ~x732 & ~x771 & ~x774;
assign c66 =  x72 &  x433 &  x522 &  x550;
assign c68 =  x577 &  x605 &  x633 & ~x8 & ~x53 & ~x250 & ~x278 & ~x479 & ~x527 & ~x539 & ~x556 & ~x587 & ~x594 & ~x610 & ~x781;
assign c610 =  x397 &  x552 & ~x168;
assign c612 =  x395 &  x515 &  x555;
assign c614 =  x463 &  x551 & ~x5 & ~x10 & ~x107 & ~x226 & ~x308 & ~x364 & ~x504 & ~x707 & ~x740;
assign c616 =  x515 &  x550 & ~x3 & ~x66 & ~x196 & ~x325;
assign c618 = ~x142 & ~x166 & ~x171 & ~x202 & ~x210 & ~x221 & ~x226 & ~x301 & ~x308 & ~x333 & ~x342 & ~x360 & ~x364 & ~x426 & ~x462 & ~x502 & ~x526 & ~x553 & ~x566 & ~x567 & ~x568 & ~x611 & ~x624 & ~x638 & ~x667 & ~x672 & ~x694 & ~x771;
assign c620 = ~x204 & ~x235 & ~x317 & ~x378 & ~x434;
assign c622 =  x394 &  x556;
assign c624 =  x378 &  x577 &  x604 & ~x353;
assign c626 =  x406 &  x434 &  x551 & ~x197 & ~x644 & ~x730;
assign c628 =  x550 & ~x2 & ~x9 & ~x55 & ~x66 & ~x143 & ~x278 & ~x281 & ~x309 & ~x560 & ~x624 & ~x643 & ~x697 & ~x702 & ~x703 & ~x738 & ~x759 & ~x765;
assign c630 =  x129 &  x130 &  x158 &  x578 & ~x1 & ~x113 & ~x138 & ~x363 & ~x504 & ~x589 & ~x731 & ~x755;
assign c632 =  x302 &  x550;
assign c634 =  x324 &  x352 &  x631 &  x659 & ~x8 & ~x106 & ~x226 & ~x285 & ~x514 & ~x539 & ~x637;
assign c636 =  x389;
assign c638 =  x518 &  x609;
assign c640 = ~x8 & ~x77 & ~x95 & ~x110 & ~x142 & ~x166 & ~x192 & ~x228 & ~x230 & ~x246 & ~x279 & ~x306 & ~x308 & ~x401 & ~x444 & ~x448 & ~x450 & ~x485 & ~x549 & ~x553 & ~x585 & ~x592 & ~x594 & ~x620 & ~x664 & ~x702 & ~x707 & ~x749 & ~x754;
assign c642 =  x472 &  x636;
assign c644 =  x406 &  x434 &  x523 &  x551 & ~x0 & ~x1 & ~x2 & ~x55 & ~x79 & ~x82 & ~x110 & ~x112 & ~x114 & ~x136 & ~x137 & ~x170 & ~x195 & ~x222 & ~x223 & ~x447 & ~x758 & ~x765;
assign c646 =  x211 & ~x19 & ~x35 & ~x46 & ~x83 & ~x132 & ~x147 & ~x161 & ~x244 & ~x278 & ~x368 & ~x425 & ~x446 & ~x485 & ~x539 & ~x542 & ~x552 & ~x560 & ~x580 & ~x583 & ~x608 & ~x615 & ~x638 & ~x663 & ~x669 & ~x670 & ~x703;
assign c648 =  x237 &  x266 &  x294 &  x321 &  x406 &  x433 & ~x36 & ~x55 & ~x195 & ~x723;
assign c650 =  x186 &  x214 & ~x0 & ~x8 & ~x34 & ~x36 & ~x38 & ~x80 & ~x145 & ~x163 & ~x250 & ~x257 & ~x277 & ~x281 & ~x341 & ~x396 & ~x449 & ~x556 & ~x610 & ~x614 & ~x638 & ~x640 & ~x651 & ~x695 & ~x697 & ~x702 & ~x728 & ~x749 & ~x777;
assign c652 = ~x19 & ~x24 & ~x111 & ~x164 & ~x170 & ~x220 & ~x228 & ~x313 & ~x317 & ~x387 & ~x401 & ~x539 & ~x561 & ~x596 & ~x603 & ~x608 & ~x612 & ~x733 & ~x755 & ~x771;
assign c654 =  x103 &  x550 &  x551;
assign c656 =  x350 &  x434 & ~x19 & ~x26 & ~x51 & ~x53 & ~x79 & ~x89 & ~x109 & ~x149 & ~x165 & ~x167 & ~x171 & ~x255 & ~x283 & ~x307 & ~x348 & ~x502 & ~x562 & ~x664 & ~x672 & ~x695 & ~x702 & ~x725 & ~x758 & ~x765 & ~x766;
assign c658 =  x424 &  x452 &  x463;
assign c660 =  x575 &  x664 & ~x35 & ~x167 & ~x254;
assign c662 =  x237 &  x238 &  x350 &  x378 &  x406 &  x490 & ~x198 & ~x279 & ~x306 & ~x474 & ~x534 & ~x583 & ~x666 & ~x730 & ~x735;
assign c664 =  x267 &  x463 &  x547 &  x631 & ~x104 & ~x144 & ~x553 & ~x666 & ~x729;
assign c666 = ~x188 & ~x208 & ~x232 & ~x293 & ~x357 & ~x582;
assign c668 =  x407 &  x424 & ~x84;
assign c670 = ~x0 & ~x77 & ~x89 & ~x106 & ~x164 & ~x193 & ~x230 & ~x273 & ~x281 & ~x318 & ~x342 & ~x429 & ~x436 & ~x492 & ~x513 & ~x560 & ~x563 & ~x610 & ~x717 & ~x763;
assign c672 =  x125 &  x238 &  x350 &  x574 &  x657 & ~x622;
assign c674 =  x424 &  x493 &  x535;
assign c676 =  x130 &  x514 & ~x678;
assign c678 =  x266 &  x684 & ~x168 & ~x219 & ~x249 & ~x341 & ~x364 & ~x422 & ~x506 & ~x512 & ~x513 & ~x568 & ~x591 & ~x621 & ~x634;
assign c680 =  x211 &  x267 &  x631 &  x659 &  x687 & ~x254 & ~x522;
assign c682 =  x266 &  x294 &  x378 &  x657 &  x684 & ~x568;
assign c684 =  x488 &  x554 &  x609 & ~x6 & ~x28 & ~x33 & ~x64;
assign c686 =  x237 &  x629 &  x683 & ~x605;
assign c688 =  x211 &  x295 &  x323 &  x463 &  x575 & ~x104 & ~x105 & ~x187 & ~x190 & ~x446 & ~x503 & ~x581 & ~x757;
assign c690 =  x422 &  x562 &  x618;
assign c692 =  x577 &  x633 &  x717 & ~x1 & ~x116 & ~x165 & ~x226 & ~x248 & ~x251 & ~x305 & ~x309 & ~x333 & ~x363 & ~x395 & ~x415 & ~x455 & ~x471 & ~x526 & ~x555 & ~x586 & ~x587 & ~x589 & ~x727 & ~x759;
assign c694 =  x515 & ~x8 & ~x279 & ~x354 & ~x453 & ~x469 & ~x622 & ~x625 & ~x676 & ~x679 & ~x708 & ~x717;
assign c696 =  x184 &  x212 &  x324 &  x408 &  x605 & ~x87 & ~x107 & ~x137 & ~x191 & ~x194 & ~x281 & ~x539 & ~x610;
assign c698 = ~x19 & ~x28 & ~x35 & ~x85 & ~x91 & ~x111 & ~x193 & ~x197 & ~x203 & ~x204 & ~x223 & ~x232 & ~x257 & ~x282 & ~x288 & ~x305 & ~x341 & ~x348 & ~x388 & ~x394 & ~x422 & ~x483 & ~x502 & ~x507 & ~x534 & ~x557 & ~x560 & ~x566 & ~x569 & ~x580 & ~x583 & ~x608 & ~x610 & ~x636 & ~x640 & ~x643 & ~x670 & ~x674 & ~x702 & ~x708 & ~x757;
assign c6100 = ~x79 & ~x181 & ~x195 & ~x207 & ~x248 & ~x253 & ~x349 & ~x446 & ~x501 & ~x585 & ~x597 & ~x653 & ~x701;
assign c6102 =  x11 &  x600;
assign c6104 = ~x8 & ~x19 & ~x55 & ~x102 & ~x163 & ~x190 & ~x198 & ~x317 & ~x539 & ~x552 & ~x566 & ~x588 & ~x633 & ~x661 & ~x696 & ~x738;
assign c6106 =  x102 &  x522 &  x523 &  x550 & ~x164 & ~x192;
assign c6108 =  x184 &  x268 &  x604 &  x605 & ~x54 & ~x169 & ~x365 & ~x639 & ~x699;
assign c6110 =  x238 &  x656 & ~x193 & ~x444 & ~x514 & ~x565 & ~x637 & ~x664 & ~x665;
assign c6112 =  x214 & ~x108 & ~x210 & ~x219 & ~x220 & ~x341 & ~x359 & ~x362 & ~x364 & ~x449 & ~x474 & ~x479 & ~x527 & ~x556 & ~x702 & ~x726;
assign c6114 =  x515 &  x551 &  x578 & ~x139 & ~x708 & ~x728 & ~x777;
assign c6116 =  x692 &  x720 & ~x94;
assign c6118 =  x479 &  x675;
assign c6120 =  x351 &  x576 &  x604 & ~x169 & ~x192 & ~x219 & ~x222 & ~x256 & ~x310 & ~x337 & ~x394 & ~x448 & ~x501 & ~x532 & ~x540 & ~x609 & ~x610;
assign c6122 =  x238 &  x323 &  x658 &  x686 & ~x542;
assign c6124 =  x212 &  x324 &  x579 & ~x53;
assign c6126 =  x514 &  x515 &  x551 &  x607;
assign c6128 =  x73 &  x74 & ~x197 & ~x210 & ~x225 & ~x421 & ~x590 & ~x646 & ~x672 & ~x677 & ~x679 & ~x764 & ~x778;
assign c6130 = ~x114 & ~x175 & ~x203 & ~x277 & ~x317 & ~x390 & ~x455 & ~x471 & ~x474 & ~x485 & ~x491 & ~x539 & ~x624 & ~x697 & ~x751;
assign c6132 =  x572 &  x626 & ~x107 & ~x248 & ~x437 & ~x511 & ~x550 & ~x610;
assign c6134 =  x213 &  x434 & ~x80 & ~x135 & ~x206 & ~x308 & ~x375 & ~x532 & ~x735 & ~x748 & ~x777;
assign c6136 =  x506 &  x562 &  x674;
assign c6138 =  x277 &  x527;
assign c6140 =  x324 &  x600 &  x662 & ~x169 & ~x614 & ~x642 & ~x673;
assign c6142 =  x575 &  x627 & ~x95;
assign c6144 =  x300 &  x576 & ~x38 & ~x79 & ~x137 & ~x285;
assign c6146 =  x237 &  x378 &  x602 &  x657 & ~x162 & ~x419 & ~x423 & ~x580 & ~x594 & ~x650;
assign c6148 = ~x113 & ~x144 & ~x202 & ~x222 & ~x276 & ~x285 & ~x286 & ~x291 & ~x304 & ~x316 & ~x317 & ~x333 & ~x367 & ~x492 & ~x520 & ~x525 & ~x526 & ~x565 & ~x580 & ~x610 & ~x640 & ~x698 & ~x730;
assign c6150 =  x157 & ~x0 & ~x19 & ~x83 & ~x88 & ~x137 & ~x140 & ~x166 & ~x255 & ~x279 & ~x283 & ~x332 & ~x335 & ~x342 & ~x388 & ~x392 & ~x446 & ~x499 & ~x513 & ~x526 & ~x530 & ~x532 & ~x555 & ~x563 & ~x589 & ~x591 & ~x621 & ~x644;
assign c6152 = ~x11 & ~x13 & ~x51 & ~x53 & ~x78 & ~x145 & ~x163 & ~x195 & ~x222 & ~x238 & ~x253 & ~x256 & ~x265 & ~x278 & ~x300 & ~x309 & ~x329 & ~x378 & ~x389 & ~x391 & ~x537 & ~x562 & ~x566 & ~x567 & ~x582 & ~x585 & ~x625 & ~x729 & ~x758 & ~x760 & ~x782;
assign c6154 =  x367 &  x462 &  x524;
assign c6156 =  x323 &  x324 &  x629 & ~x145 & ~x392 & ~x494 & ~x553;
assign c6158 =  x323 & ~x4 & ~x28 & ~x36 & ~x49 & ~x58 & ~x135 & ~x151 & ~x168 & ~x217 & ~x219 & ~x230 & ~x284 & ~x285 & ~x307 & ~x313 & ~x341 & ~x342 & ~x368 & ~x393 & ~x394 & ~x396 & ~x454 & ~x475 & ~x494 & ~x534 & ~x540 & ~x553 & ~x556 & ~x560 & ~x563 & ~x564 & ~x579 & ~x589 & ~x612 & ~x613 & ~x616 & ~x618 & ~x640 & ~x676 & ~x693 & ~x695 & ~x698 & ~x724;
assign c6160 = ~x7 & ~x21 & ~x139 & ~x281 & ~x306 & ~x335 & ~x358 & ~x401 & ~x420 & ~x443 & ~x453 & ~x457 & ~x458 & ~x466 & ~x492 & ~x496 & ~x510 & ~x526 & ~x532 & ~x539 & ~x608 & ~x615 & ~x637 & ~x638 & ~x669 & ~x702;
assign c6162 =  x211 &  x576 &  x689 & ~x539;
assign c6164 =  x562;
assign c6166 =  x209 &  x265 &  x294 &  x350 & ~x364 & ~x422 & ~x636 & ~x638;
assign c6168 =  x433 & ~x16 & ~x259 & ~x340 & ~x342 & ~x353 & ~x354 & ~x358 & ~x389 & ~x471 & ~x563 & ~x580 & ~x608 & ~x622 & ~x636 & ~x707;
assign c6170 =  x294 &  x517 &  x572 &  x599 &  x600 &  x626 &  x627 & ~x112 & ~x644 & ~x756 & ~x776 & ~x778;
assign c6172 =  x267 &  x631 &  x659 &  x686 & ~x77 & ~x245 & ~x277 & ~x313 & ~x415 & ~x417 & ~x421 & ~x477 & ~x537 & ~x550 & ~x607;
assign c6174 =  x294 &  x379 &  x406 &  x603 &  x631 &  x659 & ~x733 & ~x776;
assign c6176 =  x340 &  x368 &  x424 &  x462;
assign c6178 =  x528;
assign c6180 =  x546 &  x579 &  x606 &  x607 & ~x66 & ~x93;
assign c6182 =  x368 &  x424 &  x462;
assign c6184 =  x406 &  x554;
assign c6186 =  x73 &  x157 &  x270 & ~x114 & ~x255 & ~x280 & ~x781;
assign c6188 =  x577 &  x605 &  x633 &  x661 & ~x24 & ~x96 & ~x133 & ~x164 & ~x276 & ~x308 & ~x390 & ~x391 & ~x416 & ~x472 & ~x644 & ~x762;
assign c6190 =  x629 &  x662 & ~x80 & ~x252 & ~x487 & ~x515 & ~x532;
assign c6192 =  x211 &  x267 &  x295 &  x323 &  x379 &  x463 & ~x139 & ~x189 & ~x477 & ~x504 & ~x566 & ~x590 & ~x624 & ~x708 & ~x728 & ~x730;
assign c6194 =  x389;
assign c6196 =  x579 &  x606 &  x607 & ~x38 & ~x66 & ~x194 & ~x281 & ~x363 & ~x391 & ~x476 & ~x532 & ~x698 & ~x757 & ~x763;
assign c6198 =  x600 &  x627 &  x710 & ~x84 & ~x167 & ~x443 & ~x534 & ~x579 & ~x728;
assign c6200 =  x47 &  x662;
assign c6202 =  x393 &  x611;
assign c6204 =  x296 &  x576 &  x659 &  x687 & ~x470 & ~x666;
assign c6206 =  x605 &  x691 & ~x66 & ~x94;
assign c6208 =  x605 &  x633 & ~x1 & ~x26 & ~x29 & ~x64 & ~x95 & ~x104 & ~x137 & ~x162 & ~x163 & ~x164 & ~x192 & ~x227 & ~x228 & ~x250 & ~x253 & ~x256 & ~x276 & ~x333 & ~x338 & ~x341 & ~x359 & ~x360 & ~x368 & ~x415 & ~x417 & ~x449 & ~x451 & ~x475 & ~x476 & ~x539 & ~x555 & ~x581 & ~x589 & ~x618 & ~x642;
assign c6210 = ~x86 & ~x178 & ~x207 & ~x209 & ~x350 & ~x416 & ~x592;
assign c6212 =  x509;
assign c6214 =  x238 &  x294 &  x378 &  x406 &  x574 &  x630 & ~x0 & ~x28 & ~x199 & ~x482 & ~x521 & ~x538 & ~x777;
assign c6216 = ~x0 & ~x2 & ~x8 & ~x36 & ~x39 & ~x56 & ~x80 & ~x104 & ~x111 & ~x135 & ~x139 & ~x175 & ~x202 & ~x228 & ~x232 & ~x259 & ~x330 & ~x336 & ~x342 & ~x343 & ~x345 & ~x359 & ~x391 & ~x418 & ~x425 & ~x429 & ~x501 & ~x502 & ~x522 & ~x526 & ~x538 & ~x539 & ~x552 & ~x553 & ~x560 & ~x580 & ~x582 & ~x593 & ~x608 & ~x635 & ~x673 & ~x698 & ~x702 & ~x717 & ~x728 & ~x738 & ~x748 & ~x774 & ~x781;
assign c6218 =  x618;
assign c6220 =  x328 &  x575 &  x603 & ~x108 & ~x141 & ~x194 & ~x249 & ~x279 & ~x360 & ~x474 & ~x530 & ~x590;
assign c6222 = ~x0 & ~x2 & ~x19 & ~x32 & ~x35 & ~x82 & ~x95 & ~x104 & ~x108 & ~x135 & ~x143 & ~x146 & ~x167 & ~x169 & ~x195 & ~x226 & ~x229 & ~x288 & ~x339 & ~x365 & ~x368 & ~x383 & ~x415 & ~x417 & ~x446 & ~x507 & ~x526 & ~x527 & ~x538 & ~x539 & ~x552 & ~x580 & ~x587 & ~x594 & ~x598 & ~x609 & ~x610 & ~x620 & ~x644 & ~x646 & ~x667 & ~x694 & ~x706 & ~x726 & ~x733 & ~x745 & ~x757 & ~x774 & ~x777 & ~x783;
assign c6224 =  x157 &  x298 & ~x439;
assign c6226 =  x576 &  x604 &  x659 &  x687 & ~x53 & ~x77 & ~x105 & ~x135 & ~x187 & ~x188 & ~x221 & ~x246 & ~x279 & ~x365 & ~x426 & ~x441 & ~x511 & ~x529 & ~x580 & ~x582 & ~x589 & ~x640 & ~x642 & ~x751;
assign c6228 =  x571 &  x572 &  x597 & ~x113 & ~x618;
assign c6230 =  x675;
assign c6232 =  x544 &  x571 &  x609 & ~x96;
assign c6234 =  x184 &  x212 &  x576 &  x604 & ~x78 & ~x135 & ~x161 & ~x228 & ~x368 & ~x388 & ~x393 & ~x420 & ~x452 & ~x500 & ~x563 & ~x566 & ~x585 & ~x702 & ~x708;
assign c6236 = ~x3 & ~x42 & ~x208 & ~x249 & ~x265 & ~x376 & ~x526 & ~x536 & ~x625 & ~x642 & ~x651 & ~x652 & ~x758 & ~x771;
assign c6238 =  x324 &  x576 &  x604 &  x632 & ~x0 & ~x81 & ~x86 & ~x109 & ~x134 & ~x163 & ~x221 & ~x275 & ~x278 & ~x279 & ~x280 & ~x285 & ~x451 & ~x471 & ~x503 & ~x540 & ~x558 & ~x588 & ~x591 & ~x610 & ~x621 & ~x696 & ~x762 & ~x783;
assign c6240 =  x366;
assign c6242 =  x571 &  x572 &  x598 &  x623 & ~x2;
assign c6244 =  x656 & ~x12 & ~x39 & ~x77 & ~x112 & ~x139 & ~x332 & ~x419 & ~x497 & ~x513 & ~x570 & ~x638 & ~x666;
assign c6246 =  x547 &  x636 &  x637;
assign c6248 =  x506 &  x546 &  x562;
assign c6250 = ~x118 & ~x226 & ~x230 & ~x316 & ~x330 & ~x342 & ~x492 & ~x534 & ~x539 & ~x540 & ~x562 & ~x578 & ~x679 & ~x705 & ~x733 & ~x772;
assign c6252 =  x179 &  x187 &  x216 & ~x52 & ~x389 & ~x418 & ~x424 & ~x532;
assign c6254 =  x211 &  x212 &  x323 &  x604 & ~x92 & ~x104;
assign c6256 =  x302 & ~x326;
assign c6258 =  x213 &  x578 &  x606 & ~x139 & ~x229 & ~x421 & ~x652 & ~x653 & ~x706;
assign c6260 =  x546 &  x609 &  x637 & ~x142 & ~x777;
assign c6262 =  x184 &  x212 &  x324 &  x408 &  x632 & ~x364 & ~x451 & ~x540 & ~x619;
assign c6264 =  x352 &  x662 & ~x8 & ~x32 & ~x108 & ~x278 & ~x333 & ~x454 & ~x481;
assign c6266 =  x627 &  x628 &  x629 & ~x4 & ~x81 & ~x226 & ~x367 & ~x485 & ~x528 & ~x537;
assign c6268 =  x572 &  x609 &  x637 & ~x62 & ~x66;
assign c6270 =  x493 &  x609 & ~x7 & ~x39 & ~x83 & ~x122;
assign c6272 =  x236 &  x572 &  x598 &  x599 & ~x23 & ~x54 & ~x476 & ~x618;
assign c6274 = ~x181 & ~x190 & ~x210 & ~x273 & ~x286 & ~x350 & ~x397;
assign c6276 =  x378 &  x522 &  x550 & ~x135 & ~x326 & ~x354 & ~x705;
assign c6278 =  x237 &  x489 &  x598 &  x600 &  x628 & ~x441;
assign c6280 =  x212 & ~x0 & ~x19 & ~x79 & ~x84 & ~x131 & ~x160 & ~x167 & ~x186 & ~x194 & ~x217 & ~x229 & ~x279 & ~x282 & ~x304 & ~x309 & ~x315 & ~x338 & ~x363 & ~x366 & ~x391 & ~x392 & ~x397 & ~x416 & ~x499 & ~x508 & ~x526 & ~x533 & ~x539 & ~x553 & ~x561 & ~x582 & ~x594 & ~x613 & ~x623 & ~x638 & ~x650 & ~x721 & ~x725 & ~x782;
assign c6282 =  x101 &  x129 &  x578 & ~x111 & ~x252 & ~x428 & ~x587 & ~x595;
assign c6284 =  x462 &  x571 & ~x52 & ~x124 & ~x738;
assign c6286 = ~x261 & ~x455 & ~x491 & ~x497 & ~x529 & ~x540 & ~x622 & ~x647 & ~x771;
assign c6288 =  x506;
assign c6290 =  x598 &  x664 & ~x56 & ~x167 & ~x756;
assign c6292 =  x574 &  x663 &  x664 & ~x431;
assign c6294 =  x239 &  x324 &  x547 & ~x597 & ~x624;
assign c6296 =  x157 & ~x18 & ~x19 & ~x104 & ~x105 & ~x200 & ~x229 & ~x255 & ~x281 & ~x330 & ~x333 & ~x339 & ~x342 & ~x360 & ~x394 & ~x471 & ~x508 & ~x512 & ~x526 & ~x532 & ~x539 & ~x540 & ~x562 & ~x565 & ~x610 & ~x646 & ~x681 & ~x708 & ~x728 & ~x732 & ~x758 & ~x759 & ~x778 & ~x781;
assign c6298 =  x129 &  x551 &  x578 & ~x0 & ~x54 & ~x110 & ~x733;
assign c6300 =  x378 &  x655 &  x683 & ~x3 & ~x578 & ~x592 & ~x693 & ~x703 & ~x730;
assign c6302 =  x572 &  x597 &  x598 & ~x29 & ~x61 & ~x63 & ~x64 & ~x78 & ~x79 & ~x142 & ~x144 & ~x196 & ~x197 & ~x466 & ~x475 & ~x501 & ~x532 & ~x583 & ~x618 & ~x698 & ~x760;
assign c6304 =  x473 &  x609;
assign c6306 =  x606 & ~x8 & ~x35 & ~x63 & ~x95 & ~x135 & ~x228 & ~x278 & ~x338 & ~x367 & ~x554 & ~x590 & ~x697;
assign c6308 =  x294 &  x547 &  x633 & ~x111 & ~x113 & ~x220 & ~x364 & ~x450 & ~x640 & ~x765;
assign c6310 =  x415 &  x565 & ~x777;
assign c6312 =  x266 &  x574 &  x629 &  x655 &  x657;
assign c6314 =  x463 &  x497 &  x525 & ~x138 & ~x779;
assign c6316 =  x515 &  x550 & ~x113 & ~x222 & ~x250 & ~x475 & ~x503 & ~x558 & ~x560 & ~x750;
assign c6318 = ~x137 & ~x143 & ~x198 & ~x378 & ~x379 & ~x401 & ~x470 & ~x513 & ~x534 & ~x557 & ~x568 & ~x590 & ~x609 & ~x610 & ~x642 & ~x665 & ~x674 & ~x676 & ~x694 & ~x753 & ~x757;
assign c6320 =  x214 &  x242 & ~x32 & ~x82 & ~x163 & ~x188 & ~x230 & ~x274 & ~x368 & ~x391 & ~x442 & ~x469 & ~x474 & ~x534 & ~x620 & ~x646 & ~x735;
assign c6322 =  x655 &  x683 &  x710 & ~x482 & ~x521 & ~x580;
assign c6324 =  x514 &  x541 &  x578 & ~x89 & ~x90 & ~x112;
assign c6326 =  x294 &  x574 & ~x363 & ~x464 & ~x748;
assign c6328 = ~x58 & ~x112 & ~x115 & ~x181 & ~x198 & ~x199 & ~x209 & ~x210 & ~x237 & ~x283 & ~x331 & ~x341 & ~x471 & ~x476 & ~x582 & ~x583 & ~x593 & ~x650 & ~x652 & ~x729 & ~x770;
assign c6330 =  x205 &  x237 & ~x3 & ~x7 & ~x46 & ~x54 & ~x55 & ~x110 & ~x115 & ~x139 & ~x168 & ~x201 & ~x226 & ~x251 & ~x278 & ~x308 & ~x331 & ~x363 & ~x364 & ~x415 & ~x534 & ~x589 & ~x595 & ~x610 & ~x611 & ~x621 & ~x646 & ~x676 & ~x699 & ~x733 & ~x781;
assign c6332 =  x238 &  x266 &  x294 &  x378 &  x434 &  x462 & ~x8 & ~x106 & ~x145 & ~x313 & ~x359 & ~x390 & ~x532 & ~x538 & ~x540 & ~x580 & ~x610 & ~x624;
assign c6334 = ~x58 & ~x163 & ~x181 & ~x266 & ~x323 & ~x534 & ~x568 & ~x726 & ~x781;
assign c6336 =  x294 &  x490 &  x574 & ~x436;
assign c6338 =  x212 &  x631 &  x686 & ~x60 & ~x160 & ~x200 & ~x283 & ~x302 & ~x363 & ~x368 & ~x448 & ~x468 & ~x511 & ~x556 & ~x583 & ~x608 & ~x609 & ~x617 & ~x753;
assign c6340 =  x189 &  x294 &  x378 &  x406;
assign c6342 = ~x39 & ~x81 & ~x135 & ~x181 & ~x208 & ~x209 & ~x210 & ~x228 & ~x277 & ~x312 & ~x363 & ~x388 & ~x389 & ~x396 & ~x563 & ~x675 & ~x762;
assign c6344 =  x238 &  x266 &  x406 &  x600 &  x628 & ~x514;
assign c6346 =  x268 &  x576 &  x604 &  x632 & ~x23 & ~x45 & ~x115 & ~x134 & ~x198 & ~x228 & ~x255 & ~x389;
assign c6348 =  x546 &  x609;
assign c6350 =  x241 &  x297 &  x631 & ~x111 & ~x341 & ~x396 & ~x423 & ~x446 & ~x518 & ~x529 & ~x558 & ~x566 & ~x641;
assign c6352 =  x600 &  x637 & ~x33 & ~x111 & ~x252;
assign c6354 = ~x0 & ~x26 & ~x141 & ~x218 & ~x237 & ~x258 & ~x293 & ~x360 & ~x415 & ~x447 & ~x454 & ~x528 & ~x538 & ~x563 & ~x616 & ~x624 & ~x638 & ~x639 & ~x669 & ~x704 & ~x746 & ~x756;
assign c6356 =  x321 &  x349 &  x683 &  x709 & ~x475 & ~x532 & ~x730 & ~x761;
assign c6358 =  x214 &  x550 &  x578 & ~x105 & ~x106 & ~x258 & ~x556 & ~x705;
assign c6360 =  x449;
assign c6362 = ~x54 & ~x62 & ~x77 & ~x247 & ~x276 & ~x277 & ~x290 & ~x308 & ~x345 & ~x363 & ~x370 & ~x471 & ~x554 & ~x555 & ~x623 & ~x625 & ~x639 & ~x648 & ~x677 & ~x688 & ~x748 & ~x772 & ~x777;
assign c6364 = ~x23 & ~x39 & ~x56 & ~x66 & ~x87 & ~x93 & ~x114 & ~x196 & ~x226 & ~x279 & ~x284 & ~x307 & ~x308 & ~x335 & ~x364 & ~x386 & ~x458 & ~x489 & ~x526 & ~x550 & ~x552 & ~x553 & ~x567 & ~x610 & ~x654;
assign c6366 =  x267 &  x378 &  x434 &  x462 &  x605 & ~x109 & ~x250 & ~x251 & ~x354 & ~x561;
assign c6368 =  x212 &  x324 &  x604 & ~x104 & ~x161 & ~x199 & ~x340 & ~x394 & ~x481 & ~x503 & ~x610 & ~x703;
assign c6370 =  x129 &  x157 &  x241 &  x577 & ~x77 & ~x167 & ~x245 & ~x394 & ~x446 & ~x588 & ~x611 & ~x759;
assign c6372 =  x237 &  x657 &  x683 & ~x577;
assign c6374 =  x600 &  x626 &  x627 &  x628 & ~x53 & ~x60 & ~x226 & ~x413 & ~x495 & ~x532 & ~x566 & ~x617 & ~x730;
assign c6376 =  x131 &  x132 &  x551 & ~x8;
assign c6378 =  x602 &  x630 &  x657 & ~x7 & ~x35 & ~x139 & ~x526 & ~x532 & ~x537 & ~x552 & ~x563 & ~x578 & ~x580 & ~x610 & ~x636;
assign c6380 =  x129 &  x522 & ~x55 & ~x77 & ~x109 & ~x111 & ~x197 & ~x227 & ~x283 & ~x504 & ~x560 & ~x622 & ~x709 & ~x736 & ~x756 & ~x777;
assign c6382 =  x233 &  x234 &  x631 & ~x0 & ~x168 & ~x196 & ~x226 & ~x252 & ~x276 & ~x277 & ~x284 & ~x303 & ~x414 & ~x425 & ~x449 & ~x450 & ~x610 & ~x671 & ~x676;
assign c6384 =  x434 &  x550 & ~x196 & ~x326 & ~x335 & ~x664 & ~x758;
assign c6386 =  x574 &  x664 &  x692;
assign c6388 =  x211 &  x267 &  x295 &  x323 &  x379 &  x659 & ~x102 & ~x143 & ~x252 & ~x334 & ~x337 & ~x636 & ~x647 & ~x726 & ~x781;
assign c6390 =  x156 &  x297 & ~x162 & ~x284 & ~x309 & ~x370 & ~x427 & ~x482 & ~x484 & ~x495 & ~x524 & ~x539 & ~x565 & ~x580 & ~x728;
assign c6392 =  x546 &  x636 & ~x29 & ~x57 & ~x251 & ~x671 & ~x767;
assign c6394 =  x321 &  x405 &  x433 &  x544 & ~x24 & ~x436;
assign c6396 =  x551 &  x568 &  x578 & ~x35 & ~x120 & ~x759;
assign c6398 =  x211 &  x323 &  x547 &  x575 & ~x185 & ~x482;
assign c6400 =  x179 &  x205 &  x238 &  x266 &  x294;
assign c6402 =  x628 &  x629 &  x655 &  x656 & ~x88 & ~x169 & ~x305 & ~x336 & ~x484 & ~x526 & ~x528 & ~x537 & ~x540 & ~x552 & ~x584 & ~x590 & ~x670 & ~x722;
assign c6404 =  x294 &  x574 & ~x87 & ~x313 & ~x492;
assign c6406 =  x546 &  x577 &  x636 &  x637;
assign c6408 =  x211 &  x267 &  x295 & ~x129 & ~x201 & ~x219 & ~x285 & ~x315 & ~x330 & ~x536 & ~x539 & ~x665 & ~x733 & ~x735;
assign c6410 =  x208 &  x270 & ~x8 & ~x29 & ~x32 & ~x108 & ~x136 & ~x137 & ~x163 & ~x251 & ~x282 & ~x313 & ~x368 & ~x394 & ~x423 & ~x473 & ~x587 & ~x647 & ~x667 & ~x702 & ~x726 & ~x731 & ~x759;
assign c6412 =  x324 &  x577 &  x605 &  x633 &  x688 & ~x85 & ~x196 & ~x220 & ~x306 & ~x339 & ~x415 & ~x444 & ~x471 & ~x480 & ~x676;
assign c6414 =  x691 & ~x95 & ~x139 & ~x276 & ~x458 & ~x532;
assign c6416 =  x562 &  x618 &  x646;
assign c6418 =  x295 &  x631 &  x687 & ~x0 & ~x19 & ~x54 & ~x115 & ~x163 & ~x167 & ~x199 & ~x246 & ~x363 & ~x368 & ~x394 & ~x398 & ~x419 & ~x498 & ~x500 & ~x503 & ~x509 & ~x539 & ~x552 & ~x564 & ~x580 & ~x590 & ~x759;
assign c6420 =  x491 &  x580 & ~x82 & ~x92 & ~x168 & ~x198 & ~x765;
assign c6422 =  x379 &  x658 &  x686 &  x713 & ~x0 & ~x77 & ~x106 & ~x117 & ~x246 & ~x278 & ~x361 & ~x501 & ~x507 & ~x510 & ~x527;
assign c6424 =  x491 &  x524 &  x552 &  x580;
assign c6426 =  x270 &  x575 & ~x57 & ~x79 & ~x109 & ~x170 & ~x224 & ~x246 & ~x286 & ~x336 & ~x392 & ~x413 & ~x532 & ~x557 & ~x643 & ~x646 & ~x671 & ~x676 & ~x736 & ~x782;
assign c6428 =  x367 &  x582;
assign c6430 =  x458 &  x551 & ~x27 & ~x139 & ~x298 & ~x760;
assign c6432 = ~x25 & ~x82 & ~x143 & ~x290 & ~x348 & ~x363 & ~x401 & ~x403 & ~x409 & ~x437 & ~x444 & ~x525 & ~x594 & ~x624 & ~x638 & ~x694 & ~x775;
assign c6434 = ~x148 & ~x181 & ~x208 & ~x238 & ~x263 & ~x379 & ~x504 & ~x589 & ~x681;
assign c6436 =  x238 &  x656 &  x683 &  x711 & ~x542 & ~x567;
assign c6438 =  x377 &  x653 &  x657;
assign c6440 = ~x11 & ~x19 & ~x21 & ~x33 & ~x49 & ~x51 & ~x55 & ~x80 & ~x92 & ~x102 & ~x110 & ~x119 & ~x139 & ~x159 & ~x168 & ~x196 & ~x197 & ~x200 & ~x226 & ~x228 & ~x229 & ~x231 & ~x249 & ~x275 & ~x278 & ~x281 & ~x307 & ~x310 & ~x316 & ~x341 & ~x343 & ~x358 & ~x363 & ~x368 & ~x413 & ~x420 & ~x429 & ~x443 & ~x479 & ~x482 & ~x484 & ~x501 & ~x502 & ~x504 & ~x507 & ~x511 & ~x527 & ~x529 & ~x531 & ~x534 & ~x562 & ~x567 & ~x569 & ~x580 & ~x591 & ~x593 & ~x594 & ~x610 & ~x611 & ~x618 & ~x625 & ~x642 & ~x644 & ~x645 & ~x673 & ~x677 & ~x735 & ~x778;
assign c6442 = ~x95 & ~x131 & ~x190 & ~x342 & ~x419 & ~x426 & ~x486 & ~x495 & ~x522 & ~x565 & ~x591 & ~x593 & ~x650 & ~x654 & ~x676 & ~x748;
assign c6444 =  x607 &  x693;
assign c6446 = ~x119 & ~x168 & ~x390 & ~x436 & ~x485 & ~x491 & ~x566 & ~x593 & ~x609 & ~x612 & ~x661;
assign c6448 =  x238 &  x323 &  x378 &  x379 &  x631 &  x659 &  x687 & ~x141 & ~x422 & ~x650;
assign c6450 = ~x81 & ~x201 & ~x206 & ~x208 & ~x210 & ~x317 & ~x324 & ~x532 & ~x782;
assign c6452 =  x295 &  x323 &  x547 &  x603 & ~x163 & ~x186 & ~x365 & ~x552 & ~x592;
assign c6454 =  x130 &  x298 &  x635;
assign c6456 = ~x2 & ~x39 & ~x79 & ~x87 & ~x104 & ~x133 & ~x176 & ~x196 & ~x201 & ~x228 & ~x251 & ~x279 & ~x287 & ~x308 & ~x340 & ~x360 & ~x401 & ~x447 & ~x501 & ~x513 & ~x528 & ~x532 & ~x567 & ~x569 & ~x590 & ~x592 & ~x625 & ~x646 & ~x697 & ~x716 & ~x733 & ~x749 & ~x770;
assign c6458 = ~x85 & ~x200 & ~x260 & ~x290 & ~x318 & ~x339 & ~x357 & ~x388 & ~x472 & ~x474 & ~x535 & ~x622 & ~x658 & ~x774;
assign c6460 =  x213 &  x631 & ~x165 & ~x255 & ~x312 & ~x334 & ~x340 & ~x364 & ~x388 & ~x455 & ~x487 & ~x502 & ~x533 & ~x610 & ~x780;
assign c6462 =  x602 &  x628 &  x654 &  x657 & ~x2 & ~x170;
assign c6464 =  x267 &  x604 & ~x167 & ~x227 & ~x245 & ~x284 & ~x422 & ~x512 & ~x553 & ~x557 & ~x723;
assign c6466 = ~x0 & ~x29 & ~x84 & ~x108 & ~x134 & ~x137 & ~x142 & ~x191 & ~x201 & ~x202 & ~x222 & ~x224 & ~x227 & ~x245 & ~x250 & ~x303 & ~x304 & ~x311 & ~x360 & ~x363 & ~x367 & ~x372 & ~x389 & ~x408 & ~x418 & ~x444 & ~x478 & ~x482 & ~x497 & ~x502 & ~x529 & ~x552 & ~x553 & ~x560 & ~x565 & ~x581 & ~x633 & ~x664 & ~x679 & ~x688 & ~x696 & ~x701 & ~x706 & ~x719 & ~x735 & ~x743 & ~x755 & ~x759 & ~x777;
assign c6468 =  x540;
assign c6470 =  x211 &  x379 &  x657 &  x712 & ~x257 & ~x608;
assign c6472 =  x433 &  x656 &  x683 &  x711 & ~x0 & ~x394 & ~x514 & ~x607 & ~x608 & ~x636;
assign c6474 =  x211 &  x239 &  x295 &  x379 & ~x21 & ~x58 & ~x75 & ~x108 & ~x111 & ~x226 & ~x364 & ~x391 & ~x529 & ~x537 & ~x556 & ~x568 & ~x596 & ~x616 & ~x642 & ~x646 & ~x650 & ~x665 & ~x671 & ~x679 & ~x697 & ~x699 & ~x704 & ~x752 & ~x753;
assign c6476 =  x549 & ~x39 & ~x79 & ~x87 & ~x139 & ~x144 & ~x162 & ~x191 & ~x210 & ~x248 & ~x275 & ~x282 & ~x395 & ~x471 & ~x527 & ~x610 & ~x613 & ~x643 & ~x674 & ~x759;
assign c6478 =  x499 &  x619;
assign c6480 =  x361 &  x493;
assign c6482 =  x368 &  x497 &  x525 & ~x112 & ~x139;
assign c6484 =  x434 &  x498 &  x578;
assign c6486 =  x571 &  x572 &  x635 &  x636 & ~x767;
assign c6488 =  x568 &  x577 & ~x353;
assign c6490 =  x579 &  x580 &  x607 & ~x8 & ~x52 & ~x54 & ~x79 & ~x96 & ~x167 & ~x169 & ~x195 & ~x225 & ~x728 & ~x781;
assign c6492 =  x544 &  x572 &  x600 &  x627 & ~x342 & ~x362 & ~x458 & ~x553;
assign c6494 =  x434 &  x553 & ~x110 & ~x354;
assign c6496 = ~x8 & ~x14 & ~x140 & ~x167 & ~x301 & ~x468 & ~x492 & ~x526 & ~x580 & ~x583 & ~x607 & ~x636 & ~x667 & ~x677 & ~x707 & ~x761 & ~x781;
assign c6498 = ~x134 & ~x151 & ~x186 & ~x213 & ~x317 & ~x542 & ~x595 & ~x636 & ~x688 & ~x709;
assign c61 =  x347 & ~x234 & ~x256 & ~x269;
assign c63 =  x439 &  x466 &  x467 & ~x375 & ~x406 & ~x432;
assign c65 = ~x403 & ~x460 & ~x488 & ~x517 & ~x546 & ~x627 & ~x656 & ~x684 & ~x717;
assign c67 =  x356 &  x360;
assign c69 =  x465 &  x743 & ~x146 & ~x298 & ~x303 & ~x399 & ~x457 & ~x525;
assign c611 =  x741 & ~x75 & ~x112 & ~x143 & ~x148 & ~x246 & ~x247 & ~x248 & ~x285 & ~x302 & ~x357 & ~x416 & ~x419 & ~x527 & ~x589 & ~x630 & ~x673 & ~x752;
assign c613 =  x359 &  x390 & ~x12 & ~x585;
assign c617 =  x345 &  x372 &  x400 & ~x708 & ~x771;
assign c619 =  x120 &  x232 &  x260;
assign c621 =  x67 &  x96 &  x317 & ~x75 & ~x479 & ~x725;
assign c623 =  x288 &  x314 & ~x160 & ~x539;
assign c625 =  x307;
assign c627 =  x123 &  x151 & ~x212 & ~x240 & ~x285;
assign c629 = ~x74 & ~x128 & ~x156 & ~x183 & ~x184 & ~x211 & ~x214 & ~x533 & ~x724;
assign c631 =  x356 &  x359;
assign c633 = ~x374 & ~x418 & ~x429 & ~x460 & ~x517 & ~x661;
assign c635 =  x95 &  x152 &  x290;
assign c637 =  x124 &  x127 &  x154 &  x291 & ~x160;
assign c639 =  x33;
assign c641 =  x138;
assign c643 =  x320 &  x432 & ~x39 & ~x298 & ~x333;
assign c645 =  x67 &  x96 &  x124 & ~x404;
assign c647 =  x359 & ~x465 & ~x522;
assign c649 =  x69 &  x126 & ~x460;
assign c651 =  x276;
assign c653 =  x166;
assign c655 =  x127 &  x485 &  x717 & ~x204;
assign c657 =  x403 &  x431 & ~x87 & ~x298 & ~x382 & ~x655;
assign c659 =  x320 & ~x19 & ~x134 & ~x185 & ~x191 & ~x268 & ~x269 & ~x335 & ~x422;
assign c661 =  x313 & ~x98 & ~x125 & ~x182;
assign c663 = ~x321 & ~x543;
assign c665 =  x432 & ~x70 & ~x299 & ~x318 & ~x442;
assign c667 = ~x33 & ~x47 & ~x76 & ~x240 & ~x241 & ~x242 & ~x249 & ~x253 & ~x267 & ~x269 & ~x270 & ~x272 & ~x284 & ~x285 & ~x287 & ~x297 & ~x476 & ~x538 & ~x586 & ~x638 & ~x699;
assign c669 =  x40 &  x466 & ~x48 & ~x160 & ~x188 & ~x190;
assign c671 =  x330 &  x474;
assign c673 = ~x99 & ~x126 & ~x156 & ~x269;
assign c675 =  x742 &  x743 &  x771 & ~x55 & ~x63 & ~x145 & ~x203 & ~x220 & ~x372 & ~x455 & ~x524;
assign c677 =  x109;
assign c679 = ~x103 & ~x114 & ~x162 & ~x183 & ~x184 & ~x215 & ~x241 & ~x242 & ~x421 & ~x482 & ~x678 & ~x733;
assign c681 =  x650 & ~x574;
assign c683 =  x376 &  x432 & ~x32 & ~x96 & ~x111 & ~x197 & ~x336 & ~x392 & ~x413 & ~x428 & ~x497 & ~x525 & ~x526 & ~x535 & ~x672 & ~x731 & ~x734 & ~x757;
assign c685 =  x64 &  x94;
assign c687 = ~x46 & ~x70 & ~x128 & ~x130 & ~x156 & ~x715 & ~x740;
assign c689 =  x494 & ~x331 & ~x404 & ~x433 & ~x692;
assign c691 =  x67 &  x151 & ~x320;
assign c693 =  x89;
assign c695 =  x370 & ~x161 & ~x639 & ~x715;
assign c697 =  x258 & ~x126 & ~x514;
assign c699 = ~x128 & ~x129 & ~x156 & ~x211 & ~x213 & ~x267 & ~x467 & ~x676;
assign c6101 =  x432 & ~x125 & ~x355 & ~x383 & ~x443 & ~x666 & ~x678;
assign c6103 =  x402 &  x430 & ~x227 & ~x270 & ~x288 & ~x343 & ~x611 & ~x706 & ~x733 & ~x763;
assign c6105 =  x41 &  x42 &  x71 &  x125 & ~x3 & ~x90 & ~x102 & ~x391 & ~x396 & ~x445 & ~x760;
assign c6107 =  x444 & ~x378 & ~x545;
assign c6109 =  x41 & ~x45 & ~x49 & ~x102 & ~x104 & ~x146 & ~x546 & ~x662;
assign c6111 = ~x67 & ~x516 & ~x517 & ~x545 & ~x628 & ~x629 & ~x686;
assign c6113 = ~x45 & ~x99 & ~x126 & ~x156 & ~x320;
assign c6115 =  x427 & ~x627 & ~x740 & ~x741;
assign c6117 = ~x461 & ~x548 & ~x576 & ~x601;
assign c6119 =  x495 & ~x433 & ~x435 & ~x462 & ~x476;
assign c6121 =  x278 & ~x474;
assign c6123 =  x161 & ~x125 & ~x720;
assign c6125 =  x249 & ~x473;
assign c6127 = ~x18 & ~x41 & ~x69 & ~x99 & ~x127 & ~x128 & ~x156 & ~x184;
assign c6129 =  x741 & ~x63 & ~x341 & ~x449 & ~x686;
assign c6131 =  x95 &  x123 &  x207;
assign c6133 =  x278 & ~x467 & ~x553;
assign c6135 =  x714 &  x772 & ~x86 & ~x249 & ~x275 & ~x330 & ~x440 & ~x554 & ~x646;
assign c6137 =  x133 &  x175 & ~x125 & ~x662;
assign c6139 =  x595 & ~x160 & ~x299 & ~x333 & ~x335;
assign c6141 =  x362 & ~x610;
assign c6143 =  x127 &  x182 & ~x111 & ~x193 & ~x225 & ~x241 & ~x268 & ~x269 & ~x298 & ~x304 & ~x305 & ~x324 & ~x535 & ~x559 & ~x562 & ~x644 & ~x724 & ~x781;
assign c6145 =  x201 & ~x41 & ~x98;
assign c6147 = ~x102 & ~x126 & ~x156 & ~x686 & ~x713;
assign c6149 =  x434 &  x520 & ~x41 & ~x411 & ~x666 & ~x732 & ~x745;
assign c6151 =  x111;
assign c6153 = ~x38 & ~x49 & ~x71 & ~x99 & ~x152 & ~x153 & ~x683 & ~x690;
assign c6155 = ~x462 & ~x545 & ~x546 & ~x714;
assign c6157 =  x66 &  x95 & ~x25 & ~x52 & ~x128 & ~x132 & ~x133;
assign c6159 =  x411 & ~x601;
assign c6161 =  x347 & ~x161 & ~x204 & ~x342 & ~x498 & ~x521 & ~x585;
assign c6163 =  x139;
assign c6165 =  x67 &  x124 & ~x320;
assign c6167 =  x741 & ~x162 & ~x516 & ~x661 & ~x726;
assign c6169 = ~x70 & ~x125 & ~x152 & ~x236 & ~x355 & ~x690;
assign c6171 =  x466 &  x769;
assign c6173 =  x218 &  x245 &  x246 & ~x745;
assign c6175 =  x610 & ~x71;
assign c6177 =  x154 &  x715 &  x716 &  x717 & ~x358 & ~x423 & ~x503 & ~x725 & ~x783;
assign c6179 = ~x322 & ~x377 & ~x404 & ~x406 & ~x546;
assign c6181 =  x467 &  x468 & ~x407;
assign c6183 =  x109;
assign c6185 =  x66 &  x95 &  x124 &  x262 &  x290;
assign c6187 = ~x403 & ~x404 & ~x405 & ~x435;
assign c6189 =  x127 &  x403 &  x715 & ~x579 & ~x765;
assign c6191 =  x172 & ~x71 & ~x98;
assign c6193 =  x373 & ~x39 & ~x541 & ~x740 & ~x741;
assign c6195 =  x716 &  x717 &  x747 & ~x133 & ~x161 & ~x246 & ~x395 & ~x610;
assign c6197 =  x741 &  x742 & ~x19 & ~x21 & ~x36 & ~x81 & ~x82 & ~x112 & ~x141 & ~x146 & ~x165 & ~x201 & ~x206 & ~x257 & ~x299 & ~x301 & ~x335 & ~x367 & ~x385 & ~x411 & ~x414 & ~x423 & ~x501 & ~x508 & ~x530 & ~x534 & ~x556 & ~x558 & ~x559 & ~x637 & ~x642 & ~x645 & ~x647 & ~x669 & ~x674 & ~x701 & ~x704 & ~x724 & ~x727 & ~x728;
assign c6199 =  x99 &  x431 &  x746;
assign c6201 =  x175 & ~x99 & ~x155 & ~x236;
assign c6203 = ~x23 & ~x65 & ~x392 & ~x516 & ~x545 & ~x572 & ~x574 & ~x629 & ~x656 & ~x686;
assign c6205 =  x740 &  x741 &  x742 & ~x338 & ~x365 & ~x395 & ~x534 & ~x620 & ~x637 & ~x658;
assign c6207 =  x97 &  x124 &  x345 & ~x232;
assign c6209 =  x64 &  x526 & ~x73;
assign c6211 = ~x26 & ~x115 & ~x207 & ~x223 & ~x234 & ~x516 & ~x628 & ~x629;
assign c6213 =  x326 &  x439 & ~x404;
assign c6215 =  x68 &  x126 &  x744 & ~x160 & ~x190 & ~x423;
assign c6217 =  x118 & ~x99;
assign c6219 =  x382 &  x409 &  x410 & ~x34 & ~x64 & ~x65 & ~x84 & ~x173 & ~x202 & ~x229 & ~x248 & ~x304 & ~x335;
assign c6221 =  x127 &  x290 & ~x78 & ~x148 & ~x230 & ~x231 & ~x308 & ~x563 & ~x615 & ~x669 & ~x722 & ~x754;
assign c6223 =  x149 & ~x99;
assign c6225 = ~x211 & ~x215 & ~x241 & ~x252 & ~x268 & ~x269 & ~x298 & ~x416;
assign c6227 = ~x403 & ~x404 & ~x460 & ~x515 & ~x546 & ~x573 & ~x742;
assign c6229 =  x342 & ~x41 & ~x43 & ~x738 & ~x742;
assign c6231 = ~x403 & ~x461 & ~x546 & ~x628 & ~x657;
assign c6233 =  x210 &  x516 &  x772 & ~x358 & ~x577 & ~x583;
assign c6235 =  x125 &  x319 & ~x16 & ~x44 & ~x76 & ~x625 & ~x698;
assign c6237 =  x154 &  x438 & ~x107 & ~x275 & ~x433;
assign c6239 =  x439 & ~x402 & ~x404 & ~x434;
assign c6241 =  x319 &  x371 & ~x597 & ~x653;
assign c6243 =  x391 & ~x610;
assign c6245 =  x183 &  x403 &  x431 & ~x82 & ~x357 & ~x399 & ~x449;
assign c6247 =  x437 &  x466 &  x494 & ~x8 & ~x330 & ~x460 & ~x502;
assign c6249 =  x166;
assign c6251 =  x740 &  x741 & ~x54 & ~x134 & ~x140 & ~x143 & ~x147 & ~x174 & ~x175 & ~x222 & ~x277 & ~x306 & ~x369 & ~x390 & ~x471 & ~x472 & ~x506 & ~x508 & ~x527 & ~x563 & ~x576 & ~x591 & ~x610 & ~x613 & ~x644 & ~x697;
assign c6253 =  x356 & ~x405 & ~x463;
assign c6255 =  x353 &  x439 &  x467 & ~x451;
assign c6257 =  x181 &  x376 &  x403 & ~x217 & ~x289 & ~x298;
assign c6259 =  x296 & ~x461 & ~x528 & ~x658;
assign c6261 =  x596 & ~x320 & ~x451;
assign c6263 =  x247 &  x272;
assign c6265 =  x95 &  x96 &  x316;
assign c6267 =  x399 &  x428;
assign c6269 =  x120 & ~x349;
assign c6271 = ~x404 & ~x435 & ~x740;
assign c6273 =  x741 &  x743 &  x772 & ~x289 & ~x333;
assign c6275 =  x402 &  x430 &  x485 & ~x395 & ~x496;
assign c6277 = ~x70 & ~x152 & ~x573 & ~x685 & ~x768;
assign c6279 =  x373 &  x401 &  x429 & ~x41;
assign c6281 =  x344 &  x370 & ~x496 & ~x624;
assign c6283 =  x99 &  x716 &  x744 &  x746 & ~x60 & ~x76 & ~x309 & ~x331 & ~x360 & ~x447 & ~x505 & ~x698;
assign c6285 =  x345 &  x483 & ~x229 & ~x231;
assign c6287 =  x43 &  x100 &  x743 & ~x298 & ~x299 & ~x330 & ~x562;
assign c6289 =  x403 & ~x41 & ~x673 & ~x683 & ~x709;
assign c6291 =  x382 &  x596;
assign c6293 = ~x12 & ~x32 & ~x50 & ~x119 & ~x220 & ~x268 & ~x269 & ~x270 & ~x272 & ~x298 & ~x737 & ~x738;
assign c6295 = ~x74 & ~x128 & ~x183 & ~x212 & ~x397 & ~x467 & ~x746;
assign c6297 =  x430 & ~x41 & ~x70 & ~x713 & ~x740;
assign c6299 =  x403 &  x431 &  x573 & ~x54 & ~x59 & ~x109 & ~x243 & ~x249 & ~x305 & ~x340 & ~x365 & ~x420 & ~x444 & ~x617 & ~x706 & ~x736;
assign c6301 = ~x65 & ~x375 & ~x403 & ~x431 & ~x460 & ~x486 & ~x599 & ~x600 & ~x601 & ~x615 & ~x629 & ~x685;
assign c6303 =  x436 & ~x128 & ~x156 & ~x242 & ~x360 & ~x678;
assign c6305 =  x439 &  x596 & ~x245;
assign c6307 =  x127 &  x210 &  x348 &  x432 & ~x271 & ~x468;
assign c6309 =  x219;
assign c6311 =  x466 & ~x76 & ~x214 & ~x272 & ~x302 & ~x421 & ~x430 & ~x761;
assign c6313 =  x91 & ~x155;
assign c6315 = ~x0 & ~x30 & ~x32 & ~x53 & ~x136 & ~x392 & ~x404 & ~x433 & ~x460 & ~x546 & ~x751 & ~x774 & ~x777;
assign c6317 =  x79 & ~x714;
assign c6319 =  x538;
assign c6321 = ~x122 & ~x128 & ~x647 & ~x711 & ~x745;
assign c6323 = ~x9 & ~x15 & ~x16 & ~x99 & ~x102 & ~x128 & ~x476 & ~x740 & ~x741 & ~x745 & ~x768;
assign c6325 =  x78 &  x674;
assign c6327 =  x331 &  x362 & ~x584;
assign c6329 =  x109;
assign c6331 =  x439 &  x596;
assign c6333 =  x162 & ~x278 & ~x390;
assign c6335 =  x38 &  x66 &  x95;
assign c6337 =  x154 &  x235 &  x290;
assign c6339 =  x286 & ~x19 & ~x393 & ~x713 & ~x733 & ~x740;
assign c6341 =  x749;
assign c6343 =  x347 &  x374 & ~x75 & ~x121 & ~x493 & ~x684;
assign c6345 =  x269 &  x299;
assign c6347 =  x126 &  x320 &  x347 & ~x269;
assign c6349 =  x428 &  x510 &  x591;
assign c6351 =  x176 & ~x71 & ~x82 & ~x320;
assign c6353 =  x438 &  x596 & ~x277 & ~x670;
assign c6355 =  x167;
assign c6357 = ~x22 & ~x223 & ~x320 & ~x321 & ~x356 & ~x403 & ~x433 & ~x461 & ~x516;
assign c6359 =  x65 &  x412 &  x441;
assign c6361 = ~x72 & ~x75 & ~x99 & ~x126 & ~x156 & ~x694 & ~x740 & ~x745 & ~x767;
assign c6363 =  x545 &  x743 & ~x203 & ~x234 & ~x272 & ~x358 & ~x392 & ~x481;
assign c6365 =  x165;
assign c6367 =  x347 & ~x193 & ~x234 & ~x243 & ~x269 & ~x298;
assign c6369 =  x436 & ~x64 & ~x70 & ~x272 & ~x301 & ~x429 & ~x471 & ~x581 & ~x650 & ~x748;
assign c6371 =  x594 & ~x233 & ~x250 & ~x274 & ~x343 & ~x691 & ~x713;
assign c6373 =  x128 &  x155 & ~x68 & ~x234 & ~x269 & ~x270 & ~x298 & ~x564 & ~x619 & ~x700;
assign c6375 = ~x169 & ~x488 & ~x490 & ~x516 & ~x517 & ~x602 & ~x691 & ~x718;
assign c6377 =  x133 & ~x331 & ~x690;
assign c6379 = ~x73 & ~x127 & ~x128 & ~x152 & ~x156 & ~x673;
assign c6381 =  x160 & ~x125 & ~x319 & ~x346;
assign c6383 =  x707 & ~x572;
assign c6385 =  x465 &  x625 & ~x621;
assign c6387 =  x771 & ~x399 & ~x629 & ~x631;
assign c6389 =  x127 &  x431 &  x716 & ~x63 & ~x343 & ~x383 & ~x583;
assign c6391 =  x354 &  x381 &  x439 &  x467 & ~x129;
assign c6393 =  x217 &  x243 & ~x152 & ~x180;
assign c6395 =  x468 & ~x435;
assign c6397 =  x127 &  x432 &  x716 & ~x4 & ~x148 & ~x201 & ~x412 & ~x471 & ~x619 & ~x675;
assign c6399 =  x66 &  x94 &  x206 &  x207 & ~x23 & ~x365 & ~x564 & ~x644 & ~x699 & ~x730;
assign c6401 =  x232 &  x258 &  x259 & ~x168 & ~x320 & ~x650;
assign c6403 =  x91 & ~x127;
assign c6405 =  x360 & ~x14 & ~x638;
assign c6407 =  x152 &  x319 &  x345 &  x373;
assign c6409 =  x137;
assign c6411 = ~x41 & ~x42 & ~x69 & ~x70 & ~x73 & ~x98 & ~x99 & ~x648 & ~x701 & ~x714 & ~x740 & ~x758;
assign c6413 =  x468 & ~x461;
assign c6415 =  x468 & ~x434;
assign c6417 =  x96 &  x207 & ~x321;
assign c6419 =  x89;
assign c6421 =  x68 &  x685 &  x715 & ~x117 & ~x214 & ~x423 & ~x525 & ~x677 & ~x696;
assign c6423 = ~x207 & ~x236 & ~x460 & ~x600 & ~x601;
assign c6425 =  x320 & ~x268 & ~x269 & ~x412 & ~x680;
assign c6427 =  x743 &  x771 & ~x386 & ~x528 & ~x631 & ~x667;
assign c6429 =  x134;
assign c6431 =  x740 &  x741 &  x770 & ~x611 & ~x637 & ~x660 & ~x662;
assign c6433 =  x358 & ~x73;
assign c6435 =  x111;
assign c6437 =  x122 &  x151 &  x262 &  x290 & ~x43 & ~x75 & ~x103 & ~x420 & ~x758 & ~x760;
assign c6439 =  x65 &  x66 &  x95 & ~x128;
assign c6441 =  x742 &  x743 &  x771 & ~x270 & ~x331 & ~x560;
assign c6443 = ~x37 & ~x65 & ~x461 & ~x488 & ~x546 & ~x658 & ~x685;
assign c6445 =  x144 & ~x71;
assign c6447 =  x105 & ~x97 & ~x98 & ~x633 & ~x661;
assign c6449 =  x274;
assign c6451 =  x107;
assign c6453 =  x741 & ~x25 & ~x36 & ~x302 & ~x314 & ~x391 & ~x416 & ~x426 & ~x471 & ~x475 & ~x658 & ~x661;
assign c6455 =  x743 &  x744 &  x745 & ~x277 & ~x387 & ~x393 & ~x576 & ~x578;
assign c6457 =  x385 & ~x132 & ~x435;
assign c6459 =  x454 &  x456 & ~x42 & ~x744;
assign c6461 =  x771 & ~x219 & ~x398 & ~x418 & ~x426 & ~x557 & ~x610 & ~x633 & ~x660 & ~x661;
assign c6463 =  x346 &  x347 &  x431 & ~x44 & ~x80 & ~x84 & ~x141 & ~x172 & ~x173 & ~x277 & ~x670 & ~x757 & ~x780;
assign c6465 =  x196;
assign c6467 =  x67 &  x95 &  x96 & ~x404 & ~x430 & ~x644 & ~x670;
assign c6469 =  x43 & ~x234 & ~x269;
assign c6471 =  x772 & ~x46 & ~x88 & ~x119 & ~x230 & ~x241 & ~x370 & ~x455 & ~x582 & ~x588 & ~x646 & ~x676 & ~x758;
assign c6473 =  x192;
assign c6475 =  x360 & ~x466;
assign c6477 =  x161 & ~x544;
assign c6479 =  x230 & ~x71 & ~x99;
assign c6481 = ~x17 & ~x84 & ~x104 & ~x156 & ~x160 & ~x183 & ~x184 & ~x211 & ~x212 & ~x254 & ~x308 & ~x333 & ~x498 & ~x525 & ~x616 & ~x668 & ~x700 & ~x703 & ~x723 & ~x736 & ~x764;
assign c6483 =  x119 & ~x663;
assign c6485 =  x273 &  x276;
assign c6487 =  x318 &  x346 & ~x243 & ~x269;
assign c6489 =  x122 &  x316 &  x343;
assign c6491 =  x41 & ~x3 & ~x35 & ~x55 & ~x59 & ~x81 & ~x110 & ~x130 & ~x143 & ~x145 & ~x174 & ~x197 & ~x205 & ~x246 & ~x247 & ~x272 & ~x302 & ~x305 & ~x327 & ~x339 & ~x343 & ~x384 & ~x388 & ~x395 & ~x419 & ~x441 & ~x452 & ~x559 & ~x697 & ~x723 & ~x728 & ~x734 & ~x751 & ~x763 & ~x780;
assign c6493 =  x354 &  x495 & ~x15 & ~x131;
assign c6495 =  x110;
assign c6497 =  x175 & ~x46 & ~x156 & ~x183;
assign c6499 =  x370 & ~x568;
assign c70 =  x204 & ~x384 & ~x497 & ~x508 & ~x591 & ~x650 & ~x721;
assign c72 =  x483 &  x511 & ~x55 & ~x88 & ~x117 & ~x129 & ~x132 & ~x230 & ~x231 & ~x232 & ~x338 & ~x754;
assign c74 =  x334 & ~x56 & ~x103 & ~x116 & ~x161 & ~x175 & ~x191 & ~x225 & ~x475 & ~x530 & ~x566 & ~x595 & ~x609 & ~x621 & ~x652;
assign c76 =  x249 & ~x84 & ~x424 & ~x524 & ~x568 & ~x608 & ~x613 & ~x779;
assign c78 =  x219 & ~x368 & ~x466 & ~x494 & ~x497 & ~x498 & ~x765;
assign c710 =  x263 &  x372 &  x486 & ~x10 & ~x568 & ~x651 & ~x775;
assign c712 =  x349 &  x374 &  x401 &  x511 & ~x79 & ~x147 & ~x175 & ~x202 & ~x228 & ~x310 & ~x779;
assign c714 =  x154 &  x249 & ~x417 & ~x498 & ~x523;
assign c716 =  x149 &  x454 &  x628;
assign c718 =  x203 &  x236 & ~x568 & ~x573;
assign c720 =  x317 &  x403 &  x460 & ~x85 & ~x113 & ~x483 & ~x513 & ~x557 & ~x566 & ~x571 & ~x592 & ~x738 & ~x765;
assign c722 =  x756;
assign c724 =  x55;
assign c726 =  x782;
assign c728 = ~x82 & ~x377 & ~x425 & ~x538 & ~x547 & ~x565 & ~x575 & ~x579 & ~x606 & ~x617 & ~x619 & ~x634 & ~x638 & ~x641 & ~x667 & ~x745;
assign c730 =  x26;
assign c732 =  x321 & ~x149 & ~x161 & ~x175 & ~x176 & ~x201 & ~x202 & ~x257 & ~x615 & ~x645;
assign c734 =  x447 &  x520;
assign c736 =  x448 & ~x277;
assign c738 =  x251 &  x454;
assign c740 =  x306 &  x387 & ~x62 & ~x169 & ~x496 & ~x497;
assign c742 =  x448;
assign c744 =  x404 &  x418 & ~x142 & ~x145 & ~x147 & ~x176 & ~x191 & ~x198 & ~x202 & ~x229 & ~x566 & ~x720 & ~x735;
assign c746 = ~x122 & ~x231 & ~x232 & ~x274 & ~x312 & ~x534 & ~x655 & ~x666 & ~x775;
assign c748 =  x210 &  x246 & ~x611;
assign c750 =  x27;
assign c752 =  x123 &  x274 & ~x540;
assign c754 =  x180 &  x221 & ~x77 & ~x523;
assign c756 =  x222 &  x275 &  x276;
assign c758 =  x111;
assign c760 =  x179 &  x203 & ~x446 & ~x496 & ~x498 & ~x524 & ~x527 & ~x571 & ~x573 & ~x581 & ~x582 & ~x673 & ~x696 & ~x697 & ~x712 & ~x738 & ~x753;
assign c762 =  x71 &  x150 & ~x156;
assign c764 =  x444 & ~x218 & ~x584 & ~x606 & ~x721;
assign c766 =  x350 &  x483 &  x518 &  x519 & ~x102 & ~x144 & ~x161 & ~x167 & ~x252 & ~x280 & ~x697 & ~x705 & ~x782;
assign c768 =  x446 &  x520 & ~x613;
assign c770 =  x386 & ~x655;
assign c772 =  x121 &  x152 &  x186 & ~x552;
assign c774 =  x616;
assign c776 =  x294 &  x408 &  x483 & ~x249;
assign c778 =  x391;
assign c780 =  x28;
assign c782 =  x203 &  x232 & ~x415 & ~x458 & ~x509 & ~x514;
assign c784 =  x513 &  x598 &  x710;
assign c786 =  x297 &  x454 &  x459;
assign c788 =  x455 &  x513 &  x570 & ~x278;
assign c790 =  x71 &  x97 &  x148 & ~x251 & ~x533 & ~x671;
assign c792 =  x94 &  x690 &  x739;
assign c794 =  x457 &  x485 &  x486 &  x514 &  x543 &  x572 & ~x310 & ~x778;
assign c796 =  x420;
assign c798 =  x180 &  x233 & ~x416 & ~x503 & ~x516 & ~x628;
assign c7100 =  x377 & ~x69 & ~x121 & ~x170 & ~x288 & ~x342;
assign c7102 =  x99 &  x353 &  x518 & ~x130 & ~x165 & ~x210;
assign c7104 =  x756;
assign c7106 =  x249 & ~x363 & ~x417 & ~x445 & ~x475 & ~x556 & ~x571 & ~x584 & ~x597 & ~x646 & ~x684 & ~x693 & ~x720;
assign c7108 =  x124 &  x518 & ~x231 & ~x310 & ~x773;
assign c7110 =  x643;
assign c7112 =  x1;
assign c7114 =  x319 &  x348 & ~x352 & ~x446 & ~x512 & ~x591 & ~x652 & ~x653 & ~x679 & ~x741 & ~x768;
assign c7116 =  x446 &  x525;
assign c7118 =  x616;
assign c7120 =  x352 &  x430 &  x458 & ~x13 & ~x82 & ~x117 & ~x119 & ~x163 & ~x252 & ~x775;
assign c7122 =  x342 &  x371 & ~x3 & ~x22 & ~x53 & ~x480 & ~x508 & ~x526 & ~x531 & ~x552 & ~x620;
assign c7124 =  x242 & ~x186 & ~x478 & ~x619 & ~x629 & ~x656;
assign c7126 =  x96 &  x485 &  x520 & ~x231 & ~x256;
assign c7128 =  x655 & ~x312;
assign c7130 =  x124 &  x192 & ~x555;
assign c7132 =  x112;
assign c7136 =  x111;
assign c7138 =  x454 &  x500 & ~x216;
assign c7140 =  x322 &  x427 & ~x117 & ~x199 & ~x311 & ~x685 & ~x687;
assign c7142 =  x207 & ~x456 & ~x484 & ~x542 & ~x565 & ~x569 & ~x624 & ~x702;
assign c7144 = ~x35 & ~x36 & ~x40 & ~x41 & ~x42 & ~x59 & ~x68 & ~x69 & ~x76 & ~x113 & ~x117 & ~x120 & ~x121 & ~x133 & ~x142 & ~x149 & ~x175 & ~x184 & ~x194 & ~x204 & ~x229 & ~x231 & ~x310 & ~x616 & ~x665 & ~x678 & ~x679 & ~x681 & ~x723;
assign c7146 =  x162 &  x180 & ~x479 & ~x573;
assign c7148 =  x334 & ~x5 & ~x7 & ~x21 & ~x29 & ~x32 & ~x45 & ~x71 & ~x104 & ~x112 & ~x117 & ~x160 & ~x161 & ~x169 & ~x195 & ~x224 & ~x475 & ~x523 & ~x566 & ~x594 & ~x611 & ~x638 & ~x639 & ~x643 & ~x651 & ~x659 & ~x664 & ~x674 & ~x677 & ~x679 & ~x692 & ~x694 & ~x760 & ~x761;
assign c7150 =  x313 &  x400 & ~x507 & ~x511 & ~x552 & ~x566 & ~x585 & ~x591;
assign c7152 =  x500 & ~x109 & ~x171 & ~x191 & ~x216 & ~x622 & ~x624 & ~x637 & ~x639;
assign c7154 =  x180 &  x298 &  x455 & ~x619;
assign c7156 =  x352 &  x356 & ~x12 & ~x746 & ~x747;
assign c7158 =  x350 &  x600 & ~x135 & ~x186 & ~x253 & ~x338;
assign c7160 =  x377 & ~x63 & ~x148 & ~x342 & ~x619 & ~x644 & ~x686 & ~x695 & ~x730;
assign c7162 =  x418 & ~x40 & ~x117 & ~x147 & ~x180 & ~x216 & ~x257 & ~x258 & ~x766;
assign c7164 =  x27;
assign c7166 =  x95 &  x203 & ~x438 & ~x452 & ~x523 & ~x526 & ~x586 & ~x670 & ~x761 & ~x762;
assign c7168 =  x297 &  x320 &  x520 & ~x60 & ~x198 & ~x201 & ~x701 & ~x761;
assign c7170 =  x94 &  x316;
assign c7172 =  x55;
assign c7174 = ~x19 & ~x116 & ~x486 & ~x515 & ~x525 & ~x527 & ~x536 & ~x565 & ~x573 & ~x598 & ~x608 & ~x621 & ~x776;
assign c7176 =  x456 &  x552 & ~x211 & ~x257;
assign c7178 =  x184 &  x185 &  x186 & ~x497 & ~x534 & ~x549;
assign c7180 =  x494 & ~x228 & ~x259 & ~x285 & ~x773;
assign c7182 =  x448;
assign c7184 =  x111;
assign c7186 =  x97 &  x163 & ~x456 & ~x765;
assign c7188 =  x95 &  x692 & ~x596 & ~x624;
assign c7190 =  x308;
assign c7192 =  x351 &  x510 & ~x90 & ~x117 & ~x171 & ~x231 & ~x279 & ~x281 & ~x283 & ~x698 & ~x701 & ~x752;
assign c7194 =  x756;
assign c7196 =  x184 &  x208 &  x260 & ~x494 & ~x497 & ~x522 & ~x552 & ~x570;
assign c7198 =  x27;
assign c7200 =  x390 &  x442 & ~x131 & ~x523;
assign c7202 = ~x7 & ~x19 & ~x70 & ~x79 & ~x103 & ~x105 & ~x117 & ~x140 & ~x145 & ~x196 & ~x454 & ~x507 & ~x608 & ~x612 & ~x634 & ~x674 & ~x686 & ~x709 & ~x729 & ~x743 & ~x749;
assign c7204 =  x401 &  x430 &  x459 &  x574 & ~x569 & ~x571;
assign c7206 =  x93 &  x118 & ~x497;
assign c7208 =  x219 & ~x61 & ~x484 & ~x523 & ~x554 & ~x624 & ~x642;
assign c7210 = ~x118 & ~x121 & ~x143 & ~x483 & ~x526 & ~x542 & ~x567 & ~x684 & ~x714;
assign c7212 =  x419 &  x470 &  x471 & ~x649 & ~x651;
assign c7214 =  x350 &  x351 &  x373 &  x398 & ~x747;
assign c7216 =  x417 &  x522 & ~x130 & ~x158 & ~x201 & ~x696;
assign c7218 =  x455 &  x485 &  x514 &  x571 & ~x254;
assign c7220 =  x83;
assign c7222 = ~x395 & ~x455 & ~x479 & ~x509 & ~x524 & ~x525 & ~x535 & ~x550 & ~x566 & ~x578 & ~x596 & ~x634 & ~x636 & ~x673 & ~x691 & ~x707 & ~x732 & ~x733 & ~x741 & ~x751 & ~x768;
assign c7224 = ~x58 & ~x117 & ~x196 & ~x243 & ~x425 & ~x435 & ~x492 & ~x537 & ~x566 & ~x567 & ~x637 & ~x648 & ~x649 & ~x671 & ~x754 & ~x757;
assign c7226 =  x428 &  x455 &  x485 &  x513 &  x542 & ~x222 & ~x645 & ~x702 & ~x756 & ~x773;
assign c7228 =  x353 &  x574 & ~x168 & ~x259;
assign c7230 =  x404 &  x607 & ~x200;
assign c7232 =  x495 & ~x29 & ~x135 & ~x145 & ~x160 & ~x170 & ~x189 & ~x218 & ~x606 & ~x619 & ~x738;
assign c7234 =  x203 & ~x34 & ~x295 & ~x409 & ~x416 & ~x418 & ~x419 & ~x523 & ~x636 & ~x637 & ~x723 & ~x773;
assign c7236 =  x0;
assign c7238 =  x458 &  x574 & ~x61 & ~x568 & ~x655;
assign c7240 =  x236 &  x263 &  x346 &  x349 &  x483;
assign c7242 =  x373 &  x455 &  x520 & ~x117 & ~x189;
assign c7244 =  x233 & ~x1 & ~x39 & ~x41 & ~x42 & ~x50 & ~x563 & ~x568 & ~x591 & ~x634 & ~x636 & ~x646 & ~x718 & ~x719 & ~x739 & ~x765;
assign c7246 = ~x50 & ~x53 & ~x115 & ~x227 & ~x425 & ~x450 & ~x535 & ~x560 & ~x573 & ~x594 & ~x611 & ~x636 & ~x667 & ~x697 & ~x708 & ~x773;
assign c7248 =  x387 &  x410 & ~x6 & ~x468 & ~x469 & ~x497 & ~x678 & ~x743;
assign c7250 = ~x47 & ~x64 & ~x456 & ~x483 & ~x512 & ~x534 & ~x572 & ~x581 & ~x593 & ~x608 & ~x612 & ~x624 & ~x711 & ~x768;
assign c7252 =  x227 &  x253;
assign c7254 = ~x1 & ~x3 & ~x6 & ~x111 & ~x117 & ~x432 & ~x447 & ~x493 & ~x501 & ~x508 & ~x518 & ~x561 & ~x580 & ~x591 & ~x637 & ~x716 & ~x743 & ~x744 & ~x765 & ~x775;
assign c7256 = ~x22 & ~x82 & ~x115 & ~x197 & ~x484 & ~x486 & ~x500 & ~x555 & ~x589 & ~x591 & ~x601 & ~x626 & ~x690;
assign c7258 =  x363 &  x442 & ~x501;
assign c7260 =  x149 &  x209 &  x237 & ~x538 & ~x548 & ~x722;
assign c7264 =  x416 &  x441 &  x442 & ~x32 & ~x104 & ~x610 & ~x683 & ~x735 & ~x736 & ~x740;
assign c7266 =  x656 &  x690 &  x739;
assign c7268 = ~x281 & ~x418 & ~x451 & ~x537 & ~x558 & ~x568 & ~x579 & ~x585 & ~x606 & ~x634 & ~x681 & ~x697 & ~x744 & ~x764 & ~x779 & ~x783;
assign c7270 = ~x19 & ~x22 & ~x57 & ~x352 & ~x363 & ~x390 & ~x419 & ~x497 & ~x498 & ~x523 & ~x554 & ~x571 & ~x587 & ~x594 & ~x637 & ~x665 & ~x737;
assign c7272 =  x190 &  x358 & ~x497;
assign c7274 =  x151 &  x177 &  x263 & ~x770;
assign c7276 =  x27;
assign c7278 =  x485 &  x570 &  x598 &  x710;
assign c7280 =  x294 &  x486 &  x544;
assign c7282 =  x783;
assign c7284 =  x124 &  x213 &  x317 &  x344 & ~x0 & ~x9 & ~x115 & ~x141 & ~x224 & ~x643 & ~x696;
assign c7286 =  x96 &  x100;
assign c7288 =  x124 &  x458 &  x572 &  x602;
assign c7290 =  x275 &  x345 & ~x86 & ~x481 & ~x511 & ~x594 & ~x649 & ~x650 & ~x690;
assign c7292 =  x94 &  x480 &  x766;
assign c7294 =  x615;
assign c7296 =  x25;
assign c7298 =  x139;
assign c7300 =  x176 & ~x425 & ~x457 & ~x467 & ~x496 & ~x497 & ~x498 & ~x565 & ~x626 & ~x703;
assign c7302 =  x248 &  x316 & ~x450 & ~x524;
assign c7304 =  x656 &  x689 & ~x624;
assign c7306 =  x349 &  x408 &  x455 &  x518 & ~x226 & ~x774;
assign c7308 =  x28;
assign c7310 =  x94;
assign c7312 =  x453 &  x664 &  x710;
assign c7314 =  x26;
assign c7316 =  x420 &  x532;
assign c7320 =  x350 &  x389 & ~x143 & ~x649;
assign c7322 =  x783;
assign c7324 =  x27;
assign c7326 =  x455 &  x510 &  x602 & ~x306 & ~x311 & ~x314;
assign c7328 =  x380 &  x620;
assign c7330 =  x181 &  x233 & ~x4 & ~x437 & ~x441;
assign c7332 =  x156 &  x278 & ~x526 & ~x528 & ~x552;
assign c7334 =  x727;
assign c7336 =  x459 &  x544 & ~x484 & ~x626;
assign c7338 =  x0;
assign c7340 =  x350 &  x446 &  x500 &  x525;
assign c7342 =  x485 &  x542 &  x599 &  x627 & ~x6 & ~x50 & ~x59 & ~x130 & ~x622 & ~x750;
assign c7344 =  x280;
assign c7346 = ~x7 & ~x24 & ~x72 & ~x76 & ~x79 & ~x80 & ~x113 & ~x141 & ~x143 & ~x165 & ~x216 & ~x227 & ~x409 & ~x425 & ~x485 & ~x541 & ~x582 & ~x619 & ~x653 & ~x679 & ~x682 & ~x690 & ~x709 & ~x715 & ~x720 & ~x734 & ~x746 & ~x748 & ~x752 & ~x762 & ~x766 & ~x775;
assign c7348 =  x399 &  x485 &  x513 &  x542 &  x599;
assign c7350 =  x483 &  x485 &  x544 & ~x58 & ~x114 & ~x145 & ~x228 & ~x282 & ~x283 & ~x335 & ~x772;
assign c7352 = ~x125 & ~x160 & ~x177 & ~x228 & ~x671 & ~x716 & ~x726 & ~x735 & ~x739 & ~x768;
assign c7354 =  x427 &  x428 &  x485 &  x513 &  x542 & ~x226;
assign c7356 =  x180 &  x250;
assign c7358 =  x389 &  x412 &  x413 & ~x496 & ~x497;
assign c7360 =  x55;
assign c7362 =  x26;
assign c7364 =  x426 &  x455 &  x485 &  x513 & ~x82 & ~x106 & ~x668 & ~x693 & ~x732;
assign c7366 = ~x27 & ~x94 & ~x134 & ~x149 & ~x175 & ~x204 & ~x232 & ~x255 & ~x310 & ~x312 & ~x651 & ~x708 & ~x725 & ~x743 & ~x774;
assign c7368 =  x372 &  x454 & ~x23 & ~x47 & ~x166 & ~x369 & ~x559 & ~x781;
assign c7370 =  x404 & ~x40 & ~x58 & ~x113 & ~x121 & ~x219 & ~x232 & ~x645 & ~x778;
assign c7372 = ~x12 & ~x48 & ~x73 & ~x79 & ~x83 & ~x168 & ~x324 & ~x403 & ~x474 & ~x500 & ~x531 & ~x535 & ~x549 & ~x556 & ~x558 & ~x614 & ~x618 & ~x696 & ~x709 & ~x718 & ~x773;
assign c7374 =  x476;
assign c7376 =  x548 &  x565 & ~x230 & ~x248;
assign c7378 =  x27;
assign c7380 =  x376 & ~x191 & ~x231 & ~x232 & ~x257 & ~x720 & ~x746;
assign c7382 =  x472 &  x494 & ~x159 & ~x193 & ~x280 & ~x619;
assign c7384 =  x56;
assign c7386 =  x354 &  x375 & ~x40 & ~x93 & ~x200 & ~x586;
assign c7388 =  x196 &  x643;
assign c7390 =  x334 & ~x113 & ~x232 & ~x528;
assign c7392 =  x278 & ~x390 & ~x497 & ~x510 & ~x569 & ~x626;
assign c7394 =  x165;
assign c7396 =  x756 &  x760;
assign c7398 =  x185 &  x232 &  x233 &  x260 & ~x458 & ~x550;
assign c7400 =  x95 &  x618;
assign c7402 =  x408 & ~x176 & ~x232;
assign c7404 =  x158 &  x221 & ~x479;
assign c7406 =  x483 &  x602 & ~x202 & ~x249 & ~x285 & ~x755;
assign c7408 =  x280;
assign c7410 =  x471 & ~x1 & ~x89 & ~x117 & ~x130 & ~x142 & ~x143 & ~x158 & ~x164 & ~x221 & ~x531 & ~x582 & ~x639 & ~x702;
assign c7412 =  x267 &  x269 &  x292 & ~x20 & ~x607;
assign c7414 =  x288 & ~x33 & ~x57 & ~x60 & ~x106 & ~x421 & ~x455 & ~x478 & ~x482 & ~x492 & ~x534 & ~x565 & ~x568 & ~x585 & ~x594 & ~x621 & ~x622 & ~x655 & ~x681 & ~x694 & ~x737 & ~x739;
assign c7416 =  x417 & ~x11 & ~x33 & ~x91 & ~x115 & ~x225 & ~x288 & ~x679 & ~x702 & ~x732 & ~x739 & ~x779 & ~x780;
assign c7418 =  x472 & ~x232;
assign c7420 =  x500 &  x573;
assign c7422 = ~x26 & ~x34 & ~x69 & ~x146 & ~x165 & ~x199 & ~x204 & ~x231 & ~x259 & ~x568 & ~x569 & ~x570 & ~x582 & ~x668 & ~x723 & ~x739 & ~x758 & ~x759 & ~x767 & ~x769 & ~x773;
assign c7424 =  x99 &  x246 & ~x615 & ~x649 & ~x716;
assign c7426 =  x700;
assign c7428 =  x233 & ~x271 & ~x455 & ~x552 & ~x634 & ~x635 & ~x637 & ~x666;
assign c7430 =  x27;
assign c7432 =  x353 & ~x29 & ~x32 & ~x93 & ~x104 & ~x117 & ~x118 & ~x119 & ~x142 & ~x149 & ~x216 & ~x220 & ~x257 & ~x646 & ~x693 & ~x699 & ~x721 & ~x731 & ~x775;
assign c7434 =  x334 & ~x117 & ~x142 & ~x497 & ~x499 & ~x500 & ~x524 & ~x529 & ~x556 & ~x595 & ~x653;
assign c7436 =  x350 &  x400 & ~x171 & ~x200 & ~x231 & ~x248 & ~x625;
assign c7438 =  x71 &  x486 & ~x687;
assign c7440 = ~x43 & ~x104 & ~x115 & ~x156 & ~x257 & ~x284 & ~x500 & ~x526 & ~x534 & ~x558 & ~x568 & ~x624 & ~x714 & ~x755 & ~x765 & ~x766;
assign c7442 =  x395 &  x396 & ~x53 & ~x90 & ~x113 & ~x161 & ~x187 & ~x534 & ~x613 & ~x639 & ~x663 & ~x666 & ~x669 & ~x709 & ~x738;
assign c7444 =  x236 &  x379 &  x628 &  x656 & ~x10 & ~x117 & ~x283;
assign c7446 =  x24 &  x454;
assign c7448 =  x379 &  x428 &  x510 & ~x108 & ~x220 & ~x258;
assign c7450 = ~x62 & ~x485 & ~x516 & ~x523 & ~x569 & ~x656 & ~x680 & ~x773;
assign c7452 =  x270 &  x294 &  x345 & ~x655 & ~x714;
assign c7454 = ~x87 & ~x140 & ~x197 & ~x408 & ~x472 & ~x479 & ~x510 & ~x545 & ~x566 & ~x636 & ~x719;
assign c7456 =  x305 & ~x335 & ~x472 & ~x565 & ~x654 & ~x761;
assign c7458 =  x486 &  x543 &  x544 &  x572 & ~x130 & ~x171 & ~x568 & ~x615 & ~x621 & ~x708 & ~x726 & ~x746;
assign c7460 = ~x324 & ~x444 & ~x446 & ~x458 & ~x496 & ~x497 & ~x505 & ~x516 & ~x526 & ~x534 & ~x541 & ~x582 & ~x598 & ~x640 & ~x684 & ~x714 & ~x723;
assign c7462 =  x408 &  x415 & ~x677 & ~x775;
assign c7464 =  x408 &  x483 & ~x35 & ~x117 & ~x228 & ~x286;
assign c7466 =  x167;
assign c7468 =  x615;
assign c7470 = ~x59 & ~x295 & ~x435 & ~x436 & ~x480 & ~x508 & ~x536 & ~x569 & ~x577 & ~x589 & ~x608 & ~x626 & ~x648 & ~x748;
assign c7472 =  x471 &  x520 & ~x147 & ~x249 & ~x708;
assign c7474 =  x55;
assign c7476 =  x220 & ~x456 & ~x457;
assign c7478 = ~x0 & ~x7 & ~x11 & ~x326 & ~x478 & ~x508 & ~x530 & ~x532 & ~x537 & ~x540 & ~x558 & ~x579 & ~x588 & ~x596 & ~x600 & ~x608 & ~x609 & ~x624 & ~x719;
assign c7480 =  x25;
assign c7482 =  x125 &  x273 &  x518;
assign c7484 =  x418 & ~x34 & ~x83 & ~x93 & ~x149 & ~x159 & ~x202 & ~x204 & ~x207 & ~x221 & ~x615 & ~x637 & ~x719 & ~x771 & ~x777;
assign c7486 =  x181 &  x182 &  x233 & ~x34 & ~x412 & ~x580 & ~x619;
assign c7488 =  x417 &  x520 & ~x219;
assign c7490 =  x232 &  x233 & ~x456 & ~x523 & ~x541 & ~x555 & ~x673;
assign c7492 =  x122 &  x154 &  x277 & ~x497;
assign c7494 =  x324 &  x374 &  x483 & ~x184 & ~x283;
assign c7496 =  x27;
assign c7498 =  x95 & ~x411 & ~x608;
assign c71 =  x556 & ~x54 & ~x515;
assign c73 =  x341 &  x369 & ~x206 & ~x235 & ~x262;
assign c75 = ~x26 & ~x30 & ~x58 & ~x111 & ~x165 & ~x168 & ~x216 & ~x254 & ~x275 & ~x277 & ~x301 & ~x304 & ~x359 & ~x361 & ~x367 & ~x396 & ~x397 & ~x444 & ~x445 & ~x448 & ~x473 & ~x479 & ~x506 & ~x528 & ~x536 & ~x609 & ~x614 & ~x616 & ~x619 & ~x665 & ~x670 & ~x672 & ~x699 & ~x702 & ~x724 & ~x726 & ~x735 & ~x754 & ~x755;
assign c77 =  x286 &  x549 &  x576 &  x603 & ~x24 & ~x753;
assign c79 =  x482 &  x537 & ~x4 & ~x52 & ~x81 & ~x110 & ~x167 & ~x193 & ~x632 & ~x707 & ~x763;
assign c711 =  x569 &  x595 &  x596 &  x623 &  x624 & ~x27 & ~x48 & ~x109;
assign c713 =  x489 &  x517 & ~x7 & ~x214 & ~x239 & ~x242 & ~x296 & ~x587 & ~x729;
assign c715 = ~x13 & ~x51 & ~x78 & ~x195 & ~x223 & ~x249 & ~x338 & ~x340 & ~x366 & ~x367 & ~x387 & ~x388 & ~x391 & ~x414 & ~x444 & ~x554 & ~x581 & ~x582 & ~x596 & ~x647 & ~x700 & ~x702 & ~x706 & ~x763 & ~x781;
assign c717 =  x155 &  x183 & ~x32 & ~x59 & ~x83 & ~x136 & ~x304 & ~x309 & ~x415 & ~x416 & ~x451 & ~x472 & ~x505 & ~x528 & ~x671;
assign c719 =  x594 &  x621 &  x622 & ~x23 & ~x28 & ~x57 & ~x114 & ~x198 & ~x279 & ~x672 & ~x699 & ~x764 & ~x768;
assign c721 = ~x132 & ~x203 & ~x205 & ~x254 & ~x275 & ~x334 & ~x394 & ~x415 & ~x507 & ~x589 & ~x637 & ~x677 & ~x696;
assign c723 =  x318 & ~x131 & ~x275 & ~x359 & ~x360 & ~x369 & ~x387 & ~x424 & ~x554;
assign c725 =  x312 & ~x151 & ~x234;
assign c727 =  x639 & ~x54 & ~x364 & ~x739 & ~x740;
assign c729 =  x159 &  x237 & ~x30 & ~x151 & ~x448 & ~x756;
assign c731 =  x499 &  x553 &  x581;
assign c733 =  x501 & ~x350 & ~x351 & ~x430;
assign c735 = ~x208 & ~x236 & ~x237 & ~x263 & ~x264 & ~x265 & ~x770;
assign c737 =  x550 &  x576 &  x577 &  x578 &  x603 &  x604 &  x605 & ~x32 & ~x167 & ~x781;
assign c739 =  x611 & ~x518;
assign c741 = ~x8 & ~x27 & ~x265 & ~x291 & ~x292 & ~x317 & ~x318 & ~x319 & ~x344 & ~x345 & ~x346 & ~x372 & ~x373 & ~x399 & ~x400 & ~x427;
assign c743 =  x228 &  x464 & ~x469;
assign c745 =  x409 &  x437 & ~x23 & ~x58 & ~x142 & ~x198 & ~x222 & ~x275 & ~x277 & ~x282 & ~x337 & ~x361 & ~x394 & ~x445 & ~x477 & ~x478 & ~x499 & ~x557 & ~x563 & ~x584 & ~x591 & ~x704 & ~x724 & ~x728 & ~x765;
assign c747 = ~x1 & ~x2 & ~x5 & ~x20 & ~x88 & ~x167 & ~x302 & ~x348 & ~x387 & ~x404 & ~x430 & ~x431 & ~x444 & ~x721;
assign c749 = ~x32 & ~x106 & ~x312 & ~x340 & ~x369 & ~x387 & ~x390 & ~x427 & ~x663 & ~x697 & ~x724;
assign c751 =  x332 &  x360 & ~x20 & ~x299 & ~x439;
assign c753 =  x435 &  x517 & ~x56 & ~x111 & ~x361 & ~x425 & ~x610 & ~x621 & ~x728;
assign c755 = ~x13 & ~x27 & ~x45 & ~x127 & ~x156 & ~x183 & ~x236 & ~x263 & ~x265 & ~x749 & ~x757;
assign c757 =  x170;
assign c759 =  x361 & ~x241 & ~x325 & ~x384 & ~x439;
assign c761 =  x685 &  x686 & ~x31 & ~x80 & ~x136 & ~x139 & ~x282 & ~x334 & ~x361 & ~x364 & ~x388 & ~x417 & ~x445 & ~x470 & ~x475 & ~x498 & ~x588 & ~x612 & ~x614 & ~x676 & ~x758;
assign c763 = ~x236 & ~x237 & ~x263 & ~x264 & ~x265 & ~x266 & ~x292 & ~x750;
assign c765 = ~x24 & ~x151 & ~x178 & ~x180 & ~x304 & ~x307 & ~x331 & ~x336 & ~x387 & ~x388 & ~x445 & ~x529 & ~x728 & ~x757 & ~x761 & ~x776;
assign c767 =  x743 &  x771 & ~x50 & ~x59 & ~x107 & ~x167 & ~x168 & ~x222 & ~x279 & ~x281 & ~x363 & ~x423 & ~x593;
assign c769 =  x266 & ~x253 & ~x304 & ~x305 & ~x328 & ~x388 & ~x661;
assign c771 = ~x5 & ~x16 & ~x45 & ~x53 & ~x83 & ~x84 & ~x98 & ~x155 & ~x187 & ~x210 & ~x238 & ~x239 & ~x336 & ~x468 & ~x496 & ~x526 & ~x614 & ~x640 & ~x676 & ~x697 & ~x700 & ~x705 & ~x746 & ~x750;
assign c773 = ~x236 & ~x345 & ~x371 & ~x372 & ~x373 & ~x400 & ~x427;
assign c775 =  x597 & ~x236 & ~x263 & ~x264;
assign c777 =  x216 &  x526;
assign c779 =  x341 &  x553;
assign c781 = ~x100 & ~x103 & ~x151 & ~x182 & ~x208 & ~x211 & ~x753;
assign c783 =  x509 & ~x22 & ~x72 & ~x137 & ~x267 & ~x270 & ~x326 & ~x382;
assign c785 =  x557 & ~x438;
assign c787 = ~x108 & ~x112 & ~x118 & ~x133 & ~x135 & ~x136 & ~x275 & ~x306 & ~x360 & ~x367 & ~x369 & ~x386 & ~x389 & ~x395 & ~x396 & ~x442 & ~x539 & ~x562 & ~x594 & ~x652 & ~x692 & ~x707 & ~x708;
assign c789 =  x312 &  x593;
assign c791 =  x461 &  x489 &  x568 & ~x79;
assign c793 = ~x97 & ~x151 & ~x178 & ~x349 & ~x404 & ~x459;
assign c795 =  x566 &  x593 &  x594 &  x621 & ~x45 & ~x729 & ~x758;
assign c797 =  x289 & ~x183 & ~x237 & ~x239 & ~x266 & ~x297 & ~x337;
assign c799 = ~x37 & ~x349 & ~x376 & ~x378 & ~x430 & ~x431 & ~x513 & ~x539 & ~x756;
assign c7101 =  x286 & ~x206 & ~x235 & ~x236;
assign c7103 = ~x155 & ~x180 & ~x208 & ~x235 & ~x236 & ~x439 & ~x672;
assign c7105 = ~x87 & ~x193 & ~x194 & ~x249 & ~x258 & ~x282 & ~x328 & ~x330 & ~x357 & ~x369 & ~x393 & ~x425 & ~x474 & ~x558 & ~x585 & ~x593 & ~x617 & ~x621 & ~x698 & ~x702 & ~x728 & ~x734 & ~x758 & ~x780 & ~x781;
assign c7107 = ~x39 & ~x54 & ~x96 & ~x151 & ~x167 & ~x178 & ~x387 & ~x388 & ~x390 & ~x391 & ~x444 & ~x558;
assign c7109 =  x402 &  x539 &  x566 & ~x100 & ~x394 & ~x528 & ~x615 & ~x754;
assign c7111 = ~x15 & ~x212 & ~x214 & ~x296 & ~x422 & ~x476 & ~x631 & ~x632 & ~x660;
assign c7113 =  x743 &  x744 &  x745 & ~x575;
assign c7115 =  x584 & ~x658;
assign c7117 = ~x322 & ~x349 & ~x402 & ~x404 & ~x405 & ~x430 & ~x431 & ~x459 & ~x488 & ~x513 & ~x697 & ~x728 & ~x773;
assign c7119 =  x554 &  x555 & ~x355 & ~x383;
assign c7121 =  x584 &  x611 &  x612;
assign c7123 =  x368;
assign c7125 =  x229 & ~x236 & ~x237 & ~x263 & ~x264 & ~x265;
assign c7127 =  x555 &  x582 &  x637;
assign c7129 = ~x50 & ~x144 & ~x169 & ~x407 & ~x431 & ~x439 & ~x462 & ~x463 & ~x485 & ~x491 & ~x515 & ~x518 & ~x572 & ~x652 & ~x679 & ~x757;
assign c7131 =  x603 &  x630 &  x631 & ~x31 & ~x169 & ~x334 & ~x361 & ~x440 & ~x441 & ~x450 & ~x453 & ~x478 & ~x507 & ~x538 & ~x565 & ~x586 & ~x588 & ~x621 & ~x698 & ~x779;
assign c7133 =  x717 & ~x29 & ~x76 & ~x89 & ~x135 & ~x246 & ~x391 & ~x582 & ~x731 & ~x764;
assign c7135 = ~x248 & ~x274 & ~x277 & ~x284 & ~x301 & ~x308 & ~x367 & ~x388 & ~x395 & ~x499 & ~x511 & ~x527 & ~x533 & ~x558 & ~x616 & ~x643 & ~x723 & ~x762 & ~x781;
assign c7137 = ~x20 & ~x53 & ~x79 & ~x105 & ~x107 & ~x110 & ~x135 & ~x140 & ~x165 & ~x166 & ~x253 & ~x273 & ~x303 & ~x304 & ~x307 & ~x332 & ~x336 & ~x365 & ~x369 & ~x387 & ~x417 & ~x444 & ~x446 & ~x536 & ~x589 & ~x622 & ~x639 & ~x664 & ~x700 & ~x724 & ~x731;
assign c7139 = ~x154 & ~x182 & ~x237 & ~x263 & ~x264 & ~x265 & ~x292 & ~x307;
assign c7141 = ~x18 & ~x79 & ~x136 & ~x161 & ~x195 & ~x281 & ~x302 & ~x304 & ~x306 & ~x339 & ~x536 & ~x539 & ~x616 & ~x618 & ~x755;
assign c7143 = ~x292 & ~x293 & ~x320 & ~x345 & ~x346 & ~x347 & ~x373 & ~x400 & ~x401;
assign c7145 =  x284 & ~x263 & ~x318 & ~x345;
assign c7147 =  x62 &  x91 &  x119 &  x120;
assign c7149 =  x257 & ~x319 & ~x344 & ~x345 & ~x346 & ~x400 & ~x427;
assign c7151 =  x660 &  x661 &  x687 &  x688 & ~x371 & ~x703;
assign c7153 =  x41 & ~x91 & ~x142 & ~x273 & ~x274 & ~x360 & ~x362 & ~x642;
assign c7155 =  x537 & ~x60 & ~x125 & ~x353 & ~x768;
assign c7157 =  x497 &  x524 &  x551 &  x578 & ~x81;
assign c7159 =  x567 &  x568 & ~x114 & ~x298 & ~x783;
assign c7161 =  x651 &  x678 &  x679 &  x680;
assign c7163 = ~x22 & ~x24 & ~x62 & ~x351 & ~x404 & ~x405 & ~x431 & ~x432 & ~x461 & ~x464 & ~x491 & ~x514 & ~x515 & ~x753;
assign c7165 =  x604 &  x605 &  x631 &  x632 &  x659 & ~x16 & ~x46 & ~x363 & ~x419 & ~x420 & ~x477 & ~x591 & ~x615 & ~x644 & ~x735;
assign c7167 =  x567 &  x594 &  x595 & ~x98 & ~x126;
assign c7169 =  x501 & ~x439 & ~x573;
assign c7171 = ~x37 & ~x66 & ~x67 & ~x208 & ~x236 & ~x263 & ~x264 & ~x290 & ~x446 & ~x705;
assign c7173 =  x432 &  x568 & ~x44 & ~x45 & ~x99 & ~x126 & ~x756;
assign c7175 =  x469 &  x496 &  x497 &  x524 &  x551;
assign c7177 =  x613;
assign c7179 =  x434 & ~x344 & ~x347 & ~x371 & ~x374 & ~x376 & ~x401;
assign c7181 =  x155 &  x183 &  x239 &  x267 &  x295 & ~x334 & ~x445;
assign c7183 =  x501 & ~x518 & ~x546 & ~x729;
assign c7185 =  x582 & ~x405;
assign c7187 = ~x7 & ~x14 & ~x21 & ~x27 & ~x44 & ~x73 & ~x78 & ~x84 & ~x87 & ~x103 & ~x108 & ~x114 & ~x167 & ~x183 & ~x184 & ~x185 & ~x187 & ~x239 & ~x266 & ~x567 & ~x618 & ~x723 & ~x735 & ~x782;
assign c7189 =  x714 &  x715 &  x741 &  x742 & ~x111 & ~x197 & ~x446 & ~x502 & ~x531 & ~x565 & ~x588 & ~x617 & ~x636 & ~x641 & ~x756;
assign c7191 =  x116 & ~x37 & ~x111;
assign c7193 = ~x355 & ~x381 & ~x383 & ~x433 & ~x439 & ~x491;
assign c7195 =  x332 &  x360 &  x388 & ~x14 & ~x15 & ~x383 & ~x750;
assign c7197 =  x742 & ~x0 & ~x2 & ~x54 & ~x79 & ~x86 & ~x136 & ~x143 & ~x311 & ~x366 & ~x394 & ~x395 & ~x446 & ~x551 & ~x616 & ~x636 & ~x638 & ~x668 & ~x697;
assign c7199 = ~x35 & ~x105 & ~x135 & ~x158 & ~x211 & ~x213 & ~x239 & ~x241 & ~x268 & ~x295 & ~x299 & ~x323;
assign c7201 = ~x297 & ~x349 & ~x350 & ~x354 & ~x382 & ~x383 & ~x411 & ~x439 & ~x734;
assign c7203 =  x314 &  x333 &  x343 & ~x211;
assign c7205 = ~x99 & ~x166 & ~x420 & ~x464 & ~x490 & ~x572;
assign c7207 = ~x43 & ~x102 & ~x159 & ~x236 & ~x237 & ~x264 & ~x265 & ~x365 & ~x390 & ~x394 & ~x613 & ~x701;
assign c7209 = ~x126 & ~x180 & ~x208 & ~x238 & ~x295 & ~x645;
assign c7211 =  x668 & ~x29 & ~x135;
assign c7213 =  x706 &  x707 &  x708;
assign c7215 =  x686 &  x687 & ~x2 & ~x143 & ~x276 & ~x279 & ~x304 & ~x306 & ~x310 & ~x333 & ~x444 & ~x471 & ~x558 & ~x562 & ~x699;
assign c7217 =  x624 &  x681 &  x712;
assign c7219 = ~x21 & ~x76 & ~x78 & ~x253 & ~x274 & ~x281 & ~x328 & ~x332 & ~x333 & ~x358 & ~x360 & ~x362 & ~x384 & ~x387 & ~x390 & ~x419 & ~x475 & ~x537 & ~x555 & ~x559 & ~x560 & ~x672 & ~x702;
assign c7221 =  x406 &  x462 & ~x187 & ~x239 & ~x337 & ~x554 & ~x556 & ~x754;
assign c7223 =  x312 &  x536 &  x564;
assign c7225 =  x630 & ~x346 & ~x371 & ~x372 & ~x373 & ~x400;
assign c7227 =  x537 & ~x268 & ~x297 & ~x298 & ~x640;
assign c7229 = ~x64 & ~x137 & ~x253 & ~x405 & ~x431 & ~x459 & ~x491 & ~x596;
assign c7231 = ~x24 & ~x27 & ~x31 & ~x61 & ~x91 & ~x119 & ~x195 & ~x216 & ~x247 & ~x274 & ~x277 & ~x306 & ~x308 & ~x332 & ~x334 & ~x360 & ~x369 & ~x391 & ~x393 & ~x424 & ~x425 & ~x469 & ~x479 & ~x617 & ~x618 & ~x620 & ~x734 & ~x751;
assign c7233 = ~x297 & ~x404 & ~x405 & ~x437 & ~x439 & ~x490 & ~x515;
assign c7235 =  x633 &  x634 &  x660 &  x661 &  x688 & ~x21 & ~x22 & ~x28 & ~x55 & ~x80 & ~x167 & ~x564 & ~x729 & ~x782;
assign c7237 = ~x54 & ~x81 & ~x347 & ~x348 & ~x349 & ~x350 & ~x375 & ~x402 & ~x404 & ~x430 & ~x432 & ~x514 & ~x595 & ~x650 & ~x671 & ~x700 & ~x737 & ~x764;
assign c7239 =  x432 & ~x183 & ~x237 & ~x265;
assign c7241 =  x619 &  x646 &  x647 &  x675;
assign c7243 =  x512 &  x539 &  x567 & ~x27 & ~x46 & ~x57 & ~x98 & ~x126 & ~x423 & ~x448;
assign c7245 = ~x59 & ~x91 & ~x109 & ~x137 & ~x162 & ~x167 & ~x250 & ~x306 & ~x333 & ~x365 & ~x366 & ~x369 & ~x387 & ~x389 & ~x392 & ~x394 & ~x413 & ~x425 & ~x443 & ~x444 & ~x480 & ~x507 & ~x583 & ~x647 & ~x676 & ~x752;
assign c7247 =  x433 & ~x43 & ~x155 & ~x265 & ~x266;
assign c7249 =  x314 &  x498 &  x553;
assign c7251 =  x549 & ~x263 & ~x290 & ~x446;
assign c7253 =  x539 &  x566 & ~x29 & ~x167 & ~x296 & ~x351;
assign c7255 = ~x0 & ~x9 & ~x25 & ~x33 & ~x61 & ~x86 & ~x110 & ~x113 & ~x144 & ~x145 & ~x194 & ~x306 & ~x364 & ~x365 & ~x368 & ~x393 & ~x396 & ~x423 & ~x478 & ~x490 & ~x505 & ~x729 & ~x753;
assign c7257 =  x464 & ~x80 & ~x81 & ~x109 & ~x169 & ~x309 & ~x337 & ~x361 & ~x390 & ~x419 & ~x450 & ~x478 & ~x536 & ~x555 & ~x615 & ~x646 & ~x674 & ~x755;
assign c7259 =  x622 &  x623 &  x624;
assign c7261 =  x482 &  x509 &  x537 & ~x24 & ~x52 & ~x77 & ~x111 & ~x193 & ~x195 & ~x279 & ~x660 & ~x731 & ~x738 & ~x740;
assign c7263 =  x445 & ~x26 & ~x46 & ~x515;
assign c7265 =  x745 &  x746 &  x773 & ~x50 & ~x281 & ~x306 & ~x334;
assign c7267 = ~x212 & ~x213 & ~x214 & ~x237 & ~x239 & ~x265 & ~x266 & ~x296 & ~x394;
assign c7269 =  x623 &  x624 &  x625 & ~x23 & ~x165 & ~x251 & ~x450 & ~x731 & ~x757;
assign c7271 = ~x3 & ~x33 & ~x54 & ~x88 & ~x113 & ~x191 & ~x256 & ~x258 & ~x306 & ~x312 & ~x396 & ~x401 & ~x451 & ~x500 & ~x611 & ~x664 & ~x671 & ~x752;
assign c7273 =  x687 &  x715 & ~x54 & ~x195 & ~x280 & ~x311 & ~x333 & ~x334 & ~x335 & ~x386 & ~x424 & ~x448 & ~x504 & ~x528 & ~x609 & ~x674 & ~x704 & ~x783;
assign c7275 = ~x9 & ~x12 & ~x39 & ~x110 & ~x168 & ~x297 & ~x325 & ~x352 & ~x355 & ~x392 & ~x504 & ~x670;
assign c7277 =  x347 & ~x166 & ~x195 & ~x219 & ~x253 & ~x275 & ~x334 & ~x385 & ~x389 & ~x416 & ~x424 & ~x445 & ~x468 & ~x757;
assign c7279 =  x715 & ~x167 & ~x189 & ~x195 & ~x248 & ~x304 & ~x393 & ~x421 & ~x470 & ~x471 & ~x472 & ~x496 & ~x533 & ~x585 & ~x636 & ~x669 & ~x730;
assign c7281 =  x285;
assign c7283 =  x566 &  x593 &  x594 &  x621 &  x622 &  x649 & ~x644 & ~x768;
assign c7285 = ~x13 & ~x33 & ~x82 & ~x320 & ~x349 & ~x378 & ~x405 & ~x431 & ~x458 & ~x542 & ~x596 & ~x651;
assign c7287 = ~x5 & ~x28 & ~x31 & ~x141 & ~x206 & ~x235 & ~x277 & ~x303 & ~x333 & ~x360 & ~x388 & ~x476 & ~x500 & ~x532;
assign c7289 =  x295 & ~x5 & ~x144 & ~x165 & ~x283 & ~x333 & ~x334 & ~x340 & ~x390 & ~x393 & ~x469 & ~x483 & ~x526 & ~x564 & ~x618 & ~x665 & ~x668;
assign c7291 =  x509 & ~x52 & ~x98 & ~x297 & ~x717 & ~x728 & ~x745;
assign c7293 =  x466 & ~x139 & ~x262 & ~x263 & ~x362 & ~x390 & ~x446 & ~x780;
assign c7295 =  x581 &  x608 &  x609 &  x610 &  x637;
assign c7297 =  x265 & ~x20 & ~x224 & ~x247 & ~x252 & ~x255 & ~x283 & ~x304 & ~x305 & ~x307 & ~x314 & ~x391 & ~x445 & ~x476 & ~x499 & ~x503 & ~x562 & ~x613 & ~x616 & ~x662 & ~x671;
assign c7299 =  x539 &  x566 &  x567 &  x594 &  x595 & ~x353;
assign c7301 =  x445 & ~x412 & ~x439 & ~x464 & ~x518;
assign c7303 = ~x106 & ~x167 & ~x199 & ~x216 & ~x230 & ~x277 & ~x304 & ~x365 & ~x392 & ~x419 & ~x538 & ~x560 & ~x702;
assign c7305 =  x468 &  x524 &  x576;
assign c7307 =  x205 & ~x0 & ~x13 & ~x15 & ~x101 & ~x111 & ~x155 & ~x156 & ~x237 & ~x266 & ~x365 & ~x670 & ~x722 & ~x729;
assign c7309 = ~x137 & ~x151 & ~x180 & ~x372;
assign c7311 = ~x7 & ~x195 & ~x296 & ~x349 & ~x376 & ~x404 & ~x430 & ~x698 & ~x737;
assign c7313 =  x742 &  x769 &  x770 & ~x84 & ~x107 & ~x113 & ~x306 & ~x577;
assign c7315 =  x687 & ~x81 & ~x112 & ~x137 & ~x142 & ~x170 & ~x274 & ~x275 & ~x304 & ~x331 & ~x332 & ~x333 & ~x387 & ~x502 & ~x585 & ~x617 & ~x669 & ~x670;
assign c7317 =  x576 &  x603 & ~x82 & ~x373 & ~x374 & ~x401;
assign c7319 =  x694 & ~x261;
assign c7321 =  x568 &  x595 &  x596 &  x597 &  x623 &  x624;
assign c7323 =  x539 & ~x297 & ~x353 & ~x367 & ~x448;
assign c7325 =  x567 &  x595 & ~x168 & ~x373;
assign c7327 = ~x13 & ~x293 & ~x319 & ~x345 & ~x346 & ~x347 & ~x371 & ~x372 & ~x373 & ~x400 & ~x401;
assign c7329 =  x433 &  x461 &  x488 &  x489 & ~x30 & ~x45 & ~x195;
assign c7331 =  x432 & ~x46 & ~x105 & ~x239 & ~x439 & ~x470 & ~x522;
assign c7333 =  x567 &  x568 &  x595 &  x596 & ~x5 & ~x20 & ~x101;
assign c7335 = ~x26 & ~x133 & ~x162 & ~x221 & ~x250 & ~x280 & ~x284 & ~x305 & ~x366 & ~x369 & ~x384 & ~x398 & ~x412 & ~x446 & ~x453 & ~x474 & ~x508 & ~x694;
assign c7337 = ~x1 & ~x54 & ~x349 & ~x376 & ~x378 & ~x404 & ~x430 & ~x431 & ~x488 & ~x515 & ~x541 & ~x651 & ~x736;
assign c7339 =  x717 &  x744 & ~x28 & ~x79 & ~x110 & ~x111 & ~x167 & ~x168 & ~x192 & ~x193 & ~x197 & ~x249 & ~x255 & ~x391 & ~x421 & ~x557 & ~x559 & ~x560 & ~x640 & ~x645 & ~x752;
assign c7341 =  x127 &  x155 &  x183 &  x295;
assign c7343 = ~x31 & ~x90 & ~x229 & ~x245 & ~x283 & ~x306 & ~x338 & ~x367 & ~x387 & ~x388 & ~x424 & ~x446 & ~x479 & ~x499 & ~x507 & ~x581 & ~x651 & ~x677 & ~x697;
assign c7345 =  x713 &  x714 &  x740 &  x741 & ~x79 & ~x104 & ~x137 & ~x164 & ~x165 & ~x307 & ~x419 & ~x446 & ~x448 & ~x673 & ~x726 & ~x758 & ~x783;
assign c7347 = ~x48 & ~x353 & ~x439 & ~x632;
assign c7349 =  x406 &  x433 &  x461 & ~x16 & ~x76 & ~x211 & ~x212 & ~x615 & ~x633;
assign c7351 = ~x126 & ~x154 & ~x159 & ~x213 & ~x237 & ~x239 & ~x266 & ~x505 & ~x524 & ~x617;
assign c7353 =  x537 & ~x2 & ~x23 & ~x46 & ~x56 & ~x167 & ~x295 & ~x298 & ~x552 & ~x588;
assign c7355 = ~x2 & ~x21 & ~x28 & ~x59 & ~x107 & ~x112 & ~x197 & ~x199 & ~x221 & ~x245 & ~x254 & ~x275 & ~x282 & ~x301 & ~x306 & ~x359 & ~x361 & ~x365 & ~x367 & ~x390 & ~x394 & ~x416 & ~x419 & ~x420 & ~x424 & ~x472 & ~x473 & ~x477 & ~x506 & ~x587 & ~x664 & ~x674 & ~x699 & ~x700 & ~x705 & ~x723 & ~x750 & ~x758 & ~x759 & ~x760;
assign c7357 =  x228 & ~x236 & ~x336 & ~x742 & ~x778;
assign c7359 = ~x3 & ~x109 & ~x146 & ~x168 & ~x378 & ~x404 & ~x464 & ~x487 & ~x520 & ~x546 & ~x624 & ~x670 & ~x708 & ~x750;
assign c7361 =  x507 & ~x151 & ~x377 & ~x683;
assign c7363 =  x155 &  x183 & ~x23 & ~x168 & ~x196 & ~x247 & ~x252 & ~x302 & ~x304 & ~x309 & ~x334 & ~x361 & ~x391 & ~x420 & ~x449 & ~x476 & ~x530 & ~x617;
assign c7365 =  x482 & ~x14 & ~x23 & ~x31 & ~x294 & ~x295 & ~x297 & ~x323 & ~x394 & ~x767;
assign c7367 = ~x8 & ~x37 & ~x84 & ~x169 & ~x328 & ~x349 & ~x375 & ~x376 & ~x378 & ~x404 & ~x405 & ~x430 & ~x431 & ~x460;
assign c7369 =  x606 &  x633 & ~x27 & ~x319 & ~x347;
assign c7371 =  x524 &  x581 &  x610;
assign c7373 =  x549 &  x575 &  x576 &  x603 &  x630;
assign c7375 = ~x67 & ~x319 & ~x320 & ~x347 & ~x348 & ~x349 & ~x374 & ~x430 & ~x431 & ~x485;
assign c7377 =  x687 & ~x30 & ~x55 & ~x75 & ~x79 & ~x135 & ~x195 & ~x362 & ~x391 & ~x418 & ~x419 & ~x499 & ~x552 & ~x556 & ~x580 & ~x610 & ~x729 & ~x752 & ~x759 & ~x782;
assign c7379 =  x295 & ~x316 & ~x317 & ~x344 & ~x345 & ~x371 & ~x372 & ~x399 & ~x400;
assign c7381 = ~x151 & ~x179 & ~x187 & ~x208 & ~x237 & ~x496 & ~x651;
assign c7383 =  x630 &  x631 &  x632 &  x657 &  x658 & ~x166 & ~x418 & ~x439 & ~x530 & ~x589;
assign c7385 =  x369 & ~x29 & ~x61 & ~x167 & ~x404 & ~x432 & ~x489 & ~x542 & ~x707;
assign c7387 =  x434 &  x461 & ~x239;
assign c7389 =  x461 &  x462 &  x489 &  x568 & ~x32 & ~x50 & ~x75 & ~x761 & ~x780;
assign c7391 = ~x50 & ~x62 & ~x110 & ~x111 & ~x139 & ~x195 & ~x197 & ~x224 & ~x338 & ~x368 & ~x369 & ~x387 & ~x391 & ~x398 & ~x412 & ~x420 & ~x421 & ~x472 & ~x529 & ~x583 & ~x597 & ~x608 & ~x669 & ~x671 & ~x723;
assign c7393 =  x551 &  x578 &  x605 &  x606 &  x632;
assign c7395 =  x676 &  x677 &  x704;
assign c7397 =  x684 &  x685 &  x686 & ~x195 & ~x360 & ~x361 & ~x387 & ~x469 & ~x673;
assign c7399 =  x183 &  x347 & ~x30 & ~x51 & ~x139 & ~x141 & ~x200 & ~x221 & ~x255 & ~x307 & ~x362 & ~x390 & ~x396 & ~x421 & ~x422 & ~x448 & ~x729;
assign c7401 =  x501 & ~x438 & ~x439 & ~x464 & ~x490 & ~x517 & ~x573 & ~x629;
assign c7403 = ~x23 & ~x50 & ~x78 & ~x108 & ~x111 & ~x135 & ~x162 & ~x169 & ~x194 & ~x230 & ~x247 & ~x277 & ~x281 & ~x306 & ~x334 & ~x335 & ~x339 & ~x359 & ~x361 & ~x362 & ~x367 & ~x370 & ~x415 & ~x476 & ~x512 & ~x536 & ~x582 & ~x584 & ~x641 & ~x645 & ~x665 & ~x699 & ~x756;
assign c7405 = ~x0 & ~x2 & ~x22 & ~x30 & ~x35 & ~x48 & ~x53 & ~x101 & ~x102 & ~x141 & ~x182 & ~x195 & ~x345 & ~x346 & ~x372 & ~x373 & ~x400 & ~x401 & ~x429 & ~x587 & ~x643 & ~x673 & ~x730 & ~x763;
assign c7407 =  x340 &  x582;
assign c7409 =  x332 &  x360 & ~x357 & ~x439;
assign c7411 =  x595 & ~x399;
assign c7413 =  x230 & ~x151 & ~x180 & ~x208;
assign c7415 =  x383 &  x384 &  x439 & ~x21 & ~x53 & ~x54 & ~x79 & ~x107 & ~x135 & ~x136 & ~x140 & ~x251 & ~x281 & ~x418 & ~x446 & ~x642 & ~x672 & ~x754 & ~x756;
assign c7417 = ~x51 & ~x320 & ~x346 & ~x347 & ~x373 & ~x376 & ~x399 & ~x400 & ~x427 & ~x428 & ~x482;
assign c7419 =  x529 & ~x546;
assign c7421 =  x146 &  x174 & ~x97 & ~x123 & ~x151 & ~x167;
assign c7423 = ~x3 & ~x8 & ~x27 & ~x55 & ~x56 & ~x58 & ~x74 & ~x172 & ~x247 & ~x304 & ~x306 & ~x361 & ~x389 & ~x401 & ~x614 & ~x636 & ~x642 & ~x698 & ~x758;
assign c7425 = ~x52 & ~x99 & ~x127 & ~x128 & ~x155 & ~x184 & ~x211 & ~x212 & ~x239 & ~x267 & ~x393 & ~x468 & ~x551 & ~x648 & ~x667 & ~x759;
assign c7427 =  x41 & ~x32 & ~x57 & ~x79 & ~x107 & ~x247 & ~x284 & ~x306 & ~x362 & ~x475 & ~x643;
assign c7429 =  x482 & ~x151 & ~x179 & ~x206 & ~x421;
assign c7431 =  x498 &  x526 &  x554 & ~x630 & ~x760;
assign c7433 = ~x166 & ~x167 & ~x302 & ~x304 & ~x307 & ~x340 & ~x341 & ~x387 & ~x396 & ~x422 & ~x424 & ~x446 & ~x449 & ~x471 & ~x476 & ~x564 & ~x595 & ~x619 & ~x700 & ~x762;
assign c7435 =  x629 &  x630 &  x657 & ~x15 & ~x110 & ~x360 & ~x362 & ~x387 & ~x388 & ~x412 & ~x471 & ~x502 & ~x644 & ~x732;
assign c7437 =  x553 &  x581 &  x609 & ~x28 & ~x52 & ~x767;
assign c7439 =  x555 & ~x434;
assign c7441 =  x584 &  x611 &  x612;
assign c7443 = ~x59 & ~x109 & ~x189 & ~x257 & ~x273 & ~x276 & ~x304 & ~x308 & ~x332 & ~x336 & ~x358 & ~x359 & ~x369 & ~x386 & ~x387 & ~x394 & ~x416 & ~x424 & ~x504 & ~x554 & ~x563 & ~x587 & ~x637 & ~x774;
assign c7445 = ~x235 & ~x236 & ~x263 & ~x264 & ~x290 & ~x318 & ~x393 & ~x417;
assign c7447 =  x582 & ~x487 & ~x559;
assign c7449 =  x409 &  x464 & ~x25 & ~x52 & ~x56 & ~x280 & ~x281 & ~x307 & ~x363 & ~x387 & ~x390 & ~x473 & ~x474 & ~x501 & ~x502 & ~x532 & ~x552 & ~x557 & ~x560 & ~x561 & ~x612 & ~x696 & ~x697 & ~x708 & ~x760 & ~x777;
assign c7451 =  x117 & ~x64 & ~x644;
assign c7453 = ~x67 & ~x154 & ~x208 & ~x236 & ~x264 & ~x265;
assign c7455 =  x432 &  x433 & ~x21 & ~x80 & ~x131 & ~x134 & ~x213 & ~x241 & ~x422 & ~x474 & ~x476 & ~x530 & ~x559 & ~x669 & ~x672 & ~x675 & ~x700 & ~x702 & ~x703 & ~x733;
assign c7457 =  x295 & ~x55 & ~x218 & ~x247 & ~x275 & ~x308 & ~x334 & ~x387 & ~x388 & ~x446 & ~x452;
assign c7459 =  x229 &  x537;
assign c7461 = ~x64 & ~x183 & ~x211 & ~x213 & ~x239 & ~x241 & ~x267 & ~x271 & ~x295 & ~x297 & ~x323;
assign c7463 =  x536 &  x592 & ~x27 & ~x55 & ~x689 & ~x783;
assign c7465 = ~x58 & ~x137 & ~x297 & ~x405 & ~x432 & ~x436 & ~x459 & ~x488 & ~x570 & ~x677 & ~x727;
assign c7467 =  x745 &  x746 &  x772 & ~x50 & ~x165 & ~x308 & ~x419 & ~x727 & ~x783;
assign c7469 =  x575 & ~x167 & ~x290 & ~x317 & ~x344 & ~x345 & ~x371 & ~x373 & ~x398 & ~x400 & ~x427;
assign c7471 =  x651 &  x652 & ~x3 & ~x30 & ~x53 & ~x166 & ~x281 & ~x420 & ~x484 & ~x668 & ~x703;
assign c7473 =  x501 & ~x35 & ~x353 & ~x383 & ~x411;
assign c7475 =  x706 &  x709;
assign c7477 = ~x156 & ~x237 & ~x265 & ~x292 & ~x293 & ~x320 & ~x694;
assign c7479 =  x332 &  x360 & ~x239 & ~x296;
assign c7481 =  x127 &  x155 & ~x55 & ~x243 & ~x281 & ~x304 & ~x503 & ~x504 & ~x615 & ~x672;
assign c7483 = ~x23 & ~x24 & ~x28 & ~x49 & ~x51 & ~x79 & ~x83 & ~x111 & ~x165 & ~x246 & ~x275 & ~x328 & ~x360 & ~x369 & ~x386 & ~x387 & ~x390 & ~x424 & ~x526;
assign c7485 = ~x57 & ~x265 & ~x292 & ~x320 & ~x347 & ~x348 & ~x349 & ~x375 & ~x376 & ~x405 & ~x431 & ~x707;
assign c7487 = ~x304 & ~x306 & ~x343 & ~x367 & ~x439 & ~x539 & ~x700;
assign c7489 =  x468 &  x496 &  x523 &  x524 &  x551 & ~x445;
assign c7491 =  x293 & ~x60 & ~x190 & ~x274 & ~x337 & ~x390 & ~x398 & ~x424 & ~x445 & ~x587 & ~x642 & ~x780;
assign c7493 =  x596 &  x624 &  x625 & ~x20 & ~x21 & ~x24 & ~x29 & ~x79 & ~x140 & ~x168 & ~x393 & ~x421 & ~x702 & ~x727;
assign c7495 = ~x15 & ~x24 & ~x351 & ~x378 & ~x404 & ~x405 & ~x407 & ~x431 & ~x459 & ~x464 & ~x513 & ~x601 & ~x760;
assign c7497 =  x42 &  x70 & ~x0 & ~x31 & ~x33 & ~x50 & ~x57 & ~x58 & ~x85 & ~x113 & ~x137 & ~x170 & ~x194 & ~x221 & ~x224 & ~x225 & ~x249 & ~x281 & ~x304 & ~x339 & ~x420 & ~x443 & ~x445 & ~x446 & ~x474 & ~x528 & ~x529 & ~x530 & ~x586 & ~x587 & ~x620 & ~x672;
assign c7499 =  x304 &  x388 & ~x464;
assign c80 =  x455 &  x511 &  x624 & ~x172 & ~x490 & ~x572;
assign c82 =  x454 &  x593 & ~x42 & ~x46 & ~x88 & ~x199 & ~x284 & ~x518;
assign c84 =  x373 &  x652 & ~x31 & ~x53 & ~x58 & ~x60 & ~x61 & ~x82 & ~x89 & ~x141 & ~x144 & ~x145 & ~x281 & ~x335 & ~x364 & ~x392 & ~x518 & ~x519 & ~x545 & ~x546 & ~x576;
assign c86 =  x618 &  x645 & ~x408;
assign c88 = ~x86 & ~x125 & ~x151 & ~x206 & ~x275 & ~x299 & ~x319 & ~x623;
assign c810 =  x738 &  x744 & ~x398 & ~x481 & ~x497 & ~x606;
assign c812 =  x462 &  x463 &  x488 &  x689 & ~x164 & ~x329 & ~x342 & ~x415 & ~x496 & ~x499;
assign c814 =  x378 &  x406 & ~x369 & ~x519 & ~x572;
assign c816 =  x320 &  x347 & ~x2 & ~x26 & ~x31 & ~x83 & ~x90 & ~x146 & ~x162 & ~x199 & ~x278 & ~x337 & ~x519 & ~x546 & ~x571 & ~x573;
assign c818 =  x497 & ~x21 & ~x100 & ~x115 & ~x325 & ~x353 & ~x354 & ~x389 & ~x491 & ~x519 & ~x578;
assign c820 =  x322 &  x350 &  x462 & ~x1 & ~x57 & ~x90 & ~x198 & ~x221 & ~x327 & ~x328 & ~x329 & ~x336 & ~x440 & ~x578 & ~x606;
assign c822 =  x452 &  x505 & ~x332 & ~x362 & ~x487 & ~x780;
assign c824 =  x378 &  x687 &  x689 & ~x172 & ~x201 & ~x217 & ~x424;
assign c826 =  x14 &  x404 &  x431 &  x459;
assign c828 =  x397 & ~x29 & ~x135 & ~x306 & ~x331 & ~x358 & ~x487 & ~x488 & ~x653 & ~x667;
assign c830 = ~x3 & ~x4 & ~x6 & ~x28 & ~x56 & ~x111 & ~x224 & ~x253 & ~x325 & ~x332 & ~x363 & ~x379 & ~x381 & ~x397 & ~x449 & ~x476 & ~x491 & ~x546 & ~x559 & ~x704 & ~x745;
assign c832 = ~x37 & ~x147 & ~x175 & ~x225 & ~x231 & ~x254 & ~x336 & ~x342 & ~x371 & ~x416 & ~x518 & ~x530 & ~x546 & ~x587 & ~x615 & ~x671 & ~x713 & ~x733 & ~x774;
assign c834 =  x480 &  x505 & ~x461;
assign c836 =  x479 & ~x50 & ~x75 & ~x275 & ~x350 & ~x362 & ~x446 & ~x471 & ~x708;
assign c838 =  x546 &  x739 &  x743 & ~x370 & ~x400 & ~x443;
assign c840 =  x511 & ~x109 & ~x195 & ~x280 & ~x311 & ~x337 & ~x340 & ~x385 & ~x470 & ~x519 & ~x546 & ~x571 & ~x572 & ~x682;
assign c842 =  x537 &  x565 & ~x1 & ~x87 & ~x128 & ~x199 & ~x655 & ~x729;
assign c844 =  x746 & ~x685;
assign c846 =  x399 &  x455 &  x511 &  x623 &  x679 & ~x570;
assign c848 =  x767 & ~x497;
assign c850 =  x540 &  x680 & ~x8 & ~x34 & ~x89 & ~x118 & ~x146 & ~x312 & ~x452 & ~x732;
assign c852 =  x15 &  x431 & ~x24 & ~x138 & ~x144 & ~x256 & ~x258 & ~x367 & ~x695 & ~x782;
assign c854 =  x428 &  x619 & ~x451 & ~x475 & ~x505 & ~x729;
assign c856 =  x376 & ~x3 & ~x81 & ~x116 & ~x175 & ~x197 & ~x199 & ~x252 & ~x253 & ~x367 & ~x395 & ~x437 & ~x547 & ~x548 & ~x576 & ~x760;
assign c858 =  x407 &  x435 & ~x14 & ~x77 & ~x189 & ~x274 & ~x334 & ~x355 & ~x710 & ~x769;
assign c860 =  x376 &  x462 & ~x21 & ~x84 & ~x109 & ~x112 & ~x175 & ~x253 & ~x259 & ~x284 & ~x357 & ~x369 & ~x399 & ~x413 & ~x483 & ~x496 & ~x498 & ~x553 & ~x615 & ~x724 & ~x728;
assign c862 =  x377 & ~x119 & ~x287 & ~x371 & ~x505 & ~x521 & ~x544 & ~x546 & ~x615;
assign c864 =  x397 &  x453 &  x481 &  x509 &  x593 &  x621 &  x649 & ~x162 & ~x199 & ~x487 & ~x757;
assign c866 =  x406 & ~x339 & ~x383 & ~x682;
assign c868 =  x351 &  x459 &  x463;
assign c870 =  x240 &  x436 &  x744 & ~x22 & ~x110 & ~x229 & ~x444 & ~x473 & ~x551 & ~x587;
assign c872 =  x245 &  x273 &  x329 &  x413 & ~x256;
assign c874 =  x14 &  x42 &  x459 & ~x194 & ~x256 & ~x259 & ~x286 & ~x336 & ~x363 & ~x370 & ~x468 & ~x782;
assign c876 =  x511 &  x735;
assign c878 =  x187 &  x215 &  x271 &  x439;
assign c880 =  x545 &  x743 & ~x121 & ~x659;
assign c882 =  x710 &  x716 &  x717 & ~x60 & ~x106 & ~x173 & ~x175 & ~x253 & ~x257 & ~x286 & ~x387 & ~x440 & ~x528 & ~x591 & ~x701 & ~x727 & ~x758;
assign c884 =  x457 &  x597 & ~x8 & ~x88 & ~x169 & ~x202 & ~x223 & ~x225 & ~x226 & ~x229 & ~x230 & ~x277 & ~x338 & ~x365 & ~x369 & ~x394 & ~x447 & ~x734;
assign c886 =  x453 &  x507 & ~x10 & ~x28 & ~x29 & ~x50 & ~x88 & ~x106 & ~x193 & ~x254 & ~x324 & ~x407 & ~x408 & ~x435 & ~x519;
assign c888 =  x548 &  x744 & ~x553 & ~x578;
assign c890 =  x425 &  x533 & ~x135 & ~x433;
assign c892 = ~x22 & ~x26 & ~x33 & ~x37 & ~x45 & ~x57 & ~x71 & ~x81 & ~x82 & ~x98 & ~x99 & ~x100 & ~x127 & ~x128 & ~x138 & ~x156 & ~x164 & ~x195 & ~x304 & ~x335 & ~x405 & ~x656 & ~x684 & ~x696 & ~x711 & ~x744 & ~x759 & ~x760 & ~x778;
assign c894 =  x423 & ~x618;
assign c896 = ~x36 & ~x64 & ~x109 & ~x129 & ~x163 & ~x275 & ~x362 & ~x545 & ~x546 & ~x669 & ~x679 & ~x684 & ~x685 & ~x711 & ~x718 & ~x741 & ~x769;
assign c898 =  x720 &  x721 & ~x4 & ~x111 & ~x302 & ~x303 & ~x359 & ~x362 & ~x392 & ~x498 & ~x610 & ~x632 & ~x640;
assign c8100 =  x378 &  x406 &  x688 & ~x175 & ~x498;
assign c8102 =  x457 &  x736 & ~x31 & ~x335 & ~x336 & ~x471;
assign c8104 =  x349 &  x377 & ~x4 & ~x314 & ~x343 & ~x369 & ~x478 & ~x534 & ~x550 & ~x573;
assign c8106 =  x347 &  x374 & ~x50 & ~x54 & ~x113 & ~x258 & ~x341 & ~x393 & ~x472 & ~x504 & ~x519 & ~x726 & ~x748;
assign c8108 =  x374 &  x681 & ~x9 & ~x145 & ~x546 & ~x548;
assign c8110 =  x128 &  x156 &  x212 &  x352 &  x436 & ~x52 & ~x109 & ~x202 & ~x230 & ~x329 & ~x331 & ~x674 & ~x698;
assign c8112 =  x455 &  x482 &  x483 & ~x0 & ~x29 & ~x30 & ~x91 & ~x195 & ~x222 & ~x225 & ~x336 & ~x435 & ~x463 & ~x517;
assign c8114 = ~x5 & ~x8 & ~x19 & ~x64 & ~x92 & ~x172 & ~x202 & ~x222 & ~x229 & ~x254 & ~x287 & ~x342 & ~x369 & ~x408 & ~x417 & ~x418 & ~x436 & ~x445 & ~x491 & ~x576 & ~x728;
assign c8116 =  x373 & ~x46 & ~x57 & ~x109 & ~x199 & ~x285 & ~x307 & ~x337 & ~x365 & ~x490 & ~x519 & ~x546 & ~x573 & ~x576;
assign c8118 =  x152 &  x376 & ~x121 & ~x205 & ~x259 & ~x717;
assign c8120 =  x403 &  x653 & ~x111 & ~x231 & ~x259 & ~x283 & ~x371 & ~x427;
assign c8122 =  x481 &  x536 & ~x50 & ~x71 & ~x78 & ~x105 & ~x107 & ~x108 & ~x143 & ~x167 & ~x192 & ~x336 & ~x359 & ~x361 & ~x680;
assign c8124 =  x152 & ~x178 & ~x261 & ~x287 & ~x289 & ~x369 & ~x523;
assign c8126 =  x520 &  x544 &  x546;
assign c8128 =  x452 &  x533 & ~x402 & ~x432 & ~x751;
assign c8130 =  x351 &  x433 &  x626 & ~x118 & ~x536 & ~x564 & ~x668;
assign c8132 =  x157 &  x185 &  x213 &  x270 &  x297 &  x298 & ~x145 & ~x163 & ~x254;
assign c8134 =  x295 &  x407 &  x435 &  x463 &  x489 & ~x31 & ~x57 & ~x133 & ~x277 & ~x415 & ~x440 & ~x449 & ~x471 & ~x497 & ~x667;
assign c8136 =  x185 &  x297 &  x353 & ~x24 & ~x53 & ~x77 & ~x220 & ~x604 & ~x780;
assign c8138 =  x481 &  x508 &  x509 &  x524 & ~x416 & ~x435;
assign c8140 = ~x39 & ~x41 & ~x43 & ~x70 & ~x72 & ~x78 & ~x111 & ~x125 & ~x135 & ~x136 & ~x137 & ~x152 & ~x159 & ~x163 & ~x189 & ~x194 & ~x219 & ~x220 & ~x224 & ~x247 & ~x250 & ~x348 & ~x357 & ~x363 & ~x386 & ~x432 & ~x433 & ~x474 & ~x488 & ~x573 & ~x710 & ~x738 & ~x779;
assign c8142 =  x505 & ~x589;
assign c8144 =  x406 & ~x32 & ~x341 & ~x398 & ~x479 & ~x491 & ~x543 & ~x546;
assign c8146 =  x151 &  x351 &  x430;
assign c8148 =  x511 & ~x25 & ~x52 & ~x53 & ~x89 & ~x110 & ~x170 & ~x194 & ~x257 & ~x369 & ~x532 & ~x691 & ~x727;
assign c8150 = ~x2 & ~x13 & ~x41 & ~x46 & ~x49 & ~x50 & ~x117 & ~x217 & ~x226 & ~x277 & ~x322 & ~x360 & ~x386 & ~x402 & ~x433 & ~x458 & ~x707 & ~x771;
assign c8152 =  x401 &  x457 &  x652 & ~x145;
assign c8154 =  x15 &  x404 & ~x32 & ~x83 & ~x163 & ~x170 & ~x310 & ~x343 & ~x501;
assign c8156 =  x484 & ~x198 & ~x340 & ~x369 & ~x435 & ~x491 & ~x504 & ~x519 & ~x546 & ~x572 & ~x573 & ~x684 & ~x734 & ~x768;
assign c8158 =  x351 &  x352 &  x436 &  x491 & ~x219;
assign c8160 =  x452 &  x561 & ~x197 & ~x220 & ~x222 & ~x363 & ~x389 & ~x394 & ~x416 & ~x419 & ~x475;
assign c8162 =  x351 &  x463 &  x491 & ~x576;
assign c8164 =  x459 &  x491 &  x681;
assign c8166 =  x151 &  x375 & ~x22 & ~x54 & ~x62 & ~x63 & ~x107 & ~x196 & ~x342 & ~x397 & ~x398 & ~x419 & ~x575 & ~x587 & ~x778;
assign c8168 =  x344 &  x428 &  x484 &  x568 & ~x109 & ~x114 & ~x462 & ~x546;
assign c8170 =  x480 &  x507 &  x534 & ~x21 & ~x435 & ~x518 & ~x546;
assign c8172 =  x423 & ~x66 & ~x75 & ~x94 & ~x161 & ~x165 & ~x220 & ~x247 & ~x331 & ~x333 & ~x376;
assign c8174 =  x537 & ~x43 & ~x142 & ~x361 & ~x413 & ~x441 & ~x546 & ~x771;
assign c8176 =  x245 &  x273 &  x329 & ~x271;
assign c8178 =  x507 &  x621 & ~x404;
assign c8180 =  x455 &  x511 & ~x82 & ~x113 & ~x138 & ~x196 & ~x220 & ~x388 & ~x389 & ~x422 & ~x516 & ~x517 & ~x518 & ~x543 & ~x549 & ~x725 & ~x727 & ~x783;
assign c8182 =  x534 & ~x14 & ~x135 & ~x163 & ~x387 & ~x488 & ~x694;
assign c8184 =  x451 & ~x3 & ~x14 & ~x135 & ~x162 & ~x192 & ~x275 & ~x308 & ~x334 & ~x377 & ~x385 & ~x405 & ~x462 & ~x488;
assign c8186 =  x431 &  x458 & ~x26 & ~x51 & ~x60 & ~x88 & ~x102 & ~x109 & ~x171 & ~x172 & ~x252 & ~x259 & ~x273 & ~x284 & ~x302 & ~x308 & ~x369 & ~x396 & ~x414 & ~x420 & ~x427 & ~x443 & ~x496 & ~x503 & ~x532 & ~x586 & ~x640 & ~x642 & ~x646 & ~x647 & ~x667 & ~x752 & ~x781 & ~x782;
assign c8188 =  x351 &  x435 &  x488 & ~x23 & ~x25 & ~x60 & ~x165 & ~x259 & ~x341 & ~x367 & ~x427 & ~x498 & ~x503 & ~x507 & ~x524 & ~x565 & ~x702;
assign c8190 =  x398 &  x509 &  x510 &  x594 &  x622 & ~x487;
assign c8192 =  x239 &  x351 &  x375 &  x435 &  x487 & ~x453 & ~x471;
assign c8194 =  x128 &  x240 &  x380 &  x408 &  x436 & ~x50 & ~x275 & ~x360 & ~x603 & ~x604;
assign c8196 =  x322 &  x378 &  x406 &  x434 & ~x3 & ~x88 & ~x184 & ~x189 & ~x215 & ~x226 & ~x241 & ~x244 & ~x355 & ~x474;
assign c8198 =  x403 &  x431 &  x626 & ~x1 & ~x361 & ~x396 & ~x397 & ~x427 & ~x643;
assign c8200 =  x207 &  x375 &  x431 & ~x2 & ~x24 & ~x52 & ~x75 & ~x91 & ~x110 & ~x136 & ~x142 & ~x144 & ~x167 & ~x174 & ~x226 & ~x232 & ~x233 & ~x258 & ~x260 & ~x288 & ~x336 & ~x338 & ~x365 & ~x418 & ~x445 & ~x447 & ~x449 & ~x473 & ~x502 & ~x530 & ~x756 & ~x781 & ~x783;
assign c8202 =  x373 &  x540 & ~x491 & ~x544 & ~x546;
assign c8204 =  x722 & ~x424 & ~x576;
assign c8206 = ~x29 & ~x38 & ~x45 & ~x48 & ~x53 & ~x87 & ~x88 & ~x89 & ~x109 & ~x141 & ~x143 & ~x174 & ~x222 & ~x227 & ~x255 & ~x259 & ~x278 & ~x283 & ~x286 & ~x335 & ~x339 & ~x362 & ~x364 & ~x369 & ~x394 & ~x436 & ~x475 & ~x477 & ~x491 & ~x504 & ~x519 & ~x520 & ~x546 & ~x547 & ~x548 & ~x615 & ~x746 & ~x759;
assign c8208 =  x407 & ~x75 & ~x180 & ~x381 & ~x382 & ~x555 & ~x684;
assign c8210 =  x322 &  x434 &  x741 & ~x685;
assign c8212 =  x477 & ~x375 & ~x456;
assign c8214 =  x403 &  x431 & ~x54 & ~x135 & ~x149 & ~x203 & ~x250 & ~x314 & ~x315 & ~x316 & ~x335 & ~x392 & ~x463 & ~x761 & ~x774;
assign c8216 =  x457 &  x679 & ~x397;
assign c8218 =  x215 &  x243 &  x411 & ~x491 & ~x519 & ~x547;
assign c8220 =  x619 & ~x20 & ~x53 & ~x87 & ~x108 & ~x118 & ~x138 & ~x199 & ~x396 & ~x435;
assign c8222 =  x720 & ~x57 & ~x115 & ~x144 & ~x163 & ~x195 & ~x275 & ~x336 & ~x396 & ~x604 & ~x605 & ~x606 & ~x634 & ~x657 & ~x698;
assign c8224 =  x402 &  x430 &  x458 & ~x0 & ~x5 & ~x7 & ~x29 & ~x33 & ~x35 & ~x59 & ~x83 & ~x85 & ~x117 & ~x139 & ~x147 & ~x167 & ~x195 & ~x203 & ~x223 & ~x225 & ~x250 & ~x256 & ~x341 & ~x367 & ~x369 & ~x421 & ~x443 & ~x533 & ~x548 & ~x752 & ~x782;
assign c8226 =  x185 &  x353 &  x409;
assign c8228 =  x512 &  x735 & ~x88 & ~x136 & ~x139 & ~x165 & ~x172;
assign c8230 =  x42 &  x322 &  x431 & ~x171 & ~x244;
assign c8232 =  x506 & ~x87 & ~x361 & ~x591;
assign c8234 =  x546 &  x710 &  x744 & ~x299 & ~x425;
assign c8236 =  x433 &  x434 &  x625 & ~x35 & ~x91 & ~x414 & ~x426 & ~x475 & ~x477;
assign c8238 =  x434 &  x461 & ~x59 & ~x191 & ~x274 & ~x278 & ~x286 & ~x328 & ~x339 & ~x343 & ~x364 & ~x400;
assign c8240 =  x320 &  x376 & ~x89 & ~x173 & ~x183 & ~x286 & ~x334 & ~x369 & ~x475 & ~x578 & ~x630;
assign c8242 =  x424 &  x452 &  x505 & ~x278 & ~x430 & ~x457;
assign c8244 =  x434 &  x739 &  x742 & ~x661;
assign c8246 =  x373 & ~x3 & ~x49 & ~x87 & ~x137 & ~x171 & ~x251 & ~x307 & ~x332 & ~x362 & ~x491 & ~x502 & ~x516 & ~x519 & ~x520 & ~x546 & ~x548 & ~x576 & ~x602 & ~x657 & ~x700 & ~x724 & ~x731 & ~x757 & ~x759 & ~x777 & ~x782;
assign c8248 =  x536 &  x563 &  x705;
assign c8250 = ~x43 & ~x104 & ~x163 & ~x274 & ~x277 & ~x328 & ~x544 & ~x684 & ~x687 & ~x712;
assign c8252 =  x324 &  x436 &  x461;
assign c8254 =  x453 &  x534 & ~x724;
assign c8256 = ~x21 & ~x43 & ~x72 & ~x189 & ~x282 & ~x328 & ~x546 & ~x686 & ~x707 & ~x715 & ~x726;
assign c8258 = ~x173 & ~x315 & ~x363 & ~x381 & ~x491 & ~x519 & ~x546 & ~x738 & ~x739 & ~x741;
assign c8260 =  x128 &  x296 &  x431 & ~x190 & ~x387 & ~x549;
assign c8262 =  x398 &  x534 & ~x81 & ~x88 & ~x141 & ~x226 & ~x252 & ~x335 & ~x433 & ~x749;
assign c8264 =  x218 &  x330;
assign c8266 = ~x299 & ~x571;
assign c8268 =  x509 &  x617 &  x622;
assign c8270 =  x536 & ~x1 & ~x25 & ~x75 & ~x107 & ~x131 & ~x248 & ~x417 & ~x431 & ~x460 & ~x470 & ~x573 & ~x764;
assign c8272 =  x351 &  x406 & ~x131 & ~x172 & ~x202 & ~x220 & ~x275 & ~x329 & ~x334 & ~x498 & ~x587 & ~x630 & ~x671;
assign c8274 =  x397 &  x561 & ~x166;
assign c8276 =  x564 &  x733;
assign c8278 =  x477 & ~x330 & ~x374 & ~x702;
assign c8280 =  x491 &  x544 & ~x160 & ~x162 & ~x174 & ~x190 & ~x248 & ~x255 & ~x281 & ~x342 & ~x386 & ~x398 & ~x497 & ~x501 & ~x524 & ~x535 & ~x554 & ~x559 & ~x565 & ~x579 & ~x670 & ~x724;
assign c8282 =  x342 & ~x14 & ~x41 & ~x132 & ~x245 & ~x374 & ~x388 & ~x706;
assign c8284 = ~x3 & ~x6 & ~x18 & ~x44 & ~x128 & ~x143 & ~x165 & ~x201 & ~x202 & ~x250 & ~x259 & ~x307 & ~x313 & ~x392 & ~x424 & ~x465 & ~x491 & ~x519;
assign c8286 = ~x3 & ~x14 & ~x18 & ~x36 & ~x72 & ~x218 & ~x355 & ~x360 & ~x461 & ~x691 & ~x694 & ~x706 & ~x740;
assign c8288 = ~x10 & ~x156 & ~x240 & ~x255 & ~x268 & ~x390 & ~x392 & ~x408 & ~x435 & ~x437 & ~x473 & ~x519 & ~x520 & ~x728 & ~x740;
assign c8290 =  x482 & ~x7 & ~x23 & ~x88 & ~x108 & ~x136 & ~x193 & ~x247 & ~x282 & ~x304 & ~x361 & ~x407 & ~x435 & ~x491 & ~x520 & ~x546 & ~x572 & ~x577 & ~x604 & ~x605 & ~x758 & ~x767 & ~x783;
assign c8292 =  x370 & ~x75 & ~x276 & ~x361 & ~x402 & ~x475 & ~x501 & ~x572 & ~x664 & ~x692;
assign c8294 = ~x41 & ~x47 & ~x101 & ~x178 & ~x206 & ~x253 & ~x275 & ~x344 & ~x552;
assign c8296 =  x368 & ~x14 & ~x47 & ~x97 & ~x126 & ~x162 & ~x328 & ~x337 & ~x487 & ~x599 & ~x616 & ~x769 & ~x773;
assign c8298 =  x127 &  x295 &  x407 &  x460 &  x461 & ~x80 & ~x116 & ~x302 & ~x328;
assign c8300 =  x99 &  x238 &  x322 &  x431 & ~x62 & ~x104 & ~x175 & ~x203 & ~x216 & ~x273 & ~x329 & ~x339 & ~x411 & ~x451 & ~x581;
assign c8302 =  x433 &  x654 & ~x62 & ~x206 & ~x283;
assign c8304 = ~x1 & ~x19 & ~x22 & ~x65 & ~x147 & ~x167 & ~x253 & ~x286 & ~x287 & ~x315 & ~x392 & ~x408 & ~x576 & ~x744;
assign c8306 =  x539 &  x567 & ~x2 & ~x26 & ~x32 & ~x47 & ~x49 & ~x79 & ~x99 & ~x166 & ~x174 & ~x225 & ~x283 & ~x335 & ~x337 & ~x390 & ~x422 & ~x518 & ~x544 & ~x738 & ~x779;
assign c8308 =  x427 &  x537 &  x623 & ~x515 & ~x546;
assign c8310 =  x428 &  x455 &  x456 & ~x172 & ~x255 & ~x366 & ~x436 & ~x462 & ~x518 & ~x546 & ~x571 & ~x572;
assign c8312 =  x397 &  x425 & ~x14 & ~x69 & ~x529;
assign c8314 =  x484 &  x652 & ~x109 & ~x519 & ~x544 & ~x572;
assign c8316 =  x315 &  x343 &  x344 &  x372 &  x455 &  x511 &  x539 &  x567 & ~x546;
assign c8318 =  x510 &  x592 &  x619 & ~x46 & ~x55 & ~x109 & ~x435 & ~x518 & ~x519 & ~x546;
assign c8320 =  x410 &  x564 & ~x84 & ~x163 & ~x222 & ~x336 & ~x435 & ~x519 & ~x547 & ~x548 & ~x576 & ~x772;
assign c8322 =  x397 & ~x141 & ~x275 & ~x304 & ~x376 & ~x458 & ~x460 & ~x546 & ~x702 & ~x707 & ~x716 & ~x735 & ~x739;
assign c8324 =  x484 &  x624 & ~x53 & ~x284 & ~x338 & ~x491 & ~x546 & ~x733 & ~x778 & ~x782;
assign c8326 =  x212 &  x240 &  x268 &  x380 &  x408 &  x436 & ~x30 & ~x85 & ~x109 & ~x279 & ~x310 & ~x578 & ~x604 & ~x613;
assign c8328 =  x739 &  x742 &  x743 &  x745 & ~x77 & ~x161 & ~x199 & ~x329 & ~x368 & ~x414 & ~x441 & ~x497 & ~x538 & ~x617;
assign c8330 =  x258 &  x398 &  x454 &  x482 &  x566 &  x594 & ~x71 & ~x731;
assign c8332 =  x592 &  x734;
assign c8334 =  x380 &  x408 &  x436 & ~x7 & ~x24 & ~x56 & ~x96 & ~x110 & ~x133 & ~x169 & ~x216 & ~x222 & ~x271 & ~x327 & ~x337 & ~x360 & ~x388 & ~x578;
assign c8336 =  x402 &  x597 & ~x259 & ~x365 & ~x443 & ~x684;
assign c8338 =  x404 &  x653 & ~x63 & ~x205 & ~x287;
assign c8340 =  x620 & ~x1 & ~x59 & ~x89 & ~x162 & ~x163 & ~x239 & ~x252 & ~x365 & ~x445 & ~x492 & ~x764;
assign c8342 =  x520 &  x545 &  x710;
assign c8344 =  x433 &  x682;
assign c8346 =  x434 &  x626 & ~x111 & ~x142 & ~x172 & ~x287 & ~x344 & ~x371 & ~x426 & ~x679 & ~x691 & ~x707;
assign c8348 =  x407 &  x435 &  x463 & ~x52 & ~x271 & ~x327 & ~x355 & ~x684;
assign c8350 =  x425 & ~x14 & ~x113 & ~x223 & ~x253 & ~x376 & ~x377 & ~x406 & ~x417 & ~x418 & ~x623 & ~x693 & ~x757 & ~x772;
assign c8352 =  x436 &  x492 & ~x41 & ~x178 & ~x220 & ~x273 & ~x319;
assign c8354 =  x588 & ~x391;
assign c8356 =  x16 &  x404 & ~x111 & ~x453;
assign c8358 =  x508 &  x509 &  x677;
assign c8360 =  x747 & ~x443 & ~x661;
assign c8362 =  x505 & ~x618;
assign c8364 =  x183 &  x407 &  x432 &  x460 & ~x398;
assign c8366 =  x15 &  x377 &  x488 & ~x455;
assign c8368 =  x594 & ~x21 & ~x23 & ~x55 & ~x117 & ~x136 & ~x173 & ~x310 & ~x312 & ~x335 & ~x367 & ~x436 & ~x492 & ~x577 & ~x599 & ~x615 & ~x775;
assign c8370 =  x426 &  x565 &  x593 &  x678 & ~x653;
assign c8372 =  x481 &  x509 & ~x15 & ~x79 & ~x99 & ~x225 & ~x404 & ~x413 & ~x433 & ~x625;
assign c8374 =  x451 & ~x80 & ~x101 & ~x252 & ~x303 & ~x376 & ~x405 & ~x513 & ~x779;
assign c8376 =  x463 &  x544 &  x746 & ~x425 & ~x582 & ~x606 & ~x640;
assign c8378 =  x566 &  x590;
assign c8380 =  x737 &  x747;
assign c8382 =  x746 & ~x275 & ~x384 & ~x413 & ~x415 & ~x470 & ~x498 & ~x527 & ~x657 & ~x659 & ~x661 & ~x664;
assign c8384 = ~x3 & ~x33 & ~x112 & ~x144 & ~x167 & ~x240 & ~x288 & ~x337 & ~x381 & ~x423 & ~x447 & ~x466 & ~x491 & ~x492 & ~x547 & ~x604 & ~x717 & ~x719;
assign c8386 = ~x18 & ~x29 & ~x30 & ~x54 & ~x57 & ~x59 & ~x105 & ~x193 & ~x223 & ~x247 & ~x275 & ~x281 & ~x301 & ~x309 & ~x358 & ~x360 & ~x387 & ~x418 & ~x435 & ~x444 & ~x447 & ~x491 & ~x546 & ~x558 & ~x697 & ~x698 & ~x707 & ~x729 & ~x730 & ~x738 & ~x741 & ~x759 & ~x769 & ~x777;
assign c8388 =  x459 &  x681 & ~x91 & ~x427 & ~x483 & ~x509;
assign c8390 =  x402 &  x458 &  x597 & ~x21 & ~x252 & ~x314;
assign c8392 =  x151 &  x402 &  x430 & ~x27 & ~x30 & ~x55 & ~x56 & ~x57 & ~x58 & ~x60 & ~x91 & ~x116 & ~x120 & ~x138 & ~x143 & ~x145 & ~x170 & ~x227 & ~x285 & ~x307 & ~x308 & ~x311 & ~x313 & ~x341 & ~x363 & ~x396 & ~x756;
assign c8394 =  x425 &  x505 & ~x303 & ~x445;
assign c8396 =  x15 &  x405 & ~x32 & ~x52 & ~x55 & ~x106 & ~x115 & ~x144 & ~x223 & ~x276 & ~x305 & ~x341 & ~x362 & ~x369 & ~x370 & ~x388 & ~x400 & ~x451 & ~x536;
assign c8398 =  x407 &  x488 &  x716 & ~x328;
assign c8400 =  x487 &  x737;
assign c8402 =  x739 &  x744 & ~x582 & ~x684;
assign c8404 =  x401 &  x652 & ~x27 & ~x197 & ~x363 & ~x369 & ~x420 & ~x450 & ~x546;
assign c8406 =  x315 &  x343 &  x371 &  x399 &  x455 &  x483 &  x511 &  x539 &  x567 &  x623 & ~x54 & ~x62 & ~x85 & ~x110 & ~x310 & ~x335 & ~x363 & ~x390;
assign c8408 = ~x3 & ~x21 & ~x109 & ~x259 & ~x369 & ~x492 & ~x518 & ~x545 & ~x546 & ~x572 & ~x733 & ~x746 & ~x747 & ~x780;
assign c8410 =  x372 &  x428 &  x652 & ~x518 & ~x544 & ~x572;
assign c8412 =  x406 &  x433 & ~x92 & ~x188 & ~x204 & ~x259 & ~x299 & ~x394 & ~x398 & ~x444 & ~x454 & ~x637;
assign c8414 =  x708 & ~x23 & ~x311 & ~x369 & ~x492 & ~x519 & ~x630;
assign c8416 =  x735 & ~x108 & ~x190 & ~x508 & ~x684;
assign c8418 =  x701;
assign c8420 =  x743 &  x768 & ~x526 & ~x633 & ~x684 & ~x688;
assign c8422 =  x295 &  x462 &  x488 &  x716 & ~x137 & ~x276 & ~x312 & ~x370 & ~x451;
assign c8424 =  x341 &  x508 & ~x43 & ~x75 & ~x101 & ~x404 & ~x702;
assign c8426 =  x664 & ~x59 & ~x117 & ~x222 & ~x283 & ~x386 & ~x472 & ~x475 & ~x548 & ~x587 & ~x605 & ~x628 & ~x758;
assign c8428 =  x213 &  x242 &  x270 &  x297 &  x353 & ~x282 & ~x575;
assign c8430 =  x540 & ~x3 & ~x22 & ~x60 & ~x79 & ~x119 & ~x147 & ~x169 & ~x280 & ~x369 & ~x396 & ~x465 & ~x491 & ~x519 & ~x546 & ~x733 & ~x773 & ~x774;
assign c8432 =  x767 & ~x259 & ~x329 & ~x684 & ~x687;
assign c8434 =  x719 &  x736 & ~x217 & ~x498;
assign c8436 =  x266 &  x350 &  x378 &  x406 &  x434 &  x461 & ~x109 & ~x170 & ~x259 & ~x311 & ~x440 & ~x451 & ~x732 & ~x736;
assign c8438 =  x376 & ~x156 & ~x205 & ~x225 & ~x255 & ~x258 & ~x449;
assign c8440 =  x433 & ~x1 & ~x41 & ~x289;
assign c8442 =  x321 &  x653 & ~x173 & ~x202 & ~x478;
assign c8444 =  x482 &  x618 &  x622 & ~x283;
assign c8446 =  x492 &  x747 & ~x142;
assign c8448 =  x379 &  x407 &  x463 &  x491 & ~x125 & ~x578;
assign c8450 = ~x274 & ~x329 & ~x405;
assign c8452 =  x508 &  x509 &  x535 &  x536 &  x590 & ~x417;
assign c8454 =  x491 &  x744 & ~x343 & ~x429 & ~x440 & ~x578 & ~x607;
assign c8456 =  x407 &  x461 & ~x75 & ~x90 & ~x109 & ~x161 & ~x200 & ~x214 & ~x247 & ~x283 & ~x328 & ~x369 & ~x389 & ~x442 & ~x498 & ~x619 & ~x779;
assign c8458 =  x706 & ~x1 & ~x109 & ~x135 & ~x195 & ~x326 & ~x760;
assign c8460 =  x491 &  x544 &  x743 & ~x219 & ~x396 & ~x523 & ~x526 & ~x551 & ~x582;
assign c8462 =  x491 &  x710 &  x745;
assign c8464 =  x539 &  x735 & ~x507 & ~x628;
assign c8466 =  x428 &  x456 &  x735;
assign c8468 = ~x6 & ~x50 & ~x58 & ~x60 & ~x77 & ~x107 & ~x110 & ~x112 & ~x115 & ~x135 & ~x140 & ~x199 & ~x218 & ~x219 & ~x231 & ~x248 & ~x314 & ~x340 & ~x446 & ~x449 & ~x465 & ~x473 & ~x474 & ~x491 & ~x520 & ~x546 & ~x739 & ~x745;
assign c8470 =  x457 &  x607 & ~x115 & ~x533;
assign c8472 =  x396 &  x477 & ~x387 & ~x401 & ~x430;
assign c8474 =  x735 & ~x87;
assign c8476 =  x347 &  x403 &  x624 & ~x63 & ~x88 & ~x253 & ~x370 & ~x425;
assign c8478 = ~x60 & ~x79 & ~x88 & ~x99 & ~x144 & ~x145 & ~x156 & ~x194 & ~x202 & ~x224 & ~x297 & ~x339 & ~x369 & ~x391 & ~x436 & ~x548 & ~x549 & ~x576 & ~x578 & ~x606 & ~x728;
assign c8480 =  x351 &  x407 & ~x111 & ~x114 & ~x158 & ~x169 & ~x215 & ~x242 & ~x271 & ~x279 & ~x302 & ~x328 & ~x330 & ~x332 & ~x684;
assign c8482 =  x509 &  x537 & ~x14 & ~x44 & ~x52 & ~x310 & ~x332 & ~x337 & ~x362 & ~x488 & ~x498 & ~x544 & ~x570 & ~x571 & ~x600 & ~x730 & ~x775;
assign c8484 =  x397 & ~x1 & ~x28 & ~x54 & ~x61 & ~x74 & ~x75 & ~x137 & ~x273 & ~x364 & ~x743 & ~x775;
assign c8486 = ~x33 & ~x36 & ~x37 & ~x57 & ~x67 & ~x75 & ~x142 & ~x144 & ~x151 & ~x299 & ~x309 & ~x327 & ~x334 & ~x400 & ~x411 & ~x420 & ~x472 & ~x617 & ~x618 & ~x684 & ~x696 & ~x769;
assign c8488 =  x398 &  x538 &  x563 &  x594;
assign c8490 =  x617 &  x678 & ~x450;
assign c8492 =  x320 &  x663 & ~x498 & ~x573;
assign c8494 =  x718 &  x719 & ~x222 & ~x244 & ~x498 & ~x600 & ~x657;
assign c8496 =  x425 &  x506 & ~x334 & ~x404 & ~x430 & ~x518;
assign c8498 =  x433 & ~x121 & ~x136 & ~x159 & ~x192 & ~x205 & ~x287 & ~x288 & ~x318 & ~x369 & ~x371 & ~x400 & ~x401;
assign c81 =  x388 & ~x645 & ~x650;
assign c83 =  x388;
assign c85 =  x496 &  x579;
assign c87 = ~x106 & ~x209 & ~x221 & ~x369 & ~x394 & ~x422 & ~x547 & ~x619 & ~x628 & ~x761 & ~x777;
assign c89 =  x174 &  x595;
assign c811 =  x550 &  x578 & ~x511 & ~x537;
assign c813 =  x259 &  x514 & ~x208 & ~x209;
assign c815 = ~x95 & ~x444 & ~x482 & ~x510 & ~x511 & ~x514 & ~x537 & ~x562 & ~x567 & ~x569 & ~x594 & ~x624 & ~x639 & ~x664 & ~x665 & ~x754;
assign c817 =  x138;
assign c819 =  x684 & ~x143 & ~x160 & ~x452 & ~x480 & ~x554 & ~x610 & ~x635 & ~x637 & ~x664 & ~x678 & ~x689;
assign c821 =  x686 &  x713 & ~x122;
assign c823 =  x603 &  x659 & ~x567;
assign c825 =  x446;
assign c827 =  x345 & ~x240 & ~x568 & ~x582 & ~x733 & ~x759 & ~x779;
assign c829 =  x40 &  x97 &  x627 &  x655;
assign c831 =  x48;
assign c833 =  x417;
assign c835 =  x554 &  x582 &  x610 & ~x208;
assign c837 =  x69 &  x627 &  x683 & ~x527 & ~x591 & ~x637;
assign c839 =  x628 & ~x194 & ~x555;
assign c841 =  x96 & ~x164 & ~x171 & ~x197 & ~x240 & ~x312 & ~x501 & ~x527 & ~x536 & ~x587 & ~x593 & ~x610 & ~x635 & ~x637 & ~x649 & ~x665 & ~x677 & ~x723 & ~x761;
assign c843 =  x173 & ~x209;
assign c845 = ~x131 & ~x253 & ~x280 & ~x511 & ~x536 & ~x566 & ~x567 & ~x572 & ~x582 & ~x595 & ~x619 & ~x648 & ~x669 & ~x760 & ~x771;
assign c847 = ~x30 & ~x167 & ~x179 & ~x194 & ~x208 & ~x209 & ~x236 & ~x237 & ~x238 & ~x239 & ~x281 & ~x619 & ~x646 & ~x694 & ~x727 & ~x775;
assign c849 = ~x139 & ~x213 & ~x267 & ~x302 & ~x308 & ~x567 & ~x593 & ~x616 & ~x621 & ~x635 & ~x642 & ~x673 & ~x704 & ~x732 & ~x759 & ~x760 & ~x761;
assign c851 =  x356 &  x382 & ~x133 & ~x694;
assign c853 =  x467 & ~x16 & ~x139 & ~x161 & ~x502 & ~x592 & ~x720;
assign c855 = ~x88 & ~x145 & ~x173 & ~x226 & ~x356 & ~x476 & ~x511 & ~x541 & ~x567 & ~x581 & ~x585 & ~x591 & ~x592 & ~x593 & ~x610 & ~x620 & ~x717 & ~x774;
assign c857 =  x69 &  x467 & ~x694;
assign c859 = ~x265 & ~x266 & ~x267 & ~x294 & ~x296 & ~x449 & ~x555 & ~x727 & ~x752;
assign c861 =  x68 &  x97 & ~x679 & ~x720;
assign c863 =  x388 & ~x293;
assign c865 =  x314 &  x542;
assign c867 = ~x12 & ~x95 & ~x112 & ~x142 & ~x382 & ~x409 & ~x539 & ~x555 & ~x567 & ~x576 & ~x622 & ~x623 & ~x650 & ~x654 & ~x677 & ~x709 & ~x720;
assign c869 =  x571 &  x656;
assign c871 =  x356 &  x357 & ~x132 & ~x694;
assign c873 =  x334;
assign c875 = ~x510 & ~x592 & ~x598 & ~x619 & ~x621 & ~x641 & ~x678 & ~x741 & ~x760;
assign c877 =  x284 & ~x153;
assign c879 = ~x111 & ~x430 & ~x481 & ~x512 & ~x525 & ~x562 & ~x589 & ~x594 & ~x613 & ~x650 & ~x664 & ~x672 & ~x678 & ~x697;
assign c881 =  x521 &  x578 & ~x19 & ~x163 & ~x591 & ~x673;
assign c883 =  x70 &  x265 & ~x74 & ~x161 & ~x387 & ~x415 & ~x505 & ~x536 & ~x641 & ~x663;
assign c885 =  x494 &  x551 & ~x28 & ~x429 & ~x452 & ~x503;
assign c887 =  x627 &  x685 &  x713;
assign c889 =  x326 &  x357;
assign c891 =  x580 & ~x138 & ~x197 & ~x227 & ~x388 & ~x444 & ~x472 & ~x556 & ~x612 & ~x617 & ~x629 & ~x646 & ~x729;
assign c893 =  x154 &  x155 &  x181 &  x292 & ~x143 & ~x269 & ~x423 & ~x532;
assign c895 = ~x168 & ~x238 & ~x266 & ~x267 & ~x269 & ~x296 & ~x540 & ~x567 & ~x595 & ~x614;
assign c897 =  x107 & ~x246;
assign c899 =  x175 &  x204 & ~x373 & ~x474 & ~x619;
assign c8101 =  x199;
assign c8103 =  x604 & ~x591;
assign c8105 =  x388;
assign c8107 =  x382 & ~x0 & ~x102 & ~x130 & ~x172 & ~x188 & ~x452 & ~x532 & ~x583 & ~x585 & ~x611 & ~x621 & ~x660 & ~x673 & ~x694;
assign c8109 = ~x65 & ~x95 & ~x151 & ~x209 & ~x210 & ~x236 & ~x238 & ~x264 & ~x265 & ~x266 & ~x466 & ~x644 & ~x669 & ~x728;
assign c8111 =  x333;
assign c8113 =  x759;
assign c8115 =  x522 &  x551 & ~x242 & ~x446 & ~x481;
assign c8117 = ~x24 & ~x33 & ~x59 & ~x106 & ~x139 & ~x208 & ~x209 & ~x235 & ~x236 & ~x251 & ~x254 & ~x256 & ~x306 & ~x307 & ~x373 & ~x393 & ~x417 & ~x421 & ~x475 & ~x476 & ~x505 & ~x506 & ~x533 & ~x534 & ~x561 & ~x591 & ~x620 & ~x669 & ~x674 & ~x723;
assign c8119 =  x385 &  x386 & ~x84 & ~x302 & ~x761;
assign c8121 =  x446;
assign c8123 =  x467 &  x493 &  x495;
assign c8125 =  x288 & ~x175 & ~x620 & ~x650 & ~x676;
assign c8127 =  x362;
assign c8129 =  x341 &  x541 & ~x372;
assign c8131 =  x137;
assign c8133 =  x209 &  x571 &  x627 & ~x575;
assign c8135 =  x89 &  x300;
assign c8137 =  x386 & ~x133;
assign c8139 =  x98 & ~x593 & ~x595 & ~x597;
assign c8141 =  x205 &  x629;
assign c8143 =  x204 & ~x98 & ~x100 & ~x166 & ~x591 & ~x645;
assign c8145 =  x302 &  x389;
assign c8147 = ~x16 & ~x32 & ~x113 & ~x223 & ~x307 & ~x470 & ~x486 & ~x551 & ~x555 & ~x607 & ~x622 & ~x650 & ~x663 & ~x677 & ~x719 & ~x754 & ~x774;
assign c8149 =  x173 & ~x236;
assign c8151 =  x362;
assign c8153 =  x386 & ~x59 & ~x78;
assign c8155 =  x190 & ~x52 & ~x152 & ~x281 & ~x386 & ~x448 & ~x616 & ~x644;
assign c8157 =  x388;
assign c8159 =  x518 &  x630 & ~x567;
assign c8161 =  x334 &  x335;
assign c8163 =  x118;
assign c8165 = ~x0 & ~x194 & ~x384 & ~x439 & ~x480 & ~x499 & ~x511 & ~x542 & ~x591 & ~x592 & ~x623 & ~x624 & ~x665 & ~x666 & ~x740 & ~x770;
assign c8167 =  x232 & ~x8 & ~x75 & ~x111 & ~x132 & ~x364 & ~x495 & ~x631;
assign c8169 =  x226;
assign c8171 =  x106 &  x285;
assign c8173 =  x386 &  x415 & ~x193 & ~x219;
assign c8175 =  x412 & ~x242 & ~x666;
assign c8177 =  x118 &  x119 & ~x154;
assign c8179 =  x326 &  x604;
assign c8181 =  x267 &  x602 &  x630 & ~x466 & ~x606 & ~x607 & ~x619 & ~x641;
assign c8183 =  x391;
assign c8185 =  x683 &  x711 & ~x105 & ~x160 & ~x621 & ~x637 & ~x678 & ~x704;
assign c8187 =  x523 & ~x287 & ~x454 & ~x616;
assign c8189 =  x148 &  x177 & ~x238 & ~x266;
assign c8191 =  x109;
assign c8193 =  x202 &  x231 & ~x70 & ~x501 & ~x589;
assign c8195 =  x77;
assign c8197 =  x237 &  x264 &  x265 &  x686;
assign c8199 =  x237 &  x599 &  x714;
assign c8201 = ~x17 & ~x60 & ~x167 & ~x173 & ~x251 & ~x513 & ~x567 & ~x595 & ~x596 & ~x616 & ~x623 & ~x645 & ~x646 & ~x677 & ~x678 & ~x699 & ~x739 & ~x740 & ~x747 & ~x760;
assign c8203 =  x178 &  x180 &  x181 & ~x261;
assign c8205 = ~x5 & ~x21 & ~x30 & ~x51 & ~x62 & ~x86 & ~x88 & ~x110 & ~x138 & ~x199 & ~x201 & ~x229 & ~x230 & ~x314 & ~x331 & ~x341 & ~x385 & ~x411 & ~x438 & ~x441 & ~x442 & ~x444 & ~x455 & ~x458 & ~x485 & ~x507 & ~x530 & ~x562 & ~x563 & ~x567 & ~x585 & ~x593 & ~x613 & ~x620 & ~x621 & ~x622 & ~x647 & ~x649 & ~x651 & ~x665 & ~x666 & ~x670 & ~x677 & ~x678 & ~x679 & ~x745 & ~x753 & ~x779;
assign c8207 =  x499 &  x527 &  x555 & ~x277 & ~x697;
assign c8209 =  x658 &  x686 & ~x579 & ~x620 & ~x622;
assign c8211 =  x437 &  x438 & ~x18 & ~x54 & ~x133 & ~x242 & ~x338 & ~x392 & ~x420 & ~x423 & ~x449 & ~x534 & ~x563 & ~x648;
assign c8213 =  x522 & ~x223 & ~x456 & ~x502 & ~x563 & ~x602 & ~x621;
assign c8215 =  x97 &  x98 &  x126 & ~x179 & ~x645;
assign c8217 =  x355 &  x356 & ~x27 & ~x81 & ~x111 & ~x112 & ~x197 & ~x250 & ~x337 & ~x665 & ~x693 & ~x694 & ~x695 & ~x730;
assign c8219 =  x172 & ~x236;
assign c8221 =  x89;
assign c8223 = ~x0 & ~x18 & ~x58 & ~x64 & ~x108 & ~x139 & ~x140 & ~x156 & ~x218 & ~x300 & ~x328 & ~x426 & ~x460 & ~x499 & ~x555 & ~x585 & ~x591 & ~x593 & ~x614 & ~x620 & ~x644 & ~x647 & ~x666 & ~x755 & ~x757;
assign c8225 =  x136;
assign c8227 =  x657 &  x686 &  x714 & ~x662;
assign c8229 =  x395 &  x640;
assign c8231 =  x192;
assign c8233 =  x144;
assign c8235 = ~x57 & ~x93 & ~x102 & ~x254 & ~x366 & ~x367 & ~x413 & ~x554 & ~x567 & ~x594 & ~x596 & ~x597 & ~x600 & ~x621 & ~x678 & ~x703 & ~x706;
assign c8237 =  x120 &  x121 &  x150 & ~x726;
assign c8239 =  x523 & ~x721;
assign c8241 =  x498 &  x553 & ~x82 & ~x532 & ~x560 & ~x617;
assign c8243 =  x576 &  x605;
assign c8245 =  x124 &  x125 &  x771 & ~x650 & ~x663;
assign c8247 = ~x81 & ~x269 & ~x293 & ~x555 & ~x583 & ~x595 & ~x620 & ~x621 & ~x642 & ~x644 & ~x780;
assign c8249 =  x551 & ~x242 & ~x563 & ~x591 & ~x776;
assign c8251 =  x317 &  x600 &  x627 & ~x617;
assign c8253 =  x305;
assign c8255 =  x71 &  x601 &  x629 &  x657 & ~x333;
assign c8257 =  x346 & ~x94 & ~x179 & ~x541 & ~x595;
assign c8259 = ~x52 & ~x74 & ~x93 & ~x171 & ~x230 & ~x285 & ~x340 & ~x366 & ~x451 & ~x494 & ~x550 & ~x552 & ~x554 & ~x566 & ~x568 & ~x598 & ~x625 & ~x642 & ~x645 & ~x650 & ~x701 & ~x709;
assign c8261 =  x288 & ~x154 & ~x210 & ~x266 & ~x267 & ~x634;
assign c8263 = ~x146 & ~x225 & ~x233 & ~x251 & ~x442 & ~x449 & ~x479 & ~x507 & ~x512 & ~x513 & ~x537 & ~x567 & ~x617 & ~x641 & ~x648 & ~x649 & ~x666 & ~x678 & ~x700 & ~x706;
assign c8265 =  x86;
assign c8267 =  x116 & ~x179 & ~x659;
assign c8269 =  x79;
assign c8271 =  x360 & ~x191;
assign c8273 =  x272 & ~x83 & ~x104 & ~x363 & ~x383 & ~x477;
assign c8275 =  x117 & ~x266;
assign c8277 =  x602 &  x686;
assign c8279 =  x216;
assign c8281 =  x389;
assign c8283 = ~x4 & ~x5 & ~x134 & ~x157 & ~x163 & ~x238 & ~x266 & ~x267 & ~x269 & ~x526 & ~x554 & ~x609 & ~x643 & ~x644 & ~x648 & ~x728 & ~x753 & ~x765;
assign c8285 = ~x3 & ~x8 & ~x50 & ~x54 & ~x63 & ~x89 & ~x110 & ~x117 & ~x160 & ~x193 & ~x277 & ~x278 & ~x315 & ~x342 & ~x442 & ~x480 & ~x484 & ~x499 & ~x507 & ~x530 & ~x534 & ~x555 & ~x563 & ~x591 & ~x598 & ~x618 & ~x620 & ~x622 & ~x640 & ~x648 & ~x650 & ~x663 & ~x691 & ~x703 & ~x706 & ~x747 & ~x752;
assign c8287 =  x123 &  x124 &  x125 & ~x187 & ~x365 & ~x554 & ~x616 & ~x620 & ~x621 & ~x622 & ~x703;
assign c8289 =  x123 &  x125 & ~x620 & ~x621 & ~x649;
assign c8291 =  x634 & ~x513 & ~x588 & ~x591;
assign c8293 =  x97 &  x99 &  x126 & ~x179;
assign c8295 =  x418;
assign c8297 = ~x4 & ~x23 & ~x170 & ~x210 & ~x277 & ~x281 & ~x480 & ~x498 & ~x504 & ~x526 & ~x529 & ~x562 & ~x565 & ~x593 & ~x603 & ~x610 & ~x621 & ~x635 & ~x666 & ~x671 & ~x734 & ~x759;
assign c8299 =  x181 &  x184 & ~x1 & ~x27 & ~x616 & ~x653 & ~x768;
assign c8301 =  x603 & ~x538;
assign c8303 =  x149 &  x178 &  x179 & ~x164;
assign c8305 =  x603 &  x632;
assign c8307 =  x285;
assign c8309 =  x118 & ~x41 & ~x154;
assign c8311 =  x286 &  x610 & ~x589;
assign c8313 =  x496 &  x497 &  x525 &  x553 & ~x361 & ~x386;
assign c8315 =  x571 &  x634 & ~x616;
assign c8317 =  x199;
assign c8319 =  x175 &  x176 &  x205 & ~x70;
assign c8321 =  x331 &  x389;
assign c8323 =  x133 &  x173;
assign c8325 =  x98 &  x100 &  x126 & ~x255 & ~x493 & ~x501 & ~x559 & ~x672 & ~x699;
assign c8327 =  x601 &  x629 & ~x1 & ~x3 & ~x56 & ~x80 & ~x83 & ~x107 & ~x108 & ~x109 & ~x169 & ~x219 & ~x308 & ~x364 & ~x418 & ~x504 & ~x526 & ~x550 & ~x551 & ~x553 & ~x555 & ~x562 & ~x639 & ~x642 & ~x643 & ~x753 & ~x757 & ~x780 & ~x782;
assign c8329 =  x683 &  x771 & ~x241 & ~x650;
assign c8331 =  x300 & ~x440 & ~x504 & ~x724;
assign c8333 =  x146 & ~x761;
assign c8335 =  x580 &  x608 & ~x0 & ~x94 & ~x474 & ~x484;
assign c8337 = ~x0 & ~x39 & ~x479 & ~x503 & ~x507 & ~x567 & ~x568 & ~x593 & ~x594 & ~x595 & ~x598 & ~x622 & ~x648 & ~x650 & ~x678;
assign c8339 = ~x24 & ~x32 & ~x83 & ~x115 & ~x172 & ~x225 & ~x282 & ~x309 & ~x415 & ~x440 & ~x465 & ~x469 & ~x471 & ~x482 & ~x496 & ~x497 & ~x511 & ~x566 & ~x595 & ~x621 & ~x644 & ~x650 & ~x678 & ~x682 & ~x692 & ~x721 & ~x734 & ~x759;
assign c8341 = ~x38 & ~x95 & ~x181 & ~x208 & ~x236 & ~x237 & ~x238 & ~x264 & ~x293 & ~x540 & ~x574;
assign c8343 =  x178 &  x603;
assign c8345 =  x181 &  x627 &  x655 &  x715;
assign c8347 =  x69 &  x683 &  x712 & ~x640 & ~x663;
assign c8349 =  x332 & ~x555;
assign c8351 =  x514 &  x541 &  x595 & ~x683;
assign c8353 =  x311 &  x339;
assign c8355 =  x95 &  x96 & ~x242 & ~x594 & ~x648 & ~x733;
assign c8357 =  x410 &  x412 & ~x291;
assign c8359 =  x498 & ~x58 & ~x227 & ~x449 & ~x533 & ~x562 & ~x616 & ~x700 & ~x729;
assign c8361 =  x468 &  x577;
assign c8363 =  x333 &  x418;
assign c8365 =  x260 & ~x181 & ~x209 & ~x210 & ~x213 & ~x620 & ~x641;
assign c8367 =  x121 &  x124;
assign c8369 =  x579 & ~x29 & ~x58 & ~x304 & ~x424 & ~x427 & ~x429 & ~x451 & ~x479 & ~x507 & ~x561 & ~x562 & ~x676;
assign c8371 =  x265 &  x429 & ~x493 & ~x680;
assign c8373 =  x498 & ~x27 & ~x113 & ~x131 & ~x196 & ~x272 & ~x505 & ~x616 & ~x618 & ~x670 & ~x728;
assign c8375 =  x204 &  x205 &  x206;
assign c8377 =  x389 & ~x678;
assign c8379 =  x237 &  x715;
assign c8381 =  x203 & ~x8 & ~x111 & ~x227 & ~x254 & ~x336 & ~x391 & ~x400 & ~x505 & ~x530 & ~x590 & ~x641 & ~x642 & ~x646;
assign c8383 =  x125 & ~x18 & ~x204 & ~x595 & ~x650 & ~x768;
assign c8385 =  x390 &  x391;
assign c8387 =  x146 &  x176 & ~x762;
assign c8389 = ~x39 & ~x205 & ~x208 & ~x236 & ~x238 & ~x291 & ~x365 & ~x620 & ~x674;
assign c8391 =  x389 &  x446;
assign c8393 =  x73 &  x101 & ~x10 & ~x280 & ~x336 & ~x615 & ~x653 & ~x700 & ~x740 & ~x764 & ~x768;
assign c8395 = ~x95 & ~x236 & ~x237 & ~x465 & ~x526 & ~x677 & ~x697 & ~x722;
assign c8397 =  x204 &  x206 & ~x168 & ~x696;
assign c8399 =  x602 &  x658;
assign c8401 =  x97 &  x627 &  x684 &  x713;
assign c8403 =  x334;
assign c8405 =  x551 & ~x227 & ~x359 & ~x387 & ~x448 & ~x455 & ~x531 & ~x590 & ~x616 & ~x749;
assign c8407 =  x383 & ~x209 & ~x621;
assign c8409 =  x41 & ~x49 & ~x283 & ~x433 & ~x535 & ~x621 & ~x637 & ~x723 & ~x736;
assign c8411 =  x170;
assign c8413 =  x233 &  x628;
assign c8415 =  x656 &  x684 &  x713 & ~x665;
assign c8417 =  x219 & ~x96 & ~x387;
assign c8419 =  x603 &  x632 & ~x511;
assign c8421 =  x424;
assign c8423 =  x384 & ~x208 & ~x217 & ~x685 & ~x748;
assign c8425 =  x657 &  x684 & ~x608 & ~x616 & ~x665;
assign c8427 =  x264 & ~x160 & ~x173 & ~x358 & ~x420 & ~x470 & ~x509 & ~x554 & ~x568 & ~x589 & ~x592 & ~x594 & ~x595 & ~x652 & ~x678 & ~x721 & ~x764;
assign c8429 =  x474;
assign c8431 =  x122 &  x124 &  x125 & ~x649;
assign c8433 =  x166;
assign c8435 = ~x10 & ~x118 & ~x267 & ~x269 & ~x555 & ~x563 & ~x591 & ~x620 & ~x678 & ~x700;
assign c8437 =  x528 &  x584;
assign c8439 = ~x45 & ~x46 & ~x80 & ~x85 & ~x105 & ~x147 & ~x161 & ~x203 & ~x217 & ~x220 & ~x247 & ~x279 & ~x302 & ~x314 & ~x330 & ~x368 & ~x413 & ~x454 & ~x481 & ~x502 & ~x534 & ~x535 & ~x539 & ~x540 & ~x593 & ~x594 & ~x595 & ~x596 & ~x611 & ~x613 & ~x616 & ~x618 & ~x620 & ~x621 & ~x643 & ~x645 & ~x648 & ~x650 & ~x679 & ~x726 & ~x734 & ~x737 & ~x780;
assign c8441 =  x285 &  x582 &  x611;
assign c8443 =  x182 &  x210 &  x265 & ~x77 & ~x344 & ~x351 & ~x474 & ~x709;
assign c8445 =  x274 & ~x555;
assign c8447 =  x205 &  x206 &  x207 & ~x534 & ~x619;
assign c8449 = ~x51 & ~x91 & ~x109 & ~x306 & ~x454 & ~x508 & ~x511 & ~x542 & ~x543 & ~x544 & ~x555 & ~x562 & ~x568 & ~x594 & ~x595 & ~x596 & ~x620 & ~x622 & ~x668;
assign c8451 =  x554 &  x610 & ~x645 & ~x670;
assign c8453 =  x601 &  x629 & ~x18 & ~x309 & ~x584 & ~x609 & ~x643 & ~x724 & ~x770;
assign c8455 =  x278;
assign c8457 =  x437 & ~x242 & ~x267 & ~x296;
assign c8459 =  x137;
assign c8461 =  x361 &  x446;
assign c8463 =  x203 & ~x138 & ~x390 & ~x455 & ~x501 & ~x507 & ~x562;
assign c8465 =  x494 &  x551 & ~x534 & ~x719;
assign c8467 =  x199 & ~x179;
assign c8469 =  x203 &  x541;
assign c8471 =  x331;
assign c8473 =  x172;
assign c8475 =  x547 &  x576 &  x633 & ~x452 & ~x503 & ~x508 & ~x558;
assign c8477 = ~x57 & ~x123 & ~x493 & ~x542 & ~x595 & ~x598 & ~x625 & ~x648 & ~x650 & ~x696 & ~x729;
assign c8479 =  x357 & ~x162;
assign c8481 =  x341 &  x638 & ~x616;
assign c8483 =  x334;
assign c8485 =  x159 &  x186 & ~x18 & ~x372 & ~x526;
assign c8487 =  x137;
assign c8489 =  x220;
assign c8491 =  x356 & ~x562 & ~x665;
assign c8493 =  x306;
assign c8495 =  x577 & ~x507 & ~x511 & ~x537 & ~x616 & ~x619;
assign c8497 =  x171;
assign c8499 =  x367 &  x648;
assign c90 =  x413 &  x737 & ~x268 & ~x580;
assign c92 =  x741 & ~x6 & ~x18 & ~x212 & ~x216 & ~x324;
assign c94 =  x59 & ~x585 & ~x611;
assign c96 =  x109 & ~x124 & ~x178;
assign c98 =  x685;
assign c910 =  x379 & ~x36 & ~x49 & ~x183 & ~x211 & ~x238 & ~x242 & ~x524 & ~x535 & ~x558 & ~x560 & ~x592 & ~x647 & ~x765 & ~x767 & ~x769 & ~x774 & ~x778;
assign c912 =  x413 & ~x0 & ~x15 & ~x21 & ~x160 & ~x218 & ~x241 & ~x246 & ~x252 & ~x274 & ~x279 & ~x296 & ~x324 & ~x325 & ~x503 & ~x580 & ~x611;
assign c914 =  x327 & ~x44 & ~x46 & ~x71 & ~x102 & ~x181 & ~x309 & ~x426 & ~x777;
assign c916 =  x438 &  x694;
assign c918 =  x485 &  x568 &  x650 & ~x612;
assign c920 = ~x9 & ~x150 & ~x186 & ~x205 & ~x210 & ~x238 & ~x400 & ~x550 & ~x610 & ~x646;
assign c922 =  x118 &  x405 & ~x47 & ~x68 & ~x69 & ~x125 & ~x311 & ~x336 & ~x420 & ~x534 & ~x674;
assign c924 = ~x213 & ~x298 & ~x342 & ~x402 & ~x421 & ~x511 & ~x551 & ~x625 & ~x650;
assign c926 =  x738 &  x739 &  x741 & ~x210 & ~x239 & ~x269 & ~x270 & ~x524 & ~x606 & ~x620 & ~x668;
assign c928 =  x170 & ~x80 & ~x617;
assign c930 =  x324 &  x351 &  x636;
assign c932 =  x572 &  x740 & ~x210 & ~x593;
assign c934 =  x459 & ~x17 & ~x40 & ~x181 & ~x212 & ~x237 & ~x453 & ~x471 & ~x475 & ~x478 & ~x527 & ~x532 & ~x593 & ~x697;
assign c936 =  x681 &  x685 &  x712 &  x715 & ~x501 & ~x553;
assign c938 =  x125 &  x546 &  x742 & ~x105 & ~x324 & ~x540;
assign c940 =  x294 &  x464 & ~x4 & ~x234 & ~x274 & ~x304 & ~x317 & ~x475 & ~x530 & ~x617 & ~x625 & ~x632 & ~x654 & ~x681;
assign c942 =  x746 &  x747 &  x748 & ~x584 & ~x636 & ~x646 & ~x651 & ~x677 & ~x735;
assign c944 =  x134 &  x238;
assign c946 =  x552 &  x723;
assign c948 =  x518 & ~x50 & ~x54 & ~x241 & ~x299 & ~x471 & ~x585 & ~x597;
assign c950 =  x109 &  x239 & ~x304 & ~x305;
assign c952 = ~x7 & ~x24 & ~x43 & ~x46 & ~x54 & ~x127 & ~x155 & ~x182 & ~x184 & ~x187 & ~x238 & ~x239 & ~x343 & ~x390 & ~x392 & ~x393 & ~x428 & ~x468 & ~x472 & ~x478 & ~x482 & ~x506 & ~x536 & ~x617 & ~x640 & ~x676 & ~x696 & ~x704 & ~x724 & ~x730 & ~x758 & ~x772 & ~x773 & ~x779;
assign c954 =  x212 &  x411 &  x525;
assign c956 =  x357 & ~x4 & ~x24 & ~x50 & ~x133 & ~x241 & ~x268 & ~x366 & ~x443 & ~x454 & ~x524 & ~x551 & ~x582 & ~x590;
assign c958 =  x242 &  x320 & ~x359 & ~x502 & ~x602 & ~x608 & ~x617;
assign c960 =  x438 &  x537 & ~x390 & ~x542 & ~x597 & ~x746;
assign c962 =  x268 &  x482 & ~x235 & ~x301;
assign c964 =  x324 & ~x59 & ~x101 & ~x387 & ~x418 & ~x585 & ~x687 & ~x713 & ~x715 & ~x740 & ~x763 & ~x767 & ~x772 & ~x773;
assign c966 = ~x56 & ~x131 & ~x155 & ~x186 & ~x262 & ~x347 & ~x374 & ~x402 & ~x528 & ~x652 & ~x674;
assign c968 =  x467 &  x553 &  x695;
assign c970 =  x441 &  x469 & ~x302 & ~x632;
assign c972 =  x301 &  x406 & ~x161 & ~x241 & ~x468;
assign c974 =  x441 &  x493 & ~x308 & ~x324;
assign c976 =  x429 &  x457 &  x539 & ~x35 & ~x279 & ~x477 & ~x617;
assign c978 =  x485 & ~x18 & ~x40 & ~x97 & ~x290 & ~x418 & ~x421 & ~x563 & ~x643 & ~x767;
assign c980 =  x434 &  x489 &  x517 & ~x33 & ~x128 & ~x263 & ~x478 & ~x618 & ~x737;
assign c982 =  x409 &  x495;
assign c984 = ~x52 & ~x73 & ~x76 & ~x131 & ~x132 & ~x213 & ~x218 & ~x239 & ~x244 & ~x343 & ~x402 & ~x449 & ~x456 & ~x483 & ~x564 & ~x585 & ~x594 & ~x640 & ~x676 & ~x708 & ~x724;
assign c986 =  x79 &  x704 & ~x178;
assign c988 =  x485 & ~x125 & ~x126 & ~x198 & ~x263 & ~x589 & ~x591 & ~x618 & ~x738;
assign c990 =  x605 &  x609 & ~x565;
assign c992 =  x295 &  x494 & ~x273 & ~x500 & ~x570 & ~x584 & ~x680 & ~x689 & ~x713;
assign c994 =  x711 &  x716 &  x744 &  x745 & ~x18 & ~x75 & ~x211 & ~x501 & ~x509 & ~x582 & ~x674;
assign c996 =  x300 &  x301 &  x354 &  x406 & ~x131 & ~x447;
assign c998 =  x525 &  x668;
assign c9100 =  x122 &  x517 & ~x187 & ~x605 & ~x763;
assign c9102 = ~x18 & ~x44 & ~x317 & ~x426 & ~x491 & ~x590;
assign c9104 =  x744 & ~x44 & ~x73 & ~x105 & ~x353 & ~x507 & ~x585 & ~x610 & ~x735 & ~x752;
assign c9106 = ~x7 & ~x37 & ~x129 & ~x187 & ~x235 & ~x362 & ~x400 & ~x444 & ~x589 & ~x669 & ~x684 & ~x713 & ~x740;
assign c9108 = ~x19 & ~x46 & ~x127 & ~x158 & ~x213 & ~x241 & ~x309 & ~x399 & ~x401 & ~x402 & ~x430 & ~x498 & ~x501 & ~x564 & ~x582 & ~x763;
assign c9110 =  x115 & ~x71 & ~x644;
assign c9112 =  x738 &  x741 & ~x46 & ~x297 & ~x551 & ~x577 & ~x661 & ~x676;
assign c9114 = ~x17 & ~x241 & ~x268 & ~x319 & ~x373 & ~x428 & ~x534 & ~x566 & ~x614 & ~x763;
assign c9116 =  x242 &  x584 & ~x694;
assign c9118 =  x329 &  x382 &  x407 & ~x17 & ~x18 & ~x136 & ~x160 & ~x240 & ~x337 & ~x444 & ~x510 & ~x581 & ~x592 & ~x676;
assign c9120 =  x207 &  x235 & ~x538 & ~x540 & ~x633;
assign c9122 =  x423 &  x673;
assign c9124 =  x730;
assign c9126 = ~x14 & ~x18 & ~x49 & ~x101 & ~x239 & ~x309 & ~x338 & ~x342 & ~x368 & ~x387 & ~x399 & ~x588 & ~x648 & ~x649 & ~x739 & ~x757;
assign c9128 =  x212 & ~x151;
assign c9130 =  x191 &  x350;
assign c9132 =  x709 &  x739 &  x740 & ~x72 & ~x268 & ~x522 & ~x605 & ~x614;
assign c9134 =  x431 & ~x152 & ~x359 & ~x390 & ~x411 & ~x465 & ~x535 & ~x545 & ~x585;
assign c9136 =  x496 &  x610 & ~x636;
assign c9138 =  x137 &  x646;
assign c9140 =  x413 & ~x305 & ~x376 & ~x581 & ~x752;
assign c9142 = ~x97 & ~x101 & ~x127 & ~x210 & ~x421 & ~x427 & ~x468 & ~x509 & ~x534 & ~x563 & ~x684;
assign c9144 =  x135 &  x268;
assign c9146 =  x731 & ~x290 & ~x607 & ~x693;
assign c9148 =  x546 &  x574 &  x744 & ~x81 & ~x134 & ~x163 & ~x214 & ~x215 & ~x593 & ~x609 & ~x610 & ~x649 & ~x650;
assign c9150 =  x118 & ~x17 & ~x74 & ~x99 & ~x103 & ~x104 & ~x254 & ~x282 & ~x307 & ~x338 & ~x363 & ~x442 & ~x530 & ~x534 & ~x555 & ~x585 & ~x587 & ~x672 & ~x753 & ~x765 & ~x767;
assign c9152 =  x125 &  x179 & ~x215 & ~x594 & ~x610;
assign c9154 =  x29;
assign c9156 =  x633 & ~x66 & ~x187 & ~x240;
assign c9158 =  x238 &  x324 & ~x361 & ~x364 & ~x393 & ~x501 & ~x585 & ~x613 & ~x671 & ~x689 & ~x713 & ~x745;
assign c9160 =  x206 &  x385 & ~x133 & ~x195 & ~x212 & ~x554 & ~x608 & ~x619;
assign c9162 =  x497 &  x611 & ~x625;
assign c9164 =  x519 &  x741 &  x772 & ~x238 & ~x566 & ~x650 & ~x735;
assign c9166 =  x441 &  x498 & ~x571;
assign c9168 =  x495 & ~x290 & ~x334 & ~x364 & ~x571 & ~x654 & ~x708 & ~x775;
assign c9170 =  x136 &  x239;
assign c9172 =  x484 & ~x23 & ~x235 & ~x276 & ~x388 & ~x643 & ~x689 & ~x773;
assign c9174 =  x88 & ~x11 & ~x68 & ~x367 & ~x582;
assign c9176 =  x711 &  x713 &  x716 & ~x16 & ~x49 & ~x212 & ~x550 & ~x553 & ~x639;
assign c9178 =  x494 & ~x417 & ~x560 & ~x654 & ~x743;
assign c9180 =  x206 &  x489 &  x517 & ~x132 & ~x456;
assign c9182 =  x386 &  x740 &  x744;
assign c9184 =  x494 &  x521 & ~x179 & ~x277 & ~x318 & ~x330 & ~x446 & ~x633 & ~x661 & ~x688;
assign c9186 = ~x83 & ~x183 & ~x235 & ~x289 & ~x318 & ~x425 & ~x526 & ~x536 & ~x720;
assign c9188 =  x410 & ~x335 & ~x365 & ~x447 & ~x458 & ~x558 & ~x569 & ~x597 & ~x605 & ~x651 & ~x782;
assign c9190 =  x267 &  x323 &  x538 & ~x391;
assign c9192 =  x403 & ~x14 & ~x55 & ~x125 & ~x126 & ~x180 & ~x212 & ~x371 & ~x411 & ~x412 & ~x438 & ~x449 & ~x464 & ~x492 & ~x528 & ~x556 & ~x611 & ~x648 & ~x760;
assign c9194 =  x239 & ~x168 & ~x234 & ~x235 & ~x577 & ~x597 & ~x605 & ~x614 & ~x632 & ~x633 & ~x653 & ~x654;
assign c9196 =  x712 &  x716 & ~x50 & ~x370 & ~x587 & ~x632 & ~x767;
assign c9198 = ~x17 & ~x18 & ~x49 & ~x55 & ~x70 & ~x128 & ~x130 & ~x490 & ~x491 & ~x495 & ~x498 & ~x509 & ~x524 & ~x532 & ~x554 & ~x602 & ~x644 & ~x752;
assign c9200 =  x115 & ~x134 & ~x605;
assign c9202 =  x739 &  x742 &  x744 & ~x163 & ~x251 & ~x551 & ~x553 & ~x606 & ~x609;
assign c9204 = ~x73 & ~x87 & ~x97 & ~x101 & ~x234 & ~x235 & ~x365 & ~x442 & ~x481 & ~x505 & ~x651 & ~x707 & ~x736 & ~x763;
assign c9206 =  x265 &  x565 & ~x578 & ~x597 & ~x626 & ~x710;
assign c9208 = ~x68 & ~x76 & ~x187 & ~x341 & ~x368 & ~x427 & ~x456 & ~x476 & ~x506 & ~x538 & ~x560 & ~x614 & ~x707 & ~x708 & ~x714;
assign c9210 = ~x14 & ~x101 & ~x112 & ~x130 & ~x131 & ~x133 & ~x186 & ~x210 & ~x212 & ~x238 & ~x283 & ~x400 & ~x427 & ~x453 & ~x469 & ~x527 & ~x590 & ~x647 & ~x706 & ~x761 & ~x781;
assign c9212 =  x268 & ~x124 & ~x281 & ~x290 & ~x331 & ~x361 & ~x387 & ~x615 & ~x683 & ~x690 & ~x713 & ~x745 & ~x763 & ~x775;
assign c9214 =  x739 &  x740 & ~x18 & ~x128 & ~x215 & ~x238 & ~x242 & ~x527 & ~x577 & ~x578 & ~x581 & ~x609 & ~x631 & ~x760;
assign c9216 =  x711 &  x739 &  x740 & ~x16 & ~x70 & ~x98 & ~x100 & ~x127 & ~x604 & ~x605;
assign c9218 =  x136 & ~x275;
assign c9220 =  x572 &  x710 & ~x238 & ~x578;
assign c9222 =  x715 & ~x130 & ~x238 & ~x240 & ~x256 & ~x425 & ~x448 & ~x456 & ~x757;
assign c9224 =  x211;
assign c9226 =  x610 & ~x663;
assign c9228 =  x709 &  x739 &  x742 & ~x607;
assign c9230 = ~x11 & ~x45 & ~x98 & ~x99 & ~x111 & ~x125 & ~x155 & ~x238 & ~x241 & ~x395 & ~x427 & ~x444 & ~x533 & ~x584 & ~x589 & ~x644 & ~x676;
assign c9232 =  x378 &  x484 & ~x152 & ~x329 & ~x359 & ~x590;
assign c9234 = ~x101 & ~x126 & ~x130 & ~x155 & ~x261 & ~x263 & ~x312 & ~x421 & ~x426 & ~x453 & ~x582;
assign c9236 =  x409 &  x564 & ~x416 & ~x596 & ~x604 & ~x660 & ~x707 & ~x721;
assign c9238 =  x567 &  x595 & ~x126 & ~x128 & ~x156 & ~x309 & ~x366 & ~x395 & ~x415 & ~x481 & ~x503 & ~x591;
assign c9240 =  x382 & ~x278 & ~x430 & ~x431 & ~x458 & ~x540 & ~x557 & ~x559 & ~x577 & ~x596 & ~x636;
assign c9242 =  x199 & ~x163 & ~x192 & ~x539;
assign c9244 =  x273 & ~x105 & ~x127 & ~x132 & ~x155 & ~x161 & ~x184 & ~x444 & ~x479 & ~x500 & ~x504 & ~x588 & ~x619 & ~x640 & ~x646 & ~x674 & ~x733;
assign c9246 =  x376 & ~x11 & ~x16 & ~x75 & ~x98 & ~x99 & ~x130 & ~x212 & ~x371 & ~x470 & ~x561 & ~x564 & ~x619 & ~x647 & ~x725;
assign c9248 =  x265 &  x565 & ~x560 & ~x575 & ~x585 & ~x596 & ~x609;
assign c9250 =  x496 &  x668;
assign c9252 = ~x82 & ~x210 & ~x239 & ~x401 & ~x456 & ~x564 & ~x584 & ~x604 & ~x605;
assign c9254 =  x545 & ~x238;
assign c9256 =  x459 & ~x54 & ~x163 & ~x186 & ~x208 & ~x414 & ~x453 & ~x616 & ~x773;
assign c9258 = ~x9 & ~x90 & ~x136 & ~x186 & ~x270 & ~x272 & ~x528 & ~x531 & ~x532 & ~x561 & ~x565 & ~x566 & ~x684 & ~x769;
assign c9260 =  x78 &  x239;
assign c9262 = ~x4 & ~x18 & ~x31 & ~x57 & ~x61 & ~x76 & ~x142 & ~x158 & ~x163 & ~x164 & ~x198 & ~x216 & ~x240 & ~x241 & ~x252 & ~x270 & ~x272 & ~x307 & ~x402 & ~x421 & ~x429 & ~x446 & ~x456 & ~x483 & ~x504 & ~x554 & ~x563 & ~x566 & ~x590 & ~x592 & ~x613 & ~x649 & ~x737 & ~x764;
assign c9264 =  x744 &  x745 & ~x46 & ~x160 & ~x240 & ~x373 & ~x400 & ~x429 & ~x510 & ~x582 & ~x666;
assign c9266 = ~x68 & ~x267 & ~x427 & ~x507 & ~x523 & ~x652 & ~x674 & ~x732 & ~x763;
assign c9268 =  x143 & ~x106 & ~x535 & ~x589 & ~x781;
assign c9270 =  x123 &  x150 & ~x155 & ~x290 & ~x477;
assign c9272 =  x409 &  x552 & ~x690;
assign c9274 =  x142 & ~x7 & ~x418;
assign c9276 =  x357 &  x410 & ~x213 & ~x267 & ~x511;
assign c9278 =  x459 &  x595 &  x623 & ~x18 & ~x111 & ~x308 & ~x614 & ~x640 & ~x696 & ~x756 & ~x763 & ~x764;
assign c9280 =  x330 &  x435 & ~x7 & ~x105 & ~x185 & ~x365 & ~x589;
assign c9282 = ~x38 & ~x155 & ~x212 & ~x267 & ~x400 & ~x644 & ~x647 & ~x772;
assign c9284 =  x739 &  x742 & ~x26 & ~x213 & ~x238 & ~x240 & ~x272 & ~x325 & ~x554 & ~x759;
assign c9286 =  x546 &  x741 &  x745 &  x747 & ~x610;
assign c9288 = ~x1 & ~x7 & ~x22 & ~x40 & ~x49 & ~x71 & ~x73 & ~x101 & ~x124 & ~x136 & ~x154 & ~x164 & ~x344 & ~x370 & ~x396 & ~x420 & ~x479 & ~x506 & ~x563 & ~x674 & ~x731;
assign c9290 =  x351 &  x494 & ~x362 & ~x390 & ~x448 & ~x474 & ~x633 & ~x682 & ~x713;
assign c9292 =  x81 & ~x221;
assign c9294 =  x519 & ~x16 & ~x131 & ~x166 & ~x212 & ~x297 & ~x458 & ~x483 & ~x538 & ~x554 & ~x558 & ~x563 & ~x566;
assign c9296 = ~x2 & ~x19 & ~x72 & ~x97 & ~x101 & ~x110 & ~x152 & ~x336 & ~x424 & ~x441 & ~x444 & ~x479 & ~x534 & ~x535 & ~x563 & ~x616 & ~x654 & ~x684 & ~x714 & ~x765 & ~x774;
assign c9298 =  x740 &  x744 & ~x44 & ~x109 & ~x160 & ~x189 & ~x448 & ~x449 & ~x510 & ~x530 & ~x589 & ~x605 & ~x612 & ~x666;
assign c9300 =  x171 & ~x121 & ~x554;
assign c9302 =  x81;
assign c9304 = ~x40 & ~x68 & ~x84 & ~x106 & ~x127 & ~x163 & ~x235 & ~x240 & ~x340 & ~x413 & ~x446 & ~x527 & ~x644 & ~x767;
assign c9306 =  x743 &  x772 &  x773 & ~x569 & ~x595;
assign c9308 =  x81;
assign c9310 =  x272 &  x351 & ~x159 & ~x414 & ~x417 & ~x476;
assign c9312 =  x692 & ~x500 & ~x552 & ~x554 & ~x610 & ~x613 & ~x647 & ~x705 & ~x707 & ~x764;
assign c9314 =  x494 & ~x14 & ~x37 & ~x55 & ~x90 & ~x193 & ~x219 & ~x329 & ~x448 & ~x488 & ~x532 & ~x533;
assign c9316 =  x494 & ~x112 & ~x242 & ~x328 & ~x557 & ~x661 & ~x713 & ~x744;
assign c9318 =  x405 & ~x40 & ~x44 & ~x182 & ~x209 & ~x212 & ~x238 & ~x395 & ~x443 & ~x450 & ~x565 & ~x617 & ~x673 & ~x674 & ~x698;
assign c9320 =  x458 &  x595 & ~x154 & ~x155 & ~x225 & ~x692;
assign c9322 =  x212 &  x439 &  x537 & ~x263 & ~x632;
assign c9324 =  x438 & ~x77 & ~x164 & ~x184 & ~x193 & ~x213 & ~x214 & ~x215 & ~x216 & ~x269 & ~x445 & ~x447 & ~x448 & ~x456 & ~x509 & ~x535 & ~x558 & ~x566 & ~x673;
assign c9326 =  x137 &  x240 & ~x124;
assign c9328 =  x380 & ~x101 & ~x121 & ~x135 & ~x209 & ~x235 & ~x239 & ~x263 & ~x414 & ~x536 & ~x537 & ~x683 & ~x772;
assign c9330 =  x594 & ~x171 & ~x235 & ~x290 & ~x478 & ~x615 & ~x689 & ~x713 & ~x717 & ~x763;
assign c9332 = ~x9 & ~x14 & ~x16 & ~x21 & ~x48 & ~x76 & ~x77 & ~x81 & ~x99 & ~x101 & ~x127 & ~x130 & ~x153 & ~x154 & ~x155 & ~x158 & ~x212 & ~x234 & ~x366 & ~x368 & ~x451 & ~x453 & ~x477 & ~x480 & ~x481 & ~x497 & ~x530 & ~x535 & ~x588 & ~x616 & ~x647 & ~x699 & ~x723 & ~x727 & ~x760 & ~x775 & ~x779;
assign c9334 =  x659 &  x660 & ~x68 & ~x94 & ~x444 & ~x648 & ~x672 & ~x759 & ~x772;
assign c9336 =  x321 & ~x153 & ~x154 & ~x368 & ~x426 & ~x622 & ~x674 & ~x772 & ~x773;
assign c9338 =  x178 & ~x17 & ~x290 & ~x346 & ~x442 & ~x480 & ~x605 & ~x706 & ~x737;
assign c9340 =  x414 &  x742 & ~x189 & ~x551 & ~x554 & ~x605;
assign c9342 =  x521 &  x649 & ~x227 & ~x660 & ~x715;
assign c9344 =  x737 &  x769 & ~x240;
assign c9346 =  x413 &  x470 &  x584 & ~x608;
assign c9348 =  x97 &  x741 &  x744 &  x745 & ~x511 & ~x650;
assign c9350 =  x235 &  x742 & ~x133 & ~x239;
assign c9352 =  x610 &  x667 & ~x385;
assign c9354 =  x301 &  x407 & ~x22 & ~x75 & ~x78 & ~x107 & ~x131 & ~x135 & ~x160 & ~x162 & ~x163 & ~x213 & ~x416 & ~x417 & ~x554 & ~x559 & ~x729;
assign c9356 =  x358 &  x384 &  x437 & ~x133 & ~x214 & ~x218;
assign c9358 =  x235 &  x491 &  x745;
assign c9360 =  x469 &  x526 &  x612;
assign c9362 =  x207 &  x517 & ~x73 & ~x163 & ~x213 & ~x216 & ~x523 & ~x610 & ~x632;
assign c9364 =  x461 & ~x46 & ~x182 & ~x240 & ~x593 & ~x605 & ~x650;
assign c9366 =  x191 &  x324 & ~x738;
assign c9368 =  x81 &  x702;
assign c9370 =  x324 & ~x19 & ~x25 & ~x29 & ~x84 & ~x328 & ~x387 & ~x670 & ~x714 & ~x715 & ~x716 & ~x717 & ~x735 & ~x737 & ~x745 & ~x773;
assign c9372 =  x267 &  x296;
assign c9374 =  x118 &  x145 &  x348 &  x376 & ~x68 & ~x281 & ~x561;
assign c9376 =  x386 &  x740 &  x741 &  x743 & ~x607 & ~x610;
assign c9378 =  x646;
assign c9380 =  x439 &  x732;
assign c9382 =  x739 &  x740 &  x742 &  x743 &  x744 & ~x296;
assign c9384 =  x302 & ~x6 & ~x13 & ~x16 & ~x26 & ~x29 & ~x44 & ~x45 & ~x79 & ~x130 & ~x132 & ~x138 & ~x212 & ~x240 & ~x241 & ~x417 & ~x524 & ~x583 & ~x586 & ~x674 & ~x757;
assign c9386 =  x239 &  x565 & ~x234 & ~x302 & ~x634;
assign c9388 =  x235 &  x574 &  x744 & ~x620 & ~x633 & ~x661;
assign c9390 =  x427 &  x536 & ~x474 & ~x551 & ~x558 & ~x607;
assign c9392 =  x494 &  x509 & ~x561;
assign c9394 =  x239 & ~x235 & ~x261 & ~x290 & ~x317 & ~x605 & ~x738 & ~x739 & ~x767;
assign c9396 =  x295 & ~x46 & ~x302 & ~x333 & ~x390 & ~x443 & ~x473 & ~x501 & ~x586 & ~x616 & ~x680 & ~x709 & ~x710 & ~x712 & ~x740 & ~x741;
assign c9398 =  x218 &  x323 &  x324 & ~x333 & ~x385 & ~x443;
assign c9400 =  x137 &  x212;
assign c9402 =  x191 & ~x82 & ~x101 & ~x303 & ~x336 & ~x360 & ~x418 & ~x737 & ~x763;
assign c9404 =  x358 &  x410 & ~x187 & ~x339 & ~x420 & ~x469;
assign c9406 =  x709 &  x715 & ~x16 & ~x240 & ~x265 & ~x294 & ~x554 & ~x582 & ~x607 & ~x619;
assign c9408 =  x468 &  x611 &  x668;
assign c9410 =  x58;
assign c9412 = ~x6 & ~x12 & ~x25 & ~x44 & ~x45 & ~x46 & ~x57 & ~x68 & ~x72 & ~x104 & ~x109 & ~x124 & ~x127 & ~x137 & ~x139 & ~x386 & ~x413 & ~x416 & ~x440 & ~x473 & ~x475 & ~x480 & ~x507 & ~x527 & ~x530 & ~x557 & ~x616 & ~x726 & ~x728 & ~x735 & ~x737 & ~x759 & ~x760;
assign c9414 = ~x171 & ~x188 & ~x214 & ~x240 & ~x375 & ~x395 & ~x400 & ~x401 & ~x402 & ~x484 & ~x511 & ~x513 & ~x553 & ~x565 & ~x612 & ~x763;
assign c9416 =  x660 & ~x132 & ~x212 & ~x468 & ~x501 & ~x619 & ~x647 & ~x713 & ~x739 & ~x740;
assign c9418 =  x510 & ~x58 & ~x234 & ~x290 & ~x304 & ~x389 & ~x444 & ~x445 & ~x504 & ~x558 & ~x632 & ~x717 & ~x735 & ~x775;
assign c9420 =  x273 &  x351 & ~x368 & ~x412 & ~x443 & ~x526 & ~x619;
assign c9422 = ~x36 & ~x46 & ~x74 & ~x77 & ~x102 & ~x109 & ~x124 & ~x127 & ~x129 & ~x152 & ~x183 & ~x421 & ~x444 & ~x585 & ~x593 & ~x666 & ~x679 & ~x699 & ~x703 & ~x737;
assign c9424 =  x681 &  x739 &  x740;
assign c9426 =  x206 &  x517 &  x740 & ~x240 & ~x554;
assign c9428 = ~x24 & ~x68 & ~x77 & ~x127 & ~x153 & ~x393 & ~x469 & ~x529 & ~x555 & ~x680 & ~x682 & ~x705 & ~x779;
assign c9430 =  x143 & ~x586 & ~x605 & ~x613;
assign c9432 =  x742 &  x743 & ~x173 & ~x312 & ~x324 & ~x339 & ~x511 & ~x581 & ~x605 & ~x632;
assign c9434 = ~x9 & ~x26 & ~x44 & ~x46 & ~x68 & ~x80 & ~x94 & ~x99 & ~x121 & ~x127 & ~x128 & ~x149 & ~x237 & ~x239 & ~x293 & ~x452 & ~x533 & ~x563 & ~x582 & ~x584 & ~x614 & ~x705 & ~x732 & ~x769;
assign c9436 =  x468 &  x639;
assign c9438 =  x412 & ~x252 & ~x307 & ~x331 & ~x360 & ~x361 & ~x417 & ~x561 & ~x597 & ~x661 & ~x689 & ~x762;
assign c9440 =  x432 & ~x43 & ~x73 & ~x127 & ~x142 & ~x143 & ~x155 & ~x182 & ~x209 & ~x211 & ~x339 & ~x362 & ~x395 & ~x427 & ~x444 & ~x452 & ~x503 & ~x584 & ~x585 & ~x587 & ~x592 & ~x675 & ~x776;
assign c9442 =  x137 & ~x248;
assign c9444 = ~x127 & ~x175 & ~x186 & ~x216 & ~x235 & ~x236 & ~x763;
assign c9446 =  x274 & ~x127 & ~x159 & ~x239 & ~x443 & ~x477 & ~x554;
assign c9448 = ~x9 & ~x46 & ~x71 & ~x96 & ~x97 & ~x121 & ~x152 & ~x182 & ~x187 & ~x234 & ~x236 & ~x420 & ~x475 & ~x533 & ~x536 & ~x703 & ~x736 & ~x759 & ~x776;
assign c9450 =  x518 &  x716 & ~x402;
assign c9452 =  x69 & ~x77 & ~x164 & ~x238 & ~x593 & ~x607;
assign c9454 =  x740 &  x742 &  x744 & ~x16 & ~x189 & ~x458 & ~x513 & ~x578;
assign c9456 =  x519 &  x742 &  x745 & ~x222 & ~x310 & ~x325 & ~x485 & ~x619;
assign c9458 =  x275 &  x379 & ~x105 & ~x130 & ~x136 & ~x158 & ~x163 & ~x212 & ~x240 & ~x442 & ~x476 & ~x497 & ~x498;
assign c9460 =  x438 & ~x246 & ~x276 & ~x317 & ~x530 & ~x579 & ~x686 & ~x747 & ~x767;
assign c9462 =  x681 &  x712 & ~x182 & ~x223 & ~x392 & ~x523 & ~x554;
assign c9464 =  x438 &  x537 & ~x206 & ~x533 & ~x541;
assign c9466 =  x731;
assign c9468 =  x172 & ~x121 & ~x477 & ~x492 & ~x558;
assign c9470 =  x410 & ~x186 & ~x273 & ~x457 & ~x458 & ~x503;
assign c9472 =  x414 & ~x29 & ~x448 & ~x524 & ~x577;
assign c9474 = ~x74 & ~x101 & ~x155 & ~x210 & ~x212 & ~x240 & ~x241 & ~x430 & ~x470 & ~x511 & ~x533 & ~x622 & ~x650 & ~x728 & ~x739 & ~x758;
assign c9476 =  x352 &  x693 & ~x414 & ~x697 & ~x707;
assign c9478 = ~x53 & ~x76 & ~x183 & ~x190 & ~x210 & ~x212 & ~x240 & ~x241 & ~x339 & ~x401 & ~x429 & ~x456 & ~x534 & ~x538 & ~x558 & ~x610 & ~x614 & ~x618 & ~x636;
assign c9480 =  x273 &  x325 &  x326 & ~x16 & ~x102 & ~x130 & ~x212 & ~x385 & ~x703;
assign c9482 =  x376 & ~x40 & ~x50 & ~x74 & ~x100 & ~x124 & ~x154 & ~x446 & ~x536 & ~x560 & ~x641 & ~x671 & ~x729 & ~x750;
assign c9484 =  x438 & ~x197 & ~x278 & ~x362 & ~x605 & ~x681 & ~x684 & ~x713 & ~x714;
assign c9486 =  x267 &  x409 &  x495 & ~x597;
assign c9488 =  x440 &  x526 & ~x607 & ~x637;
assign c9490 =  x349 &  x460 & ~x76 & ~x182 & ~x414 & ~x773;
assign c9492 =  x609 & ~x735;
assign c9494 =  x716 & ~x346 & ~x400 & ~x511 & ~x605 & ~x644;
assign c9496 =  x468 & ~x7 & ~x55 & ~x476 & ~x478 & ~x571 & ~x597 & ~x636 & ~x652 & ~x662;
assign c9498 =  x207 &  x744 & ~x9 & ~x55 & ~x73 & ~x483 & ~x581;
assign c91 =  x333 & ~x719;
assign c93 =  x205 &  x230 &  x257;
assign c95 =  x576 & ~x5 & ~x83 & ~x447 & ~x476 & ~x487 & ~x502 & ~x514 & ~x532 & ~x582 & ~x610 & ~x724;
assign c97 =  x264 &  x543 & ~x145 & ~x204 & ~x574;
assign c99 =  x98 &  x209;
assign c911 =  x361 & ~x720;
assign c913 =  x94 &  x176 &  x203 &  x204 & ~x417 & ~x666 & ~x697 & ~x699;
assign c915 =  x204 &  x231 &  x257 &  x259 &  x285 & ~x224;
assign c917 =  x529;
assign c919 =  x520 &  x549 &  x576 & ~x81 & ~x333 & ~x526 & ~x645 & ~x696 & ~x727 & ~x757;
assign c921 = ~x3 & ~x138 & ~x141 & ~x281 & ~x387 & ~x434 & ~x435 & ~x460 & ~x461 & ~x462 & ~x479 & ~x575;
assign c923 =  x558;
assign c925 =  x189 & ~x295 & ~x349 & ~x392;
assign c927 =  x100 & ~x527;
assign c929 =  x133 & ~x320 & ~x484 & ~x648;
assign c931 =  x98 &  x237 &  x542 & ~x388;
assign c933 =  x562;
assign c935 =  x160 & ~x377;
assign c937 =  x461 & ~x36 & ~x79 & ~x122 & ~x123 & ~x147 & ~x150 & ~x172 & ~x173 & ~x175 & ~x218 & ~x245 & ~x363 & ~x498 & ~x751 & ~x760 & ~x777;
assign c939 =  x229 &  x506;
assign c941 =  x428 & ~x78 & ~x109 & ~x114 & ~x116 & ~x145 & ~x147 & ~x302 & ~x362 & ~x494 & ~x495 & ~x520;
assign c943 =  x549 &  x682 & ~x724 & ~x758;
assign c945 =  x270 &  x271 & ~x114 & ~x405 & ~x432 & ~x433;
assign c947 = ~x80 & ~x145 & ~x188 & ~x231 & ~x245 & ~x264 & ~x287 & ~x342 & ~x386 & ~x448 & ~x455 & ~x658;
assign c949 =  x602 &  x629 &  x655 &  x656 &  x682;
assign c951 = ~x405 & ~x406 & ~x408 & ~x434 & ~x462 & ~x464 & ~x546 & ~x657;
assign c953 =  x314 &  x318 &  x319 & ~x0 & ~x26 & ~x383 & ~x753;
assign c955 =  x147 &  x174 &  x203 &  x257 & ~x112 & ~x753;
assign c957 =  x555 & ~x327;
assign c959 =  x306 &  x389;
assign c961 =  x529;
assign c963 =  x315 &  x343;
assign c965 =  x259 &  x343 &  x426;
assign c967 =  x513 &  x515 & ~x29 & ~x80 & ~x108 & ~x115 & ~x117 & ~x118 & ~x172 & ~x173 & ~x248 & ~x303 & ~x331 & ~x587 & ~x755;
assign c969 =  x513 &  x514 &  x515 & ~x89 & ~x106 & ~x116 & ~x135 & ~x173 & ~x195 & ~x221 & ~x229 & ~x360 & ~x416 & ~x507;
assign c971 =  x543 &  x570 & ~x4 & ~x48 & ~x60 & ~x86 & ~x110 & ~x118 & ~x159 & ~x172 & ~x192 & ~x220 & ~x254 & ~x303 & ~x305 & ~x362 & ~x414 & ~x417 & ~x444 & ~x559 & ~x727 & ~x757;
assign c973 =  x379 & ~x64 & ~x93 & ~x114 & ~x116 & ~x137 & ~x143 & ~x172 & ~x174 & ~x282 & ~x287 & ~x303 & ~x311 & ~x313 & ~x315 & ~x339 & ~x384 & ~x498 & ~x618 & ~x695 & ~x701 & ~x728;
assign c975 =  x11 &  x542;
assign c977 =  x478;
assign c979 = ~x83 & ~x162 & ~x168 & ~x178 & ~x206 & ~x227 & ~x436 & ~x547 & ~x575;
assign c981 =  x548 &  x687;
assign c983 = ~x327;
assign c985 = ~x31 & ~x113 & ~x149 & ~x172 & ~x173 & ~x174 & ~x205 & ~x284 & ~x562 & ~x579 & ~x746;
assign c987 = ~x113 & ~x406 & ~x433 & ~x434 & ~x460 & ~x461 & ~x462 & ~x470 & ~x489 & ~x546 & ~x627 & ~x628 & ~x756;
assign c989 =  x398 &  x426 &  x454 & ~x641;
assign c991 =  x314 &  x342 &  x426 & ~x82;
assign c993 =  x474;
assign c995 =  x369 &  x480 &  x508;
assign c997 = ~x1 & ~x87 & ~x355 & ~x382 & ~x383 & ~x634 & ~x693 & ~x716 & ~x721 & ~x742;
assign c999 =  x638 &  x664 & ~x222;
assign c9101 =  x314 &  x315 &  x316 &  x317 &  x318;
assign c9103 =  x188 & ~x486;
assign c9105 = ~x12 & ~x57 & ~x168 & ~x208 & ~x292 & ~x382 & ~x439 & ~x486 & ~x514 & ~x719;
assign c9107 =  x581 &  x608 & ~x85 & ~x139 & ~x250 & ~x307;
assign c9109 = ~x5 & ~x6 & ~x22 & ~x62 & ~x82 & ~x89 & ~x116 & ~x137 & ~x149 & ~x150 & ~x189 & ~x206 & ~x226 & ~x231 & ~x248 & ~x259 & ~x272 & ~x277 & ~x280 & ~x286 & ~x303 & ~x312 & ~x331 & ~x332 & ~x339 & ~x441 & ~x502 & ~x554 & ~x728 & ~x750;
assign c9111 =  x181 &  x349 &  x543 & ~x479 & ~x602;
assign c9113 =  x68 &  x463 &  x488 & ~x172;
assign c9115 =  x408 &  x409 & ~x202 & ~x355;
assign c9117 =  x213 &  x241 & ~x172 & ~x257;
assign c9119 = ~x28 & ~x113 & ~x138 & ~x399 & ~x526 & ~x555 & ~x698 & ~x724 & ~x726 & ~x761;
assign c9121 =  x155 & ~x62 & ~x220 & ~x224 & ~x254 & ~x257 & ~x359 & ~x426 & ~x482 & ~x588 & ~x726;
assign c9123 =  x264 &  x487 & ~x206;
assign c9125 = ~x57 & ~x64 & ~x79 & ~x149 & ~x155 & ~x199 & ~x200 & ~x260 & ~x287 & ~x385 & ~x389 & ~x443 & ~x632;
assign c9127 =  x287 &  x288 &  x289 &  x290 & ~x130 & ~x141 & ~x252 & ~x422 & ~x700;
assign c9129 =  x359;
assign c9131 =  x473;
assign c9133 =  x527 &  x554 & ~x221;
assign c9135 =  x407 &  x408 &  x430 & ~x1 & ~x47 & ~x57 & ~x60 & ~x134 & ~x137 & ~x141 & ~x142 & ~x160 & ~x172 & ~x248 & ~x331 & ~x389 & ~x415 & ~x594 & ~x613 & ~x617;
assign c9137 =  x189 & ~x459 & ~x474;
assign c9139 = ~x59 & ~x90 & ~x172 & ~x181 & ~x246 & ~x254 & ~x299 & ~x383 & ~x464 & ~x479 & ~x672 & ~x700 & ~x727 & ~x732 & ~x733 & ~x750 & ~x752 & ~x783;
assign c9141 =  x526 & ~x114 & ~x214 & ~x383 & ~x723;
assign c9143 = ~x47 & ~x62 & ~x89 & ~x171 & ~x172 & ~x200 & ~x270 & ~x271 & ~x299 & ~x327 & ~x382 & ~x438 & ~x465 & ~x474 & ~x495 & ~x576;
assign c9145 =  x550 & ~x45 & ~x112 & ~x113 & ~x366 & ~x398 & ~x555 & ~x643 & ~x670 & ~x723 & ~x732 & ~x750 & ~x752 & ~x755 & ~x762;
assign c9147 =  x554 & ~x52 & ~x71 & ~x165 & ~x333;
assign c9149 =  x662 & ~x56 & ~x60 & ~x172 & ~x173 & ~x227 & ~x501 & ~x749;
assign c9151 =  x160 &  x188 & ~x376;
assign c9153 =  x72 & ~x21 & ~x196 & ~x284 & ~x341 & ~x427 & ~x508 & ~x557 & ~x729;
assign c9155 =  x388 & ~x741 & ~x745;
assign c9157 = ~x406 & ~x434 & ~x461 & ~x462;
assign c9159 = ~x53 & ~x86 & ~x103 & ~x136 & ~x204 & ~x215 & ~x231 & ~x245 & ~x248 & ~x274 & ~x275 & ~x303 & ~x337 & ~x338 & ~x387 & ~x441 & ~x475 & ~x518 & ~x545 & ~x557 & ~x559 & ~x591 & ~x609 & ~x675;
assign c9161 =  x691 &  x719 & ~x5 & ~x62 & ~x76 & ~x86 & ~x89 & ~x113 & ~x131 & ~x361 & ~x613;
assign c9163 =  x393 & ~x79 & ~x716;
assign c9165 =  x375 &  x397 &  x426;
assign c9167 =  x104 & ~x321 & ~x486;
assign c9169 =  x231 &  x257 &  x259 &  x285 & ~x114;
assign c9171 = ~x50 & ~x53 & ~x81 & ~x92 & ~x133 & ~x196 & ~x200 & ~x248 & ~x463 & ~x573 & ~x574 & ~x615 & ~x638 & ~x703;
assign c9173 = ~x164 & ~x166 & ~x172 & ~x177 & ~x178 & ~x200 & ~x271 & ~x315 & ~x356 & ~x564 & ~x665 & ~x695 & ~x720;
assign c9175 =  x213 &  x241 & ~x31 & ~x55 & ~x59 & ~x85 & ~x136 & ~x161 & ~x191 & ~x197 & ~x336;
assign c9177 =  x634 &  x662 & ~x117 & ~x221 & ~x224 & ~x226 & ~x250 & ~x445;
assign c9179 = ~x2 & ~x5 & ~x24 & ~x27 & ~x34 & ~x83 & ~x93 & ~x109 & ~x114 & ~x173 & ~x177 & ~x190 & ~x193 & ~x230 & ~x245 & ~x252 & ~x273 & ~x339 & ~x395 & ~x526 & ~x659 & ~x673 & ~x698 & ~x705 & ~x723;
assign c9181 =  x303 & ~x434;
assign c9183 =  x102 &  x104;
assign c9185 =  x563 & ~x19 & ~x379;
assign c9187 = ~x57 & ~x233 & ~x406 & ~x433 & ~x434 & ~x461 & ~x462 & ~x518 & ~x630 & ~x657;
assign c9189 =  x205 &  x208 & ~x645;
assign c9191 =  x581 & ~x45 & ~x57 & ~x78 & ~x111 & ~x138 & ~x250 & ~x644 & ~x724 & ~x729 & ~x752 & ~x778;
assign c9193 =  x161 & ~x403 & ~x457;
assign c9195 = ~x1 & ~x23 & ~x130 & ~x149 & ~x168 & ~x172 & ~x173 & ~x177 & ~x338 & ~x672 & ~x705 & ~x747 & ~x766;
assign c9197 =  x606 & ~x172;
assign c9199 =  x634 &  x662 & ~x88 & ~x114 & ~x200 & ~x306 & ~x447;
assign c9201 =  x262 & ~x27 & ~x92 & ~x108 & ~x110 & ~x197 & ~x224 & ~x243 & ~x454 & ~x461 & ~x703 & ~x778;
assign c9203 =  x543 & ~x6 & ~x74 & ~x143 & ~x221 & ~x275 & ~x305 & ~x333 & ~x652;
assign c9205 =  x119 &  x147 &  x148 &  x203 & ~x83;
assign c9207 =  x94 &  x208 &  x236;
assign c9209 =  x488 &  x514 &  x515 &  x714 & ~x249 & ~x361 & ~x389;
assign c9211 =  x463 &  x542 &  x543 & ~x164 & ~x166 & ~x173 & ~x199 & ~x228 & ~x229 & ~x254 & ~x274 & ~x331 & ~x332 & ~x367 & ~x642;
assign c9213 =  x342;
assign c9215 =  x161 & ~x405;
assign c9217 =  x71 &  x99 & ~x91 & ~x256 & ~x312 & ~x415;
assign c9219 =  x500 & ~x279;
assign c9221 =  x664 &  x691 & ~x5 & ~x142 & ~x196 & ~x222 & ~x253 & ~x279 & ~x281 & ~x305 & ~x361;
assign c9223 =  x244 & ~x83 & ~x323 & ~x514 & ~x616 & ~x765 & ~x778 & ~x783;
assign c9225 = ~x142 & ~x143 & ~x383 & ~x438 & ~x493 & ~x500 & ~x570 & ~x755 & ~x763;
assign c9227 =  x154 & ~x53 & ~x73 & ~x112 & ~x172 & ~x285 & ~x330 & ~x398 & ~x453 & ~x482 & ~x499 & ~x508 & ~x536 & ~x670 & ~x753 & ~x781;
assign c9229 = ~x3 & ~x8 & ~x58 & ~x62 & ~x379 & ~x382 & ~x463 & ~x702 & ~x713 & ~x754;
assign c9231 =  x183 & ~x174 & ~x284 & ~x286 & ~x453 & ~x509;
assign c9233 =  x443 & ~x742;
assign c9235 =  x678 & ~x406 & ~x434 & ~x489;
assign c9237 =  x619 & ~x82 & ~x166 & ~x435 & ~x729;
assign c9239 =  x176 &  x203 &  x228 &  x229;
assign c9241 =  x677 & ~x57 & ~x462 & ~x490 & ~x517 & ~x600;
assign c9243 =  x343 &  x483 & ~x424;
assign c9245 =  x239 & ~x20 & ~x22 & ~x58 & ~x117 & ~x134 & ~x135 & ~x142 & ~x172 & ~x258 & ~x287 & ~x309 & ~x311 & ~x315 & ~x500 & ~x535 & ~x756;
assign c9247 =  x102 & ~x54 & ~x459 & ~x486 & ~x590 & ~x615;
assign c9249 =  x607 & ~x196 & ~x406 & ~x757 & ~x778;
assign c9251 =  x221 &  x305;
assign c9253 =  x236 &  x405 &  x571 & ~x172 & ~x201 & ~x228;
assign c9255 =  x550 &  x578 & ~x406;
assign c9257 =  x288 &  x344 &  x372 & ~x438;
assign c9259 =  x398 &  x426 &  x454 & ~x10;
assign c9261 =  x35 &  x631;
assign c9263 =  x231 &  x259 &  x287 &  x315 & ~x742;
assign c9265 =  x291 &  x408 &  x430 & ~x359;
assign c9267 = ~x35 & ~x88 & ~x140 & ~x144 & ~x242 & ~x382 & ~x464 & ~x494 & ~x632;
assign c9269 =  x117 &  x313;
assign c9271 = ~x50 & ~x64 & ~x119 & ~x172 & ~x221 & ~x246 & ~x255 & ~x283 & ~x287 & ~x311 & ~x341 & ~x383 & ~x420 & ~x442 & ~x469 & ~x495 & ~x500 & ~x603 & ~x725;
assign c9273 =  x473;
assign c9275 =  x288 &  x400 & ~x62 & ~x89 & ~x170 & ~x726 & ~x778;
assign c9277 = ~x19 & ~x141 & ~x280 & ~x461 & ~x462 & ~x489 & ~x490 & ~x630 & ~x655 & ~x657 & ~x689 & ~x721;
assign c9279 = ~x81 & ~x173 & ~x175 & ~x205 & ~x235 & ~x284 & ~x481 & ~x506 & ~x603 & ~x630;
assign c9281 =  x533;
assign c9283 =  x264 &  x317 & ~x5 & ~x56 & ~x57 & ~x116 & ~x118 & ~x284;
assign c9285 =  x416 & ~x743;
assign c9287 = ~x715;
assign c9289 =  x472;
assign c9291 = ~x35 & ~x57 & ~x59 & ~x89 & ~x436 & ~x437 & ~x462 & ~x518 & ~x547 & ~x630 & ~x658;
assign c9293 =  x444 & ~x715;
assign c9295 =  x550 & ~x19 & ~x24 & ~x84 & ~x86 & ~x116 & ~x191 & ~x366 & ~x427 & ~x531 & ~x639 & ~x641 & ~x693 & ~x701 & ~x758;
assign c9297 =  x176 &  x230 &  x257 & ~x355 & ~x664;
assign c9299 =  x505;
assign c9301 =  x241;
assign c9303 = ~x2 & ~x44 & ~x99 & ~x107 & ~x114 & ~x165 & ~x166 & ~x193 & ~x362 & ~x461 & ~x462 & ~x487 & ~x489 & ~x490 & ~x625 & ~x726 & ~x754;
assign c9305 =  x664 & ~x378 & ~x461;
assign c9307 =  x550 & ~x32 & ~x56 & ~x434 & ~x435 & ~x461 & ~x462 & ~x463 & ~x781;
assign c9309 =  x576 &  x688 & ~x4 & ~x85 & ~x114 & ~x613 & ~x643 & ~x672;
assign c9311 =  x289 &  x292 & ~x405;
assign c9313 =  x152 &  x430;
assign c9315 =  x293 & ~x147 & ~x172 & ~x355 & ~x482;
assign c9317 = ~x19 & ~x22 & ~x31 & ~x35 & ~x47 & ~x119 & ~x158 & ~x189 & ~x223 & ~x236 & ~x279 & ~x303 & ~x307 & ~x335 & ~x355 & ~x366 & ~x383 & ~x384 & ~x393 & ~x449 & ~x452 & ~x468 & ~x502 & ~x552 & ~x587 & ~x613 & ~x643 & ~x644 & ~x652 & ~x672 & ~x695 & ~x729 & ~x749 & ~x761;
assign c9319 =  x44 & ~x147;
assign c9321 =  x520 &  x631 & ~x433;
assign c9323 =  x714 & ~x5 & ~x91 & ~x103 & ~x173 & ~x204 & ~x228 & ~x383 & ~x386 & ~x529 & ~x592;
assign c9325 = ~x23 & ~x26 & ~x75 & ~x85 & ~x112 & ~x134 & ~x142 & ~x147 & ~x162 & ~x189 & ~x203 & ~x217 & ~x224 & ~x228 & ~x286 & ~x287 & ~x288 & ~x327 & ~x357 & ~x507 & ~x509 & ~x587 & ~x674;
assign c9327 =  x244 & ~x225 & ~x323;
assign c9329 =  x213 &  x353 & ~x250 & ~x511 & ~x562;
assign c9331 =  x221 &  x305;
assign c9333 =  x233 &  x344 &  x372 & ~x72 & ~x224 & ~x783;
assign c9335 =  x64 &  x92 &  x93 &  x121 &  x149;
assign c9337 =  x151 &  x428 & ~x5 & ~x332 & ~x415 & ~x500 & ~x527 & ~x535 & ~x562 & ~x696;
assign c9339 = ~x80 & ~x143 & ~x364 & ~x377 & ~x387 & ~x393 & ~x405 & ~x406 & ~x479 & ~x547 & ~x755;
assign c9341 =  x361;
assign c9343 =  x582 & ~x15 & ~x83 & ~x102 & ~x108 & ~x135 & ~x189 & ~x191 & ~x221 & ~x250 & ~x394;
assign c9345 = ~x104 & ~x110 & ~x122 & ~x166 & ~x195 & ~x203 & ~x221 & ~x225 & ~x231 & ~x248 & ~x252 & ~x279 & ~x287 & ~x481 & ~x559 & ~x575 & ~x594 & ~x722;
assign c9347 =  x445;
assign c9349 =  x306 &  x390;
assign c9351 = ~x3 & ~x59 & ~x64 & ~x81 & ~x82 & ~x114 & ~x168 & ~x194 & ~x216 & ~x224 & ~x308 & ~x327 & ~x364 & ~x382 & ~x438 & ~x439 & ~x466 & ~x493 & ~x494 & ~x528 & ~x549 & ~x584 & ~x643 & ~x645 & ~x726 & ~x759;
assign c9353 =  x154 &  x210 & ~x33 & ~x76 & ~x143 & ~x281 & ~x385 & ~x386;
assign c9355 =  x41 &  x487 & ~x77 & ~x202 & ~x222;
assign c9357 = ~x25 & ~x36 & ~x48 & ~x49 & ~x52 & ~x57 & ~x63 & ~x76 & ~x106 & ~x133 & ~x137 & ~x139 & ~x171 & ~x173 & ~x196 & ~x221 & ~x247 & ~x248 & ~x278 & ~x287 & ~x313 & ~x314 & ~x369 & ~x370 & ~x371 & ~x451 & ~x474 & ~x480 & ~x481 & ~x485 & ~x507 & ~x531 & ~x616 & ~x646 & ~x674 & ~x675 & ~x676 & ~x728 & ~x729 & ~x752;
assign c9359 = ~x29 & ~x144 & ~x165 & ~x223 & ~x435 & ~x461 & ~x462 & ~x489 & ~x517 & ~x628 & ~x685;
assign c9361 = ~x57 & ~x86 & ~x168 & ~x379 & ~x406 & ~x435 & ~x436 & ~x518 & ~x587 & ~x689;
assign c9363 = ~x19 & ~x54 & ~x80 & ~x138 & ~x205 & ~x462 & ~x489 & ~x490 & ~x576 & ~x600 & ~x601 & ~x603 & ~x657;
assign c9365 =  x550 &  x578 & ~x77 & ~x197 & ~x200 & ~x225 & ~x228 & ~x249 & ~x254;
assign c9367 = ~x205 & ~x233 & ~x359 & ~x379 & ~x406 & ~x434 & ~x436 & ~x546 & ~x547;
assign c9369 =  x556;
assign c9371 =  x638 &  x664;
assign c9373 =  x119 &  x120 &  x148 &  x149 &  x575;
assign c9375 =  x305 & ~x611 & ~x637 & ~x720;
assign c9377 =  x155 & ~x0 & ~x86 & ~x117 & ~x172 & ~x415 & ~x474 & ~x508 & ~x528 & ~x529 & ~x609 & ~x720 & ~x753 & ~x777;
assign c9379 =  x180 &  x208 &  x430 & ~x201;
assign c9381 =  x317 &  x342;
assign c9383 =  x343 &  x454;
assign c9385 = ~x280 & ~x379 & ~x406 & ~x432 & ~x433 & ~x434 & ~x657 & ~x762;
assign c9387 = ~x27 & ~x51 & ~x56 & ~x80 & ~x83 & ~x406 & ~x434 & ~x436 & ~x461 & ~x462 & ~x463 & ~x575 & ~x576 & ~x629;
assign c9389 = ~x2 & ~x30 & ~x33 & ~x49 & ~x53 & ~x103 & ~x117 & ~x129 & ~x134 & ~x135 & ~x139 & ~x141 & ~x147 & ~x159 & ~x166 & ~x172 & ~x188 & ~x196 & ~x199 & ~x219 & ~x221 & ~x227 & ~x229 & ~x251 & ~x252 & ~x254 & ~x270 & ~x276 & ~x278 & ~x286 & ~x302 & ~x311 & ~x312 & ~x314 & ~x340 & ~x363 & ~x367 & ~x389 & ~x393 & ~x414 & ~x444 & ~x468 & ~x471 & ~x479 & ~x509 & ~x533 & ~x588 & ~x602 & ~x619 & ~x647 & ~x669 & ~x672 & ~x700 & ~x727 & ~x730 & ~x759 & ~x778 & ~x782;
assign c9391 =  x550 & ~x109 & ~x282 & ~x372 & ~x394;
assign c9393 =  x533;
assign c9395 =  x183 & ~x64 & ~x133 & ~x172 & ~x202 & ~x284;
assign c9397 =  x174 &  x229 &  x230 & ~x406 & ~x435;
assign c9399 =  x305 & ~x326 & ~x383 & ~x690;
assign c9401 =  x428 &  x435 & ~x133 & ~x147 & ~x172 & ~x387 & ~x467;
assign c9403 = ~x64 & ~x141 & ~x161 & ~x165 & ~x190 & ~x226 & ~x433 & ~x434 & ~x435 & ~x441 & ~x726;
assign c9405 =  x151 &  x152 &  x175 &  x204 & ~x140 & ~x280 & ~x361 & ~x477 & ~x505 & ~x642 & ~x696 & ~x725 & ~x726 & ~x730;
assign c9407 =  x355 & ~x166 & ~x435 & ~x436 & ~x462 & ~x489;
assign c9409 =  x241 &  x270 & ~x24 & ~x78 & ~x103 & ~x115 & ~x166 & ~x755;
assign c9411 = ~x0 & ~x24 & ~x62 & ~x88 & ~x115 & ~x174 & ~x177 & ~x193 & ~x194 & ~x200 & ~x203 & ~x223 & ~x229 & ~x248 & ~x255 & ~x259 & ~x260 & ~x286 & ~x360 & ~x481 & ~x482 & ~x621 & ~x665 & ~x666 & ~x675 & ~x730 & ~x778;
assign c9413 = ~x97 & ~x142 & ~x147 & ~x172 & ~x203 & ~x233;
assign c9415 =  x216 & ~x56 & ~x321 & ~x529;
assign c9417 =  x288 &  x428 & ~x17 & ~x705;
assign c9419 =  x539 &  x540 & ~x1 & ~x131 & ~x307 & ~x389 & ~x576;
assign c9421 =  x94 &  x233 & ~x200 & ~x777;
assign c9423 = ~x31 & ~x82 & ~x110 & ~x360 & ~x379 & ~x406 & ~x421 & ~x423 & ~x432 & ~x433 & ~x434 & ~x450 & ~x470 & ~x471 & ~x560 & ~x576 & ~x604 & ~x727 & ~x754;
assign c9425 =  x577 & ~x580 & ~x718 & ~x750;
assign c9427 =  x520 &  x631 & ~x30 & ~x31 & ~x196 & ~x253 & ~x668 & ~x721;
assign c9429 =  x361;
assign c9431 =  x154 &  x210 & ~x31 & ~x139 & ~x172 & ~x219 & ~x221 & ~x229 & ~x287;
assign c9433 =  x608 & ~x53 & ~x351;
assign c9435 =  x473;
assign c9437 =  x408 & ~x116 & ~x119 & ~x137 & ~x142 & ~x147 & ~x164 & ~x172 & ~x173 & ~x176 & ~x188 & ~x194 & ~x199 & ~x246 & ~x256 & ~x287 & ~x315 & ~x331 & ~x481 & ~x728 & ~x775;
assign c9439 = ~x33 & ~x55 & ~x59 & ~x61 & ~x65 & ~x82 & ~x116 & ~x192 & ~x196 & ~x198 & ~x200 & ~x221 & ~x227 & ~x230 & ~x245 & ~x247 & ~x248 & ~x254 & ~x259 & ~x287 & ~x304 & ~x328 & ~x359 & ~x371 & ~x384 & ~x394 & ~x423 & ~x443 & ~x447 & ~x471 & ~x481 & ~x560 & ~x581 & ~x587 & ~x590 & ~x640 & ~x650 & ~x692 & ~x704 & ~x723 & ~x724 & ~x755 & ~x762;
assign c9441 =  x152 &  x153 &  x355 & ~x171 & ~x697;
assign c9443 =  x555 & ~x221 & ~x384;
assign c9445 =  x352 & ~x62 & ~x149 & ~x172 & ~x204 & ~x257 & ~x260 & ~x366;
assign c9447 =  x608 &  x647;
assign c9449 = ~x52 & ~x57 & ~x166 & ~x204 & ~x435 & ~x461 & ~x462 & ~x656;
assign c9451 =  x217 & ~x25 & ~x252 & ~x461;
assign c9453 =  x266 & ~x86 & ~x91 & ~x105 & ~x108 & ~x122 & ~x135 & ~x188 & ~x189 & ~x199 & ~x255 & ~x259 & ~x273 & ~x414 & ~x420 & ~x442 & ~x455 & ~x564 & ~x669 & ~x732;
assign c9455 =  x233 &  x575 &  x603 & ~x280 & ~x720 & ~x778;
assign c9457 =  x42 &  x99 & ~x442;
assign c9459 =  x375 & ~x92 & ~x258 & ~x273 & ~x287 & ~x315;
assign c9461 = ~x58 & ~x64 & ~x74 & ~x93 & ~x102 & ~x117 & ~x172 & ~x173 & ~x193 & ~x202 & ~x204 & ~x222 & ~x245 & ~x248 & ~x253 & ~x257 & ~x275 & ~x288 & ~x414 & ~x482 & ~x567 & ~x592 & ~x594 & ~x632 & ~x696 & ~x721 & ~x730 & ~x732 & ~x775;
assign c9463 =  x374 &  x375 &  x408 & ~x116 & ~x229 & ~x274 & ~x315;
assign c9465 =  x12 & ~x45;
assign c9467 =  x687 & ~x4 & ~x25 & ~x30 & ~x32 & ~x59 & ~x86 & ~x225 & ~x247 & ~x255 & ~x276 & ~x283 & ~x609 & ~x615 & ~x640 & ~x645 & ~x655 & ~x670 & ~x726 & ~x729 & ~x731 & ~x732 & ~x733 & ~x750;
assign c9469 = ~x29 & ~x34 & ~x80 & ~x83 & ~x86 & ~x117 & ~x122 & ~x131 & ~x134 & ~x172 & ~x173 & ~x195 & ~x233 & ~x255 & ~x260 & ~x287 & ~x303 & ~x456 & ~x470 & ~x499 & ~x618 & ~x649 & ~x734 & ~x755;
assign c9471 =  x293 & ~x53 & ~x62 & ~x91 & ~x103 & ~x116 & ~x147 & ~x161 & ~x172 & ~x225 & ~x230 & ~x254 & ~x258 & ~x311 & ~x670 & ~x721 & ~x752;
assign c9473 =  x578 &  x606 & ~x141 & ~x376 & ~x389 & ~x721 & ~x725 & ~x777;
assign c9475 =  x236 &  x260 &  x288 & ~x30 & ~x161 & ~x197 & ~x778;
assign c9477 =  x70 &  x98 & ~x203;
assign c9479 =  x68 &  x208 &  x264;
assign c9481 =  x375 & ~x32 & ~x147 & ~x166 & ~x172 & ~x173 & ~x383;
assign c9483 =  x293 & ~x118 & ~x494 & ~x693;
assign c9485 =  x173 & ~x389 & ~x432 & ~x433;
assign c9487 =  x258 &  x314 &  x342 &  x371 & ~x23 & ~x554 & ~x667;
assign c9489 =  x294 & ~x119 & ~x314 & ~x339 & ~x355 & ~x383;
assign c9491 =  x547 &  x548 &  x631 & ~x142 & ~x746;
assign c9493 =  x619 &  x638;
assign c9495 =  x298 & ~x83 & ~x86 & ~x136 & ~x140 & ~x249 & ~x275 & ~x359 & ~x395 & ~x433 & ~x727;
assign c9497 =  x73 & ~x198 & ~x543;
assign c9499 =  x606 &  x661 & ~x23 & ~x142 & ~x167 & ~x191 & ~x363 & ~x376;

endmodule