module tm( x0,x1,x2,x3,x4,x5,x6,x7,x8,x9,x10,x11,x12,x13,x14,x15,x16,x17,x18,x19,x20,x21,x22,x23,x24,x25,x26,x27,x28,x29,x30,x31,x32,x33,x34,x35,x36,x37,x38,x39,x40,x41,x42,x43,x44,x45,x46,x47,x48,x49,x50,x51,x52,x53,x54,x55,x56,x57,x58,x59,x60,x61,x62,x63,x64,x65,x66,x67,x68,x69,x70,x71,x72,x73,x74,x75,x76,x77,x78,x79,x80,x81,x82,x83,x84,x85,x86,x87,x88,x89,x90,x91,x92,x93,x94,x95,x96,x97,x98,x99,x100,x101,x102,x103,x104,x105,x106,x107,x108,x109,x110,x111,x112,x113,x114,x115,x116,x117,x118,x119,x120,x121,x122,x123,x124,x125,x126,x127,x128,x129,x130,x131,x132,x133,x134,x135,x136,x137,x138,x139,x140,x141,x142,x143,x144,x145,x146,x147,x148,x149,x150,x151,x152,x153,x154,x155,x156,x157,x158,x159,x160,x161,x162,x163,x164,x165,x166,x167,x168,x169,x170,x171,x172,x173,x174,x175,x176,x177,x178,x179,x180,x181,x182,x183,x184,x185,x186,x187,x188,x189,x190,x191,x192,x193,x194,x195,x196,x197,x198,x199,x200,x201,x202,x203,x204,x205,x206,x207,x208,x209,x210,x211,x212,x213,x214,x215,x216,x217,x218,x219,x220,x221,x222,x223,x224,x225,x226,x227,x228,x229,x230,x231,x232,x233,x234,x235,x236,x237,x238,x239,x240,x241,x242,x243,x244,x245,x246,x247,x248,x249,x250,x251,x252,x253,x254,x255,x256,x257,x258,x259,x260,x261,x262,x263,x264,x265,x266,x267,x268,x269,x270,x271,x272,x273,x274,x275,x276,x277,x278,x279,x280,x281,x282,x283,x284,x285,x286,x287,x288,x289,x290,x291,x292,x293,x294,x295,x296,x297,x298,x299,x300,x301,x302,x303,x304,x305,x306,x307,x308,x309,x310,x311,x312,x313,x314,x315,x316,x317,x318,x319,x320,x321,x322,x323,x324,x325,x326,x327,x328,x329,x330,x331,x332,x333,x334,x335,x336,x337,x338,x339,x340,x341,x342,x343,x344,x345,x346,x347,x348,x349,x350,x351,x352,x353,x354,x355,x356,x357,x358,x359,x360,x361,x362,x363,x364,x365,x366,x367,x368,x369,x370,x371,x372,x373,x374,x375,x376,x377,x378,x379,x380,x381,x382,x383,x384,x385,x386,x387,x388,x389,x390,x391,x392,x393,x394,x395,x396,x397,x398,x399,x400,x401,x402,x403,x404,x405,x406,x407,x408,x409,x410,x411,x412,x413,x414,x415,x416,x417,x418,x419,x420,x421,x422,x423,x424,x425,x426,x427,x428,x429,x430,x431,x432,x433,x434,x435,x436,x437,x438,x439,x440,x441,x442,x443,x444,x445,x446,x447,x448,x449,x450,x451,x452,x453,x454,x455,x456,x457,x458,x459,x460,x461,x462,x463,x464,x465,x466,x467,x468,x469,x470,x471,x472,x473,x474,x475,x476,x477,x478,x479,x480,x481,x482,x483,x484,x485,x486,x487,x488,x489,x490,x491,x492,x493,x494,x495,x496,x497,x498,x499,x500,x501,x502,x503,x504,x505,x506,x507,x508,x509,x510,x511,x512,x513,x514,x515,x516,x517,x518,x519,x520,x521,x522,x523,x524,x525,x526,x527,x528,x529,x530,x531,x532,x533,x534,x535,x536,x537,x538,x539,x540,x541,x542,x543,x544,x545,x546,x547,x548,x549,x550,x551,x552,x553,x554,x555,x556,x557,x558,x559,x560,x561,x562,x563,x564,x565,x566,x567,x568,x569,x570,x571,x572,x573,x574,x575,x576,x577,x578,x579,x580,x581,x582,x583,x584,x585,x586,x587,x588,x589,x590,x591,x592,x593,x594,x595,x596,x597,x598,x599,x600,x601,x602,x603,x604,x605,x606,x607,x608,x609,x610,x611,x612,x613,x614,x615,x616,x617,x618,x619,x620,x621,x622,x623,x624,x625,x626,x627,x628,x629,x630,x631,x632,x633,x634,x635,x636,x637,x638,x639,x640,x641,x642,x643,x644,x645,x646,x647,x648,x649,x650,x651,x652,x653,x654,x655,x656,x657,x658,x659,x660,x661,x662,x663,x664,x665,x666,x667,x668,x669,x670,x671,x672,x673,x674,x675,x676,x677,x678,x679,x680,x681,x682,x683,x684,x685,x686,x687,x688,x689,x690,x691,x692,x693,x694,x695,x696,x697,x698,x699,x700,x701,x702,x703,x704,x705,x706,x707,x708,x709,x710,x711,x712,x713,x714,x715,x716,x717,x718,x719,x720,x721,x722,x723,x724,x725,x726,x727,x728,x729,x730,x731,x732,x733,x734,x735,x736,x737,x738,x739,x740,x741,x742,x743,x744,x745,x746,x747,x748,x749,x750,x751,x752,x753,x754,x755,x756,x757,x758,x759,x760,x761,x762,x763,x764,x765,x766,x767,x768,x769,x770,x771,x772,x773,x774,x775,x776,x777,x778,x779,x780,x781,x782,x783,c589,c358,c9206,c9145,c0266,c4450,c4198,c866,c238,c4366,c46,c4200,c4245,c2300,c3445,c853,c1158,c8460,c6341,c8426,c1136,c8154,c6181,c4255,c7131,c2379,c6176,c5374,c4234,c5105,c8371,c556,c6487,c9484,c013,c6146,c4168,c1223,c1188,c6142,c1103,c8326,c7248,c4437,c8354,c0395,c436,c3197,c4364,c6104,c2369,c6359,c3356,c5328,c0263,c1201,c4120,c5144,c9406,c9148,c060,c6351,c444,c8373,c1347,c7318,c0427,c1408,c4339,c322,c3119,c170,c1303,c7147,c8374,c5122,c3241,c366,c5248,c3420,c9414,c8477,c7490,c3255,c522,c8203,c8257,c464,c1340,c735,c257,c8343,c5241,c3310,c4227,c6238,c917,c9370,c9472,c7339,c1395,c7259,c193,c382,c4337,c3279,c154,c3144,c3386,c4203,c4469,c656,c4386,c9162,c9386,c7185,c7300,c1239,c7260,c8107,c6321,c4359,c467,c05,c3299,c1266,c6375,c5138,c0216,c8166,c2295,c7448,c7310,c3428,c558,c5312,c1454,c7342,c9300,c138,c6133,c9280,c2135,c985,c198,c4361,c3315,c5239,c1229,c8486,c3271,c21,c6335,c4135,c4340,c6305,c1345,c2340,c3160,c2107,c7438,c9363,c3141,c3475,c1321,c2333,c945,c1270,c5311,c7221,c1221,c3457,c6271,c8199,c8481,c0259,c0445,c4147,c7333,c8234,c958,c2471,c3125,c2271,c7236,c3341,c1182,c5378,c1278,c2472,c6132,c1189,c139,c1210,c9368,c0375,c225,c1152,c9102,c26,c4451,c5371,c8182,c3198,c8494,c3246,c9244,c062,c4257,c7328,c159,c4300,c5207,c2294,c4122,c9413,c6371,c0223,c7369,c1373,c3196,c758,c0440,c454,c9242,c6463,c3109,c2397,c9197,c4299,c2415,c734,c1234,c9402,c5247,c6431,c18,c1301,c9364,c037,c4474,c221,c3164,c8312,c3371,c0424,c3161,c2202,c7110,c9417,c9170,c5411,c3214,c3333,c44,c4150,c8489,c2342,c9291,c4490,c5304,c2368,c9313,c5391,c819,c8475,c2498,c5359,c5481,c399,c4156,c6319,c799,c4144,c622,c3330,c2386,c6159,c9105,c5268,c0264,c6157,c8324,c89,c4455,c379,c8216,c317,c0116,c9201,c7184,c854,c5394,c2217,c920,c3339,c6189,c883,c6410,c0250,c0277,c2289,c9371,c6265,c3469,c3297,c6420,c5271,c9344,c0207,c045,c2444,c3413,c4113,c0385,c649,c8122,c870,c0157,c5178,c3408,c3184,c0473,c4205,c1350,c9274,c7442,c6414,c5159,c6389,c9412,c1416,c2388,c9432,c0342,c0186,c529,c671,c3298,c7365,c4402,c0370,c2182,c9378,c5305,c7351,c0299,c9311,c7439,c0413,c4355,c0396,c7467,c0346,c9114,c8280,c0195,c2452,c6120,c1330,c3238,c5353,c9230,c2218,c1241,c5262,c9196,c6151,c061,c6369,c5367,c0188,c5284,c8193,c49,c0106,c0338,c8104,c5339,c1410,c9222,c5297,c7194,c09,c9106,c867,c5167,c6273,c6210,c8283,c3499,c10,c9192,c4470,c6459,c6179,c891,c4466,c473,c2175,c2164,c433,c772,c4492,c244,c2367,c5211,c1101,c9250,c0241,c339,c2328,c5434,c8248,c478,c7232,c9257,c1110,c886,c67,c7322,c7116,c6388,c7413,c1319,c3273,c2149,c7319,c4212,c2381,c7266,c6400,c5377,c091,c1276,c5116,c3376,c579,c1339,c447,c5379,c6158,c1230,c4426,c2339,c7235,c3100,c3192,c6144,c7405,c6274,c1124,c0465,c0171,c0466,c547,c41,c7454,c158,c1310,c9182,c3444,c7287,c3105,c115,c3169,c6308,c6390,c3433,c1277,c9316,c4454,c022,c2222,c4127,c6342,c0365,c5149,c6366,c3322,c2301,c0148,c1362,c0129,c7384,c1121,c1199,c195,c6428,c4447,c0391,c7227,c192,c6258,c7483,c4171,c9403,c6486,c0232,c0136,c2267,c822,c4435,c0107,c7479,c923,c9171,c8204,c9237,c8398,c514,c1462,c2338,c6154,c6395,c8279,c2396,c6290,c4248,c455,c3128,c1443,c5356,c8288,c1120,c685,c775,c6294,c6362,c4190,c5404,c850,c9463,c581,c8289,c657,c79,c1445,c3436,c0209,c4219,c5263,c8227,c181,c7278,c9129,c4380,c6165,c9465,c5321,c4411,c6278,c6227,c8410,c392,c6344,c7226,c4174,c611,c4397,c8125,c8316,c911,c641,c9352,c5101,c9252,c252,c0360,c9308,c9430,c5476,c285,c0435,c6222,c9419,c3139,c9477,c8113,c5276,c6328,c0336,c2305,c0316,c4475,c7499,c7299,c8442,c6111,c8146,c0423,c6424,c5484,c7453,c2211,c4347,c7421,c1132,c7228,c8269,c3344,c0459,c542,c5322,c227,c8483,c5117,c8386,c1272,c2306,c5383,c8273,c0450,c827,c027,c0282,c5425,c4464,c7320,c4157,c9392,c345,c5317,c2195,c8425,c3275,c6364,c0302,c2291,c9442,c0133,c9218,c6141,c2303,c3449,c4365,c3200,c9464,c6195,c8328,c1313,c162,c1459,c549,c7166,c6322,c4181,c5290,c452,c928,c6445,c2242,c2167,c9101,c1258,c2349,c3257,c1232,c3248,c184,c7494,c5226,c816,c2274,c2102,c0353,c4356,c124,c6438,c9122,c8159,c1105,c4104,c2470,c237,c0397,c8195,c8349,c9333,c3290,c3425,c173,c6262,c4210,c258,c331,c386,c7482,c6163,c6481,c270,c562,c80,c5454,c95,c2207,c215,c0230,c8201,c8402,c3423,c8119,c145,c25,c8342,c2214,c5196,c6303,c640,c8361,c924,c2170,c3254,c2282,c7231,c0235,c9358,c4211,c8152,c1325,c0412,c6356,c487,c4324,c341,c0415,c3353,c1418,c1176,c5292,c058,c1100,c5291,c066,c052,c5361,c9314,c164,c678,c969,c1337,c986,c1379,c3461,c2288,c9318,c8352,c873,c7106,c4155,c28,c6187,c034,c990,c981,c8242,c7269,c463,c155,c5435,c5181,c4213,c3447,c9429,c1141,c8191,c7493,c9362,c5243,c1288,c3217,c8330,c863,c9359,c185,c4379,c362,c0482,c9306,c5352,c4390,c5384,c7476,c1218,c0165,c3334,c4363,c9469,c729,c17,c7271,c9110,c537,c1102,c6310,c2419,c2357,c5256,c4348,c43,c6145,c7464,c451,c8169,c8416,c2276,c2356,c5465,c5183,c7216,c3486,c1284,c367,c2421,c5238,c2151,c594,c4271,c1185,c661,c7262,c177,c1336,c9381,c1329,c0348,c438,c8311,c2366,c672,c2255,c5137,c4407,c3230,c9294,c3368,c2162,c6429,c9135,c127,c471,c8215,c948,c913,c1430,c9437,c8480,c3153,c773,c9273,c180,c4246,c5209,c8190,c5233,c8112,c0152,c1449,c6138,c5408,c9158,c7425,c5327,c6462,c7414,c5429,c1131,c5331,c0254,c4459,c6396,c1363,c5237,c6108,c1151,c4121,c183,c415,c9346,c1499,c6134,c4375,c9144,c2476,c4336,c1178,c9277,c1314,c1403,c0406,c218,c043,c7282,c893,c2129,c019,c683,c075,c621,c7441,c7422,c0287,c0301,c1437,c6323,c134,c6409,c0199,c2484,c9271,c565,c6149,c3207,c7459,c6105,c9130,c9492,c297,c0341,c414,c6192,c0490,c9104,c5494,c3314,c8116,c6401,c8213,c8249,c7160,c7465,c699,c298,c6218,c798,c0221,c2375,c4373,c6427,c140,c6169,c1296,c3189,c15,c088,c0382,c1381,c876,c6374,c1334,c482,c9426,c5451,c0326,c835,c8235,c0184,c4116,c64,c456,c7186,c0108,c3464,c3490,c9431,c378,c1451,c3243,c7100,c214,c7325,c4258,c9498,c3406,c8222,c5457,c6307,c8239,c9441,c2469,c75,c384,c9168,c4305,c1448,c4184,c4270,c561,c5169,c3131,c1485,c1260,c336,c494,c6360,c3427,c2461,c7156,c6152,c9157,c7433,c0163,c9155,c5370,c5388,c32,c9276,c849,c8180,c0357,c9217,c1190,c9467,c462,c6117,c453,c1414,c4341,c8210,c7280,c4484,c0121,c6119,c217,c1328,c4416,c83,c5333,c5498,c3276,c3385,c8189,c1467,c7449,c7143,c3201,c1281,c9375,c9478,c829,c2206,c8315,c4272,c66,c6408,c8382,c3155,c9137,c4256,c7332,c91,c5264,c7212,c833,c2464,c7387,c755,c2401,c7230,c9350,c4408,c1349,c5336,c06,c031,c728,c3326,c9483,c9440,c5344,c4240,c9423,c3381,c5376,c9332,c5395,c8135,c4228,c023,c691,c7406,c4206,c8114,c5398,c5401,c970,c8132,c3263,c796,c0364,c9156,c8344,c6340,c3389,c8117,c9424,c8131,c2361,c4225,c6256,c840,c914,c6475,c090,c9113,c1366,c0238,c7289,c3234,c3317,c3283,c1423,c7305,c7265,c8446,c4449,c3231,c086,c618,c2402,c2299,c5278,c523,c288,c3468,c3233,c9160,c0283,c4215,c5469,c1469,c1364,c9215,c588,c2408,c3439,c814,c5309,c5488,c6407,c7373,c4362,c3471,c9287,c5269,c2191,c1205,c8261,c788,c3250,c7334,c4382,c7285,c3411,c5135,c1390,c3154,c4441,c347,c8493,c0334,c0102,c499,c6276,c7213,c5208,c9210,c489,c96,c8142,c879,c0434,c2387,c9216,c6302,c2181,c0272,c951,c882,c2380,c2293,c3440,c8453,c5382,c1356,c0322,c6337,c5121,c655,c7119,c9163,c042,c6196,c1487,c493,c0208,c5141,c6259,c0497,c531,c8276,c9147,c9126,c2481,c5157,c6136,c3467,c432,c637,c9108,c2235,c2185,c4247,c2443,c6251,c369,c8424,c9283,c9482,c6143,c488,c3208,c4180,c3302,c6211,c570,c3218,c1386,c0476,c9260,c8441,c2404,c7208,c6468,c5172,c6365,c745,c2395,c5282,c8285,c5258,c1464,c20,c0320,c1139,c6288,c8338,c2315,c5217,c5340,c3492,c8270,c8259,c8336,c0369,c7209,c38,c0442,c0297,c169,c643,c0131,c0202,c659,c064,c370,c4401,c5129,c1119,c4141,c5330,c716,c5179,c4413,c2492,c7402,c448,c4383,c860,c2103,c8457,c1442,c1252,c0246,c3289,c3390,c4499,c3476,c2418,c789,c0194,c2493,c0444,c54,c3366,c7331,c563,c7171,c8452,c1153,c4478,c082,c6406,c248,c0408,c4238,c4126,c517,c3260,c5474,c8167,c7376,c2341,c6197,c4387,c6405,c1248,c6411,c0352,c3282,c2374,c3143,c7254,c832,c093,c0256,c2482,c5493,c27,c636,c780,c5274,c8110,c9384,c7327,c3113,c3288,c0261,c111,c0340,c5492,c3338,c597,c5369,c8439,c0447,c3117,c4360,c9136,c892,c4376,c437,c7218,c2264,c9462,c711,c4163,c3474,c7257,c0167,c5446,c8357,c8440,c7272,c865,c1179,c398,c4152,c7153,c3280,c0495,c2101,c5130,c1377,c6373,c0144,c2497,c8395,c3194,c190,c1491,c626,c495,c8293,c5229,c8109,c5485,c275,c9220,c5146,c8474,c995,c1419,c686,c6284,c8447,c3478,c4302,c8103,c9154,c9427,c063,c0178,c2156,c1365,c0237,c7313,c2158,c2209,c2355,c7463,c669,c8495,c0123,c0298,c2358,c4400,c9443,c974,c271,c1480,c2163,c7484,c653,c239,c0253,c165,c4403,c4396,c7233,c9118,c443,c548,c6147,c3309,c0337,c5176,c2337,c1173,c4280,c3183,c898,c8368,c3195,c45,c8198,c038,c360,c2463,c1374,c329,c0127,c5273,c146,c3300,c2316,c7137,c9336,c6190,c4453,c0488,c7193,c191,c8144,c29,c8484,c1264,c0117,c025,c3348,c6301,c080,c5473,c615,c2168,c6416,c7154,c1461,c4137,c4119,c1285,c6343,c9111,c1392,c6399,c0425,c0489,c3272,c2194,c4105,c4217,c7237,c6432,c697,c593,c9416,c823,c7337,c5109,c627,c2430,c7316,c256,c5477,c4175,c7105,c1287,c6476,c0471,c587,c4315,c0234,c2383,c1441,c0174,c3228,c2286,c2221,c187,c0168,c4434,c33,c0191,c355,c017,c3479,c8304,c6398,c8174,c5350,c7182,c2216,c5286,c6137,c676,c1492,c6208,c2309,c6126,c6131,c16,c9225,c4368,c3335,c8462,c3343,c7240,c2204,c7377,c9164,c4263,c9188,c4294,c6267,c2332,c774,c90,c6451,c782,c1208,c7368,c026,c5392,c9194,c5120,c9174,c4351,c2105,c5161,c5405,c6306,c8435,c4457,c6404,c771,c8260,c9327,c2153,c2499,c6317,c532,c9328,c6107,c9309,c3375,c6252,c7255,c8228,c815,c059,c8365,c7419,c9349,c5449,c1114,c4209,c830,c5188,c1335,c5442,c116,c3393,c721,c3212,c4494,c60,c4128,c797,c5200,c349,c3454,c0113,c88,c7437,c1169,c5266,c1460,c069,c5242,c2119,c2258,c0393,c9399,c6254,c2160,c979,c3173,c7381,c481,c1145,c7190,c00,c0120,c8267,c3104,c446,c0363,c2307,c5110,c1473,c630,c0491,c3421,c7288,c2475,c0362,c6241,c0244,c240,c0147,c5108,c0245,c6223,c2377,c9199,c4381,c8124,c7429,c9361,c474,c4448,c5173,c5125,c2399,c1409,c468,c614,c262,c5486,c2249,c4409,c9481,c3351,c8299,c1407,c7128,c8472,c8369,c7149,c5190,c3211,c2314,c673,c2370,c0179,c7261,c714,c2428,c3110,c3266,c690,c1295,c596,c739,c3424,c1495,c0333,c7430,c612,c4224,c521,c3239,c7452,c5275,c4214,c5366,c2416,c1217,c8298,c0343,c178,c2127,c0452,c1163,c2478,c1375,c3443,c3402,c174,c572,c524,c3190,c9224,c3213,c634,c0104,c1125,c0458,c2424,c266,c4233,c790,c8364,c2269,c7163,c7164,c1393,c9304,c123,c2362,c1297,c577,c2347,c1341,c8391,c1164,c2229,c3354,c143,c999,c824,c752,c694,c8467,c076,c2308,c2327,c4140,c235,c2465,c7343,c5417,c1438,c7108,c6495,c8188,c6353,c7124,c9382,c0124,c4405,c2155,c665,c6293,c0187,c3301,c032,c8466,c2186,c692,c4118,c6332,c0390,c9339,c7440,c759,c591,c3415,c6478,c2261,c555,c961,c4308,c7121,c6140,c677,c6326,c374,c942,c5131,c982,c1150,c1257,c130,c559,c4471,c6499,c0453,c1113,c3320,c8347,c7353,c2391,c7456,c439,c613,c617,c3145,c567,c5496,c743,c6245,c0463,c3414,c4309,c6118,c122,c246,c4151,c7344,c3456,c151,c6412,c9421,c2118,c9263,c5418,c650,c6419,c3223,c6494,c754,c7392,c4249,c3484,c7161,c7145,c4178,c8170,c1420,c7391,c8412,c5365,c7196,c9385,c4133,c3380,c5221,c0206,c3357,c65,c828,c0479,c8471,c3199,c9259,c2210,c1177,c267,c7400,c2384,c0419,c0140,c5112,c8305,c8448,c6191,c2169,c861,c3364,c9470,c7291,c9496,c660,c1138,c6123,c1213,c1225,c6460,c2233,c4139,c9191,c012,c2462,c1293,c520,c2489,c321,c5142,c9337,c2277,c0428,c9181,c817,c4143,c8225,c6183,c2285,c9301,c2146,c2494,c8383,c550,c6283,c0319,c0295,c5354,c5466,c469,c318,c7349,c3129,c2433,c337,c2198,c2265,c5342,c6376,c8179,c8417,c1496,c4106,c9373,c1427,c0486,c7357,c8303,c429,c0407,c324,c7431,c5414,c7385,c8476,c2310,c4235,c1466,c380,c6447,c0314,c7371,c4307,c6272,c960,c3132,c3347,c6232,c2224,c9117,c9310,c820,c9367,c5368,c0399,c4433,c0252,c8385,c8301,c0323,c393,c9267,c3107,c3379,c8129,c7223,c3442,c420,c1343,c6433,c4262,c1250,c4378,c7222,c8149,c7220,c9334,c5180,c3358,c9321,c5206,c585,c7292,c3497,c196,c9420,c7296,c160,c1109,c395,c8229,c4129,c255,c623,c2250,c4111,c5467,c925,c4176,c6383,c0233,c0303,c4424,c742,c5213,c0331,c1247,c9366,c1421,c8379,c5447,c4146,c440,c7246,c7315,c5204,c1453,c364,c047,c6479,c397,c9407,c5482,c7103,c53,c295,c5127,c738,c7200,c050,c9374,c1299,c0197,c1497,c0296,c4281,c5410,c4218,c0222,c3121,c070,c8292,c4237,c8105,c9132,c910,c9172,c786,c411,c741,c8237,c2459,c6361,c7273,c4292,c7297,c7408,c7481,c6129,c9100,c281,c6497,c2263,c8214,c765,c1388,c4417,c9228,c137,c0304,c0205,c3399,c4244,c6455,c4193,c2420,c9329,c0487,c7335,c089,c536,c0388,c3101,c6171,c8372,c1481,c6110,c4173,c8297,c5428,c4350,c9209,c357,c6423,c0443,c81,c3345,c6248,c053,c8246,c3321,c8405,c989,c5390,c9322,c2422,c4289,c5261,c2256,c4167,c8381,c0291,c654,c3158,c4115,c4458,c56,c6454,c7435,c8458,c7397,c8422,c6357,c1259,c9452,c6352,c9279,c114,c4136,c449,c316,c0135,c4110,c6346,c368,c6275,c7118,c9139,c2311,c4242,c7215,c4185,c9341,c132,c6168,c6164,c855,c5308,c9324,c2350,c1352,c7109,c0255,c2190,c3489,c9232,c0225,c4239,c2426,c8100,c0330,c2456,c8226,c5113,c1311,c3270,c4431,c8240,c1195,c2230,c6370,c390,c6325,c152,c3494,c6441,c9184,c35,c9115,c6239,c0321,c647,c6299,c1166,c553,c0403,c0351,c4283,c0156,c0139,c7293,c6381,c1360,c1144,c7139,c3446,c6484,c8490,c1317,c2150,c9236,c3258,c5307,c278,c5348,c6443,c9494,c1171,c2154,c4125,c422,c168,c5423,c8232,c0477,c9121,c3176,c7330,c9365,c0381,c5140,c1478,c4236,c7239,c5236,c0455,c4243,c4204,c8403,c2205,c793,c845,c1413,c4498,c6347,c769,c0276,c03,c7311,c0226,c167,c4349,c4130,c2466,c3222,c4399,c8337,c750,c4467,c1236,c4463,c2365,c6219,c7136,c2364,c2215,c8335,c0418,c0496,c8101,c7270,c930,c730,c8323,c2241,c0284,c6235,c344,c2227,c0173,c1127,c9167,c8221,c2373,c7480,c4311,c213,c4428,c2460,c4290,c1249,c3455,c1498,c5363,c3182,c3124,c3483,c9458,c0122,c1187,c7126,c9377,c3174,c5427,c687,c9454,c4221,c946,c1400,c1397,c2346,c5364,c2398,c5231,c7129,c3259,c0185,c8444,c844,c6329,c5478,c484,c099,c9265,c8492,c371,c4439,c6100,c2245,c4354,c054,c9317,c718,c2454,c7245,c8133,c1372,c2442,c9112,c497,c9444,c5316,c980,c9177,c6348,c0204,c4385,c5212,c6156,c7195,c6304,c4486,c8171,c8115,c4432,c7317,c9241,c5346,c0267,c492,c1389,c0378,c9459,c4429,c7411,c1161,c6139,c0105,c1251,c8384,c8429,c94,c5160,c3453,c818,c2319,c4323,c927,c7307,c5349,c166,c0414,c2304,c9240,c2121,c6173,c9315,c3306,c1353,c4197,c282,c9150,c3383,c0166,c6277,c1263,c3264,c1231,c0311,c0196,c2266,c3405,c7214,c991,c3287,c5184,c3392,c9248,c4196,c9468,c0361,c0126,c3127,c0141,c5495,c9298,c1378,c632,c7192,c1261,c9253,c9408,c2111,c5437,c949,c7360,c247,c0373,c6377,c9493,c887,c9233,c962,c568,c0438,c2248,c9124,c4377,c0273,c8238,c719,c0114,c1361,c8211,c3281,c1107,c778,c6437,c3328,c1143,c624,c5338,c0483,c1206,c04,c7367,c3171,c7249,c582,c9140,c3391,c4343,c767,c3232,c2125,c939,c2145,c1402,c2326,c9251,c725,c952,c2480,c7138,c8351,c0137,c0271,c445,c230,c314,c0324,c7135,c6220,c635,c3116,c4158,c4443,c3284,c8419,c083,c1398,c5326,c9405,c8243,c9219,c8375,c9395,c744,c396,c651,c0309,c1455,c1122,c0405,c2243,c389,c5432,c8310,c2120,c6242,c332,c9235,c5228,c9179,c8284,c6279,c3175,c6198,c9119,c8332,c69,c3115,c323,c5244,c0354,c1271,c2405,c897,c5416,c997,c7243,c7468,c9340,c3204,c1246,c670,c6102,c326,c9446,c3378,c4328,c186,c5298,c527,c9355,c2446,c573,c0437,c9134,c1180,c8287,c9166,c4358,c4123,c956,c1117,c2262,c8140,c4329,c5185,c5214,c8253,c3477,c0467,c4436,c896,c8404,c6393,c2268,c2435,c0379,c515,c5313,c6128,c513,c736,c3462,c4268,c6379,c491,c7345,c6237,c519,c78,c6349,c7378,c0462,c1183,c584,c4172,c4177,c2313,c3112,c642,c8136,c85,c6449,c2130,c4166,c5170,c7386,c1318,c890,c667,c8244,c1128,c141,c2174,c3495,c6266,c3267,c6368,c028,c5202,c6461,c992,c3432,c77,c7341,c3350,c6295,c7361,c3193,c7460,c461,c2112,c3370,c5280,c0177,c6338,c388,c3481,c0200,c2439,c4357,c6413,c4223,c014,c352,c6384,c8130,c1290,c2113,c1394,c0317,c959,c07,c039,c9379,c4254,c5436,c2485,c2344,c9143,c6394,c988,c8156,c9449,c1468,c2110,c8207,c610,c0410,c6327,c7252,c5162,c3418,c39,c770,c7113,c62,c8327,c847,c4326,c7306,c0101,c766,c1493,c6233,c8498,c0332,c9151,c1146,c6101,c0315,c8163,c0201,c8165,c9221,c6440,c1108,c3325,c762,c7210,c4496,c4296,c3369,c0429,c4389,c226,c7275,c1412,c881,c61,c9331,c2179,c5166,c0110,c040,c2417,c5303,c5443,c862,c1227,c1494,c757,c5153,c2188,c2231,c6113,c92,c2197,c8223,c937,c161,c2192,c5192,c2240,c8437,c2474,c9448,c2226,c2390,c2491,c8183,c3373,c4427,c342,c7451,c2292,c020,c7338,c9489,c6217,c7415,c1415,c2176,c7276,c9266,c327,c3295,c7224,c274,c441,c4202,c0150,c8331,c6418,c1126,c8141,c0153,c056,c0169,c2161,c3459,c3488,c9497,c6285,c7347,c3146,c2132,c5490,c2290,c9270,c3387,c2279,c7173,c0262,c8454,c0356,c751,c8290,c7486,c8418,c7478,c5285,c8485,c3311,c3319,c5463,c934,c1192,c2140,c5216,c8317,c3388,c6312,c5415,c4282,c9203,c7323,c9495,c1483,c9438,c8274,c9425,c044,c3316,c525,c7498,c5422,c6260,c276,c8247,c1387,c416,c551,c9293,c5409,c787,c7181,c3332,c425,c8450,c3224,c5281,c4488,c1214,c675,c9435,c9487,c8230,c1175,c2109,c423,c6316,c4461,c0394,c5253,c885,c546,c7446,c6180,c8496,c8377,c0281,c884,c2189,c1216,c1159,c0251,c5421,c5351,c5223,c7418,c8306,c713,c2302,c3466,c9281,c7492,c1140,c7466,c3496,c4481,c674,c7141,c1160,c8318,c6103,c4421,c3185,c3384,c4288,c2208,c932,c0210,c812,c9123,c6280,c0224,c966,c4131,c5224,c7238,c391,c5193,c834,c311,c0402,c6243,c0344,c0454,c7458,c365,c7417,c1253,c746,c916,c2436,c2148,c5375,c9288,c7157,c260,c530,c6182,c620,c197,c2213,c8363,c3416,c8464,c7403,c6314,c8161,c912,c3285,c3470,c2128,c5396,c8463,c6367,c1331,c8459,c0151,c99,c1165,c9434,c7295,c4231,c6363,c3216,c7107,c8320,c7134,c0481,c8120,c733,c3156,c7219,c6320,c8296,c1358,c662,c5480,c6135,c8151,c1170,c2336,c7247,c8173,c4208,c7168,c024,c511,c8209,c9109,c545,c3434,c1269,c7180,c3170,c1439,c0451,c8212,c3142,c6477,c0366,c6230,c727,c7374,c2486,c4480,c2296,c4372,c9173,c0243,c4164,c1327,c1115,c7201,c841,c6444,c7286,c3163,c125,c2257,c7179,c590,c4330,c9387,c0411,c5174,c1354,c4253,c955,c2440,c3219,c0214,c5107,c0203,c046,c6313,c8262,c5372,c0325,c9372,c2166,c2177,c7443,c933,c7355,c0358,c0193,c1436,c9289,c0374,c426,c8389,c3293,c4293,c5100,c574,c5407,c4485,c0265,c8258,c6309,c8314,c0431,c5397,c8397,c3177,c679,c1282,c0145,c8387,c8252,c0492,c0318,c9107,c9307,c8482,c2199,c2447,c2320,c1191,c2468,c6115,c3159,c8218,c4335,c4191,c9187,c9245,c4444,c385,c6350,c9131,c7150,c6496,c9256,c5148,c2318,c3329,c5497,c5270,c3111,c6446,c1431,c3202,c4412,c795,c737,c71,c7142,c0306,c3346,c485,c6333,c543,c4487,c6355,c72,c9175,c7244,c7101,c5385,c2144,c9491,c348,c7277,c5154,c5195,c9299,c1200,c557,c5487,c7203,c6206,c9223,c3227,c2219,c4327,c578,c121,c6397,c7303,c4265,c015,c2172,c6386,c4260,c1417,c2431,c8353,c8333,c2467,c1482,c3123,c0484,c7301,c2393,c6194,c3118,c628,c1338,c24,c8157,c4319,c7178,c4321,c8455,c889,c6224,c899,c1244,c6127,c693,c724,c9214,c3397,c6124,c0242,c3114,c6253,c682,c0383,c3179,c5234,c3152,c4497,c5357,c6286,c216,c664,c055,c943,c1324,c5300,c7326,c6448,c9485,c6287,c8147,c5114,c575,c4199,c684,c7336,c8106,c1411,c983,c2473,c552,c1149,c071,c480,c8436,c418,c5119,c953,c1474,c7485,c6422,c5453,c1359,c954,c098,c7366,c2142,c7167,c334,c496,c6185,c7380,c8185,c9127,c0132,c0494,c0274,c135,c1489,c4279,c02,c0236,c564,c4179,c0172,c0142,c3465,c3149,c8264,c7497,c1396,c3365,c5134,c0111,c5470,c9204,c73,c5360,c296,c8313,c4313,c836,c129,c7352,c335,c6229,c888,c5445,c858,c1104,c6473,c794,c261,c7382,c5186,c5155,c220,c1267,c291,c0240,c6249,c2200,c8366,c852,c6457,c6380,c781,c4367,c273,c1196,c5272,c571,c3296,c3400,c0384,c3168,c6247,c0100,c4132,c8340,c4423,c4338,c6472,c150,c7423,c6493,c554,c8358,c7469,c9190,c9409,c087,c5106,c569,c646,c4274,c8341,c7383,c110,c4489,c3102,c994,c7491,c9302,c3236,c1174,c0231,c0347,c9356,c0130,c2458,c4425,c6450,c9480,c1384,c0387,c7474,c1315,c9268,c0430,c4304,c3205,c224,c5462,c475,c232,c55,c666,c8362,c5265,c6209,c6385,c97,c0456,c7390,c3165,c3396,c6244,c0161,c4422,c539,c2225,c619,c2371,c2223,c5215,c3210,c4226,c1348,c430,c4394,c9476,c971,c3361,c8206,c1168,c6268,c5296,c3491,c7302,c5430,c2322,c560,c0190,c2159,c287,c3448,c3367,c011,c1220,c0175,c0170,c5230,c696,c2331,c8456,c3186,c0441,c535,c6172,c0307,c918,c292,c8241,c8148,c330,c2143,c4101,c1198,c9398,c4160,c1357,c5460,c147,c6467,c8487,c8478,c6109,c1401,c8250,c5240,c9400,c848,c9353,c6466,c40,c2187,c1262,c6199,c5128,c0310,c5334,c6174,c4114,c7475,c4353,c6184,c7146,c7455,c3120,c5301,c376,c7472,c3180,c9338,c4220,c3349,c5143,c5419,c8348,c3498,c747,c3151,c284,c7364,c236,c7379,c698,c859,c5201,c779,c7148,c2329,c9290,c7409,c2410,c5295,c8411,c0345,c9159,c4342,c3360,c8162,c1283,c9335,c0469,c663,c6257,c2104,c8445,c6296,c6203,c7362,c926,c8123,c9473,c1286,c878,c1254,c5145,c8449,c3404,c785,c5205,c5426,c6112,c82,c777,c7125,c030,c1432,c8281,c9345,c4391,c0433,c120,c9433,c1292,c9138,c5345,c5220,c3265,c6300,c7151,c1294,c8200,c6255,c1477,c4162,c1162,c8278,c8370,c720,c1355,c0217,c1435,c4194,c8194,c3294,c8160,c2389,c645,c9243,c533,c251,c7274,c4317,c0118,c0219,c3122,c4479,c5439,c8309,c5461,c5163,c435,c680,c2228,c3188,c2352,c6490,c8461,c9343,c7199,c996,c2400,c756,c241,c8277,c466,c4259,c085,c8134,c8164,c8378,c1383,c9254,c265,c6177,c0420,c6482,c86,c2238,c9246,c5133,c760,c7198,c2147,c14,c51,c0278,c977,c13,c142,c5399,c9285,c095,c4188,c0257,c87,c0290,c9213,c9439,c9428,c2157,c0329,c3226,c6391,c7434,c312,c3451,c2429,c2330,c5252,c8390,c3374,c7298,c723,c710,c2427,c7445,c1342,c1463,c1157,c629,c1447,c2236,c4276,c3412,c7473,c8322,c1194,c3229,c8271,c8205,c6458,c6298,c978,c3308,c8308,c7197,c1202,c1193,c7290,c0279,c1326,c3291,c4201,c7175,c1446,c128,c5324,c188,c783,c3352,c1488,c631,c9369,c1452,c7471,c5413,c1369,c1245,c156,c950,c153,c36,c875,c7127,c1300,c6442,c4301,c6372,c0372,c7170,c7144,c3355,c0249,c5210,c8468,c7304,c1370,c598,c2345,c5412,c9410,c3377,c4462,c1433,c350,c8376,c2237,c0474,c5335,c2437,c5250,c242,c0109,c9238,c6261,c5343,c0212,c1426,c1405,c7177,c8427,c264,c375,c2457,c4419,c6270,c0115,c8451,c2477,c6392,c7263,c2479,c6498,c6345,c4153,c5171,c1256,c2385,c387,c0260,c5151,c7358,c9415,c9319,c1312,c1203,c4370,c7487,c2114,c0181,c7206,c072,c0125,c0192,c880,c57,c6250,c361,c171,c1472,c7388,c3318,c7211,c9312,c4477,c472,c5329,c753,c4159,c0227,c7426,c1197,c2283,c8491,c6334,c8396,c5306,c5222,c8192,c3493,c9347,c7267,c424,c7241,c5386,c356,c7410,c30,c9457,c23,c9202,c4303,c8128,c0149,c7395,c1450,c5194,c4138,c2423,c3292,c1490,c975,c6421,c0349,c1215,c4266,c6311,c5402,c6452,c3394,c7123,c7359,c412,c3382,c8367,c6453,c4186,c5197,c6439,c761,c3209,c5455,c5294,c290,c259,c7488,c2298,c2407,c3419,c0448,c163,c915,c7188,c018,c417,c4275,c3452,c394,c6212,c1280,c0213,c0355,c074,c776,c7189,c2122,c681,c6204,c5187,c648,c9142,c3136,c9120,c1406,c7162,c3438,c2406,c5393,c4165,c2165,c1106,c119,c9389,c229,c5115,c9286,c0380,c9165,c8138,c2259,c4222,c5314,c6456,c5472,c5255,c3303,c3359,c3395,c2323,c5124,c1444,c4482,c1385,c1155,c2441,c5302,c842,c021,c6387,c372,c3215,c3472,c748,c7279,c9295,c9396,c7130,c9261,c9226,c1228,c7398,c442,c633,c48,c688,c2409,c8172,c2239,c4440,c6489,c1137,c2376,c1306,c9460,c9205,c8356,c1134,c5424,c2312,c3261,c3429,c029,c3130,c0143,c3450,c3401,c987,c2115,c658,c8217,c4392,c9284,c4261,c7204,c9186,c792,c9200,c2378,c383,c599,c3441,c2425,c294,c3147,c0308,c041,c8121,c4318,c077,c544,c4108,c486,c7172,c63,c7496,c8118,c6382,c7294,c1142,c9330,c346,c5380,c7169,c243,c1309,c8150,c3268,c7329,c1279,c2152,c3437,c1476,c3305,c5403,c319,c5245,c1428,c6153,c5219,c2244,c921,c7396,c58,c6426,c1130,c3252,c6207,c112,c6471,c8102,c5293,c3422,c1211,c457,c0293,c2173,c6483,c9269,c0154,c1308,c2413,c465,c8282,c895,c6166,c6205,c831,c5475,c7420,c4352,c7462,c7268,c7187,c7225,c8346,c0416,c5251,c3148,c4420,c1268,c957,c1298,c1346,c035,c0288,c2412,c3426,c1382,c7155,c9445,c2334,c490,c5118,c9411,c763,c431,c968,c9278,c1265,c864,c4117,c6434,c9471,c4369,c0269,c0198,c338,c419,c067,c2117,c0398,c3253,c6297,c289,c2455,c5168,c0119,c2351,c2234,c2201,c9388,c460,c944,c8469,c1344,c8414,c2382,c1471,c3480,c5132,c3286,c3172,c9185,c113,c1289,c8307,c9125,c5257,c3463,c3269,c5406,c3262,c9227,c2275,c6417,c8430,c7363,c117,c6150,c9180,c3409,c0134,c172,c073,c3435,c2449,c1425,c2193,c0128,c1116,c1135,c1184,c4250,c8219,c4393,c1371,c872,c7165,c9303,c470,c381,c1484,c6167,c3126,c0228,c5318,c8181,c7207,c8393,c0189,c8155,c1399,c2108,c8400,c9234,c7389,c9418,c427,c4473,c839,c4109,c47,c516,c74,c2325,c2134,c5440,c6465,c9323,c4445,c7183,c5358,c7217,c7122,c6354,c4468,c1226,c0313,c668,c6234,c9229,c652,c5499,c0176,c212,c4232,c8434,c5152,c9249,c7102,c0328,c4107,c7251,c9474,c3372,c6425,c9297,c4230,c7354,c9275,c8432,c1224,c479,c5471,c9128,c5103,c5158,c936,c4298,c5156,c4297,c3240,c2116,c7324,c4414,c857,c7284,c31,c0138,c8168,c1181,c9456,c8470,c8202,c8158,c6200,c3178,c3220,c7394,c4207,c2450,c5433,c5147,c2273,c639,c2490,c211,c6114,c9351,c19,c4320,c8392,c7477,c0268,c428,c1404,c269,c9212,c1212,c1274,c5479,c0229,c315,c963,c9393,c0285,c93,c2297,c9193,c4456,c5381,c313,c6339,c1424,c2203,c0155,c7404,c2392,c1147,c7234,c8254,c1154,c328,c9258,c4182,c8176,c458,c6221,c2247,c8497,c3460,c9264,c3485,c4241,c4295,c5279,c4103,c5450,c068,c084,c5203,c9455,c272,c8184,c6148,c7120,c4460,c9152,c3166,c3487,c051,c9255,c4374,c7112,c52,c8394,c7308,c7457,c837,c6282,c3140,c223,c5320,c2360,c5136,c0280,c7399,c1367,c2432,c351,c1275,c2232,c144,c9189,c5389,c8388,c0460,c6228,c8178,c7432,c976,c3304,c9436,c9296,c148,c0400,c9390,c343,c2139,c4100,c984,c4491,c76,c1316,c5341,c353,c9262,c9153,c8196,c2434,c6402,c644,c5235,c2253,c3157,c715,c5456,c3191,c5448,c7132,c3336,c6436,c2496,c919,c3162,c6491,c1368,c2184,c1351,c6430,c0220,c131,c0401,c4442,c625,c9357,c0446,c250,c0376,c231,c4371,c249,c228,c8245,c9282,c580,c9451,c4384,c3187,c940,c3458,c8236,c7159,c5347,c5191,c149,c6469,c5111,c3430,c4438,c194,c0392,c967,c5483,c0103,c5139,c5373,c3242,c68,c0493,c6291,c5458,c9479,c6415,c583,c9475,c5325,c5452,c3249,c279,c0461,c097,c540,c1129,c538,c726,c3103,c3323,c7229,c1458,c851,c9208,c9383,c0359,c941,c9394,c5175,c096,c3221,c016,c4334,c6116,c126,c3274,c1322,c712,c2141,c6130,c175,c0464,c7470,c5489,c0158,c4415,c1255,c0480,c157,c8325,c4154,c222,c4388,c5387,c3363,c7444,c22,c9391,c4195,c3340,c3277,c5189,c9305,c0312,c0112,c8409,c7250,c8380,c8275,c4344,c874,c0389,c7264,c8428,c8272,c8255,c0270,c3482,c2403,c6485,c5299,c4418,c2414,c3247,c0286,c3106,c065,c3256,c8126,c2348,c0182,c9272,c8319,c6263,c8355,c3337,c1237,c512,c4316,c5283,c2353,c7375,c8399,c7205,c9103,c0215,c8256,c354,c9499,c1186,c286,c7115,c9146,c5198,c2124,c2394,c8145,c0432,c3181,c2287,c3407,c0485,c1204,c3417,c5199,c7340,c4149,c6231,c938,c6202,c7253,c3134,c9466,c922,c768,c8197,c4410,c0478,c5182,c0468,c1304,c7104,c6358,c6281,c0183,c4277,c9149,c592,c2123,c7283,c9141,c4483,c8265,c5123,c34,c6464,c9195,c9176,c2321,c0475,c84,c0300,c6186,c3150,c7489,c7450,c9486,c764,c1273,c199,c8407,c9325,c868,c3206,c3203,c7356,c2445,c9348,c9133,c1112,c5225,c8406,c695,c8401,c0377,c277,c3167,c3225,c8345,c6403,c6175,c8286,c2171,c1172,c0180,c6188,c8360,c722,c0422,c2138,c9292,c7372,c6236,c638,c4169,c5438,c6214,c1422,c0305,c8479,c6264,c4269,c0275,c1233,c359,c3237,c4291,c1219,c6292,c6213,c0472,c01,c6324,c0294,c4331,c5288,c811,c092,c4267,c732,c1486,c5441,c5444,c856,c0368,c3362,c4170,c3133,c2272,c7350,c1307,c8111,c8359,c9376,c5420,c810,c717,c7424,c4284,c254,c7346,c4345,c5126,c7258,c877,c1209,c2133,c421,c1465,c4406,c057,c081,c0247,c1440,c2251,c9397,c5277,c4278,c4145,c9239,c2438,c4446,c6155,c6160,c9354,c0350,c5362,c6178,c8420,c6470,c7242,c253,c826,c079,c179,c6269,c6378,c5232,c1156,c6315,c7202,c42,c3108,c8334,c3313,c4192,c3324,c8224,c0289,c5227,c5218,c8465,c9488,c7191,c182,c5468,c0371,c6289,c7370,c5249,c498,c2106,c7461,c8231,c8421,c998,c3251,c1457,c2343,c3431,c1133,c947,c7321,c4333,c4287,c5254,c1238,c5315,c3403,c1305,c510,c791,c310,c9161,c8300,c9380,c7428,c9247,c8321,c234,c0439,c869,c8329,c5260,c8208,c9490,c476,c6330,c7111,c2137,c4476,c4465,c3398,c4124,c3342,c5289,c2100,c1376,c9198,c325,c9326,c2196,c1323,c9207,c6480,c0499,c1242,c5337,c4102,c7176,c2372,c6226,c5355,c7312,c1434,c7256,c6125,c4189,c541,c3235,c9320,c333,c566,c8408,c340,c576,c5319,c4273,c1302,c70,c2483,c4187,c2317,c4322,c993,c4310,c0211,c12,c078,c373,c0162,c0335,c9178,c245,c11,c5459,c8139,c3245,c483,c9169,c7174,c0159,c2280,c377,c3327,c0436,c846,c5332,c6121,c3410,c1391,c8350,c0386,c3331,c7281,c595,c9404,c9461,c4346,c6246,c8175,c8251,c6225,c0248,c6161,c0292,c2212,c7117,c4452,c2354,c4216,c7412,c8302,c98,c6201,c8233,c740,c894,c2488,c825,c263,c8266,c5177,c4398,c964,c9450,c7140,c5150,c3307,c8413,c2260,c4285,c0239,c2136,c036,c9183,c0421,c2220,c5323,c8499,c935,c0164,c4495,c871,c0470,c1332,c8473,c7436,c3244,c4314,c210,c1167,c843,c136,c0417,c233,c2180,c1291,c1429,c6240,c929,c4148,c8443,c1479,c4183,c133,c8143,c0146,c410,c299,c8268,c1240,c4430,c7158,c1243,c283,c931,c8431,c4332,c4286,c5464,c6474,c4404,c9453,c59,c0367,c219,c2359,c972,c1111,c9422,c450,c4493,c689,c1207,c4395,c9401,c6488,c0258,c784,c2324,c7133,c4472,c6336,c2411,c1320,c4251,c4312,c0160,c0404,c413,c049,c5310,c7309,c2281,c9342,c0449,c7407,c2254,c5102,c9116,c459,c3312,c5164,c534,c8137,c8220,c973,c3135,c8263,c8294,c8423,c2448,c4142,c37,c363,c0339,c0426,c616,c2487,c6216,c2278,c1222,c5431,c731,c1380,c0327,c2131,c8488,c189,c8295,c2270,c2252,c2284,c1123,c1475,c280,c320,c838,c9211,c094,c1456,c586,c2451,c2453,c2495,c50,c2363,c7393,c3473,c8438,c6492,c8108,c8433,c813,c7114,c118,c8127,c5246,c6318,c3278,c8291,c6331,c7152,c6122,c033,c1470,c2246,c4229,c528,c0498,c526,c5267,c8415,c8187,c4134,c8186,c8177,c2178,c2335,c4264,c9231,c8339,c965,c4306,c5287,c5259,c3137,c6215,c518,c7447,c268,c3138,c293,c1118,c4161,c8153,c6193,c6162,c9360,c1235,c5491,c4112,c7495,c5104,c5165,c08,c1333,c4325,c0457,c7314,c0218,c477,c6435,c7416,c010,c2126,c749,c9447,c5400,c4252,c048,c0409,c434,c7348,c1148,c6106,c7427,c821,c2183,c176,c6170,c7401 );

input x0;
input x1;
input x2;
input x3;
input x4;
input x5;
input x6;
input x7;
input x8;
input x9;
input x10;
input x11;
input x12;
input x13;
input x14;
input x15;
input x16;
input x17;
input x18;
input x19;
input x20;
input x21;
input x22;
input x23;
input x24;
input x25;
input x26;
input x27;
input x28;
input x29;
input x30;
input x31;
input x32;
input x33;
input x34;
input x35;
input x36;
input x37;
input x38;
input x39;
input x40;
input x41;
input x42;
input x43;
input x44;
input x45;
input x46;
input x47;
input x48;
input x49;
input x50;
input x51;
input x52;
input x53;
input x54;
input x55;
input x56;
input x57;
input x58;
input x59;
input x60;
input x61;
input x62;
input x63;
input x64;
input x65;
input x66;
input x67;
input x68;
input x69;
input x70;
input x71;
input x72;
input x73;
input x74;
input x75;
input x76;
input x77;
input x78;
input x79;
input x80;
input x81;
input x82;
input x83;
input x84;
input x85;
input x86;
input x87;
input x88;
input x89;
input x90;
input x91;
input x92;
input x93;
input x94;
input x95;
input x96;
input x97;
input x98;
input x99;
input x100;
input x101;
input x102;
input x103;
input x104;
input x105;
input x106;
input x107;
input x108;
input x109;
input x110;
input x111;
input x112;
input x113;
input x114;
input x115;
input x116;
input x117;
input x118;
input x119;
input x120;
input x121;
input x122;
input x123;
input x124;
input x125;
input x126;
input x127;
input x128;
input x129;
input x130;
input x131;
input x132;
input x133;
input x134;
input x135;
input x136;
input x137;
input x138;
input x139;
input x140;
input x141;
input x142;
input x143;
input x144;
input x145;
input x146;
input x147;
input x148;
input x149;
input x150;
input x151;
input x152;
input x153;
input x154;
input x155;
input x156;
input x157;
input x158;
input x159;
input x160;
input x161;
input x162;
input x163;
input x164;
input x165;
input x166;
input x167;
input x168;
input x169;
input x170;
input x171;
input x172;
input x173;
input x174;
input x175;
input x176;
input x177;
input x178;
input x179;
input x180;
input x181;
input x182;
input x183;
input x184;
input x185;
input x186;
input x187;
input x188;
input x189;
input x190;
input x191;
input x192;
input x193;
input x194;
input x195;
input x196;
input x197;
input x198;
input x199;
input x200;
input x201;
input x202;
input x203;
input x204;
input x205;
input x206;
input x207;
input x208;
input x209;
input x210;
input x211;
input x212;
input x213;
input x214;
input x215;
input x216;
input x217;
input x218;
input x219;
input x220;
input x221;
input x222;
input x223;
input x224;
input x225;
input x226;
input x227;
input x228;
input x229;
input x230;
input x231;
input x232;
input x233;
input x234;
input x235;
input x236;
input x237;
input x238;
input x239;
input x240;
input x241;
input x242;
input x243;
input x244;
input x245;
input x246;
input x247;
input x248;
input x249;
input x250;
input x251;
input x252;
input x253;
input x254;
input x255;
input x256;
input x257;
input x258;
input x259;
input x260;
input x261;
input x262;
input x263;
input x264;
input x265;
input x266;
input x267;
input x268;
input x269;
input x270;
input x271;
input x272;
input x273;
input x274;
input x275;
input x276;
input x277;
input x278;
input x279;
input x280;
input x281;
input x282;
input x283;
input x284;
input x285;
input x286;
input x287;
input x288;
input x289;
input x290;
input x291;
input x292;
input x293;
input x294;
input x295;
input x296;
input x297;
input x298;
input x299;
input x300;
input x301;
input x302;
input x303;
input x304;
input x305;
input x306;
input x307;
input x308;
input x309;
input x310;
input x311;
input x312;
input x313;
input x314;
input x315;
input x316;
input x317;
input x318;
input x319;
input x320;
input x321;
input x322;
input x323;
input x324;
input x325;
input x326;
input x327;
input x328;
input x329;
input x330;
input x331;
input x332;
input x333;
input x334;
input x335;
input x336;
input x337;
input x338;
input x339;
input x340;
input x341;
input x342;
input x343;
input x344;
input x345;
input x346;
input x347;
input x348;
input x349;
input x350;
input x351;
input x352;
input x353;
input x354;
input x355;
input x356;
input x357;
input x358;
input x359;
input x360;
input x361;
input x362;
input x363;
input x364;
input x365;
input x366;
input x367;
input x368;
input x369;
input x370;
input x371;
input x372;
input x373;
input x374;
input x375;
input x376;
input x377;
input x378;
input x379;
input x380;
input x381;
input x382;
input x383;
input x384;
input x385;
input x386;
input x387;
input x388;
input x389;
input x390;
input x391;
input x392;
input x393;
input x394;
input x395;
input x396;
input x397;
input x398;
input x399;
input x400;
input x401;
input x402;
input x403;
input x404;
input x405;
input x406;
input x407;
input x408;
input x409;
input x410;
input x411;
input x412;
input x413;
input x414;
input x415;
input x416;
input x417;
input x418;
input x419;
input x420;
input x421;
input x422;
input x423;
input x424;
input x425;
input x426;
input x427;
input x428;
input x429;
input x430;
input x431;
input x432;
input x433;
input x434;
input x435;
input x436;
input x437;
input x438;
input x439;
input x440;
input x441;
input x442;
input x443;
input x444;
input x445;
input x446;
input x447;
input x448;
input x449;
input x450;
input x451;
input x452;
input x453;
input x454;
input x455;
input x456;
input x457;
input x458;
input x459;
input x460;
input x461;
input x462;
input x463;
input x464;
input x465;
input x466;
input x467;
input x468;
input x469;
input x470;
input x471;
input x472;
input x473;
input x474;
input x475;
input x476;
input x477;
input x478;
input x479;
input x480;
input x481;
input x482;
input x483;
input x484;
input x485;
input x486;
input x487;
input x488;
input x489;
input x490;
input x491;
input x492;
input x493;
input x494;
input x495;
input x496;
input x497;
input x498;
input x499;
input x500;
input x501;
input x502;
input x503;
input x504;
input x505;
input x506;
input x507;
input x508;
input x509;
input x510;
input x511;
input x512;
input x513;
input x514;
input x515;
input x516;
input x517;
input x518;
input x519;
input x520;
input x521;
input x522;
input x523;
input x524;
input x525;
input x526;
input x527;
input x528;
input x529;
input x530;
input x531;
input x532;
input x533;
input x534;
input x535;
input x536;
input x537;
input x538;
input x539;
input x540;
input x541;
input x542;
input x543;
input x544;
input x545;
input x546;
input x547;
input x548;
input x549;
input x550;
input x551;
input x552;
input x553;
input x554;
input x555;
input x556;
input x557;
input x558;
input x559;
input x560;
input x561;
input x562;
input x563;
input x564;
input x565;
input x566;
input x567;
input x568;
input x569;
input x570;
input x571;
input x572;
input x573;
input x574;
input x575;
input x576;
input x577;
input x578;
input x579;
input x580;
input x581;
input x582;
input x583;
input x584;
input x585;
input x586;
input x587;
input x588;
input x589;
input x590;
input x591;
input x592;
input x593;
input x594;
input x595;
input x596;
input x597;
input x598;
input x599;
input x600;
input x601;
input x602;
input x603;
input x604;
input x605;
input x606;
input x607;
input x608;
input x609;
input x610;
input x611;
input x612;
input x613;
input x614;
input x615;
input x616;
input x617;
input x618;
input x619;
input x620;
input x621;
input x622;
input x623;
input x624;
input x625;
input x626;
input x627;
input x628;
input x629;
input x630;
input x631;
input x632;
input x633;
input x634;
input x635;
input x636;
input x637;
input x638;
input x639;
input x640;
input x641;
input x642;
input x643;
input x644;
input x645;
input x646;
input x647;
input x648;
input x649;
input x650;
input x651;
input x652;
input x653;
input x654;
input x655;
input x656;
input x657;
input x658;
input x659;
input x660;
input x661;
input x662;
input x663;
input x664;
input x665;
input x666;
input x667;
input x668;
input x669;
input x670;
input x671;
input x672;
input x673;
input x674;
input x675;
input x676;
input x677;
input x678;
input x679;
input x680;
input x681;
input x682;
input x683;
input x684;
input x685;
input x686;
input x687;
input x688;
input x689;
input x690;
input x691;
input x692;
input x693;
input x694;
input x695;
input x696;
input x697;
input x698;
input x699;
input x700;
input x701;
input x702;
input x703;
input x704;
input x705;
input x706;
input x707;
input x708;
input x709;
input x710;
input x711;
input x712;
input x713;
input x714;
input x715;
input x716;
input x717;
input x718;
input x719;
input x720;
input x721;
input x722;
input x723;
input x724;
input x725;
input x726;
input x727;
input x728;
input x729;
input x730;
input x731;
input x732;
input x733;
input x734;
input x735;
input x736;
input x737;
input x738;
input x739;
input x740;
input x741;
input x742;
input x743;
input x744;
input x745;
input x746;
input x747;
input x748;
input x749;
input x750;
input x751;
input x752;
input x753;
input x754;
input x755;
input x756;
input x757;
input x758;
input x759;
input x760;
input x761;
input x762;
input x763;
input x764;
input x765;
input x766;
input x767;
input x768;
input x769;
input x770;
input x771;
input x772;
input x773;
input x774;
input x775;
input x776;
input x777;
input x778;
input x779;
input x780;
input x781;
input x782;
input x783;
output c589;
output c358;
output c9206;
output c9145;
output c0266;
output c4450;
output c4198;
output c866;
output c238;
output c4366;
output c46;
output c4200;
output c4245;
output c2300;
output c3445;
output c853;
output c1158;
output c8460;
output c6341;
output c8426;
output c1136;
output c8154;
output c6181;
output c4255;
output c7131;
output c2379;
output c6176;
output c5374;
output c4234;
output c5105;
output c8371;
output c556;
output c6487;
output c9484;
output c013;
output c6146;
output c4168;
output c1223;
output c1188;
output c6142;
output c1103;
output c8326;
output c7248;
output c4437;
output c8354;
output c0395;
output c436;
output c3197;
output c4364;
output c6104;
output c2369;
output c6359;
output c3356;
output c5328;
output c0263;
output c1201;
output c4120;
output c5144;
output c9406;
output c9148;
output c060;
output c6351;
output c444;
output c8373;
output c1347;
output c7318;
output c0427;
output c1408;
output c4339;
output c322;
output c3119;
output c170;
output c1303;
output c7147;
output c8374;
output c5122;
output c3241;
output c366;
output c5248;
output c3420;
output c9414;
output c8477;
output c7490;
output c3255;
output c522;
output c8203;
output c8257;
output c464;
output c1340;
output c735;
output c257;
output c8343;
output c5241;
output c3310;
output c4227;
output c6238;
output c917;
output c9370;
output c9472;
output c7339;
output c1395;
output c7259;
output c193;
output c382;
output c4337;
output c3279;
output c154;
output c3144;
output c3386;
output c4203;
output c4469;
output c656;
output c4386;
output c9162;
output c9386;
output c7185;
output c7300;
output c1239;
output c7260;
output c8107;
output c6321;
output c4359;
output c467;
output c05;
output c3299;
output c1266;
output c6375;
output c5138;
output c0216;
output c8166;
output c2295;
output c7448;
output c7310;
output c3428;
output c558;
output c5312;
output c1454;
output c7342;
output c9300;
output c138;
output c6133;
output c9280;
output c2135;
output c985;
output c198;
output c4361;
output c3315;
output c5239;
output c1229;
output c8486;
output c3271;
output c21;
output c6335;
output c4135;
output c4340;
output c6305;
output c1345;
output c2340;
output c3160;
output c2107;
output c7438;
output c9363;
output c3141;
output c3475;
output c1321;
output c2333;
output c945;
output c1270;
output c5311;
output c7221;
output c1221;
output c3457;
output c6271;
output c8199;
output c8481;
output c0259;
output c0445;
output c4147;
output c7333;
output c8234;
output c958;
output c2471;
output c3125;
output c2271;
output c7236;
output c3341;
output c1182;
output c5378;
output c1278;
output c2472;
output c6132;
output c1189;
output c139;
output c1210;
output c9368;
output c0375;
output c225;
output c1152;
output c9102;
output c26;
output c4451;
output c5371;
output c8182;
output c3198;
output c8494;
output c3246;
output c9244;
output c062;
output c4257;
output c7328;
output c159;
output c4300;
output c5207;
output c2294;
output c4122;
output c9413;
output c6371;
output c0223;
output c7369;
output c1373;
output c3196;
output c758;
output c0440;
output c454;
output c9242;
output c6463;
output c3109;
output c2397;
output c9197;
output c4299;
output c2415;
output c734;
output c1234;
output c9402;
output c5247;
output c6431;
output c18;
output c1301;
output c9364;
output c037;
output c4474;
output c221;
output c3164;
output c8312;
output c3371;
output c0424;
output c3161;
output c2202;
output c7110;
output c9417;
output c9170;
output c5411;
output c3214;
output c3333;
output c44;
output c4150;
output c8489;
output c2342;
output c9291;
output c4490;
output c5304;
output c2368;
output c9313;
output c5391;
output c819;
output c8475;
output c2498;
output c5359;
output c5481;
output c399;
output c4156;
output c6319;
output c799;
output c4144;
output c622;
output c3330;
output c2386;
output c6159;
output c9105;
output c5268;
output c0264;
output c6157;
output c8324;
output c89;
output c4455;
output c379;
output c8216;
output c317;
output c0116;
output c9201;
output c7184;
output c854;
output c5394;
output c2217;
output c920;
output c3339;
output c6189;
output c883;
output c6410;
output c0250;
output c0277;
output c2289;
output c9371;
output c6265;
output c3469;
output c3297;
output c6420;
output c5271;
output c9344;
output c0207;
output c045;
output c2444;
output c3413;
output c4113;
output c0385;
output c649;
output c8122;
output c870;
output c0157;
output c5178;
output c3408;
output c3184;
output c0473;
output c4205;
output c1350;
output c9274;
output c7442;
output c6414;
output c5159;
output c6389;
output c9412;
output c1416;
output c2388;
output c9432;
output c0342;
output c0186;
output c529;
output c671;
output c3298;
output c7365;
output c4402;
output c0370;
output c2182;
output c9378;
output c5305;
output c7351;
output c0299;
output c9311;
output c7439;
output c0413;
output c4355;
output c0396;
output c7467;
output c0346;
output c9114;
output c8280;
output c0195;
output c2452;
output c6120;
output c1330;
output c3238;
output c5353;
output c9230;
output c2218;
output c1241;
output c5262;
output c9196;
output c6151;
output c061;
output c6369;
output c5367;
output c0188;
output c5284;
output c8193;
output c49;
output c0106;
output c0338;
output c8104;
output c5339;
output c1410;
output c9222;
output c5297;
output c7194;
output c09;
output c9106;
output c867;
output c5167;
output c6273;
output c6210;
output c8283;
output c3499;
output c10;
output c9192;
output c4470;
output c6459;
output c6179;
output c891;
output c4466;
output c473;
output c2175;
output c2164;
output c433;
output c772;
output c4492;
output c244;
output c2367;
output c5211;
output c1101;
output c9250;
output c0241;
output c339;
output c2328;
output c5434;
output c8248;
output c478;
output c7232;
output c9257;
output c1110;
output c886;
output c67;
output c7322;
output c7116;
output c6388;
output c7413;
output c1319;
output c3273;
output c2149;
output c7319;
output c4212;
output c2381;
output c7266;
output c6400;
output c5377;
output c091;
output c1276;
output c5116;
output c3376;
output c579;
output c1339;
output c447;
output c5379;
output c6158;
output c1230;
output c4426;
output c2339;
output c7235;
output c3100;
output c3192;
output c6144;
output c7405;
output c6274;
output c1124;
output c0465;
output c0171;
output c0466;
output c547;
output c41;
output c7454;
output c158;
output c1310;
output c9182;
output c3444;
output c7287;
output c3105;
output c115;
output c3169;
output c6308;
output c6390;
output c3433;
output c1277;
output c9316;
output c4454;
output c022;
output c2222;
output c4127;
output c6342;
output c0365;
output c5149;
output c6366;
output c3322;
output c2301;
output c0148;
output c1362;
output c0129;
output c7384;
output c1121;
output c1199;
output c195;
output c6428;
output c4447;
output c0391;
output c7227;
output c192;
output c6258;
output c7483;
output c4171;
output c9403;
output c6486;
output c0232;
output c0136;
output c2267;
output c822;
output c4435;
output c0107;
output c7479;
output c923;
output c9171;
output c8204;
output c9237;
output c8398;
output c514;
output c1462;
output c2338;
output c6154;
output c6395;
output c8279;
output c2396;
output c6290;
output c4248;
output c455;
output c3128;
output c1443;
output c5356;
output c8288;
output c1120;
output c685;
output c775;
output c6294;
output c6362;
output c4190;
output c5404;
output c850;
output c9463;
output c581;
output c8289;
output c657;
output c79;
output c1445;
output c3436;
output c0209;
output c4219;
output c5263;
output c8227;
output c181;
output c7278;
output c9129;
output c4380;
output c6165;
output c9465;
output c5321;
output c4411;
output c6278;
output c6227;
output c8410;
output c392;
output c6344;
output c7226;
output c4174;
output c611;
output c4397;
output c8125;
output c8316;
output c911;
output c641;
output c9352;
output c5101;
output c9252;
output c252;
output c0360;
output c9308;
output c9430;
output c5476;
output c285;
output c0435;
output c6222;
output c9419;
output c3139;
output c9477;
output c8113;
output c5276;
output c6328;
output c0336;
output c2305;
output c0316;
output c4475;
output c7499;
output c7299;
output c8442;
output c6111;
output c8146;
output c0423;
output c6424;
output c5484;
output c7453;
output c2211;
output c4347;
output c7421;
output c1132;
output c7228;
output c8269;
output c3344;
output c0459;
output c542;
output c5322;
output c227;
output c8483;
output c5117;
output c8386;
output c1272;
output c2306;
output c5383;
output c8273;
output c0450;
output c827;
output c027;
output c0282;
output c5425;
output c4464;
output c7320;
output c4157;
output c9392;
output c345;
output c5317;
output c2195;
output c8425;
output c3275;
output c6364;
output c0302;
output c2291;
output c9442;
output c0133;
output c9218;
output c6141;
output c2303;
output c3449;
output c4365;
output c3200;
output c9464;
output c6195;
output c8328;
output c1313;
output c162;
output c1459;
output c549;
output c7166;
output c6322;
output c4181;
output c5290;
output c452;
output c928;
output c6445;
output c2242;
output c2167;
output c9101;
output c1258;
output c2349;
output c3257;
output c1232;
output c3248;
output c184;
output c7494;
output c5226;
output c816;
output c2274;
output c2102;
output c0353;
output c4356;
output c124;
output c6438;
output c9122;
output c8159;
output c1105;
output c4104;
output c2470;
output c237;
output c0397;
output c8195;
output c8349;
output c9333;
output c3290;
output c3425;
output c173;
output c6262;
output c4210;
output c258;
output c331;
output c386;
output c7482;
output c6163;
output c6481;
output c270;
output c562;
output c80;
output c5454;
output c95;
output c2207;
output c215;
output c0230;
output c8201;
output c8402;
output c3423;
output c8119;
output c145;
output c25;
output c8342;
output c2214;
output c5196;
output c6303;
output c640;
output c8361;
output c924;
output c2170;
output c3254;
output c2282;
output c7231;
output c0235;
output c9358;
output c4211;
output c8152;
output c1325;
output c0412;
output c6356;
output c487;
output c4324;
output c341;
output c0415;
output c3353;
output c1418;
output c1176;
output c5292;
output c058;
output c1100;
output c5291;
output c066;
output c052;
output c5361;
output c9314;
output c164;
output c678;
output c969;
output c1337;
output c986;
output c1379;
output c3461;
output c2288;
output c9318;
output c8352;
output c873;
output c7106;
output c4155;
output c28;
output c6187;
output c034;
output c990;
output c981;
output c8242;
output c7269;
output c463;
output c155;
output c5435;
output c5181;
output c4213;
output c3447;
output c9429;
output c1141;
output c8191;
output c7493;
output c9362;
output c5243;
output c1288;
output c3217;
output c8330;
output c863;
output c9359;
output c185;
output c4379;
output c362;
output c0482;
output c9306;
output c5352;
output c4390;
output c5384;
output c7476;
output c1218;
output c0165;
output c3334;
output c4363;
output c9469;
output c729;
output c17;
output c7271;
output c9110;
output c537;
output c1102;
output c6310;
output c2419;
output c2357;
output c5256;
output c4348;
output c43;
output c6145;
output c7464;
output c451;
output c8169;
output c8416;
output c2276;
output c2356;
output c5465;
output c5183;
output c7216;
output c3486;
output c1284;
output c367;
output c2421;
output c5238;
output c2151;
output c594;
output c4271;
output c1185;
output c661;
output c7262;
output c177;
output c1336;
output c9381;
output c1329;
output c0348;
output c438;
output c8311;
output c2366;
output c672;
output c2255;
output c5137;
output c4407;
output c3230;
output c9294;
output c3368;
output c2162;
output c6429;
output c9135;
output c127;
output c471;
output c8215;
output c948;
output c913;
output c1430;
output c9437;
output c8480;
output c3153;
output c773;
output c9273;
output c180;
output c4246;
output c5209;
output c8190;
output c5233;
output c8112;
output c0152;
output c1449;
output c6138;
output c5408;
output c9158;
output c7425;
output c5327;
output c6462;
output c7414;
output c5429;
output c1131;
output c5331;
output c0254;
output c4459;
output c6396;
output c1363;
output c5237;
output c6108;
output c1151;
output c4121;
output c183;
output c415;
output c9346;
output c1499;
output c6134;
output c4375;
output c9144;
output c2476;
output c4336;
output c1178;
output c9277;
output c1314;
output c1403;
output c0406;
output c218;
output c043;
output c7282;
output c893;
output c2129;
output c019;
output c683;
output c075;
output c621;
output c7441;
output c7422;
output c0287;
output c0301;
output c1437;
output c6323;
output c134;
output c6409;
output c0199;
output c2484;
output c9271;
output c565;
output c6149;
output c3207;
output c7459;
output c6105;
output c9130;
output c9492;
output c297;
output c0341;
output c414;
output c6192;
output c0490;
output c9104;
output c5494;
output c3314;
output c8116;
output c6401;
output c8213;
output c8249;
output c7160;
output c7465;
output c699;
output c298;
output c6218;
output c798;
output c0221;
output c2375;
output c4373;
output c6427;
output c140;
output c6169;
output c1296;
output c3189;
output c15;
output c088;
output c0382;
output c1381;
output c876;
output c6374;
output c1334;
output c482;
output c9426;
output c5451;
output c0326;
output c835;
output c8235;
output c0184;
output c4116;
output c64;
output c456;
output c7186;
output c0108;
output c3464;
output c3490;
output c9431;
output c378;
output c1451;
output c3243;
output c7100;
output c214;
output c7325;
output c4258;
output c9498;
output c3406;
output c8222;
output c5457;
output c6307;
output c8239;
output c9441;
output c2469;
output c75;
output c384;
output c9168;
output c4305;
output c1448;
output c4184;
output c4270;
output c561;
output c5169;
output c3131;
output c1485;
output c1260;
output c336;
output c494;
output c6360;
output c3427;
output c2461;
output c7156;
output c6152;
output c9157;
output c7433;
output c0163;
output c9155;
output c5370;
output c5388;
output c32;
output c9276;
output c849;
output c8180;
output c0357;
output c9217;
output c1190;
output c9467;
output c462;
output c6117;
output c453;
output c1414;
output c4341;
output c8210;
output c7280;
output c4484;
output c0121;
output c6119;
output c217;
output c1328;
output c4416;
output c83;
output c5333;
output c5498;
output c3276;
output c3385;
output c8189;
output c1467;
output c7449;
output c7143;
output c3201;
output c1281;
output c9375;
output c9478;
output c829;
output c2206;
output c8315;
output c4272;
output c66;
output c6408;
output c8382;
output c3155;
output c9137;
output c4256;
output c7332;
output c91;
output c5264;
output c7212;
output c833;
output c2464;
output c7387;
output c755;
output c2401;
output c7230;
output c9350;
output c4408;
output c1349;
output c5336;
output c06;
output c031;
output c728;
output c3326;
output c9483;
output c9440;
output c5344;
output c4240;
output c9423;
output c3381;
output c5376;
output c9332;
output c5395;
output c8135;
output c4228;
output c023;
output c691;
output c7406;
output c4206;
output c8114;
output c5398;
output c5401;
output c970;
output c8132;
output c3263;
output c796;
output c0364;
output c9156;
output c8344;
output c6340;
output c3389;
output c8117;
output c9424;
output c8131;
output c2361;
output c4225;
output c6256;
output c840;
output c914;
output c6475;
output c090;
output c9113;
output c1366;
output c0238;
output c7289;
output c3234;
output c3317;
output c3283;
output c1423;
output c7305;
output c7265;
output c8446;
output c4449;
output c3231;
output c086;
output c618;
output c2402;
output c2299;
output c5278;
output c523;
output c288;
output c3468;
output c3233;
output c9160;
output c0283;
output c4215;
output c5469;
output c1469;
output c1364;
output c9215;
output c588;
output c2408;
output c3439;
output c814;
output c5309;
output c5488;
output c6407;
output c7373;
output c4362;
output c3471;
output c9287;
output c5269;
output c2191;
output c1205;
output c8261;
output c788;
output c3250;
output c7334;
output c4382;
output c7285;
output c3411;
output c5135;
output c1390;
output c3154;
output c4441;
output c347;
output c8493;
output c0334;
output c0102;
output c499;
output c6276;
output c7213;
output c5208;
output c9210;
output c489;
output c96;
output c8142;
output c879;
output c0434;
output c2387;
output c9216;
output c6302;
output c2181;
output c0272;
output c951;
output c882;
output c2380;
output c2293;
output c3440;
output c8453;
output c5382;
output c1356;
output c0322;
output c6337;
output c5121;
output c655;
output c7119;
output c9163;
output c042;
output c6196;
output c1487;
output c493;
output c0208;
output c5141;
output c6259;
output c0497;
output c531;
output c8276;
output c9147;
output c9126;
output c2481;
output c5157;
output c6136;
output c3467;
output c432;
output c637;
output c9108;
output c2235;
output c2185;
output c4247;
output c2443;
output c6251;
output c369;
output c8424;
output c9283;
output c9482;
output c6143;
output c488;
output c3208;
output c4180;
output c3302;
output c6211;
output c570;
output c3218;
output c1386;
output c0476;
output c9260;
output c8441;
output c2404;
output c7208;
output c6468;
output c5172;
output c6365;
output c745;
output c2395;
output c5282;
output c8285;
output c5258;
output c1464;
output c20;
output c0320;
output c1139;
output c6288;
output c8338;
output c2315;
output c5217;
output c5340;
output c3492;
output c8270;
output c8259;
output c8336;
output c0369;
output c7209;
output c38;
output c0442;
output c0297;
output c169;
output c643;
output c0131;
output c0202;
output c659;
output c064;
output c370;
output c4401;
output c5129;
output c1119;
output c4141;
output c5330;
output c716;
output c5179;
output c4413;
output c2492;
output c7402;
output c448;
output c4383;
output c860;
output c2103;
output c8457;
output c1442;
output c1252;
output c0246;
output c3289;
output c3390;
output c4499;
output c3476;
output c2418;
output c789;
output c0194;
output c2493;
output c0444;
output c54;
output c3366;
output c7331;
output c563;
output c7171;
output c8452;
output c1153;
output c4478;
output c082;
output c6406;
output c248;
output c0408;
output c4238;
output c4126;
output c517;
output c3260;
output c5474;
output c8167;
output c7376;
output c2341;
output c6197;
output c4387;
output c6405;
output c1248;
output c6411;
output c0352;
output c3282;
output c2374;
output c3143;
output c7254;
output c832;
output c093;
output c0256;
output c2482;
output c5493;
output c27;
output c636;
output c780;
output c5274;
output c8110;
output c9384;
output c7327;
output c3113;
output c3288;
output c0261;
output c111;
output c0340;
output c5492;
output c3338;
output c597;
output c5369;
output c8439;
output c0447;
output c3117;
output c4360;
output c9136;
output c892;
output c4376;
output c437;
output c7218;
output c2264;
output c9462;
output c711;
output c4163;
output c3474;
output c7257;
output c0167;
output c5446;
output c8357;
output c8440;
output c7272;
output c865;
output c1179;
output c398;
output c4152;
output c7153;
output c3280;
output c0495;
output c2101;
output c5130;
output c1377;
output c6373;
output c0144;
output c2497;
output c8395;
output c3194;
output c190;
output c1491;
output c626;
output c495;
output c8293;
output c5229;
output c8109;
output c5485;
output c275;
output c9220;
output c5146;
output c8474;
output c995;
output c1419;
output c686;
output c6284;
output c8447;
output c3478;
output c4302;
output c8103;
output c9154;
output c9427;
output c063;
output c0178;
output c2156;
output c1365;
output c0237;
output c7313;
output c2158;
output c2209;
output c2355;
output c7463;
output c669;
output c8495;
output c0123;
output c0298;
output c2358;
output c4400;
output c9443;
output c974;
output c271;
output c1480;
output c2163;
output c7484;
output c653;
output c239;
output c0253;
output c165;
output c4403;
output c4396;
output c7233;
output c9118;
output c443;
output c548;
output c6147;
output c3309;
output c0337;
output c5176;
output c2337;
output c1173;
output c4280;
output c3183;
output c898;
output c8368;
output c3195;
output c45;
output c8198;
output c038;
output c360;
output c2463;
output c1374;
output c329;
output c0127;
output c5273;
output c146;
output c3300;
output c2316;
output c7137;
output c9336;
output c6190;
output c4453;
output c0488;
output c7193;
output c191;
output c8144;
output c29;
output c8484;
output c1264;
output c0117;
output c025;
output c3348;
output c6301;
output c080;
output c5473;
output c615;
output c2168;
output c6416;
output c7154;
output c1461;
output c4137;
output c4119;
output c1285;
output c6343;
output c9111;
output c1392;
output c6399;
output c0425;
output c0489;
output c3272;
output c2194;
output c4105;
output c4217;
output c7237;
output c6432;
output c697;
output c593;
output c9416;
output c823;
output c7337;
output c5109;
output c627;
output c2430;
output c7316;
output c256;
output c5477;
output c4175;
output c7105;
output c1287;
output c6476;
output c0471;
output c587;
output c4315;
output c0234;
output c2383;
output c1441;
output c0174;
output c3228;
output c2286;
output c2221;
output c187;
output c0168;
output c4434;
output c33;
output c0191;
output c355;
output c017;
output c3479;
output c8304;
output c6398;
output c8174;
output c5350;
output c7182;
output c2216;
output c5286;
output c6137;
output c676;
output c1492;
output c6208;
output c2309;
output c6126;
output c6131;
output c16;
output c9225;
output c4368;
output c3335;
output c8462;
output c3343;
output c7240;
output c2204;
output c7377;
output c9164;
output c4263;
output c9188;
output c4294;
output c6267;
output c2332;
output c774;
output c90;
output c6451;
output c782;
output c1208;
output c7368;
output c026;
output c5392;
output c9194;
output c5120;
output c9174;
output c4351;
output c2105;
output c5161;
output c5405;
output c6306;
output c8435;
output c4457;
output c6404;
output c771;
output c8260;
output c9327;
output c2153;
output c2499;
output c6317;
output c532;
output c9328;
output c6107;
output c9309;
output c3375;
output c6252;
output c7255;
output c8228;
output c815;
output c059;
output c8365;
output c7419;
output c9349;
output c5449;
output c1114;
output c4209;
output c830;
output c5188;
output c1335;
output c5442;
output c116;
output c3393;
output c721;
output c3212;
output c4494;
output c60;
output c4128;
output c797;
output c5200;
output c349;
output c3454;
output c0113;
output c88;
output c7437;
output c1169;
output c5266;
output c1460;
output c069;
output c5242;
output c2119;
output c2258;
output c0393;
output c9399;
output c6254;
output c2160;
output c979;
output c3173;
output c7381;
output c481;
output c1145;
output c7190;
output c00;
output c0120;
output c8267;
output c3104;
output c446;
output c0363;
output c2307;
output c5110;
output c1473;
output c630;
output c0491;
output c3421;
output c7288;
output c2475;
output c0362;
output c6241;
output c0244;
output c240;
output c0147;
output c5108;
output c0245;
output c6223;
output c2377;
output c9199;
output c4381;
output c8124;
output c7429;
output c9361;
output c474;
output c4448;
output c5173;
output c5125;
output c2399;
output c1409;
output c468;
output c614;
output c262;
output c5486;
output c2249;
output c4409;
output c9481;
output c3351;
output c8299;
output c1407;
output c7128;
output c8472;
output c8369;
output c7149;
output c5190;
output c3211;
output c2314;
output c673;
output c2370;
output c0179;
output c7261;
output c714;
output c2428;
output c3110;
output c3266;
output c690;
output c1295;
output c596;
output c739;
output c3424;
output c1495;
output c0333;
output c7430;
output c612;
output c4224;
output c521;
output c3239;
output c7452;
output c5275;
output c4214;
output c5366;
output c2416;
output c1217;
output c8298;
output c0343;
output c178;
output c2127;
output c0452;
output c1163;
output c2478;
output c1375;
output c3443;
output c3402;
output c174;
output c572;
output c524;
output c3190;
output c9224;
output c3213;
output c634;
output c0104;
output c1125;
output c0458;
output c2424;
output c266;
output c4233;
output c790;
output c8364;
output c2269;
output c7163;
output c7164;
output c1393;
output c9304;
output c123;
output c2362;
output c1297;
output c577;
output c2347;
output c1341;
output c8391;
output c1164;
output c2229;
output c3354;
output c143;
output c999;
output c824;
output c752;
output c694;
output c8467;
output c076;
output c2308;
output c2327;
output c4140;
output c235;
output c2465;
output c7343;
output c5417;
output c1438;
output c7108;
output c6495;
output c8188;
output c6353;
output c7124;
output c9382;
output c0124;
output c4405;
output c2155;
output c665;
output c6293;
output c0187;
output c3301;
output c032;
output c8466;
output c2186;
output c692;
output c4118;
output c6332;
output c0390;
output c9339;
output c7440;
output c759;
output c591;
output c3415;
output c6478;
output c2261;
output c555;
output c961;
output c4308;
output c7121;
output c6140;
output c677;
output c6326;
output c374;
output c942;
output c5131;
output c982;
output c1150;
output c1257;
output c130;
output c559;
output c4471;
output c6499;
output c0453;
output c1113;
output c3320;
output c8347;
output c7353;
output c2391;
output c7456;
output c439;
output c613;
output c617;
output c3145;
output c567;
output c5496;
output c743;
output c6245;
output c0463;
output c3414;
output c4309;
output c6118;
output c122;
output c246;
output c4151;
output c7344;
output c3456;
output c151;
output c6412;
output c9421;
output c2118;
output c9263;
output c5418;
output c650;
output c6419;
output c3223;
output c6494;
output c754;
output c7392;
output c4249;
output c3484;
output c7161;
output c7145;
output c4178;
output c8170;
output c1420;
output c7391;
output c8412;
output c5365;
output c7196;
output c9385;
output c4133;
output c3380;
output c5221;
output c0206;
output c3357;
output c65;
output c828;
output c0479;
output c8471;
output c3199;
output c9259;
output c2210;
output c1177;
output c267;
output c7400;
output c2384;
output c0419;
output c0140;
output c5112;
output c8305;
output c8448;
output c6191;
output c2169;
output c861;
output c3364;
output c9470;
output c7291;
output c9496;
output c660;
output c1138;
output c6123;
output c1213;
output c1225;
output c6460;
output c2233;
output c4139;
output c9191;
output c012;
output c2462;
output c1293;
output c520;
output c2489;
output c321;
output c5142;
output c9337;
output c2277;
output c0428;
output c9181;
output c817;
output c4143;
output c8225;
output c6183;
output c2285;
output c9301;
output c2146;
output c2494;
output c8383;
output c550;
output c6283;
output c0319;
output c0295;
output c5354;
output c5466;
output c469;
output c318;
output c7349;
output c3129;
output c2433;
output c337;
output c2198;
output c2265;
output c5342;
output c6376;
output c8179;
output c8417;
output c1496;
output c4106;
output c9373;
output c1427;
output c0486;
output c7357;
output c8303;
output c429;
output c0407;
output c324;
output c7431;
output c5414;
output c7385;
output c8476;
output c2310;
output c4235;
output c1466;
output c380;
output c6447;
output c0314;
output c7371;
output c4307;
output c6272;
output c960;
output c3132;
output c3347;
output c6232;
output c2224;
output c9117;
output c9310;
output c820;
output c9367;
output c5368;
output c0399;
output c4433;
output c0252;
output c8385;
output c8301;
output c0323;
output c393;
output c9267;
output c3107;
output c3379;
output c8129;
output c7223;
output c3442;
output c420;
output c1343;
output c6433;
output c4262;
output c1250;
output c4378;
output c7222;
output c8149;
output c7220;
output c9334;
output c5180;
output c3358;
output c9321;
output c5206;
output c585;
output c7292;
output c3497;
output c196;
output c9420;
output c7296;
output c160;
output c1109;
output c395;
output c8229;
output c4129;
output c255;
output c623;
output c2250;
output c4111;
output c5467;
output c925;
output c4176;
output c6383;
output c0233;
output c0303;
output c4424;
output c742;
output c5213;
output c0331;
output c1247;
output c9366;
output c1421;
output c8379;
output c5447;
output c4146;
output c440;
output c7246;
output c7315;
output c5204;
output c1453;
output c364;
output c047;
output c6479;
output c397;
output c9407;
output c5482;
output c7103;
output c53;
output c295;
output c5127;
output c738;
output c7200;
output c050;
output c9374;
output c1299;
output c0197;
output c1497;
output c0296;
output c4281;
output c5410;
output c4218;
output c0222;
output c3121;
output c070;
output c8292;
output c4237;
output c8105;
output c9132;
output c910;
output c9172;
output c786;
output c411;
output c741;
output c8237;
output c2459;
output c6361;
output c7273;
output c4292;
output c7297;
output c7408;
output c7481;
output c6129;
output c9100;
output c281;
output c6497;
output c2263;
output c8214;
output c765;
output c1388;
output c4417;
output c9228;
output c137;
output c0304;
output c0205;
output c3399;
output c4244;
output c6455;
output c4193;
output c2420;
output c9329;
output c0487;
output c7335;
output c089;
output c536;
output c0388;
output c3101;
output c6171;
output c8372;
output c1481;
output c6110;
output c4173;
output c8297;
output c5428;
output c4350;
output c9209;
output c357;
output c6423;
output c0443;
output c81;
output c3345;
output c6248;
output c053;
output c8246;
output c3321;
output c8405;
output c989;
output c5390;
output c9322;
output c2422;
output c4289;
output c5261;
output c2256;
output c4167;
output c8381;
output c0291;
output c654;
output c3158;
output c4115;
output c4458;
output c56;
output c6454;
output c7435;
output c8458;
output c7397;
output c8422;
output c6357;
output c1259;
output c9452;
output c6352;
output c9279;
output c114;
output c4136;
output c449;
output c316;
output c0135;
output c4110;
output c6346;
output c368;
output c6275;
output c7118;
output c9139;
output c2311;
output c4242;
output c7215;
output c4185;
output c9341;
output c132;
output c6168;
output c6164;
output c855;
output c5308;
output c9324;
output c2350;
output c1352;
output c7109;
output c0255;
output c2190;
output c3489;
output c9232;
output c0225;
output c4239;
output c2426;
output c8100;
output c0330;
output c2456;
output c8226;
output c5113;
output c1311;
output c3270;
output c4431;
output c8240;
output c1195;
output c2230;
output c6370;
output c390;
output c6325;
output c152;
output c3494;
output c6441;
output c9184;
output c35;
output c9115;
output c6239;
output c0321;
output c647;
output c6299;
output c1166;
output c553;
output c0403;
output c0351;
output c4283;
output c0156;
output c0139;
output c7293;
output c6381;
output c1360;
output c1144;
output c7139;
output c3446;
output c6484;
output c8490;
output c1317;
output c2150;
output c9236;
output c3258;
output c5307;
output c278;
output c5348;
output c6443;
output c9494;
output c1171;
output c2154;
output c4125;
output c422;
output c168;
output c5423;
output c8232;
output c0477;
output c9121;
output c3176;
output c7330;
output c9365;
output c0381;
output c5140;
output c1478;
output c4236;
output c7239;
output c5236;
output c0455;
output c4243;
output c4204;
output c8403;
output c2205;
output c793;
output c845;
output c1413;
output c4498;
output c6347;
output c769;
output c0276;
output c03;
output c7311;
output c0226;
output c167;
output c4349;
output c4130;
output c2466;
output c3222;
output c4399;
output c8337;
output c750;
output c4467;
output c1236;
output c4463;
output c2365;
output c6219;
output c7136;
output c2364;
output c2215;
output c8335;
output c0418;
output c0496;
output c8101;
output c7270;
output c930;
output c730;
output c8323;
output c2241;
output c0284;
output c6235;
output c344;
output c2227;
output c0173;
output c1127;
output c9167;
output c8221;
output c2373;
output c7480;
output c4311;
output c213;
output c4428;
output c2460;
output c4290;
output c1249;
output c3455;
output c1498;
output c5363;
output c3182;
output c3124;
output c3483;
output c9458;
output c0122;
output c1187;
output c7126;
output c9377;
output c3174;
output c5427;
output c687;
output c9454;
output c4221;
output c946;
output c1400;
output c1397;
output c2346;
output c5364;
output c2398;
output c5231;
output c7129;
output c3259;
output c0185;
output c8444;
output c844;
output c6329;
output c5478;
output c484;
output c099;
output c9265;
output c8492;
output c371;
output c4439;
output c6100;
output c2245;
output c4354;
output c054;
output c9317;
output c718;
output c2454;
output c7245;
output c8133;
output c1372;
output c2442;
output c9112;
output c497;
output c9444;
output c5316;
output c980;
output c9177;
output c6348;
output c0204;
output c4385;
output c5212;
output c6156;
output c7195;
output c6304;
output c4486;
output c8171;
output c8115;
output c4432;
output c7317;
output c9241;
output c5346;
output c0267;
output c492;
output c1389;
output c0378;
output c9459;
output c4429;
output c7411;
output c1161;
output c6139;
output c0105;
output c1251;
output c8384;
output c8429;
output c94;
output c5160;
output c3453;
output c818;
output c2319;
output c4323;
output c927;
output c7307;
output c5349;
output c166;
output c0414;
output c2304;
output c9240;
output c2121;
output c6173;
output c9315;
output c3306;
output c1353;
output c4197;
output c282;
output c9150;
output c3383;
output c0166;
output c6277;
output c1263;
output c3264;
output c1231;
output c0311;
output c0196;
output c2266;
output c3405;
output c7214;
output c991;
output c3287;
output c5184;
output c3392;
output c9248;
output c4196;
output c9468;
output c0361;
output c0126;
output c3127;
output c0141;
output c5495;
output c9298;
output c1378;
output c632;
output c7192;
output c1261;
output c9253;
output c9408;
output c2111;
output c5437;
output c949;
output c7360;
output c247;
output c0373;
output c6377;
output c9493;
output c887;
output c9233;
output c962;
output c568;
output c0438;
output c2248;
output c9124;
output c4377;
output c0273;
output c8238;
output c719;
output c0114;
output c1361;
output c8211;
output c3281;
output c1107;
output c778;
output c6437;
output c3328;
output c1143;
output c624;
output c5338;
output c0483;
output c1206;
output c04;
output c7367;
output c3171;
output c7249;
output c582;
output c9140;
output c3391;
output c4343;
output c767;
output c3232;
output c2125;
output c939;
output c2145;
output c1402;
output c2326;
output c9251;
output c725;
output c952;
output c2480;
output c7138;
output c8351;
output c0137;
output c0271;
output c445;
output c230;
output c314;
output c0324;
output c7135;
output c6220;
output c635;
output c3116;
output c4158;
output c4443;
output c3284;
output c8419;
output c083;
output c1398;
output c5326;
output c9405;
output c8243;
output c9219;
output c8375;
output c9395;
output c744;
output c396;
output c651;
output c0309;
output c1455;
output c1122;
output c0405;
output c2243;
output c389;
output c5432;
output c8310;
output c2120;
output c6242;
output c332;
output c9235;
output c5228;
output c9179;
output c8284;
output c6279;
output c3175;
output c6198;
output c9119;
output c8332;
output c69;
output c3115;
output c323;
output c5244;
output c0354;
output c1271;
output c2405;
output c897;
output c5416;
output c997;
output c7243;
output c7468;
output c9340;
output c3204;
output c1246;
output c670;
output c6102;
output c326;
output c9446;
output c3378;
output c4328;
output c186;
output c5298;
output c527;
output c9355;
output c2446;
output c573;
output c0437;
output c9134;
output c1180;
output c8287;
output c9166;
output c4358;
output c4123;
output c956;
output c1117;
output c2262;
output c8140;
output c4329;
output c5185;
output c5214;
output c8253;
output c3477;
output c0467;
output c4436;
output c896;
output c8404;
output c6393;
output c2268;
output c2435;
output c0379;
output c515;
output c5313;
output c6128;
output c513;
output c736;
output c3462;
output c4268;
output c6379;
output c491;
output c7345;
output c6237;
output c519;
output c78;
output c6349;
output c7378;
output c0462;
output c1183;
output c584;
output c4172;
output c4177;
output c2313;
output c3112;
output c642;
output c8136;
output c85;
output c6449;
output c2130;
output c4166;
output c5170;
output c7386;
output c1318;
output c890;
output c667;
output c8244;
output c1128;
output c141;
output c2174;
output c3495;
output c6266;
output c3267;
output c6368;
output c028;
output c5202;
output c6461;
output c992;
output c3432;
output c77;
output c7341;
output c3350;
output c6295;
output c7361;
output c3193;
output c7460;
output c461;
output c2112;
output c3370;
output c5280;
output c0177;
output c6338;
output c388;
output c3481;
output c0200;
output c2439;
output c4357;
output c6413;
output c4223;
output c014;
output c352;
output c6384;
output c8130;
output c1290;
output c2113;
output c1394;
output c0317;
output c959;
output c07;
output c039;
output c9379;
output c4254;
output c5436;
output c2485;
output c2344;
output c9143;
output c6394;
output c988;
output c8156;
output c9449;
output c1468;
output c2110;
output c8207;
output c610;
output c0410;
output c6327;
output c7252;
output c5162;
output c3418;
output c39;
output c770;
output c7113;
output c62;
output c8327;
output c847;
output c4326;
output c7306;
output c0101;
output c766;
output c1493;
output c6233;
output c8498;
output c0332;
output c9151;
output c1146;
output c6101;
output c0315;
output c8163;
output c0201;
output c8165;
output c9221;
output c6440;
output c1108;
output c3325;
output c762;
output c7210;
output c4496;
output c4296;
output c3369;
output c0429;
output c4389;
output c226;
output c7275;
output c1412;
output c881;
output c61;
output c9331;
output c2179;
output c5166;
output c0110;
output c040;
output c2417;
output c5303;
output c5443;
output c862;
output c1227;
output c1494;
output c757;
output c5153;
output c2188;
output c2231;
output c6113;
output c92;
output c2197;
output c8223;
output c937;
output c161;
output c2192;
output c5192;
output c2240;
output c8437;
output c2474;
output c9448;
output c2226;
output c2390;
output c2491;
output c8183;
output c3373;
output c4427;
output c342;
output c7451;
output c2292;
output c020;
output c7338;
output c9489;
output c6217;
output c7415;
output c1415;
output c2176;
output c7276;
output c9266;
output c327;
output c3295;
output c7224;
output c274;
output c441;
output c4202;
output c0150;
output c8331;
output c6418;
output c1126;
output c8141;
output c0153;
output c056;
output c0169;
output c2161;
output c3459;
output c3488;
output c9497;
output c6285;
output c7347;
output c3146;
output c2132;
output c5490;
output c2290;
output c9270;
output c3387;
output c2279;
output c7173;
output c0262;
output c8454;
output c0356;
output c751;
output c8290;
output c7486;
output c8418;
output c7478;
output c5285;
output c8485;
output c3311;
output c3319;
output c5463;
output c934;
output c1192;
output c2140;
output c5216;
output c8317;
output c3388;
output c6312;
output c5415;
output c4282;
output c9203;
output c7323;
output c9495;
output c1483;
output c9438;
output c8274;
output c9425;
output c044;
output c3316;
output c525;
output c7498;
output c5422;
output c6260;
output c276;
output c8247;
output c1387;
output c416;
output c551;
output c9293;
output c5409;
output c787;
output c7181;
output c3332;
output c425;
output c8450;
output c3224;
output c5281;
output c4488;
output c1214;
output c675;
output c9435;
output c9487;
output c8230;
output c1175;
output c2109;
output c423;
output c6316;
output c4461;
output c0394;
output c5253;
output c885;
output c546;
output c7446;
output c6180;
output c8496;
output c8377;
output c0281;
output c884;
output c2189;
output c1216;
output c1159;
output c0251;
output c5421;
output c5351;
output c5223;
output c7418;
output c8306;
output c713;
output c2302;
output c3466;
output c9281;
output c7492;
output c1140;
output c7466;
output c3496;
output c4481;
output c674;
output c7141;
output c1160;
output c8318;
output c6103;
output c4421;
output c3185;
output c3384;
output c4288;
output c2208;
output c932;
output c0210;
output c812;
output c9123;
output c6280;
output c0224;
output c966;
output c4131;
output c5224;
output c7238;
output c391;
output c5193;
output c834;
output c311;
output c0402;
output c6243;
output c0344;
output c0454;
output c7458;
output c365;
output c7417;
output c1253;
output c746;
output c916;
output c2436;
output c2148;
output c5375;
output c9288;
output c7157;
output c260;
output c530;
output c6182;
output c620;
output c197;
output c2213;
output c8363;
output c3416;
output c8464;
output c7403;
output c6314;
output c8161;
output c912;
output c3285;
output c3470;
output c2128;
output c5396;
output c8463;
output c6367;
output c1331;
output c8459;
output c0151;
output c99;
output c1165;
output c9434;
output c7295;
output c4231;
output c6363;
output c3216;
output c7107;
output c8320;
output c7134;
output c0481;
output c8120;
output c733;
output c3156;
output c7219;
output c6320;
output c8296;
output c1358;
output c662;
output c5480;
output c6135;
output c8151;
output c1170;
output c2336;
output c7247;
output c8173;
output c4208;
output c7168;
output c024;
output c511;
output c8209;
output c9109;
output c545;
output c3434;
output c1269;
output c7180;
output c3170;
output c1439;
output c0451;
output c8212;
output c3142;
output c6477;
output c0366;
output c6230;
output c727;
output c7374;
output c2486;
output c4480;
output c2296;
output c4372;
output c9173;
output c0243;
output c4164;
output c1327;
output c1115;
output c7201;
output c841;
output c6444;
output c7286;
output c3163;
output c125;
output c2257;
output c7179;
output c590;
output c4330;
output c9387;
output c0411;
output c5174;
output c1354;
output c4253;
output c955;
output c2440;
output c3219;
output c0214;
output c5107;
output c0203;
output c046;
output c6313;
output c8262;
output c5372;
output c0325;
output c9372;
output c2166;
output c2177;
output c7443;
output c933;
output c7355;
output c0358;
output c0193;
output c1436;
output c9289;
output c0374;
output c426;
output c8389;
output c3293;
output c4293;
output c5100;
output c574;
output c5407;
output c4485;
output c0265;
output c8258;
output c6309;
output c8314;
output c0431;
output c5397;
output c8397;
output c3177;
output c679;
output c1282;
output c0145;
output c8387;
output c8252;
output c0492;
output c0318;
output c9107;
output c9307;
output c8482;
output c2199;
output c2447;
output c2320;
output c1191;
output c2468;
output c6115;
output c3159;
output c8218;
output c4335;
output c4191;
output c9187;
output c9245;
output c4444;
output c385;
output c6350;
output c9131;
output c7150;
output c6496;
output c9256;
output c5148;
output c2318;
output c3329;
output c5497;
output c5270;
output c3111;
output c6446;
output c1431;
output c3202;
output c4412;
output c795;
output c737;
output c71;
output c7142;
output c0306;
output c3346;
output c485;
output c6333;
output c543;
output c4487;
output c6355;
output c72;
output c9175;
output c7244;
output c7101;
output c5385;
output c2144;
output c9491;
output c348;
output c7277;
output c5154;
output c5195;
output c9299;
output c1200;
output c557;
output c5487;
output c7203;
output c6206;
output c9223;
output c3227;
output c2219;
output c4327;
output c578;
output c121;
output c6397;
output c7303;
output c4265;
output c015;
output c2172;
output c6386;
output c4260;
output c1417;
output c2431;
output c8353;
output c8333;
output c2467;
output c1482;
output c3123;
output c0484;
output c7301;
output c2393;
output c6194;
output c3118;
output c628;
output c1338;
output c24;
output c8157;
output c4319;
output c7178;
output c4321;
output c8455;
output c889;
output c6224;
output c899;
output c1244;
output c6127;
output c693;
output c724;
output c9214;
output c3397;
output c6124;
output c0242;
output c3114;
output c6253;
output c682;
output c0383;
output c3179;
output c5234;
output c3152;
output c4497;
output c5357;
output c6286;
output c216;
output c664;
output c055;
output c943;
output c1324;
output c5300;
output c7326;
output c6448;
output c9485;
output c6287;
output c8147;
output c5114;
output c575;
output c4199;
output c684;
output c7336;
output c8106;
output c1411;
output c983;
output c2473;
output c552;
output c1149;
output c071;
output c480;
output c8436;
output c418;
output c5119;
output c953;
output c1474;
output c7485;
output c6422;
output c5453;
output c1359;
output c954;
output c098;
output c7366;
output c2142;
output c7167;
output c334;
output c496;
output c6185;
output c7380;
output c8185;
output c9127;
output c0132;
output c0494;
output c0274;
output c135;
output c1489;
output c4279;
output c02;
output c0236;
output c564;
output c4179;
output c0172;
output c0142;
output c3465;
output c3149;
output c8264;
output c7497;
output c1396;
output c3365;
output c5134;
output c0111;
output c5470;
output c9204;
output c73;
output c5360;
output c296;
output c8313;
output c4313;
output c836;
output c129;
output c7352;
output c335;
output c6229;
output c888;
output c5445;
output c858;
output c1104;
output c6473;
output c794;
output c261;
output c7382;
output c5186;
output c5155;
output c220;
output c1267;
output c291;
output c0240;
output c6249;
output c2200;
output c8366;
output c852;
output c6457;
output c6380;
output c781;
output c4367;
output c273;
output c1196;
output c5272;
output c571;
output c3296;
output c3400;
output c0384;
output c3168;
output c6247;
output c0100;
output c4132;
output c8340;
output c4423;
output c4338;
output c6472;
output c150;
output c7423;
output c6493;
output c554;
output c8358;
output c7469;
output c9190;
output c9409;
output c087;
output c5106;
output c569;
output c646;
output c4274;
output c8341;
output c7383;
output c110;
output c4489;
output c3102;
output c994;
output c7491;
output c9302;
output c3236;
output c1174;
output c0231;
output c0347;
output c9356;
output c0130;
output c2458;
output c4425;
output c6450;
output c9480;
output c1384;
output c0387;
output c7474;
output c1315;
output c9268;
output c0430;
output c4304;
output c3205;
output c224;
output c5462;
output c475;
output c232;
output c55;
output c666;
output c8362;
output c5265;
output c6209;
output c6385;
output c97;
output c0456;
output c7390;
output c3165;
output c3396;
output c6244;
output c0161;
output c4422;
output c539;
output c2225;
output c619;
output c2371;
output c2223;
output c5215;
output c3210;
output c4226;
output c1348;
output c430;
output c4394;
output c9476;
output c971;
output c3361;
output c8206;
output c1168;
output c6268;
output c5296;
output c3491;
output c7302;
output c5430;
output c2322;
output c560;
output c0190;
output c2159;
output c287;
output c3448;
output c3367;
output c011;
output c1220;
output c0175;
output c0170;
output c5230;
output c696;
output c2331;
output c8456;
output c3186;
output c0441;
output c535;
output c6172;
output c0307;
output c918;
output c292;
output c8241;
output c8148;
output c330;
output c2143;
output c4101;
output c1198;
output c9398;
output c4160;
output c1357;
output c5460;
output c147;
output c6467;
output c8487;
output c8478;
output c6109;
output c1401;
output c8250;
output c5240;
output c9400;
output c848;
output c9353;
output c6466;
output c40;
output c2187;
output c1262;
output c6199;
output c5128;
output c0310;
output c5334;
output c6174;
output c4114;
output c7475;
output c4353;
output c6184;
output c7146;
output c7455;
output c3120;
output c5301;
output c376;
output c7472;
output c3180;
output c9338;
output c4220;
output c3349;
output c5143;
output c5419;
output c8348;
output c3498;
output c747;
output c3151;
output c284;
output c7364;
output c236;
output c7379;
output c698;
output c859;
output c5201;
output c779;
output c7148;
output c2329;
output c9290;
output c7409;
output c2410;
output c5295;
output c8411;
output c0345;
output c9159;
output c4342;
output c3360;
output c8162;
output c1283;
output c9335;
output c0469;
output c663;
output c6257;
output c2104;
output c8445;
output c6296;
output c6203;
output c7362;
output c926;
output c8123;
output c9473;
output c1286;
output c878;
output c1254;
output c5145;
output c8449;
output c3404;
output c785;
output c5205;
output c5426;
output c6112;
output c82;
output c777;
output c7125;
output c030;
output c1432;
output c8281;
output c9345;
output c4391;
output c0433;
output c120;
output c9433;
output c1292;
output c9138;
output c5345;
output c5220;
output c3265;
output c6300;
output c7151;
output c1294;
output c8200;
output c6255;
output c1477;
output c4162;
output c1162;
output c8278;
output c8370;
output c720;
output c1355;
output c0217;
output c1435;
output c4194;
output c8194;
output c3294;
output c8160;
output c2389;
output c645;
output c9243;
output c533;
output c251;
output c7274;
output c4317;
output c0118;
output c0219;
output c3122;
output c4479;
output c5439;
output c8309;
output c5461;
output c5163;
output c435;
output c680;
output c2228;
output c3188;
output c2352;
output c6490;
output c8461;
output c9343;
output c7199;
output c996;
output c2400;
output c756;
output c241;
output c8277;
output c466;
output c4259;
output c085;
output c8134;
output c8164;
output c8378;
output c1383;
output c9254;
output c265;
output c6177;
output c0420;
output c6482;
output c86;
output c2238;
output c9246;
output c5133;
output c760;
output c7198;
output c2147;
output c14;
output c51;
output c0278;
output c977;
output c13;
output c142;
output c5399;
output c9285;
output c095;
output c4188;
output c0257;
output c87;
output c0290;
output c9213;
output c9439;
output c9428;
output c2157;
output c0329;
output c3226;
output c6391;
output c7434;
output c312;
output c3451;
output c2429;
output c2330;
output c5252;
output c8390;
output c3374;
output c7298;
output c723;
output c710;
output c2427;
output c7445;
output c1342;
output c1463;
output c1157;
output c629;
output c1447;
output c2236;
output c4276;
output c3412;
output c7473;
output c8322;
output c1194;
output c3229;
output c8271;
output c8205;
output c6458;
output c6298;
output c978;
output c3308;
output c8308;
output c7197;
output c1202;
output c1193;
output c7290;
output c0279;
output c1326;
output c3291;
output c4201;
output c7175;
output c1446;
output c128;
output c5324;
output c188;
output c783;
output c3352;
output c1488;
output c631;
output c9369;
output c1452;
output c7471;
output c5413;
output c1369;
output c1245;
output c156;
output c950;
output c153;
output c36;
output c875;
output c7127;
output c1300;
output c6442;
output c4301;
output c6372;
output c0372;
output c7170;
output c7144;
output c3355;
output c0249;
output c5210;
output c8468;
output c7304;
output c1370;
output c598;
output c2345;
output c5412;
output c9410;
output c3377;
output c4462;
output c1433;
output c350;
output c8376;
output c2237;
output c0474;
output c5335;
output c2437;
output c5250;
output c242;
output c0109;
output c9238;
output c6261;
output c5343;
output c0212;
output c1426;
output c1405;
output c7177;
output c8427;
output c264;
output c375;
output c2457;
output c4419;
output c6270;
output c0115;
output c8451;
output c2477;
output c6392;
output c7263;
output c2479;
output c6498;
output c6345;
output c4153;
output c5171;
output c1256;
output c2385;
output c387;
output c0260;
output c5151;
output c7358;
output c9415;
output c9319;
output c1312;
output c1203;
output c4370;
output c7487;
output c2114;
output c0181;
output c7206;
output c072;
output c0125;
output c0192;
output c880;
output c57;
output c6250;
output c361;
output c171;
output c1472;
output c7388;
output c3318;
output c7211;
output c9312;
output c4477;
output c472;
output c5329;
output c753;
output c4159;
output c0227;
output c7426;
output c1197;
output c2283;
output c8491;
output c6334;
output c8396;
output c5306;
output c5222;
output c8192;
output c3493;
output c9347;
output c7267;
output c424;
output c7241;
output c5386;
output c356;
output c7410;
output c30;
output c9457;
output c23;
output c9202;
output c4303;
output c8128;
output c0149;
output c7395;
output c1450;
output c5194;
output c4138;
output c2423;
output c3292;
output c1490;
output c975;
output c6421;
output c0349;
output c1215;
output c4266;
output c6311;
output c5402;
output c6452;
output c3394;
output c7123;
output c7359;
output c412;
output c3382;
output c8367;
output c6453;
output c4186;
output c5197;
output c6439;
output c761;
output c3209;
output c5455;
output c5294;
output c290;
output c259;
output c7488;
output c2298;
output c2407;
output c3419;
output c0448;
output c163;
output c915;
output c7188;
output c018;
output c417;
output c4275;
output c3452;
output c394;
output c6212;
output c1280;
output c0213;
output c0355;
output c074;
output c776;
output c7189;
output c2122;
output c681;
output c6204;
output c5187;
output c648;
output c9142;
output c3136;
output c9120;
output c1406;
output c7162;
output c3438;
output c2406;
output c5393;
output c4165;
output c2165;
output c1106;
output c119;
output c9389;
output c229;
output c5115;
output c9286;
output c0380;
output c9165;
output c8138;
output c2259;
output c4222;
output c5314;
output c6456;
output c5472;
output c5255;
output c3303;
output c3359;
output c3395;
output c2323;
output c5124;
output c1444;
output c4482;
output c1385;
output c1155;
output c2441;
output c5302;
output c842;
output c021;
output c6387;
output c372;
output c3215;
output c3472;
output c748;
output c7279;
output c9295;
output c9396;
output c7130;
output c9261;
output c9226;
output c1228;
output c7398;
output c442;
output c633;
output c48;
output c688;
output c2409;
output c8172;
output c2239;
output c4440;
output c6489;
output c1137;
output c2376;
output c1306;
output c9460;
output c9205;
output c8356;
output c1134;
output c5424;
output c2312;
output c3261;
output c3429;
output c029;
output c3130;
output c0143;
output c3450;
output c3401;
output c987;
output c2115;
output c658;
output c8217;
output c4392;
output c9284;
output c4261;
output c7204;
output c9186;
output c792;
output c9200;
output c2378;
output c383;
output c599;
output c3441;
output c2425;
output c294;
output c3147;
output c0308;
output c041;
output c8121;
output c4318;
output c077;
output c544;
output c4108;
output c486;
output c7172;
output c63;
output c7496;
output c8118;
output c6382;
output c7294;
output c1142;
output c9330;
output c346;
output c5380;
output c7169;
output c243;
output c1309;
output c8150;
output c3268;
output c7329;
output c1279;
output c2152;
output c3437;
output c1476;
output c3305;
output c5403;
output c319;
output c5245;
output c1428;
output c6153;
output c5219;
output c2244;
output c921;
output c7396;
output c58;
output c6426;
output c1130;
output c3252;
output c6207;
output c112;
output c6471;
output c8102;
output c5293;
output c3422;
output c1211;
output c457;
output c0293;
output c2173;
output c6483;
output c9269;
output c0154;
output c1308;
output c2413;
output c465;
output c8282;
output c895;
output c6166;
output c6205;
output c831;
output c5475;
output c7420;
output c4352;
output c7462;
output c7268;
output c7187;
output c7225;
output c8346;
output c0416;
output c5251;
output c3148;
output c4420;
output c1268;
output c957;
output c1298;
output c1346;
output c035;
output c0288;
output c2412;
output c3426;
output c1382;
output c7155;
output c9445;
output c2334;
output c490;
output c5118;
output c9411;
output c763;
output c431;
output c968;
output c9278;
output c1265;
output c864;
output c4117;
output c6434;
output c9471;
output c4369;
output c0269;
output c0198;
output c338;
output c419;
output c067;
output c2117;
output c0398;
output c3253;
output c6297;
output c289;
output c2455;
output c5168;
output c0119;
output c2351;
output c2234;
output c2201;
output c9388;
output c460;
output c944;
output c8469;
output c1344;
output c8414;
output c2382;
output c1471;
output c3480;
output c5132;
output c3286;
output c3172;
output c9185;
output c113;
output c1289;
output c8307;
output c9125;
output c5257;
output c3463;
output c3269;
output c5406;
output c3262;
output c9227;
output c2275;
output c6417;
output c8430;
output c7363;
output c117;
output c6150;
output c9180;
output c3409;
output c0134;
output c172;
output c073;
output c3435;
output c2449;
output c1425;
output c2193;
output c0128;
output c1116;
output c1135;
output c1184;
output c4250;
output c8219;
output c4393;
output c1371;
output c872;
output c7165;
output c9303;
output c470;
output c381;
output c1484;
output c6167;
output c3126;
output c0228;
output c5318;
output c8181;
output c7207;
output c8393;
output c0189;
output c8155;
output c1399;
output c2108;
output c8400;
output c9234;
output c7389;
output c9418;
output c427;
output c4473;
output c839;
output c4109;
output c47;
output c516;
output c74;
output c2325;
output c2134;
output c5440;
output c6465;
output c9323;
output c4445;
output c7183;
output c5358;
output c7217;
output c7122;
output c6354;
output c4468;
output c1226;
output c0313;
output c668;
output c6234;
output c9229;
output c652;
output c5499;
output c0176;
output c212;
output c4232;
output c8434;
output c5152;
output c9249;
output c7102;
output c0328;
output c4107;
output c7251;
output c9474;
output c3372;
output c6425;
output c9297;
output c4230;
output c7354;
output c9275;
output c8432;
output c1224;
output c479;
output c5471;
output c9128;
output c5103;
output c5158;
output c936;
output c4298;
output c5156;
output c4297;
output c3240;
output c2116;
output c7324;
output c4414;
output c857;
output c7284;
output c31;
output c0138;
output c8168;
output c1181;
output c9456;
output c8470;
output c8202;
output c8158;
output c6200;
output c3178;
output c3220;
output c7394;
output c4207;
output c2450;
output c5433;
output c5147;
output c2273;
output c639;
output c2490;
output c211;
output c6114;
output c9351;
output c19;
output c4320;
output c8392;
output c7477;
output c0268;
output c428;
output c1404;
output c269;
output c9212;
output c1212;
output c1274;
output c5479;
output c0229;
output c315;
output c963;
output c9393;
output c0285;
output c93;
output c2297;
output c9193;
output c4456;
output c5381;
output c313;
output c6339;
output c1424;
output c2203;
output c0155;
output c7404;
output c2392;
output c1147;
output c7234;
output c8254;
output c1154;
output c328;
output c9258;
output c4182;
output c8176;
output c458;
output c6221;
output c2247;
output c8497;
output c3460;
output c9264;
output c3485;
output c4241;
output c4295;
output c5279;
output c4103;
output c5450;
output c068;
output c084;
output c5203;
output c9455;
output c272;
output c8184;
output c6148;
output c7120;
output c4460;
output c9152;
output c3166;
output c3487;
output c051;
output c9255;
output c4374;
output c7112;
output c52;
output c8394;
output c7308;
output c7457;
output c837;
output c6282;
output c3140;
output c223;
output c5320;
output c2360;
output c5136;
output c0280;
output c7399;
output c1367;
output c2432;
output c351;
output c1275;
output c2232;
output c144;
output c9189;
output c5389;
output c8388;
output c0460;
output c6228;
output c8178;
output c7432;
output c976;
output c3304;
output c9436;
output c9296;
output c148;
output c0400;
output c9390;
output c343;
output c2139;
output c4100;
output c984;
output c4491;
output c76;
output c1316;
output c5341;
output c353;
output c9262;
output c9153;
output c8196;
output c2434;
output c6402;
output c644;
output c5235;
output c2253;
output c3157;
output c715;
output c5456;
output c3191;
output c5448;
output c7132;
output c3336;
output c6436;
output c2496;
output c919;
output c3162;
output c6491;
output c1368;
output c2184;
output c1351;
output c6430;
output c0220;
output c131;
output c0401;
output c4442;
output c625;
output c9357;
output c0446;
output c250;
output c0376;
output c231;
output c4371;
output c249;
output c228;
output c8245;
output c9282;
output c580;
output c9451;
output c4384;
output c3187;
output c940;
output c3458;
output c8236;
output c7159;
output c5347;
output c5191;
output c149;
output c6469;
output c5111;
output c3430;
output c4438;
output c194;
output c0392;
output c967;
output c5483;
output c0103;
output c5139;
output c5373;
output c3242;
output c68;
output c0493;
output c6291;
output c5458;
output c9479;
output c6415;
output c583;
output c9475;
output c5325;
output c5452;
output c3249;
output c279;
output c0461;
output c097;
output c540;
output c1129;
output c538;
output c726;
output c3103;
output c3323;
output c7229;
output c1458;
output c851;
output c9208;
output c9383;
output c0359;
output c941;
output c9394;
output c5175;
output c096;
output c3221;
output c016;
output c4334;
output c6116;
output c126;
output c3274;
output c1322;
output c712;
output c2141;
output c6130;
output c175;
output c0464;
output c7470;
output c5489;
output c0158;
output c4415;
output c1255;
output c0480;
output c157;
output c8325;
output c4154;
output c222;
output c4388;
output c5387;
output c3363;
output c7444;
output c22;
output c9391;
output c4195;
output c3340;
output c3277;
output c5189;
output c9305;
output c0312;
output c0112;
output c8409;
output c7250;
output c8380;
output c8275;
output c4344;
output c874;
output c0389;
output c7264;
output c8428;
output c8272;
output c8255;
output c0270;
output c3482;
output c2403;
output c6485;
output c5299;
output c4418;
output c2414;
output c3247;
output c0286;
output c3106;
output c065;
output c3256;
output c8126;
output c2348;
output c0182;
output c9272;
output c8319;
output c6263;
output c8355;
output c3337;
output c1237;
output c512;
output c4316;
output c5283;
output c2353;
output c7375;
output c8399;
output c7205;
output c9103;
output c0215;
output c8256;
output c354;
output c9499;
output c1186;
output c286;
output c7115;
output c9146;
output c5198;
output c2124;
output c2394;
output c8145;
output c0432;
output c3181;
output c2287;
output c3407;
output c0485;
output c1204;
output c3417;
output c5199;
output c7340;
output c4149;
output c6231;
output c938;
output c6202;
output c7253;
output c3134;
output c9466;
output c922;
output c768;
output c8197;
output c4410;
output c0478;
output c5182;
output c0468;
output c1304;
output c7104;
output c6358;
output c6281;
output c0183;
output c4277;
output c9149;
output c592;
output c2123;
output c7283;
output c9141;
output c4483;
output c8265;
output c5123;
output c34;
output c6464;
output c9195;
output c9176;
output c2321;
output c0475;
output c84;
output c0300;
output c6186;
output c3150;
output c7489;
output c7450;
output c9486;
output c764;
output c1273;
output c199;
output c8407;
output c9325;
output c868;
output c3206;
output c3203;
output c7356;
output c2445;
output c9348;
output c9133;
output c1112;
output c5225;
output c8406;
output c695;
output c8401;
output c0377;
output c277;
output c3167;
output c3225;
output c8345;
output c6403;
output c6175;
output c8286;
output c2171;
output c1172;
output c0180;
output c6188;
output c8360;
output c722;
output c0422;
output c2138;
output c9292;
output c7372;
output c6236;
output c638;
output c4169;
output c5438;
output c6214;
output c1422;
output c0305;
output c8479;
output c6264;
output c4269;
output c0275;
output c1233;
output c359;
output c3237;
output c4291;
output c1219;
output c6292;
output c6213;
output c0472;
output c01;
output c6324;
output c0294;
output c4331;
output c5288;
output c811;
output c092;
output c4267;
output c732;
output c1486;
output c5441;
output c5444;
output c856;
output c0368;
output c3362;
output c4170;
output c3133;
output c2272;
output c7350;
output c1307;
output c8111;
output c8359;
output c9376;
output c5420;
output c810;
output c717;
output c7424;
output c4284;
output c254;
output c7346;
output c4345;
output c5126;
output c7258;
output c877;
output c1209;
output c2133;
output c421;
output c1465;
output c4406;
output c057;
output c081;
output c0247;
output c1440;
output c2251;
output c9397;
output c5277;
output c4278;
output c4145;
output c9239;
output c2438;
output c4446;
output c6155;
output c6160;
output c9354;
output c0350;
output c5362;
output c6178;
output c8420;
output c6470;
output c7242;
output c253;
output c826;
output c079;
output c179;
output c6269;
output c6378;
output c5232;
output c1156;
output c6315;
output c7202;
output c42;
output c3108;
output c8334;
output c3313;
output c4192;
output c3324;
output c8224;
output c0289;
output c5227;
output c5218;
output c8465;
output c9488;
output c7191;
output c182;
output c5468;
output c0371;
output c6289;
output c7370;
output c5249;
output c498;
output c2106;
output c7461;
output c8231;
output c8421;
output c998;
output c3251;
output c1457;
output c2343;
output c3431;
output c1133;
output c947;
output c7321;
output c4333;
output c4287;
output c5254;
output c1238;
output c5315;
output c3403;
output c1305;
output c510;
output c791;
output c310;
output c9161;
output c8300;
output c9380;
output c7428;
output c9247;
output c8321;
output c234;
output c0439;
output c869;
output c8329;
output c5260;
output c8208;
output c9490;
output c476;
output c6330;
output c7111;
output c2137;
output c4476;
output c4465;
output c3398;
output c4124;
output c3342;
output c5289;
output c2100;
output c1376;
output c9198;
output c325;
output c9326;
output c2196;
output c1323;
output c9207;
output c6480;
output c0499;
output c1242;
output c5337;
output c4102;
output c7176;
output c2372;
output c6226;
output c5355;
output c7312;
output c1434;
output c7256;
output c6125;
output c4189;
output c541;
output c3235;
output c9320;
output c333;
output c566;
output c8408;
output c340;
output c576;
output c5319;
output c4273;
output c1302;
output c70;
output c2483;
output c4187;
output c2317;
output c4322;
output c993;
output c4310;
output c0211;
output c12;
output c078;
output c373;
output c0162;
output c0335;
output c9178;
output c245;
output c11;
output c5459;
output c8139;
output c3245;
output c483;
output c9169;
output c7174;
output c0159;
output c2280;
output c377;
output c3327;
output c0436;
output c846;
output c5332;
output c6121;
output c3410;
output c1391;
output c8350;
output c0386;
output c3331;
output c7281;
output c595;
output c9404;
output c9461;
output c4346;
output c6246;
output c8175;
output c8251;
output c6225;
output c0248;
output c6161;
output c0292;
output c2212;
output c7117;
output c4452;
output c2354;
output c4216;
output c7412;
output c8302;
output c98;
output c6201;
output c8233;
output c740;
output c894;
output c2488;
output c825;
output c263;
output c8266;
output c5177;
output c4398;
output c964;
output c9450;
output c7140;
output c5150;
output c3307;
output c8413;
output c2260;
output c4285;
output c0239;
output c2136;
output c036;
output c9183;
output c0421;
output c2220;
output c5323;
output c8499;
output c935;
output c0164;
output c4495;
output c871;
output c0470;
output c1332;
output c8473;
output c7436;
output c3244;
output c4314;
output c210;
output c1167;
output c843;
output c136;
output c0417;
output c233;
output c2180;
output c1291;
output c1429;
output c6240;
output c929;
output c4148;
output c8443;
output c1479;
output c4183;
output c133;
output c8143;
output c0146;
output c410;
output c299;
output c8268;
output c1240;
output c4430;
output c7158;
output c1243;
output c283;
output c931;
output c8431;
output c4332;
output c4286;
output c5464;
output c6474;
output c4404;
output c9453;
output c59;
output c0367;
output c219;
output c2359;
output c972;
output c1111;
output c9422;
output c450;
output c4493;
output c689;
output c1207;
output c4395;
output c9401;
output c6488;
output c0258;
output c784;
output c2324;
output c7133;
output c4472;
output c6336;
output c2411;
output c1320;
output c4251;
output c4312;
output c0160;
output c0404;
output c413;
output c049;
output c5310;
output c7309;
output c2281;
output c9342;
output c0449;
output c7407;
output c2254;
output c5102;
output c9116;
output c459;
output c3312;
output c5164;
output c534;
output c8137;
output c8220;
output c973;
output c3135;
output c8263;
output c8294;
output c8423;
output c2448;
output c4142;
output c37;
output c363;
output c0339;
output c0426;
output c616;
output c2487;
output c6216;
output c2278;
output c1222;
output c5431;
output c731;
output c1380;
output c0327;
output c2131;
output c8488;
output c189;
output c8295;
output c2270;
output c2252;
output c2284;
output c1123;
output c1475;
output c280;
output c320;
output c838;
output c9211;
output c094;
output c1456;
output c586;
output c2451;
output c2453;
output c2495;
output c50;
output c2363;
output c7393;
output c3473;
output c8438;
output c6492;
output c8108;
output c8433;
output c813;
output c7114;
output c118;
output c8127;
output c5246;
output c6318;
output c3278;
output c8291;
output c6331;
output c7152;
output c6122;
output c033;
output c1470;
output c2246;
output c4229;
output c528;
output c0498;
output c526;
output c5267;
output c8415;
output c8187;
output c4134;
output c8186;
output c8177;
output c2178;
output c2335;
output c4264;
output c9231;
output c8339;
output c965;
output c4306;
output c5287;
output c5259;
output c3137;
output c6215;
output c518;
output c7447;
output c268;
output c3138;
output c293;
output c1118;
output c4161;
output c8153;
output c6193;
output c6162;
output c9360;
output c1235;
output c5491;
output c4112;
output c7495;
output c5104;
output c5165;
output c08;
output c1333;
output c4325;
output c0457;
output c7314;
output c0218;
output c477;
output c6435;
output c7416;
output c010;
output c2126;
output c749;
output c9447;
output c5400;
output c4252;
output c048;
output c0409;
output c434;
output c7348;
output c1148;
output c6106;
output c7427;
output c821;
output c2183;
output c176;
output c6170;
output c7401;

assign c00 =  x41 & ~x118 & ~x487 & ~x490 & ~x589 & ~x609;
assign c02 =  x70 &  x603 &  x626 &  x627 &  x629 &  x683 &  x765 &  x769 &  x770 & ~x2 & ~x4 & ~x5 & ~x22 & ~x55 & ~x141 & ~x169 & ~x198 & ~x224 & ~x336 & ~x337 & ~x366 & ~x421 & ~x447 & ~x449 & ~x450 & ~x470 & ~x473 & ~x482 & ~x528 & ~x529 & ~x530 & ~x534 & ~x557 & ~x565 & ~x584 & ~x587 & ~x646 & ~x667 & ~x671 & ~x675 & ~x696 & ~x703 & ~x753;
assign c04 = ~x5 & ~x24 & ~x28 & ~x30 & ~x31 & ~x34 & ~x51 & ~x54 & ~x55 & ~x56 & ~x59 & ~x79 & ~x84 & ~x85 & ~x138 & ~x139 & ~x168 & ~x197 & ~x205 & ~x207 & ~x223 & ~x252 & ~x278 & ~x279 & ~x307 & ~x310 & ~x333 & ~x334 & ~x339 & ~x368 & ~x370 & ~x390 & ~x392 & ~x393 & ~x395 & ~x416 & ~x425 & ~x426 & ~x448 & ~x450 & ~x454 & ~x469 & ~x473 & ~x479 & ~x480 & ~x482 & ~x497 & ~x498 & ~x499 & ~x500 & ~x501 & ~x502 & ~x504 & ~x505 & ~x507 & ~x510 & ~x525 & ~x526 & ~x528 & ~x531 & ~x533 & ~x537 & ~x554 & ~x556 & ~x557 & ~x558 & ~x560 & ~x563 & ~x565 & ~x583 & ~x584 & ~x585 & ~x587 & ~x589 & ~x591 & ~x613 & ~x614 & ~x616 & ~x617 & ~x621 & ~x638 & ~x641 & ~x646 & ~x647 & ~x667 & ~x669 & ~x670 & ~x673 & ~x674 & ~x676 & ~x698 & ~x723 & ~x727 & ~x728 & ~x729 & ~x752 & ~x754 & ~x757 & ~x759 & ~x761 & ~x778 & ~x781 & ~x783;
assign c06 = ~x336 & ~x344 & ~x372 & ~x520 & ~x632 & ~x658 & ~x732;
assign c08 =  x40 &  x41 &  x42 &  x44 & ~x2 & ~x4 & ~x5 & ~x7 & ~x13 & ~x14 & ~x25 & ~x28 & ~x31 & ~x33 & ~x58 & ~x80 & ~x112 & ~x115 & ~x140 & ~x168 & ~x195 & ~x223 & ~x332 & ~x334 & ~x338 & ~x361 & ~x363 & ~x365 & ~x367 & ~x393 & ~x417 & ~x427 & ~x455 & ~x470 & ~x476 & ~x478 & ~x481 & ~x503 & ~x532 & ~x557 & ~x560 & ~x561 & ~x563 & ~x565 & ~x566 & ~x584 & ~x588 & ~x591 & ~x594 & ~x614 & ~x615 & ~x617 & ~x622 & ~x644 & ~x645 & ~x646 & ~x650 & ~x668 & ~x670 & ~x674 & ~x676 & ~x678 & ~x695 & ~x702 & ~x703 & ~x704 & ~x724 & ~x734 & ~x752 & ~x756 & ~x757 & ~x761 & ~x762;
assign c010 = ~x279 & ~x363 & ~x417 & ~x419 & ~x445 & ~x455 & ~x483 & ~x594 & ~x709 & ~x710 & ~x711 & ~x713 & ~x750 & ~x751;
assign c012 =  x42 &  x285 &  x736 & ~x3 & ~x20 & ~x21 & ~x23 & ~x24 & ~x26 & ~x52 & ~x57 & ~x59 & ~x81 & ~x82 & ~x83 & ~x84 & ~x86 & ~x114 & ~x169 & ~x279 & ~x306 & ~x308 & ~x335 & ~x389 & ~x394 & ~x395 & ~x422 & ~x450 & ~x476 & ~x477 & ~x504 & ~x505 & ~x506 & ~x530 & ~x533 & ~x560 & ~x561 & ~x562 & ~x586 & ~x614 & ~x642 & ~x667 & ~x673 & ~x674 & ~x695 & ~x697 & ~x700 & ~x703 & ~x723 & ~x724 & ~x725 & ~x755 & ~x756 & ~x757 & ~x759 & ~x779 & ~x781;
assign c014 =  x711 & ~x1 & ~x25 & ~x29 & ~x30 & ~x32 & ~x52 & ~x54 & ~x84 & ~x167 & ~x168 & ~x279 & ~x308 & ~x364 & ~x494 & ~x501 & ~x502 & ~x529 & ~x530 & ~x558 & ~x559 & ~x588 & ~x589 & ~x591 & ~x614 & ~x615 & ~x671 & ~x672 & ~x727 & ~x728 & ~x729 & ~x782;
assign c016 =  x565 &  x707 &  x713 & ~x32 & ~x723 & ~x726 & ~x751;
assign c018 =  x227 &  x255;
assign c020 =  x432 & ~x1 & ~x5 & ~x9 & ~x55 & ~x81 & ~x96 & ~x111 & ~x137 & ~x138 & ~x251 & ~x448 & ~x478 & ~x507 & ~x528 & ~x557 & ~x558 & ~x613 & ~x616 & ~x618 & ~x644 & ~x674 & ~x759;
assign c022 =  x430 & ~x0 & ~x1 & ~x3 & ~x11 & ~x12 & ~x13 & ~x14 & ~x15 & ~x16 & ~x17 & ~x23 & ~x25 & ~x26 & ~x28 & ~x29 & ~x30 & ~x41 & ~x42 & ~x53 & ~x54 & ~x55 & ~x57 & ~x58 & ~x81 & ~x83 & ~x84 & ~x85 & ~x86 & ~x110 & ~x111 & ~x113 & ~x114 & ~x136 & ~x137 & ~x138 & ~x139 & ~x140 & ~x141 & ~x166 & ~x167 & ~x168 & ~x197 & ~x198 & ~x224 & ~x225 & ~x250 & ~x279 & ~x282 & ~x307 & ~x309 & ~x310 & ~x333 & ~x335 & ~x336 & ~x337 & ~x361 & ~x363 & ~x364 & ~x390 & ~x391 & ~x393 & ~x418 & ~x420 & ~x421 & ~x446 & ~x447 & ~x448 & ~x451 & ~x474 & ~x475 & ~x476 & ~x477 & ~x478 & ~x502 & ~x503 & ~x504 & ~x505 & ~x506 & ~x531 & ~x532 & ~x558 & ~x559 & ~x560 & ~x586 & ~x587 & ~x588 & ~x589 & ~x590 & ~x616 & ~x617 & ~x618 & ~x642 & ~x643 & ~x644 & ~x645 & ~x671 & ~x674 & ~x700 & ~x702 & ~x726 & ~x727 & ~x728 & ~x729 & ~x757 & ~x758 & ~x759 & ~x782;
assign c024 = ~x1 & ~x32 & ~x126 & ~x128 & ~x424 & ~x441 & ~x443 & ~x454 & ~x469 & ~x470 & ~x482 & ~x498 & ~x510 & ~x528 & ~x553 & ~x593 & ~x641 & ~x749;
assign c026 =  x274 &  x571 &  x576 & ~x1 & ~x4 & ~x7 & ~x8 & ~x20 & ~x22 & ~x24 & ~x26 & ~x27 & ~x29 & ~x31 & ~x32 & ~x33 & ~x58 & ~x60 & ~x82 & ~x86 & ~x87 & ~x109 & ~x115 & ~x137 & ~x166 & ~x168 & ~x169 & ~x194 & ~x197 & ~x198 & ~x221 & ~x223 & ~x225 & ~x250 & ~x253 & ~x305 & ~x308 & ~x336 & ~x362 & ~x363 & ~x365 & ~x391 & ~x394 & ~x418 & ~x422 & ~x423 & ~x450 & ~x451 & ~x474 & ~x477 & ~x478 & ~x504 & ~x505 & ~x507 & ~x530 & ~x532 & ~x533 & ~x558 & ~x561 & ~x562 & ~x591 & ~x594 & ~x612 & ~x616 & ~x620 & ~x621 & ~x648 & ~x649 & ~x667 & ~x668 & ~x698 & ~x701 & ~x703 & ~x705 & ~x706 & ~x723 & ~x726 & ~x728 & ~x729 & ~x730 & ~x731 & ~x733 & ~x734 & ~x750 & ~x751 & ~x754 & ~x779;
assign c028 = ~x5 & ~x14 & ~x24 & ~x94 & ~x124 & ~x125 & ~x127 & ~x335 & ~x478 & ~x481 & ~x501 & ~x528 & ~x534 & ~x537 & ~x554 & ~x556 & ~x584 & ~x586 & ~x593 & ~x640 & ~x644 & ~x649 & ~x669 & ~x674 & ~x697 & ~x701 & ~x704 & ~x726 & ~x752 & ~x761 & ~x762;
assign c030 =  x70 &  x520 &  x573 &  x628 &  x629 &  x659 & ~x4 & ~x9 & ~x21 & ~x27 & ~x29 & ~x50 & ~x53 & ~x56 & ~x57 & ~x112 & ~x139 & ~x143 & ~x169 & ~x195 & ~x223 & ~x228 & ~x249 & ~x250 & ~x308 & ~x368 & ~x384 & ~x390 & ~x395 & ~x444 & ~x447 & ~x475 & ~x480 & ~x502 & ~x506 & ~x526 & ~x527 & ~x563 & ~x586 & ~x609 & ~x613 & ~x614 & ~x619 & ~x639 & ~x644 & ~x646 & ~x668 & ~x693 & ~x694 & ~x696 & ~x749 & ~x752 & ~x754 & ~x757 & ~x783;
assign c032 =  x94 &  x126 &  x215 &  x238 &  x293 &  x317 &  x355 &  x405 &  x576 &  x601 &  x686 &  x690 &  x719 &  x747 & ~x6 & ~x113 & ~x116 & ~x226 & ~x246 & ~x309 & ~x394 & ~x450 & ~x477 & ~x480 & ~x536 & ~x555 & ~x589 & ~x613 & ~x616 & ~x617;
assign c034 = ~x58 & ~x109 & ~x113 & ~x135 & ~x390 & ~x398 & ~x416 & ~x441 & ~x446 & ~x450 & ~x455 & ~x468 & ~x503 & ~x525 & ~x538 & ~x558 & ~x584 & ~x611 & ~x642 & ~x669 & ~x695 & ~x706 & ~x708 & ~x723 & ~x733 & ~x750 & ~x763 & ~x766 & ~x767 & ~x772 & ~x773 & ~x776 & ~x779;
assign c036 =  x539 &  x595 & ~x12 & ~x14 & ~x15 & ~x68 & ~x84 & ~x309 & ~x334 & ~x757 & ~x783;
assign c038 =  x209 &  x237 &  x266 &  x269 &  x289 &  x290 &  x317 &  x464 &  x513 &  x630 &  x686 &  x712 &  x713 &  x769 & ~x55 & ~x57 & ~x135 & ~x139 & ~x169 & ~x202 & ~x229 & ~x247 & ~x443 & ~x474 & ~x530 & ~x560 & ~x644 & ~x646;
assign c040 =  x77 &  x78 & ~x0 & ~x54 & ~x223 & ~x280 & ~x309 & ~x365 & ~x391 & ~x422 & ~x616 & ~x640 & ~x642 & ~x669 & ~x702 & ~x756 & ~x783;
assign c042 = ~x343 & ~x389 & ~x419 & ~x445 & ~x473 & ~x594 & ~x608 & ~x655 & ~x678;
assign c044 =  x41 &  x42 &  x43 &  x258 & ~x4 & ~x6 & ~x7 & ~x8 & ~x22 & ~x23 & ~x31 & ~x32 & ~x33 & ~x51 & ~x53 & ~x55 & ~x58 & ~x60 & ~x81 & ~x114 & ~x115 & ~x136 & ~x139 & ~x141 & ~x142 & ~x169 & ~x170 & ~x194 & ~x196 & ~x223 & ~x250 & ~x251 & ~x309 & ~x363 & ~x398 & ~x414 & ~x418 & ~x420 & ~x424 & ~x426 & ~x444 & ~x448 & ~x450 & ~x471 & ~x473 & ~x474 & ~x477 & ~x480 & ~x481 & ~x482 & ~x503 & ~x507 & ~x510 & ~x526 & ~x530 & ~x531 & ~x534 & ~x535 & ~x538 & ~x554 & ~x555 & ~x556 & ~x557 & ~x561 & ~x562 & ~x563 & ~x585 & ~x587 & ~x588 & ~x589 & ~x592 & ~x610 & ~x612 & ~x613 & ~x614 & ~x615 & ~x616 & ~x617 & ~x621 & ~x622 & ~x638 & ~x639 & ~x644 & ~x646 & ~x647 & ~x648 & ~x649 & ~x650 & ~x669 & ~x670 & ~x671 & ~x677 & ~x694 & ~x695 & ~x696 & ~x699 & ~x701 & ~x702 & ~x703 & ~x704 & ~x705 & ~x706 & ~x722 & ~x723 & ~x725 & ~x727 & ~x730 & ~x731 & ~x752 & ~x753 & ~x755 & ~x757 & ~x760 & ~x761 & ~x778 & ~x780 & ~x781 & ~x782;
assign c046 =  x94 &  x123 &  x157 &  x378 & ~x8 & ~x21 & ~x34 & ~x51 & ~x52 & ~x54 & ~x61 & ~x81 & ~x114 & ~x139 & ~x141 & ~x195 & ~x245 & ~x255 & ~x284 & ~x306 & ~x315 & ~x333 & ~x363 & ~x364 & ~x365 & ~x371 & ~x389 & ~x413 & ~x447 & ~x449 & ~x473 & ~x536 & ~x589 & ~x615 & ~x616 & ~x697 & ~x725 & ~x726 & ~x728 & ~x733 & ~x750 & ~x783;
assign c048 = ~x14 & ~x404 & ~x461 & ~x502 & ~x508 & ~x529 & ~x558 & ~x583 & ~x593 & ~x698 & ~x704 & ~x723 & ~x732;
assign c050 = ~x1 & ~x10 & ~x11 & ~x15 & ~x19 & ~x28 & ~x39 & ~x40 & ~x41 & ~x44 & ~x56 & ~x57 & ~x84 & ~x112 & ~x137 & ~x139 & ~x140 & ~x167 & ~x335 & ~x475 & ~x502 & ~x529 & ~x559 & ~x560 & ~x729 & ~x731 & ~x757;
assign c052 =  x206 &  x325 &  x406 &  x518 &  x573 &  x598 & ~x28 & ~x91 & ~x119 & ~x146 & ~x175 & ~x255 & ~x310 & ~x385 & ~x394 & ~x442 & ~x503 & ~x586 & ~x673 & ~x753;
assign c054 = ~x384 & ~x418 & ~x435 & ~x440 & ~x447 & ~x494 & ~x501 & ~x582 & ~x733;
assign c056 =  x49 & ~x1 & ~x25 & ~x113 & ~x415 & ~x534 & ~x564 & ~x612 & ~x676 & ~x696 & ~x698 & ~x725 & ~x729;
assign c058 =  x64 & ~x3 & ~x4 & ~x6 & ~x23 & ~x24 & ~x26 & ~x29 & ~x30 & ~x54 & ~x55 & ~x85 & ~x141 & ~x168 & ~x196 & ~x222 & ~x224 & ~x279 & ~x281 & ~x336 & ~x363 & ~x419 & ~x448 & ~x476 & ~x522 & ~x531 & ~x671 & ~x757 & ~x759 & ~x779 & ~x780;
assign c060 =  x63 & ~x4 & ~x22 & ~x23 & ~x27 & ~x34 & ~x54 & ~x55 & ~x112 & ~x194 & ~x223 & ~x253 & ~x254 & ~x339 & ~x360 & ~x361 & ~x363 & ~x364 & ~x370 & ~x389 & ~x395 & ~x426 & ~x445 & ~x453 & ~x532 & ~x537 & ~x559 & ~x560 & ~x562 & ~x584 & ~x586 & ~x612 & ~x615 & ~x616 & ~x668 & ~x671 & ~x672 & ~x696 & ~x697 & ~x701 & ~x704 & ~x732 & ~x760;
assign c062 =  x567 &  x568 &  x596 &  x651 &  x652 &  x654 &  x657 &  x678 &  x679 &  x680 &  x706 &  x707 &  x708 &  x714 &  x736 & ~x11 & ~x13 & ~x14 & ~x15 & ~x16 & ~x25 & ~x54 & ~x82 & ~x334 & ~x587 & ~x616 & ~x757;
assign c064 =  x125 &  x130 &  x157 &  x158 &  x214 &  x240 &  x289 &  x320 &  x321 &  x345 &  x349 &  x433 &  x437 &  x461 &  x462 &  x465 &  x488 &  x492 &  x516 &  x517 &  x518 &  x520 &  x549 &  x569 &  x572 &  x578 &  x600 &  x602 &  x603 &  x605 &  x606 &  x625 &  x629 &  x632 &  x656 &  x659 &  x660 & ~x23 & ~x29 & ~x30 & ~x50 & ~x80 & ~x113 & ~x115 & ~x140 & ~x164 & ~x165 & ~x170 & ~x197 & ~x222 & ~x249 & ~x250 & ~x278 & ~x284 & ~x304 & ~x305 & ~x337 & ~x360 & ~x385 & ~x394 & ~x413 & ~x424 & ~x446 & ~x447 & ~x470 & ~x476 & ~x478 & ~x503 & ~x538 & ~x553 & ~x558 & ~x561 & ~x582 & ~x590 & ~x591 & ~x611 & ~x640 & ~x641 & ~x642 & ~x644 & ~x645 & ~x646 & ~x668 & ~x696 & ~x723 & ~x753 & ~x754 & ~x757 & ~x761 & ~x780;
assign c066 = ~x371 & ~x418 & ~x473 & ~x483 & ~x705 & ~x709 & ~x710 & ~x711 & ~x729 & ~x741;
assign c068 =  x130 &  x157 &  x270 &  x298 &  x488 &  x568 &  x575 &  x603 & ~x6 & ~x22 & ~x28 & ~x51 & ~x52 & ~x54 & ~x59 & ~x79 & ~x86 & ~x110 & ~x114 & ~x165 & ~x223 & ~x227 & ~x248 & ~x304 & ~x305 & ~x309 & ~x333 & ~x336 & ~x361 & ~x362 & ~x390 & ~x393 & ~x419 & ~x440 & ~x446 & ~x468 & ~x475 & ~x476 & ~x477 & ~x506 & ~x530 & ~x558 & ~x561 & ~x589 & ~x621 & ~x642 & ~x643 & ~x644 & ~x647 & ~x674 & ~x675 & ~x677 & ~x700 & ~x702 & ~x703 & ~x705 & ~x722 & ~x723 & ~x729 & ~x732 & ~x752 & ~x756 & ~x759 & ~x779 & ~x780 & ~x781;
assign c070 =  x143;
assign c072 =  x227 & ~x22 & ~x27 & ~x83 & ~x224 & ~x307 & ~x588 & ~x616 & ~x759 & ~x782 & ~x783;
assign c074 =  x133 &  x146 &  x188 &  x573 &  x607 & ~x3 & ~x24 & ~x82 & ~x86 & ~x108 & ~x141 & ~x143 & ~x170 & ~x335 & ~x337 & ~x419 & ~x447 & ~x449 & ~x455 & ~x697 & ~x703 & ~x723 & ~x724 & ~x758 & ~x760 & ~x781;
assign c076 =  x271 &  x413 &  x574 &  x682 &  x690 &  x747 &  x749 & ~x366 & ~x394 & ~x506 & ~x671 & ~x757;
assign c078 = ~x0 & ~x2 & ~x5 & ~x7 & ~x8 & ~x22 & ~x23 & ~x25 & ~x26 & ~x27 & ~x29 & ~x31 & ~x55 & ~x58 & ~x59 & ~x60 & ~x84 & ~x85 & ~x108 & ~x112 & ~x113 & ~x137 & ~x142 & ~x143 & ~x166 & ~x168 & ~x169 & ~x170 & ~x193 & ~x194 & ~x196 & ~x197 & ~x221 & ~x223 & ~x224 & ~x225 & ~x252 & ~x279 & ~x280 & ~x307 & ~x308 & ~x336 & ~x337 & ~x350 & ~x363 & ~x365 & ~x366 & ~x389 & ~x392 & ~x395 & ~x417 & ~x419 & ~x421 & ~x426 & ~x441 & ~x446 & ~x447 & ~x469 & ~x475 & ~x476 & ~x477 & ~x482 & ~x505 & ~x510 & ~x526 & ~x527 & ~x533 & ~x536 & ~x558 & ~x561 & ~x563 & ~x584 & ~x588 & ~x589 & ~x590 & ~x593 & ~x610 & ~x612 & ~x614 & ~x615 & ~x618 & ~x619 & ~x620 & ~x638 & ~x644 & ~x646 & ~x649 & ~x650 & ~x666 & ~x668 & ~x669 & ~x670 & ~x671 & ~x672 & ~x673 & ~x674 & ~x678 & ~x695 & ~x698 & ~x700 & ~x702 & ~x704 & ~x706 & ~x728 & ~x729 & ~x730 & ~x732 & ~x734 & ~x750 & ~x751 & ~x753 & ~x754 & ~x756 & ~x758 & ~x760 & ~x762 & ~x777 & ~x778 & ~x779 & ~x782;
assign c080 =  x133 & ~x7 & ~x25 & ~x33 & ~x35 & ~x55 & ~x61 & ~x87 & ~x138 & ~x169 & ~x198 & ~x223 & ~x224 & ~x251 & ~x252 & ~x306 & ~x337 & ~x422 & ~x423 & ~x446 & ~x475 & ~x479 & ~x502 & ~x530 & ~x533 & ~x560 & ~x564 & ~x582 & ~x591 & ~x610 & ~x614 & ~x640 & ~x644 & ~x668 & ~x673 & ~x697 & ~x704 & ~x723 & ~x729 & ~x751 & ~x756 & ~x761 & ~x762 & ~x777 & ~x779;
assign c082 =  x270 &  x465 &  x603 &  x606 &  x625 &  x658 &  x681 &  x684 &  x691 &  x742 &  x766 &  x767 &  x769 &  x770 &  x771 &  x773 & ~x2 & ~x80 & ~x114 & ~x138 & ~x139 & ~x196 & ~x224 & ~x225 & ~x278 & ~x279 & ~x282 & ~x283 & ~x365 & ~x389 & ~x397 & ~x414 & ~x418 & ~x442 & ~x447 & ~x476 & ~x480 & ~x504 & ~x508 & ~x526 & ~x561 & ~x565 & ~x583 & ~x585 & ~x588 & ~x591 & ~x618 & ~x639 & ~x640 & ~x648 & ~x673 & ~x677 & ~x703 & ~x731 & ~x732 & ~x760 & ~x780;
assign c084 =  x290 &  x549 &  x599 &  x603 &  x625 & ~x9 & ~x36 & ~x141 & ~x280 & ~x391 & ~x555 & ~x679 & ~x700;
assign c086 =  x289 &  x317 &  x570 &  x712 &  x736 & ~x0 & ~x1 & ~x8 & ~x9 & ~x21 & ~x27 & ~x35 & ~x36 & ~x54 & ~x56 & ~x80 & ~x81 & ~x85 & ~x88 & ~x113 & ~x143 & ~x281 & ~x282 & ~x309 & ~x337 & ~x359 & ~x362 & ~x389 & ~x394 & ~x415 & ~x417 & ~x419 & ~x420 & ~x446 & ~x450 & ~x451 & ~x470 & ~x471 & ~x475 & ~x479 & ~x498 & ~x499 & ~x503 & ~x504 & ~x528 & ~x534 & ~x562 & ~x586 & ~x590 & ~x615 & ~x639 & ~x640 & ~x644 & ~x669 & ~x696 & ~x700 & ~x703 & ~x704 & ~x752 & ~x754 & ~x761 & ~x783;
assign c088 =  x490 &  x770 & ~x147 & ~x371 & ~x619 & ~x752 & ~x759 & ~x780;
assign c090 = ~x456 & ~x583 & ~x593 & ~x610 & ~x646 & ~x710 & ~x721 & ~x737 & ~x751 & ~x772;
assign c092 =  x198;
assign c094 =  x325 & ~x334 & ~x362 & ~x416 & ~x734 & ~x738 & ~x762;
assign c096 =  x90 &  x94 &  x97 &  x147 &  x158 &  x177 &  x548 &  x689 & ~x22 & ~x52 & ~x55 & ~x82 & ~x85 & ~x168 & ~x196 & ~x393 & ~x448 & ~x531 & ~x560 & ~x594 & ~x645 & ~x648 & ~x673 & ~x676 & ~x754 & ~x755 & ~x757 & ~x759;
assign c098 =  x310 &  x311 & ~x29;
assign c0100 =  x339 & ~x29 & ~x49 & ~x137 & ~x139 & ~x559 & ~x643 & ~x759;
assign c0102 =  x204 &  x232 &  x322 &  x457 &  x542 &  x599 &  x624 &  x686 &  x738 &  x742 &  x763 & ~x83 & ~x505 & ~x783;
assign c0104 =  x107 & ~x168 & ~x252 & ~x395 & ~x477 & ~x560 & ~x590 & ~x614 & ~x642 & ~x669 & ~x703 & ~x758;
assign c0106 =  x123 &  x128 &  x424 & ~x22 & ~x26 & ~x110 & ~x138 & ~x141 & ~x142 & ~x166 & ~x223 & ~x224 & ~x225 & ~x250 & ~x251 & ~x280 & ~x559 & ~x757 & ~x758 & ~x779;
assign c0108 =  x77 &  x228 & ~x56 & ~x82 & ~x112 & ~x223 & ~x224 & ~x307 & ~x482 & ~x732;
assign c0110 = ~x50 & ~x128 & ~x277 & ~x306 & ~x334 & ~x338 & ~x362 & ~x390 & ~x393 & ~x440 & ~x441 & ~x443 & ~x444 & ~x449 & ~x454 & ~x468 & ~x501 & ~x502 & ~x529 & ~x530 & ~x555 & ~x557 & ~x566 & ~x608 & ~x609 & ~x636 & ~x642 & ~x666 & ~x673 & ~x721 & ~x750 & ~x756 & ~x761;
assign c0112 =  x16 &  x76 &  x124 & ~x5 & ~x307;
assign c0114 =  x40 &  x768 &  x769 &  x771 & ~x0 & ~x3 & ~x4 & ~x5 & ~x7 & ~x8 & ~x27 & ~x29 & ~x53 & ~x57 & ~x58 & ~x79 & ~x81 & ~x83 & ~x108 & ~x111 & ~x120 & ~x140 & ~x141 & ~x166 & ~x193 & ~x197 & ~x198 & ~x222 & ~x223 & ~x225 & ~x249 & ~x251 & ~x278 & ~x308 & ~x339 & ~x362 & ~x365 & ~x415 & ~x425 & ~x444 & ~x445 & ~x472 & ~x474 & ~x475 & ~x476 & ~x477 & ~x480 & ~x481 & ~x500 & ~x509 & ~x510 & ~x528 & ~x530 & ~x532 & ~x533 & ~x534 & ~x535 & ~x536 & ~x554 & ~x558 & ~x565 & ~x566 & ~x582 & ~x584 & ~x585 & ~x586 & ~x587 & ~x588 & ~x589 & ~x593 & ~x611 & ~x618 & ~x620 & ~x621 & ~x638 & ~x639 & ~x641 & ~x645 & ~x670 & ~x674 & ~x675 & ~x676 & ~x695 & ~x697 & ~x699 & ~x704 & ~x723 & ~x726 & ~x727 & ~x731 & ~x733 & ~x750 & ~x751 & ~x755 & ~x780 & ~x782 & ~x783;
assign c0116 =  x79;
assign c0118 =  x98 &  x155 &  x312 &  x460 &  x515 &  x547 &  x598 &  x601 &  x682 &  x715 & ~x3 & ~x54 & ~x60 & ~x254 & ~x419 & ~x559 & ~x704;
assign c0120 =  x71 &  x461 &  x630 & ~x0 & ~x85 & ~x133 & ~x196 & ~x249 & ~x362 & ~x399 & ~x419 & ~x446 & ~x449 & ~x455 & ~x530 & ~x536 & ~x582 & ~x593 & ~x614 & ~x618 & ~x640 & ~x650 & ~x706;
assign c0122 =  x542 &  x551 &  x579 &  x662 &  x712 &  x714 &  x748 &  x749 & ~x10 & ~x14 & ~x195 & ~x252 & ~x334 & ~x392 & ~x587 & ~x588 & ~x757 & ~x758;
assign c0124 =  x144 & ~x6 & ~x25 & ~x26 & ~x27 & ~x29 & ~x51 & ~x56 & ~x85 & ~x141 & ~x309 & ~x450 & ~x476 & ~x589 & ~x642 & ~x702 & ~x731 & ~x757 & ~x759;
assign c0126 = ~x2 & ~x4 & ~x13 & ~x14 & ~x15 & ~x27 & ~x59 & ~x73 & ~x80 & ~x86 & ~x87 & ~x96 & ~x109 & ~x112 & ~x137 & ~x141 & ~x166 & ~x168 & ~x196 & ~x197 & ~x222 & ~x251 & ~x253 & ~x278 & ~x279 & ~x307 & ~x308 & ~x446 & ~x472 & ~x478 & ~x500 & ~x501 & ~x502 & ~x504 & ~x506 & ~x530 & ~x532 & ~x535 & ~x536 & ~x556 & ~x558 & ~x560 & ~x561 & ~x562 & ~x584 & ~x586 & ~x589 & ~x614 & ~x615 & ~x617 & ~x618 & ~x619 & ~x641 & ~x644 & ~x646 & ~x669 & ~x670 & ~x671 & ~x673 & ~x674 & ~x675 & ~x698 & ~x701 & ~x731 & ~x759 & ~x783;
assign c0128 =  x204 &  x409 &  x545 &  x741 & ~x27 & ~x55 & ~x56 & ~x62 & ~x106 & ~x163 & ~x201 & ~x229 & ~x256 & ~x307 & ~x421 & ~x561 & ~x584 & ~x588 & ~x615 & ~x616 & ~x641 & ~x642 & ~x670 & ~x672 & ~x781;
assign c0130 =  x177 &  x233 &  x289 &  x298 &  x402 &  x429 &  x571 &  x573 &  x575 &  x596 &  x600 &  x603 & ~x24 & ~x29 & ~x162 & ~x168 & ~x225 & ~x278 & ~x399 & ~x527 & ~x559 & ~x565 & ~x585 & ~x640 & ~x647 & ~x649 & ~x780 & ~x782;
assign c0132 =  x351 & ~x180 & ~x309 & ~x364 & ~x385 & ~x413 & ~x441 & ~x442 & ~x469 & ~x470 & ~x498 & ~x505 & ~x527 & ~x583 & ~x672 & ~x675 & ~x703 & ~x781;
assign c0134 = ~x2 & ~x7 & ~x30 & ~x84 & ~x85 & ~x86 & ~x104 & ~x113 & ~x114 & ~x132 & ~x133 & ~x140 & ~x156 & ~x157 & ~x160 & ~x166 & ~x225 & ~x226 & ~x306 & ~x307 & ~x311 & ~x334 & ~x336 & ~x337 & ~x366 & ~x390 & ~x396 & ~x398 & ~x415 & ~x416 & ~x423 & ~x425 & ~x441 & ~x445 & ~x450 & ~x451 & ~x454 & ~x469 & ~x471 & ~x474 & ~x476 & ~x497 & ~x509 & ~x525 & ~x531 & ~x555 & ~x561 & ~x582 & ~x583 & ~x591 & ~x593 & ~x611 & ~x638 & ~x646 & ~x647 & ~x648 & ~x649 & ~x669 & ~x670 & ~x671 & ~x677 & ~x700 & ~x704 & ~x705 & ~x726 & ~x728 & ~x753 & ~x778 & ~x781 & ~x782;
assign c0136 =  x233 &  x263 &  x267 &  x270 &  x289 &  x297 &  x457 &  x488 &  x493 &  x545 &  x548 &  x570 &  x572 &  x577 &  x578 &  x596 &  x603 &  x624 &  x625 &  x629 &  x630 &  x657 &  x661 &  x662 &  x681 & ~x2 & ~x4 & ~x5 & ~x29 & ~x55 & ~x56 & ~x63 & ~x83 & ~x85 & ~x87 & ~x109 & ~x140 & ~x144 & ~x165 & ~x171 & ~x191 & ~x198 & ~x200 & ~x248 & ~x249 & ~x252 & ~x254 & ~x277 & ~x280 & ~x282 & ~x305 & ~x306 & ~x363 & ~x388 & ~x419 & ~x420 & ~x447 & ~x472 & ~x507 & ~x508 & ~x530 & ~x531 & ~x534 & ~x583 & ~x586 & ~x592 & ~x611 & ~x612 & ~x614 & ~x616 & ~x619 & ~x648 & ~x668 & ~x677 & ~x699 & ~x701 & ~x704 & ~x728 & ~x732 & ~x761 & ~x780;
assign c0138 =  x282;
assign c0140 = ~x22 & ~x252 & ~x392 & ~x418 & ~x445 & ~x448 & ~x473 & ~x477 & ~x500 & ~x529 & ~x532 & ~x535 & ~x558 & ~x563 & ~x583 & ~x612 & ~x618 & ~x621 & ~x640 & ~x667 & ~x670 & ~x696 & ~x701 & ~x704 & ~x706 & ~x709 & ~x710 & ~x713 & ~x720 & ~x722 & ~x752 & ~x762;
assign c0142 = ~x0 & ~x2 & ~x170 & ~x178 & ~x180 & ~x194 & ~x339 & ~x361 & ~x413 & ~x416 & ~x418 & ~x442 & ~x443 & ~x446 & ~x473 & ~x477 & ~x498 & ~x502 & ~x510 & ~x528 & ~x538 & ~x564 & ~x566 & ~x583 & ~x612 & ~x616 & ~x619 & ~x641 & ~x645 & ~x667 & ~x670 & ~x671 & ~x699 & ~x706 & ~x725 & ~x751 & ~x756 & ~x762;
assign c0144 =  x76 &  x105 &  x232 &  x573 &  x604 &  x626 &  x627 &  x628 &  x654 &  x655 &  x684 & ~x6 & ~x28 & ~x84 & ~x335 & ~x365 & ~x390 & ~x423 & ~x448 & ~x451 & ~x477 & ~x531 & ~x619 & ~x621 & ~x639 & ~x667 & ~x671 & ~x696 & ~x698 & ~x702 & ~x728 & ~x733 & ~x734 & ~x752;
assign c0146 = ~x25 & ~x95 & ~x126 & ~x333 & ~x481 & ~x483 & ~x530 & ~x554 & ~x566 & ~x668 & ~x695 & ~x750 & ~x752;
assign c0148 = ~x300 & ~x390 & ~x492 & ~x705 & ~x723 & ~x733 & ~x750;
assign c0150 =  x91 &  x443;
assign c0152 = ~x102 & ~x198 & ~x333 & ~x412 & ~x415 & ~x419 & ~x421 & ~x446 & ~x469 & ~x470 & ~x498 & ~x506 & ~x510 & ~x551 & ~x552 & ~x676 & ~x723 & ~x732 & ~x750 & ~x751;
assign c0154 =  x144 &  x255 & ~x84 & ~x168 & ~x280 & ~x364 & ~x643;
assign c0156 =  x212 &  x270 &  x298 &  x462 &  x572 &  x629 &  x630 & ~x2 & ~x21 & ~x23 & ~x59 & ~x110 & ~x136 & ~x138 & ~x142 & ~x198 & ~x221 & ~x312 & ~x328 & ~x360 & ~x361 & ~x384 & ~x392 & ~x394 & ~x445 & ~x451 & ~x496 & ~x506 & ~x530 & ~x555 & ~x559 & ~x560 & ~x590 & ~x591 & ~x613 & ~x615 & ~x640 & ~x642 & ~x666 & ~x667 & ~x675 & ~x725 & ~x726 & ~x727 & ~x756 & ~x757 & ~x777;
assign c0158 =  x42 &  x128 &  x201 &  x258 & ~x0 & ~x3 & ~x52 & ~x61 & ~x82 & ~x111 & ~x165 & ~x279 & ~x503 & ~x588 & ~x676 & ~x677 & ~x705 & ~x732 & ~x755;
assign c0160 =  x78 & ~x1 & ~x5 & ~x23 & ~x56 & ~x82 & ~x111 & ~x195 & ~x196 & ~x279 & ~x336 & ~x360 & ~x362 & ~x366 & ~x367 & ~x391 & ~x393 & ~x419 & ~x421 & ~x447 & ~x501 & ~x503 & ~x530 & ~x531 & ~x617 & ~x645 & ~x674 & ~x699 & ~x700 & ~x702 & ~x724 & ~x727 & ~x728 & ~x754 & ~x755 & ~x758;
assign c0162 =  x510 &  x708 &  x735 &  x739 & ~x0 & ~x12 & ~x13 & ~x15;
assign c0164 =  x270 &  x437 & ~x165 & ~x393 & ~x414 & ~x421 & ~x445 & ~x526 & ~x645 & ~x646 & ~x673 & ~x772 & ~x773 & ~x779;
assign c0166 =  x203 & ~x1 & ~x2 & ~x3 & ~x5 & ~x10 & ~x23 & ~x24 & ~x25 & ~x26 & ~x27 & ~x28 & ~x29 & ~x32 & ~x51 & ~x52 & ~x54 & ~x55 & ~x56 & ~x57 & ~x59 & ~x79 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x108 & ~x110 & ~x111 & ~x112 & ~x138 & ~x139 & ~x141 & ~x164 & ~x167 & ~x168 & ~x169 & ~x194 & ~x196 & ~x197 & ~x198 & ~x223 & ~x225 & ~x226 & ~x251 & ~x252 & ~x253 & ~x279 & ~x280 & ~x281 & ~x282 & ~x304 & ~x305 & ~x306 & ~x307 & ~x308 & ~x309 & ~x332 & ~x333 & ~x335 & ~x336 & ~x338 & ~x361 & ~x362 & ~x364 & ~x365 & ~x366 & ~x389 & ~x390 & ~x391 & ~x392 & ~x393 & ~x395 & ~x418 & ~x419 & ~x420 & ~x421 & ~x422 & ~x445 & ~x447 & ~x448 & ~x449 & ~x473 & ~x474 & ~x475 & ~x476 & ~x477 & ~x478 & ~x501 & ~x502 & ~x503 & ~x504 & ~x524 & ~x532 & ~x558 & ~x559 & ~x560 & ~x586 & ~x587 & ~x588 & ~x613 & ~x615 & ~x617 & ~x618 & ~x643 & ~x646 & ~x668 & ~x671 & ~x672 & ~x673 & ~x695 & ~x696 & ~x697 & ~x698 & ~x699 & ~x701 & ~x703 & ~x723 & ~x724 & ~x725 & ~x726 & ~x729 & ~x730 & ~x731 & ~x751 & ~x753 & ~x755 & ~x756 & ~x758 & ~x777 & ~x779 & ~x781 & ~x782 & ~x783;
assign c0168 =  x396 &  x537 & ~x10 & ~x336 & ~x391 & ~x588;
assign c0170 =  x233 &  x265 &  x298 &  x318 &  x380 &  x406 &  x463 &  x607 & ~x7 & ~x21 & ~x24 & ~x29 & ~x33 & ~x51 & ~x58 & ~x83 & ~x108 & ~x109 & ~x136 & ~x138 & ~x140 & ~x197 & ~x226 & ~x249 & ~x254 & ~x279 & ~x308 & ~x313 & ~x329 & ~x332 & ~x360 & ~x365 & ~x371 & ~x386 & ~x392 & ~x393 & ~x399 & ~x413 & ~x414 & ~x447 & ~x452 & ~x473 & ~x474 & ~x476 & ~x480 & ~x497 & ~x500 & ~x501 & ~x502 & ~x503 & ~x507 & ~x525 & ~x529 & ~x532 & ~x533 & ~x534 & ~x554 & ~x561 & ~x562 & ~x586 & ~x594 & ~x612 & ~x614 & ~x617 & ~x622 & ~x639 & ~x667 & ~x671 & ~x675 & ~x677 & ~x695 & ~x706 & ~x726 & ~x752 & ~x757 & ~x759 & ~x783;
assign c0172 =  x115;
assign c0174 =  x102 &  x176 &  x204 &  x651 &  x653 &  x710 &  x743 & ~x52 & ~x112 & ~x137 & ~x141 & ~x144 & ~x164 & ~x169 & ~x219 & ~x223 & ~x283 & ~x419 & ~x445 & ~x448 & ~x477 & ~x480 & ~x499 & ~x500 & ~x503 & ~x504 & ~x532 & ~x535 & ~x588 & ~x612 & ~x613 & ~x668 & ~x669 & ~x674 & ~x727 & ~x756 & ~x781;
assign c0176 =  x8;
assign c0178 =  x233 &  x298 &  x405 &  x462 &  x519 &  x573 &  x575 &  x631 &  x632 &  x633 &  x656 &  x660 &  x663 & ~x60 & ~x86 & ~x303 & ~x306 & ~x342 & ~x343 & ~x357 & ~x363 & ~x371 & ~x399 & ~x422 & ~x479 & ~x480 & ~x553 & ~x594 & ~x612 & ~x704 & ~x733 & ~x760;
assign c0180 =  x264 &  x344 &  x596 &  x622 &  x629 &  x650 &  x736 &  x739 & ~x23 & ~x394 & ~x477 & ~x478 & ~x502 & ~x530 & ~x562 & ~x642;
assign c0182 =  x204 &  x260 &  x316 &  x320 &  x512 &  x682 &  x740 &  x763 & ~x141 & ~x167 & ~x421 & ~x673 & ~x698;
assign c0184 = ~x2 & ~x13 & ~x25 & ~x118 & ~x151 & ~x277 & ~x310 & ~x362 & ~x394 & ~x395 & ~x423 & ~x441 & ~x477 & ~x504 & ~x529 & ~x533 & ~x537 & ~x561 & ~x590 & ~x619 & ~x698 & ~x700 & ~x753 & ~x758;
assign c0186 =  x200 & ~x52 & ~x80 & ~x82 & ~x138 & ~x250 & ~x251 & ~x252 & ~x279 & ~x364 & ~x391 & ~x553 & ~x695 & ~x696 & ~x698 & ~x724 & ~x726 & ~x750 & ~x751 & ~x752 & ~x753 & ~x780;
assign c0188 =  x596 &  x623 &  x680 & ~x11 & ~x12 & ~x14 & ~x15 & ~x56 & ~x201 & ~x249 & ~x311 & ~x393 & ~x504 & ~x507 & ~x528 & ~x534 & ~x615 & ~x755 & ~x782;
assign c0190 =  x39 &  x44 &  x598 &  x652 & ~x1 & ~x4 & ~x5 & ~x6 & ~x7 & ~x8 & ~x19 & ~x20 & ~x21 & ~x22 & ~x23 & ~x24 & ~x25 & ~x26 & ~x30 & ~x32 & ~x34 & ~x49 & ~x51 & ~x52 & ~x53 & ~x54 & ~x55 & ~x56 & ~x57 & ~x58 & ~x59 & ~x60 & ~x61 & ~x79 & ~x80 & ~x82 & ~x83 & ~x84 & ~x85 & ~x86 & ~x87 & ~x109 & ~x113 & ~x115 & ~x138 & ~x141 & ~x142 & ~x143 & ~x166 & ~x167 & ~x169 & ~x170 & ~x171 & ~x198 & ~x222 & ~x225 & ~x251 & ~x252 & ~x253 & ~x254 & ~x279 & ~x281 & ~x305 & ~x306 & ~x307 & ~x308 & ~x334 & ~x335 & ~x336 & ~x337 & ~x339 & ~x362 & ~x363 & ~x364 & ~x365 & ~x366 & ~x367 & ~x385 & ~x386 & ~x387 & ~x388 & ~x389 & ~x392 & ~x393 & ~x396 & ~x414 & ~x415 & ~x416 & ~x418 & ~x419 & ~x420 & ~x421 & ~x422 & ~x425 & ~x445 & ~x447 & ~x448 & ~x450 & ~x452 & ~x470 & ~x475 & ~x477 & ~x478 & ~x479 & ~x480 & ~x498 & ~x500 & ~x502 & ~x503 & ~x505 & ~x506 & ~x509 & ~x526 & ~x527 & ~x529 & ~x530 & ~x531 & ~x532 & ~x534 & ~x535 & ~x536 & ~x537 & ~x538 & ~x554 & ~x557 & ~x558 & ~x559 & ~x560 & ~x563 & ~x564 & ~x565 & ~x583 & ~x585 & ~x586 & ~x588 & ~x590 & ~x592 & ~x593 & ~x594 & ~x610 & ~x612 & ~x615 & ~x616 & ~x617 & ~x618 & ~x619 & ~x620 & ~x621 & ~x638 & ~x639 & ~x640 & ~x641 & ~x643 & ~x644 & ~x646 & ~x649 & ~x667 & ~x669 & ~x670 & ~x672 & ~x677 & ~x694 & ~x695 & ~x696 & ~x697 & ~x699 & ~x701 & ~x704 & ~x722 & ~x723 & ~x725 & ~x726 & ~x727 & ~x728 & ~x730 & ~x731 & ~x732 & ~x733 & ~x750 & ~x752 & ~x755 & ~x756 & ~x757 & ~x760 & ~x778 & ~x779 & ~x780 & ~x781;
assign c0192 =  x68 &  x73 &  x285 &  x568 &  x629 & ~x4 & ~x23 & ~x24 & ~x31 & ~x85 & ~x111 & ~x138 & ~x168 & ~x196 & ~x280 & ~x362 & ~x393 & ~x503 & ~x504 & ~x615 & ~x642 & ~x672 & ~x699 & ~x703 & ~x758;
assign c0194 =  x41 &  x42 &  x44 &  x748 & ~x0 & ~x2 & ~x3 & ~x4 & ~x5 & ~x6 & ~x7 & ~x8 & ~x9 & ~x19 & ~x20 & ~x22 & ~x23 & ~x24 & ~x25 & ~x26 & ~x27 & ~x28 & ~x29 & ~x30 & ~x31 & ~x33 & ~x34 & ~x50 & ~x51 & ~x52 & ~x53 & ~x55 & ~x56 & ~x57 & ~x58 & ~x59 & ~x79 & ~x80 & ~x81 & ~x82 & ~x84 & ~x85 & ~x86 & ~x88 & ~x108 & ~x109 & ~x110 & ~x111 & ~x112 & ~x114 & ~x115 & ~x116 & ~x136 & ~x137 & ~x138 & ~x139 & ~x141 & ~x143 & ~x165 & ~x166 & ~x167 & ~x168 & ~x170 & ~x171 & ~x195 & ~x196 & ~x197 & ~x198 & ~x221 & ~x222 & ~x223 & ~x224 & ~x226 & ~x250 & ~x251 & ~x252 & ~x253 & ~x278 & ~x280 & ~x281 & ~x306 & ~x307 & ~x308 & ~x309 & ~x336 & ~x337 & ~x363 & ~x364 & ~x365 & ~x366 & ~x369 & ~x386 & ~x387 & ~x389 & ~x391 & ~x392 & ~x393 & ~x394 & ~x395 & ~x396 & ~x398 & ~x414 & ~x415 & ~x416 & ~x418 & ~x419 & ~x420 & ~x422 & ~x425 & ~x426 & ~x442 & ~x444 & ~x445 & ~x446 & ~x448 & ~x449 & ~x450 & ~x451 & ~x452 & ~x453 & ~x454 & ~x470 & ~x471 & ~x472 & ~x473 & ~x474 & ~x475 & ~x476 & ~x477 & ~x478 & ~x479 & ~x480 & ~x481 & ~x498 & ~x499 & ~x500 & ~x501 & ~x502 & ~x503 & ~x504 & ~x505 & ~x506 & ~x507 & ~x509 & ~x527 & ~x528 & ~x530 & ~x531 & ~x532 & ~x534 & ~x535 & ~x536 & ~x553 & ~x554 & ~x555 & ~x556 & ~x557 & ~x559 & ~x560 & ~x561 & ~x562 & ~x563 & ~x565 & ~x582 & ~x583 & ~x584 & ~x585 & ~x586 & ~x587 & ~x588 & ~x590 & ~x591 & ~x593 & ~x594 & ~x610 & ~x611 & ~x612 & ~x613 & ~x614 & ~x615 & ~x616 & ~x618 & ~x619 & ~x620 & ~x621 & ~x622 & ~x638 & ~x639 & ~x640 & ~x642 & ~x643 & ~x644 & ~x647 & ~x648 & ~x649 & ~x650 & ~x666 & ~x668 & ~x669 & ~x670 & ~x671 & ~x673 & ~x674 & ~x675 & ~x676 & ~x677 & ~x678 & ~x694 & ~x695 & ~x696 & ~x698 & ~x700 & ~x701 & ~x702 & ~x703 & ~x704 & ~x705 & ~x706 & ~x722 & ~x723 & ~x724 & ~x725 & ~x726 & ~x728 & ~x729 & ~x730 & ~x731 & ~x732 & ~x733 & ~x734 & ~x749 & ~x750 & ~x751 & ~x752 & ~x753 & ~x754 & ~x755 & ~x756 & ~x757 & ~x758 & ~x759 & ~x760 & ~x761 & ~x762 & ~x778 & ~x780 & ~x782 & ~x783;
assign c0196 =  x213 &  x214 &  x215 &  x233 &  x236 &  x242 &  x268 &  x290 &  x323 &  x345 &  x405 &  x408 &  x429 &  x430 &  x462 &  x463 &  x465 &  x485 &  x519 &  x542 &  x548 &  x577 &  x597 &  x601 &  x602 &  x605 &  x626 &  x628 &  x632 &  x659 &  x681 & ~x50 & ~x62 & ~x89 & ~x115 & ~x140 & ~x146 & ~x168 & ~x170 & ~x193 & ~x225 & ~x282 & ~x339 & ~x360 & ~x393 & ~x417 & ~x450 & ~x451 & ~x528 & ~x529 & ~x558 & ~x585 & ~x586 & ~x591 & ~x611 & ~x614 & ~x616 & ~x671 & ~x699 & ~x701 & ~x702 & ~x753;
assign c0198 =  x97 &  x214 &  x266 &  x269 &  x354 &  x401 &  x434 &  x464 &  x517 &  x599 &  x602 &  x605 &  x625 &  x629 &  x631 &  x655 &  x658 &  x660 & ~x3 & ~x5 & ~x23 & ~x24 & ~x53 & ~x85 & ~x107 & ~x140 & ~x166 & ~x250 & ~x255 & ~x278 & ~x281 & ~x339 & ~x386 & ~x396 & ~x397 & ~x413 & ~x441 & ~x445 & ~x446 & ~x447 & ~x450 & ~x470 & ~x478 & ~x497 & ~x502 & ~x525 & ~x557 & ~x561 & ~x610 & ~x637 & ~x638 & ~x646 & ~x722 & ~x750 & ~x756 & ~x781 & ~x783;
assign c0200 = ~x56 & ~x165 & ~x291 & ~x295 & ~x306 & ~x468 & ~x525 & ~x553 & ~x559 & ~x732 & ~x733 & ~x750 & ~x751;
assign c0202 =  x271 &  x299 &  x323 &  x405 &  x434 &  x437 &  x462 &  x465 &  x490 &  x546 &  x572 &  x579 &  x600 &  x634 &  x655 & ~x29 & ~x84 & ~x114 & ~x138 & ~x391 & ~x393 & ~x425 & ~x480 & ~x499 & ~x526 & ~x527 & ~x530 & ~x538 & ~x584 & ~x589 & ~x594 & ~x639 & ~x641 & ~x707 & ~x780;
assign c0204 =  x159 &  x177 &  x180 &  x259 &  x600 & ~x37 & ~x62 & ~x78 & ~x224 & ~x280 & ~x535 & ~x583 & ~x611 & ~x695 & ~x729;
assign c0206 =  x125 &  x242 &  x243 &  x354 &  x401 &  x457 &  x544 &  x572 &  x598 &  x602 &  x657 &  x769 &  x771 & ~x58 & ~x80 & ~x107 & ~x116 & ~x254 & ~x307 & ~x333 & ~x339 & ~x363 & ~x368 & ~x392 & ~x421 & ~x441 & ~x445 & ~x446 & ~x474 & ~x476 & ~x510 & ~x554 & ~x584 & ~x592 & ~x616 & ~x643 & ~x644 & ~x668 & ~x671 & ~x674 & ~x676 & ~x723 & ~x727 & ~x755 & ~x780;
assign c0208 = ~x93 & ~x102 & ~x129 & ~x334 & ~x566 & ~x610 & ~x658;
assign c0210 =  x231 &  x345 &  x748 & ~x20 & ~x51 & ~x81 & ~x84 & ~x142 & ~x251 & ~x253 & ~x338 & ~x361 & ~x365 & ~x369 & ~x389 & ~x392 & ~x416 & ~x417 & ~x444 & ~x472 & ~x475 & ~x482 & ~x501 & ~x510 & ~x532 & ~x537 & ~x558 & ~x618 & ~x620 & ~x640 & ~x646 & ~x674 & ~x678 & ~x702 & ~x723 & ~x726 & ~x728 & ~x729 & ~x730 & ~x732 & ~x755 & ~x760;
assign c0212 =  x736 &  x737 & ~x14 & ~x297;
assign c0214 = ~x94 & ~x413 & ~x418 & ~x441 & ~x538 & ~x577 & ~x583 & ~x605 & ~x610 & ~x752;
assign c0216 =  x204 &  x289 &  x568 & ~x5 & ~x8 & ~x33 & ~x52 & ~x79 & ~x138 & ~x169 & ~x281 & ~x304 & ~x333 & ~x448 & ~x478 & ~x496 & ~x561 & ~x647 & ~x671 & ~x695 & ~x699 & ~x700 & ~x702 & ~x722 & ~x781;
assign c0218 =  x129 &  x482 & ~x24 & ~x31 & ~x54 & ~x82 & ~x364 & ~x562 & ~x583 & ~x724;
assign c0220 = ~x205 & ~x322 & ~x565 & ~x614 & ~x638 & ~x667 & ~x733 & ~x750;
assign c0222 =  x39 &  x71 &  x215 & ~x197 & ~x308 & ~x336 & ~x363 & ~x587 & ~x623 & ~x704 & ~x706 & ~x724;
assign c0224 =  x297 & ~x58 & ~x156 & ~x415 & ~x453 & ~x502 & ~x528 & ~x565 & ~x593;
assign c0226 =  x198;
assign c0228 =  x257 &  x597 & ~x0 & ~x2 & ~x4 & ~x5 & ~x8 & ~x20 & ~x24 & ~x26 & ~x27 & ~x28 & ~x29 & ~x30 & ~x31 & ~x50 & ~x51 & ~x53 & ~x57 & ~x78 & ~x84 & ~x85 & ~x86 & ~x107 & ~x109 & ~x112 & ~x114 & ~x136 & ~x137 & ~x139 & ~x195 & ~x197 & ~x223 & ~x251 & ~x280 & ~x308 & ~x335 & ~x445 & ~x447 & ~x450 & ~x451 & ~x474 & ~x476 & ~x477 & ~x478 & ~x479 & ~x480 & ~x481 & ~x499 & ~x500 & ~x501 & ~x502 & ~x507 & ~x529 & ~x533 & ~x554 & ~x555 & ~x556 & ~x557 & ~x560 & ~x561 & ~x564 & ~x583 & ~x584 & ~x585 & ~x587 & ~x592 & ~x593 & ~x611 & ~x612 & ~x614 & ~x618 & ~x620 & ~x640 & ~x641 & ~x645 & ~x647 & ~x666 & ~x667 & ~x668 & ~x670 & ~x671 & ~x673 & ~x694 & ~x698 & ~x699 & ~x701 & ~x702 & ~x704 & ~x705 & ~x722 & ~x729 & ~x732 & ~x750 & ~x754 & ~x756 & ~x757 & ~x759 & ~x760 & ~x761 & ~x778 & ~x779 & ~x782 & ~x783;
assign c0230 =  x47 &  x372 &  x651 &  x735 & ~x110 & ~x223 & ~x225 & ~x360 & ~x415 & ~x500 & ~x501 & ~x531 & ~x534 & ~x560 & ~x584 & ~x587 & ~x647 & ~x674 & ~x753;
assign c0232 =  x193;
assign c0234 =  x226;
assign c0236 =  x130 &  x154 &  x157 &  x237 &  x289 &  x298 &  x574 &  x631 &  x659 &  x664 &  x691 & ~x27 & ~x33 & ~x89 & ~x134 & ~x162 & ~x190 & ~x250 & ~x508 & ~x509 & ~x588 & ~x704;
assign c0238 =  x16 &  x373 &  x598 & ~x0 & ~x1 & ~x2 & ~x3 & ~x4 & ~x5 & ~x21 & ~x23 & ~x27 & ~x28 & ~x29 & ~x30 & ~x32 & ~x54 & ~x56 & ~x58 & ~x59 & ~x82 & ~x84 & ~x85 & ~x113 & ~x140 & ~x141 & ~x169 & ~x278 & ~x280 & ~x281 & ~x308 & ~x336 & ~x337 & ~x364 & ~x390 & ~x391 & ~x393 & ~x394 & ~x419 & ~x420 & ~x421 & ~x422 & ~x445 & ~x446 & ~x448 & ~x449 & ~x450 & ~x474 & ~x478 & ~x506 & ~x530 & ~x532 & ~x533 & ~x534 & ~x561 & ~x562 & ~x587 & ~x588 & ~x592 & ~x593 & ~x611 & ~x613 & ~x615 & ~x639 & ~x641 & ~x642 & ~x647 & ~x648 & ~x666 & ~x668 & ~x673 & ~x674 & ~x675 & ~x676 & ~x696 & ~x698 & ~x699 & ~x700 & ~x701 & ~x703 & ~x704 & ~x724 & ~x725 & ~x727 & ~x728 & ~x729 & ~x731 & ~x751 & ~x752 & ~x753 & ~x755 & ~x756 & ~x757 & ~x760 & ~x761 & ~x779 & ~x782 & ~x783;
assign c0240 =  x233 &  x352 &  x403 &  x596 &  x659 & ~x58 & ~x111 & ~x119 & ~x172 & ~x202 & ~x229 & ~x246 & ~x390 & ~x445 & ~x565 & ~x619 & ~x726;
assign c0242 =  x77 &  x231 & ~x0 & ~x3 & ~x4 & ~x5 & ~x7 & ~x8 & ~x22 & ~x23 & ~x24 & ~x26 & ~x28 & ~x31 & ~x32 & ~x53 & ~x54 & ~x55 & ~x83 & ~x86 & ~x109 & ~x110 & ~x138 & ~x139 & ~x140 & ~x142 & ~x168 & ~x169 & ~x170 & ~x195 & ~x223 & ~x224 & ~x252 & ~x280 & ~x308 & ~x309 & ~x333 & ~x334 & ~x335 & ~x337 & ~x338 & ~x339 & ~x362 & ~x394 & ~x419 & ~x420 & ~x421 & ~x423 & ~x449 & ~x475 & ~x477 & ~x478 & ~x502 & ~x503 & ~x505 & ~x506 & ~x533 & ~x558 & ~x559 & ~x586 & ~x643 & ~x646 & ~x666 & ~x671 & ~x672 & ~x674 & ~x695 & ~x696 & ~x699 & ~x701 & ~x704 & ~x723 & ~x724 & ~x725 & ~x726 & ~x730 & ~x731 & ~x751 & ~x752 & ~x756 & ~x757 & ~x781;
assign c0244 = ~x58 & ~x94 & ~x120 & ~x126 & ~x129 & ~x158 & ~x333 & ~x528 & ~x553 & ~x726;
assign c0246 = ~x372 & ~x485 & ~x657 & ~x659;
assign c0248 =  x40 &  x217 &  x236 &  x246 &  x599 & ~x21 & ~x23 & ~x26 & ~x28 & ~x51 & ~x82 & ~x85 & ~x110 & ~x111 & ~x168 & ~x196 & ~x280 & ~x282 & ~x390 & ~x444 & ~x450 & ~x473 & ~x562 & ~x642 & ~x669 & ~x672 & ~x693 & ~x725 & ~x757 & ~x782;
assign c0250 =  x48 & ~x0 & ~x1 & ~x3 & ~x7 & ~x22 & ~x23 & ~x25 & ~x27 & ~x28 & ~x30 & ~x31 & ~x55 & ~x56 & ~x58 & ~x83 & ~x84 & ~x85 & ~x113 & ~x139 & ~x141 & ~x167 & ~x168 & ~x169 & ~x170 & ~x194 & ~x224 & ~x225 & ~x254 & ~x278 & ~x279 & ~x280 & ~x282 & ~x283 & ~x306 & ~x307 & ~x308 & ~x310 & ~x333 & ~x334 & ~x335 & ~x336 & ~x337 & ~x338 & ~x361 & ~x362 & ~x363 & ~x388 & ~x390 & ~x391 & ~x393 & ~x421 & ~x422 & ~x445 & ~x446 & ~x447 & ~x448 & ~x450 & ~x451 & ~x476 & ~x479 & ~x504 & ~x506 & ~x528 & ~x529 & ~x531 & ~x534 & ~x535 & ~x561 & ~x562 & ~x585 & ~x586 & ~x587 & ~x588 & ~x591 & ~x592 & ~x613 & ~x615 & ~x616 & ~x617 & ~x620 & ~x643 & ~x669 & ~x671 & ~x673 & ~x674 & ~x675 & ~x695 & ~x697 & ~x702 & ~x703 & ~x723 & ~x725 & ~x727 & ~x729 & ~x730 & ~x731 & ~x751 & ~x753 & ~x756 & ~x757 & ~x758 & ~x759 & ~x760 & ~x775 & ~x778 & ~x780 & ~x783;
assign c0252 =  x231 &  x736 & ~x5 & ~x58 & ~x83 & ~x87 & ~x112 & ~x167 & ~x168 & ~x250 & ~x252 & ~x306 & ~x309 & ~x313 & ~x330 & ~x358 & ~x361 & ~x363 & ~x369 & ~x389 & ~x395 & ~x396 & ~x397 & ~x422 & ~x443 & ~x448 & ~x453 & ~x473 & ~x477 & ~x479 & ~x526 & ~x536 & ~x562 & ~x564 & ~x585 & ~x592 & ~x593 & ~x594 & ~x616 & ~x620 & ~x639 & ~x644 & ~x645 & ~x669 & ~x674 & ~x676 & ~x699 & ~x701 & ~x705 & ~x724 & ~x752 & ~x781;
assign c0254 =  x339 &  x359;
assign c0256 =  x172 & ~x26 & ~x54 & ~x58 & ~x84 & ~x85 & ~x141 & ~x169 & ~x197 & ~x390 & ~x413 & ~x732 & ~x758;
assign c0258 =  x455 &  x599 & ~x56 & ~x168 & ~x335 & ~x533 & ~x534 & ~x558 & ~x562 & ~x583 & ~x588 & ~x591 & ~x617 & ~x619 & ~x645 & ~x672 & ~x699 & ~x701 & ~x731 & ~x756 & ~x768 & ~x775 & ~x778;
assign c0260 = ~x1 & ~x2 & ~x3 & ~x4 & ~x5 & ~x6 & ~x7 & ~x21 & ~x22 & ~x23 & ~x25 & ~x26 & ~x28 & ~x29 & ~x52 & ~x54 & ~x58 & ~x59 & ~x81 & ~x82 & ~x87 & ~x88 & ~x110 & ~x113 & ~x114 & ~x115 & ~x139 & ~x141 & ~x142 & ~x143 & ~x167 & ~x168 & ~x170 & ~x171 & ~x193 & ~x194 & ~x197 & ~x198 & ~x221 & ~x223 & ~x224 & ~x225 & ~x251 & ~x252 & ~x255 & ~x277 & ~x278 & ~x279 & ~x281 & ~x307 & ~x308 & ~x311 & ~x334 & ~x335 & ~x336 & ~x337 & ~x338 & ~x366 & ~x388 & ~x389 & ~x390 & ~x391 & ~x392 & ~x393 & ~x394 & ~x395 & ~x396 & ~x399 & ~x415 & ~x416 & ~x417 & ~x419 & ~x420 & ~x422 & ~x424 & ~x445 & ~x446 & ~x447 & ~x449 & ~x450 & ~x451 & ~x453 & ~x472 & ~x476 & ~x477 & ~x478 & ~x479 & ~x483 & ~x497 & ~x499 & ~x501 & ~x504 & ~x505 & ~x506 & ~x507 & ~x508 & ~x509 & ~x511 & ~x525 & ~x526 & ~x528 & ~x529 & ~x530 & ~x531 & ~x534 & ~x535 & ~x537 & ~x539 & ~x555 & ~x560 & ~x561 & ~x562 & ~x564 & ~x565 & ~x566 & ~x567 & ~x583 & ~x591 & ~x592 & ~x593 & ~x594 & ~x615 & ~x616 & ~x619 & ~x620 & ~x621 & ~x622 & ~x623 & ~x639 & ~x644 & ~x647 & ~x648 & ~x650 & ~x667 & ~x668 & ~x672 & ~x675 & ~x676 & ~x678 & ~x695 & ~x701 & ~x704 & ~x705 & ~x706 & ~x707 & ~x723 & ~x724 & ~x726 & ~x727 & ~x728 & ~x729 & ~x731 & ~x732 & ~x733 & ~x734 & ~x752 & ~x754 & ~x758 & ~x759 & ~x760 & ~x761 & ~x780 & ~x783;
assign c0262 =  x171 & ~x392 & ~x559 & ~x615 & ~x757;
assign c0264 =  x164 & ~x535;
assign c0266 =  x214 &  x236 &  x267 &  x323 &  x346 &  x433 &  x434 &  x462 &  x488 &  x489 & ~x15 & ~x22 & ~x52 & ~x54 & ~x59 & ~x80 & ~x87 & ~x110 & ~x141 & ~x166 & ~x167 & ~x169 & ~x170 & ~x172 & ~x221 & ~x250 & ~x251 & ~x252 & ~x280 & ~x281 & ~x304 & ~x308 & ~x310 & ~x311 & ~x332 & ~x335 & ~x337 & ~x364 & ~x389 & ~x391 & ~x394 & ~x450 & ~x472 & ~x475 & ~x505 & ~x506 & ~x532 & ~x533 & ~x535 & ~x560 & ~x585 & ~x611 & ~x615 & ~x616 & ~x618 & ~x642 & ~x646 & ~x647 & ~x674 & ~x731 & ~x755 & ~x758 & ~x759 & ~x763 & ~x765 & ~x775 & ~x778 & ~x780;
assign c0268 = ~x3 & ~x14 & ~x81 & ~x104 & ~x133 & ~x160 & ~x162 & ~x164 & ~x167 & ~x197 & ~x302 & ~x332 & ~x384 & ~x426 & ~x444 & ~x450 & ~x473 & ~x482 & ~x497 & ~x504 & ~x508 & ~x528 & ~x532 & ~x553 & ~x558 & ~x586 & ~x589 & ~x616 & ~x669 & ~x671 & ~x703 & ~x705 & ~x723 & ~x726 & ~x732 & ~x733 & ~x774 & ~x778;
assign c0270 =  x286 &  x330 &  x340 &  x369 &  x387 &  x396 &  x656 &  x681 & ~x559 & ~x728;
assign c0272 =  x39 &  x40 &  x41 &  x42 &  x43 &  x44 &  x601 & ~x3 & ~x5 & ~x7 & ~x20 & ~x21 & ~x24 & ~x25 & ~x26 & ~x27 & ~x31 & ~x32 & ~x33 & ~x50 & ~x52 & ~x53 & ~x55 & ~x56 & ~x57 & ~x59 & ~x82 & ~x84 & ~x85 & ~x86 & ~x112 & ~x114 & ~x115 & ~x137 & ~x142 & ~x143 & ~x166 & ~x169 & ~x170 & ~x195 & ~x197 & ~x198 & ~x221 & ~x224 & ~x225 & ~x226 & ~x250 & ~x251 & ~x253 & ~x277 & ~x279 & ~x305 & ~x307 & ~x308 & ~x335 & ~x336 & ~x339 & ~x362 & ~x363 & ~x365 & ~x366 & ~x367 & ~x368 & ~x369 & ~x370 & ~x386 & ~x388 & ~x389 & ~x392 & ~x393 & ~x395 & ~x396 & ~x397 & ~x416 & ~x417 & ~x420 & ~x426 & ~x441 & ~x442 & ~x445 & ~x447 & ~x449 & ~x450 & ~x451 & ~x452 & ~x453 & ~x469 & ~x471 & ~x472 & ~x478 & ~x479 & ~x480 & ~x481 & ~x497 & ~x498 & ~x499 & ~x503 & ~x504 & ~x506 & ~x507 & ~x509 & ~x510 & ~x527 & ~x529 & ~x531 & ~x532 & ~x534 & ~x538 & ~x554 & ~x556 & ~x558 & ~x561 & ~x563 & ~x564 & ~x565 & ~x566 & ~x581 & ~x582 & ~x583 & ~x585 & ~x586 & ~x588 & ~x590 & ~x591 & ~x592 & ~x593 & ~x594 & ~x609 & ~x614 & ~x618 & ~x619 & ~x620 & ~x638 & ~x639 & ~x640 & ~x641 & ~x645 & ~x649 & ~x665 & ~x666 & ~x668 & ~x670 & ~x671 & ~x672 & ~x673 & ~x674 & ~x675 & ~x677 & ~x678 & ~x693 & ~x695 & ~x696 & ~x700 & ~x701 & ~x702 & ~x705 & ~x706 & ~x721 & ~x729 & ~x730 & ~x749 & ~x752 & ~x753 & ~x754 & ~x755 & ~x756 & ~x757 & ~x760 & ~x761 & ~x763 & ~x777 & ~x778 & ~x780 & ~x782;
assign c0274 =  x38 &  x69 &  x76 &  x130 &  x131 &  x317 &  x459 &  x545 &  x575 &  x603 &  x633 & ~x1 & ~x4 & ~x7 & ~x22 & ~x29 & ~x53 & ~x139 & ~x140 & ~x142 & ~x167 & ~x168 & ~x170 & ~x196 & ~x222 & ~x250 & ~x311 & ~x360 & ~x363 & ~x397 & ~x417 & ~x446 & ~x451 & ~x475 & ~x479 & ~x507 & ~x530 & ~x589 & ~x593 & ~x612 & ~x618 & ~x620 & ~x639 & ~x643 & ~x672 & ~x700 & ~x754 & ~x758 & ~x760 & ~x780;
assign c0276 = ~x19 & ~x26 & ~x28 & ~x29 & ~x33 & ~x52 & ~x54 & ~x108 & ~x113 & ~x115 & ~x142 & ~x168 & ~x195 & ~x225 & ~x327 & ~x361 & ~x362 & ~x367 & ~x390 & ~x416 & ~x438 & ~x445 & ~x447 & ~x472 & ~x475 & ~x480 & ~x497 & ~x502 & ~x525 & ~x526 & ~x529 & ~x534 & ~x553 & ~x554 & ~x555 & ~x561 & ~x581 & ~x587 & ~x609 & ~x610 & ~x611 & ~x612 & ~x616 & ~x618 & ~x638 & ~x669 & ~x670 & ~x673 & ~x674 & ~x695 & ~x696 & ~x700 & ~x732 & ~x751 & ~x754 & ~x755 & ~x756 & ~x778;
assign c0278 =  x78 & ~x0 & ~x4 & ~x28 & ~x29 & ~x85 & ~x196 & ~x393 & ~x422 & ~x476 & ~x477 & ~x505 & ~x532 & ~x560 & ~x566 & ~x587 & ~x615 & ~x671 & ~x674 & ~x723 & ~x724 & ~x729 & ~x731;
assign c0280 = ~x4 & ~x51 & ~x80 & ~x107 & ~x111 & ~x141 & ~x195 & ~x197 & ~x198 & ~x237 & ~x238 & ~x239 & ~x280 & ~x334 & ~x337 & ~x361 & ~x395 & ~x417 & ~x419 & ~x441 & ~x450 & ~x452 & ~x454 & ~x482 & ~x502 & ~x506 & ~x554 & ~x560 & ~x564 & ~x566 & ~x609 & ~x615 & ~x622 & ~x642 & ~x668 & ~x695 & ~x697 & ~x702 & ~x703 & ~x704 & ~x722 & ~x730 & ~x733 & ~x753 & ~x759 & ~x762 & ~x777;
assign c0282 =  x215 &  x542 &  x543 &  x548 &  x568 &  x575 &  x596 & ~x12 & ~x13 & ~x30 & ~x88 & ~x89 & ~x112 & ~x135 & ~x138 & ~x173 & ~x192 & ~x193 & ~x201 & ~x250 & ~x254 & ~x275 & ~x390 & ~x416 & ~x422 & ~x449 & ~x477 & ~x501 & ~x503 & ~x536 & ~x562 & ~x586 & ~x591 & ~x645 & ~x668 & ~x730 & ~x731 & ~x753 & ~x782;
assign c0284 =  x79;
assign c0286 = ~x30 & ~x81 & ~x102 & ~x119 & ~x123 & ~x124 & ~x128 & ~x147 & ~x167 & ~x307 & ~x390 & ~x421 & ~x449 & ~x452 & ~x471 & ~x475 & ~x476 & ~x477 & ~x500 & ~x501 & ~x506 & ~x533 & ~x535 & ~x537 & ~x589 & ~x640 & ~x726;
assign c0288 =  x45 &  x162 &  x218 & ~x1 & ~x2 & ~x8 & ~x19 & ~x22 & ~x25 & ~x27 & ~x33 & ~x34 & ~x54 & ~x79 & ~x81 & ~x82 & ~x84 & ~x86 & ~x87 & ~x109 & ~x113 & ~x114 & ~x140 & ~x307 & ~x335 & ~x337 & ~x363 & ~x364 & ~x391 & ~x394 & ~x450 & ~x501 & ~x502 & ~x505 & ~x529 & ~x531 & ~x533 & ~x586 & ~x588 & ~x592 & ~x610 & ~x611 & ~x614 & ~x619 & ~x638 & ~x642 & ~x643 & ~x647 & ~x666 & ~x667 & ~x670 & ~x672 & ~x675 & ~x696 & ~x699 & ~x702 & ~x724 & ~x727 & ~x728 & ~x754 & ~x755 & ~x758 & ~x778 & ~x780 & ~x781 & ~x782;
assign c0290 =  x736 & ~x7 & ~x349 & ~x730;
assign c0292 =  x40 &  x44 &  x45 &  x218 & ~x1 & ~x5 & ~x6 & ~x7 & ~x22 & ~x27 & ~x28 & ~x32 & ~x33 & ~x53 & ~x81 & ~x85 & ~x86 & ~x109 & ~x138 & ~x139 & ~x142 & ~x171 & ~x193 & ~x196 & ~x198 & ~x251 & ~x252 & ~x279 & ~x305 & ~x310 & ~x333 & ~x361 & ~x391 & ~x418 & ~x449 & ~x475 & ~x476 & ~x478 & ~x502 & ~x506 & ~x531 & ~x558 & ~x562 & ~x588 & ~x590 & ~x614 & ~x619 & ~x641 & ~x642 & ~x646 & ~x666 & ~x668 & ~x669 & ~x676 & ~x694 & ~x695 & ~x696 & ~x699 & ~x702 & ~x726 & ~x729 & ~x730 & ~x755 & ~x759 & ~x778 & ~x780 & ~x781 & ~x783;
assign c0294 =  x98 &  x179 &  x180 &  x233 &  x263 &  x289 &  x298 &  x317 &  x402 &  x598 &  x599 &  x628 &  x653 &  x654 &  x685 &  x687 &  x716 & ~x6 & ~x33 & ~x78 & ~x138 & ~x191 & ~x225 & ~x247 & ~x277 & ~x309 & ~x417 & ~x565 & ~x587 & ~x591 & ~x617 & ~x638 & ~x697 & ~x759 & ~x761;
assign c0296 =  x13 &  x624 & ~x6 & ~x7 & ~x28 & ~x29 & ~x54 & ~x82 & ~x196 & ~x281 & ~x282 & ~x364 & ~x390 & ~x393 & ~x502 & ~x504 & ~x558 & ~x561 & ~x587 & ~x593 & ~x618 & ~x621 & ~x650 & ~x705 & ~x724 & ~x729 & ~x731 & ~x734 & ~x752 & ~x755 & ~x758;
assign c0298 = ~x0 & ~x4 & ~x34 & ~x52 & ~x54 & ~x82 & ~x86 & ~x136 & ~x140 & ~x166 & ~x168 & ~x223 & ~x227 & ~x393 & ~x418 & ~x445 & ~x473 & ~x474 & ~x483 & ~x502 & ~x529 & ~x557 & ~x588 & ~x594 & ~x676 & ~x704 & ~x707 & ~x710 & ~x731 & ~x733 & ~x734 & ~x751 & ~x753 & ~x762 & ~x766 & ~x768 & ~x769 & ~x771 & ~x772 & ~x782;
assign c0300 = ~x97 & ~x100 & ~x103 & ~x446 & ~x499 & ~x733 & ~x766 & ~x772;
assign c0302 =  x289 &  x373 &  x457 &  x461 & ~x0 & ~x5 & ~x6 & ~x21 & ~x30 & ~x31 & ~x54 & ~x58 & ~x81 & ~x86 & ~x108 & ~x113 & ~x116 & ~x137 & ~x138 & ~x141 & ~x168 & ~x170 & ~x194 & ~x197 & ~x198 & ~x199 & ~x220 & ~x226 & ~x248 & ~x254 & ~x276 & ~x280 & ~x281 & ~x304 & ~x307 & ~x308 & ~x311 & ~x334 & ~x338 & ~x362 & ~x384 & ~x393 & ~x412 & ~x419 & ~x420 & ~x421 & ~x422 & ~x423 & ~x446 & ~x450 & ~x451 & ~x454 & ~x469 & ~x472 & ~x478 & ~x501 & ~x506 & ~x525 & ~x526 & ~x532 & ~x533 & ~x534 & ~x560 & ~x561 & ~x565 & ~x582 & ~x587 & ~x588 & ~x591 & ~x615 & ~x618 & ~x619 & ~x622 & ~x641 & ~x642 & ~x643 & ~x644 & ~x669 & ~x670 & ~x673 & ~x695 & ~x696 & ~x697 & ~x698 & ~x706 & ~x722 & ~x726 & ~x728 & ~x732 & ~x749 & ~x751 & ~x760 & ~x778 & ~x779 & ~x781 & ~x782;
assign c0304 =  x135 & ~x7 & ~x33 & ~x113 & ~x114 & ~x137 & ~x140 & ~x142 & ~x167 & ~x194 & ~x224 & ~x280 & ~x479 & ~x564 & ~x619 & ~x641 & ~x669 & ~x673 & ~x675 & ~x700 & ~x703 & ~x728;
assign c0306 = ~x566 & ~x604 & ~x606 & ~x607;
assign c0308 = ~x14 & ~x23 & ~x55 & ~x79 & ~x110 & ~x112 & ~x142 & ~x166 & ~x248 & ~x255 & ~x306 & ~x311 & ~x332 & ~x334 & ~x388 & ~x446 & ~x468 & ~x475 & ~x476 & ~x530 & ~x555 & ~x585 & ~x609 & ~x614 & ~x638 & ~x647 & ~x669 & ~x671 & ~x694 & ~x695 & ~x698 & ~x721 & ~x733 & ~x751 & ~x771 & ~x773 & ~x774;
assign c0310 = ~x57 & ~x279 & ~x516 & ~x575 & ~x621 & ~x631 & ~x666 & ~x722;
assign c0312 =  x164 & ~x589 & ~x615;
assign c0314 =  x569 &  x570 & ~x2 & ~x5 & ~x18 & ~x36 & ~x112 & ~x140 & ~x142 & ~x167 & ~x171 & ~x198 & ~x223 & ~x225 & ~x254 & ~x277 & ~x280 & ~x310 & ~x311 & ~x334 & ~x336 & ~x342 & ~x360 & ~x362 & ~x368 & ~x413 & ~x415 & ~x418 & ~x423 & ~x425 & ~x442 & ~x447 & ~x448 & ~x451 & ~x453 & ~x474 & ~x477 & ~x481 & ~x482 & ~x483 & ~x497 & ~x503 & ~x504 & ~x507 & ~x508 & ~x554 & ~x560 & ~x566 & ~x583 & ~x587 & ~x611 & ~x615 & ~x617 & ~x620 & ~x641 & ~x644 & ~x649 & ~x669 & ~x671 & ~x676 & ~x725 & ~x728 & ~x731 & ~x749 & ~x750 & ~x758 & ~x759 & ~x760 & ~x762 & ~x777 & ~x778 & ~x783;
assign c0316 = ~x440 & ~x494 & ~x522 & ~x602 & ~x609;
assign c0318 =  x290 &  x351 &  x376 &  x517 &  x770 & ~x22 & ~x27 & ~x35 & ~x58 & ~x119 & ~x140 & ~x147 & ~x166 & ~x199 & ~x280 & ~x281 & ~x305 & ~x420 & ~x474 & ~x477 & ~x500 & ~x558 & ~x559 & ~x646 & ~x727;
assign c0320 =  x43 &  x78 & ~x6 & ~x365 & ~x367 & ~x391 & ~x475 & ~x476 & ~x617 & ~x619 & ~x673 & ~x675 & ~x697 & ~x759;
assign c0322 =  x43 &  x44 & ~x52 & ~x56 & ~x59 & ~x83 & ~x110 & ~x165 & ~x169 & ~x251 & ~x268 & ~x308 & ~x362 & ~x392 & ~x394 & ~x424 & ~x475 & ~x558 & ~x592 & ~x617 & ~x668 & ~x676 & ~x706 & ~x723 & ~x726 & ~x756;
assign c0324 = ~x4 & ~x52 & ~x109 & ~x336 & ~x393 & ~x417 & ~x445 & ~x450 & ~x454 & ~x458 & ~x462 & ~x470 & ~x471 & ~x477 & ~x482 & ~x498 & ~x501 & ~x534 & ~x583 & ~x618 & ~x638 & ~x647 & ~x650 & ~x668 & ~x675 & ~x706 & ~x723 & ~x751 & ~x752 & ~x753 & ~x778;
assign c0326 = ~x91 & ~x152 & ~x328 & ~x472 & ~x563 & ~x564 & ~x592 & ~x609 & ~x733 & ~x752;
assign c0328 = ~x92 & ~x130 & ~x180 & ~x362 & ~x469 & ~x497 & ~x525 & ~x529 & ~x536 & ~x538 & ~x557 & ~x638 & ~x694 & ~x723;
assign c0330 =  x42 &  x44 &  x737 &  x740 &  x745 &  x767 &  x768 &  x769 &  x770 &  x771 &  x772 & ~x0 & ~x1 & ~x2 & ~x26 & ~x55 & ~x57 & ~x58 & ~x59 & ~x86 & ~x109 & ~x110 & ~x195 & ~x281 & ~x309 & ~x334 & ~x337 & ~x366 & ~x391 & ~x395 & ~x427 & ~x445 & ~x446 & ~x447 & ~x448 & ~x452 & ~x455 & ~x474 & ~x475 & ~x499 & ~x530 & ~x532 & ~x533 & ~x557 & ~x560 & ~x584 & ~x590 & ~x611 & ~x614 & ~x615 & ~x619 & ~x620 & ~x645 & ~x648 & ~x668 & ~x670 & ~x698 & ~x724 & ~x752 & ~x756 & ~x757;
assign c0332 = ~x383 & ~x495 & ~x522 & ~x576 & ~x607 & ~x694 & ~x750;
assign c0334 =  x73 &  x93 &  x98 &  x127 &  x187 &  x293 &  x327 &  x355 &  x516 &  x551 &  x569 &  x653 &  x716 &  x746 &  x747 &  x749 & ~x88 & ~x252 & ~x254;
assign c0336 = ~x6 & ~x22 & ~x98 & ~x141 & ~x195 & ~x414 & ~x425 & ~x451 & ~x453 & ~x473 & ~x477 & ~x500 & ~x507 & ~x526 & ~x528 & ~x537 & ~x558 & ~x585 & ~x610 & ~x643 & ~x697 & ~x751 & ~x766 & ~x767 & ~x773 & ~x781 & ~x783;
assign c0338 =  x9 &  x46 &  x627 & ~x223 & ~x225 & ~x280 & ~x310 & ~x416 & ~x478 & ~x533 & ~x589 & ~x672 & ~x760;
assign c0340 =  x179 &  x205 &  x242 &  x351 &  x353 &  x462 &  x601 &  x602 & ~x1 & ~x6 & ~x21 & ~x30 & ~x33 & ~x53 & ~x78 & ~x86 & ~x105 & ~x106 & ~x108 & ~x144 & ~x146 & ~x161 & ~x164 & ~x165 & ~x169 & ~x189 & ~x196 & ~x202 & ~x255 & ~x331 & ~x336 & ~x339 & ~x360 & ~x390 & ~x444 & ~x477 & ~x478 & ~x505 & ~x528 & ~x529 & ~x556 & ~x560 & ~x588 & ~x612 & ~x616 & ~x669 & ~x698 & ~x700 & ~x753;
assign c0342 = ~x2 & ~x111 & ~x344 & ~x391 & ~x502 & ~x508 & ~x627 & ~x709 & ~x710 & ~x750;
assign c0344 = ~x343 & ~x371 & ~x479 & ~x649 & ~x706 & ~x740 & ~x746;
assign c0346 =  x43 &  x99 &  x178 &  x290 &  x353 &  x381 &  x402 &  x404 &  x430 &  x431 &  x436 &  x437 &  x544 &  x570 &  x573 &  x599 &  x600 &  x629 &  x656 &  x714 & ~x0 & ~x7 & ~x21 & ~x23 & ~x24 & ~x28 & ~x29 & ~x30 & ~x51 & ~x55 & ~x58 & ~x60 & ~x79 & ~x82 & ~x86 & ~x88 & ~x110 & ~x113 & ~x115 & ~x136 & ~x139 & ~x143 & ~x144 & ~x164 & ~x165 & ~x166 & ~x167 & ~x193 & ~x195 & ~x196 & ~x198 & ~x221 & ~x250 & ~x254 & ~x277 & ~x278 & ~x281 & ~x282 & ~x283 & ~x305 & ~x307 & ~x311 & ~x336 & ~x339 & ~x362 & ~x419 & ~x420 & ~x445 & ~x446 & ~x449 & ~x479 & ~x504 & ~x531 & ~x533 & ~x556 & ~x557 & ~x558 & ~x561 & ~x564 & ~x581 & ~x584 & ~x586 & ~x587 & ~x617 & ~x637 & ~x638 & ~x665 & ~x666 & ~x671 & ~x677 & ~x693 & ~x694 & ~x699 & ~x701 & ~x721 & ~x722 & ~x725 & ~x727 & ~x730 & ~x731 & ~x750 & ~x751 & ~x752 & ~x754 & ~x755 & ~x759 & ~x760 & ~x777;
assign c0348 = ~x102 & ~x129 & ~x177 & ~x180 & ~x444 & ~x482 & ~x497 & ~x612 & ~x732;
assign c0350 =  x41 &  x42 &  x43 &  x44 &  x520 & ~x0 & ~x1 & ~x2 & ~x3 & ~x4 & ~x5 & ~x6 & ~x7 & ~x8 & ~x9 & ~x18 & ~x19 & ~x20 & ~x21 & ~x22 & ~x23 & ~x24 & ~x25 & ~x26 & ~x27 & ~x28 & ~x29 & ~x30 & ~x31 & ~x33 & ~x34 & ~x35 & ~x49 & ~x50 & ~x51 & ~x52 & ~x53 & ~x54 & ~x55 & ~x56 & ~x57 & ~x58 & ~x59 & ~x60 & ~x79 & ~x80 & ~x81 & ~x82 & ~x83 & ~x84 & ~x86 & ~x87 & ~x88 & ~x108 & ~x109 & ~x110 & ~x111 & ~x112 & ~x113 & ~x114 & ~x115 & ~x137 & ~x140 & ~x141 & ~x142 & ~x165 & ~x166 & ~x168 & ~x169 & ~x171 & ~x193 & ~x194 & ~x195 & ~x196 & ~x197 & ~x198 & ~x221 & ~x223 & ~x224 & ~x225 & ~x226 & ~x250 & ~x251 & ~x252 & ~x253 & ~x279 & ~x280 & ~x281 & ~x307 & ~x308 & ~x309 & ~x334 & ~x335 & ~x336 & ~x337 & ~x338 & ~x339 & ~x362 & ~x363 & ~x364 & ~x365 & ~x366 & ~x367 & ~x368 & ~x389 & ~x390 & ~x391 & ~x392 & ~x393 & ~x394 & ~x395 & ~x396 & ~x397 & ~x413 & ~x414 & ~x415 & ~x416 & ~x417 & ~x418 & ~x419 & ~x420 & ~x421 & ~x422 & ~x423 & ~x442 & ~x446 & ~x447 & ~x448 & ~x449 & ~x450 & ~x451 & ~x452 & ~x453 & ~x470 & ~x472 & ~x473 & ~x474 & ~x475 & ~x476 & ~x478 & ~x479 & ~x498 & ~x499 & ~x501 & ~x502 & ~x503 & ~x504 & ~x505 & ~x507 & ~x510 & ~x528 & ~x529 & ~x530 & ~x531 & ~x532 & ~x533 & ~x534 & ~x536 & ~x537 & ~x554 & ~x556 & ~x558 & ~x559 & ~x560 & ~x561 & ~x562 & ~x564 & ~x581 & ~x582 & ~x584 & ~x586 & ~x587 & ~x588 & ~x589 & ~x590 & ~x592 & ~x593 & ~x609 & ~x610 & ~x611 & ~x612 & ~x613 & ~x614 & ~x615 & ~x616 & ~x617 & ~x618 & ~x619 & ~x620 & ~x621 & ~x622 & ~x638 & ~x639 & ~x640 & ~x641 & ~x642 & ~x644 & ~x645 & ~x646 & ~x647 & ~x648 & ~x649 & ~x667 & ~x669 & ~x670 & ~x671 & ~x672 & ~x673 & ~x674 & ~x675 & ~x676 & ~x678 & ~x694 & ~x695 & ~x696 & ~x697 & ~x698 & ~x699 & ~x700 & ~x701 & ~x703 & ~x704 & ~x705 & ~x722 & ~x723 & ~x724 & ~x725 & ~x727 & ~x728 & ~x729 & ~x730 & ~x731 & ~x732 & ~x733 & ~x734 & ~x750 & ~x751 & ~x752 & ~x753 & ~x754 & ~x755 & ~x757 & ~x758 & ~x759 & ~x760 & ~x761 & ~x762 & ~x778 & ~x779 & ~x780 & ~x781 & ~x782 & ~x783;
assign c0352 =  x177 &  x179 &  x183 &  x202 &  x687 & ~x254 & ~x643 & ~x705 & ~x782;
assign c0354 =  x238 &  x461 &  x518 &  x607 & ~x63 & ~x119 & ~x217 & ~x257;
assign c0356 =  x737 &  x740 &  x741 &  x743 &  x744 &  x745 &  x746 & ~x24 & ~x54 & ~x139 & ~x151 & ~x391 & ~x422 & ~x643 & ~x645 & ~x672 & ~x674;
assign c0358 =  x269 &  x296 &  x353 &  x486 &  x490 &  x544 &  x545 &  x570 &  x574 &  x605 &  x655 & ~x1 & ~x2 & ~x4 & ~x13 & ~x27 & ~x37 & ~x59 & ~x60 & ~x85 & ~x86 & ~x113 & ~x116 & ~x223 & ~x501 & ~x504 & ~x507 & ~x528 & ~x529 & ~x563 & ~x584 & ~x586 & ~x592 & ~x612 & ~x640 & ~x641 & ~x646 & ~x668 & ~x673 & ~x697 & ~x700 & ~x703 & ~x761;
assign c0360 =  x116 & ~x58 & ~x139 & ~x141 & ~x563 & ~x646;
assign c0362 = ~x24 & ~x52 & ~x67 & ~x72 & ~x73 & ~x74 & ~x397 & ~x414 & ~x415 & ~x446 & ~x470 & ~x479 & ~x536 & ~x565 & ~x583 & ~x621 & ~x648 & ~x700 & ~x754 & ~x778;
assign c0364 =  x236 &  x512 &  x567 &  x628 &  x776 & ~x368 & ~x452 & ~x558 & ~x699;
assign c0366 =  x77 &  x220 & ~x83 & ~x84 & ~x85 & ~x168 & ~x335 & ~x588 & ~x675 & ~x699;
assign c0368 =  x69 &  x134 &  x146 &  x190 &  x247 &  x550 &  x661 &  x720 &  x748 & ~x28 & ~x55 & ~x60 & ~x110 & ~x141 & ~x194 & ~x195 & ~x477 & ~x559 & ~x588;
assign c0370 = ~x488 & ~x686 & ~x750;
assign c0372 =  x313 &  x367 & ~x224;
assign c0374 =  x137;
assign c0376 =  x261 &  x267 &  x271 &  x289 &  x290 &  x317 &  x408 &  x550 &  x598 &  x600 &  x605 & ~x28 & ~x37 & ~x86 & ~x168 & ~x334 & ~x337 & ~x362 & ~x475 & ~x527 & ~x529 & ~x562 & ~x585 & ~x612 & ~x617 & ~x695 & ~x700 & ~x726 & ~x760 & ~x761;
assign c0378 =  x39 &  x40 &  x41 &  x42 &  x43 &  x44 &  x600 &  x628 &  x634 &  x709 &  x748 & ~x0 & ~x1 & ~x2 & ~x4 & ~x5 & ~x22 & ~x23 & ~x26 & ~x28 & ~x31 & ~x51 & ~x52 & ~x57 & ~x61 & ~x82 & ~x84 & ~x85 & ~x86 & ~x87 & ~x110 & ~x111 & ~x112 & ~x113 & ~x114 & ~x116 & ~x137 & ~x138 & ~x141 & ~x142 & ~x168 & ~x169 & ~x196 & ~x197 & ~x251 & ~x252 & ~x253 & ~x280 & ~x282 & ~x308 & ~x309 & ~x334 & ~x335 & ~x336 & ~x337 & ~x362 & ~x363 & ~x366 & ~x392 & ~x419 & ~x421 & ~x422 & ~x447 & ~x448 & ~x449 & ~x450 & ~x474 & ~x475 & ~x476 & ~x477 & ~x503 & ~x505 & ~x533 & ~x559 & ~x560 & ~x587 & ~x588 & ~x645 & ~x671 & ~x672 & ~x673 & ~x674 & ~x699 & ~x700 & ~x704 & ~x724 & ~x726 & ~x728 & ~x730 & ~x731 & ~x733 & ~x753 & ~x755 & ~x756 & ~x757 & ~x759 & ~x760 & ~x780 & ~x781 & ~x782 & ~x783;
assign c0380 =  x507 & ~x29 & ~x253;
assign c0382 =  x191 & ~x29 & ~x56 & ~x84 & ~x140 & ~x304 & ~x306 & ~x308 & ~x334 & ~x363 & ~x390 & ~x392 & ~x393 & ~x418 & ~x473 & ~x478 & ~x501 & ~x505 & ~x534 & ~x587 & ~x615 & ~x616 & ~x641 & ~x642 & ~x668 & ~x672 & ~x674 & ~x698 & ~x699 & ~x700 & ~x703 & ~x731 & ~x751 & ~x779;
assign c0384 = ~x27 & ~x81 & ~x92 & ~x154 & ~x337 & ~x363 & ~x387 & ~x451 & ~x482 & ~x499 & ~x536 & ~x560 & ~x668 & ~x676 & ~x678 & ~x705 & ~x749 & ~x766;
assign c0386 = ~x140 & ~x444 & ~x520 & ~x521 & ~x547 & ~x609 & ~x621 & ~x639 & ~x750 & ~x756 & ~x762 & ~x778;
assign c0388 =  x482 & ~x13 & ~x14 & ~x40 & ~x41;
assign c0390 =  x388 &  x422 &  x472;
assign c0392 = ~x399 & ~x469 & ~x626 & ~x627 & ~x629 & ~x632;
assign c0394 =  x289 &  x375 &  x378 &  x461 &  x514 &  x573 &  x578 &  x626 &  x630 &  x658 & ~x2 & ~x22 & ~x25 & ~x30 & ~x61 & ~x79 & ~x139 & ~x173 & ~x224 & ~x255 & ~x258 & ~x281 & ~x282 & ~x363 & ~x365 & ~x385 & ~x395 & ~x397 & ~x419 & ~x441 & ~x472 & ~x525 & ~x532 & ~x553 & ~x586 & ~x591 & ~x610 & ~x617 & ~x645 & ~x699 & ~x723 & ~x730 & ~x757 & ~x783;
assign c0396 =  x214 &  x603 &  x607 &  x662 &  x689 & ~x91 & ~x371 & ~x530 & ~x566 & ~x669 & ~x734;
assign c0398 = ~x19 & ~x26 & ~x61 & ~x81 & ~x87 & ~x308 & ~x333 & ~x334 & ~x384 & ~x394 & ~x450 & ~x451 & ~x483 & ~x501 & ~x504 & ~x533 & ~x553 & ~x564 & ~x581 & ~x592 & ~x649 & ~x664 & ~x665 & ~x666 & ~x674 & ~x691 & ~x695 & ~x704 & ~x723 & ~x725 & ~x729 & ~x772 & ~x773;
assign c0400 =  x298 & ~x2 & ~x24 & ~x32 & ~x82 & ~x83 & ~x111 & ~x129 & ~x196 & ~x307 & ~x308 & ~x366 & ~x421 & ~x444 & ~x450 & ~x500 & ~x501 & ~x510 & ~x531 & ~x533 & ~x535 & ~x558 & ~x559 & ~x564 & ~x585 & ~x591 & ~x613 & ~x615 & ~x618 & ~x641 & ~x646 & ~x672 & ~x675 & ~x699 & ~x756;
assign c0402 =  x229 &  x339 &  x359 &  x395;
assign c0404 =  x102 &  x126 &  x129 &  x149 &  x151 &  x152 &  x156 &  x177 &  x181 &  x183 &  x187 &  x206 &  x214 &  x233 &  x237 &  x266 &  x290 &  x291 &  x292 &  x298 &  x317 &  x321 &  x325 &  x346 &  x347 &  x348 &  x353 &  x402 &  x403 &  x404 &  x429 &  x432 &  x433 &  x437 &  x457 &  x460 &  x464 &  x465 &  x485 &  x488 &  x490 &  x492 &  x514 &  x516 &  x517 &  x518 &  x519 &  x544 &  x546 &  x548 &  x570 &  x571 &  x574 &  x597 &  x598 &  x600 &  x602 &  x603 &  x604 &  x605 &  x606 &  x629 &  x630 &  x632 &  x653 &  x655 & ~x3 & ~x4 & ~x22 & ~x54 & ~x57 & ~x58 & ~x60 & ~x78 & ~x84 & ~x112 & ~x114 & ~x138 & ~x141 & ~x144 & ~x169 & ~x196 & ~x223 & ~x249 & ~x278 & ~x280 & ~x281 & ~x308 & ~x334 & ~x336 & ~x363 & ~x364 & ~x368 & ~x395 & ~x421 & ~x445 & ~x446 & ~x475 & ~x477 & ~x479 & ~x500 & ~x505 & ~x506 & ~x527 & ~x529 & ~x531 & ~x556 & ~x562 & ~x582 & ~x583 & ~x584 & ~x586 & ~x594 & ~x611 & ~x612 & ~x614 & ~x615 & ~x618 & ~x641 & ~x666 & ~x667 & ~x672 & ~x695 & ~x696 & ~x700 & ~x702 & ~x726 & ~x730 & ~x752 & ~x755 & ~x759 & ~x760 & ~x780;
assign c0406 = ~x507 & ~x556 & ~x557 & ~x584 & ~x645 & ~x709 & ~x723 & ~x733 & ~x734 & ~x741 & ~x742 & ~x743 & ~x744 & ~x762 & ~x766 & ~x768 & ~x772 & ~x783;
assign c0408 =  x127 &  x208 &  x241 &  x269 &  x319 &  x348 &  x349 &  x350 &  x377 &  x403 &  x435 &  x465 &  x489 &  x490 &  x541 &  x548 &  x602 &  x625 &  x716 &  x771 & ~x51 & ~x57 & ~x81 & ~x87 & ~x163 & ~x172 & ~x253 & ~x303 & ~x308 & ~x310 & ~x385 & ~x390 & ~x416 & ~x419 & ~x501 & ~x504 & ~x558 & ~x559 & ~x583 & ~x590 & ~x620 & ~x643 & ~x675 & ~x696 & ~x698 & ~x750 & ~x779;
assign c0410 =  x46 &  x76 &  x77 &  x245 & ~x0 & ~x1 & ~x2 & ~x3 & ~x4 & ~x5 & ~x6 & ~x22 & ~x23 & ~x24 & ~x25 & ~x26 & ~x27 & ~x28 & ~x29 & ~x30 & ~x31 & ~x56 & ~x57 & ~x58 & ~x83 & ~x85 & ~x113 & ~x139 & ~x140 & ~x141 & ~x168 & ~x195 & ~x196 & ~x198 & ~x252 & ~x253 & ~x278 & ~x279 & ~x281 & ~x306 & ~x307 & ~x308 & ~x309 & ~x336 & ~x339 & ~x362 & ~x365 & ~x366 & ~x391 & ~x392 & ~x393 & ~x418 & ~x420 & ~x422 & ~x448 & ~x502 & ~x503 & ~x531 & ~x533 & ~x559 & ~x586 & ~x588 & ~x616 & ~x617 & ~x618 & ~x668 & ~x673 & ~x674 & ~x696 & ~x700 & ~x702 & ~x724 & ~x729 & ~x753 & ~x755 & ~x756 & ~x758 & ~x777 & ~x779 & ~x781 & ~x782;
assign c0412 =  x289 &  x298 &  x607 &  x628 &  x653 & ~x3 & ~x110 & ~x190 & ~x191 & ~x199 & ~x279 & ~x362 & ~x371 & ~x478 & ~x483 & ~x565 & ~x589 & ~x594 & ~x618 & ~x730 & ~x753;
assign c0414 =  x115;
assign c0416 =  x229 &  x230 &  x332 &  x359 &  x360 & ~x2 & ~x4 & ~x29 & ~x166 & ~x222 & ~x252 & ~x559 & ~x730 & ~x783;
assign c0418 =  x310;
assign c0420 =  x550 &  x624 &  x764 &  x774 & ~x195 & ~x252 & ~x554 & ~x559 & ~x587 & ~x610;
assign c0422 =  x274 &  x288 &  x318 &  x402 &  x574 &  x624 &  x635 &  x735 & ~x390 & ~x587 & ~x646 & ~x703 & ~x728;
assign c0424 =  x580 &  x608 &  x693 &  x720 &  x722 & ~x13 & ~x14 & ~x28;
assign c0426 = ~x5 & ~x74 & ~x102 & ~x197 & ~x226 & ~x254 & ~x306 & ~x336 & ~x384 & ~x387 & ~x388 & ~x392 & ~x396 & ~x412 & ~x414 & ~x415 & ~x421 & ~x451 & ~x497 & ~x504 & ~x525 & ~x553 & ~x563 & ~x580 & ~x609 & ~x620 & ~x636 & ~x664 & ~x666 & ~x751;
assign c0428 =  x38 &  x102 &  x523 &  x541 &  x596 &  x606 &  x629 &  x633 &  x663 &  x709 &  x710 &  x737 &  x742 &  x745 & ~x1 & ~x3 & ~x26 & ~x27 & ~x29 & ~x31 & ~x51 & ~x56 & ~x83 & ~x84 & ~x85 & ~x86 & ~x143 & ~x170 & ~x196 & ~x224 & ~x252 & ~x278 & ~x279 & ~x280 & ~x306 & ~x308 & ~x309 & ~x335 & ~x337 & ~x365 & ~x390 & ~x392 & ~x393 & ~x418 & ~x419 & ~x421 & ~x504 & ~x525 & ~x531 & ~x532 & ~x533 & ~x560 & ~x588 & ~x675 & ~x700 & ~x701 & ~x726 & ~x729 & ~x731 & ~x732 & ~x733 & ~x753 & ~x755 & ~x760;
assign c0430 =  x354 &  x607 &  x630 & ~x1 & ~x140 & ~x147 & ~x307 & ~x483 & ~x525 & ~x588 & ~x706;
assign c0432 =  x510 &  x654 &  x706 &  x708 & ~x11 & ~x12 & ~x13;
assign c0434 = ~x15 & ~x60 & ~x280 & ~x281 & ~x307 & ~x308 & ~x362 & ~x371 & ~x447 & ~x558 & ~x584 & ~x590 & ~x686 & ~x687 & ~x703;
assign c0436 =  x205 &  x263 &  x271 &  x289 &  x292 &  x298 &  x299 &  x402 &  x435 &  x463 &  x490 &  x495 &  x521 &  x522 &  x542 &  x545 &  x547 &  x574 &  x602 &  x605 &  x606 &  x607 &  x627 &  x630 &  x656 &  x658 & ~x0 & ~x6 & ~x21 & ~x22 & ~x135 & ~x139 & ~x141 & ~x142 & ~x146 & ~x168 & ~x172 & ~x173 & ~x196 & ~x306 & ~x312 & ~x417 & ~x453 & ~x477 & ~x535 & ~x557 & ~x589 & ~x620 & ~x645 & ~x700 & ~x755;
assign c0438 =  x39 &  x229 &  x572 &  x603 &  x625 &  x653 &  x743 & ~x0 & ~x3 & ~x31 & ~x51 & ~x54 & ~x109 & ~x114 & ~x167 & ~x169 & ~x197 & ~x281 & ~x311 & ~x361 & ~x364 & ~x474 & ~x476 & ~x501 & ~x506 & ~x558 & ~x560 & ~x614 & ~x615 & ~x649 & ~x666 & ~x667 & ~x673 & ~x676 & ~x697 & ~x703 & ~x724 & ~x728 & ~x730 & ~x731 & ~x732 & ~x751 & ~x752 & ~x754 & ~x759 & ~x761 & ~x782;
assign c0440 =  x44 &  x457 &  x597 & ~x3 & ~x20 & ~x54 & ~x56 & ~x59 & ~x112 & ~x170 & ~x225 & ~x244 & ~x306 & ~x333 & ~x447 & ~x526 & ~x529 & ~x534 & ~x566 & ~x586 & ~x590 & ~x615 & ~x618 & ~x638 & ~x650 & ~x667 & ~x704 & ~x755;
assign c0442 =  x177 &  x268 &  x270 &  x573 &  x630 & ~x7 & ~x91 & ~x115 & ~x147 & ~x224 & ~x338 & ~x387 & ~x727 & ~x782;
assign c0444 =  x191 &  x411 &  x579 &  x603 &  x662 &  x719 &  x720 & ~x50 & ~x109 & ~x167 & ~x391 & ~x534 & ~x559 & ~x587 & ~x676 & ~x757 & ~x780;
assign c0446 =  x96 &  x97 &  x99 & ~x111 & ~x239 & ~x447 & ~x614 & ~x724;
assign c0448 =  x624 &  x659 &  x717 &  x774 & ~x76;
assign c0450 =  x229 &  x247 &  x255 &  x256 &  x283 & ~x56 & ~x85 & ~x756;
assign c0452 =  x229 &  x513 &  x519 &  x655 &  x656 & ~x2 & ~x5 & ~x56 & ~x57 & ~x60 & ~x80 & ~x85 & ~x88 & ~x139 & ~x143 & ~x167 & ~x195 & ~x223 & ~x251 & ~x279 & ~x363 & ~x477 & ~x479 & ~x500 & ~x503 & ~x504 & ~x508 & ~x554 & ~x560 & ~x562 & ~x586 & ~x611 & ~x619 & ~x621 & ~x643 & ~x695 & ~x699 & ~x704 & ~x706 & ~x733 & ~x751 & ~x755 & ~x781 & ~x782;
assign c0454 =  x130 &  x210 &  x322 &  x325 &  x345 &  x430 &  x546 &  x602 &  x657 &  x689 & ~x20 & ~x134 & ~x197 & ~x198 & ~x230 & ~x286 & ~x302 & ~x341 & ~x342 & ~x385 & ~x417 & ~x422 & ~x501 & ~x560 & ~x668 & ~x703 & ~x757;
assign c0456 =  x45 & ~x353;
assign c0458 =  x369 &  x471 &  x508 &  x708 & ~x196;
assign c0460 = ~x293 & ~x483 & ~x597 & ~x709;
assign c0462 = ~x344 & ~x362 & ~x469 & ~x525 & ~x564 & ~x667 & ~x711 & ~x713;
assign c0464 = ~x471 & ~x632 & ~x633 & ~x634 & ~x686 & ~x722 & ~x750;
assign c0466 =  x595 &  x707 &  x708 & ~x4 & ~x12 & ~x13 & ~x15 & ~x41 & ~x43 & ~x54 & ~x58 & ~x110 & ~x335 & ~x588;
assign c0470 = ~x686;
assign c0472 =  x243 &  x289 &  x294 &  x355 &  x378 &  x401 &  x430 &  x432 &  x433 &  x437 &  x464 &  x494 &  x518 &  x519 &  x522 &  x569 &  x603 &  x607 &  x634 &  x635 &  x655 &  x658 &  x662 &  x681 &  x685 &  x690 &  x713 & ~x4 & ~x21 & ~x22 & ~x50 & ~x56 & ~x81 & ~x83 & ~x84 & ~x86 & ~x87 & ~x111 & ~x113 & ~x137 & ~x138 & ~x139 & ~x140 & ~x168 & ~x195 & ~x226 & ~x252 & ~x308 & ~x343 & ~x360 & ~x421 & ~x446 & ~x474 & ~x476 & ~x478 & ~x504 & ~x507 & ~x529 & ~x534 & ~x537 & ~x555 & ~x557 & ~x562 & ~x588 & ~x593 & ~x648 & ~x672 & ~x674 & ~x676 & ~x703 & ~x723 & ~x732 & ~x759 & ~x761 & ~x779;
assign c0474 =  x125 &  x126 &  x152 &  x178 &  x205 &  x209 &  x299 &  x346 &  x355 &  x401 &  x406 &  x514 &  x572 &  x578 &  x603 &  x607 &  x625 &  x691 &  x713 & ~x32 & ~x114 & ~x171 & ~x227 & ~x253 & ~x279 & ~x335 & ~x363 & ~x455 & ~x469 & ~x475 & ~x537 & ~x566 & ~x667 & ~x671 & ~x675 & ~x729;
assign c0476 =  x142;
assign c0478 =  x543 &  x567 &  x623 &  x710 & ~x12 & ~x15 & ~x41 & ~x42 & ~x55 & ~x57 & ~x85 & ~x420 & ~x671 & ~x729;
assign c0480 = ~x139 & ~x166 & ~x320 & ~x322 & ~x454 & ~x471 & ~x477 & ~x509 & ~x528 & ~x535 & ~x555 & ~x558 & ~x560 & ~x564 & ~x582 & ~x585 & ~x589 & ~x621 & ~x638 & ~x650 & ~x667 & ~x703 & ~x723 & ~x751 & ~x752 & ~x762;
assign c0482 =  x171;
assign c0484 =  x483 &  x539 &  x596 &  x624 &  x656 &  x657 &  x685 &  x707 &  x712 & ~x11 & ~x13 & ~x14 & ~x26 & ~x55 & ~x111 & ~x168 & ~x308 & ~x309 & ~x333 & ~x393 & ~x422 & ~x446 & ~x532 & ~x533 & ~x558 & ~x561 & ~x586 & ~x587 & ~x672 & ~x727 & ~x754 & ~x755 & ~x758;
assign c0486 =  x220 &  x341 & ~x5 & ~x85 & ~x364;
assign c0488 = ~x164 & ~x384 & ~x525 & ~x553 & ~x590 & ~x618 & ~x631 & ~x633 & ~x635 & ~x637 & ~x638 & ~x732;
assign c0490 =  x312 & ~x10 & ~x11 & ~x12 & ~x16 & ~x84 & ~x278 & ~x280 & ~x756;
assign c0492 =  x41 &  x43 &  x768 &  x769 &  x773 &  x774 & ~x0 & ~x53 & ~x57 & ~x84 & ~x111 & ~x113 & ~x169 & ~x197 & ~x223 & ~x251 & ~x252 & ~x309 & ~x337 & ~x392 & ~x449 & ~x474 & ~x478 & ~x503 & ~x505 & ~x532 & ~x559 & ~x562 & ~x588 & ~x638 & ~x643 & ~x649 & ~x675 & ~x698 & ~x701 & ~x702 & ~x703 & ~x704 & ~x780 & ~x781;
assign c0494 =  x735 & ~x5 & ~x27 & ~x94;
assign c0496 =  x105 &  x126 &  x343 &  x596 & ~x3 & ~x88 & ~x363 & ~x648 & ~x699;
assign c0498 = ~x456 & ~x598 & ~x601;
assign c01 =  x26;
assign c03 =  x252;
assign c05 =  x42 &  x123 &  x711 & ~x6 & ~x77 & ~x84 & ~x89 & ~x142 & ~x163 & ~x191 & ~x201 & ~x285 & ~x303 & ~x446 & ~x451 & ~x505 & ~x564 & ~x693 & ~x721;
assign c07 =  x392;
assign c09 = ~x17 & ~x95 & ~x152 & ~x742;
assign c011 =  x504;
assign c013 = ~x94 & ~x680 & ~x717;
assign c015 =  x224;
assign c017 =  x555 & ~x134;
assign c019 =  x43 &  x723;
assign c021 =  x141;
assign c023 =  x148 &  x681 & ~x25 & ~x78 & ~x117 & ~x173 & ~x192 & ~x310 & ~x363 & ~x533 & ~x619 & ~x665 & ~x707;
assign c025 =  x756;
assign c027 =  x1;
assign c029 =  x195;
assign c031 =  x279;
assign c033 =  x37 &  x74 &  x129 &  x178 &  x179 &  x182 &  x213 &  x235 &  x270 &  x295 &  x296 &  x352 &  x379 &  x407 &  x429 &  x458 &  x466 &  x468 &  x496 &  x551 &  x552 &  x576 &  x599 & ~x23 & ~x30 & ~x32 & ~x56 & ~x87 & ~x137 & ~x198 & ~x221 & ~x277 & ~x333 & ~x535 & ~x558 & ~x641 & ~x728 & ~x756 & ~x777 & ~x783;
assign c037 =  x51;
assign c039 =  x44 &  x237 &  x372 &  x384 & ~x108 & ~x228 & ~x254 & ~x275 & ~x276;
assign c041 =  x180 &  x211 &  x239 &  x295 &  x711 &  x712 &  x719 & ~x173 & ~x256 & ~x344 & ~x442;
assign c043 = ~x201 & ~x256 & ~x434 & ~x630;
assign c045 =  x746 & ~x284 & ~x287 & ~x299 & ~x443;
assign c047 =  x723;
assign c049 =  x307;
assign c051 =  x45 &  x694 &  x705;
assign c053 =  x420;
assign c055 = ~x1 & ~x3 & ~x11 & ~x16 & ~x36 & ~x46 & ~x47 & ~x63 & ~x76 & ~x161 & ~x189 & ~x191 & ~x199 & ~x201 & ~x245 & ~x276 & ~x282 & ~x310 & ~x673;
assign c057 =  x13 & ~x77 & ~x174 & ~x312;
assign c059 =  x40 & ~x1 & ~x2 & ~x25 & ~x26 & ~x29 & ~x33 & ~x51 & ~x52 & ~x56 & ~x58 & ~x59 & ~x62 & ~x77 & ~x79 & ~x81 & ~x82 & ~x85 & ~x87 & ~x88 & ~x90 & ~x105 & ~x106 & ~x107 & ~x109 & ~x111 & ~x113 & ~x115 & ~x116 & ~x118 & ~x134 & ~x135 & ~x137 & ~x138 & ~x139 & ~x143 & ~x145 & ~x163 & ~x164 & ~x165 & ~x168 & ~x169 & ~x172 & ~x173 & ~x191 & ~x196 & ~x199 & ~x200 & ~x224 & ~x226 & ~x229 & ~x247 & ~x248 & ~x250 & ~x252 & ~x256 & ~x274 & ~x275 & ~x278 & ~x279 & ~x282 & ~x284 & ~x285 & ~x304 & ~x305 & ~x306 & ~x311 & ~x331 & ~x332 & ~x333 & ~x336 & ~x337 & ~x340 & ~x360 & ~x361 & ~x362 & ~x363 & ~x364 & ~x367 & ~x368 & ~x387 & ~x389 & ~x392 & ~x393 & ~x395 & ~x396 & ~x415 & ~x416 & ~x418 & ~x422 & ~x424 & ~x444 & ~x445 & ~x446 & ~x447 & ~x448 & ~x451 & ~x452 & ~x471 & ~x474 & ~x479 & ~x500 & ~x501 & ~x506 & ~x531 & ~x533 & ~x535 & ~x559 & ~x560 & ~x563 & ~x586 & ~x589 & ~x590 & ~x618 & ~x639 & ~x640 & ~x642 & ~x643 & ~x644 & ~x645 & ~x646 & ~x647 & ~x671 & ~x673 & ~x674 & ~x675 & ~x698 & ~x700 & ~x703 & ~x704 & ~x727 & ~x728 & ~x729 & ~x730 & ~x753 & ~x756 & ~x757 & ~x758 & ~x764 & ~x765 & ~x779 & ~x782;
assign c061 =  x279;
assign c063 =  x41 &  x131 &  x158 &  x211 &  x267 &  x270 &  x292 &  x430 &  x436 &  x466 &  x495 &  x542 &  x569 &  x577 &  x606 &  x717 & ~x26 & ~x50 & ~x79 & ~x82 & ~x87 & ~x116 & ~x117 & ~x139 & ~x165 & ~x220 & ~x223 & ~x224 & ~x226 & ~x278 & ~x280 & ~x310 & ~x333 & ~x360 & ~x361 & ~x387 & ~x388 & ~x424 & ~x449 & ~x451 & ~x474 & ~x501 & ~x504 & ~x527 & ~x586 & ~x588 & ~x616 & ~x617 & ~x647 & ~x667 & ~x672 & ~x674 & ~x699 & ~x722 & ~x777 & ~x778;
assign c065 =  x280;
assign c067 =  x85;
assign c069 =  x755;
assign c071 =  x307;
assign c073 =  x29;
assign c075 =  x443 &  x677;
assign c077 =  x783;
assign c079 =  x122 &  x239 &  x263 &  x268 &  x350 &  x375 &  x382 &  x437 &  x487 &  x521 &  x551 &  x599 &  x627 &  x632 &  x633 &  x716 &  x736 & ~x59 & ~x79 & ~x86 & ~x111 & ~x116 & ~x143 & ~x163 & ~x167 & ~x225 & ~x228 & ~x255 & ~x257 & ~x281 & ~x285 & ~x303 & ~x304 & ~x340 & ~x418 & ~x504 & ~x562 & ~x593 & ~x611 & ~x619 & ~x621 & ~x677 & ~x696 & ~x704 & ~x754 & ~x759 & ~x763 & ~x781;
assign c081 =  x158 &  x292 &  x745 & ~x145 & ~x167 & ~x248 & ~x623;
assign c083 = ~x65 & ~x122 & ~x232 & ~x261;
assign c085 =  x588;
assign c087 =  x42 &  x98 &  x209 &  x237 & ~x145 & ~x218;
assign c089 = ~x402 & ~x493;
assign c091 = ~x275 & ~x406 & ~x434 & ~x574;
assign c093 =  x196;
assign c095 =  x391;
assign c097 = ~x43 & ~x96 & ~x123 & ~x233 & ~x235;
assign c099 =  x59;
assign c0101 = ~x11 & ~x47 & ~x144 & ~x204 & ~x232 & ~x313 & ~x341 & ~x722;
assign c0103 =  x296 &  x371 &  x479 &  x525 &  x538 &  x566;
assign c0105 =  x292 &  x739 & ~x144 & ~x201 & ~x256 & ~x277 & ~x532 & ~x651 & ~x678;
assign c0107 =  x738 & ~x7 & ~x48 & ~x90 & ~x115 & ~x138 & ~x163 & ~x531 & ~x587 & ~x636 & ~x651 & ~x724 & ~x748 & ~x776;
assign c0109 =  x757;
assign c0111 =  x154 &  x464 & ~x90 & ~x162 & ~x285 & ~x623;
assign c0113 =  x782;
assign c0115 =  x224;
assign c0117 = ~x261 & ~x289 & ~x683;
assign c0119 =  x731;
assign c0121 =  x41 &  x68 &  x291 &  x318 &  x404 &  x410 &  x466 &  x579 &  x598 &  x688 & ~x9 & ~x24 & ~x32 & ~x49 & ~x54 & ~x106 & ~x113 & ~x137 & ~x163 & ~x227 & ~x248 & ~x251 & ~x282 & ~x283 & ~x368 & ~x418 & ~x559 & ~x700 & ~x723 & ~x728;
assign c0123 =  x412 & ~x9 & ~x36 & ~x49 & ~x201 & ~x227 & ~x367;
assign c0125 =  x1;
assign c0127 =  x675 & ~x540;
assign c0129 =  x56;
assign c0131 =  x23;
assign c0133 =  x279;
assign c0135 =  x759;
assign c0137 =  x363;
assign c0139 =  x632 & ~x133 & ~x623 & ~x664;
assign c0141 =  x711 & ~x145 & ~x258 & ~x260 & ~x271;
assign c0143 =  x97 &  x179 &  x207 &  x213 &  x238 &  x325 &  x400 &  x466 &  x550 &  x663 & ~x33 & ~x34 & ~x35 & ~x49 & ~x54 & ~x89 & ~x111 & ~x164 & ~x254 & ~x278 & ~x338 & ~x340 & ~x393 & ~x560 & ~x584 & ~x616 & ~x722 & ~x723 & ~x728 & ~x729;
assign c0145 =  x181 &  x404 &  x717 & ~x110 & ~x162 & ~x201 & ~x608 & ~x637;
assign c0147 =  x123 &  x128 &  x152 &  x185 &  x241 &  x265 &  x319 &  x324 &  x379 &  x402 &  x407 &  x431 &  x460 &  x466 &  x494 &  x513 &  x541 &  x547 &  x577 &  x599 &  x605 &  x625 &  x655 &  x660 &  x688 &  x737 & ~x6 & ~x26 & ~x29 & ~x50 & ~x57 & ~x81 & ~x83 & ~x84 & ~x85 & ~x87 & ~x113 & ~x115 & ~x134 & ~x144 & ~x163 & ~x164 & ~x166 & ~x168 & ~x169 & ~x171 & ~x172 & ~x173 & ~x195 & ~x197 & ~x223 & ~x228 & ~x253 & ~x255 & ~x277 & ~x278 & ~x279 & ~x303 & ~x305 & ~x308 & ~x309 & ~x313 & ~x332 & ~x334 & ~x338 & ~x339 & ~x364 & ~x366 & ~x368 & ~x388 & ~x395 & ~x447 & ~x448 & ~x478 & ~x504 & ~x528 & ~x529 & ~x533 & ~x534 & ~x535 & ~x556 & ~x561 & ~x586 & ~x587 & ~x589 & ~x641 & ~x646 & ~x647 & ~x649 & ~x697 & ~x701 & ~x704 & ~x705 & ~x723 & ~x725 & ~x730 & ~x752 & ~x753 & ~x756 & ~x757 & ~x762 & ~x778;
assign c0149 =  x559;
assign c0151 = ~x41 & ~x69 & ~x71 & ~x315;
assign c0153 =  x26;
assign c0155 = ~x134 & ~x743;
assign c0157 =  x384 & ~x90 & ~x161 & ~x331;
assign c0159 =  x675;
assign c0161 =  x84;
assign c0163 =  x237 &  x403 &  x632 &  x744 &  x746 & ~x26 & ~x35 & ~x54 & ~x106 & ~x168 & ~x172 & ~x191 & ~x250 & ~x276 & ~x334 & ~x335 & ~x336 & ~x341 & ~x499 & ~x500 & ~x504 & ~x509 & ~x641 & ~x693 & ~x758;
assign c0165 = ~x77 & ~x80 & ~x163 & ~x218 & ~x368 & ~x623 & ~x680 & ~x735 & ~x763;
assign c0167 =  x782;
assign c0169 =  x29;
assign c0171 =  x111;
assign c0173 = ~x187 & ~x216 & ~x271 & ~x288;
assign c0175 =  x343 &  x344 & ~x62 & ~x338 & ~x736 & ~x764;
assign c0177 =  x391;
assign c0179 = ~x45 & ~x202 & ~x666;
assign c0181 =  x210 &  x324 &  x711 &  x740 & ~x77 & ~x218;
assign c0183 =  x73 &  x123 &  x209 & ~x90 & ~x104 & ~x117 & ~x118 & ~x135 & ~x255 & ~x284 & ~x359;
assign c0185 =  x588;
assign c0187 =  x230 &  x240 &  x296 &  x351 &  x413 &  x425 &  x466 &  x482 &  x511 & ~x762;
assign c0189 = ~x429 & ~x690;
assign c0191 =  x26;
assign c0193 =  x709 & ~x145 & ~x229 & ~x232 & ~x257 & ~x260 & ~x271 & ~x287;
assign c0195 =  x112;
assign c0197 =  x65 &  x67 &  x94 &  x95 &  x127 &  x128 &  x207 &  x231 &  x238 &  x240 &  x267 &  x381 &  x402 &  x403 &  x407 &  x409 &  x432 &  x433 &  x439 &  x464 &  x494 &  x544 &  x598 &  x603 &  x604 &  x605 &  x635 &  x746 & ~x30 & ~x111 & ~x142 & ~x144 & ~x165 & ~x192 & ~x221 & ~x281 & ~x363 & ~x394 & ~x395 & ~x477 & ~x502 & ~x587 & ~x590 & ~x643 & ~x670 & ~x699 & ~x776;
assign c0199 =  x111;
assign c0201 =  x235 &  x273 &  x371 &  x380 &  x440 &  x469 &  x470 &  x482 &  x483 &  x566 & ~x762;
assign c0203 =  x620 & ~x738;
assign c0205 =  x40 &  x676;
assign c0207 =  x363;
assign c0209 =  x555 &  x610 & ~x8;
assign c0211 =  x57;
assign c0213 =  x783;
assign c0215 =  x717 & ~x224 & ~x246 & ~x423 & ~x679 & ~x692 & ~x698 & ~x779;
assign c0217 = ~x46 & ~x76 & ~x179 & ~x184 & ~x208 & ~x262;
assign c0219 = ~x87 & ~x175 & ~x202 & ~x204 & ~x215 & ~x218 & ~x229 & ~x244 & ~x247 & ~x248 & ~x273 & ~x275 & ~x287 & ~x302 & ~x314;
assign c0221 =  x430 & ~x163 & ~x244 & ~x260 & ~x300 & ~x329 & ~x344;
assign c0225 =  x41 &  x66 &  x182 & ~x1 & ~x4 & ~x22 & ~x23 & ~x26 & ~x27 & ~x28 & ~x29 & ~x30 & ~x32 & ~x49 & ~x58 & ~x59 & ~x76 & ~x78 & ~x79 & ~x82 & ~x84 & ~x86 & ~x88 & ~x89 & ~x108 & ~x111 & ~x112 & ~x135 & ~x136 & ~x137 & ~x138 & ~x143 & ~x163 & ~x165 & ~x168 & ~x169 & ~x170 & ~x192 & ~x193 & ~x197 & ~x220 & ~x221 & ~x222 & ~x225 & ~x227 & ~x248 & ~x250 & ~x253 & ~x276 & ~x277 & ~x278 & ~x279 & ~x282 & ~x305 & ~x308 & ~x310 & ~x359 & ~x364 & ~x365 & ~x366 & ~x393 & ~x396 & ~x417 & ~x420 & ~x422 & ~x445 & ~x447 & ~x473 & ~x479 & ~x505 & ~x529 & ~x530 & ~x531 & ~x533 & ~x557 & ~x558 & ~x563 & ~x589 & ~x591 & ~x615 & ~x616 & ~x617 & ~x619 & ~x640 & ~x643 & ~x644 & ~x645 & ~x669 & ~x671 & ~x672 & ~x674 & ~x698 & ~x699 & ~x700 & ~x702 & ~x703 & ~x725 & ~x727 & ~x729 & ~x753 & ~x754 & ~x757 & ~x760 & ~x775 & ~x779 & ~x780 & ~x783;
assign c0227 =  x28;
assign c0229 =  x534;
assign c0233 =  x356 &  x375 &  x408 &  x508 & ~x136 & ~x670;
assign c0235 =  x39 &  x155 &  x182 &  x208 &  x211 & ~x146 & ~x190 & ~x331;
assign c0237 = ~x273 & ~x720;
assign c0239 =  x727;
assign c0243 =  x103 & ~x35 & ~x78 & ~x106 & ~x145 & ~x251 & ~x499 & ~x529 & ~x535 & ~x650 & ~x678 & ~x693 & ~x725 & ~x734 & ~x749;
assign c0245 =  x186 &  x740 & ~x48 & ~x735 & ~x748;
assign c0247 = ~x46 & ~x267 & ~x313;
assign c0249 =  x16 &  x648;
assign c0251 =  x380 &  x413 &  x468 &  x524 &  x527 & ~x23 & ~x136 & ~x673;
assign c0253 =  x67 &  x73 &  x128 &  x182 &  x431 & ~x36 & ~x63 & ~x77 & ~x144 & ~x202 & ~x340 & ~x503;
assign c0255 =  x525 & ~x20 & ~x24 & ~x35 & ~x48 & ~x49 & ~x59 & ~x77 & ~x78 & ~x79 & ~x107 & ~x117 & ~x139 & ~x143 & ~x249 & ~x256 & ~x276 & ~x303 & ~x331 & ~x447 & ~x675 & ~x727 & ~x753 & ~x756;
assign c0257 =  x195;
assign c0259 =  x5;
assign c0261 =  x296 &  x357 &  x412 &  x468 &  x472 &  x496 & ~x778;
assign c0263 =  x729;
assign c0265 =  x39 &  x72 &  x96 &  x128 &  x182 &  x183 &  x207 &  x208 &  x213 &  x264 &  x348 &  x515 &  x576 & ~x5 & ~x19 & ~x29 & ~x30 & ~x50 & ~x139 & ~x141 & ~x143 & ~x221 & ~x248 & ~x276 & ~x303 & ~x304 & ~x310 & ~x312 & ~x338 & ~x366 & ~x391 & ~x395 & ~x474 & ~x535 & ~x563 & ~x640 & ~x779;
assign c0267 =  x15 & ~x77 & ~x172 & ~x200 & ~x201 & ~x391;
assign c0269 =  x27;
assign c0271 =  x140;
assign c0273 =  x279;
assign c0275 =  x29;
assign c0277 =  x42 &  x208 &  x324 &  x748 & ~x9 & ~x27 & ~x33 & ~x87 & ~x141 & ~x163 & ~x164 & ~x198 & ~x199 & ~x220 & ~x277 & ~x310 & ~x338 & ~x361 & ~x561;
assign c0279 =  x534;
assign c0281 =  x113;
assign c0283 = ~x77 & ~x176 & ~x268;
assign c0285 =  x334;
assign c0287 =  x167;
assign c0289 =  x40 &  x72 &  x148 &  x209 &  x352 &  x438 &  x626 &  x690 &  x709 & ~x227 & ~x303 & ~x312 & ~x331 & ~x452 & ~x700 & ~x706;
assign c0291 =  x76 &  x709 & ~x14 & ~x144 & ~x191 & ~x305 & ~x312 & ~x332 & ~x526 & ~x593;
assign c0293 =  x588;
assign c0295 = ~x20 & ~x135 & ~x176 & ~x200 & ~x230 & ~x231 & ~x271 & ~x272 & ~x283 & ~x285 & ~x287 & ~x315;
assign c0297 =  x372 &  x400 & ~x11 & ~x19 & ~x23 & ~x47 & ~x48 & ~x49 & ~x51 & ~x76 & ~x89 & ~x105 & ~x136 & ~x163 & ~x254 & ~x255 & ~x278 & ~x335 & ~x418 & ~x558 & ~x559 & ~x615 & ~x674 & ~x781;
assign c0299 = ~x292 & ~x551;
assign c0301 =  x166;
assign c0303 =  x727;
assign c0305 = ~x16 & ~x47 & ~x48 & ~x49 & ~x176 & ~x189 & ~x274 & ~x277 & ~x305 & ~x613;
assign c0307 =  x666 &  x677;
assign c0309 = ~x11 & ~x35 & ~x46 & ~x285 & ~x717;
assign c0311 = ~x144 & ~x230 & ~x243 & ~x246 & ~x259 & ~x260 & ~x271 & ~x273 & ~x330 & ~x414 & ~x443 & ~x780;
assign c0313 =  x728;
assign c0315 =  x504;
assign c0317 = ~x77 & ~x144 & ~x286 & ~x326 & ~x330 & ~x457;
assign c0319 =  x196;
assign c0321 =  x421;
assign c0323 =  x560;
assign c0325 = ~x191 & ~x227 & ~x228 & ~x518 & ~x574 & ~x742;
assign c0327 =  x65 &  x71 &  x72 &  x73 &  x74 &  x127 &  x263 &  x320 &  x323 &  x404 &  x407 &  x430 &  x437 &  x488 &  x521 &  x661 &  x682 &  x683 & ~x136 & ~x139 & ~x168 & ~x193 & ~x219 & ~x220 & ~x221 & ~x222 & ~x253 & ~x283 & ~x331 & ~x339 & ~x392 & ~x396 & ~x420 & ~x446 & ~x452 & ~x508 & ~x534 & ~x589 & ~x614 & ~x675 & ~x677 & ~x698 & ~x706 & ~x730 & ~x731 & ~x733;
assign c0329 = ~x16 & ~x71 & ~x233 & ~x260;
assign c0331 =  x726;
assign c0333 =  x477;
assign c0335 =  x588;
assign c0337 =  x739 & ~x64 & ~x736;
assign c0339 =  x72 &  x73 &  x94 &  x95 &  x97 &  x132 &  x154 &  x183 &  x211 &  x237 &  x263 &  x403 &  x435 &  x438 &  x542 &  x577 &  x627 &  x681 &  x684 &  x711 &  x712 &  x738 & ~x28 & ~x82 & ~x110 & ~x135 & ~x144 & ~x194 & ~x197 & ~x226 & ~x280 & ~x363 & ~x397 & ~x452 & ~x476 & ~x557 & ~x592 & ~x612 & ~x666 & ~x676 & ~x699;
assign c0341 =  x40 &  x424 &  x676;
assign c0343 =  x168;
assign c0345 =  x695 & ~x108;
assign c0349 =  x756;
assign c0351 =  x278;
assign c0353 =  x84 &  x223;
assign c0355 = ~x75 & ~x245 & ~x261 & ~x287;
assign c0357 =  x112;
assign c0359 = ~x124 & ~x296 & ~x661;
assign c0361 = ~x38 & ~x260;
assign c0363 =  x57;
assign c0365 =  x757;
assign c0367 = ~x204 & ~x230 & ~x260 & ~x271 & ~x301 & ~x316 & ~x357 & ~x386;
assign c0369 =  x666 & ~x164 & ~x172 & ~x221 & ~x473 & ~x590;
assign c0371 =  x279;
assign c0373 =  x29;
assign c0375 =  x425 & ~x726 & ~x773;
assign c0377 =  x783;
assign c0381 =  x308;
assign c0383 =  x616;
assign c0385 =  x383 &  x440 &  x524 &  x566 &  x607 &  x637 & ~x19 & ~x250 & ~x335 & ~x670 & ~x701 & ~x754;
assign c0387 =  x307;
assign c0389 =  x501;
assign c0391 =  x54;
assign c0393 =  x44 & ~x9 & ~x220;
assign c0395 =  x57;
assign c0397 =  x74 &  x101 &  x160 &  x203 &  x207 &  x351 &  x374 &  x408 &  x436 &  x464 &  x488 &  x551 &  x572 &  x603 &  x604 & ~x30 & ~x52 & ~x53 & ~x142 & ~x200 & ~x249 & ~x250 & ~x284 & ~x308 & ~x333 & ~x339 & ~x362 & ~x419 & ~x528 & ~x585 & ~x586 & ~x725 & ~x762 & ~x777 & ~x782;
assign c0399 =  x584;
assign c0401 =  x757;
assign c0403 =  x26;
assign c0405 =  x616;
assign c0407 =  x643;
assign c0409 =  x56;
assign c0411 = ~x204 & ~x242 & ~x256;
assign c0413 =  x113;
assign c0415 =  x223;
assign c0417 =  x593 & ~x172;
assign c0419 =  x198;
assign c0421 = ~x69 & ~x260 & ~x287;
assign c0423 =  x307;
assign c0425 = ~x76 & ~x152 & ~x548 & ~x735;
assign c0427 =  x505;
assign c0429 =  x361 &  x413;
assign c0433 =  x422;
assign c0435 =  x364;
assign c0437 =  x28;
assign c0439 =  x67 &  x71 &  x73 &  x74 &  x95 &  x102 &  x131 &  x213 &  x264 &  x381 &  x521 &  x718 & ~x2 & ~x26 & ~x59 & ~x60 & ~x77 & ~x85 & ~x86 & ~x198 & ~x249 & ~x340 & ~x387 & ~x390 & ~x391 & ~x422 & ~x450 & ~x452 & ~x473 & ~x506 & ~x531 & ~x534 & ~x557 & ~x562 & ~x648 & ~x675 & ~x695 & ~x697 & ~x732 & ~x778;
assign c0441 =  x271 &  x416 & ~x701;
assign c0443 =  x92 &  x212 &  x322 &  x376 &  x381 &  x466 &  x709 &  x717 & ~x2 & ~x23 & ~x90 & ~x112 & ~x113 & ~x170 & ~x191 & ~x309 & ~x446 & ~x620 & ~x666 & ~x667 & ~x671 & ~x694 & ~x724 & ~x778;
assign c0445 = ~x2 & ~x3 & ~x6 & ~x8 & ~x11 & ~x17 & ~x20 & ~x31 & ~x33 & ~x35 & ~x36 & ~x47 & ~x48 & ~x56 & ~x59 & ~x61 & ~x76 & ~x82 & ~x85 & ~x88 & ~x89 & ~x90 & ~x104 & ~x105 & ~x106 & ~x110 & ~x116 & ~x135 & ~x136 & ~x142 & ~x144 & ~x145 & ~x162 & ~x163 & ~x164 & ~x172 & ~x174 & ~x198 & ~x200 & ~x201 & ~x219 & ~x221 & ~x222 & ~x251 & ~x256 & ~x334 & ~x337 & ~x449 & ~x532 & ~x563 & ~x613 & ~x614 & ~x643 & ~x646 & ~x700 & ~x751 & ~x757;
assign c0447 =  x102 &  x745 & ~x106 & ~x170 & ~x190 & ~x679;
assign c0449 =  x587;
assign c0451 =  x57;
assign c0453 =  x112;
assign c0455 =  x42 &  x95 &  x356 &  x438 & ~x78 & ~x79 & ~x80 & ~x82 & ~x106 & ~x108 & ~x191 & ~x221 & ~x337 & ~x366 & ~x473 & ~x560 & ~x614 & ~x640 & ~x645 & ~x698 & ~x726;
assign c0457 =  x758;
assign c0459 =  x55;
assign c0461 =  x222;
assign c0463 =  x503;
assign c0465 =  x676 & ~x762;
assign c0467 =  x758;
assign c0469 =  x538 & ~x64;
assign c0471 = ~x105 & ~x171 & ~x175 & ~x310 & ~x741;
assign c0473 =  x195;
assign c0475 = ~x163 & ~x436;
assign c0477 =  x195;
assign c0479 = ~x204 & ~x241 & ~x286 & ~x302;
assign c0481 =  x167 &  x587;
assign c0483 = ~x50 & ~x134 & ~x231 & ~x246 & ~x258 & ~x299 & ~x301 & ~x420 & ~x482 & ~x586 & ~x612;
assign c0485 =  x280;
assign c0487 = ~x99 & ~x179 & ~x599 & ~x744;
assign c0489 =  x128 &  x571 & ~x115 & ~x216 & ~x230 & ~x244 & ~x272;
assign c0491 =  x42 &  x399 &  x400 & ~x77 & ~x90 & ~x106;
assign c0493 =  x440 &  x441 &  x537 & ~x9;
assign c0497 =  x258 &  x324 &  x342 &  x372 &  x380 &  x386 &  x442 &  x482 &  x483 & ~x702 & ~x762;
assign c0499 =  x14 & ~x50 & ~x76 & ~x117 & ~x756;
assign c10 =  x296 &  x374 &  x457 &  x767 & ~x19 & ~x50 & ~x245 & ~x589 & ~x665;
assign c12 =  x240 &  x323 &  x348 &  x351 &  x376 &  x405 &  x491 & ~x0 & ~x2 & ~x25 & ~x26 & ~x29 & ~x30 & ~x33 & ~x35 & ~x47 & ~x48 & ~x51 & ~x54 & ~x58 & ~x62 & ~x83 & ~x87 & ~x88 & ~x104 & ~x106 & ~x108 & ~x112 & ~x115 & ~x117 & ~x133 & ~x140 & ~x141 & ~x146 & ~x159 & ~x161 & ~x164 & ~x172 & ~x187 & ~x188 & ~x197 & ~x201 & ~x226 & ~x247 & ~x253 & ~x273 & ~x274 & ~x276 & ~x279 & ~x282 & ~x285 & ~x288 & ~x308 & ~x312 & ~x327 & ~x341 & ~x360 & ~x367 & ~x368 & ~x371 & ~x372 & ~x391 & ~x397 & ~x401 & ~x417 & ~x422 & ~x429 & ~x441 & ~x442 & ~x445 & ~x449 & ~x454 & ~x466 & ~x468 & ~x474 & ~x494 & ~x495 & ~x498 & ~x502 & ~x508 & ~x511 & ~x512 & ~x532 & ~x537 & ~x554 & ~x556 & ~x558 & ~x559 & ~x565 & ~x582 & ~x584 & ~x587 & ~x588 & ~x596 & ~x607 & ~x609 & ~x615 & ~x619 & ~x623 & ~x642 & ~x672 & ~x673 & ~x691 & ~x696 & ~x700 & ~x703 & ~x721 & ~x724 & ~x726 & ~x727 & ~x736 & ~x747 & ~x749 & ~x750 & ~x752 & ~x761 & ~x764 & ~x776;
assign c14 =  x660 &  x738 & ~x194 & ~x250 & ~x556 & ~x658 & ~x676 & ~x714;
assign c16 = ~x36 & ~x80 & ~x86 & ~x160 & ~x162 & ~x188 & ~x216 & ~x231 & ~x246 & ~x261 & ~x272 & ~x274 & ~x278 & ~x287 & ~x300 & ~x304 & ~x309 & ~x316 & ~x337 & ~x358 & ~x365 & ~x454 & ~x456 & ~x458 & ~x467 & ~x469 & ~x497 & ~x504 & ~x539 & ~x558 & ~x580 & ~x582 & ~x585 & ~x608 & ~x613 & ~x618 & ~x625 & ~x651 & ~x652 & ~x655 & ~x664 & ~x673 & ~x694 & ~x706 & ~x709 & ~x764 & ~x766;
assign c18 =  x560;
assign c110 =  x718 & ~x276 & ~x658 & ~x686 & ~x742;
assign c112 =  x294 &  x319 &  x572 &  x600 &  x627 &  x682 &  x767 & ~x0 & ~x58 & ~x76 & ~x112 & ~x133 & ~x171 & ~x190 & ~x193 & ~x195 & ~x201 & ~x246 & ~x274 & ~x277 & ~x283 & ~x310 & ~x312 & ~x391 & ~x446 & ~x503 & ~x506 & ~x592 & ~x619 & ~x674 & ~x769;
assign c114 =  x320 &  x377 &  x521 &  x551 &  x572 &  x628 &  x634 &  x712 &  x739 &  x774 & ~x1 & ~x28 & ~x55 & ~x170 & ~x222 & ~x224 & ~x255 & ~x337 & ~x390 & ~x477 & ~x501 & ~x529 & ~x587 & ~x770 & ~x781;
assign c116 =  x226;
assign c118 =  x458 & ~x490 & ~x574 & ~x630 & ~x686 & ~x742;
assign c120 =  x45 &  x128 &  x408 &  x712 & ~x220 & ~x714;
assign c122 =  x20 & ~x711;
assign c124 =  x73 &  x74 &  x209 &  x238 &  x293 &  x355 &  x379 &  x407 &  x411 &  x436 &  x458 &  x515 &  x521 &  x625 &  x635 &  x710 &  x738 & ~x24 & ~x29 & ~x62 & ~x79 & ~x107 & ~x144 & ~x163 & ~x167 & ~x172 & ~x198 & ~x200 & ~x220 & ~x246 & ~x248 & ~x256 & ~x309 & ~x313 & ~x336 & ~x362 & ~x445 & ~x473 & ~x562 & ~x646 & ~x674 & ~x698 & ~x730;
assign c126 =  x407 &  x547 & ~x2 & ~x23 & ~x29 & ~x33 & ~x36 & ~x55 & ~x57 & ~x62 & ~x112 & ~x113 & ~x135 & ~x138 & ~x140 & ~x145 & ~x146 & ~x147 & ~x164 & ~x173 & ~x192 & ~x220 & ~x223 & ~x231 & ~x243 & ~x246 & ~x247 & ~x303 & ~x342 & ~x365 & ~x371 & ~x398 & ~x426 & ~x438 & ~x456 & ~x472 & ~x478 & ~x479 & ~x481 & ~x484 & ~x498 & ~x500 & ~x525 & ~x528 & ~x530 & ~x536 & ~x537 & ~x553 & ~x560 & ~x588 & ~x596 & ~x609 & ~x613 & ~x643 & ~x647 & ~x648 & ~x651 & ~x664 & ~x666 & ~x676 & ~x680 & ~x694 & ~x695 & ~x700 & ~x717 & ~x719 & ~x721 & ~x726 & ~x729 & ~x781 & ~x783;
assign c128 =  x154 &  x182 &  x211 &  x267 &  x268 &  x408 &  x520 &  x548 &  x576 &  x577 &  x656 & ~x0 & ~x6 & ~x22 & ~x25 & ~x33 & ~x34 & ~x51 & ~x57 & ~x58 & ~x60 & ~x62 & ~x77 & ~x79 & ~x85 & ~x86 & ~x88 & ~x107 & ~x108 & ~x114 & ~x116 & ~x117 & ~x137 & ~x140 & ~x142 & ~x145 & ~x146 & ~x162 & ~x169 & ~x173 & ~x190 & ~x191 & ~x194 & ~x217 & ~x218 & ~x219 & ~x220 & ~x221 & ~x223 & ~x226 & ~x228 & ~x229 & ~x230 & ~x254 & ~x275 & ~x276 & ~x278 & ~x280 & ~x281 & ~x283 & ~x301 & ~x305 & ~x307 & ~x308 & ~x311 & ~x312 & ~x363 & ~x364 & ~x369 & ~x386 & ~x389 & ~x390 & ~x391 & ~x394 & ~x397 & ~x414 & ~x418 & ~x427 & ~x441 & ~x449 & ~x454 & ~x468 & ~x469 & ~x473 & ~x476 & ~x477 & ~x481 & ~x498 & ~x500 & ~x507 & ~x509 & ~x510 & ~x511 & ~x524 & ~x526 & ~x529 & ~x531 & ~x538 & ~x562 & ~x584 & ~x585 & ~x589 & ~x593 & ~x610 & ~x612 & ~x616 & ~x618 & ~x639 & ~x644 & ~x646 & ~x669 & ~x674 & ~x692 & ~x693 & ~x694 & ~x697 & ~x698 & ~x701 & ~x723 & ~x726 & ~x728 & ~x733 & ~x735 & ~x753 & ~x759 & ~x760 & ~x764 & ~x765 & ~x770 & ~x777;
assign c130 =  x44 &  x154 &  x179 &  x186 &  x187 &  x211 &  x215 &  x237 &  x262 &  x268 &  x270 &  x325 &  x382 &  x437 &  x457 & ~x34 & ~x35 & ~x50 & ~x52 & ~x53 & ~x56 & ~x61 & ~x77 & ~x106 & ~x137 & ~x146 & ~x167 & ~x168 & ~x170 & ~x229 & ~x254 & ~x280 & ~x301 & ~x330 & ~x331 & ~x334 & ~x342 & ~x370 & ~x390 & ~x444 & ~x452 & ~x476 & ~x480 & ~x499 & ~x510 & ~x527 & ~x531 & ~x536 & ~x558 & ~x559 & ~x593 & ~x618 & ~x620 & ~x697 & ~x700 & ~x729 & ~x758 & ~x762 & ~x763;
assign c132 =  x576 & ~x3 & ~x6 & ~x20 & ~x21 & ~x26 & ~x29 & ~x32 & ~x33 & ~x48 & ~x49 & ~x64 & ~x87 & ~x104 & ~x107 & ~x113 & ~x135 & ~x136 & ~x138 & ~x142 & ~x146 & ~x165 & ~x200 & ~x201 & ~x202 & ~x216 & ~x220 & ~x221 & ~x227 & ~x249 & ~x250 & ~x259 & ~x260 & ~x289 & ~x305 & ~x307 & ~x309 & ~x312 & ~x314 & ~x315 & ~x317 & ~x327 & ~x328 & ~x336 & ~x342 & ~x361 & ~x365 & ~x367 & ~x385 & ~x394 & ~x398 & ~x399 & ~x412 & ~x421 & ~x424 & ~x449 & ~x453 & ~x467 & ~x482 & ~x485 & ~x496 & ~x500 & ~x501 & ~x507 & ~x510 & ~x512 & ~x523 & ~x531 & ~x536 & ~x539 & ~x540 & ~x551 & ~x553 & ~x559 & ~x560 & ~x563 & ~x565 & ~x569 & ~x582 & ~x586 & ~x587 & ~x593 & ~x595 & ~x608 & ~x609 & ~x611 & ~x616 & ~x617 & ~x621 & ~x623 & ~x624 & ~x637 & ~x644 & ~x647 & ~x654 & ~x668 & ~x673 & ~x675 & ~x677 & ~x678 & ~x692 & ~x696 & ~x699 & ~x704 & ~x705 & ~x706 & ~x710 & ~x730 & ~x731 & ~x735 & ~x737 & ~x753 & ~x754 & ~x756 & ~x759 & ~x780 & ~x782;
assign c134 = ~x12 & ~x63 & ~x68 & ~x80 & ~x116 & ~x142 & ~x146 & ~x190 & ~x199 & ~x243 & ~x282 & ~x302 & ~x343 & ~x344 & ~x362 & ~x370 & ~x383 & ~x413 & ~x421 & ~x427 & ~x453 & ~x466 & ~x467 & ~x468 & ~x482 & ~x494 & ~x495 & ~x508 & ~x565 & ~x567 & ~x580 & ~x594 & ~x608 & ~x644 & ~x645 & ~x674 & ~x693 & ~x726 & ~x751 & ~x757 & ~x769 & ~x776;
assign c136 =  x22;
assign c138 =  x39 &  x95 &  x295 &  x491 &  x659 &  x687 & ~x1 & ~x22 & ~x27 & ~x35 & ~x49 & ~x52 & ~x76 & ~x77 & ~x104 & ~x110 & ~x113 & ~x142 & ~x161 & ~x166 & ~x171 & ~x188 & ~x197 & ~x226 & ~x227 & ~x244 & ~x246 & ~x272 & ~x278 & ~x287 & ~x300 & ~x301 & ~x302 & ~x309 & ~x314 & ~x328 & ~x333 & ~x335 & ~x337 & ~x356 & ~x357 & ~x383 & ~x384 & ~x385 & ~x398 & ~x399 & ~x427 & ~x443 & ~x451 & ~x467 & ~x469 & ~x470 & ~x475 & ~x483 & ~x507 & ~x508 & ~x509 & ~x555 & ~x559 & ~x566 & ~x581 & ~x583 & ~x590 & ~x612 & ~x613 & ~x635 & ~x648 & ~x652 & ~x662 & ~x676 & ~x705 & ~x735 & ~x753;
assign c140 =  x265 &  x632 & ~x1 & ~x5 & ~x7 & ~x8 & ~x9 & ~x25 & ~x26 & ~x27 & ~x30 & ~x35 & ~x37 & ~x48 & ~x50 & ~x52 & ~x54 & ~x57 & ~x58 & ~x63 & ~x64 & ~x65 & ~x79 & ~x89 & ~x90 & ~x91 & ~x92 & ~x104 & ~x105 & ~x106 & ~x107 & ~x109 & ~x110 & ~x112 & ~x114 & ~x115 & ~x117 & ~x120 & ~x132 & ~x138 & ~x143 & ~x146 & ~x147 & ~x148 & ~x169 & ~x172 & ~x173 & ~x176 & ~x188 & ~x191 & ~x192 & ~x193 & ~x195 & ~x196 & ~x199 & ~x202 & ~x203 & ~x204 & ~x216 & ~x217 & ~x221 & ~x224 & ~x225 & ~x226 & ~x227 & ~x228 & ~x244 & ~x245 & ~x249 & ~x250 & ~x251 & ~x252 & ~x259 & ~x260 & ~x261 & ~x272 & ~x273 & ~x274 & ~x276 & ~x277 & ~x279 & ~x280 & ~x281 & ~x282 & ~x300 & ~x304 & ~x306 & ~x307 & ~x308 & ~x309 & ~x311 & ~x312 & ~x313 & ~x317 & ~x328 & ~x333 & ~x336 & ~x337 & ~x338 & ~x359 & ~x360 & ~x361 & ~x362 & ~x363 & ~x364 & ~x366 & ~x368 & ~x370 & ~x373 & ~x392 & ~x394 & ~x396 & ~x397 & ~x398 & ~x399 & ~x401 & ~x412 & ~x413 & ~x415 & ~x416 & ~x419 & ~x422 & ~x423 & ~x424 & ~x425 & ~x428 & ~x441 & ~x443 & ~x446 & ~x447 & ~x449 & ~x450 & ~x456 & ~x457 & ~x467 & ~x468 & ~x469 & ~x476 & ~x477 & ~x480 & ~x481 & ~x485 & ~x495 & ~x500 & ~x501 & ~x502 & ~x505 & ~x506 & ~x513 & ~x526 & ~x532 & ~x534 & ~x536 & ~x537 & ~x538 & ~x541 & ~x552 & ~x561 & ~x562 & ~x567 & ~x581 & ~x584 & ~x585 & ~x586 & ~x589 & ~x591 & ~x595 & ~x596 & ~x597 & ~x607 & ~x609 & ~x615 & ~x618 & ~x619 & ~x620 & ~x636 & ~x637 & ~x638 & ~x641 & ~x643 & ~x644 & ~x648 & ~x649 & ~x650 & ~x651 & ~x652 & ~x663 & ~x665 & ~x669 & ~x672 & ~x673 & ~x674 & ~x675 & ~x680 & ~x682 & ~x692 & ~x694 & ~x696 & ~x698 & ~x699 & ~x700 & ~x703 & ~x704 & ~x706 & ~x707 & ~x708 & ~x709 & ~x719 & ~x722 & ~x728 & ~x730 & ~x731 & ~x732 & ~x733 & ~x734 & ~x737 & ~x751 & ~x756 & ~x760 & ~x761 & ~x762 & ~x766 & ~x777 & ~x781;
assign c142 =  x255;
assign c144 = ~x36 & ~x56 & ~x186 & ~x225 & ~x230 & ~x257 & ~x259 & ~x285 & ~x306 & ~x312 & ~x314 & ~x334 & ~x371 & ~x411 & ~x412 & ~x415 & ~x480 & ~x496 & ~x595 & ~x616 & ~x620 & ~x675 & ~x695 & ~x714 & ~x728;
assign c146 =  x20;
assign c148 =  x131 & ~x116 & ~x390 & ~x490 & ~x546 & ~x630 & ~x714;
assign c150 =  x348 &  x626 &  x739 & ~x33 & ~x62 & ~x85 & ~x144 & ~x169 & ~x200 & ~x313 & ~x361 & ~x476 & ~x477 & ~x531 & ~x646 & ~x701 & ~x741;
assign c152 =  x45 &  x177 &  x298 &  x318 & ~x36 & ~x64 & ~x108 & ~x173 & ~x301 & ~x483 & ~x507 & ~x525 & ~x529 & ~x609 & ~x664 & ~x672 & ~x695 & ~x702 & ~x704 & ~x734 & ~x755;
assign c154 =  x2 & ~x156;
assign c156 =  x239 &  x240 &  x291 &  x341 &  x374 &  x509 &  x678;
assign c158 =  x672;
assign c160 =  x20 &  x343;
assign c162 = ~x0 & ~x8 & ~x20 & ~x36 & ~x47 & ~x86 & ~x116 & ~x117 & ~x132 & ~x140 & ~x141 & ~x142 & ~x159 & ~x160 & ~x162 & ~x168 & ~x172 & ~x192 & ~x201 & ~x226 & ~x230 & ~x246 & ~x257 & ~x280 & ~x300 & ~x302 & ~x309 & ~x313 & ~x336 & ~x339 & ~x340 & ~x355 & ~x361 & ~x368 & ~x387 & ~x388 & ~x391 & ~x412 & ~x413 & ~x414 & ~x421 & ~x439 & ~x446 & ~x448 & ~x466 & ~x471 & ~x473 & ~x474 & ~x500 & ~x501 & ~x502 & ~x510 & ~x522 & ~x552 & ~x559 & ~x563 & ~x583 & ~x584 & ~x612 & ~x617 & ~x621 & ~x634 & ~x635 & ~x642 & ~x648 & ~x651 & ~x667 & ~x669 & ~x672 & ~x677 & ~x678 & ~x700 & ~x701 & ~x705 & ~x717 & ~x731 & ~x736 & ~x750 & ~x752 & ~x754 & ~x774 & ~x777;
assign c164 =  x4;
assign c166 =  x684 & ~x110 & ~x137 & ~x166 & ~x193 & ~x245 & ~x280 & ~x329 & ~x367 & ~x405 & ~x433 & ~x529 & ~x565 & ~x589 & ~x592 & ~x594 & ~x641 & ~x676 & ~x679 & ~x706 & ~x707 & ~x762;
assign c168 =  x42 &  x44 &  x72 &  x98 &  x129 &  x151 &  x156 &  x179 &  x186 &  x233 &  x265 &  x269 &  x270 &  x291 &  x298 &  x344 &  x374 &  x465 &  x494 &  x739 &  x771 & ~x5 & ~x6 & ~x21 & ~x33 & ~x56 & ~x89 & ~x110 & ~x116 & ~x117 & ~x141 & ~x145 & ~x165 & ~x192 & ~x201 & ~x219 & ~x227 & ~x248 & ~x281 & ~x304 & ~x312 & ~x335 & ~x338 & ~x390 & ~x398 & ~x419 & ~x453 & ~x469 & ~x530 & ~x536 & ~x559 & ~x591 & ~x611 & ~x613 & ~x696 & ~x753 & ~x760;
assign c170 =  x514 & ~x78 & ~x517 & ~x545 & ~x714 & ~x742;
assign c172 =  x569 & ~x253 & ~x574 & ~x629 & ~x658 & ~x686;
assign c174 =  x348 &  x352 &  x378 &  x403 &  x430 &  x542 &  x684 &  x771 & ~x86 & ~x189 & ~x278 & ~x413 & ~x480 & ~x483 & ~x505 & ~x531 & ~x555 & ~x637 & ~x665 & ~x701 & ~x705 & ~x706 & ~x769 & ~x776;
assign c176 =  x19 & ~x461;
assign c178 =  x28;
assign c180 =  x0;
assign c182 =  x325 &  x351 &  x456 &  x540 &  x661 &  x689 &  x747 & ~x171 & ~x308 & ~x387 & ~x505 & ~x531 & ~x558 & ~x727 & ~x728 & ~x770;
assign c184 =  x71 &  x154 &  x183 &  x211 &  x234 &  x290 &  x487 &  x627 &  x655 & ~x1 & ~x3 & ~x5 & ~x9 & ~x23 & ~x33 & ~x36 & ~x48 & ~x60 & ~x62 & ~x77 & ~x85 & ~x89 & ~x105 & ~x106 & ~x111 & ~x134 & ~x144 & ~x145 & ~x162 & ~x169 & ~x174 & ~x191 & ~x202 & ~x228 & ~x230 & ~x231 & ~x248 & ~x250 & ~x274 & ~x275 & ~x281 & ~x344 & ~x358 & ~x363 & ~x369 & ~x386 & ~x389 & ~x397 & ~x400 & ~x416 & ~x443 & ~x445 & ~x447 & ~x454 & ~x468 & ~x474 & ~x500 & ~x534 & ~x536 & ~x556 & ~x567 & ~x581 & ~x583 & ~x585 & ~x609 & ~x610 & ~x616 & ~x635 & ~x643 & ~x648 & ~x665 & ~x666 & ~x671 & ~x672 & ~x678 & ~x724 & ~x725 & ~x731 & ~x748 & ~x757 & ~x760;
assign c186 =  x572 & ~x456 & ~x597 & ~x603 & ~x710;
assign c188 = ~x323 & ~x489 & ~x517 & ~x545 & ~x546 & ~x603 & ~x630 & ~x659 & ~x714 & ~x715 & ~x742;
assign c190 =  x739 & ~x29 & ~x49 & ~x52 & ~x146 & ~x199 & ~x259 & ~x283 & ~x284 & ~x315 & ~x329 & ~x366 & ~x392 & ~x417 & ~x423 & ~x426 & ~x469 & ~x473 & ~x498 & ~x530 & ~x561 & ~x585 & ~x595 & ~x615 & ~x673 & ~x674 & ~x742 & ~x755;
assign c192 =  x239 &  x269 &  x408 & ~x0 & ~x20 & ~x21 & ~x56 & ~x57 & ~x58 & ~x105 & ~x106 & ~x133 & ~x169 & ~x172 & ~x191 & ~x216 & ~x224 & ~x257 & ~x274 & ~x303 & ~x305 & ~x306 & ~x308 & ~x309 & ~x316 & ~x356 & ~x384 & ~x415 & ~x420 & ~x421 & ~x422 & ~x427 & ~x440 & ~x473 & ~x476 & ~x485 & ~x496 & ~x506 & ~x540 & ~x552 & ~x554 & ~x558 & ~x564 & ~x567 & ~x593 & ~x596 & ~x608 & ~x624 & ~x645 & ~x665 & ~x670 & ~x673 & ~x677 & ~x694 & ~x696 & ~x701 & ~x707 & ~x728 & ~x731 & ~x734 & ~x751 & ~x754 & ~x780;
assign c194 =  x14 & ~x357 & ~x436;
assign c196 =  x409 &  x605 & ~x54 & ~x56 & ~x66 & ~x147 & ~x250 & ~x332 & ~x442 & ~x480 & ~x508 & ~x526 & ~x615 & ~x640 & ~x733 & ~x751 & ~x757;
assign c198 =  x594 & ~x629 & ~x740;
assign c1100 =  x342 &  x763 & ~x768;
assign c1102 =  x68 &  x96 &  x265 &  x267 &  x268 &  x297 &  x323 &  x346 &  x376 &  x548 &  x576 & ~x1 & ~x5 & ~x23 & ~x24 & ~x26 & ~x32 & ~x52 & ~x54 & ~x62 & ~x86 & ~x89 & ~x105 & ~x116 & ~x117 & ~x146 & ~x188 & ~x193 & ~x223 & ~x279 & ~x284 & ~x312 & ~x333 & ~x334 & ~x369 & ~x442 & ~x453 & ~x455 & ~x467 & ~x469 & ~x478 & ~x480 & ~x495 & ~x504 & ~x510 & ~x511 & ~x528 & ~x531 & ~x579 & ~x583 & ~x590 & ~x596 & ~x609 & ~x621 & ~x635 & ~x636 & ~x641 & ~x643 & ~x664 & ~x669 & ~x670 & ~x680 & ~x693 & ~x695 & ~x696 & ~x699 & ~x706 & ~x708 & ~x725 & ~x728 & ~x729 & ~x732 & ~x747 & ~x758 & ~x759 & ~x775;
assign c1104 =  x718 & ~x68 & ~x244 & ~x316 & ~x328;
assign c1106 =  x616;
assign c1108 =  x13 &  x15 &  x16 &  x17 &  x130 &  x326 &  x464 & ~x78 & ~x109 & ~x114 & ~x134 & ~x190 & ~x224 & ~x302 & ~x306 & ~x332 & ~x385 & ~x470 & ~x481 & ~x482 & ~x637 & ~x702 & ~x730;
assign c1110 =  x616;
assign c1112 =  x14 &  x45 &  x66 &  x214 & ~x2 & ~x21 & ~x22 & ~x30 & ~x33 & ~x78 & ~x84 & ~x85 & ~x88 & ~x91 & ~x133 & ~x137 & ~x144 & ~x145 & ~x163 & ~x170 & ~x173 & ~x175 & ~x189 & ~x191 & ~x192 & ~x198 & ~x203 & ~x218 & ~x220 & ~x221 & ~x224 & ~x225 & ~x230 & ~x246 & ~x251 & ~x252 & ~x257 & ~x259 & ~x274 & ~x276 & ~x278 & ~x285 & ~x286 & ~x287 & ~x303 & ~x312 & ~x313 & ~x314 & ~x329 & ~x338 & ~x340 & ~x341 & ~x343 & ~x359 & ~x361 & ~x367 & ~x385 & ~x386 & ~x387 & ~x391 & ~x392 & ~x395 & ~x396 & ~x416 & ~x422 & ~x424 & ~x425 & ~x427 & ~x441 & ~x442 & ~x446 & ~x472 & ~x474 & ~x475 & ~x500 & ~x502 & ~x507 & ~x508 & ~x530 & ~x532 & ~x533 & ~x538 & ~x539 & ~x553 & ~x558 & ~x564 & ~x567 & ~x581 & ~x585 & ~x587 & ~x588 & ~x593 & ~x609 & ~x611 & ~x613 & ~x617 & ~x618 & ~x619 & ~x649 & ~x650 & ~x666 & ~x671 & ~x694 & ~x695 & ~x702 & ~x704 & ~x721 & ~x731 & ~x735 & ~x749 & ~x754 & ~x755 & ~x781;
assign c1114 =  x13 &  x17 &  x18 & ~x6 & ~x53 & ~x60 & ~x136 & ~x305 & ~x528 & ~x648 & ~x667 & ~x720 & ~x722 & ~x749 & ~x750 & ~x777;
assign c1116 =  x11 &  x185 &  x325 &  x353 & ~x49 & ~x58 & ~x63 & ~x109 & ~x120 & ~x147 & ~x176 & ~x218 & ~x223 & ~x253 & ~x282 & ~x312 & ~x334 & ~x414 & ~x449 & ~x594 & ~x647 & ~x677 & ~x757 & ~x759;
assign c1118 =  x73 &  x154 &  x213 &  x242 &  x262 &  x269 &  x318 &  x354 &  x741 & ~x21 & ~x35 & ~x80 & ~x86 & ~x114 & ~x116 & ~x136 & ~x146 & ~x190 & ~x201 & ~x254 & ~x285 & ~x333 & ~x361 & ~x365 & ~x370 & ~x397 & ~x417 & ~x426 & ~x444 & ~x469 & ~x482 & ~x483 & ~x525 & ~x567 & ~x588 & ~x613 & ~x642 & ~x643 & ~x645 & ~x665 & ~x668 & ~x672 & ~x694 & ~x706 & ~x727 & ~x753 & ~x755 & ~x756 & ~x757 & ~x763 & ~x777;
assign c1120 =  x127 &  x154 &  x183 &  x240 &  x320 &  x324 &  x435 &  x491 &  x519 & ~x104 & ~x120 & ~x142 & ~x169 & ~x194 & ~x216 & ~x228 & ~x275 & ~x287 & ~x300 & ~x327 & ~x344 & ~x355 & ~x360 & ~x369 & ~x401 & ~x427 & ~x428 & ~x429 & ~x444 & ~x457 & ~x468 & ~x505 & ~x526 & ~x624 & ~x648 & ~x651 & ~x653 & ~x662 & ~x668 & ~x680 & ~x700 & ~x707 & ~x709 & ~x735 & ~x737 & ~x749 & ~x751 & ~x755;
assign c1122 =  x10 &  x13 &  x38 & ~x3 & ~x56 & ~x76 & ~x78 & ~x112 & ~x115 & ~x118 & ~x139 & ~x142 & ~x145 & ~x170 & ~x172 & ~x175 & ~x194 & ~x203 & ~x217 & ~x223 & ~x230 & ~x250 & ~x273 & ~x274 & ~x286 & ~x302 & ~x307 & ~x314 & ~x329 & ~x338 & ~x359 & ~x362 & ~x384 & ~x389 & ~x412 & ~x426 & ~x452 & ~x454 & ~x468 & ~x478 & ~x500 & ~x504 & ~x529 & ~x557 & ~x559 & ~x581 & ~x586 & ~x591 & ~x594 & ~x672 & ~x679 & ~x693 & ~x700 & ~x706 & ~x707 & ~x721 & ~x752 & ~x759 & ~x778;
assign c1124 =  x656 & ~x2 & ~x29 & ~x52 & ~x63 & ~x78 & ~x89 & ~x141 & ~x161 & ~x162 & ~x171 & ~x189 & ~x196 & ~x198 & ~x201 & ~x217 & ~x218 & ~x227 & ~x231 & ~x246 & ~x250 & ~x273 & ~x286 & ~x308 & ~x309 & ~x313 & ~x331 & ~x334 & ~x341 & ~x342 & ~x357 & ~x358 & ~x370 & ~x415 & ~x419 & ~x422 & ~x444 & ~x446 & ~x448 & ~x472 & ~x475 & ~x478 & ~x480 & ~x498 & ~x501 & ~x536 & ~x537 & ~x556 & ~x557 & ~x563 & ~x585 & ~x587 & ~x613 & ~x616 & ~x618 & ~x620 & ~x639 & ~x643 & ~x648 & ~x658 & ~x667 & ~x672 & ~x686 & ~x702 & ~x726 & ~x762 & ~x770 & ~x781;
assign c1126 =  x234 &  x236 &  x238 &  x268 &  x296 &  x373 &  x432 &  x598 &  x605 &  x626 &  x656 &  x709 &  x737 &  x745 & ~x23 & ~x24 & ~x50 & ~x85 & ~x89 & ~x110 & ~x111 & ~x251 & ~x281 & ~x304 & ~x389 & ~x391 & ~x419 & ~x503 & ~x504 & ~x505 & ~x614 & ~x645 & ~x701 & ~x769;
assign c1128 =  x576 &  x684 & ~x0 & ~x1 & ~x2 & ~x3 & ~x4 & ~x6 & ~x7 & ~x9 & ~x19 & ~x20 & ~x21 & ~x22 & ~x23 & ~x26 & ~x27 & ~x28 & ~x29 & ~x34 & ~x35 & ~x36 & ~x48 & ~x49 & ~x50 & ~x51 & ~x52 & ~x53 & ~x56 & ~x57 & ~x58 & ~x60 & ~x62 & ~x63 & ~x76 & ~x77 & ~x78 & ~x79 & ~x80 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x90 & ~x92 & ~x105 & ~x106 & ~x108 & ~x109 & ~x110 & ~x112 & ~x113 & ~x114 & ~x115 & ~x117 & ~x118 & ~x119 & ~x120 & ~x132 & ~x133 & ~x134 & ~x137 & ~x138 & ~x143 & ~x144 & ~x145 & ~x147 & ~x148 & ~x160 & ~x161 & ~x163 & ~x165 & ~x168 & ~x169 & ~x170 & ~x171 & ~x172 & ~x174 & ~x176 & ~x189 & ~x190 & ~x192 & ~x193 & ~x194 & ~x199 & ~x200 & ~x203 & ~x216 & ~x217 & ~x219 & ~x220 & ~x221 & ~x222 & ~x223 & ~x224 & ~x226 & ~x230 & ~x244 & ~x246 & ~x247 & ~x248 & ~x249 & ~x250 & ~x252 & ~x254 & ~x255 & ~x256 & ~x258 & ~x259 & ~x260 & ~x272 & ~x276 & ~x279 & ~x281 & ~x283 & ~x284 & ~x285 & ~x286 & ~x287 & ~x300 & ~x301 & ~x303 & ~x304 & ~x306 & ~x307 & ~x308 & ~x309 & ~x310 & ~x313 & ~x315 & ~x329 & ~x330 & ~x331 & ~x332 & ~x333 & ~x335 & ~x336 & ~x337 & ~x339 & ~x341 & ~x344 & ~x356 & ~x358 & ~x359 & ~x360 & ~x361 & ~x363 & ~x365 & ~x366 & ~x367 & ~x370 & ~x371 & ~x384 & ~x385 & ~x386 & ~x387 & ~x388 & ~x389 & ~x390 & ~x391 & ~x393 & ~x395 & ~x396 & ~x397 & ~x398 & ~x400 & ~x411 & ~x412 & ~x413 & ~x414 & ~x415 & ~x416 & ~x418 & ~x419 & ~x420 & ~x423 & ~x425 & ~x426 & ~x427 & ~x439 & ~x440 & ~x441 & ~x443 & ~x444 & ~x445 & ~x446 & ~x448 & ~x450 & ~x451 & ~x453 & ~x454 & ~x456 & ~x468 & ~x470 & ~x472 & ~x473 & ~x475 & ~x477 & ~x478 & ~x479 & ~x482 & ~x484 & ~x496 & ~x498 & ~x499 & ~x500 & ~x501 & ~x503 & ~x504 & ~x506 & ~x507 & ~x508 & ~x509 & ~x511 & ~x525 & ~x526 & ~x527 & ~x528 & ~x529 & ~x530 & ~x536 & ~x537 & ~x538 & ~x552 & ~x553 & ~x554 & ~x555 & ~x556 & ~x557 & ~x559 & ~x560 & ~x563 & ~x564 & ~x567 & ~x568 & ~x580 & ~x581 & ~x582 & ~x583 & ~x584 & ~x585 & ~x587 & ~x588 & ~x589 & ~x593 & ~x594 & ~x595 & ~x596 & ~x608 & ~x610 & ~x613 & ~x615 & ~x616 & ~x617 & ~x619 & ~x620 & ~x621 & ~x623 & ~x624 & ~x625 & ~x636 & ~x638 & ~x640 & ~x642 & ~x643 & ~x645 & ~x646 & ~x648 & ~x650 & ~x651 & ~x652 & ~x664 & ~x665 & ~x666 & ~x667 & ~x669 & ~x670 & ~x671 & ~x674 & ~x675 & ~x676 & ~x677 & ~x678 & ~x679 & ~x692 & ~x693 & ~x694 & ~x695 & ~x696 & ~x697 & ~x705 & ~x706 & ~x719 & ~x721 & ~x722 & ~x724 & ~x726 & ~x728 & ~x729 & ~x730 & ~x731 & ~x734 & ~x735 & ~x736 & ~x748 & ~x749 & ~x750 & ~x752 & ~x753 & ~x756 & ~x757 & ~x759 & ~x761 & ~x762 & ~x764 & ~x765 & ~x770 & ~x777 & ~x778 & ~x779 & ~x780 & ~x781;
assign c1130 =  x127 &  x238 &  x323 &  x379 &  x407 &  x435 &  x463 &  x547 &  x603 &  x687 &  x715 & ~x59 & ~x77 & ~x88 & ~x111 & ~x196 & ~x226 & ~x253 & ~x254 & ~x283 & ~x340 & ~x358 & ~x453 & ~x477 & ~x498 & ~x503 & ~x504 & ~x506 & ~x509 & ~x615 & ~x648 & ~x649 & ~x668 & ~x672 & ~x673 & ~x675 & ~x678 & ~x689 & ~x704 & ~x745;
assign c1132 =  x632 &  x716 & ~x35 & ~x43 & ~x52 & ~x56 & ~x91 & ~x105 & ~x109 & ~x134 & ~x144 & ~x148 & ~x200 & ~x202 & ~x203 & ~x220 & ~x224 & ~x227 & ~x230 & ~x231 & ~x253 & ~x258 & ~x260 & ~x273 & ~x274 & ~x282 & ~x284 & ~x303 & ~x313 & ~x315 & ~x336 & ~x360 & ~x361 & ~x392 & ~x396 & ~x422 & ~x424 & ~x425 & ~x441 & ~x449 & ~x455 & ~x473 & ~x482 & ~x499 & ~x502 & ~x553 & ~x555 & ~x556 & ~x562 & ~x564 & ~x585 & ~x586 & ~x594 & ~x610 & ~x618 & ~x620 & ~x643 & ~x647 & ~x650 & ~x668 & ~x696 & ~x699 & ~x706 & ~x754 & ~x755 & ~x760 & ~x770 & ~x783;
assign c1134 =  x39 &  x290 &  x323 &  x325 & ~x5 & ~x86 & ~x147 & ~x161 & ~x164 & ~x165 & ~x204 & ~x220 & ~x224 & ~x313 & ~x316 & ~x344 & ~x385 & ~x387 & ~x497 & ~x498 & ~x525 & ~x562 & ~x563 & ~x635 & ~x733 & ~x754;
assign c1136 = ~x12 & ~x31 & ~x46 & ~x55 & ~x56 & ~x104 & ~x110 & ~x113 & ~x173 & ~x188 & ~x205 & ~x228 & ~x301 & ~x307 & ~x315 & ~x330 & ~x342 & ~x386 & ~x391 & ~x410 & ~x413 & ~x418 & ~x429 & ~x439 & ~x446 & ~x479 & ~x484 & ~x496 & ~x497 & ~x523 & ~x531 & ~x541 & ~x562 & ~x563 & ~x569 & ~x583 & ~x595 & ~x621 & ~x634 & ~x636 & ~x662 & ~x671 & ~x699 & ~x700 & ~x720 & ~x727 & ~x729 & ~x761 & ~x769 & ~x774;
assign c1138 =  x101 &  x128 &  x237 &  x349 &  x408 &  x431 &  x439 &  x521 &  x568 &  x624 &  x718 &  x736 &  x738 & ~x81 & ~x111 & ~x145 & ~x507 & ~x557 & ~x566 & ~x696 & ~x701;
assign c1140 =  x152 &  x210 &  x236 &  x242 &  x266 &  x269 &  x288 &  x291 &  x293 &  x294 &  x296 &  x371 &  x375 &  x382 &  x437 &  x484 &  x493 &  x523 &  x539 &  x567 &  x568 &  x569 &  x579 &  x596 &  x607 &  x624 &  x652 &  x679 &  x709 & ~x32 & ~x52 & ~x59 & ~x84 & ~x195 & ~x252 & ~x278 & ~x781;
assign c1142 =  x782;
assign c1146 =  x45 &  x126 &  x241 &  x290 & ~x259 & ~x273 & ~x281 & ~x365 & ~x444 & ~x468 & ~x585 & ~x708;
assign c1148 = ~x26 & ~x31 & ~x48 & ~x51 & ~x54 & ~x55 & ~x58 & ~x62 & ~x63 & ~x80 & ~x86 & ~x87 & ~x90 & ~x104 & ~x106 & ~x111 & ~x117 & ~x192 & ~x194 & ~x197 & ~x200 & ~x202 & ~x219 & ~x220 & ~x226 & ~x228 & ~x252 & ~x256 & ~x258 & ~x260 & ~x279 & ~x306 & ~x312 & ~x329 & ~x337 & ~x338 & ~x342 & ~x364 & ~x366 & ~x385 & ~x389 & ~x414 & ~x417 & ~x420 & ~x423 & ~x424 & ~x447 & ~x449 & ~x450 & ~x452 & ~x468 & ~x472 & ~x482 & ~x483 & ~x490 & ~x498 & ~x504 & ~x507 & ~x508 & ~x509 & ~x511 & ~x526 & ~x528 & ~x529 & ~x530 & ~x538 & ~x557 & ~x560 & ~x562 & ~x564 & ~x568 & ~x611 & ~x615 & ~x640 & ~x642 & ~x646 & ~x665 & ~x668 & ~x673 & ~x696 & ~x705 & ~x706 & ~x723 & ~x729 & ~x736 & ~x751 & ~x753 & ~x754 & ~x759 & ~x778 & ~x779;
assign c1150 =  x267 &  x379 & ~x3 & ~x27 & ~x28 & ~x33 & ~x59 & ~x75 & ~x84 & ~x86 & ~x104 & ~x111 & ~x132 & ~x134 & ~x135 & ~x173 & ~x174 & ~x188 & ~x189 & ~x190 & ~x199 & ~x201 & ~x225 & ~x259 & ~x279 & ~x303 & ~x306 & ~x317 & ~x327 & ~x333 & ~x341 & ~x344 & ~x367 & ~x373 & ~x396 & ~x417 & ~x426 & ~x442 & ~x446 & ~x454 & ~x455 & ~x467 & ~x473 & ~x476 & ~x495 & ~x508 & ~x512 & ~x523 & ~x524 & ~x529 & ~x560 & ~x611 & ~x622 & ~x625 & ~x644 & ~x649 & ~x675 & ~x678 & ~x725 & ~x727 & ~x728 & ~x729 & ~x732 & ~x738 & ~x755 & ~x758 & ~x760 & ~x764;
assign c1152 =  x605 & ~x224 & ~x278 & ~x336 & ~x602 & ~x630 & ~x658 & ~x686 & ~x714 & ~x759 & ~x770;
assign c1154 =  x100 &  x240 &  x269 &  x297 &  x325 &  x375 &  x432 &  x629 &  x713 & ~x61 & ~x245 & ~x285 & ~x306 & ~x419 & ~x425 & ~x468 & ~x482 & ~x540 & ~x555 & ~x642 & ~x650 & ~x663 & ~x706 & ~x719 & ~x732 & ~x733 & ~x765;
assign c1156 =  x43 &  x69 &  x233 &  x242 &  x317 &  x326 &  x382 & ~x63 & ~x64 & ~x245 & ~x427 & ~x503 & ~x507 & ~x587 & ~x589 & ~x650 & ~x733;
assign c1158 =  x70 &  x72 &  x98 &  x151 &  x153 &  x178 &  x213 &  x236 &  x269 &  x293 &  x408 &  x741 & ~x61 & ~x62 & ~x63 & ~x82 & ~x112 & ~x118 & ~x144 & ~x161 & ~x168 & ~x189 & ~x202 & ~x223 & ~x225 & ~x248 & ~x277 & ~x304 & ~x336 & ~x337 & ~x366 & ~x384 & ~x387 & ~x388 & ~x390 & ~x416 & ~x419 & ~x427 & ~x440 & ~x451 & ~x471 & ~x480 & ~x483 & ~x498 & ~x503 & ~x510 & ~x524 & ~x535 & ~x552 & ~x560 & ~x619 & ~x620 & ~x639 & ~x641 & ~x669 & ~x675 & ~x676 & ~x679 & ~x691 & ~x693 & ~x695 & ~x705 & ~x708 & ~x722 & ~x734 & ~x749 & ~x759 & ~x777 & ~x781 & ~x783;
assign c1160 =  x211 &  x716 & ~x19 & ~x29 & ~x32 & ~x35 & ~x57 & ~x61 & ~x62 & ~x63 & ~x80 & ~x83 & ~x89 & ~x104 & ~x105 & ~x108 & ~x119 & ~x132 & ~x134 & ~x139 & ~x141 & ~x142 & ~x143 & ~x175 & ~x189 & ~x193 & ~x194 & ~x196 & ~x217 & ~x228 & ~x231 & ~x248 & ~x254 & ~x257 & ~x273 & ~x279 & ~x283 & ~x286 & ~x302 & ~x330 & ~x332 & ~x336 & ~x338 & ~x341 & ~x342 & ~x359 & ~x390 & ~x414 & ~x425 & ~x426 & ~x428 & ~x452 & ~x456 & ~x479 & ~x480 & ~x481 & ~x483 & ~x499 & ~x503 & ~x505 & ~x509 & ~x538 & ~x540 & ~x553 & ~x554 & ~x558 & ~x582 & ~x583 & ~x591 & ~x592 & ~x594 & ~x596 & ~x609 & ~x619 & ~x623 & ~x647 & ~x652 & ~x670 & ~x671 & ~x705 & ~x720 & ~x723 & ~x725 & ~x733 & ~x734 & ~x735 & ~x736 & ~x754 & ~x762 & ~x763 & ~x764 & ~x765 & ~x770;
assign c1162 =  x14 &  x41 &  x604 & ~x0 & ~x1 & ~x2 & ~x3 & ~x6 & ~x21 & ~x22 & ~x23 & ~x30 & ~x31 & ~x33 & ~x34 & ~x51 & ~x52 & ~x53 & ~x54 & ~x58 & ~x59 & ~x60 & ~x62 & ~x63 & ~x77 & ~x80 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x86 & ~x87 & ~x89 & ~x105 & ~x106 & ~x108 & ~x109 & ~x115 & ~x118 & ~x119 & ~x132 & ~x135 & ~x137 & ~x139 & ~x141 & ~x142 & ~x143 & ~x144 & ~x145 & ~x146 & ~x160 & ~x162 & ~x163 & ~x164 & ~x165 & ~x166 & ~x169 & ~x170 & ~x172 & ~x175 & ~x188 & ~x190 & ~x191 & ~x198 & ~x199 & ~x200 & ~x201 & ~x203 & ~x217 & ~x218 & ~x219 & ~x221 & ~x222 & ~x223 & ~x228 & ~x245 & ~x246 & ~x247 & ~x249 & ~x251 & ~x256 & ~x257 & ~x258 & ~x272 & ~x273 & ~x274 & ~x275 & ~x276 & ~x278 & ~x279 & ~x281 & ~x282 & ~x283 & ~x284 & ~x285 & ~x286 & ~x287 & ~x288 & ~x300 & ~x301 & ~x304 & ~x305 & ~x306 & ~x307 & ~x308 & ~x309 & ~x311 & ~x312 & ~x315 & ~x328 & ~x329 & ~x330 & ~x331 & ~x332 & ~x333 & ~x336 & ~x337 & ~x338 & ~x340 & ~x342 & ~x343 & ~x356 & ~x357 & ~x358 & ~x360 & ~x363 & ~x365 & ~x366 & ~x369 & ~x370 & ~x383 & ~x385 & ~x388 & ~x389 & ~x390 & ~x391 & ~x392 & ~x395 & ~x396 & ~x397 & ~x398 & ~x411 & ~x412 & ~x414 & ~x415 & ~x416 & ~x417 & ~x418 & ~x419 & ~x420 & ~x421 & ~x422 & ~x423 & ~x424 & ~x425 & ~x426 & ~x427 & ~x439 & ~x441 & ~x442 & ~x444 & ~x445 & ~x446 & ~x447 & ~x448 & ~x450 & ~x451 & ~x453 & ~x454 & ~x456 & ~x467 & ~x469 & ~x470 & ~x471 & ~x472 & ~x473 & ~x474 & ~x477 & ~x480 & ~x481 & ~x496 & ~x498 & ~x499 & ~x501 & ~x503 & ~x505 & ~x506 & ~x507 & ~x524 & ~x525 & ~x527 & ~x528 & ~x532 & ~x533 & ~x534 & ~x535 & ~x536 & ~x537 & ~x538 & ~x552 & ~x554 & ~x555 & ~x557 & ~x558 & ~x559 & ~x561 & ~x562 & ~x565 & ~x567 & ~x580 & ~x581 & ~x582 & ~x583 & ~x584 & ~x585 & ~x586 & ~x589 & ~x590 & ~x591 & ~x593 & ~x595 & ~x608 & ~x609 & ~x610 & ~x611 & ~x612 & ~x613 & ~x617 & ~x620 & ~x621 & ~x622 & ~x636 & ~x637 & ~x638 & ~x639 & ~x641 & ~x642 & ~x643 & ~x648 & ~x651 & ~x664 & ~x665 & ~x666 & ~x667 & ~x668 & ~x670 & ~x672 & ~x673 & ~x674 & ~x676 & ~x677 & ~x678 & ~x679 & ~x680 & ~x692 & ~x693 & ~x694 & ~x695 & ~x697 & ~x700 & ~x703 & ~x705 & ~x706 & ~x707 & ~x720 & ~x721 & ~x722 & ~x723 & ~x724 & ~x725 & ~x726 & ~x728 & ~x729 & ~x731 & ~x732 & ~x733 & ~x751 & ~x754 & ~x756 & ~x758 & ~x759 & ~x762 & ~x776;
assign c1164 =  x57;
assign c1166 =  x544 & ~x13 & ~x41 & ~x146 & ~x162 & ~x285 & ~x416 & ~x565 & ~x611 & ~x667 & ~x694 & ~x770;
assign c1168 =  x516 &  x657 & ~x91 & ~x166 & ~x215 & ~x253 & ~x307 & ~x503 & ~x615 & ~x626 & ~x704 & ~x757 & ~x779;
assign c1170 =  x407 &  x435 &  x488 &  x628 &  x684 & ~x0 & ~x15 & ~x32 & ~x33 & ~x56 & ~x63 & ~x79 & ~x107 & ~x115 & ~x137 & ~x145 & ~x219 & ~x221 & ~x247 & ~x255 & ~x274 & ~x276 & ~x280 & ~x307 & ~x330 & ~x332 & ~x366 & ~x386 & ~x389 & ~x418 & ~x422 & ~x424 & ~x475 & ~x478 & ~x481 & ~x504 & ~x507 & ~x531 & ~x610 & ~x620 & ~x640 & ~x648 & ~x649 & ~x666 & ~x669 & ~x686 & ~x703 & ~x704 & ~x723 & ~x778;
assign c1172 =  x265 &  x410 &  x540 &  x605 &  x624 &  x632 &  x652 & ~x192 & ~x277 & ~x444 & ~x725 & ~x769;
assign c1174 =  x45 &  x122 &  x373 &  x384 &  x410 &  x439 &  x494 &  x596 &  x607 &  x624 & ~x24 & ~x30 & ~x80 & ~x82 & ~x113 & ~x171 & ~x221 & ~x250 & ~x362 & ~x420 & ~x585 & ~x590 & ~x700 & ~x758 & ~x781;
assign c1176 =  x50;
assign c1178 =  x10 &  x38 &  x661 & ~x36 & ~x106 & ~x148 & ~x200 & ~x256 & ~x260 & ~x342 & ~x496 & ~x564 & ~x679 & ~x754;
assign c1180 =  x128 &  x210 &  x459 & ~x25 & ~x26 & ~x336 & ~x546 & ~x574 & ~x602 & ~x614;
assign c1182 =  x376 &  x405 & ~x3 & ~x6 & ~x21 & ~x22 & ~x33 & ~x48 & ~x60 & ~x79 & ~x88 & ~x89 & ~x92 & ~x106 & ~x107 & ~x108 & ~x171 & ~x173 & ~x174 & ~x194 & ~x203 & ~x223 & ~x228 & ~x246 & ~x247 & ~x259 & ~x272 & ~x276 & ~x277 & ~x281 & ~x341 & ~x355 & ~x361 & ~x367 & ~x385 & ~x390 & ~x391 & ~x398 & ~x401 & ~x443 & ~x446 & ~x452 & ~x456 & ~x457 & ~x467 & ~x478 & ~x480 & ~x500 & ~x511 & ~x513 & ~x523 & ~x524 & ~x534 & ~x558 & ~x613 & ~x624 & ~x637 & ~x640 & ~x647 & ~x650 & ~x681 & ~x693 & ~x695 & ~x697 & ~x698 & ~x705 & ~x709 & ~x722 & ~x733 & ~x753 & ~x756 & ~x758 & ~x761 & ~x770;
assign c1184 =  x22 & ~x627;
assign c1186 =  x82;
assign c1188 =  x105 &  x314 &  x399 &  x651;
assign c1190 =  x717 & ~x27 & ~x76 & ~x77 & ~x161 & ~x225 & ~x390 & ~x393 & ~x415 & ~x527 & ~x609 & ~x637 & ~x643 & ~x658 & ~x665 & ~x686 & ~x714;
assign c1192 =  x151 &  x179 &  x210 & ~x199 & ~x518 & ~x546;
assign c1194 =  x339;
assign c1196 =  x47 &  x103 &  x154 &  x176 &  x179 &  x209 &  x232 &  x267 &  x271 &  x289 &  x577 &  x681 &  x709;
assign c1198 =  x151 &  x154 &  x182 &  x207 &  x212 &  x239 &  x324 &  x347 &  x348 &  x432 & ~x1 & ~x21 & ~x31 & ~x37 & ~x51 & ~x59 & ~x65 & ~x82 & ~x89 & ~x115 & ~x116 & ~x132 & ~x134 & ~x140 & ~x146 & ~x148 & ~x162 & ~x175 & ~x188 & ~x191 & ~x193 & ~x194 & ~x196 & ~x201 & ~x216 & ~x223 & ~x229 & ~x231 & ~x244 & ~x245 & ~x254 & ~x257 & ~x259 & ~x272 & ~x273 & ~x274 & ~x279 & ~x284 & ~x307 & ~x310 & ~x313 & ~x327 & ~x328 & ~x331 & ~x335 & ~x338 & ~x360 & ~x383 & ~x384 & ~x385 & ~x394 & ~x399 & ~x400 & ~x412 & ~x427 & ~x428 & ~x451 & ~x467 & ~x472 & ~x477 & ~x484 & ~x502 & ~x524 & ~x529 & ~x534 & ~x551 & ~x552 & ~x554 & ~x555 & ~x557 & ~x568 & ~x585 & ~x607 & ~x612 & ~x619 & ~x624 & ~x635 & ~x642 & ~x644 & ~x652 & ~x678 & ~x680 & ~x703 & ~x705 & ~x708 & ~x724 & ~x734 & ~x736 & ~x748 & ~x759 & ~x761 & ~x762 & ~x776 & ~x777 & ~x780 & ~x781;
assign c1200 =  x97 &  x203 &  x231 &  x343 &  x596 & ~x767;
assign c1202 =  x263 &  x348 &  x573 & ~x24 & ~x36 & ~x52 & ~x82 & ~x87 & ~x88 & ~x90 & ~x92 & ~x106 & ~x109 & ~x135 & ~x142 & ~x163 & ~x165 & ~x166 & ~x192 & ~x197 & ~x198 & ~x255 & ~x272 & ~x285 & ~x288 & ~x289 & ~x302 & ~x303 & ~x311 & ~x328 & ~x336 & ~x338 & ~x345 & ~x359 & ~x362 & ~x373 & ~x398 & ~x400 & ~x401 & ~x416 & ~x419 & ~x422 & ~x447 & ~x485 & ~x525 & ~x527 & ~x540 & ~x554 & ~x611 & ~x622 & ~x625 & ~x637 & ~x638 & ~x652 & ~x654 & ~x665 & ~x666 & ~x678 & ~x681 & ~x682 & ~x695 & ~x698 & ~x701 & ~x702 & ~x705 & ~x706 & ~x707 & ~x708 & ~x710 & ~x719 & ~x720 & ~x722 & ~x779;
assign c1204 =  x73 &  x154 &  x235 &  x237 &  x268 &  x298 &  x344 &  x349 &  x375 &  x407 &  x429 &  x437 &  x579 &  x595 &  x596 &  x653 &  x707 &  x735 &  x736 & ~x23 & ~x25 & ~x30 & ~x54 & ~x55 & ~x108 & ~x109 & ~x114 & ~x141 & ~x220 & ~x221 & ~x251 & ~x277 & ~x279 & ~x307 & ~x395 & ~x422 & ~x447 & ~x559 & ~x561 & ~x589 & ~x613 & ~x642 & ~x644 & ~x670 & ~x698 & ~x726;
assign c1206 =  x179 &  x181 &  x182 &  x269 &  x297 &  x318 &  x575 &  x576 &  x603 &  x604 &  x628 &  x631 &  x685 & ~x0 & ~x30 & ~x52 & ~x61 & ~x79 & ~x83 & ~x142 & ~x167 & ~x171 & ~x225 & ~x274 & ~x276 & ~x302 & ~x329 & ~x370 & ~x388 & ~x389 & ~x416 & ~x423 & ~x426 & ~x453 & ~x478 & ~x525 & ~x553 & ~x566 & ~x586 & ~x619 & ~x623 & ~x650 & ~x674 & ~x693 & ~x750 & ~x752 & ~x759 & ~x770 & ~x778;
assign c1208 =  x521 & ~x80 & ~x81 & ~x142 & ~x224 & ~x308 & ~x331 & ~x337 & ~x394 & ~x476 & ~x506 & ~x574 & ~x589 & ~x602 & ~x630 & ~x644 & ~x658 & ~x686 & ~x714 & ~x770;
assign c1210 =  x435 &  x463 &  x491 &  x682 &  x771 & ~x23 & ~x26 & ~x31 & ~x51 & ~x60 & ~x77 & ~x80 & ~x86 & ~x91 & ~x104 & ~x107 & ~x112 & ~x119 & ~x132 & ~x137 & ~x146 & ~x148 & ~x161 & ~x162 & ~x168 & ~x170 & ~x171 & ~x174 & ~x187 & ~x188 & ~x189 & ~x192 & ~x198 & ~x229 & ~x271 & ~x273 & ~x276 & ~x279 & ~x280 & ~x283 & ~x309 & ~x313 & ~x327 & ~x329 & ~x331 & ~x356 & ~x357 & ~x360 & ~x361 & ~x367 & ~x371 & ~x384 & ~x388 & ~x412 & ~x414 & ~x415 & ~x441 & ~x443 & ~x444 & ~x450 & ~x470 & ~x478 & ~x480 & ~x497 & ~x502 & ~x504 & ~x505 & ~x508 & ~x529 & ~x530 & ~x533 & ~x535 & ~x537 & ~x554 & ~x555 & ~x564 & ~x592 & ~x611 & ~x638 & ~x641 & ~x649 & ~x650 & ~x665 & ~x671 & ~x678 & ~x695 & ~x704 & ~x723 & ~x753 & ~x756 & ~x769 & ~x778 & ~x782;
assign c1212 =  x95 &  x151 &  x262 &  x270 &  x289 &  x298 &  x344 &  x353 &  x484 &  x579 &  x597 &  x607 &  x624 &  x656 &  x662 & ~x52 & ~x63 & ~x106 & ~x139 & ~x170 & ~x173 & ~x305 & ~x306 & ~x397 & ~x477 & ~x754;
assign c1214 =  x514 & ~x223 & ~x306 & ~x517 & ~x573 & ~x601 & ~x685 & ~x741;
assign c1216 =  x20;
assign c1218 = ~x0 & ~x1 & ~x2 & ~x3 & ~x4 & ~x5 & ~x6 & ~x7 & ~x8 & ~x9 & ~x18 & ~x19 & ~x20 & ~x21 & ~x22 & ~x23 & ~x24 & ~x25 & ~x26 & ~x27 & ~x28 & ~x29 & ~x30 & ~x31 & ~x32 & ~x33 & ~x34 & ~x35 & ~x36 & ~x48 & ~x49 & ~x50 & ~x51 & ~x52 & ~x53 & ~x54 & ~x55 & ~x56 & ~x57 & ~x58 & ~x59 & ~x60 & ~x61 & ~x62 & ~x63 & ~x64 & ~x76 & ~x77 & ~x78 & ~x79 & ~x80 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x86 & ~x87 & ~x88 & ~x89 & ~x90 & ~x91 & ~x92 & ~x104 & ~x105 & ~x106 & ~x107 & ~x108 & ~x109 & ~x110 & ~x111 & ~x112 & ~x113 & ~x114 & ~x115 & ~x116 & ~x117 & ~x118 & ~x119 & ~x120 & ~x132 & ~x133 & ~x134 & ~x135 & ~x136 & ~x137 & ~x138 & ~x139 & ~x140 & ~x141 & ~x142 & ~x143 & ~x144 & ~x145 & ~x146 & ~x147 & ~x148 & ~x160 & ~x161 & ~x162 & ~x163 & ~x164 & ~x165 & ~x166 & ~x167 & ~x168 & ~x169 & ~x170 & ~x171 & ~x172 & ~x173 & ~x174 & ~x175 & ~x188 & ~x189 & ~x190 & ~x191 & ~x192 & ~x193 & ~x194 & ~x195 & ~x196 & ~x197 & ~x198 & ~x199 & ~x200 & ~x201 & ~x202 & ~x203 & ~x204 & ~x215 & ~x216 & ~x217 & ~x218 & ~x219 & ~x220 & ~x221 & ~x222 & ~x223 & ~x224 & ~x225 & ~x226 & ~x227 & ~x228 & ~x229 & ~x230 & ~x231 & ~x232 & ~x243 & ~x244 & ~x245 & ~x246 & ~x247 & ~x248 & ~x249 & ~x250 & ~x251 & ~x252 & ~x253 & ~x254 & ~x255 & ~x256 & ~x257 & ~x258 & ~x259 & ~x260 & ~x272 & ~x273 & ~x274 & ~x275 & ~x276 & ~x277 & ~x278 & ~x279 & ~x280 & ~x281 & ~x282 & ~x283 & ~x284 & ~x285 & ~x286 & ~x287 & ~x288 & ~x299 & ~x300 & ~x301 & ~x302 & ~x303 & ~x304 & ~x305 & ~x306 & ~x307 & ~x308 & ~x309 & ~x310 & ~x311 & ~x312 & ~x313 & ~x314 & ~x315 & ~x316 & ~x328 & ~x329 & ~x330 & ~x331 & ~x332 & ~x333 & ~x334 & ~x335 & ~x336 & ~x337 & ~x338 & ~x339 & ~x340 & ~x341 & ~x342 & ~x343 & ~x355 & ~x356 & ~x357 & ~x358 & ~x359 & ~x360 & ~x361 & ~x362 & ~x363 & ~x364 & ~x365 & ~x366 & ~x367 & ~x368 & ~x369 & ~x370 & ~x371 & ~x372 & ~x383 & ~x384 & ~x385 & ~x386 & ~x387 & ~x388 & ~x389 & ~x390 & ~x391 & ~x392 & ~x393 & ~x394 & ~x395 & ~x396 & ~x397 & ~x398 & ~x399 & ~x400 & ~x411 & ~x412 & ~x413 & ~x414 & ~x415 & ~x416 & ~x417 & ~x418 & ~x419 & ~x420 & ~x421 & ~x422 & ~x423 & ~x424 & ~x425 & ~x426 & ~x427 & ~x428 & ~x439 & ~x440 & ~x441 & ~x442 & ~x443 & ~x444 & ~x445 & ~x446 & ~x447 & ~x448 & ~x449 & ~x450 & ~x451 & ~x452 & ~x453 & ~x454 & ~x455 & ~x456 & ~x467 & ~x468 & ~x469 & ~x470 & ~x471 & ~x472 & ~x473 & ~x474 & ~x475 & ~x476 & ~x477 & ~x478 & ~x479 & ~x480 & ~x481 & ~x482 & ~x483 & ~x484 & ~x495 & ~x496 & ~x497 & ~x498 & ~x499 & ~x500 & ~x501 & ~x502 & ~x503 & ~x504 & ~x505 & ~x506 & ~x507 & ~x508 & ~x509 & ~x510 & ~x511 & ~x512 & ~x523 & ~x524 & ~x525 & ~x526 & ~x527 & ~x528 & ~x529 & ~x531 & ~x532 & ~x533 & ~x534 & ~x535 & ~x536 & ~x537 & ~x539 & ~x540 & ~x551 & ~x552 & ~x553 & ~x554 & ~x555 & ~x556 & ~x557 & ~x558 & ~x559 & ~x560 & ~x561 & ~x562 & ~x563 & ~x564 & ~x565 & ~x566 & ~x567 & ~x568 & ~x579 & ~x580 & ~x581 & ~x582 & ~x583 & ~x584 & ~x585 & ~x586 & ~x587 & ~x588 & ~x589 & ~x590 & ~x591 & ~x592 & ~x593 & ~x594 & ~x595 & ~x596 & ~x606 & ~x607 & ~x608 & ~x609 & ~x610 & ~x611 & ~x612 & ~x613 & ~x614 & ~x615 & ~x616 & ~x617 & ~x618 & ~x619 & ~x620 & ~x621 & ~x622 & ~x623 & ~x624 & ~x636 & ~x637 & ~x638 & ~x639 & ~x640 & ~x641 & ~x642 & ~x643 & ~x644 & ~x645 & ~x646 & ~x647 & ~x648 & ~x649 & ~x650 & ~x651 & ~x652 & ~x663 & ~x664 & ~x665 & ~x666 & ~x667 & ~x668 & ~x669 & ~x670 & ~x671 & ~x672 & ~x673 & ~x674 & ~x675 & ~x676 & ~x677 & ~x678 & ~x679 & ~x680 & ~x692 & ~x693 & ~x694 & ~x695 & ~x696 & ~x697 & ~x698 & ~x699 & ~x700 & ~x701 & ~x702 & ~x703 & ~x704 & ~x705 & ~x706 & ~x707 & ~x708 & ~x709 & ~x720 & ~x721 & ~x722 & ~x723 & ~x724 & ~x725 & ~x726 & ~x727 & ~x728 & ~x729 & ~x730 & ~x731 & ~x732 & ~x733 & ~x736 & ~x748 & ~x749 & ~x750 & ~x751 & ~x752 & ~x753 & ~x754 & ~x755 & ~x756 & ~x757 & ~x758 & ~x759 & ~x760 & ~x761 & ~x762 & ~x763 & ~x764 & ~x765 & ~x766 & ~x774 & ~x775 & ~x776 & ~x777 & ~x778 & ~x779 & ~x780 & ~x781 & ~x782 & ~x783;
assign c1220 =  x396;
assign c1222 =  x644 &  x696;
assign c1224 = ~x59 & ~x88 & ~x115 & ~x165 & ~x166 & ~x304 & ~x389 & ~x434 & ~x462 & ~x489 & ~x490 & ~x503 & ~x518 & ~x545 & ~x546 & ~x562 & ~x574 & ~x601 & ~x602 & ~x629 & ~x630 & ~x657 & ~x658 & ~x685 & ~x686 & ~x713 & ~x741 & ~x742 & ~x769 & ~x770;
assign c1226 =  x26;
assign c1228 =  x40 &  x42 &  x44 &  x68 &  x69 &  x73 &  x98 &  x100 &  x124 &  x126 &  x127 &  x151 &  x155 &  x158 &  x180 &  x181 &  x182 &  x183 &  x186 &  x211 &  x212 &  x213 &  x234 &  x235 &  x240 &  x291 &  x297 &  x324 &  x352 &  x375 &  x403 &  x409 &  x515 &  x576 &  x713 & ~x0 & ~x2 & ~x3 & ~x7 & ~x8 & ~x31 & ~x51 & ~x52 & ~x54 & ~x56 & ~x59 & ~x77 & ~x81 & ~x84 & ~x87 & ~x90 & ~x107 & ~x115 & ~x117 & ~x119 & ~x140 & ~x164 & ~x169 & ~x170 & ~x171 & ~x172 & ~x190 & ~x191 & ~x193 & ~x195 & ~x197 & ~x201 & ~x219 & ~x220 & ~x226 & ~x227 & ~x230 & ~x246 & ~x250 & ~x253 & ~x254 & ~x258 & ~x279 & ~x282 & ~x285 & ~x302 & ~x309 & ~x311 & ~x335 & ~x365 & ~x367 & ~x369 & ~x370 & ~x389 & ~x396 & ~x413 & ~x416 & ~x420 & ~x421 & ~x427 & ~x441 & ~x445 & ~x453 & ~x454 & ~x469 & ~x474 & ~x476 & ~x482 & ~x483 & ~x497 & ~x501 & ~x508 & ~x511 & ~x531 & ~x533 & ~x553 & ~x560 & ~x562 & ~x565 & ~x589 & ~x591 & ~x615 & ~x616 & ~x617 & ~x620 & ~x623 & ~x637 & ~x641 & ~x645 & ~x647 & ~x649 & ~x672 & ~x679 & ~x694 & ~x698 & ~x703 & ~x704 & ~x705 & ~x707 & ~x720 & ~x721 & ~x733 & ~x735 & ~x753 & ~x757 & ~x758 & ~x776 & ~x778 & ~x779 & ~x782;
assign c1230 =  x39 &  x234 &  x262 & ~x1 & ~x37 & ~x50 & ~x61 & ~x63 & ~x65 & ~x77 & ~x79 & ~x84 & ~x88 & ~x90 & ~x91 & ~x110 & ~x116 & ~x146 & ~x174 & ~x196 & ~x217 & ~x224 & ~x226 & ~x229 & ~x250 & ~x257 & ~x275 & ~x277 & ~x279 & ~x302 & ~x304 & ~x308 & ~x309 & ~x367 & ~x370 & ~x386 & ~x388 & ~x397 & ~x444 & ~x446 & ~x447 & ~x476 & ~x479 & ~x484 & ~x499 & ~x502 & ~x527 & ~x533 & ~x536 & ~x552 & ~x553 & ~x557 & ~x562 & ~x580 & ~x581 & ~x584 & ~x585 & ~x592 & ~x608 & ~x610 & ~x621 & ~x636 & ~x638 & ~x640 & ~x644 & ~x646 & ~x648 & ~x650 & ~x652 & ~x666 & ~x667 & ~x671 & ~x704 & ~x705 & ~x721 & ~x728 & ~x748 & ~x758 & ~x761;
assign c1232 =  x11 &  x13 &  x70 &  x155 &  x206 &  x262 &  x264 &  x318 &  x324 &  x379 &  x604 &  x688 & ~x5 & ~x104 & ~x107 & ~x118 & ~x163 & ~x164 & ~x217 & ~x226 & ~x256 & ~x311 & ~x389 & ~x420 & ~x477 & ~x537 & ~x616 & ~x698;
assign c1234 =  x45 &  x74 &  x126 &  x156 &  x208 &  x209 &  x210 &  x237 &  x242 &  x263 &  x266 &  x268 &  x290 &  x291 &  x294 &  x295 &  x323 &  x345 &  x347 &  x349 &  x351 &  x355 &  x373 &  x400 &  x407 &  x411 &  x428 &  x429 &  x432 &  x435 &  x463 &  x484 &  x495 &  x512 &  x519 &  x523 &  x540 &  x547 &  x568 &  x624 &  x635 &  x680 &  x681 & ~x1 & ~x3 & ~x23 & ~x27 & ~x32 & ~x51 & ~x53 & ~x54 & ~x56 & ~x57 & ~x58 & ~x59 & ~x62 & ~x79 & ~x87 & ~x107 & ~x109 & ~x110 & ~x114 & ~x115 & ~x164 & ~x167 & ~x169 & ~x170 & ~x171 & ~x192 & ~x194 & ~x198 & ~x199 & ~x248 & ~x251 & ~x252 & ~x254 & ~x306 & ~x307 & ~x310 & ~x311 & ~x332 & ~x333 & ~x334 & ~x338 & ~x362 & ~x363 & ~x365 & ~x366 & ~x396 & ~x416 & ~x419 & ~x420 & ~x423 & ~x424 & ~x449 & ~x473 & ~x478 & ~x500 & ~x502 & ~x504 & ~x506 & ~x507 & ~x531 & ~x534 & ~x562 & ~x584 & ~x587 & ~x588 & ~x590 & ~x612 & ~x614 & ~x615 & ~x617 & ~x618 & ~x643 & ~x647 & ~x648 & ~x675 & ~x676 & ~x696 & ~x703 & ~x724 & ~x726 & ~x728 & ~x755 & ~x756 & ~x757 & ~x758 & ~x778 & ~x779 & ~x781 & ~x783;
assign c1236 =  x13 &  x17 &  x90;
assign c1238 =  x268 &  x292 &  x293 &  x431 &  x458 &  x487 &  x493 &  x543 &  x576 &  x605 &  x683 &  x684 &  x687 &  x715 &  x739 &  x744 &  x767 &  x768 &  x772 & ~x0 & ~x1 & ~x2 & ~x24 & ~x25 & ~x26 & ~x51 & ~x52 & ~x53 & ~x55 & ~x61 & ~x62 & ~x76 & ~x77 & ~x79 & ~x80 & ~x81 & ~x84 & ~x85 & ~x90 & ~x91 & ~x104 & ~x106 & ~x110 & ~x111 & ~x113 & ~x115 & ~x117 & ~x118 & ~x119 & ~x133 & ~x134 & ~x135 & ~x136 & ~x140 & ~x141 & ~x143 & ~x145 & ~x160 & ~x163 & ~x165 & ~x166 & ~x168 & ~x170 & ~x172 & ~x174 & ~x175 & ~x188 & ~x189 & ~x192 & ~x193 & ~x194 & ~x195 & ~x198 & ~x199 & ~x200 & ~x216 & ~x220 & ~x221 & ~x222 & ~x226 & ~x229 & ~x230 & ~x231 & ~x244 & ~x247 & ~x248 & ~x251 & ~x254 & ~x255 & ~x258 & ~x275 & ~x277 & ~x279 & ~x281 & ~x283 & ~x286 & ~x302 & ~x304 & ~x305 & ~x313 & ~x314 & ~x315 & ~x328 & ~x329 & ~x331 & ~x332 & ~x334 & ~x337 & ~x339 & ~x342 & ~x357 & ~x361 & ~x362 & ~x363 & ~x366 & ~x370 & ~x386 & ~x389 & ~x391 & ~x395 & ~x398 & ~x399 & ~x413 & ~x414 & ~x417 & ~x419 & ~x421 & ~x422 & ~x426 & ~x427 & ~x440 & ~x441 & ~x442 & ~x448 & ~x449 & ~x450 & ~x453 & ~x454 & ~x455 & ~x473 & ~x474 & ~x475 & ~x481 & ~x483 & ~x497 & ~x498 & ~x503 & ~x504 & ~x505 & ~x525 & ~x526 & ~x527 & ~x530 & ~x531 & ~x532 & ~x553 & ~x554 & ~x555 & ~x558 & ~x561 & ~x563 & ~x564 & ~x566 & ~x582 & ~x583 & ~x584 & ~x588 & ~x589 & ~x594 & ~x611 & ~x613 & ~x617 & ~x619 & ~x621 & ~x638 & ~x639 & ~x641 & ~x646 & ~x647 & ~x667 & ~x669 & ~x670 & ~x675 & ~x678 & ~x697 & ~x698 & ~x702 & ~x723 & ~x724 & ~x728 & ~x730 & ~x731 & ~x734 & ~x751 & ~x753 & ~x754 & ~x761 & ~x763 & ~x776 & ~x782 & ~x783;
assign c1240 =  x560;
assign c1242 =  x73 &  x267 &  x408 &  x521 &  x569 &  x595 &  x651 & ~x334 & ~x769;
assign c1244 =  x103 &  x748 & ~x490 & ~x574 & ~x602 & ~x743;
assign c1246 = ~x2 & ~x8 & ~x19 & ~x57 & ~x60 & ~x77 & ~x83 & ~x85 & ~x86 & ~x87 & ~x88 & ~x106 & ~x110 & ~x112 & ~x115 & ~x117 & ~x132 & ~x134 & ~x142 & ~x162 & ~x166 & ~x190 & ~x191 & ~x199 & ~x200 & ~x201 & ~x220 & ~x223 & ~x226 & ~x231 & ~x248 & ~x250 & ~x254 & ~x256 & ~x257 & ~x259 & ~x272 & ~x273 & ~x275 & ~x276 & ~x284 & ~x285 & ~x302 & ~x305 & ~x306 & ~x307 & ~x309 & ~x328 & ~x330 & ~x333 & ~x338 & ~x340 & ~x357 & ~x363 & ~x364 & ~x365 & ~x366 & ~x371 & ~x389 & ~x412 & ~x418 & ~x419 & ~x426 & ~x427 & ~x440 & ~x447 & ~x448 & ~x451 & ~x462 & ~x468 & ~x471 & ~x474 & ~x479 & ~x481 & ~x483 & ~x495 & ~x497 & ~x499 & ~x502 & ~x505 & ~x508 & ~x518 & ~x527 & ~x529 & ~x535 & ~x538 & ~x568 & ~x582 & ~x593 & ~x608 & ~x619 & ~x620 & ~x624 & ~x644 & ~x645 & ~x664 & ~x668 & ~x669 & ~x673 & ~x692 & ~x697 & ~x699 & ~x701 & ~x707 & ~x720 & ~x724 & ~x751 & ~x752 & ~x754 & ~x781;
assign c1248 =  x39 &  x68 &  x241 &  x572 &  x768 & ~x9 & ~x105 & ~x132 & ~x146 & ~x216 & ~x229 & ~x300 & ~x556 & ~x615 & ~x734;
assign c1250 =  x236 &  x320 &  x351 &  x402 &  x435 &  x459 &  x571 &  x627 &  x683 &  x767 &  x771 & ~x3 & ~x24 & ~x31 & ~x51 & ~x59 & ~x61 & ~x62 & ~x88 & ~x105 & ~x116 & ~x118 & ~x136 & ~x137 & ~x140 & ~x162 & ~x170 & ~x173 & ~x201 & ~x219 & ~x222 & ~x225 & ~x246 & ~x251 & ~x256 & ~x275 & ~x312 & ~x314 & ~x337 & ~x395 & ~x414 & ~x420 & ~x422 & ~x426 & ~x442 & ~x443 & ~x446 & ~x471 & ~x476 & ~x483 & ~x531 & ~x555 & ~x563 & ~x581 & ~x587 & ~x591 & ~x609 & ~x610 & ~x619 & ~x645 & ~x647 & ~x649 & ~x693 & ~x695 & ~x705 & ~x722 & ~x747 & ~x782 & ~x783;
assign c1252 =  x39 &  x745 & ~x26 & ~x115 & ~x163 & ~x172 & ~x247 & ~x253 & ~x284 & ~x304 & ~x444 & ~x445 & ~x447 & ~x474 & ~x527 & ~x584 & ~x621 & ~x658 & ~x686 & ~x701 & ~x742 & ~x757 & ~x759 & ~x760 & ~x770;
assign c1254 =  x238 &  x464 & ~x421 & ~x459;
assign c1256 = ~x133 & ~x241 & ~x245 & ~x246 & ~x252 & ~x272 & ~x276 & ~x297 & ~x336 & ~x367 & ~x383 & ~x409 & ~x453 & ~x465 & ~x466 & ~x480 & ~x502 & ~x552 & ~x776;
assign c1258 =  x44 &  x73 &  x99 &  x126 &  x153 &  x179 &  x180 &  x209 &  x212 &  x234 &  x237 &  x238 &  x261 &  x263 &  x266 &  x267 &  x290 &  x293 &  x295 &  x318 &  x322 &  x326 &  x344 &  x345 &  x346 &  x347 &  x349 &  x354 &  x375 &  x378 &  x381 &  x400 &  x405 &  x407 &  x409 &  x456 &  x457 &  x458 &  x460 &  x463 &  x466 &  x484 &  x485 &  x493 &  x549 &  x568 &  x569 &  x577 &  x596 &  x607 &  x652 &  x654 &  x680 &  x681 &  x715 & ~x1 & ~x3 & ~x6 & ~x27 & ~x32 & ~x34 & ~x56 & ~x58 & ~x59 & ~x61 & ~x82 & ~x85 & ~x110 & ~x114 & ~x117 & ~x138 & ~x143 & ~x164 & ~x165 & ~x172 & ~x193 & ~x197 & ~x198 & ~x221 & ~x222 & ~x223 & ~x226 & ~x284 & ~x304 & ~x305 & ~x306 & ~x310 & ~x335 & ~x364 & ~x365 & ~x366 & ~x368 & ~x390 & ~x391 & ~x393 & ~x418 & ~x419 & ~x444 & ~x501 & ~x502 & ~x535 & ~x536 & ~x556 & ~x560 & ~x561 & ~x584 & ~x588 & ~x614 & ~x619 & ~x640 & ~x645 & ~x671 & ~x673 & ~x676 & ~x702 & ~x703 & ~x704 & ~x725 & ~x727 & ~x729 & ~x760 & ~x779 & ~x780 & ~x782;
assign c1260 =  x39 &  x100 &  x124 &  x152 &  x155 &  x179 &  x213 &  x240 &  x291 &  x346 &  x402 &  x548 &  x712 & ~x48 & ~x55 & ~x76 & ~x88 & ~x90 & ~x107 & ~x142 & ~x144 & ~x146 & ~x168 & ~x172 & ~x217 & ~x230 & ~x256 & ~x273 & ~x329 & ~x338 & ~x362 & ~x370 & ~x387 & ~x419 & ~x427 & ~x453 & ~x511 & ~x609 & ~x616 & ~x640 & ~x648 & ~x699 & ~x708 & ~x755 & ~x783;
assign c1262 =  x254 &  x588;
assign c1264 =  x95 &  x96 &  x98 &  x100 &  x128 &  x151 &  x155 &  x156 &  x179 &  x210 &  x268 &  x297 &  x298 &  x326 &  x381 &  x465 &  x487 &  x685 & ~x3 & ~x19 & ~x36 & ~x56 & ~x76 & ~x77 & ~x78 & ~x87 & ~x117 & ~x132 & ~x140 & ~x162 & ~x170 & ~x193 & ~x200 & ~x252 & ~x276 & ~x308 & ~x334 & ~x335 & ~x392 & ~x420 & ~x447 & ~x474 & ~x482 & ~x501 & ~x534 & ~x553 & ~x561 & ~x584 & ~x587 & ~x588 & ~x594 & ~x639 & ~x641 & ~x645 & ~x647 & ~x649 & ~x670 & ~x706 & ~x758 & ~x780;
assign c1266 =  x46 &  x123 &  x212 &  x238 &  x356 &  x399 &  x457 &  x467 &  x652 &  x653 & ~x28 & ~x248 & ~x417 & ~x423 & ~x672;
assign c1268 =  x9 & ~x34 & ~x49 & ~x57 & ~x77 & ~x105 & ~x106 & ~x117 & ~x144 & ~x168 & ~x197 & ~x274 & ~x276 & ~x305 & ~x358 & ~x418 & ~x421 & ~x498 & ~x500 & ~x612;
assign c1270 =  x43 &  x44 &  x47 &  x72 &  x154 &  x155 &  x159 &  x186 &  x242 &  x299 & ~x60 & ~x61 & ~x79 & ~x84 & ~x193 & ~x391 & ~x417 & ~x422 & ~x444 & ~x505 & ~x506 & ~x640 & ~x722 & ~x748 & ~x750 & ~x751 & ~x755 & ~x760 & ~x776;
assign c1272 = ~x629;
assign c1274 =  x2;
assign c1276 =  x598 & ~x1 & ~x3 & ~x5 & ~x27 & ~x28 & ~x33 & ~x54 & ~x80 & ~x82 & ~x86 & ~x88 & ~x107 & ~x110 & ~x111 & ~x114 & ~x115 & ~x136 & ~x141 & ~x145 & ~x163 & ~x167 & ~x172 & ~x191 & ~x193 & ~x199 & ~x219 & ~x221 & ~x227 & ~x249 & ~x252 & ~x253 & ~x276 & ~x279 & ~x282 & ~x306 & ~x308 & ~x312 & ~x331 & ~x332 & ~x334 & ~x336 & ~x337 & ~x360 & ~x362 & ~x388 & ~x392 & ~x395 & ~x418 & ~x420 & ~x444 & ~x446 & ~x447 & ~x452 & ~x472 & ~x474 & ~x476 & ~x502 & ~x504 & ~x505 & ~x506 & ~x508 & ~x535 & ~x560 & ~x561 & ~x562 & ~x563 & ~x584 & ~x587 & ~x601 & ~x613 & ~x616 & ~x617 & ~x619 & ~x629 & ~x640 & ~x646 & ~x647 & ~x667 & ~x668 & ~x670 & ~x671 & ~x676 & ~x695 & ~x696 & ~x700 & ~x702 & ~x724 & ~x726 & ~x727 & ~x731 & ~x741 & ~x751 & ~x754 & ~x758 & ~x762 & ~x769 & ~x780 & ~x783;
assign c1278 = ~x90 & ~x100 & ~x167 & ~x175 & ~x188 & ~x230 & ~x249 & ~x304 & ~x325 & ~x344 & ~x368 & ~x411 & ~x468 & ~x607 & ~x669 & ~x720 & ~x723 & ~x725 & ~x765;
assign c1280 = ~x2 & ~x8 & ~x23 & ~x33 & ~x62 & ~x63 & ~x108 & ~x136 & ~x140 & ~x162 & ~x166 & ~x190 & ~x203 & ~x219 & ~x220 & ~x224 & ~x229 & ~x246 & ~x248 & ~x252 & ~x255 & ~x259 & ~x260 & ~x272 & ~x283 & ~x285 & ~x286 & ~x287 & ~x299 & ~x300 & ~x302 & ~x329 & ~x337 & ~x342 & ~x345 & ~x356 & ~x357 & ~x370 & ~x387 & ~x389 & ~x392 & ~x400 & ~x401 & ~x411 & ~x425 & ~x427 & ~x429 & ~x445 & ~x446 & ~x447 & ~x455 & ~x457 & ~x472 & ~x474 & ~x479 & ~x480 & ~x482 & ~x495 & ~x506 & ~x508 & ~x523 & ~x528 & ~x542 & ~x552 & ~x558 & ~x560 & ~x562 & ~x563 & ~x564 & ~x566 & ~x567 & ~x583 & ~x586 & ~x588 & ~x593 & ~x609 & ~x616 & ~x626 & ~x643 & ~x649 & ~x662 & ~x674 & ~x679 & ~x681 & ~x694 & ~x695 & ~x705 & ~x718 & ~x722 & ~x726 & ~x754 & ~x774;
assign c1282 =  x25;
assign c1284 =  x571 & ~x117 & ~x249 & ~x283 & ~x361 & ~x497 & ~x545 & ~x581 & ~x629 & ~x685 & ~x693 & ~x713 & ~x741 & ~x783;
assign c1286 =  x154 &  x209 &  x240 &  x493 &  x605 & ~x3 & ~x21 & ~x57 & ~x62 & ~x87 & ~x135 & ~x203 & ~x389 & ~x417 & ~x475 & ~x497 & ~x502 & ~x539 & ~x574 & ~x587 & ~x595 & ~x652 & ~x761;
assign c1288 =  x150 &  x155 &  x430 & ~x5 & ~x52 & ~x278 & ~x338 & ~x362 & ~x517;
assign c1290 =  x48 &  x764;
assign c1292 =  x283 &  x765;
assign c1294 =  x154 &  x210 &  x599 & ~x7 & ~x26 & ~x60 & ~x62 & ~x139 & ~x163 & ~x370 & ~x418 & ~x420 & ~x450 & ~x480 & ~x509 & ~x530 & ~x602 & ~x643 & ~x651 & ~x671 & ~x673 & ~x694 & ~x699 & ~x761 & ~x776;
assign c1296 =  x57;
assign c1298 =  x644;
assign c1300 =  x593 & ~x602 & ~x629;
assign c1302 =  x373 &  x541 &  x547 &  x603 & ~x56 & ~x103 & ~x104 & ~x132 & ~x284 & ~x479 & ~x554 & ~x769;
assign c1304 =  x338;
assign c1306 =  x12 &  x14 &  x15 &  x16 &  x17 &  x96 &  x99 &  x205 &  x318 & ~x32 & ~x60 & ~x108 & ~x136 & ~x143 & ~x165 & ~x167 & ~x222 & ~x277 & ~x363 & ~x391 & ~x422 & ~x501 & ~x505 & ~x528 & ~x559 & ~x562 & ~x590 & ~x618 & ~x695 & ~x702 & ~x777;
assign c1308 =  x211 &  x240 &  x263 &  x295 &  x322 &  x347 &  x381 &  x409 &  x431 &  x432 &  x435 &  x464 &  x487 &  x493 &  x600 &  x603 &  x627 &  x628 &  x656 &  x683 &  x684 &  x687 &  x689 &  x716 &  x744 &  x768 &  x772 &  x773 & ~x3 & ~x26 & ~x27 & ~x31 & ~x34 & ~x78 & ~x83 & ~x87 & ~x106 & ~x115 & ~x118 & ~x145 & ~x161 & ~x165 & ~x167 & ~x193 & ~x196 & ~x197 & ~x203 & ~x217 & ~x247 & ~x283 & ~x305 & ~x314 & ~x336 & ~x393 & ~x395 & ~x416 & ~x417 & ~x421 & ~x423 & ~x451 & ~x473 & ~x476 & ~x500 & ~x508 & ~x533 & ~x538 & ~x553 & ~x560 & ~x589 & ~x592 & ~x593 & ~x638 & ~x702 & ~x705 & ~x727 & ~x728 & ~x751 & ~x757;
assign c1310 =  x95 &  x208 &  x211 &  x262 &  x403 &  x458 &  x543 &  x655 &  x683 &  x711 & ~x0 & ~x3 & ~x24 & ~x85 & ~x89 & ~x109 & ~x110 & ~x146 & ~x168 & ~x169 & ~x171 & ~x189 & ~x196 & ~x200 & ~x202 & ~x225 & ~x227 & ~x257 & ~x273 & ~x278 & ~x284 & ~x335 & ~x361 & ~x389 & ~x392 & ~x416 & ~x475 & ~x501 & ~x503 & ~x505 & ~x564 & ~x592 & ~x618 & ~x642 & ~x643 & ~x648 & ~x692 & ~x693 & ~x723 & ~x724 & ~x730 & ~x769 & ~x780;
assign c1312 = ~x0 & ~x1 & ~x3 & ~x4 & ~x7 & ~x8 & ~x19 & ~x22 & ~x25 & ~x30 & ~x31 & ~x34 & ~x35 & ~x49 & ~x51 & ~x53 & ~x55 & ~x56 & ~x58 & ~x59 & ~x60 & ~x80 & ~x84 & ~x85 & ~x86 & ~x87 & ~x90 & ~x91 & ~x103 & ~x104 & ~x105 & ~x109 & ~x110 & ~x112 & ~x113 & ~x115 & ~x116 & ~x132 & ~x133 & ~x135 & ~x136 & ~x140 & ~x141 & ~x142 & ~x143 & ~x144 & ~x160 & ~x161 & ~x163 & ~x166 & ~x167 & ~x168 & ~x171 & ~x172 & ~x173 & ~x175 & ~x188 & ~x190 & ~x191 & ~x194 & ~x200 & ~x201 & ~x202 & ~x203 & ~x218 & ~x219 & ~x220 & ~x221 & ~x222 & ~x224 & ~x225 & ~x227 & ~x228 & ~x230 & ~x231 & ~x245 & ~x248 & ~x249 & ~x250 & ~x251 & ~x253 & ~x254 & ~x257 & ~x258 & ~x259 & ~x260 & ~x276 & ~x277 & ~x278 & ~x282 & ~x283 & ~x285 & ~x286 & ~x287 & ~x288 & ~x301 & ~x302 & ~x306 & ~x307 & ~x308 & ~x311 & ~x312 & ~x313 & ~x316 & ~x328 & ~x330 & ~x333 & ~x334 & ~x335 & ~x337 & ~x338 & ~x339 & ~x342 & ~x343 & ~x356 & ~x358 & ~x365 & ~x366 & ~x368 & ~x369 & ~x370 & ~x372 & ~x385 & ~x386 & ~x387 & ~x390 & ~x391 & ~x394 & ~x395 & ~x398 & ~x399 & ~x400 & ~x412 & ~x413 & ~x414 & ~x417 & ~x419 & ~x423 & ~x427 & ~x441 & ~x444 & ~x445 & ~x446 & ~x452 & ~x455 & ~x468 & ~x469 & ~x472 & ~x474 & ~x475 & ~x476 & ~x478 & ~x480 & ~x483 & ~x497 & ~x498 & ~x500 & ~x501 & ~x502 & ~x503 & ~x504 & ~x506 & ~x507 & ~x508 & ~x510 & ~x523 & ~x524 & ~x526 & ~x529 & ~x530 & ~x532 & ~x534 & ~x538 & ~x540 & ~x551 & ~x553 & ~x555 & ~x556 & ~x557 & ~x562 & ~x563 & ~x565 & ~x568 & ~x582 & ~x584 & ~x586 & ~x588 & ~x589 & ~x592 & ~x593 & ~x594 & ~x595 & ~x606 & ~x607 & ~x609 & ~x611 & ~x612 & ~x614 & ~x615 & ~x617 & ~x618 & ~x623 & ~x624 & ~x634 & ~x637 & ~x638 & ~x639 & ~x640 & ~x641 & ~x642 & ~x643 & ~x644 & ~x645 & ~x648 & ~x649 & ~x650 & ~x652 & ~x664 & ~x665 & ~x667 & ~x668 & ~x669 & ~x670 & ~x671 & ~x672 & ~x675 & ~x676 & ~x677 & ~x678 & ~x680 & ~x690 & ~x692 & ~x695 & ~x699 & ~x700 & ~x701 & ~x702 & ~x703 & ~x705 & ~x719 & ~x722 & ~x724 & ~x725 & ~x727 & ~x730 & ~x733 & ~x735 & ~x750 & ~x751 & ~x754 & ~x756 & ~x758 & ~x759 & ~x762 & ~x764 & ~x765 & ~x769 & ~x775 & ~x776 & ~x778 & ~x779;
assign c1314 =  x209 &  x431 &  x487 &  x543 &  x571 &  x605 &  x627 &  x632 &  x660 &  x683 &  x684 &  x711 &  x717 & ~x0 & ~x1 & ~x3 & ~x4 & ~x6 & ~x7 & ~x8 & ~x21 & ~x22 & ~x23 & ~x24 & ~x27 & ~x30 & ~x32 & ~x33 & ~x48 & ~x49 & ~x50 & ~x51 & ~x52 & ~x53 & ~x56 & ~x58 & ~x59 & ~x61 & ~x64 & ~x77 & ~x78 & ~x79 & ~x82 & ~x83 & ~x85 & ~x86 & ~x87 & ~x88 & ~x89 & ~x104 & ~x105 & ~x107 & ~x109 & ~x112 & ~x113 & ~x114 & ~x115 & ~x116 & ~x117 & ~x119 & ~x133 & ~x135 & ~x136 & ~x137 & ~x138 & ~x140 & ~x141 & ~x142 & ~x145 & ~x160 & ~x164 & ~x165 & ~x166 & ~x167 & ~x172 & ~x189 & ~x191 & ~x193 & ~x195 & ~x197 & ~x199 & ~x200 & ~x201 & ~x202 & ~x218 & ~x222 & ~x224 & ~x225 & ~x226 & ~x229 & ~x230 & ~x244 & ~x246 & ~x247 & ~x248 & ~x249 & ~x250 & ~x252 & ~x253 & ~x254 & ~x255 & ~x256 & ~x257 & ~x273 & ~x274 & ~x275 & ~x277 & ~x278 & ~x281 & ~x282 & ~x284 & ~x285 & ~x301 & ~x302 & ~x303 & ~x308 & ~x309 & ~x310 & ~x311 & ~x314 & ~x329 & ~x330 & ~x333 & ~x334 & ~x335 & ~x338 & ~x341 & ~x342 & ~x359 & ~x360 & ~x362 & ~x363 & ~x364 & ~x365 & ~x366 & ~x367 & ~x368 & ~x369 & ~x388 & ~x390 & ~x391 & ~x394 & ~x395 & ~x396 & ~x398 & ~x415 & ~x417 & ~x418 & ~x419 & ~x420 & ~x421 & ~x422 & ~x423 & ~x424 & ~x425 & ~x442 & ~x444 & ~x448 & ~x452 & ~x470 & ~x471 & ~x472 & ~x474 & ~x475 & ~x478 & ~x481 & ~x501 & ~x502 & ~x503 & ~x504 & ~x505 & ~x508 & ~x526 & ~x527 & ~x528 & ~x529 & ~x532 & ~x533 & ~x534 & ~x535 & ~x536 & ~x557 & ~x558 & ~x559 & ~x564 & ~x566 & ~x582 & ~x584 & ~x585 & ~x588 & ~x589 & ~x590 & ~x591 & ~x593 & ~x612 & ~x614 & ~x615 & ~x618 & ~x619 & ~x621 & ~x638 & ~x640 & ~x642 & ~x643 & ~x644 & ~x648 & ~x649 & ~x667 & ~x668 & ~x669 & ~x670 & ~x671 & ~x674 & ~x675 & ~x679 & ~x695 & ~x697 & ~x698 & ~x699 & ~x701 & ~x704 & ~x705 & ~x707 & ~x723 & ~x724 & ~x725 & ~x726 & ~x727 & ~x728 & ~x729 & ~x730 & ~x750 & ~x751 & ~x756 & ~x757 & ~x759 & ~x761 & ~x770 & ~x778 & ~x779 & ~x781 & ~x783;
assign c1316 =  x128 &  x210 &  x212 &  x213 &  x235 &  x236 &  x237 &  x239 &  x241 &  x269 &  x325 &  x376 &  x685 &  x741 & ~x27 & ~x28 & ~x36 & ~x53 & ~x56 & ~x57 & ~x58 & ~x59 & ~x85 & ~x110 & ~x117 & ~x119 & ~x136 & ~x144 & ~x147 & ~x167 & ~x175 & ~x176 & ~x219 & ~x227 & ~x228 & ~x229 & ~x231 & ~x252 & ~x255 & ~x259 & ~x282 & ~x288 & ~x303 & ~x304 & ~x311 & ~x315 & ~x316 & ~x357 & ~x359 & ~x360 & ~x367 & ~x372 & ~x388 & ~x391 & ~x392 & ~x399 & ~x415 & ~x416 & ~x424 & ~x428 & ~x442 & ~x444 & ~x449 & ~x453 & ~x454 & ~x456 & ~x508 & ~x509 & ~x512 & ~x513 & ~x525 & ~x534 & ~x536 & ~x553 & ~x555 & ~x561 & ~x589 & ~x595 & ~x596 & ~x643 & ~x652 & ~x678 & ~x680 & ~x708 & ~x730 & ~x731 & ~x748 & ~x754;
assign c1318 =  x588;
assign c1320 =  x13 &  x19 & ~x79;
assign c1322 =  x238 &  x294 &  x463 &  x598 &  x710 & ~x26 & ~x52 & ~x55 & ~x58 & ~x88 & ~x110 & ~x168 & ~x169 & ~x193 & ~x196 & ~x199 & ~x227 & ~x305 & ~x308 & ~x310 & ~x418 & ~x473 & ~x474 & ~x529 & ~x531 & ~x562 & ~x590 & ~x614 & ~x615 & ~x641 & ~x686 & ~x702 & ~x756 & ~x770;
assign c1324 =  x765 & ~x329 & ~x388 & ~x445 & ~x769;
assign c1326 =  x45 &  x210 &  x294 &  x355 &  x662 &  x747 &  x748;
assign c1328 =  x279;
assign c1330 =  x27;
assign c1332 =  x103 &  x131 & ~x574 & ~x602 & ~x658 & ~x713;
assign c1334 =  x238 &  x408 & ~x136 & ~x144 & ~x249 & ~x305 & ~x310 & ~x518 & ~x546 & ~x574 & ~x602 & ~x771;
assign c1336 =  x43 &  x44 &  x73 &  x127 &  x129 &  x177 &  x242 &  x271 &  x296 &  x298 &  x317 &  x327 &  x345 &  x430 &  x551 &  x738 & ~x27 & ~x88 & ~x107 & ~x144 & ~x161 & ~x164 & ~x172 & ~x246 & ~x363 & ~x502 & ~x508 & ~x510 & ~x565 & ~x645 & ~x730;
assign c1338 = ~x353 & ~x437 & ~x465 & ~x571 & ~x627 & ~x739;
assign c1340 =  x10 &  x12 &  x127 & ~x24 & ~x63 & ~x106 & ~x134 & ~x145 & ~x170 & ~x245 & ~x303 & ~x359 & ~x613 & ~x673;
assign c1342 =  x11 &  x14 &  x213 & ~x52 & ~x54 & ~x64 & ~x287 & ~x339 & ~x363 & ~x368 & ~x504 & ~x562 & ~x615 & ~x647 & ~x752 & ~x779;
assign c1344 =  x69 & ~x171 & ~x173 & ~x585 & ~x711 & ~x722 & ~x767;
assign c1346 =  x20 &  x231 &  x343 &  x356;
assign c1348 =  x38 &  x42 &  x121 &  x205 &  x233 & ~x48 & ~x77 & ~x104 & ~x114 & ~x132 & ~x141 & ~x145 & ~x163 & ~x173 & ~x189 & ~x190 & ~x217 & ~x218 & ~x244 & ~x315 & ~x331 & ~x338 & ~x339 & ~x385 & ~x419 & ~x480 & ~x537 & ~x556 & ~x559 & ~x616 & ~x648 & ~x673 & ~x695 & ~x723 & ~x729 & ~x731 & ~x755;
assign c1350 =  x10 &  x12 & ~x216 & ~x217 & ~x255 & ~x277 & ~x283 & ~x385 & ~x478 & ~x498 & ~x780;
assign c1352 =  x98 &  x578 &  x662 & ~x558 & ~x574;
assign c1354 =  x747 & ~x686 & ~x714 & ~x742;
assign c1356 =  x184 &  x207 &  x483 &  x516 &  x524 &  x680 &  x681 &  x735;
assign c1358 =  x622 & ~x601 & ~x629 & ~x658 & ~x741 & ~x769;
assign c1360 =  x42 &  x45 &  x102 &  x213 &  x629 &  x713 & ~x1 & ~x6 & ~x7 & ~x8 & ~x20 & ~x21 & ~x28 & ~x30 & ~x31 & ~x32 & ~x34 & ~x53 & ~x57 & ~x58 & ~x78 & ~x79 & ~x81 & ~x83 & ~x86 & ~x108 & ~x114 & ~x115 & ~x120 & ~x134 & ~x142 & ~x162 & ~x164 & ~x165 & ~x167 & ~x168 & ~x171 & ~x190 & ~x192 & ~x197 & ~x218 & ~x221 & ~x247 & ~x253 & ~x254 & ~x256 & ~x258 & ~x277 & ~x307 & ~x309 & ~x310 & ~x335 & ~x336 & ~x360 & ~x361 & ~x368 & ~x387 & ~x391 & ~x398 & ~x425 & ~x426 & ~x443 & ~x447 & ~x449 & ~x452 & ~x453 & ~x470 & ~x475 & ~x481 & ~x482 & ~x483 & ~x497 & ~x501 & ~x504 & ~x505 & ~x508 & ~x510 & ~x532 & ~x534 & ~x555 & ~x582 & ~x592 & ~x620 & ~x623 & ~x638 & ~x643 & ~x645 & ~x650 & ~x651 & ~x666 & ~x667 & ~x668 & ~x672 & ~x674 & ~x676 & ~x678 & ~x679 & ~x692 & ~x696 & ~x700 & ~x703 & ~x706 & ~x707 & ~x726 & ~x727 & ~x729 & ~x735 & ~x748 & ~x756 & ~x760 & ~x762;
assign c1362 =  x560;
assign c1364 =  x637 & ~x571;
assign c1366 =  x42 &  x241 &  x351 &  x576 & ~x2 & ~x3 & ~x34 & ~x57 & ~x80 & ~x82 & ~x91 & ~x107 & ~x119 & ~x135 & ~x143 & ~x167 & ~x170 & ~x172 & ~x175 & ~x195 & ~x219 & ~x223 & ~x226 & ~x228 & ~x231 & ~x252 & ~x259 & ~x300 & ~x308 & ~x312 & ~x336 & ~x344 & ~x363 & ~x368 & ~x391 & ~x413 & ~x414 & ~x419 & ~x420 & ~x421 & ~x422 & ~x423 & ~x426 & ~x440 & ~x453 & ~x454 & ~x468 & ~x470 & ~x482 & ~x484 & ~x523 & ~x533 & ~x556 & ~x559 & ~x566 & ~x568 & ~x589 & ~x635 & ~x638 & ~x663 & ~x668 & ~x670 & ~x680 & ~x701 & ~x707 & ~x708 & ~x719 & ~x727 & ~x729 & ~x751 & ~x753 & ~x755 & ~x774 & ~x778;
assign c1368 =  x69 &  x71 &  x72 &  x99 &  x100 &  x123 &  x128 &  x154 &  x179 &  x209 &  x212 &  x236 &  x240 &  x242 &  x264 &  x265 &  x266 &  x321 &  x325 &  x348 &  x352 &  x353 &  x377 &  x380 &  x409 &  x437 &  x464 &  x521 &  x633 & ~x3 & ~x4 & ~x7 & ~x27 & ~x28 & ~x36 & ~x52 & ~x53 & ~x55 & ~x58 & ~x61 & ~x63 & ~x80 & ~x85 & ~x89 & ~x105 & ~x106 & ~x107 & ~x110 & ~x111 & ~x113 & ~x114 & ~x117 & ~x118 & ~x119 & ~x134 & ~x139 & ~x146 & ~x162 & ~x164 & ~x165 & ~x168 & ~x169 & ~x174 & ~x189 & ~x192 & ~x195 & ~x196 & ~x197 & ~x202 & ~x217 & ~x219 & ~x221 & ~x222 & ~x225 & ~x226 & ~x228 & ~x248 & ~x251 & ~x252 & ~x256 & ~x258 & ~x274 & ~x275 & ~x276 & ~x280 & ~x283 & ~x329 & ~x332 & ~x334 & ~x338 & ~x363 & ~x368 & ~x387 & ~x388 & ~x393 & ~x414 & ~x415 & ~x419 & ~x427 & ~x442 & ~x443 & ~x445 & ~x446 & ~x447 & ~x448 & ~x449 & ~x452 & ~x453 & ~x454 & ~x468 & ~x473 & ~x477 & ~x482 & ~x496 & ~x497 & ~x501 & ~x503 & ~x504 & ~x508 & ~x511 & ~x526 & ~x527 & ~x528 & ~x529 & ~x533 & ~x535 & ~x536 & ~x539 & ~x552 & ~x553 & ~x555 & ~x557 & ~x563 & ~x582 & ~x584 & ~x586 & ~x587 & ~x590 & ~x593 & ~x610 & ~x611 & ~x620 & ~x623 & ~x637 & ~x641 & ~x643 & ~x644 & ~x664 & ~x665 & ~x670 & ~x672 & ~x673 & ~x674 & ~x677 & ~x678 & ~x692 & ~x693 & ~x698 & ~x699 & ~x701 & ~x702 & ~x704 & ~x720 & ~x727 & ~x728 & ~x729 & ~x749 & ~x750 & ~x757 & ~x758 & ~x759 & ~x763 & ~x777 & ~x779 & ~x781;
assign c1370 =  x211 &  x351 &  x405 &  x407 &  x435 &  x463 &  x486 &  x491 &  x519 &  x547 &  x549 &  x570 &  x598 &  x603 &  x604 &  x605 &  x628 &  x661 &  x682 &  x688 &  x710 &  x717 &  x738 &  x740 &  x744 &  x772 & ~x0 & ~x1 & ~x2 & ~x3 & ~x4 & ~x5 & ~x6 & ~x7 & ~x20 & ~x21 & ~x22 & ~x23 & ~x24 & ~x25 & ~x27 & ~x28 & ~x29 & ~x30 & ~x34 & ~x48 & ~x50 & ~x52 & ~x54 & ~x55 & ~x56 & ~x57 & ~x59 & ~x60 & ~x61 & ~x77 & ~x78 & ~x79 & ~x80 & ~x81 & ~x82 & ~x84 & ~x86 & ~x87 & ~x88 & ~x90 & ~x91 & ~x105 & ~x107 & ~x108 & ~x109 & ~x110 & ~x111 & ~x112 & ~x115 & ~x116 & ~x118 & ~x133 & ~x134 & ~x136 & ~x137 & ~x138 & ~x139 & ~x140 & ~x141 & ~x142 & ~x144 & ~x146 & ~x161 & ~x163 & ~x164 & ~x165 & ~x166 & ~x167 & ~x169 & ~x170 & ~x171 & ~x173 & ~x174 & ~x189 & ~x190 & ~x191 & ~x192 & ~x193 & ~x194 & ~x195 & ~x197 & ~x198 & ~x199 & ~x202 & ~x217 & ~x218 & ~x219 & ~x222 & ~x225 & ~x226 & ~x227 & ~x228 & ~x229 & ~x230 & ~x245 & ~x249 & ~x250 & ~x251 & ~x253 & ~x254 & ~x255 & ~x256 & ~x257 & ~x258 & ~x274 & ~x275 & ~x277 & ~x279 & ~x280 & ~x281 & ~x282 & ~x283 & ~x284 & ~x285 & ~x286 & ~x302 & ~x303 & ~x304 & ~x305 & ~x306 & ~x310 & ~x313 & ~x314 & ~x329 & ~x330 & ~x332 & ~x333 & ~x335 & ~x336 & ~x339 & ~x340 & ~x341 & ~x342 & ~x358 & ~x359 & ~x361 & ~x362 & ~x364 & ~x365 & ~x367 & ~x369 & ~x386 & ~x387 & ~x389 & ~x390 & ~x391 & ~x393 & ~x394 & ~x396 & ~x397 & ~x398 & ~x415 & ~x417 & ~x418 & ~x420 & ~x421 & ~x422 & ~x425 & ~x426 & ~x442 & ~x444 & ~x445 & ~x446 & ~x447 & ~x448 & ~x449 & ~x450 & ~x451 & ~x453 & ~x471 & ~x472 & ~x473 & ~x478 & ~x479 & ~x481 & ~x482 & ~x498 & ~x499 & ~x500 & ~x505 & ~x507 & ~x508 & ~x509 & ~x510 & ~x526 & ~x529 & ~x530 & ~x531 & ~x532 & ~x533 & ~x534 & ~x535 & ~x536 & ~x537 & ~x538 & ~x554 & ~x555 & ~x557 & ~x559 & ~x560 & ~x563 & ~x564 & ~x581 & ~x582 & ~x585 & ~x587 & ~x588 & ~x589 & ~x590 & ~x591 & ~x592 & ~x593 & ~x594 & ~x610 & ~x611 & ~x612 & ~x613 & ~x614 & ~x615 & ~x618 & ~x619 & ~x620 & ~x622 & ~x639 & ~x640 & ~x641 & ~x643 & ~x645 & ~x650 & ~x666 & ~x667 & ~x668 & ~x669 & ~x670 & ~x671 & ~x673 & ~x674 & ~x675 & ~x694 & ~x698 & ~x700 & ~x701 & ~x702 & ~x704 & ~x705 & ~x722 & ~x723 & ~x724 & ~x725 & ~x726 & ~x727 & ~x728 & ~x729 & ~x730 & ~x731 & ~x732 & ~x751 & ~x752 & ~x753 & ~x756 & ~x757 & ~x758 & ~x759 & ~x760 & ~x761 & ~x762 & ~x763 & ~x770 & ~x776 & ~x779 & ~x780 & ~x783;
assign c1372 =  x478 &  x534;
assign c1374 =  x10 & ~x321;
assign c1376 = ~x12 & ~x71 & ~x191 & ~x301 & ~x382 & ~x387 & ~x397 & ~x580 & ~x664 & ~x770;
assign c1378 =  x260 &  x291 &  x440 & ~x52 & ~x80;
assign c1380 =  x42 &  x126 &  x155 &  x261 &  x267 &  x289 &  x438 &  x519 & ~x21 & ~x29 & ~x55 & ~x60 & ~x61 & ~x63 & ~x77 & ~x118 & ~x136 & ~x142 & ~x173 & ~x199 & ~x225 & ~x226 & ~x247 & ~x301 & ~x302 & ~x336 & ~x392 & ~x394 & ~x426 & ~x481 & ~x553 & ~x564 & ~x566 & ~x584 & ~x666 & ~x667 & ~x758 & ~x763 & ~x778;
assign c1382 =  x146 & ~x165 & ~x517 & ~x546 & ~x574 & ~x629 & ~x658 & ~x686 & ~x712 & ~x714 & ~x741 & ~x768;
assign c1384 =  x68 &  x156 &  x289 &  x298 &  x373 &  x633 & ~x217 & ~x594 & ~x764;
assign c1386 =  x72 &  x269 &  x295 &  x326 &  x437 &  x577 & ~x32 & ~x77 & ~x118 & ~x136 & ~x164 & ~x224 & ~x227 & ~x245 & ~x334 & ~x341 & ~x385 & ~x386 & ~x390 & ~x440 & ~x483 & ~x534 & ~x553 & ~x563 & ~x608 & ~x624 & ~x644 & ~x692 & ~x708 & ~x726;
assign c1388 =  x756;
assign c1390 =  x20 &  x97 &  x286;
assign c1392 = ~x1 & ~x8 & ~x22 & ~x32 & ~x50 & ~x57 & ~x84 & ~x108 & ~x117 & ~x135 & ~x138 & ~x143 & ~x165 & ~x170 & ~x171 & ~x173 & ~x174 & ~x190 & ~x195 & ~x197 & ~x199 & ~x200 & ~x217 & ~x221 & ~x227 & ~x245 & ~x247 & ~x253 & ~x255 & ~x272 & ~x273 & ~x277 & ~x304 & ~x330 & ~x331 & ~x336 & ~x357 & ~x390 & ~x397 & ~x398 & ~x415 & ~x420 & ~x423 & ~x441 & ~x501 & ~x532 & ~x538 & ~x539 & ~x552 & ~x558 & ~x559 & ~x561 & ~x566 & ~x591 & ~x595 & ~x613 & ~x614 & ~x619 & ~x621 & ~x630 & ~x639 & ~x640 & ~x641 & ~x651 & ~x658 & ~x664 & ~x665 & ~x670 & ~x676 & ~x677 & ~x692 & ~x696 & ~x698 & ~x705 & ~x707 & ~x720 & ~x724 & ~x734 & ~x742 & ~x761 & ~x770 & ~x777 & ~x779;
assign c1394 =  x767 &  x771 &  x772 &  x773 & ~x192 & ~x769;
assign c1396 = ~x175 & ~x328 & ~x494 & ~x568 & ~x741;
assign c1398 =  x68 &  x125 &  x236 &  x263 &  x348 &  x376 & ~x9 & ~x20 & ~x47 & ~x49 & ~x55 & ~x57 & ~x61 & ~x77 & ~x83 & ~x89 & ~x92 & ~x105 & ~x107 & ~x108 & ~x109 & ~x110 & ~x111 & ~x115 & ~x116 & ~x138 & ~x142 & ~x147 & ~x148 & ~x163 & ~x169 & ~x191 & ~x196 & ~x198 & ~x200 & ~x220 & ~x222 & ~x223 & ~x225 & ~x227 & ~x230 & ~x259 & ~x273 & ~x279 & ~x281 & ~x282 & ~x283 & ~x284 & ~x300 & ~x309 & ~x312 & ~x313 & ~x316 & ~x317 & ~x330 & ~x338 & ~x340 & ~x367 & ~x383 & ~x384 & ~x389 & ~x392 & ~x393 & ~x396 & ~x400 & ~x415 & ~x416 & ~x425 & ~x428 & ~x441 & ~x447 & ~x456 & ~x468 & ~x474 & ~x475 & ~x476 & ~x483 & ~x495 & ~x507 & ~x513 & ~x524 & ~x525 & ~x527 & ~x532 & ~x534 & ~x537 & ~x556 & ~x566 & ~x567 & ~x569 & ~x581 & ~x584 & ~x586 & ~x592 & ~x614 & ~x616 & ~x622 & ~x636 & ~x667 & ~x669 & ~x673 & ~x677 & ~x679 & ~x703 & ~x719 & ~x729 & ~x731 & ~x733 & ~x759 & ~x760 & ~x764 & ~x775 & ~x776;
assign c1400 =  x605 & ~x78 & ~x80 & ~x87 & ~x109 & ~x305 & ~x307 & ~x331 & ~x395 & ~x427 & ~x441 & ~x563 & ~x630 & ~x658 & ~x676 & ~x686 & ~x714;
assign c1402 =  x0;
assign c1404 =  x46 &  x74 &  x102 &  x156 &  x180 &  x298 &  x327 &  x344 &  x372 &  x485 &  x569 &  x578 &  x681 & ~x21 & ~x22 & ~x28 & ~x49 & ~x51 & ~x162 & ~x201 & ~x282 & ~x285 & ~x303 & ~x330 & ~x341 & ~x391 & ~x396 & ~x478 & ~x583 & ~x705 & ~x763;
assign c1406 =  x643;
assign c1408 =  x408 & ~x573 & ~x574 & ~x602;
assign c1410 =  x683 & ~x129 & ~x172 & ~x228 & ~x275 & ~x286 & ~x315 & ~x363 & ~x397 & ~x442 & ~x469 & ~x552 & ~x590 & ~x615 & ~x639 & ~x750 & ~x781;
assign c1412 = ~x5 & ~x21 & ~x22 & ~x28 & ~x32 & ~x52 & ~x77 & ~x83 & ~x87 & ~x134 & ~x138 & ~x143 & ~x160 & ~x172 & ~x194 & ~x221 & ~x229 & ~x230 & ~x231 & ~x232 & ~x259 & ~x275 & ~x288 & ~x305 & ~x306 & ~x311 & ~x312 & ~x328 & ~x334 & ~x362 & ~x368 & ~x369 & ~x372 & ~x383 & ~x390 & ~x392 & ~x399 & ~x401 & ~x413 & ~x414 & ~x425 & ~x428 & ~x439 & ~x440 & ~x441 & ~x451 & ~x452 & ~x456 & ~x457 & ~x467 & ~x473 & ~x484 & ~x501 & ~x512 & ~x523 & ~x524 & ~x525 & ~x532 & ~x533 & ~x534 & ~x538 & ~x541 & ~x552 & ~x562 & ~x569 & ~x581 & ~x582 & ~x586 & ~x587 & ~x588 & ~x594 & ~x595 & ~x607 & ~x612 & ~x616 & ~x635 & ~x640 & ~x642 & ~x652 & ~x663 & ~x664 & ~x669 & ~x679 & ~x690 & ~x705 & ~x721 & ~x725 & ~x765 & ~x770 & ~x778;
assign c1414 =  x407 &  x435 &  x491 & ~x0 & ~x2 & ~x3 & ~x4 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x34 & ~x36 & ~x49 & ~x51 & ~x54 & ~x55 & ~x57 & ~x58 & ~x62 & ~x63 & ~x76 & ~x78 & ~x79 & ~x83 & ~x84 & ~x88 & ~x89 & ~x90 & ~x106 & ~x107 & ~x111 & ~x142 & ~x143 & ~x144 & ~x145 & ~x160 & ~x162 & ~x163 & ~x164 & ~x166 & ~x169 & ~x172 & ~x175 & ~x176 & ~x189 & ~x190 & ~x193 & ~x195 & ~x199 & ~x200 & ~x201 & ~x202 & ~x219 & ~x220 & ~x223 & ~x224 & ~x231 & ~x244 & ~x245 & ~x249 & ~x251 & ~x253 & ~x254 & ~x260 & ~x272 & ~x276 & ~x278 & ~x280 & ~x283 & ~x286 & ~x299 & ~x306 & ~x307 & ~x308 & ~x310 & ~x312 & ~x313 & ~x315 & ~x328 & ~x333 & ~x335 & ~x337 & ~x339 & ~x356 & ~x357 & ~x359 & ~x360 & ~x362 & ~x366 & ~x367 & ~x369 & ~x382 & ~x383 & ~x386 & ~x388 & ~x390 & ~x392 & ~x399 & ~x400 & ~x401 & ~x412 & ~x418 & ~x420 & ~x422 & ~x425 & ~x427 & ~x441 & ~x444 & ~x448 & ~x450 & ~x455 & ~x457 & ~x466 & ~x468 & ~x472 & ~x474 & ~x478 & ~x482 & ~x485 & ~x494 & ~x497 & ~x503 & ~x504 & ~x506 & ~x508 & ~x512 & ~x528 & ~x531 & ~x534 & ~x536 & ~x551 & ~x552 & ~x553 & ~x554 & ~x556 & ~x559 & ~x564 & ~x578 & ~x580 & ~x582 & ~x583 & ~x586 & ~x587 & ~x588 & ~x589 & ~x590 & ~x591 & ~x607 & ~x608 & ~x609 & ~x610 & ~x611 & ~x613 & ~x614 & ~x617 & ~x620 & ~x636 & ~x637 & ~x640 & ~x648 & ~x650 & ~x651 & ~x665 & ~x667 & ~x668 & ~x670 & ~x673 & ~x674 & ~x675 & ~x691 & ~x693 & ~x698 & ~x701 & ~x703 & ~x704 & ~x706 & ~x719 & ~x720 & ~x721 & ~x723 & ~x726 & ~x727 & ~x728 & ~x730 & ~x733 & ~x734 & ~x735 & ~x736 & ~x749 & ~x751 & ~x753 & ~x755 & ~x758 & ~x759 & ~x760 & ~x761 & ~x762 & ~x763 & ~x774 & ~x778 & ~x780 & ~x783;
assign c1416 =  x40 &  x98 &  x127 &  x185 &  x209 &  x214 &  x242 &  x264 &  x381 & ~x2 & ~x26 & ~x27 & ~x57 & ~x90 & ~x91 & ~x105 & ~x108 & ~x110 & ~x137 & ~x192 & ~x220 & ~x231 & ~x250 & ~x305 & ~x311 & ~x336 & ~x387 & ~x415 & ~x419 & ~x424 & ~x450 & ~x455 & ~x469 & ~x505 & ~x536 & ~x537 & ~x558 & ~x561 & ~x586 & ~x588 & ~x623 & ~x643 & ~x650 & ~x672 & ~x673 & ~x680 & ~x699 & ~x704 & ~x725 & ~x732 & ~x749 & ~x752 & ~x760;
assign c1418 =  x294 &  x662 &  x718 &  x736 &  x747 &  x748 & ~x742;
assign c1420 =  x238 &  x264 &  x433 &  x435 &  x686 & ~x6 & ~x8 & ~x23 & ~x24 & ~x25 & ~x30 & ~x31 & ~x47 & ~x51 & ~x61 & ~x76 & ~x77 & ~x81 & ~x83 & ~x105 & ~x109 & ~x110 & ~x117 & ~x120 & ~x132 & ~x133 & ~x140 & ~x159 & ~x163 & ~x164 & ~x165 & ~x167 & ~x170 & ~x174 & ~x193 & ~x197 & ~x204 & ~x216 & ~x220 & ~x226 & ~x231 & ~x246 & ~x253 & ~x254 & ~x255 & ~x256 & ~x260 & ~x271 & ~x273 & ~x279 & ~x281 & ~x282 & ~x288 & ~x299 & ~x300 & ~x302 & ~x306 & ~x308 & ~x314 & ~x316 & ~x327 & ~x329 & ~x330 & ~x331 & ~x332 & ~x333 & ~x342 & ~x354 & ~x355 & ~x358 & ~x359 & ~x370 & ~x383 & ~x384 & ~x387 & ~x394 & ~x400 & ~x410 & ~x412 & ~x413 & ~x414 & ~x417 & ~x422 & ~x424 & ~x425 & ~x446 & ~x450 & ~x453 & ~x454 & ~x455 & ~x469 & ~x474 & ~x475 & ~x480 & ~x484 & ~x494 & ~x495 & ~x498 & ~x499 & ~x500 & ~x505 & ~x523 & ~x524 & ~x525 & ~x528 & ~x529 & ~x531 & ~x535 & ~x539 & ~x552 & ~x555 & ~x562 & ~x565 & ~x566 & ~x580 & ~x591 & ~x592 & ~x607 & ~x609 & ~x610 & ~x614 & ~x616 & ~x621 & ~x624 & ~x636 & ~x640 & ~x641 & ~x648 & ~x651 & ~x652 & ~x671 & ~x674 & ~x677 & ~x678 & ~x680 & ~x692 & ~x697 & ~x698 & ~x701 & ~x702 & ~x703 & ~x704 & ~x705 & ~x708 & ~x719 & ~x720 & ~x721 & ~x724 & ~x749 & ~x753 & ~x756 & ~x760 & ~x761 & ~x764 & ~x765 & ~x778 & ~x780 & ~x782;
assign c1422 =  x70 &  x98 &  x123 &  x151 &  x154 &  x155 &  x180 &  x182 &  x183 &  x184 &  x206 &  x210 &  x211 &  x237 &  x238 &  x239 &  x263 &  x269 &  x271 &  x290 &  x293 &  x297 &  x320 &  x325 &  x347 &  x353 &  x375 &  x382 &  x430 &  x431 &  x437 &  x459 &  x465 &  x487 &  x493 &  x515 &  x521 &  x544 &  x549 &  x605 &  x661 &  x684 &  x717 & ~x1 & ~x25 & ~x26 & ~x54 & ~x60 & ~x78 & ~x84 & ~x86 & ~x87 & ~x108 & ~x109 & ~x110 & ~x111 & ~x113 & ~x116 & ~x136 & ~x139 & ~x143 & ~x169 & ~x170 & ~x174 & ~x193 & ~x201 & ~x222 & ~x224 & ~x246 & ~x250 & ~x253 & ~x275 & ~x277 & ~x281 & ~x282 & ~x303 & ~x304 & ~x306 & ~x307 & ~x311 & ~x314 & ~x334 & ~x336 & ~x339 & ~x341 & ~x360 & ~x387 & ~x390 & ~x395 & ~x415 & ~x418 & ~x446 & ~x449 & ~x479 & ~x504 & ~x506 & ~x528 & ~x529 & ~x534 & ~x556 & ~x585 & ~x588 & ~x589 & ~x590 & ~x618 & ~x644 & ~x646 & ~x648 & ~x669 & ~x670 & ~x671 & ~x673 & ~x675 & ~x676 & ~x703 & ~x725 & ~x726 & ~x729 & ~x731 & ~x753 & ~x759 & ~x761 & ~x777 & ~x778 & ~x779 & ~x782;
assign c1424 =  x97 &  x345 &  x375 &  x485 &  x598 & ~x2 & ~x31 & ~x50 & ~x60 & ~x77 & ~x90 & ~x107 & ~x111 & ~x135 & ~x137 & ~x139 & ~x145 & ~x189 & ~x217 & ~x227 & ~x250 & ~x257 & ~x258 & ~x273 & ~x274 & ~x303 & ~x330 & ~x336 & ~x356 & ~x357 & ~x390 & ~x392 & ~x395 & ~x423 & ~x424 & ~x426 & ~x427 & ~x441 & ~x455 & ~x469 & ~x475 & ~x483 & ~x502 & ~x509 & ~x552 & ~x553 & ~x562 & ~x645 & ~x667 & ~x692 & ~x696 & ~x701 & ~x706 & ~x720 & ~x722 & ~x733 & ~x753 & ~x761 & ~x779;
assign c1426 =  x73 &  x100 &  x234 &  x297 &  x325 &  x348 &  x354 &  x375 &  x376 &  x438 &  x466 & ~x7 & ~x91 & ~x307 & ~x329 & ~x364 & ~x368 & ~x387 & ~x415 & ~x441 & ~x455 & ~x539 & ~x553 & ~x565 & ~x586 & ~x610 & ~x618 & ~x619 & ~x620 & ~x651 & ~x666 & ~x695 & ~x706 & ~x725 & ~x776;
assign c1428 =  x646;
assign c1430 =  x39 & ~x202 & ~x276 & ~x286 & ~x329 & ~x406 & ~x475 & ~x645 & ~x721 & ~x725;
assign c1432 =  x22;
assign c1434 =  x44 &  x238 &  x267 &  x319 &  x431 &  x520 &  x631 &  x689 &  x740 &  x745 & ~x15 & ~x19 & ~x64 & ~x80 & ~x82 & ~x109 & ~x114 & ~x116 & ~x134 & ~x135 & ~x168 & ~x170 & ~x173 & ~x225 & ~x252 & ~x278 & ~x305 & ~x306 & ~x334 & ~x358 & ~x367 & ~x416 & ~x446 & ~x449 & ~x497 & ~x526 & ~x582 & ~x589 & ~x592 & ~x609 & ~x648 & ~x675 & ~x703 & ~x722 & ~x725 & ~x726 & ~x734 & ~x752 & ~x755 & ~x762 & ~x777 & ~x779;
assign c1436 =  x13 &  x17 &  x18 &  x101 & ~x5 & ~x27 & ~x85 & ~x107 & ~x108 & ~x115 & ~x138 & ~x333 & ~x336 & ~x446 & ~x474 & ~x532 & ~x647 & ~x670 & ~x671 & ~x695 & ~x730 & ~x751;
assign c1438 =  x263 & ~x20 & ~x47 & ~x60 & ~x87 & ~x110 & ~x140 & ~x188 & ~x327 & ~x334 & ~x438 & ~x466 & ~x468 & ~x469 & ~x531 & ~x536 & ~x606 & ~x618 & ~x635 & ~x698 & ~x702 & ~x746 & ~x747;
assign c1440 =  x178 &  x234 &  x237 &  x262 &  x264 &  x266 &  x267 &  x289 &  x292 &  x294 &  x324 &  x345 &  x347 &  x375 &  x401 &  x402 &  x432 &  x460 &  x464 &  x485 &  x513 &  x515 &  x547 &  x570 &  x577 &  x711 &  x771 & ~x1 & ~x5 & ~x7 & ~x22 & ~x28 & ~x29 & ~x31 & ~x35 & ~x56 & ~x78 & ~x85 & ~x105 & ~x106 & ~x110 & ~x116 & ~x133 & ~x137 & ~x138 & ~x141 & ~x161 & ~x162 & ~x167 & ~x168 & ~x190 & ~x199 & ~x201 & ~x219 & ~x220 & ~x248 & ~x275 & ~x278 & ~x283 & ~x302 & ~x303 & ~x329 & ~x339 & ~x359 & ~x361 & ~x365 & ~x388 & ~x392 & ~x423 & ~x424 & ~x446 & ~x472 & ~x478 & ~x482 & ~x498 & ~x503 & ~x506 & ~x509 & ~x528 & ~x534 & ~x535 & ~x554 & ~x559 & ~x561 & ~x583 & ~x585 & ~x587 & ~x611 & ~x619 & ~x643 & ~x649 & ~x667 & ~x668 & ~x677 & ~x702 & ~x705 & ~x725 & ~x726 & ~x730 & ~x731 & ~x733 & ~x752 & ~x760 & ~x780 & ~x781;
assign c1442 =  x42 &  x45 &  x72 &  x215 &  x261 &  x440 &  x523 &  x708 & ~x53 & ~x58 & ~x87 & ~x137 & ~x198 & ~x199 & ~x221 & ~x306 & ~x334 & ~x338 & ~x670 & ~x781;
assign c1444 =  x20 & ~x191 & ~x712 & ~x740;
assign c1446 = ~x127 & ~x235 & ~x272 & ~x288 & ~x302 & ~x328 & ~x329 & ~x341 & ~x399 & ~x454 & ~x467 & ~x495 & ~x511 & ~x512;
assign c1448 =  x213 &  x241 &  x269 &  x321 &  x325 &  x377 &  x381 &  x604 &  x629 &  x656 & ~x0 & ~x3 & ~x28 & ~x48 & ~x55 & ~x62 & ~x64 & ~x77 & ~x81 & ~x85 & ~x107 & ~x109 & ~x111 & ~x112 & ~x136 & ~x144 & ~x162 & ~x163 & ~x170 & ~x174 & ~x195 & ~x196 & ~x203 & ~x217 & ~x219 & ~x227 & ~x228 & ~x231 & ~x246 & ~x248 & ~x249 & ~x256 & ~x274 & ~x280 & ~x284 & ~x285 & ~x303 & ~x329 & ~x334 & ~x339 & ~x342 & ~x360 & ~x361 & ~x363 & ~x370 & ~x386 & ~x387 & ~x398 & ~x415 & ~x417 & ~x419 & ~x443 & ~x445 & ~x449 & ~x468 & ~x483 & ~x496 & ~x498 & ~x504 & ~x508 & ~x526 & ~x530 & ~x531 & ~x554 & ~x558 & ~x559 & ~x584 & ~x587 & ~x590 & ~x591 & ~x609 & ~x624 & ~x639 & ~x640 & ~x642 & ~x644 & ~x648 & ~x652 & ~x664 & ~x667 & ~x669 & ~x677 & ~x681 & ~x692 & ~x694 & ~x700 & ~x705 & ~x708 & ~x709 & ~x723 & ~x731 & ~x733 & ~x757 & ~x759;
assign c1450 = ~x15 & ~x19 & ~x33 & ~x54 & ~x56 & ~x90 & ~x91 & ~x105 & ~x111 & ~x115 & ~x118 & ~x145 & ~x146 & ~x160 & ~x171 & ~x187 & ~x193 & ~x194 & ~x200 & ~x201 & ~x202 & ~x243 & ~x254 & ~x255 & ~x271 & ~x299 & ~x304 & ~x305 & ~x306 & ~x308 & ~x333 & ~x362 & ~x370 & ~x371 & ~x382 & ~x391 & ~x398 & ~x413 & ~x426 & ~x428 & ~x439 & ~x440 & ~x455 & ~x466 & ~x472 & ~x475 & ~x480 & ~x483 & ~x494 & ~x495 & ~x496 & ~x498 & ~x505 & ~x511 & ~x530 & ~x558 & ~x579 & ~x586 & ~x590 & ~x591 & ~x607 & ~x611 & ~x613 & ~x621 & ~x645 & ~x648 & ~x650 & ~x662 & ~x673 & ~x696 & ~x707 & ~x710 & ~x718 & ~x719 & ~x736 & ~x751 & ~x761 & ~x762 & ~x764 & ~x765 & ~x774;
assign c1452 =  x663 & ~x602 & ~x714 & ~x742;
assign c1454 =  x19 &  x188 & ~x62 & ~x310;
assign c1456 =  x72 &  x100 &  x577 &  x683 &  x711 &  x712 &  x772 & ~x77 & ~x118 & ~x119 & ~x163 & ~x203 & ~x282 & ~x338 & ~x415 & ~x426 & ~x581 & ~x664 & ~x695 & ~x720;
assign c1458 =  x209 & ~x517 & ~x574 & ~x601 & ~x630 & ~x713;
assign c1460 =  x44 &  x149 &  x177 &  x318 &  x346 &  x768 & ~x21 & ~x27 & ~x36 & ~x79 & ~x87 & ~x89 & ~x119 & ~x169 & ~x170 & ~x172 & ~x195 & ~x222 & ~x370 & ~x415 & ~x418 & ~x474 & ~x504 & ~x533 & ~x535 & ~x583 & ~x669 & ~x678 & ~x697 & ~x699 & ~x726 & ~x754 & ~x764 & ~x776 & ~x781;
assign c1462 =  x209 &  x316 & ~x657;
assign c1464 =  x90;
assign c1466 =  x90 &  x368;
assign c1468 =  x31 & ~x296;
assign c1470 =  x42 &  x43 &  x177 &  x205 &  x233 &  x317 &  x322 &  x401 &  x541 &  x570 &  x626 &  x682 &  x710 & ~x1 & ~x22 & ~x23 & ~x26 & ~x27 & ~x28 & ~x30 & ~x36 & ~x53 & ~x61 & ~x80 & ~x89 & ~x106 & ~x111 & ~x112 & ~x113 & ~x117 & ~x141 & ~x169 & ~x170 & ~x174 & ~x192 & ~x195 & ~x196 & ~x200 & ~x219 & ~x221 & ~x223 & ~x247 & ~x253 & ~x274 & ~x301 & ~x304 & ~x305 & ~x311 & ~x313 & ~x331 & ~x332 & ~x333 & ~x334 & ~x341 & ~x342 & ~x366 & ~x367 & ~x368 & ~x370 & ~x389 & ~x395 & ~x398 & ~x415 & ~x416 & ~x424 & ~x426 & ~x441 & ~x443 & ~x444 & ~x445 & ~x451 & ~x453 & ~x472 & ~x482 & ~x483 & ~x502 & ~x534 & ~x553 & ~x564 & ~x586 & ~x588 & ~x593 & ~x594 & ~x612 & ~x613 & ~x615 & ~x617 & ~x641 & ~x642 & ~x669 & ~x695 & ~x725 & ~x728 & ~x734 & ~x752 & ~x755 & ~x761 & ~x762 & ~x764 & ~x776 & ~x782;
assign c1472 =  x11 &  x14 &  x39 &  x41 &  x67 &  x71 &  x72 &  x129 &  x182 &  x236 &  x269 & ~x34 & ~x53 & ~x58 & ~x60 & ~x64 & ~x79 & ~x104 & ~x106 & ~x135 & ~x140 & ~x143 & ~x146 & ~x172 & ~x188 & ~x200 & ~x218 & ~x222 & ~x283 & ~x331 & ~x384 & ~x470 & ~x478 & ~x509 & ~x525 & ~x529 & ~x536 & ~x557 & ~x609 & ~x611 & ~x620 & ~x668 & ~x673 & ~x705 & ~x724 & ~x751;
assign c1474 =  x525 &  x607 &  x608 &  x622;
assign c1476 = ~x71 & ~x382 & ~x423 & ~x439 & ~x466 & ~x467 & ~x624;
assign c1478 =  x74 &  x238 &  x427 &  x519 &  x523 &  x575 &  x624 &  x635 &  x682 &  x688 &  x709 & ~x90 & ~x173 & ~x257 & ~x471 & ~x534;
assign c1480 =  x67 &  x96 &  x182 &  x213 &  x236 &  x270 &  x289 &  x317 &  x326 &  x401 &  x437 &  x494 &  x661 &  x710 &  x739 &  x772 & ~x7 & ~x52 & ~x111 & ~x170 & ~x218 & ~x251 & ~x282 & ~x370 & ~x386 & ~x394 & ~x413 & ~x469 & ~x558 & ~x564 & ~x588 & ~x613 & ~x673 & ~x700;
assign c1482 =  x95 &  x262 &  x326 &  x374 &  x772 & ~x3 & ~x4 & ~x499 & ~x581 & ~x639 & ~x754;
assign c1484 = ~x27 & ~x50 & ~x54 & ~x56 & ~x85 & ~x135 & ~x140 & ~x162 & ~x164 & ~x170 & ~x171 & ~x195 & ~x220 & ~x260 & ~x275 & ~x277 & ~x278 & ~x281 & ~x329 & ~x373 & ~x374 & ~x439 & ~x454 & ~x527 & ~x558 & ~x595 & ~x623 & ~x652 & ~x673 & ~x680 & ~x733 & ~x739 & ~x766 & ~x767;
assign c1486 =  x97 & ~x453 & ~x459 & ~x651;
assign c1488 =  x41 & ~x77 & ~x80 & ~x145 & ~x163 & ~x245 & ~x273 & ~x282 & ~x300 & ~x329 & ~x383 & ~x444 & ~x469 & ~x489 & ~x497 & ~x554 & ~x643 & ~x647;
assign c1490 =  x8 &  x775;
assign c1492 =  x103 &  x596 &  x734;
assign c1494 =  x46 &  x47 &  x103 & ~x24 & ~x143 & ~x630 & ~x686 & ~x714;
assign c1496 =  x522 & ~x55 & ~x546 & ~x603 & ~x631;
assign c1498 =  x99 &  x153 &  x238 &  x269 &  x293 &  x344 &  x345 &  x428 &  x623 &  x635 & ~x114 & ~x279 & ~x391 & ~x757 & ~x759 & ~x781;
assign c11 = ~x66 & ~x93 & ~x98 & ~x209;
assign c13 =  x185 &  x489 &  x490 &  x514 & ~x79 & ~x339 & ~x766 & ~x768;
assign c15 =  x41 &  x407 &  x493 &  x543 &  x571 & ~x1 & ~x10 & ~x47 & ~x308 & ~x419 & ~x450 & ~x584 & ~x766 & ~x767 & ~x779;
assign c17 = ~x131 & ~x140 & ~x239 & ~x322 & ~x368 & ~x532;
assign c19 =  x350 &  x379 &  x404 &  x545 &  x600 &  x768 &  x769 &  x770 & ~x25 & ~x52 & ~x274 & ~x368 & ~x419 & ~x533 & ~x554 & ~x556 & ~x587 & ~x695 & ~x700;
assign c111 =  x436 &  x490 &  x630 &  x655 &  x740 &  x741 &  x769 &  x770 & ~x5 & ~x7 & ~x164 & ~x194 & ~x338 & ~x507 & ~x526 & ~x527 & ~x588 & ~x783;
assign c113 =  x546 &  x571 &  x689 &  x714 &  x770 & ~x197 & ~x511;
assign c115 = ~x75 & ~x102 & ~x122 & ~x124 & ~x763;
assign c117 =  x334;
assign c119 =  x97 &  x465 &  x519 &  x602 &  x627 & ~x10 & ~x22 & ~x79 & ~x114 & ~x143 & ~x175 & ~x220 & ~x223 & ~x531 & ~x730 & ~x731 & ~x754 & ~x766 & ~x783;
assign c121 =  x426 & ~x20 & ~x87 & ~x88 & ~x135 & ~x756;
assign c123 = ~x487 & ~x488 & ~x660 & ~x777;
assign c125 =  x686 &  x739 & ~x2 & ~x24 & ~x60 & ~x87 & ~x108 & ~x137 & ~x143 & ~x201 & ~x218 & ~x222 & ~x227 & ~x234 & ~x242 & ~x262 & ~x305 & ~x312 & ~x334 & ~x342 & ~x361 & ~x367 & ~x397 & ~x423 & ~x474 & ~x502 & ~x506 & ~x555 & ~x589 & ~x613 & ~x699 & ~x700 & ~x704 & ~x723;
assign c127 = ~x13 & ~x542 & ~x569 & ~x600 & ~x622;
assign c129 = ~x23 & ~x131 & ~x148 & ~x194 & ~x573 & ~x587 & ~x599 & ~x601 & ~x603 & ~x633 & ~x778;
assign c131 =  x63 &  x769;
assign c133 =  x472;
assign c135 =  x511 & ~x638 & ~x764;
assign c137 =  x487 &  x599 &  x602 &  x658 &  x714 & ~x26 & ~x190 & ~x234 & ~x645;
assign c139 =  x411 & ~x596 & ~x691;
assign c141 =  x344;
assign c143 =  x157 &  x461 &  x630 &  x659 &  x712 & ~x30 & ~x142 & ~x165 & ~x168 & ~x305 & ~x339 & ~x360 & ~x417 & ~x511 & ~x667 & ~x673 & ~x757 & ~x768;
assign c145 = ~x2 & ~x5 & ~x32 & ~x84 & ~x133 & ~x136 & ~x137 & ~x193 & ~x196 & ~x210 & ~x219 & ~x307 & ~x364 & ~x529 & ~x559;
assign c147 = ~x5 & ~x24 & ~x113 & ~x172 & ~x367 & ~x389 & ~x423 & ~x533 & ~x616 & ~x622 & ~x642 & ~x657 & ~x660 & ~x687 & ~x721 & ~x734 & ~x763 & ~x777;
assign c149 = ~x1 & ~x7 & ~x14 & ~x53 & ~x139 & ~x146 & ~x169 & ~x202 & ~x210 & ~x222 & ~x257 & ~x285 & ~x587 & ~x731;
assign c151 =  x356 & ~x26 & ~x49 & ~x59 & ~x104 & ~x110 & ~x113 & ~x776;
assign c153 =  x96 &  x97 &  x238 &  x461 &  x574 &  x658 &  x659 & ~x4 & ~x32 & ~x90 & ~x115 & ~x171 & ~x191 & ~x205 & ~x255 & ~x271 & ~x342 & ~x358 & ~x373 & ~x400 & ~x420 & ~x446 & ~x482 & ~x503 & ~x567 & ~x643 & ~x647 & ~x672 & ~x673 & ~x675 & ~x728;
assign c155 =  x135;
assign c157 =  x193;
assign c159 =  x158 &  x378 &  x468 &  x546 &  x628 &  x656 &  x740 & ~x700;
assign c161 =  x485 & ~x18 & ~x113 & ~x345 & ~x474 & ~x512 & ~x775;
assign c163 =  x43 &  x375 &  x376 &  x403 &  x405 &  x485 &  x487 & ~x32 & ~x59 & ~x108 & ~x191 & ~x193 & ~x220 & ~x275 & ~x304 & ~x390 & ~x449 & ~x500 & ~x533 & ~x535 & ~x590 & ~x619 & ~x643 & ~x729 & ~x731 & ~x766 & ~x775;
assign c165 = ~x6 & ~x19 & ~x58 & ~x80 & ~x211 & ~x266;
assign c167 = ~x408;
assign c169 =  x669;
assign c171 = ~x34 & ~x111 & ~x121 & ~x169 & ~x238 & ~x266 & ~x728;
assign c173 =  x258 & ~x642;
assign c175 =  x62;
assign c177 =  x332;
assign c179 =  x466 & ~x1 & ~x5 & ~x39 & ~x56 & ~x65 & ~x75 & ~x86 & ~x114 & ~x230 & ~x251 & ~x256 & ~x364 & ~x394 & ~x589 & ~x616 & ~x760;
assign c181 =  x769 & ~x10 & ~x24 & ~x184;
assign c183 =  x403 &  x546 &  x574 &  x686 &  x689 &  x714 &  x770 & ~x19 & ~x138 & ~x279 & ~x567 & ~x666;
assign c185 =  x434 &  x517 &  x547 &  x599 &  x689 &  x712 &  x769 &  x770 &  x771 & ~x8 & ~x20 & ~x24 & ~x84 & ~x164 & ~x223 & ~x224 & ~x225 & ~x273 & ~x281 & ~x302 & ~x451 & ~x476 & ~x498 & ~x587 & ~x617 & ~x646 & ~x751;
assign c187 =  x455 & ~x152;
assign c189 =  x677 & ~x393;
assign c191 =  x39 &  x71 &  x181 &  x184 & ~x4 & ~x7 & ~x20 & ~x24 & ~x58 & ~x59 & ~x81 & ~x84 & ~x248 & ~x279 & ~x280 & ~x445 & ~x477 & ~x479 & ~x563 & ~x730 & ~x774;
assign c193 =  x244 & ~x2 & ~x765;
assign c195 =  x380 & ~x225 & ~x238 & ~x758;
assign c197 =  x553 & ~x20 & ~x360;
assign c199 =  x518 & ~x1 & ~x56 & ~x139 & ~x164 & ~x225 & ~x255 & ~x281 & ~x362 & ~x391 & ~x394 & ~x448 & ~x616 & ~x670 & ~x700 & ~x728 & ~x729 & ~x748 & ~x757 & ~x770 & ~x771 & ~x773;
assign c1101 = ~x41 & ~x146 & ~x217 & ~x684;
assign c1103 = ~x14 & ~x599 & ~x600 & ~x605 & ~x663;
assign c1105 = ~x13 & ~x516 & ~x741 & ~x776;
assign c1107 =  x284;
assign c1109 =  x69 &  x70 &  x181 &  x208 &  x464 &  x490 & ~x14 & ~x52 & ~x55 & ~x132 & ~x148 & ~x163 & ~x195 & ~x243 & ~x250 & ~x280 & ~x310 & ~x369 & ~x480 & ~x532 & ~x536 & ~x586 & ~x591 & ~x640 & ~x650;
assign c1111 =  x65 &  x245;
assign c1113 =  x43 &  x44 & ~x6 & ~x162 & ~x336 & ~x351 & ~x443 & ~x668 & ~x674 & ~x760;
assign c1115 =  x272 & ~x635;
assign c1117 =  x405 &  x634 &  x686 &  x711 &  x745 & ~x115 & ~x137 & ~x252 & ~x283 & ~x335 & ~x670 & ~x707;
assign c1119 =  x593 & ~x709;
assign c1121 =  x372 &  x658 &  x745 & ~x12;
assign c1123 =  x127 &  x157 &  x597 & ~x15 & ~x307 & ~x344 & ~x527;
assign c1125 = ~x487 & ~x576;
assign c1127 = ~x401 & ~x460 & ~x632 & ~x735;
assign c1129 =  x43 & ~x23 & ~x102 & ~x107 & ~x189 & ~x224 & ~x351 & ~x363 & ~x666;
assign c1131 =  x72 &  x118 & ~x21 & ~x86 & ~x615;
assign c1133 =  x370;
assign c1135 =  x715 & ~x56 & ~x195 & ~x206 & ~x234 & ~x345 & ~x454 & ~x497 & ~x617 & ~x750;
assign c1137 = ~x604 & ~x628 & ~x630 & ~x661 & ~x679 & ~x687 & ~x710 & ~x735;
assign c1139 =  x124 &  x267 &  x434 &  x628 &  x657 &  x710 &  x714 &  x742 &  x746 & ~x30 & ~x54 & ~x247 & ~x280 & ~x337 & ~x383 & ~x393 & ~x399 & ~x444 & ~x456 & ~x535 & ~x564 & ~x613 & ~x617 & ~x642 & ~x730 & ~x732 & ~x751;
assign c1141 = ~x6 & ~x13 & ~x19 & ~x432 & ~x748 & ~x777;
assign c1143 =  x208 &  x739 &  x741 & ~x1 & ~x10 & ~x53 & ~x108 & ~x119 & ~x196 & ~x269 & ~x333 & ~x366 & ~x423 & ~x449;
assign c1145 =  x41 &  x433 &  x465 &  x572 & ~x55 & ~x89 & ~x114 & ~x270 & ~x338 & ~x724;
assign c1147 = ~x11 & ~x167 & ~x254 & ~x266 & ~x278 & ~x282 & ~x304 & ~x317 & ~x640 & ~x752;
assign c1149 =  x711 &  x737 &  x769 & ~x81 & ~x84 & ~x251 & ~x391 & ~x395 & ~x445 & ~x450 & ~x617 & ~x698;
assign c1151 = ~x4 & ~x6 & ~x432;
assign c1153 =  x69 &  x433 &  x434 &  x491 &  x516 &  x545 &  x570 &  x571 &  x628 &  x629 &  x683 & ~x24 & ~x25 & ~x56 & ~x168 & ~x194 & ~x588 & ~x755 & ~x772;
assign c1155 =  x95 &  x405 &  x433 &  x571 &  x574 &  x629 & ~x22 & ~x60 & ~x83 & ~x111 & ~x197 & ~x277 & ~x281 & ~x305 & ~x476 & ~x502 & ~x505 & ~x591 & ~x757 & ~x765 & ~x768;
assign c1157 =  x43 &  x68 &  x94 &  x151 & ~x7 & ~x20 & ~x29 & ~x32 & ~x58 & ~x109 & ~x110 & ~x140 & ~x141 & ~x165 & ~x167 & ~x168 & ~x248 & ~x252 & ~x276 & ~x279 & ~x284 & ~x310 & ~x340 & ~x363 & ~x366 & ~x367 & ~x391 & ~x418 & ~x444 & ~x446 & ~x472 & ~x478 & ~x501 & ~x505 & ~x529 & ~x533 & ~x534 & ~x559 & ~x560 & ~x561 & ~x588 & ~x590 & ~x613 & ~x615 & ~x642 & ~x644 & ~x671 & ~x729 & ~x773;
assign c1159 =  x388 &  x573;
assign c1161 =  x499 & ~x49;
assign c1163 =  x127 &  x154 &  x212 &  x347 &  x348 &  x433 &  x465 &  x517 &  x518 &  x599 &  x602 &  x659 &  x685 &  x714 & ~x250 & ~x252 & ~x282 & ~x331 & ~x340 & ~x373 & ~x384 & ~x399 & ~x527 & ~x534 & ~x561 & ~x753;
assign c1165 =  x42 &  x204 & ~x775;
assign c1167 =  x303;
assign c1169 =  x129 &  x378 &  x463 &  x518 &  x570 &  x576 &  x655 &  x686 &  x711 &  x741 &  x769 &  x770 & ~x26 & ~x29 & ~x59 & ~x199 & ~x222 & ~x229 & ~x368 & ~x417 & ~x423 & ~x560 & ~x614 & ~x702;
assign c1171 =  x64 &  x658 & ~x563;
assign c1173 =  x663 &  x740 &  x770;
assign c1175 = ~x436 & ~x460 & ~x491 & ~x691;
assign c1177 =  x737 &  x740 & ~x14;
assign c1179 =  x299 & ~x4 & ~x27 & ~x45 & ~x76 & ~x86 & ~x112 & ~x114 & ~x255;
assign c1181 =  x299 &  x327 & ~x73;
assign c1183 =  x741 & ~x121 & ~x161 & ~x325 & ~x586;
assign c1185 =  x64 &  x573 & ~x225 & ~x670 & ~x758;
assign c1187 = ~x603 & ~x604 & ~x605 & ~x668 & ~x683 & ~x687 & ~x749;
assign c1189 = ~x83 & ~x169 & ~x390 & ~x442 & ~x470 & ~x481 & ~x509 & ~x572 & ~x576 & ~x592 & ~x603 & ~x711 & ~x759;
assign c1191 =  x78;
assign c1193 =  x98 &  x517 &  x599 &  x709 &  x740 & ~x8 & ~x116 & ~x167 & ~x173 & ~x246 & ~x248 & ~x356 & ~x424 & ~x502 & ~x510 & ~x530 & ~x615 & ~x671 & ~x760;
assign c1195 =  x40 &  x230 & ~x1 & ~x3 & ~x21 & ~x25 & ~x30 & ~x141 & ~x252 & ~x280 & ~x309 & ~x362 & ~x586 & ~x644 & ~x646 & ~x672 & ~x781;
assign c1197 =  x267 &  x519 &  x720 &  x740 &  x769 &  x770;
assign c1199 =  x91 &  x574;
assign c1201 =  x17 &  x713 &  x714 &  x739;
assign c1203 =  x129 &  x156 &  x157 &  x293 &  x513 & ~x4 & ~x20 & ~x23 & ~x61 & ~x78 & ~x81 & ~x82 & ~x117 & ~x163 & ~x172 & ~x199 & ~x225 & ~x251 & ~x277 & ~x279 & ~x280 & ~x282 & ~x288 & ~x310 & ~x328 & ~x339 & ~x342 & ~x367 & ~x369 & ~x390 & ~x418 & ~x423 & ~x469 & ~x525 & ~x539 & ~x613 & ~x642 & ~x666 & ~x670 & ~x753 & ~x779;
assign c1205 =  x209 &  x378 &  x436 &  x491 &  x573 &  x688 &  x745 &  x769 &  x770 & ~x8 & ~x26 & ~x117 & ~x329 & ~x358 & ~x502 & ~x565 & ~x610;
assign c1207 = ~x19 & ~x21 & ~x281 & ~x323 & ~x326 & ~x406 & ~x728 & ~x730;
assign c1209 =  x69 & ~x4 & ~x11 & ~x56 & ~x113 & ~x196 & ~x291 & ~x305 & ~x752 & ~x775 & ~x776;
assign c1211 =  x267 &  x292 &  x379 &  x403 &  x431 &  x435 &  x459 &  x462 &  x488 &  x515 &  x518 &  x519 &  x520 &  x570 &  x573 &  x575 &  x631 & ~x2 & ~x4 & ~x22 & ~x28 & ~x56 & ~x57 & ~x81 & ~x88 & ~x111 & ~x112 & ~x142 & ~x198 & ~x221 & ~x223 & ~x282 & ~x284 & ~x305 & ~x308 & ~x334 & ~x361 & ~x367 & ~x390 & ~x422 & ~x450 & ~x476 & ~x502 & ~x507 & ~x534 & ~x537 & ~x588 & ~x589 & ~x615 & ~x701 & ~x727 & ~x754 & ~x756 & ~x757 & ~x758 & ~x769 & ~x771;
assign c1213 =  x680 & ~x19;
assign c1215 =  x69 &  x573 &  x575 &  x656 &  x739 & ~x11 & ~x132 & ~x136 & ~x142 & ~x308 & ~x309 & ~x314 & ~x333 & ~x357 & ~x499 & ~x506 & ~x615 & ~x730 & ~x759;
assign c1217 =  x36 &  x517 & ~x167 & ~x223;
assign c1219 =  x74 &  x92 &  x349 & ~x620 & ~x644;
assign c1221 =  x686 &  x711 & ~x2 & ~x26 & ~x31 & ~x262;
assign c1223 =  x127 &  x238 &  x435 &  x518 &  x520 &  x745 &  x769 &  x770 & ~x277 & ~x331 & ~x582 & ~x695;
assign c1225 = ~x95 & ~x101 & ~x126 & ~x129 & ~x711;
assign c1227 =  x116;
assign c1229 =  x430 & ~x20 & ~x59 & ~x106 & ~x112 & ~x115 & ~x141 & ~x251 & ~x310 & ~x360 & ~x533 & ~x560 & ~x618 & ~x641 & ~x644 & ~x700 & ~x730 & ~x755 & ~x766 & ~x767 & ~x771 & ~x773;
assign c1231 =  x97 &  x125 &  x127 &  x154 &  x266 &  x292 &  x354 &  x376 &  x433 &  x517 &  x519 &  x549 &  x570 &  x571 &  x603 &  x605 &  x625 &  x654 &  x657 &  x686 &  x689 & ~x7 & ~x29 & ~x84 & ~x143 & ~x166 & ~x197 & ~x306 & ~x335 & ~x336 & ~x368 & ~x391 & ~x504 & ~x531 & ~x556 & ~x563 & ~x615 & ~x648 & ~x756 & ~x758;
assign c1233 =  x329 & ~x20 & ~x134;
assign c1235 =  x603 &  x711;
assign c1237 =  x501;
assign c1241 =  x272 &  x602 &  x658 &  x739 &  x741;
assign c1243 =  x231 &  x244 & ~x19;
assign c1245 =  x165;
assign c1247 =  x98 &  x517 &  x520 &  x570 &  x601 & ~x62 & ~x81 & ~x115 & ~x476 & ~x587 & ~x649 & ~x699 & ~x766 & ~x767;
assign c1249 =  x522 &  x709 &  x718 &  x747 &  x770 & ~x281;
assign c1251 =  x40 &  x41 &  x42 &  x43 & ~x7 & ~x9 & ~x22 & ~x31 & ~x52 & ~x54 & ~x56 & ~x80 & ~x83 & ~x107 & ~x195 & ~x197 & ~x223 & ~x225 & ~x249 & ~x252 & ~x279 & ~x280 & ~x282 & ~x332 & ~x336 & ~x338 & ~x388 & ~x420 & ~x423 & ~x448 & ~x450 & ~x451 & ~x579 & ~x589 & ~x616 & ~x635 & ~x652 & ~x663 & ~x681 & ~x691 & ~x702 & ~x728 & ~x730 & ~x768 & ~x775 & ~x779 & ~x782;
assign c1253 =  x64 &  x130 &  x601 & ~x169;
assign c1255 =  x706 &  x712;
assign c1257 =  x406 &  x434 &  x465 &  x548 & ~x3 & ~x9 & ~x10 & ~x20 & ~x140 & ~x222 & ~x280 & ~x357 & ~x561 & ~x588 & ~x672 & ~x677 & ~x704 & ~x767;
assign c1259 =  x63 &  x741;
assign c1261 =  x43 &  x274 & ~x397 & ~x670;
assign c1263 =  x71 &  x686 &  x739 & ~x2 & ~x250;
assign c1265 =  x742 &  x747 &  x766 &  x770 & ~x80;
assign c1267 =  x154 &  x157 &  x186 &  x376 &  x409 &  x514 &  x521 &  x542 &  x602 &  x659 &  x686 &  x690 &  x709 &  x712 &  x714 &  x716 &  x718 &  x738 &  x739 &  x741 &  x745 & ~x1 & ~x59 & ~x110 & ~x114 & ~x222 & ~x250 & ~x254 & ~x363 & ~x366 & ~x475 & ~x504 & ~x506 & ~x588 & ~x700;
assign c1269 =  x737 &  x739 &  x741 &  x742 & ~x1 & ~x4 & ~x400 & ~x428 & ~x553 & ~x612 & ~x640;
assign c1271 =  x259 &  x712;
assign c1273 =  x186 &  x597 &  x740 &  x742 & ~x14;
assign c1277 =  x70 &  x127 &  x181 &  x290 &  x433 &  x434 &  x518 &  x522 &  x657 &  x661 &  x747 & ~x0 & ~x31 & ~x55 & ~x166 & ~x198 & ~x280 & ~x332 & ~x356 & ~x389 & ~x420 & ~x530 & ~x592 & ~x645 & ~x703 & ~x722 & ~x781;
assign c1279 =  x554 &  x599;
assign c1281 =  x573 &  x712 &  x739 &  x770 & ~x2 & ~x34 & ~x49 & ~x54 & ~x84 & ~x112 & ~x140 & ~x195 & ~x223 & ~x225 & ~x253 & ~x278 & ~x279 & ~x282 & ~x299 & ~x392 & ~x418 & ~x441 & ~x480 & ~x502 & ~x534 & ~x555 & ~x558 & ~x565 & ~x588 & ~x619 & ~x644 & ~x670 & ~x671 & ~x676 & ~x698 & ~x703 & ~x704 & ~x729 & ~x753 & ~x761;
assign c1283 =  x404 &  x405 &  x435 &  x459 &  x488 &  x514 &  x543 &  x546 &  x547 &  x576 &  x601 &  x630 &  x657 & ~x3 & ~x33 & ~x58 & ~x224 & ~x255 & ~x306 & ~x338 & ~x364 & ~x446 & ~x449 & ~x771 & ~x782;
assign c1285 =  x329;
assign c1287 = ~x403 & ~x491 & ~x492 & ~x493;
assign c1289 =  x375 &  x493 &  x547 & ~x7 & ~x9 & ~x19 & ~x29 & ~x31 & ~x53 & ~x60 & ~x83 & ~x114 & ~x192 & ~x196 & ~x225 & ~x254 & ~x333 & ~x449 & ~x505 & ~x533 & ~x738 & ~x755 & ~x775;
assign c1291 =  x215 &  x322 &  x431 & ~x78 & ~x222 & ~x698 & ~x766;
assign c1293 = ~x264 & ~x345 & ~x375 & ~x719;
assign c1295 =  x737 &  x739 &  x741 &  x742 &  x743 &  x746 & ~x0 & ~x1 & ~x3 & ~x6 & ~x7 & ~x14 & ~x22 & ~x23 & ~x30 & ~x31 & ~x54 & ~x55 & ~x80 & ~x82 & ~x87 & ~x109 & ~x110 & ~x111 & ~x114 & ~x115 & ~x116 & ~x141 & ~x165 & ~x168 & ~x194 & ~x198 & ~x251 & ~x252 & ~x279 & ~x306 & ~x336 & ~x368 & ~x391 & ~x392 & ~x394 & ~x420 & ~x446 & ~x448 & ~x502 & ~x503 & ~x532 & ~x534 & ~x558 & ~x587 & ~x589 & ~x619 & ~x642 & ~x643 & ~x644 & ~x645 & ~x648 & ~x673 & ~x675 & ~x700 & ~x756 & ~x757 & ~x760 & ~x777 & ~x780 & ~x781 & ~x782;
assign c1297 = ~x15 & ~x16 & ~x121 & ~x166 & ~x669 & ~x728 & ~x763;
assign c1299 = ~x154 & ~x348;
assign c1301 =  x263 &  x514 &  x516 &  x548 &  x570 &  x573 &  x574 & ~x141 & ~x226 & ~x526 & ~x581 & ~x589 & ~x767;
assign c1303 =  x630 & ~x101 & ~x196;
assign c1305 =  x46 & ~x7 & ~x199 & ~x222 & ~x261 & ~x289 & ~x309 & ~x447 & ~x563;
assign c1307 = ~x93 & ~x95 & ~x101 & ~x136 & ~x208 & ~x758 & ~x782;
assign c1309 =  x332;
assign c1311 =  x145;
assign c1313 =  x108;
assign c1315 =  x93 & ~x709 & ~x710 & ~x768;
assign c1317 =  x276;
assign c1319 =  x243 &  x655 &  x658 & ~x17;
assign c1321 = ~x18 & ~x19 & ~x27 & ~x48 & ~x49 & ~x55 & ~x137 & ~x336 & ~x408 & ~x447 & ~x735 & ~x778;
assign c1323 =  x218 & ~x442 & ~x454 & ~x510 & ~x526 & ~x566;
assign c1325 =  x378 & ~x79 & ~x707 & ~x710 & ~x741;
assign c1327 = ~x34 & ~x116 & ~x394 & ~x654 & ~x686 & ~x691 & ~x698 & ~x740;
assign c1329 =  x37 &  x38 &  x40 &  x438 & ~x1 & ~x3 & ~x20 & ~x21 & ~x28 & ~x29 & ~x30 & ~x55 & ~x57 & ~x85 & ~x88 & ~x110 & ~x111 & ~x112 & ~x113 & ~x168 & ~x193 & ~x221 & ~x309 & ~x364 & ~x393 & ~x448 & ~x449 & ~x475 & ~x477 & ~x532 & ~x534 & ~x565 & ~x583 & ~x646 & ~x647 & ~x671 & ~x702 & ~x752 & ~x760 & ~x777;
assign c1331 =  x467 & ~x6 & ~x17 & ~x132 & ~x391 & ~x394 & ~x754;
assign c1333 =  x62 &  x573;
assign c1335 =  x37 &  x75 & ~x425;
assign c1337 =  x120 & ~x650 & ~x765;
assign c1339 =  x120 &  x408 &  x548 &  x571 &  x573 &  x574 &  x713 &  x740;
assign c1341 =  x287 &  x301 & ~x19 & ~x34 & ~x48 & ~x77;
assign c1343 =  x443;
assign c1345 =  x350 &  x459 &  x463 &  x518 &  x712 &  x739 &  x745 &  x769 &  x770 & ~x4 & ~x29 & ~x53 & ~x55 & ~x61 & ~x83 & ~x84 & ~x138 & ~x143 & ~x194 & ~x335 & ~x470 & ~x475 & ~x476 & ~x498 & ~x499 & ~x502 & ~x535 & ~x556 & ~x588 & ~x590 & ~x610 & ~x648 & ~x759;
assign c1347 =  x302;
assign c1349 =  x664 & ~x384 & ~x427;
assign c1351 =  x43 & ~x408 & ~x697;
assign c1353 =  x744 &  x769 &  x770 & ~x568 & ~x587;
assign c1355 =  x40 &  x41 &  x43 &  x486 &  x658 & ~x29 & ~x90 & ~x317 & ~x364 & ~x400 & ~x441 & ~x553 & ~x559 & ~x693;
assign c1357 = ~x24 & ~x46 & ~x109 & ~x743 & ~x748 & ~x768 & ~x772;
assign c1359 =  x69 &  x124 &  x489 & ~x83 & ~x270 & ~x317 & ~x471 & ~x527 & ~x610 & ~x674 & ~x757;
assign c1361 =  x97 &  x127 &  x153 &  x156 &  x240 &  x322 &  x465 &  x521 &  x546 &  x547 &  x685 &  x714 & ~x24 & ~x25 & ~x60 & ~x81 & ~x113 & ~x114 & ~x116 & ~x144 & ~x218 & ~x248 & ~x306 & ~x317 & ~x344 & ~x367 & ~x371 & ~x416 & ~x484 & ~x614 & ~x622 & ~x673 & ~x750 & ~x752 & ~x779;
assign c1363 =  x100 &  x296 & ~x0 & ~x39 & ~x44 & ~x695 & ~x765 & ~x766;
assign c1365 =  x569 & ~x10 & ~x48 & ~x199 & ~x767;
assign c1367 =  x483 &  x515 &  x630 & ~x0 & ~x18 & ~x78;
assign c1369 =  x611 & ~x57;
assign c1371 =  x739 &  x742 & ~x110 & ~x139 & ~x169 & ~x296 & ~x335 & ~x532 & ~x668 & ~x724 & ~x755;
assign c1373 =  x40 &  x41 & ~x6 & ~x7 & ~x9 & ~x19 & ~x22 & ~x23 & ~x26 & ~x29 & ~x32 & ~x33 & ~x48 & ~x53 & ~x54 & ~x57 & ~x58 & ~x59 & ~x60 & ~x77 & ~x85 & ~x86 & ~x87 & ~x105 & ~x110 & ~x112 & ~x134 & ~x138 & ~x139 & ~x140 & ~x143 & ~x144 & ~x163 & ~x166 & ~x168 & ~x225 & ~x251 & ~x252 & ~x254 & ~x277 & ~x305 & ~x333 & ~x366 & ~x367 & ~x447 & ~x450 & ~x532 & ~x560 & ~x561 & ~x587 & ~x614 & ~x616 & ~x644 & ~x670 & ~x672 & ~x698 & ~x699 & ~x727 & ~x728 & ~x730 & ~x754 & ~x770 & ~x771 & ~x772 & ~x773 & ~x775 & ~x782;
assign c1375 =  x157 &  x654 & ~x191 & ~x205 & ~x232 & ~x300 & ~x344 & ~x358 & ~x365 & ~x371 & ~x400 & ~x456 & ~x508 & ~x527 & ~x558 & ~x671 & ~x674;
assign c1377 = ~x7 & ~x112 & ~x139 & ~x599 & ~x628 & ~x632 & ~x665 & ~x670 & ~x687 & ~x763;
assign c1379 =  x484 & ~x579;
assign c1381 =  x245 & ~x2 & ~x20 & ~x477 & ~x532 & ~x730;
assign c1383 =  x70 &  x457 & ~x0 & ~x1 & ~x6 & ~x10 & ~x17 & ~x18 & ~x20 & ~x21 & ~x25 & ~x28 & ~x31 & ~x36 & ~x47 & ~x50 & ~x56 & ~x59 & ~x60 & ~x62 & ~x80 & ~x83 & ~x85 & ~x89 & ~x90 & ~x105 & ~x117 & ~x134 & ~x138 & ~x139 & ~x140 & ~x141 & ~x142 & ~x144 & ~x165 & ~x170 & ~x171 & ~x172 & ~x173 & ~x190 & ~x191 & ~x221 & ~x226 & ~x227 & ~x247 & ~x248 & ~x249 & ~x250 & ~x254 & ~x255 & ~x275 & ~x276 & ~x279 & ~x280 & ~x281 & ~x282 & ~x283 & ~x304 & ~x306 & ~x308 & ~x312 & ~x333 & ~x335 & ~x337 & ~x339 & ~x340 & ~x365 & ~x389 & ~x394 & ~x395 & ~x396 & ~x423 & ~x444 & ~x449 & ~x450 & ~x529 & ~x557 & ~x559 & ~x560 & ~x587 & ~x590 & ~x615 & ~x644 & ~x646 & ~x647 & ~x701 & ~x754 & ~x756 & ~x757 & ~x759 & ~x760 & ~x781 & ~x782;
assign c1385 =  x91 & ~x453 & ~x481;
assign c1387 =  x466 & ~x100;
assign c1389 =  x64 &  x76 & ~x54 & ~x281 & ~x307 & ~x310 & ~x446;
assign c1391 =  x739 &  x741 &  x742 &  x745 & ~x54 & ~x129 & ~x194 & ~x218 & ~x448 & ~x450 & ~x502 & ~x697 & ~x704;
assign c1393 =  x186 &  x692 & ~x13;
assign c1395 =  x37 &  x126 &  x127 &  x683 &  x739 &  x740 & ~x587;
assign c1397 =  x322 & ~x710 & ~x743;
assign c1399 =  x411 & ~x42 & ~x67 & ~x111;
assign c1401 =  x387;
assign c1403 =  x682 & ~x19 & ~x519;
assign c1405 =  x436 &  x464 & ~x10 & ~x36 & ~x145 & ~x213 & ~x256 & ~x333 & ~x339 & ~x592 & ~x772 & ~x773;
assign c1407 =  x414 & ~x22 & ~x748;
assign c1409 =  x97 &  x124 &  x377 &  x490 &  x575 &  x656 &  x689 & ~x135 & ~x246 & ~x270 & ~x447 & ~x497 & ~x567;
assign c1411 =  x127 &  x518 &  x600 &  x601 &  x654 & ~x1 & ~x33 & ~x60 & ~x200 & ~x201 & ~x220 & ~x226 & ~x227 & ~x250 & ~x252 & ~x259 & ~x277 & ~x314 & ~x391 & ~x526 & ~x527 & ~x532 & ~x534 & ~x761 & ~x773;
assign c1413 = ~x10 & ~x23 & ~x30 & ~x58 & ~x64 & ~x76 & ~x143 & ~x174 & ~x234 & ~x250 & ~x274 & ~x390 & ~x644 & ~x664 & ~x670 & ~x701 & ~x735 & ~x752 & ~x773;
assign c1415 =  x347 &  x546 &  x603 &  x627 &  x714 & ~x10 & ~x11 & ~x171 & ~x541;
assign c1417 =  x46 &  x661 & ~x260 & ~x539;
assign c1419 =  x733 & ~x775;
assign c1421 =  x715 & ~x182;
assign c1423 =  x385 &  x441 & ~x727 & ~x775;
assign c1425 =  x158 &  x267 &  x435 &  x461 &  x521 &  x571 &  x630 &  x661 &  x740 &  x741 &  x742 & ~x53 & ~x109 & ~x135 & ~x163 & ~x277 & ~x279 & ~x334 & ~x397 & ~x399 & ~x500 & ~x617 & ~x751 & ~x760;
assign c1427 =  x272 & ~x4 & ~x19 & ~x20 & ~x49 & ~x281 & ~x311 & ~x390 & ~x473 & ~x730 & ~x759 & ~x775;
assign c1429 =  x97 &  x151 &  x518 &  x626 &  x686 &  x746 & ~x14 & ~x84 & ~x363 & ~x555 & ~x560 & ~x641 & ~x697;
assign c1431 = ~x14 & ~x23 & ~x29 & ~x33 & ~x58 & ~x140 & ~x142 & ~x192 & ~x306 & ~x391 & ~x419 & ~x500 & ~x507 & ~x530 & ~x532 & ~x547 & ~x584 & ~x618 & ~x756 & ~x777;
assign c1433 =  x681 & ~x45;
assign c1435 =  x518 &  x655 &  x746 &  x769 &  x770 & ~x11 & ~x248 & ~x673;
assign c1437 =  x200 & ~x560;
assign c1439 =  x193;
assign c1441 = ~x7 & ~x13 & ~x14 & ~x35 & ~x53 & ~x66 & ~x113 & ~x131 & ~x139 & ~x140 & ~x194 & ~x234 & ~x363 & ~x759 & ~x763 & ~x773 & ~x777;
assign c1443 =  x415;
assign c1445 = ~x57 & ~x138 & ~x181 & ~x197 & ~x655;
assign c1447 =  x611;
assign c1449 = ~x403 & ~x407 & ~x408 & ~x442;
assign c1451 = ~x86 & ~x514 & ~x575 & ~x584 & ~x587 & ~x656 & ~x657 & ~x763 & ~x777;
assign c1453 =  x40 & ~x550 & ~x626 & ~x662;
assign c1455 = ~x748 & ~x764;
assign c1457 =  x454 & ~x48;
assign c1459 =  x445;
assign c1461 =  x41 &  x157 &  x490 &  x518 &  x546 &  x683 & ~x233 & ~x670;
assign c1463 =  x770 &  x772 & ~x14 & ~x272 & ~x358 & ~x536;
assign c1465 =  x129 &  x156 &  x157 &  x625 & ~x13 & ~x167 & ~x232;
assign c1467 =  x122 &  x129 &  x180 &  x207 &  x208 &  x264 &  x378 &  x406 &  x431 &  x459 &  x462 &  x489 &  x491 &  x517 &  x518 &  x542 &  x570 &  x573 &  x576 &  x632 &  x660 &  x712 & ~x6 & ~x7 & ~x9 & ~x58 & ~x78 & ~x82 & ~x106 & ~x132 & ~x134 & ~x137 & ~x141 & ~x201 & ~x226 & ~x338 & ~x386 & ~x418 & ~x448 & ~x451 & ~x482 & ~x504 & ~x532 & ~x538 & ~x554 & ~x565 & ~x567 & ~x622 & ~x644 & ~x650 & ~x731 & ~x756 & ~x759 & ~x760;
assign c1469 =  x37 &  x493 &  x573 &  x602 & ~x194 & ~x253 & ~x423 & ~x474 & ~x502 & ~x559 & ~x566 & ~x585 & ~x732;
assign c1471 =  x362;
assign c1473 =  x172;
assign c1475 =  x130 &  x157 &  x320 &  x352 &  x491 &  x655 &  x743 &  x745 & ~x11 & ~x332 & ~x673;
assign c1477 = ~x61 & ~x391 & ~x530 & ~x584 & ~x586 & ~x644 & ~x688 & ~x712 & ~x714 & ~x715 & ~x735 & ~x741 & ~x743 & ~x754 & ~x764 & ~x773 & ~x774;
assign c1479 =  x186 &  x625 &  x742 &  x746 & ~x363 & ~x448 & ~x554 & ~x560 & ~x614;
assign c1481 =  x602 &  x633 & ~x184;
assign c1483 = ~x14 & ~x121 & ~x208;
assign c1485 =  x43 &  x546 & ~x60 & ~x78 & ~x105 & ~x134 & ~x139 & ~x143 & ~x589 & ~x765 & ~x767;
assign c1487 =  x174 &  x518;
assign c1489 =  x637 & ~x424;
assign c1491 = ~x21 & ~x150 & ~x152 & ~x209 & ~x761;
assign c1493 =  x658 &  x742 & ~x1 & ~x51 & ~x53 & ~x57 & ~x59 & ~x62 & ~x83 & ~x110 & ~x160 & ~x167 & ~x196 & ~x219 & ~x220 & ~x234 & ~x242 & ~x281 & ~x298 & ~x532;
assign c1495 =  x155 &  x181 &  x658 & ~x166 & ~x206 & ~x242 & ~x503 & ~x726;
assign c1497 =  x407 &  x434 &  x437 &  x459 &  x461 &  x488 &  x514 &  x520 &  x543 &  x547 &  x549 &  x574 &  x575 &  x576 &  x601 &  x602 &  x630 & ~x2 & ~x4 & ~x24 & ~x28 & ~x29 & ~x32 & ~x55 & ~x59 & ~x61 & ~x81 & ~x84 & ~x85 & ~x115 & ~x141 & ~x142 & ~x163 & ~x165 & ~x166 & ~x192 & ~x193 & ~x196 & ~x197 & ~x222 & ~x227 & ~x252 & ~x255 & ~x336 & ~x392 & ~x422 & ~x448 & ~x449 & ~x450 & ~x473 & ~x503 & ~x506 & ~x532 & ~x562 & ~x698 & ~x771 & ~x782;
assign c1499 =  x43 & ~x601 & ~x606;
assign c20 =  x286 &  x342 &  x370 & ~x1 & ~x4 & ~x6 & ~x8 & ~x20 & ~x23 & ~x24 & ~x25 & ~x27 & ~x28 & ~x50 & ~x55 & ~x56 & ~x59 & ~x60 & ~x81 & ~x83 & ~x107 & ~x109 & ~x112 & ~x115 & ~x139 & ~x140 & ~x193 & ~x199 & ~x221 & ~x222 & ~x223 & ~x249 & ~x251 & ~x278 & ~x281 & ~x283 & ~x304 & ~x311 & ~x334 & ~x335 & ~x336 & ~x363 & ~x366 & ~x389 & ~x392 & ~x418 & ~x420 & ~x446 & ~x475 & ~x502 & ~x504 & ~x505 & ~x534 & ~x552 & ~x562 & ~x589 & ~x590 & ~x613 & ~x614 & ~x641 & ~x643 & ~x674 & ~x697 & ~x698 & ~x730 & ~x753 & ~x754 & ~x755 & ~x767 & ~x769 & ~x771 & ~x773;
assign c22 =  x342 &  x566 &  x622 & ~x194 & ~x281 & ~x305 & ~x568 & ~x589 & ~x670 & ~x753 & ~x755;
assign c24 =  x133 &  x146 &  x147 &  x161 &  x271 &  x377 &  x379 &  x382 &  x442 &  x498 &  x550 &  x582 &  x602 &  x607 &  x625 &  x627 &  x629 &  x630 &  x632 &  x639 &  x666 & ~x3 & ~x32 & ~x53 & ~x55 & ~x60 & ~x83 & ~x86 & ~x110 & ~x140 & ~x166 & ~x196 & ~x197 & ~x224 & ~x251 & ~x254 & ~x277 & ~x281 & ~x361 & ~x418 & ~x449 & ~x450 & ~x476 & ~x562 & ~x589 & ~x614 & ~x619 & ~x670 & ~x674 & ~x700 & ~x702 & ~x727 & ~x728 & ~x731 & ~x770 & ~x776 & ~x782;
assign c26 = ~x52 & ~x69 & ~x70 & ~x71 & ~x361 & ~x645 & ~x767 & ~x774;
assign c28 =  x147 &  x161 &  x442 &  x458 &  x572 &  x778 & ~x7 & ~x58 & ~x82 & ~x85 & ~x115 & ~x136 & ~x169 & ~x170 & ~x222 & ~x224 & ~x251 & ~x473 & ~x475 & ~x477 & ~x505 & ~x558 & ~x559 & ~x615 & ~x618 & ~x671 & ~x699 & ~x752 & ~x756 & ~x771 & ~x781 & ~x782;
assign c210 =  x68 &  x98 &  x152 &  x188 &  x215 &  x217 &  x242 &  x243 &  x245 &  x272 &  x402 &  x490 &  x544 &  x576 &  x601 &  x706 &  x749 & ~x3 & ~x27 & ~x30 & ~x54 & ~x61 & ~x107 & ~x135 & ~x144 & ~x165 & ~x248 & ~x253 & ~x254 & ~x306 & ~x366 & ~x388 & ~x392 & ~x393 & ~x395 & ~x450 & ~x477 & ~x478 & ~x503 & ~x533 & ~x560 & ~x563 & ~x613 & ~x616 & ~x645 & ~x668 & ~x779 & ~x782;
assign c212 = ~x70 & ~x227 & ~x249 & ~x305 & ~x361 & ~x421 & ~x747 & ~x765 & ~x773;
assign c214 =  x750 & ~x21 & ~x34 & ~x53 & ~x55 & ~x85 & ~x254 & ~x277 & ~x305 & ~x338 & ~x391 & ~x420 & ~x501 & ~x505 & ~x532 & ~x608 & ~x673 & ~x698 & ~x700 & ~x702 & ~x727 & ~x752 & ~x753 & ~x754 & ~x757;
assign c216 =  x46 &  x257 &  x345 &  x374 &  x564 &  x603 &  x630 &  x632 &  x633 &  x657 &  x659 &  x662 &  x689 & ~x2 & ~x60 & ~x85 & ~x109 & ~x111 & ~x112 & ~x115 & ~x137 & ~x165 & ~x170 & ~x195 & ~x251 & ~x334 & ~x504 & ~x586 & ~x616 & ~x646 & ~x672 & ~x727 & ~x758;
assign c218 =  x526 &  x638 & ~x6 & ~x21 & ~x22 & ~x28 & ~x30 & ~x33 & ~x50 & ~x81 & ~x109 & ~x137 & ~x138 & ~x143 & ~x164 & ~x166 & ~x168 & ~x171 & ~x195 & ~x225 & ~x277 & ~x278 & ~x280 & ~x307 & ~x309 & ~x333 & ~x334 & ~x335 & ~x337 & ~x355 & ~x362 & ~x364 & ~x392 & ~x419 & ~x446 & ~x449 & ~x474 & ~x534 & ~x558 & ~x586 & ~x587 & ~x644 & ~x672 & ~x700 & ~x726 & ~x730 & ~x758 & ~x783;
assign c220 = ~x71 & ~x220 & ~x249 & ~x305 & ~x361 & ~x362 & ~x390 & ~x418 & ~x741;
assign c222 =  x76 &  x104 &  x161 &  x442 &  x498 &  x526 & ~x4 & ~x24 & ~x25 & ~x29 & ~x30 & ~x31 & ~x51 & ~x52 & ~x58 & ~x79 & ~x80 & ~x81 & ~x84 & ~x85 & ~x86 & ~x88 & ~x109 & ~x115 & ~x136 & ~x139 & ~x170 & ~x195 & ~x198 & ~x252 & ~x279 & ~x281 & ~x307 & ~x337 & ~x366 & ~x417 & ~x421 & ~x445 & ~x475 & ~x478 & ~x506 & ~x534 & ~x614 & ~x615 & ~x617 & ~x618 & ~x701 & ~x728 & ~x767 & ~x771;
assign c224 =  x70 &  x572 &  x714 &  x741 &  x770 &  x771 &  x774 & ~x24 & ~x31 & ~x82 & ~x108 & ~x111 & ~x113 & ~x137 & ~x192 & ~x251 & ~x449 & ~x477 & ~x531 & ~x587 & ~x589;
assign c226 =  x74 &  x149 &  x232 &  x357 &  x398 &  x399 &  x402 &  x426 &  x460 &  x462 &  x514 &  x517 &  x518 &  x545 & ~x1 & ~x3 & ~x22 & ~x23 & ~x25 & ~x28 & ~x31 & ~x34 & ~x51 & ~x54 & ~x57 & ~x60 & ~x79 & ~x80 & ~x81 & ~x82 & ~x88 & ~x107 & ~x111 & ~x113 & ~x115 & ~x137 & ~x138 & ~x140 & ~x165 & ~x169 & ~x170 & ~x194 & ~x197 & ~x198 & ~x222 & ~x225 & ~x226 & ~x227 & ~x278 & ~x279 & ~x281 & ~x282 & ~x304 & ~x306 & ~x308 & ~x338 & ~x339 & ~x363 & ~x389 & ~x390 & ~x422 & ~x475 & ~x503 & ~x530 & ~x532 & ~x559 & ~x560 & ~x561 & ~x614 & ~x617 & ~x641 & ~x642 & ~x698 & ~x701 & ~x753 & ~x766 & ~x768 & ~x769 & ~x770 & ~x775;
assign c228 =  x44 &  x119 &  x160 &  x345 &  x351 &  x406 &  x490 &  x659 & ~x7 & ~x84 & ~x111 & ~x194 & ~x197 & ~x254 & ~x255 & ~x312 & ~x332 & ~x336 & ~x340 & ~x365 & ~x388 & ~x505 & ~x506 & ~x584 & ~x699 & ~x727 & ~x730 & ~x752 & ~x756;
assign c230 =  x216 &  x348 &  x413 &  x426 &  x437 &  x441 &  x482 &  x490 &  x566 &  x706 & ~x3 & ~x33 & ~x52 & ~x78 & ~x81 & ~x82 & ~x136 & ~x137 & ~x140 & ~x141 & ~x143 & ~x166 & ~x167 & ~x170 & ~x254 & ~x279 & ~x335 & ~x336 & ~x338 & ~x364 & ~x394 & ~x419 & ~x423 & ~x448 & ~x451 & ~x501 & ~x505 & ~x563 & ~x616 & ~x620 & ~x647 & ~x670 & ~x673 & ~x697 & ~x700 & ~x701 & ~x726 & ~x727 & ~x757;
assign c232 = ~x0 & ~x1 & ~x3 & ~x4 & ~x5 & ~x8 & ~x22 & ~x31 & ~x32 & ~x52 & ~x53 & ~x59 & ~x62 & ~x77 & ~x84 & ~x85 & ~x86 & ~x107 & ~x108 & ~x109 & ~x110 & ~x112 & ~x115 & ~x118 & ~x134 & ~x135 & ~x136 & ~x137 & ~x138 & ~x139 & ~x141 & ~x143 & ~x144 & ~x166 & ~x170 & ~x171 & ~x193 & ~x195 & ~x197 & ~x220 & ~x223 & ~x224 & ~x226 & ~x227 & ~x248 & ~x249 & ~x250 & ~x253 & ~x254 & ~x275 & ~x277 & ~x278 & ~x279 & ~x280 & ~x282 & ~x305 & ~x310 & ~x332 & ~x333 & ~x334 & ~x335 & ~x388 & ~x390 & ~x391 & ~x392 & ~x393 & ~x395 & ~x419 & ~x420 & ~x423 & ~x424 & ~x446 & ~x448 & ~x449 & ~x450 & ~x451 & ~x472 & ~x475 & ~x476 & ~x477 & ~x500 & ~x501 & ~x502 & ~x506 & ~x507 & ~x550 & ~x557 & ~x562 & ~x578 & ~x586 & ~x590 & ~x615 & ~x641 & ~x643 & ~x671 & ~x673 & ~x697 & ~x699 & ~x700 & ~x727 & ~x759 & ~x782 & ~x783;
assign c234 =  x92 &  x105 &  x246 &  x302 &  x639 & ~x2 & ~x114 & ~x193 & ~x221 & ~x223 & ~x391 & ~x560 & ~x588 & ~x641 & ~x753;
assign c236 =  x357 &  x470 & ~x196 & ~x277 & ~x418 & ~x474 & ~x550 & ~x588;
assign c238 =  x38 &  x46 &  x67 &  x162 &  x247 &  x639 & ~x7 & ~x141 & ~x166 & ~x336 & ~x391 & ~x420;
assign c240 =  x389;
assign c242 =  x45 &  x148 &  x161 &  x313 &  x344 &  x414 &  x425 &  x439 &  x454 &  x600 &  x629 &  x630 &  x655 &  x681 &  x683 & ~x1 & ~x20 & ~x32 & ~x61 & ~x83 & ~x87 & ~x114 & ~x165 & ~x171 & ~x335 & ~x337 & ~x363 & ~x365 & ~x367 & ~x389 & ~x449 & ~x451 & ~x531 & ~x590 & ~x647 & ~x703 & ~x730;
assign c244 =  x98 &  x298 &  x299 &  x400 &  x433 &  x574 &  x597 &  x602 &  x654 & ~x20 & ~x22 & ~x49 & ~x57 & ~x61 & ~x112 & ~x170 & ~x221 & ~x227 & ~x248 & ~x254 & ~x275 & ~x282 & ~x303 & ~x309 & ~x311 & ~x332 & ~x333 & ~x338 & ~x362 & ~x364 & ~x393 & ~x443 & ~x448 & ~x450 & ~x474 & ~x476 & ~x480 & ~x502 & ~x507 & ~x531 & ~x556 & ~x562 & ~x589 & ~x591 & ~x697 & ~x729 & ~x730 & ~x731 & ~x751 & ~x754 & ~x782;
assign c246 =  x147 &  x230 &  x370 &  x429 &  x514 &  x666 &  x683 &  x685 &  x686 &  x750 & ~x1 & ~x2 & ~x52 & ~x82 & ~x84 & ~x113 & ~x138 & ~x139 & ~x199 & ~x220 & ~x253 & ~x337 & ~x361 & ~x364 & ~x475 & ~x584 & ~x644 & ~x646 & ~x671 & ~x698 & ~x701 & ~x726 & ~x748 & ~x755 & ~x757;
assign c248 =  x44 &  x45 &  x441 &  x526 &  x638 & ~x1 & ~x2 & ~x3 & ~x6 & ~x14 & ~x20 & ~x22 & ~x23 & ~x24 & ~x27 & ~x28 & ~x34 & ~x49 & ~x50 & ~x55 & ~x56 & ~x57 & ~x58 & ~x60 & ~x61 & ~x80 & ~x83 & ~x88 & ~x107 & ~x108 & ~x109 & ~x111 & ~x114 & ~x115 & ~x140 & ~x165 & ~x224 & ~x226 & ~x250 & ~x254 & ~x277 & ~x279 & ~x306 & ~x307 & ~x308 & ~x336 & ~x337 & ~x361 & ~x362 & ~x364 & ~x365 & ~x392 & ~x394 & ~x418 & ~x422 & ~x478 & ~x503 & ~x529 & ~x558 & ~x561 & ~x613 & ~x617 & ~x618 & ~x643 & ~x674 & ~x700 & ~x701 & ~x702 & ~x726 & ~x730 & ~x754 & ~x756 & ~x758 & ~x782 & ~x783;
assign c250 =  x561;
assign c252 =  x77 &  x527 &  x668 & ~x27 & ~x54 & ~x56 & ~x85 & ~x109 & ~x142 & ~x166 & ~x196 & ~x364 & ~x365 & ~x449 & ~x783;
assign c254 = ~x6 & ~x8 & ~x10 & ~x20 & ~x32 & ~x58 & ~x80 & ~x84 & ~x111 & ~x112 & ~x115 & ~x135 & ~x139 & ~x143 & ~x165 & ~x167 & ~x224 & ~x226 & ~x278 & ~x280 & ~x332 & ~x334 & ~x336 & ~x427 & ~x447 & ~x455 & ~x504 & ~x567 & ~x665 & ~x671 & ~x673;
assign c256 =  x107;
assign c258 =  x244 &  x260 &  x328 &  x376 &  x437 &  x458 &  x460 &  x461 &  x470 &  x483 &  x487 &  x553 &  x554 &  x571 &  x572 &  x622 &  x665 & ~x106 & ~x114 & ~x115 & ~x135 & ~x144 & ~x166 & ~x167 & ~x191 & ~x193 & ~x195 & ~x200 & ~x248 & ~x276 & ~x277 & ~x284 & ~x303 & ~x308 & ~x309 & ~x334 & ~x360 & ~x366 & ~x395 & ~x416 & ~x443 & ~x447 & ~x506 & ~x530 & ~x613 & ~x615 & ~x671 & ~x675 & ~x701 & ~x728;
assign c260 =  x69 &  x188 &  x266 &  x289 &  x316 &  x328 &  x456 &  x514 &  x517 &  x519 &  x573 &  x602 &  x629 &  x653 &  x688 &  x738 &  x772 & ~x7 & ~x29 & ~x56 & ~x83 & ~x113 & ~x136 & ~x167 & ~x221 & ~x224 & ~x225 & ~x226 & ~x279 & ~x337 & ~x366 & ~x417 & ~x671 & ~x726 & ~x730 & ~x781;
assign c262 =  x95 &  x182 &  x244 &  x410 &  x462 &  x490 &  x510 &  x538 &  x568 &  x569 &  x599 &  x605 &  x610 &  x625 &  x627 &  x632 &  x633 &  x666 &  x677 &  x705 & ~x1 & ~x29 & ~x30 & ~x52 & ~x54 & ~x55 & ~x61 & ~x79 & ~x84 & ~x108 & ~x115 & ~x116 & ~x137 & ~x141 & ~x143 & ~x168 & ~x194 & ~x223 & ~x277 & ~x282 & ~x283 & ~x306 & ~x337 & ~x361 & ~x363 & ~x395 & ~x419 & ~x448 & ~x450 & ~x451 & ~x473 & ~x503 & ~x532 & ~x535 & ~x557 & ~x562 & ~x563 & ~x642 & ~x672 & ~x698 & ~x707 & ~x728 & ~x763;
assign c264 = ~x3 & ~x9 & ~x10 & ~x18 & ~x20 & ~x22 & ~x23 & ~x31 & ~x33 & ~x49 & ~x50 & ~x59 & ~x60 & ~x62 & ~x79 & ~x80 & ~x84 & ~x88 & ~x108 & ~x110 & ~x113 & ~x117 & ~x135 & ~x167 & ~x170 & ~x172 & ~x193 & ~x197 & ~x224 & ~x228 & ~x229 & ~x248 & ~x249 & ~x252 & ~x253 & ~x255 & ~x283 & ~x284 & ~x304 & ~x306 & ~x310 & ~x312 & ~x334 & ~x337 & ~x362 & ~x365 & ~x390 & ~x393 & ~x394 & ~x417 & ~x418 & ~x422 & ~x424 & ~x444 & ~x445 & ~x447 & ~x450 & ~x474 & ~x475 & ~x476 & ~x478 & ~x479 & ~x500 & ~x502 & ~x503 & ~x504 & ~x506 & ~x529 & ~x533 & ~x535 & ~x556 & ~x563 & ~x564 & ~x584 & ~x619 & ~x620 & ~x641 & ~x644 & ~x648 & ~x672 & ~x676 & ~x699 & ~x704 & ~x729 & ~x740 & ~x742 & ~x743 & ~x744 & ~x745 & ~x758 & ~x759 & ~x769 & ~x771 & ~x773 & ~x780 & ~x781 & ~x783;
assign c266 =  x38 &  x703;
assign c268 =  x44 & ~x1 & ~x2 & ~x4 & ~x7 & ~x8 & ~x9 & ~x19 & ~x20 & ~x21 & ~x27 & ~x31 & ~x34 & ~x35 & ~x49 & ~x52 & ~x53 & ~x56 & ~x58 & ~x61 & ~x79 & ~x81 & ~x83 & ~x85 & ~x87 & ~x88 & ~x112 & ~x113 & ~x136 & ~x137 & ~x138 & ~x140 & ~x142 & ~x143 & ~x194 & ~x196 & ~x197 & ~x198 & ~x199 & ~x221 & ~x222 & ~x223 & ~x227 & ~x254 & ~x279 & ~x283 & ~x304 & ~x309 & ~x333 & ~x334 & ~x337 & ~x362 & ~x366 & ~x390 & ~x392 & ~x393 & ~x417 & ~x418 & ~x420 & ~x448 & ~x450 & ~x477 & ~x497 & ~x503 & ~x525 & ~x558 & ~x587 & ~x588 & ~x589 & ~x615 & ~x643 & ~x644 & ~x700;
assign c270 =  x644;
assign c272 =  x592 &  x596 & ~x0 & ~x3 & ~x4 & ~x5 & ~x23 & ~x24 & ~x26 & ~x27 & ~x28 & ~x29 & ~x30 & ~x31 & ~x52 & ~x53 & ~x55 & ~x58 & ~x59 & ~x82 & ~x87 & ~x109 & ~x110 & ~x111 & ~x113 & ~x140 & ~x141 & ~x142 & ~x166 & ~x168 & ~x194 & ~x195 & ~x196 & ~x197 & ~x222 & ~x225 & ~x226 & ~x250 & ~x253 & ~x278 & ~x279 & ~x281 & ~x307 & ~x308 & ~x335 & ~x336 & ~x337 & ~x362 & ~x363 & ~x393 & ~x419 & ~x421 & ~x448 & ~x449 & ~x476 & ~x504 & ~x560 & ~x589 & ~x699 & ~x700 & ~x706 & ~x729 & ~x756 & ~x757 & ~x782;
assign c274 =  x232 & ~x82 & ~x107 & ~x248 & ~x250 & ~x364 & ~x393 & ~x421 & ~x444 & ~x471 & ~x472 & ~x699 & ~x730 & ~x741 & ~x742 & ~x743 & ~x745 & ~x767 & ~x782;
assign c276 = ~x70 & ~x71 & ~x350;
assign c278 =  x450 & ~x649;
assign c280 =  x71 &  x259 &  x272 &  x314 &  x329 &  x385 &  x406 &  x426 &  x431 &  x459 &  x518 &  x523 &  x566 &  x599 &  x631 &  x658 &  x682 &  x706 &  x709 &  x711 &  x715 & ~x20 & ~x34 & ~x54 & ~x55 & ~x59 & ~x64 & ~x107 & ~x172 & ~x222 & ~x228 & ~x250 & ~x278 & ~x306 & ~x335 & ~x392 & ~x417 & ~x418 & ~x505 & ~x507 & ~x530 & ~x531 & ~x562 & ~x563 & ~x590 & ~x644 & ~x703 & ~x754 & ~x756 & ~x758;
assign c282 =  x431 &  x565 &  x593 &  x621 &  x627 &  x649 & ~x1 & ~x4 & ~x6 & ~x23 & ~x26 & ~x27 & ~x29 & ~x31 & ~x50 & ~x53 & ~x56 & ~x57 & ~x80 & ~x82 & ~x85 & ~x108 & ~x109 & ~x110 & ~x111 & ~x112 & ~x113 & ~x114 & ~x115 & ~x142 & ~x165 & ~x167 & ~x169 & ~x170 & ~x194 & ~x197 & ~x223 & ~x227 & ~x249 & ~x278 & ~x281 & ~x305 & ~x306 & ~x307 & ~x308 & ~x310 & ~x338 & ~x361 & ~x367 & ~x391 & ~x392 & ~x394 & ~x419 & ~x420 & ~x422 & ~x447 & ~x476 & ~x477 & ~x504 & ~x505 & ~x506 & ~x531 & ~x532 & ~x562 & ~x586 & ~x588 & ~x589 & ~x616 & ~x617 & ~x618 & ~x642 & ~x644 & ~x651 & ~x671 & ~x672 & ~x679 & ~x701 & ~x726 & ~x735 & ~x756 & ~x757 & ~x763 & ~x767 & ~x769 & ~x771 & ~x774 & ~x775;
assign c284 =  x192 &  x339;
assign c286 =  x734 &  x762 & ~x0 & ~x3 & ~x4 & ~x26 & ~x29 & ~x35 & ~x52 & ~x56 & ~x58 & ~x60 & ~x61 & ~x79 & ~x86 & ~x88 & ~x107 & ~x110 & ~x111 & ~x114 & ~x116 & ~x138 & ~x139 & ~x142 & ~x144 & ~x145 & ~x166 & ~x173 & ~x195 & ~x198 & ~x221 & ~x223 & ~x226 & ~x249 & ~x277 & ~x279 & ~x282 & ~x283 & ~x308 & ~x310 & ~x333 & ~x334 & ~x336 & ~x340 & ~x360 & ~x361 & ~x363 & ~x367 & ~x393 & ~x394 & ~x395 & ~x416 & ~x449 & ~x475 & ~x476 & ~x530 & ~x533 & ~x535 & ~x562 & ~x564 & ~x586 & ~x592 & ~x613 & ~x614 & ~x642 & ~x647 & ~x648 & ~x669 & ~x670 & ~x699 & ~x700 & ~x702 & ~x703 & ~x757 & ~x760 & ~x766 & ~x780;
assign c288 =  x314 &  x342 &  x398 & ~x427;
assign c290 =  x235 &  x298 &  x299 &  x517 &  x597 & ~x1 & ~x4 & ~x23 & ~x53 & ~x83 & ~x84 & ~x87 & ~x112 & ~x164 & ~x169 & ~x196 & ~x252 & ~x255 & ~x280 & ~x283 & ~x284 & ~x304 & ~x367 & ~x419 & ~x420 & ~x476 & ~x615 & ~x694 & ~x722;
assign c292 =  x367 & ~x138 & ~x677;
assign c294 =  x77 &  x430 &  x486 &  x542 & ~x81 & ~x138 & ~x169 & ~x224 & ~x475;
assign c296 = ~x0 & ~x1 & ~x2 & ~x3 & ~x4 & ~x7 & ~x8 & ~x9 & ~x12 & ~x21 & ~x24 & ~x25 & ~x28 & ~x31 & ~x34 & ~x35 & ~x49 & ~x50 & ~x53 & ~x54 & ~x55 & ~x56 & ~x58 & ~x60 & ~x61 & ~x62 & ~x77 & ~x78 & ~x79 & ~x81 & ~x82 & ~x84 & ~x85 & ~x88 & ~x89 & ~x107 & ~x108 & ~x109 & ~x115 & ~x117 & ~x135 & ~x137 & ~x140 & ~x141 & ~x164 & ~x165 & ~x166 & ~x172 & ~x192 & ~x193 & ~x194 & ~x195 & ~x196 & ~x197 & ~x198 & ~x199 & ~x200 & ~x222 & ~x224 & ~x225 & ~x248 & ~x249 & ~x250 & ~x253 & ~x254 & ~x255 & ~x278 & ~x279 & ~x280 & ~x282 & ~x283 & ~x304 & ~x306 & ~x308 & ~x311 & ~x332 & ~x333 & ~x334 & ~x336 & ~x337 & ~x361 & ~x362 & ~x363 & ~x366 & ~x367 & ~x388 & ~x389 & ~x392 & ~x393 & ~x418 & ~x419 & ~x421 & ~x422 & ~x445 & ~x446 & ~x448 & ~x450 & ~x474 & ~x477 & ~x478 & ~x479 & ~x502 & ~x503 & ~x504 & ~x505 & ~x506 & ~x529 & ~x532 & ~x533 & ~x534 & ~x559 & ~x560 & ~x562 & ~x585 & ~x586 & ~x587 & ~x589 & ~x591 & ~x614 & ~x615 & ~x616 & ~x618 & ~x619 & ~x641 & ~x642 & ~x643 & ~x644 & ~x646 & ~x647 & ~x670 & ~x671 & ~x672 & ~x673 & ~x674 & ~x675 & ~x698 & ~x702 & ~x704 & ~x727 & ~x728 & ~x729 & ~x730 & ~x754 & ~x756 & ~x757 & ~x758 & ~x760 & ~x764 & ~x765 & ~x766 & ~x768 & ~x770 & ~x771 & ~x781 & ~x782 & ~x783;
assign c298 =  x527 & ~x638;
assign c2100 = ~x77 & ~x133 & ~x425 & ~x543 & ~x573;
assign c2102 =  x95 &  x160 &  x403 &  x464 &  x468 &  x545 &  x710 &  x778 & ~x61 & ~x88 & ~x116 & ~x166 & ~x171 & ~x200 & ~x223 & ~x284 & ~x420 & ~x448 & ~x449 & ~x473 & ~x476;
assign c2104 =  x39 &  x44 &  x191 &  x527 & ~x31 & ~x32 & ~x226 & ~x250 & ~x281 & ~x310 & ~x505 & ~x534 & ~x643;
assign c2106 =  x750 & ~x7 & ~x23 & ~x28 & ~x57 & ~x107 & ~x110 & ~x111 & ~x114 & ~x144 & ~x164 & ~x168 & ~x192 & ~x194 & ~x197 & ~x220 & ~x221 & ~x252 & ~x254 & ~x278 & ~x306 & ~x334 & ~x336 & ~x337 & ~x363 & ~x364 & ~x391 & ~x416 & ~x420 & ~x446 & ~x451 & ~x473 & ~x479 & ~x527 & ~x563 & ~x617 & ~x698 & ~x726 & ~x728 & ~x758 & ~x765 & ~x768 & ~x770 & ~x771 & ~x773;
assign c2108 =  x587;
assign c2110 =  x38 &  x39 &  x469 & ~x31 & ~x138 & ~x221 & ~x334 & ~x366 & ~x389 & ~x448 & ~x473 & ~x474 & ~x585 & ~x726;
assign c2112 =  x37 &  x38 &  x145 &  x592 &  x629 & ~x0 & ~x3 & ~x24 & ~x32 & ~x57 & ~x82 & ~x141 & ~x225 & ~x281 & ~x308 & ~x419 & ~x421 & ~x447 & ~x476;
assign c2114 =  x96 &  x514 &  x626 &  x627 &  x630 &  x654 &  x655 &  x657 &  x722 &  x750 & ~x19 & ~x23 & ~x24 & ~x58 & ~x60 & ~x108 & ~x111 & ~x138 & ~x141 & ~x171 & ~x221 & ~x224 & ~x227 & ~x253 & ~x279 & ~x281 & ~x283 & ~x308 & ~x311 & ~x338 & ~x364 & ~x389 & ~x393 & ~x445 & ~x446 & ~x449 & ~x451 & ~x477 & ~x530 & ~x535 & ~x559 & ~x561 & ~x590 & ~x591 & ~x645 & ~x671 & ~x673 & ~x698 & ~x701 & ~x725 & ~x731 & ~x735 & ~x756 & ~x765 & ~x766 & ~x768 & ~x769 & ~x770 & ~x771 & ~x772;
assign c2116 =  x228 &  x452 &  x709 &  x712 &  x713 &  x717 & ~x24 & ~x33 & ~x194 & ~x363;
assign c2118 =  x201 &  x387 &  x415 & ~x1 & ~x56 & ~x87 & ~x136 & ~x171 & ~x250 & ~x255 & ~x280 & ~x307 & ~x308 & ~x310 & ~x422 & ~x446 & ~x559 & ~x561 & ~x585 & ~x614 & ~x642 & ~x646 & ~x673 & ~x725 & ~x758 & ~x783;
assign c2120 =  x131 &  x174 &  x212 & ~x4 & ~x12 & ~x15 & ~x21 & ~x57 & ~x363;
assign c2122 =  x42 & ~x29 & ~x97 & ~x98 & ~x99 & ~x164 & ~x220 & ~x337 & ~x392 & ~x421 & ~x473 & ~x501 & ~x504 & ~x559 & ~x585 & ~x615 & ~x757;
assign c2124 = ~x3 & ~x5 & ~x29 & ~x110 & ~x162 & ~x166 & ~x168 & ~x249 & ~x276 & ~x277 & ~x282 & ~x339 & ~x362 & ~x365 & ~x367 & ~x390 & ~x417 & ~x422 & ~x447 & ~x448 & ~x501 & ~x502 & ~x506 & ~x533 & ~x588 & ~x615 & ~x626 & ~x629 & ~x632 & ~x633 & ~x675 & ~x783;
assign c2126 =  x39 & ~x26 & ~x53 & ~x87 & ~x168 & ~x198 & ~x210 & ~x276 & ~x277 & ~x280 & ~x308 & ~x393 & ~x419 & ~x420 & ~x641 & ~x644;
assign c2128 =  x39 &  x358 &  x482 &  x510 &  x610 & ~x0 & ~x1 & ~x3 & ~x6 & ~x12 & ~x13 & ~x25 & ~x27 & ~x31 & ~x57 & ~x58 & ~x61 & ~x111 & ~x112 & ~x142 & ~x167 & ~x221 & ~x222 & ~x225 & ~x249 & ~x251 & ~x252 & ~x253 & ~x279 & ~x283 & ~x306 & ~x309 & ~x334 & ~x336 & ~x420 & ~x448 & ~x449 & ~x474 & ~x476 & ~x504 & ~x560 & ~x588 & ~x614 & ~x645 & ~x646 & ~x673 & ~x702 & ~x756 & ~x757;
assign c2130 =  x508 & ~x638;
assign c2132 =  x385 & ~x26 & ~x384 & ~x644;
assign c2134 =  x749 & ~x28 & ~x49 & ~x59 & ~x83 & ~x85 & ~x109 & ~x145 & ~x193 & ~x196 & ~x199 & ~x251 & ~x304 & ~x335 & ~x339 & ~x364 & ~x421 & ~x446 & ~x447 & ~x451 & ~x505 & ~x531 & ~x561 & ~x564 & ~x620 & ~x640 & ~x727 & ~x728 & ~x729 & ~x755 & ~x768 & ~x771 & ~x779 & ~x783;
assign c2136 = ~x0 & ~x1 & ~x2 & ~x4 & ~x5 & ~x6 & ~x7 & ~x21 & ~x22 & ~x27 & ~x28 & ~x34 & ~x49 & ~x52 & ~x53 & ~x55 & ~x56 & ~x61 & ~x78 & ~x82 & ~x84 & ~x85 & ~x86 & ~x87 & ~x88 & ~x105 & ~x107 & ~x108 & ~x109 & ~x115 & ~x116 & ~x135 & ~x136 & ~x137 & ~x140 & ~x141 & ~x143 & ~x164 & ~x165 & ~x167 & ~x169 & ~x171 & ~x185 & ~x186 & ~x199 & ~x200 & ~x220 & ~x222 & ~x224 & ~x225 & ~x226 & ~x227 & ~x248 & ~x249 & ~x250 & ~x251 & ~x254 & ~x276 & ~x277 & ~x278 & ~x279 & ~x280 & ~x281 & ~x282 & ~x283 & ~x305 & ~x308 & ~x309 & ~x310 & ~x311 & ~x332 & ~x333 & ~x334 & ~x336 & ~x338 & ~x339 & ~x362 & ~x363 & ~x364 & ~x365 & ~x367 & ~x388 & ~x389 & ~x390 & ~x392 & ~x393 & ~x394 & ~x395 & ~x417 & ~x418 & ~x422 & ~x423 & ~x448 & ~x449 & ~x474 & ~x475 & ~x476 & ~x477 & ~x478 & ~x501 & ~x528 & ~x530 & ~x532 & ~x533 & ~x535 & ~x557 & ~x558 & ~x560 & ~x561 & ~x584 & ~x585 & ~x588 & ~x612 & ~x614 & ~x615 & ~x617 & ~x643 & ~x646 & ~x669 & ~x672 & ~x673 & ~x674 & ~x697 & ~x702 & ~x724 & ~x728 & ~x730 & ~x753 & ~x754 & ~x755 & ~x757 & ~x764 & ~x781 & ~x783;
assign c2138 = ~x59 & ~x98 & ~x276 & ~x277 & ~x337 & ~x361 & ~x726 & ~x736 & ~x738 & ~x746;
assign c2140 =  x11 &  x16 &  x44 &  x750 & ~x1 & ~x3 & ~x6 & ~x34 & ~x54 & ~x57 & ~x82 & ~x115 & ~x138 & ~x140 & ~x166 & ~x196 & ~x221 & ~x305 & ~x308 & ~x333 & ~x506 & ~x529 & ~x533 & ~x617 & ~x730 & ~x754 & ~x763;
assign c2142 =  x45 & ~x27 & ~x59 & ~x112 & ~x114 & ~x115 & ~x166 & ~x182 & ~x197 & ~x220 & ~x252 & ~x277 & ~x281 & ~x361 & ~x362 & ~x421 & ~x474 & ~x559 & ~x616 & ~x670 & ~x782;
assign c2144 =  x11 &  x65 &  x92 &  x124 &  x147 &  x149 &  x189 &  x261 &  x343 &  x358 &  x381 &  x382 &  x406 &  x410 &  x466 &  x521 &  x607 & ~x20 & ~x59 & ~x138 & ~x167 & ~x362 & ~x364 & ~x392 & ~x478 & ~x506 & ~x530 & ~x533 & ~x558 & ~x590 & ~x617 & ~x674 & ~x701 & ~x728;
assign c2146 =  x385 & ~x31 & ~x179 & ~x334 & ~x360 & ~x363 & ~x416 & ~x418 & ~x501 & ~x557 & ~x561 & ~x585 & ~x673;
assign c2148 =  x10 &  x620 & ~x6 & ~x21 & ~x22 & ~x23 & ~x25 & ~x26 & ~x31 & ~x59 & ~x60 & ~x82 & ~x84 & ~x278 & ~x447 & ~x616;
assign c2150 =  x45 &  x95 &  x130 &  x203 &  x217 &  x498 &  x574 &  x575 &  x632 &  x634 &  x656 &  x658 &  x737 &  x742 &  x744 & ~x1 & ~x3 & ~x22 & ~x30 & ~x52 & ~x110 & ~x138 & ~x140 & ~x223 & ~x249 & ~x339 & ~x364 & ~x390 & ~x420 & ~x421 & ~x446 & ~x449 & ~x475 & ~x562 & ~x589 & ~x618 & ~x731 & ~x753 & ~x782;
assign c2152 =  x45 & ~x195 & ~x210 & ~x754;
assign c2154 = ~x31 & ~x50 & ~x54 & ~x58 & ~x80 & ~x85 & ~x86 & ~x109 & ~x113 & ~x115 & ~x138 & ~x139 & ~x141 & ~x164 & ~x192 & ~x193 & ~x227 & ~x248 & ~x251 & ~x254 & ~x277 & ~x305 & ~x335 & ~x349 & ~x350 & ~x366 & ~x389 & ~x390 & ~x395 & ~x419 & ~x448 & ~x450 & ~x473 & ~x475 & ~x478 & ~x529 & ~x531 & ~x557 & ~x561 & ~x585 & ~x587 & ~x588 & ~x614 & ~x643 & ~x697 & ~x700 & ~x701 & ~x765 & ~x767 & ~x768 & ~x769 & ~x770 & ~x771 & ~x774;
assign c2156 = ~x0 & ~x2 & ~x3 & ~x9 & ~x20 & ~x21 & ~x26 & ~x28 & ~x29 & ~x32 & ~x49 & ~x52 & ~x54 & ~x55 & ~x57 & ~x58 & ~x60 & ~x80 & ~x81 & ~x82 & ~x83 & ~x86 & ~x107 & ~x111 & ~x114 & ~x136 & ~x137 & ~x138 & ~x139 & ~x143 & ~x144 & ~x167 & ~x192 & ~x193 & ~x194 & ~x195 & ~x197 & ~x198 & ~x199 & ~x220 & ~x224 & ~x227 & ~x249 & ~x251 & ~x252 & ~x253 & ~x254 & ~x255 & ~x278 & ~x279 & ~x281 & ~x282 & ~x283 & ~x304 & ~x306 & ~x307 & ~x308 & ~x309 & ~x333 & ~x334 & ~x336 & ~x362 & ~x365 & ~x391 & ~x393 & ~x395 & ~x417 & ~x418 & ~x419 & ~x420 & ~x421 & ~x423 & ~x428 & ~x445 & ~x446 & ~x447 & ~x448 & ~x449 & ~x451 & ~x456 & ~x473 & ~x474 & ~x476 & ~x501 & ~x503 & ~x505 & ~x507 & ~x529 & ~x530 & ~x535 & ~x557 & ~x558 & ~x559 & ~x561 & ~x562 & ~x563 & ~x585 & ~x587 & ~x588 & ~x613 & ~x614 & ~x615 & ~x617 & ~x619 & ~x641 & ~x642 & ~x643 & ~x644 & ~x670 & ~x672 & ~x673 & ~x675 & ~x697 & ~x699 & ~x700 & ~x725 & ~x726 & ~x728 & ~x729 & ~x740 & ~x741 & ~x744 & ~x754 & ~x756 & ~x759 & ~x764 & ~x766 & ~x767 & ~x768 & ~x769 & ~x772 & ~x773 & ~x781;
assign c2158 =  x76 &  x163 &  x388;
assign c2160 =  x45 & ~x268;
assign c2162 =  x37 &  x46 &  x256 &  x380 & ~x363;
assign c2164 =  x77 &  x218 &  x290 &  x442 & ~x1 & ~x3 & ~x22 & ~x32 & ~x52 & ~x54 & ~x56 & ~x60 & ~x81 & ~x83 & ~x108 & ~x111 & ~x112 & ~x138 & ~x141 & ~x165 & ~x195 & ~x196 & ~x197 & ~x279 & ~x307 & ~x308 & ~x335 & ~x364 & ~x448 & ~x476 & ~x700 & ~x728;
assign c2166 = ~x0 & ~x1 & ~x2 & ~x4 & ~x7 & ~x21 & ~x22 & ~x23 & ~x26 & ~x27 & ~x30 & ~x32 & ~x33 & ~x35 & ~x50 & ~x51 & ~x52 & ~x53 & ~x54 & ~x79 & ~x80 & ~x83 & ~x89 & ~x107 & ~x108 & ~x109 & ~x116 & ~x137 & ~x138 & ~x170 & ~x171 & ~x196 & ~x199 & ~x220 & ~x221 & ~x228 & ~x250 & ~x278 & ~x306 & ~x307 & ~x308 & ~x310 & ~x338 & ~x339 & ~x361 & ~x362 & ~x389 & ~x390 & ~x391 & ~x395 & ~x417 & ~x421 & ~x422 & ~x423 & ~x445 & ~x446 & ~x448 & ~x474 & ~x477 & ~x478 & ~x502 & ~x505 & ~x507 & ~x531 & ~x533 & ~x534 & ~x535 & ~x558 & ~x560 & ~x561 & ~x562 & ~x563 & ~x585 & ~x588 & ~x591 & ~x595 & ~x615 & ~x616 & ~x617 & ~x619 & ~x642 & ~x700 & ~x701 & ~x738 & ~x739 & ~x741 & ~x743 & ~x753 & ~x754 & ~x755 & ~x758 & ~x759 & ~x766 & ~x769 & ~x770 & ~x772 & ~x773 & ~x783;
assign c2168 =  x40 &  x68 &  x72 &  x96 &  x127 &  x234 &  x268 &  x289 &  x299 &  x659 &  x710 &  x711 &  x742 & ~x0 & ~x37 & ~x55 & ~x64 & ~x85 & ~x88 & ~x117 & ~x118 & ~x140 & ~x166 & ~x167 & ~x226 & ~x252 & ~x280 & ~x311 & ~x332 & ~x338 & ~x363 & ~x395 & ~x417 & ~x419 & ~x446 & ~x614 & ~x616 & ~x645 & ~x646 & ~x670 & ~x698 & ~x699 & ~x727 & ~x728 & ~x760;
assign c2170 =  x42 &  x69 &  x71 &  x381 &  x454 &  x462 &  x464 &  x469 &  x545 &  x566 &  x573 &  x734 & ~x6 & ~x7 & ~x24 & ~x25 & ~x49 & ~x192 & ~x199 & ~x283 & ~x362 & ~x394 & ~x477 & ~x507 & ~x561 & ~x648 & ~x669 & ~x670 & ~x760;
assign c2172 = ~x244 & ~x272 & ~x382 & ~x519;
assign c2174 =  x160 &  x218 &  x274 &  x357 &  x375 &  x493 &  x604 &  x629 &  x631 &  x655 &  x662 &  x750 & ~x113 & ~x225 & ~x418 & ~x500 & ~x528 & ~x645;
assign c2176 = ~x20 & ~x21 & ~x29 & ~x30 & ~x31 & ~x57 & ~x80 & ~x81 & ~x103 & ~x104 & ~x128 & ~x131 & ~x135 & ~x141 & ~x142 & ~x158 & ~x193 & ~x196 & ~x199 & ~x220 & ~x227 & ~x248 & ~x252 & ~x304 & ~x333 & ~x338 & ~x392 & ~x395 & ~x448 & ~x450 & ~x473 & ~x477 & ~x478 & ~x507 & ~x529 & ~x530 & ~x535 & ~x557 & ~x558 & ~x563 & ~x613 & ~x616 & ~x645 & ~x646 & ~x669 & ~x728 & ~x756 & ~x758 & ~x759;
assign c2178 =  x287 &  x315 &  x779 & ~x1 & ~x108 & ~x199 & ~x311 & ~x363 & ~x364 & ~x393 & ~x473 & ~x503 & ~x505 & ~x529 & ~x531 & ~x535 & ~x588 & ~x589 & ~x590 & ~x616 & ~x641 & ~x674 & ~x702 & ~x730 & ~x753 & ~x763 & ~x769 & ~x771 & ~x773;
assign c2180 =  x44 &  x68 &  x122 &  x323 &  x484 &  x518 &  x571 &  x625 &  x634 &  x657 &  x717 &  x718 &  x737 & ~x28 & ~x50 & ~x77 & ~x165 & ~x171 & ~x192 & ~x249 & ~x251 & ~x252 & ~x562 & ~x591 & ~x614 & ~x697 & ~x731;
assign c2182 =  x408 & ~x0 & ~x22 & ~x55 & ~x111 & ~x115 & ~x137 & ~x143 & ~x164 & ~x192 & ~x224 & ~x250 & ~x253 & ~x254 & ~x310 & ~x337 & ~x361 & ~x364 & ~x390 & ~x477 & ~x478 & ~x531 & ~x562 & ~x586 & ~x587 & ~x618 & ~x624 & ~x699 & ~x701 & ~x729 & ~x738 & ~x741 & ~x743 & ~x744 & ~x746 & ~x747 & ~x759 & ~x768 & ~x774;
assign c2186 =  x542 &  x571 &  x628 &  x649 & ~x8 & ~x25 & ~x61 & ~x82 & ~x114 & ~x116 & ~x196 & ~x224 & ~x252 & ~x278 & ~x306 & ~x307 & ~x332 & ~x335 & ~x336 & ~x473 & ~x479 & ~x591 & ~x673 & ~x702 & ~x735 & ~x743 & ~x744 & ~x763 & ~x776;
assign c2188 =  x348 &  x441 &  x469 & ~x0 & ~x53 & ~x54 & ~x55 & ~x80 & ~x83 & ~x113 & ~x115 & ~x139 & ~x142 & ~x220 & ~x222 & ~x224 & ~x248 & ~x249 & ~x279 & ~x310 & ~x337 & ~x363 & ~x391 & ~x393 & ~x418 & ~x445 & ~x474 & ~x475 & ~x478 & ~x495 & ~x504 & ~x532 & ~x561 & ~x589 & ~x590 & ~x615 & ~x617 & ~x618 & ~x729 & ~x756;
assign c2190 = ~x126 & ~x418 & ~x439 & ~x467;
assign c2192 =  x385 & ~x2 & ~x3 & ~x5 & ~x6 & ~x26 & ~x29 & ~x32 & ~x50 & ~x51 & ~x52 & ~x60 & ~x80 & ~x82 & ~x84 & ~x110 & ~x113 & ~x114 & ~x136 & ~x141 & ~x165 & ~x168 & ~x170 & ~x196 & ~x197 & ~x227 & ~x251 & ~x281 & ~x283 & ~x305 & ~x308 & ~x334 & ~x337 & ~x339 & ~x355 & ~x366 & ~x392 & ~x394 & ~x421 & ~x446 & ~x448 & ~x449 & ~x475 & ~x530 & ~x559 & ~x587 & ~x588 & ~x617 & ~x643 & ~x645 & ~x673 & ~x702 & ~x728 & ~x773 & ~x783;
assign c2194 =  x264 & ~x537 & ~x649 & ~x748;
assign c2196 =  x654 &  x656 &  x659 &  x710 &  x711 &  x712 &  x713 &  x715 & ~x3 & ~x15 & ~x22 & ~x50 & ~x51 & ~x54 & ~x57 & ~x88 & ~x114 & ~x116 & ~x194 & ~x251 & ~x729 & ~x734 & ~x755;
assign c2198 = ~x1 & ~x4 & ~x6 & ~x7 & ~x22 & ~x23 & ~x27 & ~x49 & ~x83 & ~x86 & ~x87 & ~x107 & ~x108 & ~x112 & ~x135 & ~x138 & ~x140 & ~x141 & ~x171 & ~x193 & ~x195 & ~x220 & ~x226 & ~x248 & ~x253 & ~x277 & ~x278 & ~x282 & ~x306 & ~x307 & ~x334 & ~x365 & ~x417 & ~x418 & ~x420 & ~x425 & ~x448 & ~x475 & ~x501 & ~x530 & ~x534 & ~x557 & ~x558 & ~x559 & ~x562 & ~x563 & ~x585 & ~x586 & ~x612 & ~x613 & ~x617 & ~x618 & ~x643 & ~x697 & ~x699 & ~x701 & ~x730 & ~x739 & ~x740 & ~x741 & ~x742 & ~x743 & ~x744 & ~x745 & ~x746 & ~x747 & ~x755 & ~x756 & ~x767 & ~x769 & ~x772 & ~x775;
assign c2200 =  x367;
assign c2202 =  x39 &  x259 &  x260 &  x413 &  x706 & ~x32 & ~x52 & ~x53 & ~x58 & ~x107 & ~x114 & ~x139 & ~x167 & ~x170 & ~x221 & ~x225 & ~x248 & ~x338 & ~x417 & ~x508 & ~x534 & ~x645 & ~x726 & ~x753 & ~x757 & ~x781;
assign c2204 =  x582 &  x638 &  x666 & ~x23 & ~x25 & ~x27 & ~x51 & ~x56 & ~x59 & ~x80 & ~x82 & ~x85 & ~x138 & ~x165 & ~x194 & ~x195 & ~x306 & ~x333 & ~x337 & ~x365 & ~x391 & ~x446 & ~x447 & ~x502 & ~x531 & ~x557 & ~x580 & ~x590 & ~x608 & ~x614 & ~x617 & ~x645 & ~x700 & ~x754 & ~x755 & ~x770;
assign c2206 =  x727;
assign c2208 =  x71 &  x120 &  x161 &  x301 &  x314 &  x426 &  x540 &  x568 &  x581 &  x634 &  x654 &  x655 &  x660 &  x677 &  x689 &  x709 &  x711 &  x717 & ~x2 & ~x28 & ~x107 & ~x141 & ~x249 & ~x283 & ~x534 & ~x591 & ~x673 & ~x702;
assign c2210 =  x318 &  x426 & ~x523;
assign c2212 =  x456 &  x499 & ~x7 & ~x15 & ~x27 & ~x62 & ~x80 & ~x109 & ~x111 & ~x168 & ~x221;
assign c2214 = ~x356 & ~x743 & ~x744;
assign c2218 = ~x1 & ~x2 & ~x5 & ~x6 & ~x9 & ~x18 & ~x20 & ~x22 & ~x26 & ~x27 & ~x29 & ~x31 & ~x33 & ~x53 & ~x57 & ~x59 & ~x61 & ~x79 & ~x84 & ~x86 & ~x88 & ~x91 & ~x104 & ~x107 & ~x109 & ~x110 & ~x112 & ~x115 & ~x116 & ~x137 & ~x138 & ~x139 & ~x141 & ~x142 & ~x164 & ~x167 & ~x168 & ~x169 & ~x170 & ~x172 & ~x191 & ~x192 & ~x197 & ~x198 & ~x221 & ~x222 & ~x223 & ~x224 & ~x226 & ~x227 & ~x249 & ~x252 & ~x253 & ~x254 & ~x255 & ~x276 & ~x277 & ~x281 & ~x283 & ~x304 & ~x305 & ~x307 & ~x308 & ~x309 & ~x310 & ~x311 & ~x332 & ~x334 & ~x337 & ~x360 & ~x364 & ~x366 & ~x367 & ~x389 & ~x390 & ~x391 & ~x393 & ~x395 & ~x439 & ~x446 & ~x448 & ~x450 & ~x467 & ~x473 & ~x474 & ~x476 & ~x500 & ~x501 & ~x502 & ~x503 & ~x505 & ~x506 & ~x529 & ~x530 & ~x531 & ~x532 & ~x558 & ~x559 & ~x560 & ~x562 & ~x585 & ~x586 & ~x587 & ~x588 & ~x614 & ~x615 & ~x617 & ~x641 & ~x642 & ~x645 & ~x648 & ~x670 & ~x671 & ~x673 & ~x698 & ~x699 & ~x701 & ~x726 & ~x727 & ~x729 & ~x756 & ~x767 & ~x768 & ~x769 & ~x772 & ~x775;
assign c2220 = ~x0 & ~x4 & ~x5 & ~x24 & ~x27 & ~x30 & ~x31 & ~x32 & ~x52 & ~x54 & ~x55 & ~x56 & ~x80 & ~x82 & ~x83 & ~x110 & ~x111 & ~x138 & ~x141 & ~x142 & ~x167 & ~x169 & ~x198 & ~x223 & ~x224 & ~x226 & ~x250 & ~x253 & ~x254 & ~x277 & ~x278 & ~x279 & ~x280 & ~x281 & ~x306 & ~x308 & ~x356 & ~x363 & ~x365 & ~x391 & ~x393 & ~x447 & ~x475 & ~x503 & ~x532 & ~x559 & ~x560 & ~x587 & ~x616 & ~x643 & ~x672 & ~x729 & ~x739 & ~x763 & ~x766 & ~x768 & ~x772 & ~x773 & ~x775 & ~x776 & ~x777 & ~x782 & ~x783;
assign c2222 =  x299 & ~x3 & ~x4 & ~x6 & ~x8 & ~x19 & ~x22 & ~x24 & ~x28 & ~x29 & ~x30 & ~x31 & ~x33 & ~x35 & ~x48 & ~x52 & ~x53 & ~x56 & ~x57 & ~x61 & ~x63 & ~x75 & ~x76 & ~x77 & ~x85 & ~x86 & ~x89 & ~x91 & ~x104 & ~x110 & ~x111 & ~x117 & ~x134 & ~x135 & ~x137 & ~x144 & ~x145 & ~x172 & ~x173 & ~x192 & ~x198 & ~x199 & ~x220 & ~x222 & ~x227 & ~x228 & ~x247 & ~x249 & ~x251 & ~x252 & ~x253 & ~x256 & ~x275 & ~x281 & ~x304 & ~x308 & ~x310 & ~x312 & ~x331 & ~x332 & ~x333 & ~x334 & ~x336 & ~x338 & ~x339 & ~x360 & ~x366 & ~x368 & ~x388 & ~x392 & ~x393 & ~x396 & ~x416 & ~x417 & ~x419 & ~x423 & ~x424 & ~x446 & ~x447 & ~x449 & ~x450 & ~x452 & ~x472 & ~x473 & ~x477 & ~x478 & ~x479 & ~x480 & ~x502 & ~x503 & ~x506 & ~x507 & ~x529 & ~x532 & ~x533 & ~x536 & ~x558 & ~x559 & ~x560 & ~x561 & ~x587 & ~x588 & ~x589 & ~x590 & ~x613 & ~x615 & ~x617 & ~x618 & ~x619 & ~x640 & ~x643 & ~x673 & ~x675 & ~x699 & ~x758 & ~x775;
assign c2224 =  x76 &  x92 &  x146 &  x464 &  x705 & ~x27 & ~x29 & ~x85 & ~x109 & ~x110 & ~x112 & ~x138 & ~x141 & ~x165 & ~x166 & ~x169 & ~x364 & ~x391 & ~x419 & ~x447 & ~x449 & ~x474 & ~x478 & ~x505 & ~x559 & ~x588 & ~x645 & ~x673 & ~x699 & ~x701 & ~x763 & ~x782 & ~x783;
assign c2226 =  x750 & ~x3 & ~x58 & ~x88 & ~x111 & ~x112 & ~x114 & ~x116 & ~x138 & ~x169 & ~x172 & ~x196 & ~x221 & ~x224 & ~x226 & ~x255 & ~x307 & ~x310 & ~x334 & ~x335 & ~x361 & ~x419 & ~x447 & ~x448 & ~x449 & ~x474 & ~x475 & ~x479 & ~x506 & ~x533 & ~x558 & ~x563 & ~x586 & ~x587 & ~x589 & ~x613 & ~x643 & ~x647 & ~x651 & ~x701 & ~x743 & ~x744 & ~x747 & ~x755 & ~x758 & ~x763 & ~x773 & ~x783;
assign c2228 =  x686 &  x687 &  x690 &  x709 &  x710 &  x713 &  x714 &  x716 &  x762 & ~x21 & ~x30 & ~x60 & ~x80 & ~x86 & ~x88 & ~x111 & ~x166 & ~x167 & ~x193 & ~x198 & ~x225 & ~x447 & ~x450 & ~x505 & ~x557 & ~x591 & ~x641 & ~x643 & ~x669 & ~x672 & ~x697 & ~x699 & ~x702 & ~x767 & ~x770 & ~x782 & ~x783;
assign c2230 =  x36 & ~x30 & ~x85 & ~x309 & ~x726 & ~x737 & ~x739 & ~x740 & ~x741 & ~x744 & ~x757 & ~x769 & ~x772 & ~x774;
assign c2232 =  x263 & ~x30 & ~x52 & ~x108 & ~x278 & ~x280 & ~x307 & ~x361 & ~x390 & ~x478 & ~x568 & ~x698 & ~x699 & ~x726 & ~x746 & ~x767 & ~x772 & ~x773;
assign c2234 =  x441 &  x469 & ~x4 & ~x5 & ~x6 & ~x7 & ~x8 & ~x9 & ~x28 & ~x29 & ~x36 & ~x48 & ~x51 & ~x53 & ~x56 & ~x59 & ~x60 & ~x64 & ~x65 & ~x76 & ~x78 & ~x79 & ~x86 & ~x92 & ~x104 & ~x110 & ~x116 & ~x138 & ~x139 & ~x142 & ~x144 & ~x170 & ~x193 & ~x198 & ~x219 & ~x220 & ~x222 & ~x223 & ~x224 & ~x225 & ~x248 & ~x249 & ~x253 & ~x254 & ~x255 & ~x276 & ~x277 & ~x282 & ~x304 & ~x310 & ~x332 & ~x334 & ~x336 & ~x339 & ~x361 & ~x388 & ~x389 & ~x390 & ~x391 & ~x393 & ~x395 & ~x396 & ~x420 & ~x421 & ~x422 & ~x423 & ~x446 & ~x447 & ~x448 & ~x449 & ~x450 & ~x451 & ~x472 & ~x473 & ~x478 & ~x502 & ~x528 & ~x530 & ~x532 & ~x534 & ~x561 & ~x563 & ~x587 & ~x615 & ~x617 & ~x618 & ~x643 & ~x645 & ~x670 & ~x671 & ~x673 & ~x699 & ~x700 & ~x728 & ~x731 & ~x754 & ~x758 & ~x760 & ~x780 & ~x783;
assign c2236 =  x94 &  x349 &  x407 &  x575 &  x576 &  x630 &  x631 &  x655 & ~x2 & ~x4 & ~x8 & ~x23 & ~x24 & ~x31 & ~x35 & ~x49 & ~x50 & ~x53 & ~x55 & ~x57 & ~x59 & ~x60 & ~x79 & ~x80 & ~x81 & ~x83 & ~x110 & ~x115 & ~x135 & ~x136 & ~x138 & ~x140 & ~x143 & ~x144 & ~x163 & ~x164 & ~x167 & ~x169 & ~x171 & ~x172 & ~x193 & ~x194 & ~x197 & ~x198 & ~x224 & ~x225 & ~x227 & ~x248 & ~x250 & ~x251 & ~x252 & ~x278 & ~x279 & ~x304 & ~x306 & ~x307 & ~x309 & ~x310 & ~x333 & ~x335 & ~x337 & ~x360 & ~x361 & ~x362 & ~x364 & ~x366 & ~x388 & ~x389 & ~x390 & ~x392 & ~x394 & ~x395 & ~x416 & ~x417 & ~x422 & ~x444 & ~x446 & ~x449 & ~x450 & ~x451 & ~x472 & ~x473 & ~x474 & ~x475 & ~x479 & ~x505 & ~x507 & ~x528 & ~x531 & ~x559 & ~x585 & ~x588 & ~x613 & ~x617 & ~x618 & ~x643 & ~x645 & ~x669 & ~x671 & ~x673 & ~x701 & ~x726 & ~x729 & ~x738 & ~x740 & ~x741 & ~x742 & ~x743 & ~x744 & ~x745 & ~x757 & ~x764 & ~x765 & ~x766 & ~x767 & ~x768 & ~x769 & ~x770 & ~x771 & ~x773 & ~x774 & ~x780 & ~x781 & ~x782;
assign c2238 =  x116;
assign c2240 =  x44 &  x45 &  x70 &  x594 &  x622 & ~x0 & ~x1 & ~x3 & ~x5 & ~x7 & ~x21 & ~x23 & ~x24 & ~x26 & ~x27 & ~x29 & ~x33 & ~x34 & ~x50 & ~x53 & ~x55 & ~x58 & ~x59 & ~x61 & ~x78 & ~x79 & ~x81 & ~x83 & ~x86 & ~x87 & ~x89 & ~x110 & ~x111 & ~x116 & ~x136 & ~x139 & ~x140 & ~x141 & ~x165 & ~x166 & ~x167 & ~x168 & ~x169 & ~x171 & ~x194 & ~x195 & ~x221 & ~x223 & ~x225 & ~x227 & ~x251 & ~x253 & ~x281 & ~x282 & ~x308 & ~x309 & ~x311 & ~x334 & ~x337 & ~x338 & ~x339 & ~x361 & ~x362 & ~x364 & ~x366 & ~x392 & ~x394 & ~x395 & ~x417 & ~x421 & ~x446 & ~x447 & ~x449 & ~x474 & ~x476 & ~x502 & ~x503 & ~x504 & ~x506 & ~x531 & ~x534 & ~x558 & ~x561 & ~x562 & ~x586 & ~x590 & ~x614 & ~x615 & ~x617 & ~x618 & ~x642 & ~x643 & ~x644 & ~x646 & ~x671 & ~x672 & ~x673 & ~x674 & ~x698 & ~x700 & ~x701 & ~x702 & ~x727 & ~x754 & ~x755 & ~x759 & ~x783;
assign c2242 =  x449;
assign c2244 =  x609 & ~x4 & ~x6 & ~x7 & ~x19 & ~x24 & ~x26 & ~x27 & ~x34 & ~x35 & ~x48 & ~x49 & ~x59 & ~x77 & ~x78 & ~x85 & ~x87 & ~x88 & ~x143 & ~x167 & ~x193 & ~x196 & ~x200 & ~x221 & ~x227 & ~x249 & ~x250 & ~x251 & ~x254 & ~x275 & ~x303 & ~x304 & ~x308 & ~x309 & ~x310 & ~x332 & ~x361 & ~x363 & ~x387 & ~x388 & ~x417 & ~x418 & ~x423 & ~x447 & ~x448 & ~x450 & ~x471 & ~x475 & ~x477 & ~x480 & ~x532 & ~x534 & ~x556 & ~x557 & ~x559 & ~x562 & ~x583 & ~x584 & ~x589 & ~x612 & ~x615 & ~x620 & ~x639 & ~x640 & ~x648 & ~x675 & ~x696 & ~x703 & ~x723;
assign c2246 =  x131 &  x330 &  x467 & ~x4 & ~x9 & ~x10 & ~x14 & ~x15 & ~x30 & ~x58 & ~x60 & ~x78 & ~x84 & ~x86 & ~x107 & ~x138 & ~x142 & ~x169 & ~x227 & ~x254 & ~x310 & ~x337 & ~x362 & ~x390 & ~x419 & ~x421;
assign c2248 =  x38 &  x444;
assign c2252 =  x66 &  x150 &  x383 &  x453 & ~x15 & ~x20 & ~x30 & ~x34 & ~x49 & ~x78 & ~x88 & ~x110 & ~x111 & ~x143 & ~x168 & ~x196 & ~x223 & ~x337 & ~x338 & ~x366 & ~x390 & ~x447 & ~x644 & ~x782;
assign c2254 =  x63 &  x117 &  x256 &  x312 & ~x27 & ~x31 & ~x52 & ~x53 & ~x55 & ~x110 & ~x141 & ~x420;
assign c2256 = ~x1 & ~x3 & ~x4 & ~x21 & ~x25 & ~x26 & ~x52 & ~x57 & ~x82 & ~x83 & ~x85 & ~x109 & ~x111 & ~x141 & ~x143 & ~x164 & ~x166 & ~x167 & ~x223 & ~x225 & ~x227 & ~x283 & ~x305 & ~x306 & ~x334 & ~x364 & ~x390 & ~x391 & ~x392 & ~x412 & ~x417 & ~x473 & ~x476 & ~x477 & ~x478 & ~x502 & ~x505 & ~x530 & ~x531 & ~x532 & ~x558 & ~x585 & ~x590 & ~x614 & ~x616 & ~x670 & ~x671 & ~x673 & ~x698 & ~x700 & ~x739 & ~x740 & ~x743 & ~x744 & ~x745 & ~x746 & ~x755 & ~x757 & ~x758 & ~x765 & ~x766 & ~x772 & ~x773 & ~x776;
assign c2258 =  x46 &  x73 &  x133 &  x174 &  x593 &  x715 &  x716 & ~x23 & ~x142 & ~x167;
assign c2260 =  x329 &  x436 & ~x5 & ~x6 & ~x55 & ~x60 & ~x113 & ~x222 & ~x282 & ~x306 & ~x311 & ~x445 & ~x502 & ~x528 & ~x558 & ~x614 & ~x615 & ~x641 & ~x644 & ~x645 & ~x664 & ~x700 & ~x702 & ~x773;
assign c2262 = ~x23 & ~x24 & ~x28 & ~x56 & ~x58 & ~x80 & ~x84 & ~x85 & ~x112 & ~x114 & ~x141 & ~x166 & ~x170 & ~x171 & ~x172 & ~x195 & ~x197 & ~x225 & ~x248 & ~x276 & ~x277 & ~x278 & ~x283 & ~x304 & ~x305 & ~x332 & ~x334 & ~x336 & ~x337 & ~x350 & ~x361 & ~x365 & ~x389 & ~x390 & ~x395 & ~x416 & ~x418 & ~x421 & ~x445 & ~x446 & ~x449 & ~x451 & ~x472 & ~x475 & ~x500 & ~x501 & ~x502 & ~x503 & ~x504 & ~x530 & ~x533 & ~x558 & ~x584 & ~x586 & ~x588 & ~x591 & ~x644 & ~x672 & ~x697 & ~x724 & ~x726 & ~x728 & ~x756 & ~x757 & ~x765 & ~x766 & ~x767 & ~x768 & ~x769 & ~x770 & ~x771 & ~x773 & ~x775;
assign c2264 =  x144 &  x479 &  x480 & ~x28;
assign c2266 =  x174 &  x202 &  x205 &  x402 &  x414 &  x425 &  x464 &  x518 & ~x6 & ~x15 & ~x22 & ~x57 & ~x60 & ~x80 & ~x89 & ~x107 & ~x114 & ~x166 & ~x193 & ~x200 & ~x308 & ~x309 & ~x361 & ~x390 & ~x588 & ~x615 & ~x699;
assign c2268 =  x60;
assign c2270 =  x320 & ~x79 & ~x197 & ~x283 & ~x361 & ~x640 & ~x683 & ~x688 & ~x765;
assign c2272 =  x10 &  x667 & ~x28 & ~x82 & ~x83 & ~x112 & ~x114 & ~x141;
assign c2274 =  x38 &  x39 &  x45 &  x94 &  x272 &  x317 &  x375 &  x384 &  x403 &  x405 &  x460 &  x490 &  x513 &  x515 &  x516 & ~x0 & ~x1 & ~x2 & ~x6 & ~x22 & ~x26 & ~x28 & ~x29 & ~x30 & ~x33 & ~x34 & ~x52 & ~x54 & ~x56 & ~x58 & ~x59 & ~x61 & ~x79 & ~x82 & ~x83 & ~x107 & ~x108 & ~x109 & ~x110 & ~x112 & ~x113 & ~x114 & ~x115 & ~x116 & ~x137 & ~x139 & ~x140 & ~x144 & ~x164 & ~x165 & ~x167 & ~x171 & ~x192 & ~x195 & ~x199 & ~x221 & ~x222 & ~x225 & ~x226 & ~x248 & ~x250 & ~x252 & ~x253 & ~x276 & ~x282 & ~x305 & ~x306 & ~x307 & ~x310 & ~x311 & ~x333 & ~x336 & ~x337 & ~x360 & ~x361 & ~x362 & ~x390 & ~x393 & ~x417 & ~x418 & ~x419 & ~x422 & ~x446 & ~x447 & ~x449 & ~x450 & ~x451 & ~x475 & ~x478 & ~x479 & ~x505 & ~x507 & ~x531 & ~x534 & ~x558 & ~x560 & ~x561 & ~x562 & ~x585 & ~x586 & ~x587 & ~x589 & ~x590 & ~x616 & ~x641 & ~x672 & ~x697 & ~x707 & ~x725 & ~x726 & ~x753 & ~x763 & ~x781;
assign c2276 =  x348 &  x455 &  x609 &  x665 & ~x49 & ~x79 & ~x135 & ~x172 & ~x419 & ~x639 & ~x669;
assign c2278 =  x356 &  x434 &  x435 &  x546 & ~x34 & ~x83 & ~x138 & ~x275 & ~x303 & ~x452 & ~x611 & ~x670 & ~x759 & ~x780;
assign c2280 = ~x2 & ~x3 & ~x5 & ~x7 & ~x21 & ~x22 & ~x23 & ~x25 & ~x26 & ~x29 & ~x31 & ~x32 & ~x34 & ~x50 & ~x51 & ~x53 & ~x55 & ~x58 & ~x61 & ~x78 & ~x82 & ~x85 & ~x108 & ~x109 & ~x137 & ~x141 & ~x165 & ~x167 & ~x169 & ~x170 & ~x171 & ~x172 & ~x196 & ~x198 & ~x200 & ~x220 & ~x221 & ~x222 & ~x225 & ~x227 & ~x247 & ~x248 & ~x249 & ~x253 & ~x255 & ~x256 & ~x278 & ~x279 & ~x280 & ~x281 & ~x282 & ~x283 & ~x309 & ~x332 & ~x334 & ~x337 & ~x365 & ~x366 & ~x367 & ~x389 & ~x393 & ~x394 & ~x417 & ~x419 & ~x450 & ~x451 & ~x473 & ~x479 & ~x500 & ~x502 & ~x504 & ~x505 & ~x506 & ~x529 & ~x530 & ~x531 & ~x534 & ~x535 & ~x557 & ~x560 & ~x584 & ~x585 & ~x586 & ~x589 & ~x590 & ~x612 & ~x613 & ~x614 & ~x615 & ~x616 & ~x618 & ~x619 & ~x643 & ~x645 & ~x646 & ~x647 & ~x671 & ~x682 & ~x684 & ~x685 & ~x688 & ~x689 & ~x691 & ~x699 & ~x716 & ~x727 & ~x731 & ~x738 & ~x739 & ~x740 & ~x741 & ~x746 & ~x754 & ~x756 & ~x758 & ~x760 & ~x767 & ~x769 & ~x772 & ~x773;
assign c2282 = ~x0 & ~x3 & ~x5 & ~x22 & ~x25 & ~x28 & ~x30 & ~x31 & ~x33 & ~x61 & ~x76 & ~x80 & ~x105 & ~x133 & ~x138 & ~x144 & ~x193 & ~x220 & ~x256 & ~x276 & ~x279 & ~x280 & ~x281 & ~x332 & ~x335 & ~x338 & ~x339 & ~x354 & ~x366 & ~x410 & ~x417 & ~x438 & ~x447 & ~x448 & ~x449 & ~x474 & ~x476 & ~x500 & ~x505 & ~x507 & ~x558 & ~x699 & ~x700 & ~x781;
assign c2284 =  x245 &  x341 &  x369 &  x485 &  x521 &  x541 &  x544 &  x653 &  x733 & ~x86 & ~x88 & ~x114 & ~x249 & ~x281 & ~x309 & ~x337 & ~x395 & ~x531 & ~x562 & ~x644 & ~x651 & ~x701 & ~x730;
assign c2286 =  x721 & ~x1 & ~x3 & ~x4 & ~x6 & ~x7 & ~x9 & ~x18 & ~x24 & ~x27 & ~x28 & ~x31 & ~x32 & ~x34 & ~x35 & ~x51 & ~x55 & ~x58 & ~x59 & ~x61 & ~x63 & ~x64 & ~x79 & ~x80 & ~x81 & ~x84 & ~x85 & ~x87 & ~x88 & ~x89 & ~x108 & ~x109 & ~x110 & ~x111 & ~x113 & ~x115 & ~x136 & ~x140 & ~x141 & ~x143 & ~x167 & ~x168 & ~x170 & ~x171 & ~x191 & ~x192 & ~x194 & ~x195 & ~x196 & ~x198 & ~x199 & ~x200 & ~x223 & ~x225 & ~x228 & ~x249 & ~x250 & ~x251 & ~x253 & ~x256 & ~x278 & ~x303 & ~x305 & ~x307 & ~x308 & ~x309 & ~x311 & ~x332 & ~x333 & ~x334 & ~x335 & ~x336 & ~x360 & ~x362 & ~x363 & ~x365 & ~x388 & ~x389 & ~x391 & ~x395 & ~x417 & ~x418 & ~x422 & ~x424 & ~x443 & ~x444 & ~x446 & ~x448 & ~x449 & ~x451 & ~x452 & ~x472 & ~x473 & ~x475 & ~x476 & ~x477 & ~x479 & ~x501 & ~x502 & ~x504 & ~x505 & ~x507 & ~x508 & ~x529 & ~x531 & ~x558 & ~x561 & ~x562 & ~x583 & ~x585 & ~x586 & ~x614 & ~x616 & ~x618 & ~x619 & ~x644 & ~x646 & ~x669 & ~x670 & ~x671 & ~x672 & ~x675 & ~x698 & ~x699 & ~x701 & ~x702 & ~x725 & ~x727 & ~x728 & ~x729 & ~x753 & ~x756 & ~x757 & ~x759 & ~x767 & ~x768 & ~x772 & ~x775 & ~x779 & ~x780 & ~x782;
assign c2288 = ~x97 & ~x347 & ~x393 & ~x474 & ~x735;
assign c2290 =  x15 &  x94 &  x160 &  x269 &  x371 &  x470 &  x654 &  x655 &  x691 &  x706 &  x734 & ~x2 & ~x3 & ~x4 & ~x6 & ~x20 & ~x29 & ~x30 & ~x32 & ~x49 & ~x50 & ~x54 & ~x55 & ~x56 & ~x59 & ~x78 & ~x81 & ~x83 & ~x86 & ~x87 & ~x88 & ~x108 & ~x111 & ~x116 & ~x143 & ~x164 & ~x167 & ~x168 & ~x169 & ~x192 & ~x199 & ~x223 & ~x224 & ~x250 & ~x252 & ~x254 & ~x277 & ~x280 & ~x305 & ~x307 & ~x309 & ~x310 & ~x311 & ~x335 & ~x362 & ~x363 & ~x365 & ~x367 & ~x393 & ~x420 & ~x421 & ~x423 & ~x446 & ~x451 & ~x473 & ~x474 & ~x506 & ~x507 & ~x529 & ~x533 & ~x534 & ~x535 & ~x559 & ~x561 & ~x586 & ~x590 & ~x591 & ~x614 & ~x616 & ~x644 & ~x647 & ~x670 & ~x671 & ~x672 & ~x673 & ~x698 & ~x703 & ~x726 & ~x729 & ~x730 & ~x731 & ~x756 & ~x759 & ~x766 & ~x767 & ~x771 & ~x772 & ~x774 & ~x775 & ~x783;
assign c2292 =  x172 &  x647;
assign c2294 =  x450;
assign c2296 =  x204 &  x262 &  x272 &  x458 &  x512 &  x575 &  x603 & ~x5 & ~x9 & ~x12 & ~x13 & ~x21 & ~x24 & ~x25 & ~x26 & ~x29 & ~x30 & ~x31 & ~x54 & ~x83 & ~x86 & ~x88 & ~x111 & ~x116 & ~x135 & ~x139 & ~x164 & ~x166 & ~x194 & ~x198 & ~x221 & ~x222 & ~x227 & ~x250 & ~x251 & ~x252 & ~x253 & ~x306 & ~x308 & ~x310 & ~x334 & ~x361 & ~x363 & ~x390 & ~x448 & ~x757 & ~x782;
assign c2298 = ~x1 & ~x4 & ~x5 & ~x7 & ~x20 & ~x31 & ~x32 & ~x48 & ~x49 & ~x51 & ~x52 & ~x53 & ~x55 & ~x58 & ~x59 & ~x61 & ~x76 & ~x78 & ~x82 & ~x83 & ~x84 & ~x107 & ~x108 & ~x110 & ~x113 & ~x114 & ~x115 & ~x116 & ~x143 & ~x164 & ~x167 & ~x168 & ~x171 & ~x195 & ~x197 & ~x200 & ~x221 & ~x226 & ~x227 & ~x228 & ~x248 & ~x253 & ~x281 & ~x306 & ~x307 & ~x309 & ~x310 & ~x332 & ~x334 & ~x362 & ~x390 & ~x391 & ~x394 & ~x395 & ~x418 & ~x419 & ~x420 & ~x421 & ~x423 & ~x446 & ~x447 & ~x448 & ~x450 & ~x473 & ~x475 & ~x476 & ~x477 & ~x479 & ~x503 & ~x504 & ~x506 & ~x507 & ~x513 & ~x530 & ~x533 & ~x535 & ~x587 & ~x588 & ~x589 & ~x619 & ~x641 & ~x644 & ~x669 & ~x672 & ~x698 & ~x699 & ~x701 & ~x728 & ~x730 & ~x760 & ~x781 & ~x782;
assign c2300 =  x289 & ~x167 & ~x195 & ~x215 & ~x227 & ~x334 & ~x364 & ~x392 & ~x393 & ~x417 & ~x445 & ~x477 & ~x502 & ~x558 & ~x616 & ~x641 & ~x674 & ~x725 & ~x776;
assign c2302 =  x44 &  x70 &  x413 &  x489 &  x683 &  x746 &  x750 & ~x62 & ~x91 & ~x105 & ~x278 & ~x281 & ~x473 & ~x613 & ~x730 & ~x760;
assign c2304 =  x17 &  x553 & ~x449 & ~x528 & ~x780;
assign c2306 = ~x2 & ~x6 & ~x22 & ~x52 & ~x53 & ~x58 & ~x59 & ~x60 & ~x85 & ~x87 & ~x109 & ~x140 & ~x142 & ~x143 & ~x153 & ~x155 & ~x165 & ~x167 & ~x168 & ~x169 & ~x170 & ~x171 & ~x172 & ~x192 & ~x195 & ~x220 & ~x247 & ~x249 & ~x250 & ~x277 & ~x282 & ~x283 & ~x306 & ~x332 & ~x334 & ~x336 & ~x337 & ~x338 & ~x339 & ~x361 & ~x362 & ~x363 & ~x390 & ~x394 & ~x423 & ~x445 & ~x446 & ~x449 & ~x473 & ~x502 & ~x503 & ~x504 & ~x530 & ~x534 & ~x557 & ~x560 & ~x585 & ~x589 & ~x590 & ~x614 & ~x615 & ~x641 & ~x645 & ~x669 & ~x670 & ~x698 & ~x699 & ~x700 & ~x726 & ~x756 & ~x757 & ~x758 & ~x764 & ~x766 & ~x767 & ~x768 & ~x769 & ~x770 & ~x775 & ~x783;
assign c2308 =  x89 &  x386 & ~x0 & ~x24 & ~x26 & ~x32 & ~x52 & ~x54 & ~x55 & ~x82 & ~x83 & ~x86 & ~x109 & ~x308 & ~x531 & ~x729 & ~x756;
assign c2310 =  x636 & ~x103 & ~x118 & ~x361 & ~x363 & ~x611 & ~x675;
assign c2312 = ~x4 & ~x5 & ~x6 & ~x24 & ~x31 & ~x51 & ~x52 & ~x55 & ~x56 & ~x58 & ~x61 & ~x81 & ~x83 & ~x107 & ~x108 & ~x135 & ~x136 & ~x138 & ~x144 & ~x165 & ~x167 & ~x171 & ~x193 & ~x194 & ~x196 & ~x198 & ~x219 & ~x221 & ~x222 & ~x223 & ~x224 & ~x226 & ~x227 & ~x246 & ~x249 & ~x250 & ~x252 & ~x253 & ~x255 & ~x274 & ~x277 & ~x278 & ~x279 & ~x280 & ~x304 & ~x305 & ~x306 & ~x309 & ~x310 & ~x332 & ~x333 & ~x334 & ~x335 & ~x338 & ~x339 & ~x360 & ~x361 & ~x362 & ~x364 & ~x389 & ~x390 & ~x392 & ~x393 & ~x417 & ~x418 & ~x419 & ~x421 & ~x448 & ~x449 & ~x474 & ~x477 & ~x479 & ~x500 & ~x501 & ~x506 & ~x507 & ~x527 & ~x528 & ~x532 & ~x556 & ~x584 & ~x587 & ~x615 & ~x617 & ~x643 & ~x644 & ~x645 & ~x646 & ~x670 & ~x672 & ~x696 & ~x698 & ~x701 & ~x726 & ~x727 & ~x740 & ~x741 & ~x742 & ~x744 & ~x745 & ~x768 & ~x769 & ~x772 & ~x773 & ~x783;
assign c2314 =  x44 &  x70 &  x567 &  x595 &  x609 &  x693 &  x711 &  x716 &  x741 &  x742 &  x743 & ~x6 & ~x21 & ~x24 & ~x28 & ~x31 & ~x54 & ~x61 & ~x111 & ~x220 & ~x221 & ~x224 & ~x388 & ~x418 & ~x419 & ~x420 & ~x446 & ~x449 & ~x473 & ~x474 & ~x501 & ~x529 & ~x589 & ~x640 & ~x703;
assign c2316 =  x75 &  x300 &  x329 &  x435 &  x465 &  x482 &  x545 & ~x1 & ~x14 & ~x199 & ~x249 & ~x307 & ~x558 & ~x586 & ~x590 & ~x646 & ~x671 & ~x702 & ~x756;
assign c2318 =  x300 &  x356 &  x497 &  x511 &  x693 &  x721 &  x749 &  x777 & ~x0 & ~x2 & ~x3 & ~x4 & ~x5 & ~x6 & ~x7 & ~x22 & ~x23 & ~x25 & ~x28 & ~x31 & ~x34 & ~x48 & ~x51 & ~x52 & ~x53 & ~x55 & ~x57 & ~x58 & ~x59 & ~x60 & ~x78 & ~x79 & ~x80 & ~x81 & ~x82 & ~x88 & ~x106 & ~x107 & ~x108 & ~x109 & ~x110 & ~x111 & ~x112 & ~x136 & ~x137 & ~x138 & ~x140 & ~x141 & ~x163 & ~x166 & ~x167 & ~x168 & ~x170 & ~x171 & ~x172 & ~x194 & ~x195 & ~x197 & ~x198 & ~x199 & ~x220 & ~x227 & ~x228 & ~x247 & ~x248 & ~x249 & ~x251 & ~x254 & ~x275 & ~x277 & ~x279 & ~x281 & ~x282 & ~x283 & ~x284 & ~x303 & ~x304 & ~x305 & ~x306 & ~x307 & ~x308 & ~x309 & ~x332 & ~x333 & ~x334 & ~x336 & ~x338 & ~x339 & ~x360 & ~x363 & ~x366 & ~x388 & ~x389 & ~x390 & ~x391 & ~x393 & ~x395 & ~x419 & ~x421 & ~x422 & ~x423 & ~x447 & ~x448 & ~x449 & ~x473 & ~x476 & ~x478 & ~x479 & ~x501 & ~x502 & ~x503 & ~x507 & ~x534 & ~x561 & ~x562 & ~x585 & ~x587 & ~x589 & ~x590 & ~x613 & ~x619 & ~x642 & ~x644 & ~x669 & ~x672 & ~x673 & ~x674 & ~x699 & ~x700 & ~x701 & ~x726 & ~x727 & ~x753 & ~x754 & ~x755 & ~x757 & ~x765 & ~x767 & ~x768 & ~x770 & ~x774 & ~x781;
assign c2320 =  x751 & ~x4 & ~x22 & ~x31 & ~x32 & ~x55 & ~x58 & ~x79 & ~x83 & ~x85 & ~x86 & ~x110 & ~x115 & ~x141 & ~x166 & ~x167 & ~x195 & ~x198 & ~x224 & ~x225 & ~x253 & ~x310 & ~x334 & ~x364 & ~x366 & ~x391 & ~x419 & ~x447 & ~x506 & ~x530 & ~x531 & ~x533 & ~x558 & ~x567 & ~x586 & ~x617 & ~x644 & ~x674 & ~x728 & ~x755 & ~x764 & ~x766 & ~x767 & ~x770 & ~x776;
assign c2322 = ~x1 & ~x3 & ~x22 & ~x24 & ~x25 & ~x27 & ~x33 & ~x82 & ~x125 & ~x138 & ~x252 & ~x277 & ~x307 & ~x308 & ~x355 & ~x393 & ~x417 & ~x418 & ~x419 & ~x445 & ~x449 & ~x530 & ~x532 & ~x586 & ~x587 & ~x588 & ~x644 & ~x670 & ~x756 & ~x757 & ~x764;
assign c2324 =  x95 &  x122 &  x125 &  x158 &  x176 &  x245 &  x263 &  x328 &  x402 &  x404 &  x413 &  x458 &  x482 &  x488 &  x525 &  x539 &  x553 &  x573 &  x574 &  x581 &  x609 &  x628 &  x637 &  x693 &  x721 &  x749 & ~x0 & ~x1 & ~x7 & ~x20 & ~x25 & ~x87 & ~x109 & ~x116 & ~x117 & ~x136 & ~x137 & ~x140 & ~x144 & ~x169 & ~x171 & ~x172 & ~x192 & ~x193 & ~x199 & ~x221 & ~x226 & ~x227 & ~x248 & ~x254 & ~x255 & ~x283 & ~x337 & ~x338 & ~x360 & ~x392 & ~x418 & ~x419 & ~x447 & ~x450 & ~x476 & ~x478 & ~x479 & ~x502 & ~x529 & ~x530 & ~x533 & ~x535 & ~x562 & ~x586 & ~x587 & ~x588 & ~x613 & ~x619 & ~x640 & ~x673 & ~x675 & ~x697 & ~x699 & ~x701 & ~x730 & ~x758 & ~x780 & ~x783;
assign c2326 =  x641 &  x647;
assign c2328 =  x10 &  x16 &  x582 & ~x22 & ~x30 & ~x58 & ~x80 & ~x729;
assign c2330 =  x442 &  x498 & ~x2 & ~x24 & ~x26 & ~x28 & ~x31 & ~x55 & ~x58 & ~x85 & ~x113 & ~x115 & ~x142 & ~x223 & ~x250 & ~x251 & ~x280 & ~x281 & ~x307 & ~x308 & ~x337 & ~x389 & ~x392 & ~x394 & ~x446 & ~x450 & ~x475 & ~x503 & ~x531 & ~x637 & ~x644 & ~x670 & ~x672 & ~x727 & ~x755 & ~x758;
assign c2332 =  x596 & ~x22 & ~x56 & ~x142 & ~x164 & ~x222 & ~x223 & ~x253 & ~x417 & ~x427 & ~x754;
assign c2334 =  x95 &  x101 &  x103 &  x132 &  x217 &  x302 &  x330 &  x414 &  x433 &  x435 &  x462 &  x463 &  x470 &  x515 &  x518 &  x570 &  x598 &  x599 &  x603 &  x627 &  x657 &  x661 & ~x29 & ~x50 & ~x57 & ~x61 & ~x82 & ~x107 & ~x137 & ~x199 & ~x221 & ~x305 & ~x334 & ~x366 & ~x391 & ~x445 & ~x446 & ~x450 & ~x474 & ~x507 & ~x531 & ~x557 & ~x562 & ~x589 & ~x616 & ~x731 & ~x757;
assign c2336 =  x45 &  x273 &  x315 &  x426 &  x427 &  x492 &  x515 &  x746 &  x750 & ~x21 & ~x60 & ~x83 & ~x88 & ~x110 & ~x116 & ~x141 & ~x169 & ~x192 & ~x224 & ~x248 & ~x252 & ~x255 & ~x339 & ~x363 & ~x389 & ~x449 & ~x450 & ~x479 & ~x505 & ~x529 & ~x532 & ~x560 & ~x584 & ~x585 & ~x615 & ~x644 & ~x645 & ~x671 & ~x673 & ~x674 & ~x725 & ~x754 & ~x781;
assign c2338 =  x589;
assign c2340 =  x596 & ~x85 & ~x138 & ~x254 & ~x309 & ~x336 & ~x505 & ~x523 & ~x530 & ~x645;
assign c2342 =  x42 &  x44 &  x398 &  x594 &  x678 & ~x0 & ~x3 & ~x8 & ~x25 & ~x33 & ~x78 & ~x81 & ~x82 & ~x83 & ~x116 & ~x138 & ~x144 & ~x172 & ~x303 & ~x305 & ~x336 & ~x393 & ~x395 & ~x420 & ~x450 & ~x452 & ~x472 & ~x476 & ~x501 & ~x528 & ~x562 & ~x586 & ~x700 & ~x702 & ~x704 & ~x730;
assign c2344 =  x16 & ~x0 & ~x7 & ~x24 & ~x25 & ~x49 & ~x59 & ~x84 & ~x87 & ~x88 & ~x113 & ~x136 & ~x137 & ~x141 & ~x142 & ~x144 & ~x163 & ~x195 & ~x219 & ~x220 & ~x222 & ~x226 & ~x253 & ~x255 & ~x278 & ~x305 & ~x311 & ~x333 & ~x363 & ~x365 & ~x387 & ~x391 & ~x416 & ~x417 & ~x503 & ~x529 & ~x531 & ~x560 & ~x562 & ~x613 & ~x645 & ~x698 & ~x725 & ~x753 & ~x755 & ~x767 & ~x768 & ~x773;
assign c2346 =  x395 & ~x447 & ~x756 & ~x762;
assign c2348 =  x37 &  x92 &  x101 &  x119 &  x189 &  x300 &  x408 &  x458 &  x554 &  x569 &  x593 & ~x21 & ~x61 & ~x83 & ~x115 & ~x116 & ~x169 & ~x250 & ~x590 & ~x642;
assign c2350 =  x652 & ~x84 & ~x86 & ~x638 & ~x762;
assign c2352 =  x721 & ~x656 & ~x657 & ~x659 & ~x662;
assign c2354 =  x38 &  x43 &  x257 &  x273 &  x411 &  x733 & ~x19 & ~x25 & ~x35 & ~x56 & ~x59 & ~x137 & ~x310 & ~x334 & ~x338 & ~x390 & ~x392 & ~x394 & ~x420 & ~x446 & ~x447 & ~x474 & ~x530 & ~x532 & ~x670 & ~x700 & ~x729 & ~x757;
assign c2356 =  x10 &  x554 &  x582 &  x610 & ~x1 & ~x3 & ~x7 & ~x20 & ~x23 & ~x27 & ~x50 & ~x53 & ~x54 & ~x56 & ~x57 & ~x60 & ~x83 & ~x84 & ~x85 & ~x111 & ~x112 & ~x138 & ~x167 & ~x169 & ~x171 & ~x193 & ~x196 & ~x198 & ~x221 & ~x224 & ~x249 & ~x250 & ~x277 & ~x280 & ~x281 & ~x305 & ~x306 & ~x333 & ~x339 & ~x361 & ~x362 & ~x363 & ~x366 & ~x389 & ~x417 & ~x420 & ~x474 & ~x506 & ~x531 & ~x533 & ~x558 & ~x560 & ~x590 & ~x616 & ~x699 & ~x701 & ~x754 & ~x755 & ~x757;
assign c2358 =  x477;
assign c2360 =  x43 &  x44 &  x665 & ~x19 & ~x20 & ~x22 & ~x24 & ~x53 & ~x55 & ~x106 & ~x169 & ~x170 & ~x226 & ~x278 & ~x281 & ~x340 & ~x476 & ~x564 & ~x617 & ~x618 & ~x620 & ~x671 & ~x723 & ~x752 & ~x760 & ~x783;
assign c2362 =  x75 &  x92 &  x133 &  x287 &  x302 &  x435 &  x582 & ~x1 & ~x5 & ~x13 & ~x28 & ~x30 & ~x61 & ~x87 & ~x109 & ~x110 & ~x111 & ~x166 & ~x169 & ~x252 & ~x474 & ~x476 & ~x560 & ~x728 & ~x730;
assign c2364 =  x469 & ~x1 & ~x29 & ~x30 & ~x52 & ~x123 & ~x124 & ~x126 & ~x127 & ~x220 & ~x227 & ~x304 & ~x311 & ~x335 & ~x389 & ~x421 & ~x445 & ~x446 & ~x447 & ~x473 & ~x501 & ~x533 & ~x613 & ~x618;
assign c2366 =  x38 &  x174 &  x218 &  x301 &  x498 & ~x3 & ~x21 & ~x30 & ~x53 & ~x54 & ~x79 & ~x83 & ~x86 & ~x137 & ~x139 & ~x196 & ~x197 & ~x224 & ~x250 & ~x251 & ~x307 & ~x308 & ~x334 & ~x337 & ~x339 & ~x395 & ~x530 & ~x531 & ~x556 & ~x559 & ~x585 & ~x589 & ~x590 & ~x641 & ~x643 & ~x670 & ~x701 & ~x759 & ~x782;
assign c2368 =  x506;
assign c2370 =  x96 &  x99 &  x148 &  x205 &  x244 &  x318 &  x329 &  x371 &  x382 &  x385 &  x407 &  x430 &  x437 &  x440 &  x441 &  x459 &  x486 &  x517 &  x546 &  x567 &  x594 &  x603 &  x706 &  x721 & ~x22 & ~x29 & ~x51 & ~x59 & ~x89 & ~x108 & ~x113 & ~x138 & ~x163 & ~x167 & ~x169 & ~x170 & ~x194 & ~x197 & ~x222 & ~x223 & ~x224 & ~x226 & ~x337 & ~x338 & ~x361 & ~x362 & ~x368 & ~x424 & ~x452 & ~x475 & ~x504 & ~x529 & ~x558 & ~x559 & ~x560 & ~x616 & ~x647 & ~x697 & ~x701 & ~x729 & ~x759;
assign c2372 =  x91 &  x92 &  x119 &  x161 &  x203 &  x273 &  x385 &  x434 &  x435 &  x485 &  x492 &  x515 &  x546 & ~x4 & ~x31 & ~x61 & ~x110 & ~x141 & ~x143 & ~x164 & ~x197 & ~x309 & ~x423 & ~x445 & ~x557 & ~x558 & ~x560 & ~x588 & ~x613 & ~x614 & ~x641 & ~x669 & ~x670 & ~x698 & ~x703 & ~x731 & ~x754 & ~x759;
assign c2374 =  x200 & ~x2 & ~x12 & ~x24 & ~x756;
assign c2376 = ~x4 & ~x5 & ~x6 & ~x25 & ~x29 & ~x55 & ~x57 & ~x59 & ~x80 & ~x108 & ~x110 & ~x111 & ~x137 & ~x138 & ~x140 & ~x141 & ~x143 & ~x164 & ~x166 & ~x167 & ~x168 & ~x169 & ~x170 & ~x171 & ~x195 & ~x196 & ~x221 & ~x225 & ~x226 & ~x250 & ~x253 & ~x254 & ~x276 & ~x278 & ~x308 & ~x334 & ~x335 & ~x362 & ~x365 & ~x384 & ~x390 & ~x391 & ~x392 & ~x393 & ~x417 & ~x418 & ~x420 & ~x421 & ~x448 & ~x473 & ~x475 & ~x476 & ~x477 & ~x504 & ~x531 & ~x532 & ~x533 & ~x558 & ~x560 & ~x585 & ~x615 & ~x616 & ~x617 & ~x644 & ~x645 & ~x673 & ~x701 & ~x702 & ~x727 & ~x739 & ~x740 & ~x741 & ~x744 & ~x754 & ~x755 & ~x756 & ~x758 & ~x759 & ~x767 & ~x768 & ~x769 & ~x772 & ~x773 & ~x775;
assign c2378 =  x10 &  x11 &  x426 & ~x7 & ~x24 & ~x28 & ~x56 & ~x111;
assign c2380 =  x325 &  x357 &  x413 &  x435 &  x525 &  x750 & ~x4 & ~x6 & ~x24 & ~x30 & ~x32 & ~x54 & ~x81 & ~x88 & ~x109 & ~x138 & ~x164 & ~x165 & ~x168 & ~x171 & ~x192 & ~x198 & ~x220 & ~x221 & ~x226 & ~x279 & ~x281 & ~x282 & ~x283 & ~x307 & ~x334 & ~x364 & ~x366 & ~x394 & ~x418 & ~x419 & ~x421 & ~x447 & ~x449 & ~x475 & ~x476 & ~x477 & ~x503 & ~x532 & ~x558 & ~x559 & ~x560 & ~x590 & ~x617 & ~x643 & ~x644 & ~x674 & ~x692 & ~x698 & ~x701 & ~x720 & ~x752 & ~x757 & ~x767 & ~x769 & ~x770 & ~x772 & ~x776 & ~x783;
assign c2382 =  x203 &  x343 &  x581 &  x609 & ~x50 & ~x85 & ~x87 & ~x115 & ~x134 & ~x140 & ~x196 & ~x253 & ~x282 & ~x338 & ~x669 & ~x695 & ~x704 & ~x751 & ~x752 & ~x753 & ~x755;
assign c2384 =  x43 &  x150 &  x152 &  x203 &  x314 &  x526 &  x553 &  x566 &  x594 &  x630 &  x655 &  x666 & ~x3 & ~x23 & ~x25 & ~x26 & ~x29 & ~x52 & ~x109 & ~x113 & ~x114 & ~x135 & ~x137 & ~x139 & ~x144 & ~x224 & ~x255 & ~x277 & ~x279 & ~x281 & ~x306 & ~x311 & ~x360 & ~x367 & ~x390 & ~x391 & ~x392 & ~x393 & ~x419 & ~x528 & ~x532 & ~x533 & ~x584 & ~x587 & ~x589 & ~x590 & ~x646 & ~x647 & ~x671 & ~x675 & ~x699 & ~x703 & ~x720 & ~x731 & ~x748 & ~x752 & ~x753 & ~x759 & ~x781 & ~x782 & ~x783;
assign c2386 =  x554 & ~x3 & ~x23 & ~x24 & ~x26 & ~x51 & ~x54 & ~x80 & ~x82 & ~x112 & ~x115 & ~x140 & ~x221 & ~x225 & ~x249 & ~x250 & ~x278 & ~x308 & ~x336 & ~x362 & ~x419 & ~x468 & ~x475 & ~x476 & ~x533 & ~x557 & ~x588 & ~x614 & ~x615 & ~x756 & ~x769 & ~x782;
assign c2388 =  x229 &  x438 &  x494 &  x600 &  x621 &  x629 &  x638 &  x751 & ~x5 & ~x7 & ~x22 & ~x30 & ~x53 & ~x58 & ~x81 & ~x107 & ~x110 & ~x111 & ~x136 & ~x140 & ~x141 & ~x164 & ~x167 & ~x198 & ~x220 & ~x221 & ~x226 & ~x250 & ~x278 & ~x283 & ~x311 & ~x335 & ~x339 & ~x389 & ~x393 & ~x394 & ~x395 & ~x422 & ~x451 & ~x504 & ~x505 & ~x506 & ~x507 & ~x535 & ~x560 & ~x590 & ~x614 & ~x616 & ~x618 & ~x643 & ~x672 & ~x697 & ~x701 & ~x730 & ~x752 & ~x753 & ~x754 & ~x764 & ~x776;
assign c2390 =  x47 &  x611 &  x638 & ~x3 & ~x21 & ~x30 & ~x33 & ~x57 & ~x109 & ~x110 & ~x166 & ~x197 & ~x251 & ~x278 & ~x336 & ~x363 & ~x391 & ~x421 & ~x448 & ~x473 & ~x476 & ~x478 & ~x529 & ~x531 & ~x533 & ~x585 & ~x725 & ~x726 & ~x730 & ~x783;
assign c2392 =  x95 &  x188 &  x454 &  x511 &  x574 &  x581 &  x622 &  x706 & ~x5 & ~x8 & ~x21 & ~x22 & ~x26 & ~x35 & ~x55 & ~x59 & ~x78 & ~x80 & ~x81 & ~x87 & ~x109 & ~x117 & ~x137 & ~x142 & ~x145 & ~x168 & ~x170 & ~x195 & ~x226 & ~x248 & ~x250 & ~x254 & ~x255 & ~x333 & ~x340 & ~x363 & ~x365 & ~x367 & ~x368 & ~x416 & ~x417 & ~x418 & ~x420 & ~x445 & ~x476 & ~x501 & ~x502 & ~x508 & ~x533 & ~x559 & ~x615 & ~x617 & ~x643 & ~x645 & ~x647 & ~x648 & ~x670 & ~x675 & ~x727 & ~x754 & ~x782;
assign c2394 =  x63 &  x90 &  x106 &  x471 & ~x2 & ~x6 & ~x27 & ~x57 & ~x81 & ~x138 & ~x169 & ~x196 & ~x308 & ~x363 & ~x391 & ~x476 & ~x503 & ~x756;
assign c2396 =  x366;
assign c2398 =  x394;
assign c2400 =  x507 &  x724;
assign c2402 =  x357 &  x385 &  x463 &  x489 &  x492 & ~x1 & ~x2 & ~x3 & ~x4 & ~x5 & ~x6 & ~x19 & ~x21 & ~x22 & ~x23 & ~x24 & ~x25 & ~x26 & ~x29 & ~x30 & ~x32 & ~x49 & ~x57 & ~x58 & ~x74 & ~x78 & ~x83 & ~x88 & ~x107 & ~x108 & ~x109 & ~x111 & ~x115 & ~x136 & ~x137 & ~x138 & ~x143 & ~x164 & ~x166 & ~x167 & ~x168 & ~x170 & ~x192 & ~x193 & ~x195 & ~x197 & ~x199 & ~x220 & ~x221 & ~x224 & ~x226 & ~x227 & ~x248 & ~x249 & ~x251 & ~x252 & ~x253 & ~x255 & ~x276 & ~x278 & ~x280 & ~x281 & ~x282 & ~x304 & ~x305 & ~x306 & ~x307 & ~x308 & ~x309 & ~x310 & ~x311 & ~x333 & ~x335 & ~x336 & ~x338 & ~x361 & ~x362 & ~x363 & ~x365 & ~x366 & ~x388 & ~x390 & ~x391 & ~x393 & ~x394 & ~x419 & ~x446 & ~x475 & ~x476 & ~x502 & ~x503 & ~x504 & ~x531 & ~x533 & ~x562 & ~x587 & ~x615 & ~x645 & ~x670 & ~x672 & ~x699 & ~x700 & ~x726 & ~x728 & ~x729 & ~x756 & ~x757 & ~x764 & ~x765 & ~x766 & ~x769 & ~x770 & ~x772 & ~x774 & ~x775 & ~x780 & ~x781 & ~x782 & ~x783;
assign c2404 =  x776;
assign c2406 =  x46 &  x148 &  x205 &  x216 &  x264 &  x314 &  x315 &  x519 &  x576 &  x600 &  x602 &  x603 &  x610 &  x657 &  x683 &  x711 &  x718 & ~x1 & ~x3 & ~x4 & ~x24 & ~x27 & ~x32 & ~x53 & ~x57 & ~x59 & ~x81 & ~x83 & ~x87 & ~x108 & ~x136 & ~x141 & ~x166 & ~x167 & ~x193 & ~x195 & ~x196 & ~x197 & ~x198 & ~x225 & ~x250 & ~x278 & ~x307 & ~x333 & ~x362 & ~x363 & ~x366 & ~x394 & ~x395 & ~x418 & ~x447 & ~x501 & ~x506 & ~x532 & ~x534 & ~x587 & ~x618 & ~x642 & ~x670 & ~x702 & ~x730 & ~x754 & ~x756 & ~x758 & ~x781 & ~x783;
assign c2408 =  x375 &  x403 &  x488 &  x596 & ~x7 & ~x12 & ~x13 & ~x32 & ~x80 & ~x81 & ~x110 & ~x171 & ~x227 & ~x255 & ~x282 & ~x307 & ~x310 & ~x363 & ~x390 & ~x476 & ~x477 & ~x505 & ~x618 & ~x644 & ~x670 & ~x671 & ~x701 & ~x749;
assign c2410 = ~x0 & ~x5 & ~x7 & ~x30 & ~x52 & ~x54 & ~x61 & ~x84 & ~x99 & ~x100 & ~x112 & ~x136 & ~x143 & ~x165 & ~x168 & ~x170 & ~x196 & ~x226 & ~x227 & ~x250 & ~x281 & ~x310 & ~x335 & ~x336 & ~x338 & ~x390 & ~x418 & ~x420 & ~x422 & ~x447 & ~x450 & ~x477 & ~x502 & ~x506 & ~x531 & ~x533 & ~x534 & ~x558 & ~x588 & ~x589 & ~x644 & ~x735 & ~x758 & ~x782;
assign c2412 = ~x1 & ~x22 & ~x26 & ~x50 & ~x51 & ~x53 & ~x59 & ~x61 & ~x78 & ~x79 & ~x80 & ~x82 & ~x83 & ~x138 & ~x139 & ~x150 & ~x153 & ~x154 & ~x164 & ~x166 & ~x169 & ~x171 & ~x193 & ~x194 & ~x196 & ~x222 & ~x223 & ~x227 & ~x248 & ~x249 & ~x252 & ~x254 & ~x276 & ~x279 & ~x280 & ~x281 & ~x283 & ~x304 & ~x305 & ~x308 & ~x332 & ~x361 & ~x364 & ~x367 & ~x388 & ~x390 & ~x395 & ~x417 & ~x420 & ~x445 & ~x446 & ~x449 & ~x472 & ~x473 & ~x503 & ~x505 & ~x530 & ~x557 & ~x558 & ~x560 & ~x585 & ~x588 & ~x613 & ~x669 & ~x699 & ~x728 & ~x729 & ~x743 & ~x757 & ~x767 & ~x768 & ~x769 & ~x771 & ~x773;
assign c2414 =  x113;
assign c2416 =  x46 &  x96 &  x119 &  x146 &  x217 &  x441 &  x489 &  x521 & ~x3 & ~x20 & ~x34 & ~x80 & ~x110 & ~x171 & ~x311 & ~x446 & ~x474 & ~x477 & ~x529 & ~x535 & ~x563 & ~x588 & ~x730;
assign c2418 = ~x0 & ~x26 & ~x32 & ~x50 & ~x54 & ~x56 & ~x79 & ~x84 & ~x86 & ~x87 & ~x111 & ~x125 & ~x137 & ~x142 & ~x168 & ~x187 & ~x191 & ~x196 & ~x219 & ~x227 & ~x248 & ~x252 & ~x276 & ~x278 & ~x304 & ~x305 & ~x336 & ~x378 & ~x388 & ~x448 & ~x476 & ~x530 & ~x547 & ~x558 & ~x615 & ~x616 & ~x669 & ~x702 & ~x759 & ~x767 & ~x782 & ~x783;
assign c2420 =  x314 & ~x84 & ~x186 & ~x505;
assign c2422 =  x157 &  x217 &  x246 &  x273 &  x287 &  x302 &  x379 &  x385 &  x509 &  x516 &  x544 &  x547 &  x574 &  x603 &  x649 &  x677 &  x685 &  x705 &  x712 &  x737 &  x743 &  x744 &  x747 & ~x25 & ~x29 & ~x51 & ~x56 & ~x57 & ~x167 & ~x224 & ~x252 & ~x477 & ~x531 & ~x643 & ~x672 & ~x729;
assign c2424 =  x46 &  x173 &  x258 &  x454 &  x467 &  x471 &  x541 &  x583 &  x639 & ~x5 & ~x7 & ~x52 & ~x193 & ~x194 & ~x195 & ~x222 & ~x252 & ~x615 & ~x730;
assign c2426 =  x612;
assign c2428 = ~x677 & ~x694;
assign c2430 =  x44 & ~x77 & ~x331 & ~x410 & ~x466;
assign c2432 =  x721 & ~x31 & ~x60 & ~x551 & ~x766 & ~x768 & ~x769;
assign c2434 =  x479 & ~x677;
assign c2436 =  x104 &  x122 &  x124 &  x125 &  x128 &  x131 &  x148 &  x154 &  x157 &  x160 &  x261 &  x269 &  x272 &  x291 &  x319 &  x347 &  x402 &  x431 &  x459 &  x460 &  x487 &  x488 &  x493 &  x516 &  x519 &  x520 &  x540 &  x542 &  x546 &  x573 &  x576 &  x577 &  x598 &  x599 &  x601 &  x603 &  x625 &  x630 &  x654 &  x657 & ~x0 & ~x28 & ~x80 & ~x107 & ~x113 & ~x167 & ~x168 & ~x195 & ~x221 & ~x224 & ~x248 & ~x249 & ~x279 & ~x280 & ~x283 & ~x311 & ~x338 & ~x360 & ~x366 & ~x389 & ~x446 & ~x448 & ~x449 & ~x473 & ~x505 & ~x507 & ~x528 & ~x532 & ~x562 & ~x586 & ~x612 & ~x616 & ~x640 & ~x642 & ~x643 & ~x647 & ~x696 & ~x699 & ~x703 & ~x782 & ~x783;
assign c2438 =  x325 &  x454 &  x488 &  x522 &  x548 &  x602 &  x657 &  x706 & ~x82 & ~x110 & ~x171 & ~x222 & ~x224 & ~x586 & ~x618 & ~x671 & ~x704 & ~x768 & ~x771;
assign c2440 =  x69 &  x403 &  x462 &  x493 &  x514 &  x572 &  x576 &  x626 &  x627 &  x779 & ~x32 & ~x83 & ~x114 & ~x136 & ~x142 & ~x168 & ~x195 & ~x249 & ~x305 & ~x306 & ~x361 & ~x362 & ~x367 & ~x422 & ~x450 & ~x474 & ~x477 & ~x503 & ~x558 & ~x560 & ~x586 & ~x618 & ~x674 & ~x700 & ~x728 & ~x730 & ~x754 & ~x777;
assign c2442 =  x149 &  x178 &  x202 &  x259 &  x443 &  x715 &  x724 & ~x52 & ~x448 & ~x503 & ~x588 & ~x756;
assign c2444 =  x401 &  x451;
assign c2446 =  x673;
assign c2448 =  x39 &  x68 &  x70 &  x258 &  x286 &  x374 &  x629 &  x762 & ~x33 & ~x61 & ~x112 & ~x192 & ~x284 & ~x534 & ~x586 & ~x703 & ~x725 & ~x757 & ~x766;
assign c2450 =  x96 &  x98 &  x158 &  x175 &  x188 &  x216 &  x273 &  x301 &  x436 &  x461 &  x464 &  x494 &  x554 &  x570 &  x573 &  x575 &  x582 &  x599 &  x604 &  x610 &  x626 &  x627 &  x629 & ~x1 & ~x23 & ~x25 & ~x27 & ~x54 & ~x57 & ~x86 & ~x89 & ~x114 & ~x115 & ~x167 & ~x195 & ~x199 & ~x223 & ~x227 & ~x247 & ~x251 & ~x303 & ~x310 & ~x418 & ~x445 & ~x479 & ~x502 & ~x503 & ~x530 & ~x531 & ~x563 & ~x640 & ~x670 & ~x748 & ~x752 & ~x755 & ~x756 & ~x758 & ~x783;
assign c2452 =  x17 &  x723 & ~x20 & ~x30 & ~x225 & ~x446 & ~x449 & ~x533 & ~x557;
assign c2454 =  x116 &  x367;
assign c2456 =  x64 &  x65 &  x611 & ~x14 & ~x60 & ~x61 & ~x114 & ~x193 & ~x195 & ~x306 & ~x390 & ~x671 & ~x672;
assign c2458 = ~x3 & ~x18 & ~x24 & ~x26 & ~x75 & ~x92 & ~x104 & ~x162 & ~x279 & ~x306 & ~x333 & ~x336 & ~x340 & ~x366 & ~x391 & ~x393 & ~x417 & ~x421 & ~x500 & ~x506 & ~x536 & ~x562 & ~x584 & ~x586 & ~x639 & ~x699 & ~x704 & ~x723 & ~x775;
assign c2460 =  x70 & ~x222 & ~x678;
assign c2462 = ~x300 & ~x436 & ~x467;
assign c2464 =  x426 & ~x433 & ~x434;
assign c2466 =  x45 &  x117 &  x342 &  x442 & ~x29 & ~x168;
assign c2468 =  x440 & ~x0 & ~x6 & ~x7 & ~x8 & ~x25 & ~x34 & ~x55 & ~x88 & ~x89 & ~x110 & ~x113 & ~x115 & ~x136 & ~x137 & ~x138 & ~x197 & ~x304 & ~x307 & ~x365 & ~x390 & ~x582 & ~x694 & ~x756;
assign c2470 =  x88;
assign c2472 =  x348 & ~x0 & ~x2 & ~x3 & ~x4 & ~x7 & ~x20 & ~x21 & ~x22 & ~x23 & ~x25 & ~x29 & ~x33 & ~x50 & ~x51 & ~x53 & ~x55 & ~x56 & ~x57 & ~x58 & ~x66 & ~x83 & ~x84 & ~x86 & ~x87 & ~x107 & ~x108 & ~x109 & ~x110 & ~x113 & ~x135 & ~x136 & ~x137 & ~x138 & ~x142 & ~x143 & ~x165 & ~x166 & ~x167 & ~x168 & ~x170 & ~x192 & ~x194 & ~x195 & ~x196 & ~x199 & ~x221 & ~x222 & ~x223 & ~x224 & ~x225 & ~x226 & ~x227 & ~x248 & ~x249 & ~x252 & ~x253 & ~x255 & ~x276 & ~x277 & ~x278 & ~x281 & ~x283 & ~x306 & ~x309 & ~x310 & ~x311 & ~x334 & ~x335 & ~x336 & ~x337 & ~x339 & ~x360 & ~x362 & ~x364 & ~x388 & ~x390 & ~x391 & ~x393 & ~x417 & ~x418 & ~x420 & ~x422 & ~x445 & ~x446 & ~x447 & ~x448 & ~x449 & ~x450 & ~x473 & ~x474 & ~x475 & ~x501 & ~x504 & ~x505 & ~x532 & ~x533 & ~x557 & ~x560 & ~x586 & ~x589 & ~x613 & ~x641 & ~x642 & ~x669 & ~x670 & ~x672 & ~x728 & ~x729 & ~x756 & ~x758 & ~x759 & ~x765 & ~x766 & ~x767 & ~x769 & ~x770 & ~x771 & ~x772 & ~x773 & ~x780 & ~x781;
assign c2474 =  x46 &  x368 &  x554 &  x582 & ~x3 & ~x32 & ~x52 & ~x82 & ~x111 & ~x306 & ~x308 & ~x310 & ~x333 & ~x337 & ~x338 & ~x361 & ~x391 & ~x417 & ~x418 & ~x447 & ~x476 & ~x506 & ~x558 & ~x646 & ~x701 & ~x730 & ~x782;
assign c2476 =  x37 &  x200 & ~x5 & ~x29 & ~x194 & ~x309;
assign c2478 = ~x1 & ~x6 & ~x21 & ~x28 & ~x30 & ~x32 & ~x35 & ~x52 & ~x55 & ~x81 & ~x85 & ~x89 & ~x105 & ~x107 & ~x108 & ~x111 & ~x141 & ~x143 & ~x144 & ~x166 & ~x170 & ~x173 & ~x192 & ~x200 & ~x224 & ~x226 & ~x247 & ~x249 & ~x253 & ~x255 & ~x275 & ~x276 & ~x279 & ~x281 & ~x283 & ~x306 & ~x307 & ~x308 & ~x311 & ~x312 & ~x334 & ~x337 & ~x339 & ~x341 & ~x360 & ~x361 & ~x362 & ~x364 & ~x390 & ~x391 & ~x392 & ~x396 & ~x416 & ~x417 & ~x419 & ~x420 & ~x421 & ~x423 & ~x444 & ~x445 & ~x449 & ~x450 & ~x472 & ~x473 & ~x474 & ~x477 & ~x478 & ~x500 & ~x501 & ~x502 & ~x530 & ~x531 & ~x532 & ~x534 & ~x558 & ~x589 & ~x619 & ~x643 & ~x644 & ~x697 & ~x698 & ~x701 & ~x702 & ~x703 & ~x727 & ~x730 & ~x739 & ~x741 & ~x742 & ~x744 & ~x745 & ~x755 & ~x757 & ~x765 & ~x767 & ~x768 & ~x773;
assign c2480 =  x63 & ~x5 & ~x28 & ~x82 & ~x251 & ~x391 & ~x420 & ~x447 & ~x448 & ~x558 & ~x614 & ~x743 & ~x744 & ~x756 & ~x768 & ~x776;
assign c2482 = ~x125 & ~x418 & ~x489 & ~x517 & ~x519 & ~x663;
assign c2484 =  x300 &  x545 &  x623 &  x721 & ~x4 & ~x25 & ~x35 & ~x49 & ~x78 & ~x173 & ~x248 & ~x282 & ~x304 & ~x334 & ~x447 & ~x559 & ~x616 & ~x674 & ~x675 & ~x676 & ~x700 & ~x703 & ~x766 & ~x782;
assign c2486 =  x725 & ~x694;
assign c2488 =  x98 &  x211 &  x261 &  x262 &  x298 &  x348 &  x373 &  x435 &  x463 &  x544 &  x548 &  x571 &  x577 &  x597 &  x598 &  x601 &  x628 &  x632 &  x656 &  x682 &  x717 &  x744 & ~x0 & ~x23 & ~x29 & ~x33 & ~x64 & ~x83 & ~x84 & ~x111 & ~x113 & ~x114 & ~x139 & ~x164 & ~x257 & ~x281 & ~x306 & ~x478 & ~x503 & ~x642 & ~x670 & ~x728 & ~x755 & ~x758;
assign c2490 =  x107;
assign c2492 = ~x4 & ~x53 & ~x85 & ~x111 & ~x167 & ~x169 & ~x222 & ~x251 & ~x490 & ~x492 & ~x493 & ~x550 & ~x558 & ~x644;
assign c2494 =  x685 & ~x5 & ~x25 & ~x28 & ~x29 & ~x32 & ~x54 & ~x55 & ~x79 & ~x82 & ~x87 & ~x136 & ~x140 & ~x142 & ~x163 & ~x226 & ~x250 & ~x256 & ~x280 & ~x306 & ~x307 & ~x308 & ~x309 & ~x360 & ~x362 & ~x363 & ~x364 & ~x390 & ~x391 & ~x392 & ~x393 & ~x421 & ~x445 & ~x446 & ~x476 & ~x532 & ~x557 & ~x559 & ~x560 & ~x562 & ~x586 & ~x589 & ~x616 & ~x637 & ~x644 & ~x665 & ~x693 & ~x699 & ~x728 & ~x756 & ~x757 & ~x782 & ~x783;
assign c2496 = ~x0 & ~x2 & ~x3 & ~x5 & ~x7 & ~x22 & ~x23 & ~x24 & ~x25 & ~x26 & ~x27 & ~x28 & ~x50 & ~x51 & ~x52 & ~x56 & ~x57 & ~x58 & ~x59 & ~x60 & ~x78 & ~x80 & ~x81 & ~x83 & ~x85 & ~x87 & ~x89 & ~x107 & ~x108 & ~x109 & ~x110 & ~x111 & ~x112 & ~x114 & ~x115 & ~x116 & ~x135 & ~x137 & ~x138 & ~x139 & ~x140 & ~x141 & ~x142 & ~x143 & ~x144 & ~x163 & ~x164 & ~x167 & ~x169 & ~x170 & ~x171 & ~x172 & ~x191 & ~x192 & ~x194 & ~x195 & ~x196 & ~x197 & ~x198 & ~x199 & ~x200 & ~x220 & ~x221 & ~x222 & ~x223 & ~x224 & ~x225 & ~x226 & ~x227 & ~x228 & ~x248 & ~x249 & ~x250 & ~x251 & ~x252 & ~x253 & ~x276 & ~x277 & ~x278 & ~x280 & ~x282 & ~x283 & ~x304 & ~x305 & ~x306 & ~x307 & ~x308 & ~x309 & ~x310 & ~x311 & ~x333 & ~x335 & ~x336 & ~x337 & ~x338 & ~x360 & ~x361 & ~x362 & ~x363 & ~x364 & ~x366 & ~x367 & ~x368 & ~x388 & ~x389 & ~x392 & ~x416 & ~x417 & ~x418 & ~x419 & ~x420 & ~x421 & ~x422 & ~x423 & ~x444 & ~x447 & ~x449 & ~x451 & ~x472 & ~x473 & ~x475 & ~x476 & ~x478 & ~x479 & ~x500 & ~x501 & ~x502 & ~x503 & ~x504 & ~x529 & ~x530 & ~x532 & ~x533 & ~x534 & ~x535 & ~x556 & ~x557 & ~x559 & ~x560 & ~x561 & ~x562 & ~x584 & ~x585 & ~x587 & ~x589 & ~x590 & ~x591 & ~x612 & ~x613 & ~x614 & ~x616 & ~x617 & ~x640 & ~x643 & ~x644 & ~x645 & ~x646 & ~x647 & ~x668 & ~x669 & ~x671 & ~x672 & ~x673 & ~x675 & ~x697 & ~x699 & ~x701 & ~x702 & ~x708 & ~x710 & ~x712 & ~x713 & ~x714 & ~x715 & ~x716 & ~x717 & ~x726 & ~x727 & ~x730 & ~x731 & ~x737 & ~x738 & ~x739 & ~x740 & ~x742 & ~x745 & ~x746 & ~x747 & ~x753 & ~x754 & ~x755 & ~x756 & ~x757 & ~x758 & ~x759 & ~x764 & ~x766 & ~x767 & ~x768 & ~x769 & ~x770 & ~x771 & ~x772 & ~x773 & ~x774 & ~x776 & ~x780 & ~x782;
assign c2498 = ~x23 & ~x86 & ~x87 & ~x91 & ~x104 & ~x107 & ~x112 & ~x113 & ~x140 & ~x198 & ~x200 & ~x222 & ~x224 & ~x249 & ~x251 & ~x253 & ~x282 & ~x306 & ~x308 & ~x309 & ~x311 & ~x336 & ~x365 & ~x366 & ~x367 & ~x420 & ~x449 & ~x450 & ~x464 & ~x473 & ~x477 & ~x503 & ~x518 & ~x519 & ~x530 & ~x533 & ~x586 & ~x587 & ~x618 & ~x645 & ~x728 & ~x754 & ~x757;
assign c21 =  x140;
assign c23 =  x80;
assign c27 =  x168;
assign c29 =  x278;
assign c211 =  x364;
assign c213 =  x4;
assign c215 =  x292 &  x294 &  x313 &  x315 &  x321 &  x322 &  x327 &  x348 &  x350 &  x369 &  x376 &  x379 &  x382 &  x397 &  x402 &  x405 &  x413 &  x425 &  x429 &  x438 &  x469 &  x481 &  x488 &  x490 &  x510 &  x520 &  x522 &  x525 &  x526 &  x536 &  x546 &  x552 &  x580 &  x595 &  x609 &  x625 &  x638 &  x704 &  x706 &  x734 & ~x22 & ~x27 & ~x28 & ~x31 & ~x32 & ~x83 & ~x89 & ~x107 & ~x135 & ~x168 & ~x171 & ~x198 & ~x222 & ~x251 & ~x253 & ~x503;
assign c217 =  x2 &  x392;
assign c219 =  x140;
assign c221 = ~x42 & ~x202;
assign c223 =  x167;
assign c225 =  x336;
assign c227 =  x109 &  x197;
assign c229 =  x142;
assign c231 = ~x17 & ~x152 & ~x208;
assign c233 = ~x359 & ~x450 & ~x590 & ~x593 & ~x609 & ~x639 & ~x640 & ~x696 & ~x702 & ~x705 & ~x706;
assign c235 =  x510 & ~x0 & ~x1 & ~x2 & ~x3 & ~x7 & ~x8 & ~x10 & ~x11 & ~x17 & ~x23 & ~x26 & ~x28 & ~x31 & ~x34 & ~x35 & ~x36 & ~x37 & ~x38 & ~x46 & ~x48 & ~x51 & ~x52 & ~x55 & ~x57 & ~x59 & ~x60 & ~x62 & ~x63 & ~x64 & ~x76 & ~x77 & ~x78 & ~x79 & ~x82 & ~x84 & ~x87 & ~x89 & ~x106 & ~x109 & ~x110 & ~x112 & ~x113 & ~x115 & ~x116 & ~x137 & ~x141 & ~x142 & ~x143 & ~x144 & ~x164 & ~x167 & ~x171 & ~x191 & ~x194 & ~x195 & ~x196 & ~x223 & ~x225 & ~x251 & ~x253 & ~x254 & ~x255 & ~x256 & ~x280 & ~x305 & ~x307 & ~x311 & ~x336 & ~x364 & ~x392 & ~x419 & ~x420 & ~x448 & ~x474 & ~x475 & ~x504 & ~x532 & ~x559 & ~x560 & ~x589 & ~x615 & ~x643 & ~x725 & ~x726 & ~x727 & ~x730 & ~x754 & ~x755 & ~x756 & ~x757 & ~x759 & ~x760 & ~x775 & ~x780 & ~x782 & ~x783;
assign c237 =  x52;
assign c239 =  x83;
assign c241 = ~x38 & ~x46 & ~x289;
assign c243 =  x165;
assign c245 =  x137;
assign c247 =  x64 & ~x28 & ~x335 & ~x341 & ~x394 & ~x414 & ~x499 & ~x500 & ~x555 & ~x584 & ~x725 & ~x730 & ~x751 & ~x781;
assign c249 =  x568 &  x636 &  x663 &  x707 &  x708 &  x709 &  x719 &  x745 & ~x475 & ~x620 & ~x644 & ~x699 & ~x753;
assign c251 =  x728;
assign c253 =  x307;
assign c255 =  x64 &  x94 &  x102 &  x179 &  x181 &  x234 &  x240 &  x243 &  x266 &  x271 &  x273 &  x297 &  x378 &  x491 &  x495 &  x580 &  x635 &  x653 &  x683 &  x712 &  x740 &  x744 & ~x4 & ~x6 & ~x52 & ~x140 & ~x194 & ~x279 & ~x447 & ~x614 & ~x725;
assign c257 =  x282;
assign c259 = ~x45 & ~x147;
assign c261 =  x251;
assign c263 =  x83;
assign c265 = ~x28 & ~x33 & ~x193 & ~x337 & ~x368 & ~x395 & ~x504 & ~x636 & ~x643 & ~x648 & ~x694 & ~x695 & ~x722 & ~x723 & ~x750 & ~x778;
assign c267 =  x3;
assign c269 = ~x371 & ~x426 & ~x480;
assign c271 =  x250;
assign c273 =  x363;
assign c275 =  x136;
assign c277 = ~x356 & ~x385 & ~x582;
assign c279 = ~x11 & ~x37 & ~x38;
assign c281 =  x167;
assign c283 =  x111;
assign c285 =  x21;
assign c287 =  x93 &  x103 &  x127 &  x237 &  x240 &  x273 &  x347 &  x457 &  x599 &  x606 &  x655 &  x657 &  x659 &  x661 &  x684 &  x688 &  x690 &  x715 &  x717 &  x740 &  x746 & ~x112 & ~x138 & ~x139 & ~x169 & ~x225 & ~x337 & ~x390 & ~x531 & ~x532 & ~x533 & ~x646 & ~x648 & ~x674 & ~x676 & ~x726 & ~x729 & ~x752 & ~x756 & ~x778;
assign c289 =  x139;
assign c291 =  x65 &  x521 &  x653 &  x718 & ~x251 & ~x415 & ~x451 & ~x479 & ~x557 & ~x614 & ~x778;
assign c293 =  x22;
assign c295 =  x139;
assign c297 =  x644;
assign c299 =  x250;
assign c2101 =  x86;
assign c2103 =  x393;
assign c2105 = ~x37 & ~x39 & ~x176 & ~x772;
assign c2107 = ~x1 & ~x10 & ~x11 & ~x38 & ~x46 & ~x87 & ~x711 & ~x731 & ~x776;
assign c2109 =  x51;
assign c2113 = ~x636 & ~x637 & ~x666 & ~x679 & ~x694;
assign c2115 =  x448;
assign c2117 =  x69 & ~x38 & ~x262;
assign c2119 =  x15 &  x92 &  x175 &  x178 &  x289 &  x344 &  x355 &  x372 &  x381 &  x403 &  x441 &  x464 &  x485 &  x489 &  x498 &  x525 &  x544 & ~x4 & ~x22 & ~x27 & ~x29 & ~x30 & ~x32 & ~x33 & ~x47 & ~x56 & ~x141 & ~x142 & ~x144 & ~x164 & ~x198 & ~x250 & ~x281 & ~x335 & ~x419 & ~x501 & ~x562 & ~x588 & ~x618 & ~x643 & ~x671 & ~x674 & ~x699;
assign c2121 =  x362;
assign c2123 =  x25;
assign c2125 =  x41 &  x43 &  x93 &  x209 &  x215 &  x239 &  x260 &  x317 &  x324 &  x347 &  x349 &  x384 & ~x10 & ~x11 & ~x28 & ~x29 & ~x30 & ~x31 & ~x33 & ~x35 & ~x46 & ~x48 & ~x49 & ~x51 & ~x55 & ~x57 & ~x63 & ~x90 & ~x106 & ~x107 & ~x113 & ~x142 & ~x143 & ~x164 & ~x165 & ~x167 & ~x191 & ~x197 & ~x199 & ~x220 & ~x337 & ~x360 & ~x364 & ~x390 & ~x391 & ~x392 & ~x416 & ~x419 & ~x423 & ~x447 & ~x448 & ~x450 & ~x451 & ~x474 & ~x532 & ~x534 & ~x557 & ~x585 & ~x586 & ~x590 & ~x613 & ~x643 & ~x645 & ~x700 & ~x701 & ~x729 & ~x753 & ~x755 & ~x759 & ~x764 & ~x775;
assign c2127 =  x334;
assign c2129 =  x13 &  x15 &  x40 &  x73 &  x98 &  x101 &  x122 &  x130 &  x148 &  x158 &  x177 &  x179 &  x180 &  x184 &  x186 &  x187 &  x206 &  x209 &  x210 &  x211 &  x232 &  x237 &  x243 &  x244 &  x261 &  x262 &  x264 &  x265 &  x268 &  x288 &  x289 &  x290 &  x292 &  x294 &  x297 &  x301 &  x314 &  x316 &  x325 &  x342 &  x345 &  x348 &  x351 &  x356 &  x370 &  x371 &  x372 &  x373 &  x374 &  x379 &  x385 &  x398 &  x402 &  x406 &  x408 &  x410 &  x413 &  x430 &  x431 &  x432 &  x434 &  x435 &  x437 &  x459 &  x461 &  x464 &  x485 &  x488 &  x491 &  x492 &  x494 &  x498 &  x510 &  x513 &  x514 &  x516 &  x517 &  x526 &  x545 &  x547 &  x549 &  x550 &  x554 &  x569 & ~x5 & ~x7 & ~x8 & ~x9 & ~x18 & ~x23 & ~x24 & ~x27 & ~x29 & ~x30 & ~x32 & ~x34 & ~x35 & ~x36 & ~x49 & ~x53 & ~x54 & ~x56 & ~x59 & ~x62 & ~x84 & ~x85 & ~x109 & ~x113 & ~x114 & ~x115 & ~x135 & ~x171 & ~x192 & ~x195 & ~x196 & ~x199 & ~x220 & ~x222 & ~x225 & ~x226 & ~x250 & ~x277 & ~x309 & ~x310 & ~x336 & ~x337 & ~x338 & ~x364 & ~x365 & ~x393 & ~x449 & ~x473 & ~x475 & ~x477 & ~x502 & ~x529 & ~x531 & ~x558 & ~x559 & ~x560 & ~x585 & ~x586 & ~x615 & ~x616 & ~x642 & ~x643 & ~x670 & ~x672 & ~x700 & ~x726 & ~x727 & ~x729 & ~x754 & ~x756 & ~x764 & ~x781;
assign c2131 =  x390;
assign c2133 =  x39 &  x45 & ~x6 & ~x365 & ~x481 & ~x508 & ~x621 & ~x638 & ~x642 & ~x646 & ~x647 & ~x667 & ~x674 & ~x676 & ~x695 & ~x751 & ~x762;
assign c2135 =  x47 & ~x610;
assign c2137 =  x224;
assign c2139 =  x252;
assign c2141 =  x138;
assign c2143 =  x82;
assign c2147 =  x194;
assign c2149 =  x194;
assign c2151 =  x411 &  x495 &  x512 &  x552 &  x661 &  x692 &  x720 &  x721 &  x744 &  x747 & ~x1 & ~x23 & ~x82 & ~x225 & ~x306 & ~x310 & ~x671 & ~x672 & ~x753 & ~x757 & ~x761;
assign c2153 =  x699;
assign c2155 =  x141;
assign c2157 =  x278;
assign c2159 =  x222;
assign c2161 =  x74 &  x151 &  x184 &  x206 &  x234 &  x235 &  x236 &  x240 &  x242 &  x263 &  x295 &  x346 &  x352 &  x377 &  x380 &  x401 &  x402 &  x407 &  x410 &  x413 &  x428 &  x432 &  x433 &  x485 &  x489 &  x494 &  x513 &  x518 &  x522 &  x523 &  x540 &  x550 &  x551 &  x569 &  x571 &  x575 &  x577 &  x578 &  x580 &  x597 &  x598 &  x599 &  x605 &  x606 &  x625 &  x629 &  x632 &  x634 &  x655 &  x662 &  x708 &  x711 &  x715 & ~x2 & ~x6 & ~x23 & ~x25 & ~x32 & ~x51 & ~x57 & ~x85 & ~x110 & ~x137 & ~x138 & ~x165 & ~x169 & ~x197 & ~x224 & ~x250 & ~x279 & ~x306 & ~x308 & ~x309 & ~x336 & ~x393 & ~x418 & ~x447 & ~x588 & ~x755 & ~x756 & ~x761 & ~x778 & ~x780;
assign c2163 =  x51;
assign c2165 =  x87;
assign c2167 =  x198;
assign c2169 =  x4;
assign c2171 =  x42 &  x43 &  x96 &  x101 &  x183 &  x188 &  x203 &  x204 &  x208 &  x234 &  x259 &  x269 &  x297 &  x301 &  x313 &  x326 &  x329 &  x346 &  x372 &  x382 &  x430 &  x462 &  x481 &  x498 &  x541 &  x543 &  x545 &  x551 &  x577 &  x609 & ~x9 & ~x26 & ~x31 & ~x36 & ~x46 & ~x89 & ~x115 & ~x136 & ~x144 & ~x222 & ~x225 & ~x226 & ~x252 & ~x277 & ~x279 & ~x281 & ~x366 & ~x391 & ~x393 & ~x478 & ~x557 & ~x757 & ~x763;
assign c2173 = ~x384 & ~x398 & ~x498;
assign c2175 = ~x10 & ~x17 & ~x36 & ~x38 & ~x180 & ~x263;
assign c2177 =  x700;
assign c2179 = ~x175 & ~x341;
assign c2181 =  x56 &  x194;
assign c2183 = ~x442 & ~x651 & ~x664;
assign c2185 =  x111;
assign c2187 = ~x398 & ~x427 & ~x481;
assign c2189 = ~x440 & ~x480 & ~x498 & ~x610 & ~x724 & ~x731;
assign c2191 =  x121 &  x151 &  x214 &  x236 &  x241 &  x267 &  x315 &  x324 &  x325 &  x351 &  x354 &  x398 &  x431 &  x437 &  x457 &  x516 &  x522 &  x548 &  x662 &  x688 &  x742 & ~x5 & ~x8 & ~x18 & ~x60 & ~x78 & ~x87 & ~x106 & ~x112 & ~x114 & ~x116 & ~x143 & ~x164 & ~x169 & ~x196 & ~x225 & ~x248 & ~x249 & ~x253 & ~x281 & ~x333 & ~x364 & ~x366 & ~x418 & ~x446 & ~x501 & ~x558 & ~x590 & ~x671 & ~x672 & ~x727 & ~x730 & ~x731 & ~x753 & ~x755 & ~x761 & ~x762 & ~x776 & ~x778 & ~x779;
assign c2193 =  x84;
assign c2195 =  x224;
assign c2197 =  x12 &  x65 &  x74 &  x100 &  x130 &  x153 &  x207 &  x211 &  x242 &  x243 &  x262 &  x266 &  x274 &  x297 &  x298 &  x326 &  x350 &  x370 &  x432 &  x481 &  x488 &  x543 &  x620 &  x648 &  x694 & ~x18 & ~x33 & ~x51 & ~x60 & ~x80 & ~x82 & ~x138 & ~x197 & ~x225 & ~x227 & ~x279 & ~x532 & ~x726 & ~x781;
assign c2199 =  x38 & ~x2 & ~x6 & ~x23 & ~x27 & ~x55 & ~x59 & ~x169 & ~x308 & ~x310 & ~x362 & ~x365 & ~x387 & ~x392 & ~x415 & ~x423 & ~x444 & ~x445 & ~x448 & ~x450 & ~x472 & ~x616 & ~x619 & ~x668 & ~x672 & ~x703 & ~x705 & ~x724 & ~x732 & ~x734 & ~x753 & ~x782;
assign c2201 =  x728;
assign c2203 =  x40 &  x66 &  x68 &  x155 &  x156 &  x182 &  x185 &  x217 &  x235 &  x268 &  x269 &  x270 &  x285 &  x313 &  x316 &  x324 &  x330 &  x355 &  x357 &  x370 &  x371 &  x376 &  x378 &  x379 &  x380 &  x399 &  x413 &  x433 &  x437 &  x459 &  x464 &  x489 &  x514 &  x519 &  x526 &  x536 &  x537 &  x538 &  x541 &  x550 &  x553 &  x564 &  x565 &  x593 &  x609 &  x620 &  x637 &  x722 & ~x3 & ~x7 & ~x8 & ~x9 & ~x27 & ~x56 & ~x58 & ~x59 & ~x60 & ~x78 & ~x83 & ~x84 & ~x85 & ~x86 & ~x113 & ~x116 & ~x137 & ~x140 & ~x141 & ~x165 & ~x170 & ~x172 & ~x193 & ~x196 & ~x223 & ~x226 & ~x251 & ~x253 & ~x278 & ~x304 & ~x305 & ~x310 & ~x332 & ~x366 & ~x390 & ~x421 & ~x505 & ~x533 & ~x562 & ~x586 & ~x587 & ~x589 & ~x644 & ~x699 & ~x754 & ~x758;
assign c2205 =  x776;
assign c2207 =  x756;
assign c2211 =  x43 &  x66 &  x67 &  x188 &  x204 &  x209 &  x267 &  x268 &  x269 &  x329 &  x342 &  x350 &  x403 &  x455 &  x542 &  x543 &  x554 &  x621 &  x632 &  x638 &  x653 &  x663 &  x684 & ~x8 & ~x28 & ~x82 & ~x84 & ~x89 & ~x135 & ~x136 & ~x140 & ~x141 & ~x163 & ~x171 & ~x172 & ~x200 & ~x250 & ~x278 & ~x312 & ~x362 & ~x531 & ~x641 & ~x647 & ~x702 & ~x774 & ~x776;
assign c2213 =  x477;
assign c2215 =  x69 &  x74 &  x95 &  x100 &  x153 &  x157 &  x182 &  x185 &  x187 &  x204 &  x210 &  x211 &  x213 &  x234 &  x238 &  x241 &  x244 &  x260 &  x261 &  x271 &  x298 &  x318 &  x322 &  x324 &  x344 &  x345 &  x347 &  x351 &  x352 &  x375 &  x376 &  x379 &  x382 &  x401 &  x404 &  x407 &  x409 &  x411 &  x431 &  x433 &  x436 &  x459 &  x461 &  x465 &  x467 &  x486 &  x491 &  x492 &  x494 &  x495 &  x513 &  x514 &  x521 &  x547 &  x550 &  x552 &  x567 &  x570 &  x571 &  x580 &  x597 &  x602 &  x603 &  x606 &  x627 &  x632 &  x651 &  x653 &  x661 &  x663 &  x665 &  x681 &  x687 &  x714 & ~x3 & ~x8 & ~x19 & ~x23 & ~x25 & ~x26 & ~x27 & ~x30 & ~x56 & ~x58 & ~x80 & ~x85 & ~x110 & ~x111 & ~x137 & ~x142 & ~x226 & ~x253 & ~x278 & ~x280 & ~x282 & ~x306 & ~x361 & ~x364 & ~x366 & ~x393 & ~x419 & ~x420 & ~x447 & ~x449 & ~x450 & ~x474 & ~x503 & ~x504 & ~x558 & ~x559 & ~x616 & ~x671 & ~x672 & ~x701 & ~x702 & ~x727 & ~x728 & ~x756 & ~x759 & ~x782 & ~x783;
assign c2217 =  x251;
assign c2219 = ~x51 & ~x195 & ~x418 & ~x537 & ~x554 & ~x563 & ~x588 & ~x609 & ~x611 & ~x638 & ~x671 & ~x722 & ~x750 & ~x751 & ~x761;
assign c2221 =  x363;
assign c2223 =  x336;
assign c2225 =  x225;
assign c2227 =  x139;
assign c2229 = ~x11 & ~x45 & ~x47 & ~x48 & ~x160;
assign c2231 =  x420;
assign c2233 =  x2;
assign c2235 =  x169;
assign c2237 =  x32;
assign c2239 =  x252;
assign c2241 =  x538 &  x566 & ~x2 & ~x8 & ~x9 & ~x17 & ~x20 & ~x29 & ~x30 & ~x31 & ~x35 & ~x37 & ~x48 & ~x62 & ~x83 & ~x84 & ~x89 & ~x106 & ~x108 & ~x109 & ~x135 & ~x137 & ~x161 & ~x196 & ~x224 & ~x281 & ~x420 & ~x755;
assign c2243 =  x616;
assign c2247 =  x111;
assign c2249 =  x375 &  x467 &  x652 &  x681 & ~x285 & ~x333 & ~x676 & ~x727;
assign c2251 =  x80;
assign c2253 =  x141;
assign c2255 =  x66 & ~x57 & ~x109 & ~x196 & ~x225 & ~x282 & ~x334 & ~x414 & ~x443 & ~x479 & ~x564 & ~x592 & ~x639 & ~x647 & ~x724 & ~x725 & ~x762;
assign c2257 =  x86;
assign c2259 =  x588;
assign c2261 =  x363;
assign c2263 =  x26;
assign c2265 =  x475;
assign c2267 =  x249;
assign c2269 = ~x17 & ~x37 & ~x38 & ~x39 & ~x65 & ~x117 & ~x122;
assign c2271 =  x138;
assign c2273 =  x194 &  x644;
assign c2275 = ~x454 & ~x592;
assign c2277 =  x280;
assign c2279 =  x66 &  x179 &  x186 &  x381 &  x599 & ~x251 & ~x393 & ~x476 & ~x503 & ~x702 & ~x705 & ~x734 & ~x764;
assign c2281 = ~x21 & ~x250 & ~x397 & ~x725 & ~x732 & ~x734 & ~x762 & ~x766;
assign c2283 =  x12 &  x42 &  x91 &  x287 &  x288 &  x343 & ~x8 & ~x17 & ~x19 & ~x28 & ~x29 & ~x32 & ~x34 & ~x35 & ~x47 & ~x50 & ~x52 & ~x58 & ~x59 & ~x60 & ~x85 & ~x106 & ~x111 & ~x114 & ~x135 & ~x195 & ~x224 & ~x277 & ~x280 & ~x333 & ~x335 & ~x336 & ~x337 & ~x363 & ~x417 & ~x418 & ~x448 & ~x450 & ~x533 & ~x589 & ~x643 & ~x644 & ~x671 & ~x701 & ~x726 & ~x758 & ~x764;
assign c2285 = ~x536 & ~x592 & ~x608 & ~x638 & ~x750;
assign c2287 =  x103 &  x495 &  x664 &  x707 & ~x620;
assign c2289 =  x224;
assign c2291 =  x365;
assign c2293 =  x4;
assign c2295 =  x361;
assign c2297 =  x26 &  x757;
assign c2299 =  x4;
assign c2301 =  x51;
assign c2303 =  x169;
assign c2305 =  x248 & ~x752;
assign c2307 =  x310;
assign c2309 = ~x99;
assign c2311 =  x168;
assign c2313 =  x643;
assign c2315 =  x14 &  x66 &  x96 &  x98 &  x99 &  x122 &  x124 &  x125 &  x126 &  x127 &  x128 &  x154 &  x159 &  x178 &  x187 &  x212 &  x231 &  x232 &  x234 &  x235 &  x239 &  x240 &  x259 &  x266 &  x268 &  x269 &  x289 &  x297 &  x298 &  x318 &  x321 &  x323 &  x348 &  x351 &  x352 &  x353 &  x357 &  x374 &  x377 &  x378 &  x383 &  x385 &  x401 &  x405 &  x407 &  x408 &  x411 &  x431 &  x432 &  x457 &  x458 &  x459 &  x482 &  x485 &  x487 &  x514 &  x518 &  x519 &  x542 &  x545 &  x569 &  x573 &  x577 &  x582 &  x598 &  x599 &  x602 &  x604 &  x625 &  x633 &  x660 & ~x0 & ~x5 & ~x7 & ~x9 & ~x17 & ~x19 & ~x24 & ~x30 & ~x32 & ~x35 & ~x58 & ~x60 & ~x61 & ~x62 & ~x79 & ~x80 & ~x82 & ~x85 & ~x87 & ~x88 & ~x89 & ~x110 & ~x116 & ~x138 & ~x139 & ~x142 & ~x143 & ~x165 & ~x168 & ~x171 & ~x196 & ~x221 & ~x226 & ~x280 & ~x281 & ~x282 & ~x307 & ~x333 & ~x335 & ~x337 & ~x364 & ~x390 & ~x420 & ~x445 & ~x446 & ~x449 & ~x477 & ~x532 & ~x534 & ~x617 & ~x642 & ~x645 & ~x671 & ~x673 & ~x701 & ~x729 & ~x756 & ~x757 & ~x758 & ~x776 & ~x781 & ~x783;
assign c2317 =  x522 &  x541 &  x596 &  x651 &  x664 &  x708 & ~x55 & ~x111 & ~x334 & ~x418 & ~x452 & ~x472 & ~x479 & ~x589 & ~x641 & ~x752 & ~x755;
assign c2319 =  x23;
assign c2321 =  x24;
assign c2323 =  x27;
assign c2325 =  x447;
assign c2327 =  x363;
assign c2329 = ~x87 & ~x610 & ~x637 & ~x667 & ~x669 & ~x750 & ~x751;
assign c2333 =  x262 &  x271 &  x298 &  x314 &  x317 &  x321 &  x323 &  x344 &  x354 &  x356 &  x377 &  x378 &  x384 &  x413 &  x441 &  x458 &  x463 &  x494 &  x518 &  x522 &  x526 &  x542 &  x569 &  x570 &  x571 &  x579 &  x594 &  x595 &  x603 &  x611 &  x628 &  x630 &  x631 &  x636 &  x638 &  x657 &  x664 &  x678 &  x694 &  x695 &  x705 &  x706 & ~x18 & ~x21 & ~x22 & ~x23 & ~x27 & ~x30 & ~x136 & ~x138 & ~x168 & ~x170 & ~x253 & ~x362 & ~x364 & ~x365 & ~x419 & ~x475 & ~x476 & ~x645 & ~x783;
assign c2335 =  x141;
assign c2339 =  x112;
assign c2341 =  x510 & ~x11 & ~x46;
assign c2343 = ~x412 & ~x526;
assign c2345 = ~x230 & ~x367;
assign c2347 =  x316 &  x318 &  x319 &  x321 &  x399 &  x440 &  x485 &  x520 &  x521 &  x571 &  x629 &  x638 &  x665 & ~x20 & ~x28 & ~x46 & ~x113 & ~x142 & ~x167 & ~x227 & ~x700 & ~x748 & ~x775;
assign c2349 =  x65 &  x290 &  x294 &  x347 &  x355 &  x372 &  x437 &  x439 &  x458 &  x459 &  x468 &  x513 &  x516 &  x520 &  x544 &  x568 &  x651 &  x664 &  x692 &  x711 &  x718 &  x719 &  x720 & ~x6 & ~x23 & ~x30 & ~x53 & ~x58 & ~x81 & ~x86 & ~x140 & ~x197 & ~x221 & ~x222 & ~x249 & ~x277 & ~x281 & ~x363 & ~x365 & ~x530 & ~x587 & ~x673 & ~x780;
assign c2351 = ~x11 & ~x37 & ~x38 & ~x47 & ~x183;
assign c2353 =  x23;
assign c2355 =  x82;
assign c2357 =  x130 &  x179 &  x213 &  x234 &  x237 &  x257 &  x260 &  x261 &  x264 &  x266 &  x295 &  x300 &  x315 &  x320 &  x324 &  x341 &  x343 &  x346 &  x350 &  x353 &  x355 &  x370 &  x371 &  x372 &  x373 &  x376 &  x377 &  x378 &  x380 &  x384 &  x399 &  x401 &  x409 &  x410 &  x412 &  x414 &  x425 &  x433 &  x434 &  x436 &  x453 &  x455 &  x469 &  x493 &  x494 &  x499 &  x518 &  x521 &  x526 &  x537 &  x538 &  x542 &  x547 &  x548 &  x555 &  x566 &  x571 &  x574 &  x575 &  x582 &  x583 &  x592 &  x593 &  x601 &  x610 &  x611 &  x620 &  x627 &  x629 &  x635 & ~x1 & ~x2 & ~x6 & ~x7 & ~x8 & ~x9 & ~x18 & ~x19 & ~x27 & ~x29 & ~x32 & ~x34 & ~x36 & ~x48 & ~x50 & ~x54 & ~x55 & ~x57 & ~x58 & ~x59 & ~x63 & ~x80 & ~x81 & ~x84 & ~x86 & ~x107 & ~x109 & ~x110 & ~x112 & ~x113 & ~x140 & ~x166 & ~x169 & ~x194 & ~x223 & ~x363 & ~x364 & ~x447 & ~x503 & ~x644 & ~x700 & ~x754 & ~x756 & ~x757 & ~x758 & ~x775;
assign c2359 =  x127 &  x314 &  x342 &  x770 & ~x52 & ~x59 & ~x281 & ~x391 & ~x560 & ~x588 & ~x728 & ~x765 & ~x775;
assign c2361 =  x66 &  x121 &  x157 &  x159 &  x177 &  x180 &  x181 &  x205 &  x207 &  x215 &  x234 &  x272 &  x347 &  x351 &  x354 &  x409 &  x429 &  x469 &  x492 &  x515 &  x525 &  x597 &  x600 &  x604 &  x633 &  x662 &  x683 &  x715 &  x739 &  x741 & ~x1 & ~x23 & ~x25 & ~x29 & ~x35 & ~x54 & ~x55 & ~x82 & ~x108 & ~x114 & ~x139 & ~x166 & ~x169 & ~x194 & ~x225 & ~x254 & ~x278 & ~x279 & ~x281 & ~x334 & ~x335 & ~x336 & ~x389 & ~x445 & ~x447 & ~x448 & ~x560 & ~x561 & ~x587 & ~x588 & ~x727 & ~x729 & ~x761 & ~x762 & ~x782;
assign c2363 = ~x45 & ~x145 & ~x264;
assign c2365 =  x25;
assign c2367 = ~x17 & ~x37 & ~x45;
assign c2369 = ~x316;
assign c2371 =  x532;
assign c2373 =  x783;
assign c2375 =  x58;
assign c2377 =  x487 &  x547 & ~x42;
assign c2379 =  x14 &  x103 &  x156 &  x161 &  x181 &  x231 &  x241 &  x274 &  x300 &  x314 &  x357 &  x380 &  x415 & ~x10 & ~x27 & ~x35 & ~x36 & ~x54 & ~x77 & ~x78 & ~x111 & ~x171 & ~x394 & ~x765;
assign c2381 =  x55;
assign c2383 = ~x23 & ~x140 & ~x441 & ~x449 & ~x468 & ~x477 & ~x583 & ~x638 & ~x667 & ~x723;
assign c2385 =  x392;
assign c2387 =  x123 &  x131 &  x159 &  x203 &  x231 &  x267 &  x271 &  x329 &  x686 &  x687 & ~x22 & ~x53 & ~x58 & ~x197 & ~x420 & ~x532 & ~x589 & ~x644 & ~x648 & ~x676 & ~x732 & ~x778 & ~x779 & ~x780;
assign c2389 = ~x370 & ~x607;
assign c2391 =  x195;
assign c2393 =  x29;
assign c2395 =  x83;
assign c2397 =  x195;
assign c2399 =  x111;
assign c2401 = ~x387 & ~x470 & ~x498 & ~x499 & ~x536 & ~x563 & ~x590 & ~x621 & ~x639 & ~x641 & ~x698 & ~x723 & ~x724 & ~x777;
assign c2403 =  x86;
assign c2405 =  x40 &  x125 &  x151 &  x185 &  x210 &  x211 &  x290 &  x327 &  x345 &  x353 &  x356 &  x426 &  x458 &  x484 &  x512 &  x523 &  x569 &  x604 &  x621 &  x623 & ~x19 & ~x57 & ~x61 & ~x82 & ~x191 & ~x197 & ~x340 & ~x668 & ~x726 & ~x731;
assign c2407 = ~x175 & ~x202;
assign c2409 =  x26;
assign c2411 = ~x17 & ~x46 & ~x211;
assign c2413 =  x40 &  x42 &  x43 &  x68 &  x98 &  x123 &  x125 &  x128 &  x129 &  x152 &  x185 &  x187 &  x212 &  x214 &  x217 &  x238 &  x244 &  x258 &  x260 &  x262 &  x263 &  x264 &  x267 &  x270 &  x294 &  x299 &  x300 &  x301 &  x302 &  x315 &  x321 &  x322 &  x323 &  x324 &  x325 &  x329 &  x347 &  x353 &  x354 &  x374 &  x377 &  x378 &  x380 &  x381 &  x400 &  x405 &  x408 &  x414 &  x428 &  x432 &  x435 &  x438 &  x442 &  x460 &  x485 &  x488 &  x490 &  x493 &  x514 &  x515 &  x519 &  x521 &  x538 &  x545 &  x553 &  x570 &  x576 &  x578 &  x579 &  x601 &  x610 &  x624 &  x633 &  x634 &  x677 &  x705 &  x734 & ~x1 & ~x5 & ~x6 & ~x7 & ~x8 & ~x18 & ~x23 & ~x28 & ~x29 & ~x35 & ~x49 & ~x50 & ~x55 & ~x56 & ~x58 & ~x60 & ~x82 & ~x87 & ~x106 & ~x107 & ~x108 & ~x116 & ~x135 & ~x136 & ~x170 & ~x193 & ~x196 & ~x199 & ~x221 & ~x223 & ~x225 & ~x253 & ~x254 & ~x279 & ~x281 & ~x282 & ~x283 & ~x304 & ~x393 & ~x417 & ~x418 & ~x419 & ~x448 & ~x449 & ~x529 & ~x532 & ~x534 & ~x557 & ~x561 & ~x562 & ~x617 & ~x646 & ~x700 & ~x725 & ~x756 & ~x764 & ~x765 & ~x775;
assign c2415 = ~x39 & ~x286;
assign c2417 =  x81;
assign c2419 =  x448;
assign c2421 = ~x23 & ~x426 & ~x480 & ~x507 & ~x527 & ~x533 & ~x619 & ~x695 & ~x731 & ~x756 & ~x764 & ~x777;
assign c2423 =  x324 &  x347 &  x351 &  x359 &  x380 &  x407 &  x426 &  x441 &  x453 &  x466 &  x527 &  x569 &  x576 &  x601 &  x625 &  x649 &  x665 &  x668 &  x677 &  x693 &  x696 & ~x7 & ~x55 & ~x81 & ~x87 & ~x113 & ~x192 & ~x196 & ~x307;
assign c2425 =  x56;
assign c2427 =  x410 & ~x146 & ~x147;
assign c2429 =  x366;
assign c2431 =  x167;
assign c2433 =  x250;
assign c2437 =  x502;
assign c2439 =  x371 &  x399 &  x427 &  x510 &  x538 &  x553 &  x594 & ~x3 & ~x4 & ~x7 & ~x9 & ~x11 & ~x17 & ~x19 & ~x21 & ~x31 & ~x36 & ~x45 & ~x47 & ~x52 & ~x53 & ~x54 & ~x61 & ~x64 & ~x85 & ~x106 & ~x108 & ~x111 & ~x113 & ~x117 & ~x139 & ~x142 & ~x144 & ~x167 & ~x194 & ~x195 & ~x196 & ~x224 & ~x280 & ~x309 & ~x392 & ~x559 & ~x560 & ~x587 & ~x672 & ~x700 & ~x727 & ~x754 & ~x755 & ~x757 & ~x783;
assign c2441 =  x112 &  x251;
assign c2443 =  x336;
assign c2445 =  x194;
assign c2447 =  x729;
assign c2449 =  x166;
assign c2451 = ~x10 & ~x38 & ~x234 & ~x262 & ~x731;
assign c2453 =  x109;
assign c2455 = ~x17 & ~x38 & ~x180;
assign c2459 =  x3;
assign c2461 =  x446;
assign c2463 =  x28 &  x336;
assign c2465 =  x250;
assign c2467 =  x384 &  x482 & ~x6 & ~x7 & ~x9 & ~x21 & ~x32 & ~x37 & ~x46 & ~x54 & ~x60 & ~x64 & ~x75 & ~x77 & ~x82 & ~x84 & ~x106 & ~x108 & ~x111 & ~x114 & ~x115 & ~x117 & ~x135 & ~x142 & ~x166 & ~x169 & ~x170 & ~x171 & ~x195 & ~x196 & ~x198 & ~x200 & ~x220 & ~x223 & ~x252 & ~x255 & ~x281 & ~x283 & ~x309 & ~x339 & ~x362 & ~x395 & ~x419 & ~x423 & ~x447 & ~x532 & ~x585 & ~x587 & ~x616 & ~x618 & ~x672 & ~x674 & ~x728 & ~x731 & ~x748 & ~x755 & ~x757 & ~x759 & ~x764;
assign c2469 =  x375 &  x379 &  x385 &  x406 &  x426 &  x427 &  x433 &  x437 &  x459 &  x463 &  x468 &  x485 &  x490 &  x524 &  x538 &  x539 &  x552 &  x554 &  x566 &  x573 &  x579 &  x582 &  x594 &  x596 &  x607 &  x624 &  x626 &  x633 &  x637 &  x653 &  x654 &  x663 & ~x2 & ~x9 & ~x48 & ~x54 & ~x58 & ~x77 & ~x107 & ~x110 & ~x117 & ~x145 & ~x162 & ~x163 & ~x165 & ~x166 & ~x173 & ~x192 & ~x221 & ~x226 & ~x249 & ~x250 & ~x251 & ~x419 & ~x701 & ~x728 & ~x756 & ~x758;
assign c2471 =  x167;
assign c2473 =  x197;
assign c2477 =  x429 &  x552 & ~x90 & ~x105 & ~x162 & ~x164 & ~x174;
assign c2479 =  x40 &  x42 &  x66 &  x103 &  x566 &  x581 & ~x0 & ~x3 & ~x8 & ~x9 & ~x10 & ~x17 & ~x28 & ~x37 & ~x49 & ~x51 & ~x53 & ~x56 & ~x58 & ~x63 & ~x77 & ~x78 & ~x80 & ~x84 & ~x86 & ~x106 & ~x166 & ~x197 & ~x198 & ~x221 & ~x248 & ~x253 & ~x282 & ~x283 & ~x284 & ~x306 & ~x335 & ~x363 & ~x366 & ~x367 & ~x390 & ~x393 & ~x421 & ~x446 & ~x476 & ~x502 & ~x507 & ~x586 & ~x617 & ~x644 & ~x673 & ~x699 & ~x700 & ~x702 & ~x748 & ~x776;
assign c2481 =  x399 &  x402 &  x404 &  x410 &  x411 &  x427 &  x428 &  x439 &  x458 &  x468 &  x513 &  x522 &  x542 &  x552 &  x569 &  x597 &  x606 &  x608 &  x624 &  x650 &  x651 &  x664 &  x721 &  x722 &  x735 & ~x6 & ~x26 & ~x141 & ~x307 & ~x615 & ~x642 & ~x672 & ~x727;
assign c2483 =  x222;
assign c2485 =  x273 & ~x481 & ~x510;
assign c2487 =  x196;
assign c2489 =  x93 &  x121 &  x632 & ~x443 & ~x500 & ~x527 & ~x704;
assign c2491 =  x736 &  x747 & ~x396 & ~x415 & ~x621 & ~x668;
assign c2493 =  x82;
assign c2495 =  x40 &  x41 &  x43 &  x66 &  x71 &  x73 &  x96 &  x123 &  x154 &  x180 &  x182 &  x188 &  x203 &  x206 &  x208 &  x209 &  x212 &  x233 &  x240 &  x241 &  x261 &  x263 &  x264 &  x267 &  x268 &  x288 &  x292 &  x295 &  x299 &  x301 &  x318 &  x324 &  x327 &  x329 &  x347 &  x351 &  x357 &  x358 &  x373 &  x377 &  x380 &  x381 &  x382 &  x402 &  x414 &  x431 &  x438 &  x454 &  x458 &  x469 &  x515 &  x521 &  x522 &  x541 &  x542 &  x546 &  x570 &  x571 &  x573 &  x578 &  x593 &  x594 &  x609 &  x610 &  x627 &  x633 &  x694 &  x705 & ~x0 & ~x31 & ~x33 & ~x49 & ~x50 & ~x54 & ~x56 & ~x60 & ~x87 & ~x108 & ~x113 & ~x116 & ~x137 & ~x163 & ~x164 & ~x167 & ~x192 & ~x196 & ~x250 & ~x254 & ~x255 & ~x278 & ~x308 & ~x332 & ~x336 & ~x362 & ~x366 & ~x389 & ~x392 & ~x446 & ~x477 & ~x501 & ~x505 & ~x532 & ~x534 & ~x561 & ~x588 & ~x614 & ~x618 & ~x673 & ~x698 & ~x725 & ~x726 & ~x736 & ~x755 & ~x765 & ~x782;
assign c2497 = ~x10 & ~x37 & ~x46 & ~x47 & ~x106 & ~x208 & ~x264;
assign c2499 =  x58;
assign c30 = ~x135 & ~x146 & ~x200 & ~x239 & ~x254 & ~x330 & ~x332 & ~x333 & ~x528 & ~x580 & ~x619 & ~x636 & ~x667 & ~x694;
assign c32 =  x370 & ~x24 & ~x28 & ~x30 & ~x60 & ~x61 & ~x88 & ~x106 & ~x107 & ~x113 & ~x117 & ~x139 & ~x165 & ~x167 & ~x219 & ~x228 & ~x279 & ~x306 & ~x337 & ~x420 & ~x448 & ~x449 & ~x452 & ~x475 & ~x500 & ~x503 & ~x529 & ~x562 & ~x591 & ~x595 & ~x610 & ~x614 & ~x619 & ~x642 & ~x646 & ~x650 & ~x667 & ~x674 & ~x675 & ~x676 & ~x699 & ~x752;
assign c34 =  x626 & ~x3 & ~x23 & ~x25 & ~x29 & ~x54 & ~x55 & ~x57 & ~x87 & ~x111 & ~x136 & ~x141 & ~x197 & ~x221 & ~x251 & ~x252 & ~x277 & ~x308 & ~x317 & ~x340 & ~x389 & ~x390 & ~x392 & ~x418 & ~x472 & ~x480 & ~x500 & ~x556 & ~x560 & ~x618 & ~x646 & ~x651 & ~x665 & ~x674 & ~x678 & ~x727 & ~x750 & ~x756 & ~x762 & ~x778;
assign c36 =  x122 & ~x14 & ~x42 & ~x81 & ~x108 & ~x194 & ~x251 & ~x279 & ~x282 & ~x311 & ~x334 & ~x360 & ~x362 & ~x388 & ~x417 & ~x476 & ~x503 & ~x560 & ~x729;
assign c38 =  x750;
assign c310 =  x41 &  x46 &  x47 &  x545 &  x600 &  x658 &  x713 & ~x4 & ~x28 & ~x52 & ~x54 & ~x55 & ~x199 & ~x228 & ~x256 & ~x304 & ~x308 & ~x419 & ~x447 & ~x449 & ~x477 & ~x667 & ~x695 & ~x754 & ~x777;
assign c312 = ~x26 & ~x61 & ~x110 & ~x112 & ~x182 & ~x196 & ~x201 & ~x220 & ~x229 & ~x247 & ~x281 & ~x308 & ~x332 & ~x416 & ~x424 & ~x452 & ~x504 & ~x508 & ~x529 & ~x561 & ~x579 & ~x759;
assign c314 = ~x2 & ~x5 & ~x7 & ~x9 & ~x18 & ~x20 & ~x21 & ~x27 & ~x30 & ~x48 & ~x56 & ~x58 & ~x60 & ~x61 & ~x69 & ~x85 & ~x90 & ~x115 & ~x116 & ~x166 & ~x167 & ~x169 & ~x195 & ~x223 & ~x249 & ~x337 & ~x363 & ~x559 & ~x587 & ~x592 & ~x613 & ~x619 & ~x641 & ~x643 & ~x644 & ~x672 & ~x673 & ~x674 & ~x678 & ~x699 & ~x730 & ~x732 & ~x733 & ~x751 & ~x755 & ~x762 & ~x778;
assign c316 =  x38 &  x91 &  x386 &  x741 & ~x86 & ~x171 & ~x648 & ~x676;
assign c318 =  x65 &  x92 &  x314 &  x716 & ~x219 & ~x228 & ~x281 & ~x333 & ~x337 & ~x672 & ~x695 & ~x723 & ~x729 & ~x733 & ~x762;
assign c320 = ~x7 & ~x13 & ~x14 & ~x20 & ~x24 & ~x31 & ~x32 & ~x54 & ~x55 & ~x56 & ~x78 & ~x81 & ~x86 & ~x106 & ~x116 & ~x142 & ~x144 & ~x165 & ~x174 & ~x187 & ~x190 & ~x196 & ~x217 & ~x218 & ~x220 & ~x226 & ~x227 & ~x231 & ~x260 & ~x273 & ~x281 & ~x288 & ~x299 & ~x301 & ~x302 & ~x311 & ~x315 & ~x329 & ~x337 & ~x356 & ~x357 & ~x360 & ~x367 & ~x368 & ~x370 & ~x371 & ~x385 & ~x386 & ~x390 & ~x391 & ~x392 & ~x399 & ~x427 & ~x441 & ~x446 & ~x453 & ~x497 & ~x503 & ~x508 & ~x529 & ~x534 & ~x557 & ~x615 & ~x616 & ~x617 & ~x618 & ~x644 & ~x645 & ~x646 & ~x672 & ~x675 & ~x698 & ~x704 & ~x727 & ~x752 & ~x758 & ~x779 & ~x783;
assign c322 = ~x25 & ~x26 & ~x27 & ~x28 & ~x86 & ~x107 & ~x114 & ~x139 & ~x163 & ~x173 & ~x219 & ~x228 & ~x230 & ~x248 & ~x249 & ~x250 & ~x258 & ~x259 & ~x274 & ~x275 & ~x278 & ~x303 & ~x329 & ~x331 & ~x336 & ~x337 & ~x339 & ~x360 & ~x367 & ~x369 & ~x370 & ~x389 & ~x397 & ~x418 & ~x444 & ~x452 & ~x471 & ~x474 & ~x477 & ~x500 & ~x529 & ~x548 & ~x644 & ~x727 & ~x758 & ~x762 & ~x783;
assign c324 =  x434 &  x661 & ~x3 & ~x23 & ~x31 & ~x55 & ~x56 & ~x83 & ~x107 & ~x111 & ~x116 & ~x165 & ~x224 & ~x253 & ~x282 & ~x289 & ~x557 & ~x620 & ~x674 & ~x678 & ~x699 & ~x706;
assign c326 = ~x73 & ~x144 & ~x334 & ~x362 & ~x652 & ~x702 & ~x750 & ~x761;
assign c328 =  x10 &  x64 &  x70 &  x713 & ~x115 & ~x253 & ~x256 & ~x278 & ~x558 & ~x560 & ~x561 & ~x670;
assign c330 =  x41 &  x379 &  x434 &  x489 &  x517 &  x518 &  x546 &  x574 &  x659 &  x685 &  x741 & ~x1 & ~x10 & ~x19 & ~x22 & ~x48 & ~x52 & ~x60 & ~x80 & ~x106 & ~x113 & ~x117 & ~x139 & ~x164 & ~x173 & ~x200 & ~x201 & ~x229 & ~x275 & ~x283 & ~x308 & ~x362 & ~x366 & ~x368 & ~x414 & ~x442 & ~x447 & ~x454 & ~x501 & ~x502 & ~x530 & ~x531 & ~x558 & ~x586 & ~x614 & ~x669 & ~x670 & ~x673 & ~x725 & ~x727 & ~x755 & ~x781;
assign c332 = ~x156 & ~x257 & ~x273 & ~x549;
assign c334 =  x204 & ~x7 & ~x8 & ~x9 & ~x32 & ~x35 & ~x48 & ~x50 & ~x51 & ~x56 & ~x57 & ~x105 & ~x110 & ~x165 & ~x169 & ~x172 & ~x196 & ~x200 & ~x228 & ~x229 & ~x254 & ~x256 & ~x303 & ~x332 & ~x337 & ~x339 & ~x340 & ~x391 & ~x393 & ~x421 & ~x531 & ~x532 & ~x557 & ~x585 & ~x609 & ~x611 & ~x617 & ~x638 & ~x643 & ~x674 & ~x678 & ~x705 & ~x724 & ~x730 & ~x783;
assign c336 =  x10 &  x133 &  x684 & ~x54 & ~x87 & ~x139 & ~x169 & ~x335 & ~x364 & ~x447 & ~x617 & ~x758;
assign c338 = ~x260 & ~x299 & ~x329 & ~x342 & ~x403;
assign c340 =  x269 &  x495 & ~x28 & ~x29 & ~x84 & ~x115 & ~x141 & ~x167 & ~x197 & ~x248 & ~x279 & ~x289 & ~x333 & ~x359 & ~x365 & ~x390 & ~x419 & ~x447 & ~x449 & ~x506 & ~x613 & ~x614 & ~x645 & ~x674 & ~x698 & ~x757;
assign c342 =  x37 &  x45 &  x160 &  x272 & ~x3 & ~x24 & ~x32 & ~x59 & ~x60 & ~x62 & ~x78 & ~x86 & ~x89 & ~x117 & ~x143 & ~x169 & ~x170 & ~x193 & ~x196 & ~x197 & ~x252 & ~x282 & ~x284 & ~x362 & ~x364 & ~x395 & ~x477 & ~x616 & ~x668 & ~x676 & ~x762 & ~x783;
assign c344 =  x210 &  x378 &  x404 &  x406 &  x407 &  x459 &  x518 &  x520 &  x575 &  x714 &  x716 &  x739 &  x740 & ~x3 & ~x4 & ~x6 & ~x10 & ~x23 & ~x24 & ~x26 & ~x32 & ~x34 & ~x36 & ~x48 & ~x51 & ~x53 & ~x54 & ~x59 & ~x60 & ~x61 & ~x63 & ~x79 & ~x80 & ~x115 & ~x134 & ~x135 & ~x139 & ~x142 & ~x146 & ~x162 & ~x163 & ~x166 & ~x171 & ~x172 & ~x190 & ~x193 & ~x200 & ~x201 & ~x219 & ~x221 & ~x224 & ~x225 & ~x247 & ~x251 & ~x252 & ~x254 & ~x276 & ~x282 & ~x306 & ~x308 & ~x310 & ~x333 & ~x359 & ~x360 & ~x362 & ~x363 & ~x366 & ~x369 & ~x386 & ~x388 & ~x392 & ~x395 & ~x414 & ~x415 & ~x416 & ~x420 & ~x421 & ~x445 & ~x447 & ~x453 & ~x471 & ~x477 & ~x481 & ~x499 & ~x501 & ~x503 & ~x505 & ~x531 & ~x555 & ~x558 & ~x563 & ~x565 & ~x566 & ~x585 & ~x588 & ~x590 & ~x613 & ~x618 & ~x620 & ~x639 & ~x640 & ~x641 & ~x642 & ~x648 & ~x649 & ~x667 & ~x671 & ~x694 & ~x699 & ~x700 & ~x725 & ~x751 & ~x753 & ~x754 & ~x755 & ~x759 & ~x761 & ~x762 & ~x775 & ~x776 & ~x777 & ~x781;
assign c346 =  x446;
assign c348 = ~x97 & ~x268 & ~x478 & ~x501 & ~x507;
assign c350 =  x63 &  x741 & ~x4 & ~x52 & ~x54 & ~x86 & ~x172 & ~x198 & ~x199 & ~x220 & ~x224 & ~x248 & ~x251 & ~x253 & ~x278 & ~x311 & ~x336 & ~x338 & ~x447 & ~x476 & ~x531 & ~x616 & ~x779;
assign c352 =  x65 &  x210 &  x263 &  x436 & ~x0 & ~x3 & ~x23 & ~x111 & ~x136 & ~x139 & ~x197 & ~x220 & ~x226 & ~x248 & ~x249 & ~x253 & ~x272 & ~x277 & ~x300 & ~x315 & ~x363 & ~x364 & ~x418 & ~x504 & ~x588 & ~x644 & ~x671 & ~x700;
assign c354 =  x243 & ~x3 & ~x8 & ~x19 & ~x24 & ~x26 & ~x27 & ~x28 & ~x33 & ~x34 & ~x35 & ~x54 & ~x55 & ~x56 & ~x57 & ~x61 & ~x78 & ~x82 & ~x86 & ~x87 & ~x88 & ~x108 & ~x110 & ~x111 & ~x112 & ~x114 & ~x115 & ~x137 & ~x145 & ~x164 & ~x165 & ~x166 & ~x171 & ~x191 & ~x192 & ~x197 & ~x198 & ~x199 & ~x219 & ~x220 & ~x224 & ~x227 & ~x228 & ~x247 & ~x248 & ~x250 & ~x255 & ~x276 & ~x277 & ~x280 & ~x282 & ~x284 & ~x304 & ~x306 & ~x308 & ~x310 & ~x326 & ~x332 & ~x333 & ~x334 & ~x335 & ~x338 & ~x339 & ~x360 & ~x361 & ~x362 & ~x363 & ~x364 & ~x390 & ~x392 & ~x416 & ~x418 & ~x419 & ~x420 & ~x422 & ~x424 & ~x443 & ~x445 & ~x446 & ~x447 & ~x449 & ~x450 & ~x451 & ~x473 & ~x475 & ~x478 & ~x479 & ~x501 & ~x503 & ~x504 & ~x507 & ~x528 & ~x529 & ~x530 & ~x532 & ~x535 & ~x558 & ~x559 & ~x586 & ~x587 & ~x590 & ~x591 & ~x612 & ~x614 & ~x615 & ~x616 & ~x618 & ~x619 & ~x620 & ~x639 & ~x640 & ~x644 & ~x645 & ~x647 & ~x648 & ~x667 & ~x671 & ~x673 & ~x676 & ~x696 & ~x697 & ~x723 & ~x725 & ~x727 & ~x731 & ~x751 & ~x752 & ~x753 & ~x755 & ~x757 & ~x758 & ~x777 & ~x778 & ~x779 & ~x781 & ~x782 & ~x783;
assign c356 =  x411 & ~x19 & ~x159 & ~x224 & ~x305 & ~x339 & ~x417 & ~x452 & ~x726 & ~x758;
assign c358 =  x123 & ~x1 & ~x19 & ~x25 & ~x31 & ~x32 & ~x43 & ~x79 & ~x84 & ~x86 & ~x142 & ~x165 & ~x193 & ~x196 & ~x197 & ~x225 & ~x248 & ~x253 & ~x277 & ~x279 & ~x281 & ~x282 & ~x334 & ~x362 & ~x477 & ~x529 & ~x531 & ~x589 & ~x613 & ~x617 & ~x698 & ~x729 & ~x778;
assign c360 = ~x1 & ~x2 & ~x26 & ~x30 & ~x54 & ~x59 & ~x61 & ~x81 & ~x82 & ~x83 & ~x109 & ~x116 & ~x144 & ~x163 & ~x166 & ~x167 & ~x169 & ~x171 & ~x194 & ~x220 & ~x222 & ~x226 & ~x228 & ~x248 & ~x249 & ~x251 & ~x252 & ~x256 & ~x275 & ~x276 & ~x278 & ~x281 & ~x303 & ~x306 & ~x310 & ~x332 & ~x333 & ~x335 & ~x338 & ~x339 & ~x365 & ~x389 & ~x390 & ~x391 & ~x394 & ~x396 & ~x407 & ~x415 & ~x418 & ~x419 & ~x425 & ~x447 & ~x450 & ~x451 & ~x452 & ~x453 & ~x472 & ~x475 & ~x477 & ~x479 & ~x480 & ~x481 & ~x500 & ~x502 & ~x503 & ~x529 & ~x530 & ~x531 & ~x534 & ~x535 & ~x556 & ~x563 & ~x585 & ~x588 & ~x612 & ~x615 & ~x620 & ~x640 & ~x643 & ~x647 & ~x648 & ~x669 & ~x670 & ~x671 & ~x672 & ~x729 & ~x732 & ~x752 & ~x753 & ~x756 & ~x761 & ~x776 & ~x779 & ~x782;
assign c362 = ~x24 & ~x53 & ~x55 & ~x116 & ~x117 & ~x140 & ~x145 & ~x191 & ~x221 & ~x227 & ~x248 & ~x308 & ~x338 & ~x361 & ~x390 & ~x528 & ~x531 & ~x532 & ~x557 & ~x563 & ~x572 & ~x586 & ~x672 & ~x726 & ~x762 & ~x764 & ~x782;
assign c364 =  x292 &  x322 &  x718 & ~x25 & ~x271 & ~x365 & ~x387 & ~x426 & ~x730;
assign c366 =  x417;
assign c368 =  x406 &  x437 & ~x17 & ~x28 & ~x53 & ~x140 & ~x172 & ~x283 & ~x585 & ~x643 & ~x667 & ~x678 & ~x705 & ~x706 & ~x731;
assign c370 =  x132 &  x216 &  x246 & ~x5 & ~x82 & ~x194 & ~x197 & ~x534 & ~x639 & ~x667 & ~x669 & ~x675 & ~x704 & ~x730;
assign c372 = ~x31 & ~x84 & ~x95 & ~x140 & ~x179 & ~x201 & ~x306 & ~x360 & ~x369 & ~x414 & ~x472 & ~x508 & ~x557 & ~x580 & ~x620 & ~x694 & ~x763;
assign c374 = ~x128 & ~x288 & ~x372 & ~x611 & ~x640 & ~x672;
assign c376 =  x36 &  x42 &  x44 &  x63 & ~x2 & ~x54 & ~x110 & ~x113 & ~x169 & ~x220 & ~x228 & ~x247 & ~x248 & ~x249 & ~x275 & ~x391 & ~x500 & ~x501 & ~x532 & ~x534 & ~x588 & ~x616 & ~x755 & ~x779;
assign c378 =  x431 & ~x52 & ~x112 & ~x116 & ~x141 & ~x172 & ~x199 & ~x250 & ~x360 & ~x389 & ~x419 & ~x437 & ~x450 & ~x474 & ~x536 & ~x556 & ~x561 & ~x587 & ~x701;
assign c380 =  x155 &  x321 & ~x15 & ~x53 & ~x60 & ~x61 & ~x82 & ~x85 & ~x104 & ~x105 & ~x106 & ~x117 & ~x134 & ~x138 & ~x174 & ~x191 & ~x222 & ~x285 & ~x329 & ~x331 & ~x364 & ~x446 & ~x471 & ~x476 & ~x501 & ~x530 & ~x608 & ~x668 & ~x696 & ~x697 & ~x698 & ~x705 & ~x761 & ~x777;
assign c382 =  x746 & ~x68 & ~x131 & ~x530 & ~x534 & ~x762;
assign c384 =  x620 & ~x257;
assign c386 = ~x260 & ~x272 & ~x358 & ~x359 & ~x379 & ~x385 & ~x417 & ~x441 & ~x479 & ~x612 & ~x644;
assign c388 =  x46 &  x158 &  x689 & ~x171 & ~x254 & ~x310 & ~x424 & ~x454 & ~x505 & ~x538 & ~x595 & ~x615 & ~x705 & ~x723 & ~x732;
assign c390 =  x46 &  x66 &  x405 & ~x24 & ~x29 & ~x59 & ~x115 & ~x194 & ~x447 & ~x453 & ~x499 & ~x508 & ~x772;
assign c392 =  x153 &  x155 &  x237 &  x321 &  x347 &  x349 &  x403 &  x431 &  x464 &  x545 &  x546 &  x550 &  x596 &  x655 &  x684 & ~x27 & ~x77 & ~x80 & ~x89 & ~x105 & ~x135 & ~x167 & ~x171 & ~x225 & ~x279 & ~x280 & ~x309 & ~x331 & ~x334 & ~x361 & ~x364 & ~x392 & ~x396 & ~x448 & ~x473 & ~x530 & ~x562 & ~x565 & ~x611 & ~x613 & ~x642 & ~x731;
assign c394 = ~x4 & ~x8 & ~x49 & ~x69 & ~x71 & ~x72 & ~x82 & ~x106 & ~x115 & ~x143 & ~x220 & ~x283 & ~x305 & ~x365 & ~x447 & ~x473 & ~x530 & ~x613 & ~x703 & ~x755 & ~x757 & ~x764;
assign c396 =  x46 &  x317 & ~x2 & ~x27 & ~x115 & ~x138 & ~x141 & ~x144 & ~x225 & ~x275 & ~x278 & ~x337 & ~x421 & ~x443 & ~x756 & ~x758 & ~x761 & ~x762;
assign c398 =  x516 &  x570 &  x629 & ~x0 & ~x1 & ~x2 & ~x3 & ~x4 & ~x5 & ~x6 & ~x8 & ~x13 & ~x14 & ~x22 & ~x24 & ~x25 & ~x26 & ~x28 & ~x29 & ~x32 & ~x33 & ~x35 & ~x50 & ~x51 & ~x53 & ~x55 & ~x57 & ~x58 & ~x59 & ~x62 & ~x77 & ~x78 & ~x81 & ~x82 & ~x85 & ~x86 & ~x87 & ~x88 & ~x89 & ~x107 & ~x108 & ~x110 & ~x111 & ~x112 & ~x113 & ~x114 & ~x116 & ~x117 & ~x134 & ~x135 & ~x137 & ~x138 & ~x139 & ~x140 & ~x141 & ~x142 & ~x143 & ~x163 & ~x165 & ~x166 & ~x167 & ~x169 & ~x170 & ~x171 & ~x172 & ~x193 & ~x194 & ~x197 & ~x199 & ~x200 & ~x220 & ~x221 & ~x223 & ~x224 & ~x226 & ~x227 & ~x228 & ~x248 & ~x249 & ~x250 & ~x251 & ~x253 & ~x255 & ~x256 & ~x277 & ~x278 & ~x279 & ~x281 & ~x282 & ~x284 & ~x303 & ~x305 & ~x306 & ~x307 & ~x308 & ~x334 & ~x336 & ~x337 & ~x339 & ~x341 & ~x360 & ~x363 & ~x365 & ~x368 & ~x389 & ~x391 & ~x393 & ~x394 & ~x395 & ~x396 & ~x397 & ~x416 & ~x418 & ~x419 & ~x420 & ~x422 & ~x424 & ~x448 & ~x449 & ~x450 & ~x451 & ~x452 & ~x454 & ~x475 & ~x476 & ~x477 & ~x480 & ~x502 & ~x503 & ~x504 & ~x507 & ~x508 & ~x527 & ~x528 & ~x529 & ~x530 & ~x531 & ~x532 & ~x534 & ~x536 & ~x558 & ~x559 & ~x560 & ~x561 & ~x584 & ~x585 & ~x587 & ~x589 & ~x590 & ~x591 & ~x609 & ~x610 & ~x611 & ~x613 & ~x615 & ~x616 & ~x617 & ~x619 & ~x620 & ~x622 & ~x637 & ~x639 & ~x641 & ~x642 & ~x643 & ~x647 & ~x648 & ~x649 & ~x650 & ~x665 & ~x666 & ~x667 & ~x669 & ~x670 & ~x671 & ~x672 & ~x673 & ~x674 & ~x675 & ~x676 & ~x678 & ~x693 & ~x694 & ~x696 & ~x697 & ~x698 & ~x699 & ~x702 & ~x703 & ~x721 & ~x722 & ~x726 & ~x728 & ~x729 & ~x730 & ~x731 & ~x732 & ~x733 & ~x750 & ~x751 & ~x752 & ~x753 & ~x754 & ~x755 & ~x757 & ~x758 & ~x760 & ~x761 & ~x777 & ~x778 & ~x779 & ~x780 & ~x782;
assign c3100 =  x98 &  x124 &  x293 &  x343 &  x572 &  x740 & ~x19 & ~x25 & ~x146 & ~x163 & ~x173 & ~x197 & ~x230 & ~x309 & ~x311 & ~x395 & ~x415 & ~x474 & ~x480 & ~x530 & ~x589 & ~x591 & ~x611;
assign c3102 = ~x1 & ~x39 & ~x68 & ~x72 & ~x225 & ~x248 & ~x368 & ~x706;
assign c3104 =  x10 &  x573 &  x738 & ~x3 & ~x19 & ~x27 & ~x29 & ~x56 & ~x81 & ~x82 & ~x85 & ~x87 & ~x111 & ~x115 & ~x138 & ~x168 & ~x169 & ~x171 & ~x194 & ~x199 & ~x222 & ~x250 & ~x276 & ~x278 & ~x281 & ~x309 & ~x334 & ~x336 & ~x362 & ~x448 & ~x477 & ~x502 & ~x504 & ~x505 & ~x532 & ~x558 & ~x587 & ~x643 & ~x644 & ~x645 & ~x700 & ~x728 & ~x783;
assign c3106 = ~x77 & ~x80 & ~x88 & ~x113 & ~x140 & ~x144 & ~x163 & ~x173 & ~x249 & ~x273 & ~x306 & ~x311 & ~x362 & ~x365 & ~x380 & ~x444 & ~x448 & ~x504 & ~x533 & ~x594 & ~x617 & ~x648 & ~x664 & ~x668 & ~x693 & ~x704 & ~x705 & ~x706 & ~x729 & ~x734 & ~x756;
assign c3108 =  x299 &  x434 & ~x52 & ~x136 & ~x228 & ~x390 & ~x450 & ~x500 & ~x532 & ~x636 & ~x641 & ~x722 & ~x747;
assign c3110 =  x37 &  x39 &  x91 &  x92 &  x97 &  x236 &  x270 &  x686 &  x709 &  x737 & ~x0 & ~x164 & ~x172 & ~x220 & ~x255 & ~x279 & ~x307 & ~x420;
assign c3112 =  x11 &  x37 &  x94 &  x177 &  x235 & ~x112 & ~x142 & ~x191 & ~x198 & ~x199 & ~x221 & ~x223 & ~x252 & ~x256 & ~x276 & ~x305 & ~x339 & ~x477 & ~x615 & ~x645 & ~x670 & ~x723 & ~x752 & ~x760;
assign c3114 =  x98 &  x374 &  x524 &  x624 &  x691 &  x692 &  x707 & ~x136 & ~x167 & ~x306 & ~x780;
assign c3116 =  x517 & ~x5 & ~x51 & ~x55 & ~x60 & ~x82 & ~x86 & ~x106 & ~x107 & ~x111 & ~x112 & ~x113 & ~x162 & ~x164 & ~x166 & ~x168 & ~x170 & ~x191 & ~x193 & ~x196 & ~x199 & ~x218 & ~x223 & ~x229 & ~x247 & ~x254 & ~x284 & ~x298 & ~x307 & ~x326 & ~x333 & ~x337 & ~x361 & ~x366 & ~x395 & ~x417 & ~x418 & ~x422 & ~x424 & ~x445 & ~x452 & ~x473 & ~x502 & ~x505 & ~x506 & ~x508 & ~x558 & ~x559 & ~x560 & ~x561 & ~x588 & ~x591 & ~x616 & ~x646 & ~x671 & ~x672 & ~x676 & ~x694 & ~x700 & ~x725 & ~x727 & ~x728 & ~x730 & ~x752 & ~x780;
assign c3118 =  x216 &  x232 &  x741 & ~x0 & ~x1 & ~x8 & ~x20 & ~x21 & ~x22 & ~x24 & ~x25 & ~x26 & ~x28 & ~x29 & ~x30 & ~x51 & ~x52 & ~x53 & ~x55 & ~x57 & ~x81 & ~x82 & ~x83 & ~x85 & ~x86 & ~x105 & ~x106 & ~x107 & ~x108 & ~x114 & ~x136 & ~x138 & ~x139 & ~x142 & ~x143 & ~x165 & ~x168 & ~x169 & ~x170 & ~x192 & ~x196 & ~x197 & ~x198 & ~x200 & ~x252 & ~x253 & ~x254 & ~x255 & ~x256 & ~x276 & ~x277 & ~x278 & ~x279 & ~x280 & ~x281 & ~x282 & ~x283 & ~x284 & ~x303 & ~x308 & ~x332 & ~x336 & ~x338 & ~x340 & ~x360 & ~x361 & ~x363 & ~x366 & ~x367 & ~x390 & ~x391 & ~x393 & ~x394 & ~x417 & ~x418 & ~x420 & ~x423 & ~x444 & ~x445 & ~x446 & ~x448 & ~x449 & ~x451 & ~x471 & ~x472 & ~x474 & ~x476 & ~x478 & ~x506 & ~x529 & ~x531 & ~x532 & ~x533 & ~x537 & ~x555 & ~x557 & ~x558 & ~x559 & ~x565 & ~x566 & ~x585 & ~x589 & ~x590 & ~x612 & ~x613 & ~x614 & ~x616 & ~x618 & ~x619 & ~x621 & ~x637 & ~x638 & ~x640 & ~x642 & ~x645 & ~x650 & ~x665 & ~x667 & ~x668 & ~x672 & ~x673 & ~x674 & ~x675 & ~x676 & ~x677 & ~x693 & ~x694 & ~x697 & ~x699 & ~x700 & ~x702 & ~x704 & ~x721 & ~x722 & ~x724 & ~x726 & ~x727 & ~x730 & ~x756 & ~x758 & ~x778 & ~x781 & ~x782 & ~x783;
assign c3120 =  x325 & ~x0 & ~x25 & ~x33 & ~x111 & ~x115 & ~x168 & ~x195 & ~x204 & ~x220 & ~x222 & ~x224 & ~x228 & ~x248 & ~x249 & ~x250 & ~x277 & ~x282 & ~x307 & ~x308 & ~x332 & ~x336 & ~x343 & ~x361 & ~x365 & ~x394 & ~x395 & ~x398 & ~x414 & ~x424 & ~x452 & ~x471 & ~x472 & ~x473 & ~x474 & ~x479 & ~x503 & ~x507 & ~x528 & ~x531 & ~x535 & ~x558 & ~x583 & ~x584 & ~x587 & ~x614 & ~x619 & ~x620 & ~x647 & ~x726 & ~x755 & ~x757 & ~x759 & ~x779;
assign c3122 =  x46 &  x635 &  x663 & ~x0 & ~x55 & ~x87 & ~x227 & ~x248 & ~x252 & ~x278 & ~x316 & ~x423 & ~x473 & ~x502 & ~x529 & ~x559 & ~x612 & ~x615 & ~x647 & ~x671;
assign c3124 =  x235 &  x623 & ~x87 & ~x140 & ~x227 & ~x272 & ~x332 & ~x414 & ~x476;
assign c3126 =  x461 &  x491 & ~x1 & ~x5 & ~x10 & ~x31 & ~x87 & ~x106 & ~x118 & ~x145 & ~x222 & ~x247 & ~x277 & ~x312 & ~x400 & ~x423 & ~x500 & ~x512 & ~x534 & ~x535 & ~x556 & ~x563 & ~x647 & ~x697 & ~x733 & ~x750 & ~x756 & ~x777;
assign c3128 = ~x2 & ~x3 & ~x8 & ~x21 & ~x24 & ~x25 & ~x28 & ~x29 & ~x31 & ~x53 & ~x54 & ~x82 & ~x83 & ~x103 & ~x113 & ~x115 & ~x116 & ~x138 & ~x141 & ~x143 & ~x164 & ~x170 & ~x171 & ~x193 & ~x194 & ~x195 & ~x196 & ~x198 & ~x200 & ~x203 & ~x220 & ~x224 & ~x230 & ~x231 & ~x248 & ~x249 & ~x250 & ~x251 & ~x252 & ~x257 & ~x259 & ~x273 & ~x274 & ~x275 & ~x276 & ~x278 & ~x281 & ~x285 & ~x287 & ~x303 & ~x305 & ~x334 & ~x343 & ~x365 & ~x366 & ~x367 & ~x370 & ~x386 & ~x387 & ~x388 & ~x389 & ~x390 & ~x391 & ~x397 & ~x417 & ~x420 & ~x422 & ~x443 & ~x445 & ~x448 & ~x451 & ~x452 & ~x453 & ~x471 & ~x473 & ~x475 & ~x476 & ~x477 & ~x478 & ~x482 & ~x499 & ~x500 & ~x503 & ~x506 & ~x508 & ~x510 & ~x527 & ~x528 & ~x529 & ~x530 & ~x536 & ~x537 & ~x555 & ~x556 & ~x557 & ~x558 & ~x559 & ~x563 & ~x565 & ~x585 & ~x587 & ~x589 & ~x590 & ~x612 & ~x617 & ~x639 & ~x646 & ~x649 & ~x671 & ~x673 & ~x674 & ~x696 & ~x698 & ~x701 & ~x704 & ~x730 & ~x731 & ~x755 & ~x757 & ~x759 & ~x760 & ~x761 & ~x762 & ~x772 & ~x777 & ~x778 & ~x780;
assign c3130 =  x147 & ~x90 & ~x136 & ~x284 & ~x419 & ~x610 & ~x618 & ~x637 & ~x675;
assign c3132 = ~x78 & ~x79 & ~x87 & ~x163 & ~x171 & ~x172 & ~x206 & ~x227 & ~x234 & ~x288 & ~x289 & ~x316 & ~x329 & ~x343 & ~x344 & ~x357 & ~x358 & ~x364 & ~x386 & ~x444 & ~x469 & ~x558 & ~x648 & ~x676 & ~x696;
assign c3134 =  x460 & ~x116 & ~x170 & ~x173 & ~x221 & ~x270 & ~x276 & ~x317 & ~x364 & ~x390 & ~x473 & ~x499 & ~x508 & ~x734;
assign c3136 =  x37 &  x94 &  x206 & ~x0 & ~x2 & ~x3 & ~x5 & ~x8 & ~x13 & ~x14 & ~x21 & ~x22 & ~x23 & ~x25 & ~x26 & ~x27 & ~x28 & ~x29 & ~x30 & ~x31 & ~x32 & ~x52 & ~x53 & ~x54 & ~x55 & ~x56 & ~x57 & ~x58 & ~x59 & ~x60 & ~x79 & ~x80 & ~x81 & ~x82 & ~x83 & ~x84 & ~x86 & ~x87 & ~x88 & ~x107 & ~x108 & ~x109 & ~x110 & ~x112 & ~x113 & ~x115 & ~x116 & ~x135 & ~x136 & ~x137 & ~x139 & ~x140 & ~x141 & ~x142 & ~x143 & ~x144 & ~x164 & ~x165 & ~x166 & ~x168 & ~x169 & ~x170 & ~x171 & ~x192 & ~x193 & ~x194 & ~x195 & ~x196 & ~x197 & ~x198 & ~x199 & ~x220 & ~x221 & ~x222 & ~x223 & ~x224 & ~x225 & ~x226 & ~x227 & ~x247 & ~x249 & ~x250 & ~x251 & ~x252 & ~x253 & ~x254 & ~x255 & ~x275 & ~x276 & ~x277 & ~x278 & ~x279 & ~x281 & ~x282 & ~x283 & ~x304 & ~x305 & ~x306 & ~x307 & ~x308 & ~x309 & ~x310 & ~x311 & ~x332 & ~x333 & ~x334 & ~x335 & ~x336 & ~x337 & ~x338 & ~x339 & ~x360 & ~x361 & ~x363 & ~x364 & ~x365 & ~x366 & ~x368 & ~x389 & ~x390 & ~x391 & ~x392 & ~x393 & ~x394 & ~x417 & ~x418 & ~x419 & ~x420 & ~x421 & ~x423 & ~x444 & ~x445 & ~x449 & ~x450 & ~x451 & ~x474 & ~x475 & ~x476 & ~x477 & ~x478 & ~x479 & ~x501 & ~x502 & ~x503 & ~x504 & ~x505 & ~x506 & ~x507 & ~x528 & ~x529 & ~x530 & ~x531 & ~x532 & ~x534 & ~x535 & ~x558 & ~x559 & ~x560 & ~x561 & ~x562 & ~x585 & ~x586 & ~x587 & ~x588 & ~x589 & ~x590 & ~x615 & ~x616 & ~x618 & ~x642 & ~x643 & ~x644 & ~x645 & ~x646 & ~x647 & ~x671 & ~x673 & ~x674 & ~x699 & ~x700 & ~x701 & ~x725 & ~x726 & ~x727 & ~x728 & ~x729 & ~x730 & ~x753 & ~x754 & ~x755 & ~x756 & ~x757 & ~x758 & ~x759 & ~x760 & ~x761 & ~x762 & ~x777 & ~x778 & ~x779 & ~x780 & ~x781 & ~x782 & ~x783;
assign c3138 =  x120 & ~x2 & ~x26 & ~x27 & ~x31 & ~x58 & ~x60 & ~x61 & ~x81 & ~x85 & ~x107 & ~x110 & ~x113 & ~x114 & ~x116 & ~x117 & ~x141 & ~x169 & ~x171 & ~x173 & ~x190 & ~x196 & ~x198 & ~x199 & ~x200 & ~x220 & ~x227 & ~x248 & ~x249 & ~x253 & ~x256 & ~x277 & ~x334 & ~x337 & ~x338 & ~x361 & ~x362 & ~x390 & ~x418 & ~x449 & ~x476 & ~x503 & ~x504 & ~x507 & ~x557 & ~x558 & ~x559 & ~x586 & ~x590 & ~x615 & ~x726 & ~x752 & ~x758 & ~x777 & ~x778 & ~x779 & ~x780;
assign c3140 =  x41 &  x65 &  x120 &  x180 &  x239 &  x259 &  x322 &  x347 &  x403 &  x433 &  x630 &  x685 &  x745 & ~x26 & ~x29 & ~x50 & ~x60 & ~x82 & ~x90 & ~x118 & ~x195 & ~x640 & ~x649 & ~x674 & ~x696 & ~x702;
assign c3142 = ~x6 & ~x9 & ~x78 & ~x83 & ~x97 & ~x115 & ~x145 & ~x166 & ~x168 & ~x197 & ~x220 & ~x222 & ~x249 & ~x278 & ~x280 & ~x468 & ~x475 & ~x503 & ~x507 & ~x508 & ~x556 & ~x563 & ~x585 & ~x611 & ~x621 & ~x647 & ~x668 & ~x671 & ~x704 & ~x723 & ~x755 & ~x776;
assign c3144 =  x517 & ~x5 & ~x27 & ~x87 & ~x125 & ~x139 & ~x163 & ~x247 & ~x249 & ~x253 & ~x306 & ~x311 & ~x340 & ~x393 & ~x447 & ~x481 & ~x615 & ~x763;
assign c3146 =  x68 &  x124 &  x126 &  x128 &  x236 &  x238 &  x295 &  x323 &  x348 &  x378 &  x405 &  x437 &  x461 &  x462 &  x491 &  x516 &  x548 &  x571 &  x572 &  x577 &  x686 & ~x0 & ~x29 & ~x48 & ~x64 & ~x76 & ~x77 & ~x82 & ~x88 & ~x90 & ~x106 & ~x108 & ~x161 & ~x169 & ~x189 & ~x202 & ~x222 & ~x226 & ~x229 & ~x246 & ~x258 & ~x274 & ~x279 & ~x309 & ~x314 & ~x336 & ~x363 & ~x368 & ~x397 & ~x415 & ~x421 & ~x451 & ~x503 & ~x528 & ~x560 & ~x561 & ~x585 & ~x611 & ~x618 & ~x640 & ~x646 & ~x647 & ~x674 & ~x675 & ~x699 & ~x756 & ~x761 & ~x780 & ~x781;
assign c3148 = ~x3 & ~x5 & ~x110 & ~x111 & ~x115 & ~x188 & ~x214 & ~x242 & ~x259 & ~x260 & ~x270 & ~x271 & ~x273 & ~x304 & ~x327 & ~x329 & ~x372 & ~x397 & ~x412 & ~x413 & ~x451 & ~x455 & ~x479 & ~x497 & ~x537 & ~x590 & ~x591 & ~x610 & ~x639 & ~x671 & ~x704 & ~x762;
assign c3150 =  x536;
assign c3152 =  x261 & ~x9 & ~x51 & ~x116 & ~x200 & ~x201 & ~x228 & ~x247 & ~x276 & ~x313 & ~x340 & ~x346 & ~x394 & ~x443 & ~x475 & ~x762 & ~x779;
assign c3154 =  x40 &  x122 &  x155 &  x208 &  x351 &  x433 &  x434 &  x520 &  x545 &  x601 &  x658 &  x685 &  x742 &  x744 &  x745 & ~x6 & ~x20 & ~x21 & ~x30 & ~x32 & ~x49 & ~x52 & ~x62 & ~x76 & ~x80 & ~x84 & ~x85 & ~x105 & ~x117 & ~x164 & ~x167 & ~x190 & ~x195 & ~x219 & ~x250 & ~x256 & ~x258 & ~x285 & ~x306 & ~x308 & ~x312 & ~x333 & ~x336 & ~x341 & ~x359 & ~x363 & ~x366 & ~x389 & ~x392 & ~x394 & ~x425 & ~x446 & ~x450 & ~x535 & ~x559 & ~x590 & ~x592 & ~x612 & ~x619 & ~x641 & ~x646 & ~x649 & ~x670 & ~x679 & ~x730 & ~x781;
assign c3156 =  x568 &  x636 &  x734 &  x735 &  x736 & ~x30 & ~x82 & ~x225 & ~x250 & ~x305 & ~x332 & ~x530 & ~x728;
assign c3158 =  x311;
assign c3160 = ~x172 & ~x230 & ~x286 & ~x476 & ~x493 & ~x556 & ~x604;
assign c3162 =  x184 &  x216 &  x489 &  x490 &  x709 &  x774 & ~x78 & ~x117 & ~x163 & ~x170 & ~x173 & ~x557 & ~x674 & ~x675 & ~x676 & ~x678 & ~x730;
assign c3164 =  x354 &  x719 & ~x141 & ~x228 & ~x231 & ~x272 & ~x281 & ~x305 & ~x307 & ~x386;
assign c3166 =  x42 &  x489 & ~x4 & ~x6 & ~x17 & ~x58 & ~x226 & ~x249 & ~x254 & ~x306 & ~x354 & ~x472 & ~x502;
assign c3168 = ~x4 & ~x6 & ~x10 & ~x22 & ~x29 & ~x49 & ~x55 & ~x61 & ~x62 & ~x81 & ~x90 & ~x108 & ~x111 & ~x117 & ~x135 & ~x136 & ~x143 & ~x173 & ~x201 & ~x213 & ~x221 & ~x223 & ~x251 & ~x252 & ~x253 & ~x254 & ~x258 & ~x274 & ~x275 & ~x302 & ~x303 & ~x311 & ~x334 & ~x336 & ~x338 & ~x339 & ~x340 & ~x360 & ~x365 & ~x366 & ~x387 & ~x416 & ~x419 & ~x443 & ~x446 & ~x448 & ~x481 & ~x499 & ~x507 & ~x526 & ~x591 & ~x592 & ~x613 & ~x616 & ~x642 & ~x664 & ~x665 & ~x667 & ~x677 & ~x703 & ~x704 & ~x705 & ~x706 & ~x727 & ~x728 & ~x732 & ~x735 & ~x749 & ~x762 & ~x780;
assign c3170 =  x70 &  x95 &  x97 &  x152 &  x153 &  x156 &  x182 &  x266 &  x295 &  x348 &  x378 &  x460 &  x463 &  x465 &  x489 &  x491 &  x547 &  x574 &  x602 &  x627 &  x628 &  x655 &  x689 & ~x0 & ~x23 & ~x50 & ~x51 & ~x79 & ~x82 & ~x106 & ~x108 & ~x115 & ~x166 & ~x170 & ~x194 & ~x248 & ~x254 & ~x278 & ~x281 & ~x307 & ~x309 & ~x361 & ~x396 & ~x397 & ~x423 & ~x424 & ~x444 & ~x450 & ~x452 & ~x453 & ~x473 & ~x475 & ~x478 & ~x480 & ~x497 & ~x503 & ~x559 & ~x560 & ~x588 & ~x589 & ~x614 & ~x617 & ~x619 & ~x666 & ~x729 & ~x777;
assign c3172 =  x518 &  x630 & ~x8 & ~x25 & ~x51 & ~x88 & ~x93 & ~x168 & ~x247 & ~x251 & ~x259 & ~x361 & ~x388 & ~x397 & ~x399 & ~x444 & ~x473 & ~x498 & ~x591 & ~x614 & ~x620 & ~x671 & ~x726;
assign c3174 =  x46 &  x74 &  x91 &  x737 & ~x3 & ~x8 & ~x9 & ~x15 & ~x86 & ~x171 & ~x196 & ~x307 & ~x309 & ~x447 & ~x588;
assign c3176 =  x478;
assign c3178 =  x606 & ~x221 & ~x271 & ~x699 & ~x779;
assign c3180 =  x65 &  x120 &  x404 &  x458 &  x602 &  x631 & ~x3 & ~x25 & ~x27 & ~x29 & ~x31 & ~x35 & ~x48 & ~x56 & ~x78 & ~x81 & ~x82 & ~x84 & ~x106 & ~x107 & ~x115 & ~x141 & ~x144 & ~x163 & ~x165 & ~x192 & ~x198 & ~x199 & ~x220 & ~x224 & ~x286 & ~x304 & ~x307 & ~x313 & ~x314 & ~x334 & ~x389 & ~x390 & ~x396 & ~x448 & ~x451 & ~x481 & ~x503 & ~x529 & ~x533 & ~x613 & ~x614 & ~x618 & ~x642 & ~x645 & ~x647 & ~x695 & ~x702 & ~x723 & ~x728 & ~x732 & ~x750 & ~x752 & ~x758 & ~x780 & ~x782;
assign c3182 =  x45 &  x665;
assign c3184 = ~x35 & ~x77 & ~x78 & ~x111 & ~x163 & ~x234 & ~x303 & ~x332 & ~x373 & ~x389 & ~x390 & ~x442 & ~x452 & ~x528 & ~x563 & ~x652 & ~x694 & ~x722 & ~x734;
assign c3186 =  x10 &  x67 &  x69 &  x93 &  x349 &  x522 &  x575 &  x712 &  x714 & ~x58 & ~x82 & ~x85 & ~x141 & ~x169 & ~x200 & ~x224 & ~x252 & ~x280 & ~x558 & ~x699 & ~x759;
assign c3188 =  x350 &  x486 & ~x145 & ~x270 & ~x615 & ~x756;
assign c3190 = ~x462 & ~x599;
assign c3192 =  x322 &  x323 &  x714 & ~x298;
assign c3194 =  x396 & ~x648;
assign c3196 =  x272 &  x288 & ~x1 & ~x5 & ~x6 & ~x32 & ~x35 & ~x48 & ~x77 & ~x83 & ~x87 & ~x89 & ~x112 & ~x118 & ~x134 & ~x172 & ~x191 & ~x194 & ~x199 & ~x200 & ~x218 & ~x219 & ~x223 & ~x226 & ~x228 & ~x229 & ~x254 & ~x256 & ~x276 & ~x278 & ~x281 & ~x303 & ~x309 & ~x310 & ~x312 & ~x340 & ~x359 & ~x362 & ~x364 & ~x389 & ~x419 & ~x450 & ~x451 & ~x474 & ~x479 & ~x502 & ~x505 & ~x531 & ~x557 & ~x566 & ~x586 & ~x616 & ~x617 & ~x639 & ~x640 & ~x646 & ~x651 & ~x673 & ~x695 & ~x699 & ~x703 & ~x706 & ~x707 & ~x726 & ~x730 & ~x734 & ~x754 & ~x761 & ~x783;
assign c3198 =  x39 &  x47 &  x742 & ~x23 & ~x58 & ~x85 & ~x86 & ~x114 & ~x139 & ~x165 & ~x166 & ~x171 & ~x192 & ~x193 & ~x220 & ~x224 & ~x248 & ~x249 & ~x251 & ~x276 & ~x277 & ~x304 & ~x306 & ~x332 & ~x333 & ~x336 & ~x390 & ~x391 & ~x395 & ~x419 & ~x420 & ~x446 & ~x448 & ~x473 & ~x474 & ~x476 & ~x477 & ~x502 & ~x530 & ~x563 & ~x591 & ~x610 & ~x616 & ~x668 & ~x674 & ~x699 & ~x700 & ~x702 & ~x755 & ~x758 & ~x762 & ~x763;
assign c3200 = ~x28 & ~x56 & ~x69 & ~x144 & ~x200 & ~x391 & ~x429 & ~x505 & ~x701 & ~x761;
assign c3202 =  x300 &  x442 &  x736 &  x743 & ~x82 & ~x167 & ~x280 & ~x303 & ~x331 & ~x388 & ~x533;
assign c3204 =  x302 & ~x23 & ~x52 & ~x54 & ~x134 & ~x166 & ~x225 & ~x248 & ~x585 & ~x619 & ~x639 & ~x667 & ~x697 & ~x723 & ~x724 & ~x760;
assign c3206 = ~x96 & ~x270 & ~x372 & ~x387 & ~x699;
assign c3208 =  x155 &  x517 & ~x0 & ~x2 & ~x6 & ~x10 & ~x17 & ~x19 & ~x37 & ~x46 & ~x47 & ~x49 & ~x78 & ~x87 & ~x111 & ~x134 & ~x141 & ~x145 & ~x164 & ~x165 & ~x174 & ~x190 & ~x194 & ~x219 & ~x229 & ~x230 & ~x254 & ~x275 & ~x282 & ~x283 & ~x307 & ~x330 & ~x334 & ~x341 & ~x342 & ~x360 & ~x367 & ~x368 & ~x386 & ~x419 & ~x446 & ~x481 & ~x500 & ~x509 & ~x530 & ~x557 & ~x564 & ~x565 & ~x589 & ~x617 & ~x618 & ~x622 & ~x647 & ~x651 & ~x666 & ~x669 & ~x671 & ~x677 & ~x707 & ~x723 & ~x750 & ~x757 & ~x761 & ~x782;
assign c3210 =  x433 &  x713 & ~x19 & ~x59 & ~x141 & ~x166 & ~x190 & ~x191 & ~x195 & ~x250 & ~x256 & ~x275 & ~x333 & ~x338 & ~x361 & ~x388 & ~x421 & ~x426 & ~x440 & ~x444 & ~x445 & ~x469 & ~x480 & ~x506 & ~x509 & ~x535 & ~x537 & ~x557 & ~x561 & ~x589 & ~x618 & ~x647 & ~x755 & ~x773;
assign c3212 =  x72 &  x100 &  x122 &  x128 &  x153 &  x266 &  x294 &  x489 &  x519 &  x573 &  x686 & ~x138 & ~x259 & ~x272 & ~x307 & ~x314 & ~x362 & ~x415 & ~x420 & ~x425 & ~x534 & ~x564 & ~x617 & ~x641;
assign c3214 =  x69 &  x73 &  x95 &  x156 &  x292 &  x375 &  x462 &  x546 &  x685 &  x742 &  x744 & ~x5 & ~x28 & ~x29 & ~x62 & ~x78 & ~x81 & ~x135 & ~x138 & ~x223 & ~x283 & ~x341 & ~x364 & ~x365 & ~x425 & ~x426 & ~x443 & ~x453 & ~x473 & ~x478 & ~x527 & ~x529 & ~x566 & ~x581 & ~x593 & ~x613 & ~x621 & ~x668 & ~x698 & ~x749 & ~x781;
assign c3216 =  x154 &  x575 &  x662 & ~x8 & ~x28 & ~x85 & ~x249 & ~x250 & ~x278 & ~x289 & ~x338 & ~x448 & ~x564 & ~x672 & ~x729 & ~x757;
assign c3218 =  x210 &  x238 &  x496 &  x691 &  x694 & ~x14 & ~x20 & ~x27 & ~x57 & ~x85 & ~x139 & ~x221 & ~x561;
assign c3220 =  x41 &  x42 & ~x0 & ~x19 & ~x26 & ~x27 & ~x48 & ~x58 & ~x61 & ~x77 & ~x84 & ~x107 & ~x111 & ~x115 & ~x171 & ~x172 & ~x173 & ~x194 & ~x199 & ~x220 & ~x257 & ~x270 & ~x275 & ~x286 & ~x302 & ~x305 & ~x307 & ~x335 & ~x342 & ~x393 & ~x398 & ~x415 & ~x420 & ~x425 & ~x447 & ~x453 & ~x472 & ~x473 & ~x482 & ~x498 & ~x499 & ~x526 & ~x528 & ~x565 & ~x566 & ~x594 & ~x621 & ~x640 & ~x645 & ~x649 & ~x720 & ~x725 & ~x750 & ~x756 & ~x761 & ~x776 & ~x779;
assign c3222 =  x232 &  x321 &  x489 &  x601 &  x659 &  x713 &  x741 &  x766 & ~x6 & ~x19 & ~x78 & ~x85 & ~x107 & ~x196 & ~x197 & ~x360 & ~x362 & ~x388 & ~x423 & ~x480 & ~x503 & ~x531 & ~x589 & ~x649 & ~x667 & ~x679 & ~x695 & ~x704 & ~x733 & ~x762;
assign c3224 =  x40 &  x42 &  x99 &  x100 &  x128 &  x209 &  x210 &  x295 &  x321 &  x348 &  x350 &  x375 &  x377 &  x436 &  x461 &  x462 &  x463 &  x464 &  x487 &  x488 &  x489 &  x491 &  x517 &  x518 &  x519 &  x520 &  x521 &  x543 &  x547 &  x571 &  x574 &  x575 &  x577 &  x601 &  x603 &  x605 &  x627 &  x631 &  x658 &  x661 & ~x1 & ~x3 & ~x4 & ~x5 & ~x7 & ~x8 & ~x25 & ~x29 & ~x30 & ~x32 & ~x35 & ~x48 & ~x50 & ~x51 & ~x53 & ~x55 & ~x57 & ~x58 & ~x59 & ~x60 & ~x78 & ~x82 & ~x87 & ~x106 & ~x107 & ~x108 & ~x109 & ~x115 & ~x116 & ~x138 & ~x141 & ~x161 & ~x162 & ~x163 & ~x164 & ~x167 & ~x170 & ~x171 & ~x174 & ~x190 & ~x192 & ~x193 & ~x200 & ~x201 & ~x202 & ~x217 & ~x219 & ~x221 & ~x224 & ~x226 & ~x227 & ~x247 & ~x251 & ~x255 & ~x256 & ~x276 & ~x277 & ~x280 & ~x281 & ~x303 & ~x307 & ~x308 & ~x332 & ~x334 & ~x340 & ~x358 & ~x361 & ~x362 & ~x365 & ~x368 & ~x386 & ~x388 & ~x389 & ~x390 & ~x393 & ~x415 & ~x420 & ~x421 & ~x445 & ~x447 & ~x451 & ~x452 & ~x453 & ~x470 & ~x501 & ~x507 & ~x509 & ~x527 & ~x535 & ~x556 & ~x557 & ~x564 & ~x584 & ~x585 & ~x588 & ~x589 & ~x593 & ~x610 & ~x614 & ~x615 & ~x617 & ~x618 & ~x619 & ~x620 & ~x642 & ~x643 & ~x644 & ~x645 & ~x646 & ~x665 & ~x669 & ~x670 & ~x672 & ~x697 & ~x703 & ~x705 & ~x734 & ~x750 & ~x753 & ~x754 & ~x758 & ~x759 & ~x760 & ~x780 & ~x781;
assign c3226 =  x122 & ~x1 & ~x7 & ~x13 & ~x14 & ~x25 & ~x26 & ~x43 & ~x48 & ~x112 & ~x227 & ~x254 & ~x559 & ~x703 & ~x780;
assign c3228 =  x37 &  x45 &  x46 &  x384 &  x663 &  x737 & ~x3 & ~x111 & ~x193 & ~x197 & ~x198 & ~x200 & ~x221 & ~x304 & ~x305 & ~x309 & ~x417 & ~x418 & ~x476 & ~x504 & ~x530 & ~x586 & ~x758 & ~x777;
assign c3230 =  x517 &  x740 &  x770 & ~x7 & ~x49 & ~x50 & ~x142 & ~x169 & ~x249 & ~x251 & ~x254 & ~x276 & ~x277 & ~x370 & ~x507 & ~x553 & ~x564 & ~x586 & ~x596 & ~x623 & ~x667 & ~x695;
assign c3232 = ~x0 & ~x2 & ~x4 & ~x5 & ~x7 & ~x8 & ~x17 & ~x18 & ~x19 & ~x21 & ~x22 & ~x23 & ~x24 & ~x25 & ~x27 & ~x28 & ~x29 & ~x30 & ~x31 & ~x33 & ~x34 & ~x50 & ~x52 & ~x53 & ~x54 & ~x55 & ~x56 & ~x57 & ~x60 & ~x80 & ~x81 & ~x83 & ~x87 & ~x88 & ~x89 & ~x109 & ~x111 & ~x113 & ~x115 & ~x136 & ~x137 & ~x139 & ~x142 & ~x143 & ~x144 & ~x145 & ~x164 & ~x168 & ~x169 & ~x171 & ~x173 & ~x192 & ~x194 & ~x195 & ~x196 & ~x197 & ~x198 & ~x199 & ~x200 & ~x220 & ~x221 & ~x222 & ~x224 & ~x226 & ~x227 & ~x248 & ~x249 & ~x252 & ~x254 & ~x255 & ~x257 & ~x258 & ~x275 & ~x276 & ~x277 & ~x279 & ~x280 & ~x281 & ~x282 & ~x288 & ~x299 & ~x303 & ~x304 & ~x305 & ~x307 & ~x308 & ~x309 & ~x313 & ~x316 & ~x332 & ~x333 & ~x334 & ~x335 & ~x337 & ~x338 & ~x339 & ~x341 & ~x356 & ~x359 & ~x361 & ~x364 & ~x366 & ~x367 & ~x368 & ~x386 & ~x388 & ~x389 & ~x390 & ~x391 & ~x392 & ~x393 & ~x395 & ~x396 & ~x415 & ~x416 & ~x417 & ~x420 & ~x423 & ~x424 & ~x425 & ~x444 & ~x445 & ~x447 & ~x449 & ~x451 & ~x453 & ~x474 & ~x478 & ~x479 & ~x497 & ~x498 & ~x500 & ~x502 & ~x503 & ~x504 & ~x505 & ~x506 & ~x507 & ~x510 & ~x527 & ~x528 & ~x531 & ~x532 & ~x533 & ~x534 & ~x535 & ~x536 & ~x538 & ~x554 & ~x557 & ~x559 & ~x560 & ~x561 & ~x563 & ~x565 & ~x584 & ~x586 & ~x587 & ~x588 & ~x611 & ~x613 & ~x615 & ~x618 & ~x619 & ~x638 & ~x643 & ~x644 & ~x646 & ~x647 & ~x668 & ~x669 & ~x671 & ~x672 & ~x676 & ~x695 & ~x696 & ~x698 & ~x700 & ~x701 & ~x702 & ~x703 & ~x704 & ~x723 & ~x725 & ~x727 & ~x729 & ~x731 & ~x733 & ~x751 & ~x752 & ~x753 & ~x758 & ~x761 & ~x762 & ~x777 & ~x779 & ~x781 & ~x782 & ~x783;
assign c3234 =  x95 &  x96 &  x126 &  x127 &  x206 &  x209 &  x318 &  x319 &  x348 &  x379 &  x406 &  x458 &  x513 &  x515 &  x546 &  x681 &  x715 & ~x1 & ~x24 & ~x36 & ~x48 & ~x76 & ~x81 & ~x83 & ~x86 & ~x90 & ~x104 & ~x113 & ~x140 & ~x146 & ~x196 & ~x256 & ~x278 & ~x281 & ~x282 & ~x305 & ~x313 & ~x340 & ~x341 & ~x365 & ~x499 & ~x557 & ~x559 & ~x583 & ~x591 & ~x615 & ~x616 & ~x699 & ~x781;
assign c3236 =  x65 &  x68 &  x98 &  x127 &  x434 &  x460 & ~x28 & ~x62 & ~x90 & ~x140 & ~x144 & ~x197 & ~x226 & ~x227 & ~x230 & ~x247 & ~x252 & ~x254 & ~x257 & ~x280 & ~x306 & ~x362 & ~x394 & ~x415 & ~x416 & ~x480 & ~x503 & ~x560 & ~x584;
assign c3238 =  x434 &  x490 &  x602 &  x605 & ~x9 & ~x26 & ~x77 & ~x82 & ~x135 & ~x142 & ~x146 & ~x192 & ~x250 & ~x306 & ~x390 & ~x443 & ~x446 & ~x526 & ~x538 & ~x563 & ~x616 & ~x623 & ~x640 & ~x646 & ~x648 & ~x678 & ~x704 & ~x723 & ~x728;
assign c3240 = ~x0 & ~x8 & ~x18 & ~x20 & ~x24 & ~x32 & ~x33 & ~x50 & ~x52 & ~x59 & ~x77 & ~x78 & ~x85 & ~x87 & ~x107 & ~x111 & ~x114 & ~x115 & ~x117 & ~x135 & ~x136 & ~x137 & ~x138 & ~x141 & ~x142 & ~x145 & ~x163 & ~x164 & ~x168 & ~x173 & ~x201 & ~x218 & ~x219 & ~x220 & ~x223 & ~x228 & ~x229 & ~x248 & ~x251 & ~x253 & ~x254 & ~x276 & ~x280 & ~x284 & ~x304 & ~x305 & ~x307 & ~x309 & ~x310 & ~x334 & ~x335 & ~x336 & ~x338 & ~x361 & ~x394 & ~x415 & ~x416 & ~x417 & ~x418 & ~x421 & ~x422 & ~x425 & ~x451 & ~x473 & ~x476 & ~x477 & ~x500 & ~x501 & ~x504 & ~x506 & ~x508 & ~x531 & ~x536 & ~x542 & ~x556 & ~x557 & ~x564 & ~x587 & ~x589 & ~x593 & ~x610 & ~x613 & ~x614 & ~x618 & ~x619 & ~x620 & ~x639 & ~x644 & ~x671 & ~x672 & ~x673 & ~x674 & ~x694 & ~x696 & ~x698 & ~x701 & ~x702 & ~x703 & ~x704 & ~x723 & ~x725 & ~x728 & ~x753 & ~x760 & ~x761 & ~x762 & ~x763 & ~x777 & ~x778 & ~x779 & ~x780 & ~x781 & ~x782;
assign c3242 =  x36 &  x42 & ~x28 & ~x332 & ~x335;
assign c3244 =  x127 &  x128 &  x182 &  x352 &  x406 &  x490 &  x493 &  x515 &  x548 &  x572 & ~x2 & ~x3 & ~x5 & ~x25 & ~x27 & ~x28 & ~x32 & ~x59 & ~x79 & ~x89 & ~x143 & ~x163 & ~x167 & ~x194 & ~x195 & ~x200 & ~x220 & ~x282 & ~x308 & ~x332 & ~x334 & ~x336 & ~x365 & ~x392 & ~x421 & ~x472 & ~x473 & ~x478 & ~x501 & ~x506 & ~x512 & ~x530 & ~x588 & ~x615 & ~x669 & ~x670 & ~x695 & ~x697 & ~x704 & ~x734 & ~x762 & ~x780;
assign c3246 =  x46 &  x174 &  x182 &  x658 &  x736 & ~x168 & ~x197 & ~x762;
assign c3248 =  x271 &  x545 &  x546 & ~x5 & ~x6 & ~x20 & ~x21 & ~x23 & ~x31 & ~x52 & ~x56 & ~x58 & ~x86 & ~x87 & ~x107 & ~x108 & ~x109 & ~x117 & ~x138 & ~x139 & ~x146 & ~x162 & ~x163 & ~x164 & ~x165 & ~x196 & ~x199 & ~x200 & ~x220 & ~x222 & ~x223 & ~x224 & ~x225 & ~x226 & ~x228 & ~x254 & ~x276 & ~x277 & ~x278 & ~x280 & ~x282 & ~x304 & ~x305 & ~x309 & ~x310 & ~x331 & ~x335 & ~x336 & ~x339 & ~x361 & ~x362 & ~x390 & ~x415 & ~x416 & ~x425 & ~x426 & ~x443 & ~x446 & ~x448 & ~x449 & ~x451 & ~x452 & ~x471 & ~x476 & ~x499 & ~x502 & ~x503 & ~x506 & ~x509 & ~x531 & ~x532 & ~x533 & ~x534 & ~x552 & ~x562 & ~x565 & ~x580 & ~x584 & ~x586 & ~x590 & ~x608 & ~x611 & ~x640 & ~x643 & ~x644 & ~x666 & ~x667 & ~x669 & ~x677 & ~x678 & ~x694 & ~x697 & ~x699 & ~x706 & ~x722 & ~x723 & ~x726 & ~x727 & ~x731 & ~x734 & ~x749 & ~x755 & ~x757 & ~x760 & ~x761 & ~x762 & ~x778 & ~x781 & ~x783;
assign c3250 =  x634 & ~x14 & ~x86 & ~x121 & ~x413 & ~x427;
assign c3252 =  x433 &  x654 & ~x4 & ~x33 & ~x51 & ~x53 & ~x85 & ~x108 & ~x109 & ~x219 & ~x220 & ~x305 & ~x317 & ~x364 & ~x390 & ~x477 & ~x532 & ~x667 & ~x699 & ~x777 & ~x779 & ~x783;
assign c3254 =  x132 &  x148 &  x741 &  x743 & ~x9 & ~x20 & ~x24 & ~x31 & ~x54 & ~x107 & ~x112 & ~x138 & ~x139 & ~x196 & ~x197 & ~x223 & ~x228 & ~x253 & ~x255 & ~x257 & ~x280 & ~x282 & ~x284 & ~x305 & ~x306 & ~x309 & ~x312 & ~x332 & ~x340 & ~x361 & ~x365 & ~x368 & ~x393 & ~x396 & ~x417 & ~x421 & ~x443 & ~x445 & ~x449 & ~x452 & ~x500 & ~x501 & ~x504 & ~x531 & ~x558 & ~x562 & ~x565 & ~x585 & ~x587 & ~x612 & ~x617 & ~x639 & ~x645 & ~x647 & ~x674 & ~x700 & ~x754 & ~x760 & ~x779;
assign c3256 = ~x57 & ~x71 & ~x172 & ~x222 & ~x310 & ~x335 & ~x338 & ~x416 & ~x419 & ~x423 & ~x492 & ~x530 & ~x778 & ~x780;
assign c3258 =  x11 &  x40 &  x41 &  x44 &  x47 &  x712 & ~x28 & ~x55 & ~x87 & ~x109 & ~x112 & ~x115 & ~x221 & ~x227 & ~x281 & ~x304 & ~x309 & ~x334 & ~x340 & ~x363 & ~x390 & ~x396 & ~x448 & ~x472 & ~x502 & ~x529 & ~x530 & ~x587 & ~x615 & ~x647 & ~x673 & ~x676 & ~x697 & ~x702 & ~x704 & ~x723 & ~x727 & ~x729 & ~x757;
assign c3260 =  x180 &  x319 &  x405 &  x430 & ~x1 & ~x5 & ~x7 & ~x22 & ~x23 & ~x52 & ~x56 & ~x58 & ~x84 & ~x85 & ~x87 & ~x108 & ~x111 & ~x113 & ~x196 & ~x224 & ~x279 & ~x306 & ~x327 & ~x335 & ~x364 & ~x367 & ~x421 & ~x422 & ~x449 & ~x476 & ~x477 & ~x503 & ~x504 & ~x556 & ~x564 & ~x583 & ~x587 & ~x592 & ~x612 & ~x618 & ~x619 & ~x647 & ~x674 & ~x703 & ~x729 & ~x731 & ~x752 & ~x754 & ~x757 & ~x759 & ~x760;
assign c3262 =  x21;
assign c3264 =  x74 &  x356 &  x459 & ~x2 & ~x4 & ~x8 & ~x20 & ~x49 & ~x86 & ~x87 & ~x89 & ~x137 & ~x144 & ~x164 & ~x165 & ~x169 & ~x285 & ~x307 & ~x310 & ~x331 & ~x420 & ~x424 & ~x477 & ~x479 & ~x531 & ~x558 & ~x563 & ~x594 & ~x609 & ~x619 & ~x763 & ~x781;
assign c3266 =  x75 & ~x0 & ~x4 & ~x5 & ~x25 & ~x29 & ~x51 & ~x53 & ~x57 & ~x58 & ~x60 & ~x79 & ~x89 & ~x111 & ~x112 & ~x113 & ~x114 & ~x116 & ~x136 & ~x137 & ~x138 & ~x141 & ~x142 & ~x165 & ~x168 & ~x169 & ~x171 & ~x194 & ~x196 & ~x223 & ~x225 & ~x252 & ~x253 & ~x254 & ~x280 & ~x282 & ~x309 & ~x334 & ~x362 & ~x390 & ~x419 & ~x450 & ~x474 & ~x475 & ~x476 & ~x503 & ~x531 & ~x532 & ~x534 & ~x559 & ~x560 & ~x561 & ~x564 & ~x587 & ~x588 & ~x592 & ~x593 & ~x613 & ~x614 & ~x618 & ~x620 & ~x621 & ~x624 & ~x644 & ~x651 & ~x672 & ~x701 & ~x729 & ~x732 & ~x757 & ~x761 & ~x764 & ~x778 & ~x779 & ~x781;
assign c3268 = ~x262 & ~x371 & ~x427 & ~x455 & ~x503 & ~x510 & ~x525 & ~x567 & ~x596 & ~x775 & ~x777;
assign c3270 =  x210 &  x211 &  x434 &  x546 &  x549 &  x578 &  x633 & ~x30 & ~x55 & ~x110 & ~x115 & ~x232 & ~x363 & ~x417 & ~x423 & ~x700 & ~x727 & ~x781;
assign c3272 =  x389;
assign c3274 =  x264 &  x265 &  x653 & ~x3 & ~x56 & ~x193 & ~x204 & ~x226 & ~x248 & ~x303 & ~x386 & ~x451 & ~x471 & ~x588 & ~x618 & ~x753;
assign c3276 =  x152 &  x290 &  x348 &  x380 &  x433 &  x462 &  x486 & ~x25 & ~x26 & ~x170 & ~x260 & ~x420 & ~x558 & ~x699 & ~x757;
assign c3278 = ~x237 & ~x334 & ~x359 & ~x530 & ~x652 & ~x734;
assign c3280 =  x245 &  x601 & ~x0 & ~x21 & ~x22 & ~x24 & ~x26 & ~x28 & ~x34 & ~x55 & ~x60 & ~x83 & ~x84 & ~x134 & ~x140 & ~x143 & ~x163 & ~x171 & ~x173 & ~x191 & ~x193 & ~x195 & ~x201 & ~x228 & ~x256 & ~x282 & ~x362 & ~x393 & ~x473 & ~x474 & ~x476 & ~x556 & ~x586 & ~x592 & ~x615 & ~x620 & ~x640 & ~x650 & ~x677 & ~x695 & ~x702 & ~x728 & ~x731 & ~x758 & ~x778 & ~x782;
assign c3282 =  x11 &  x16 &  x37 & ~x307 & ~x647 & ~x672 & ~x675 & ~x783;
assign c3284 =  x63 &  x537 &  x567;
assign c3286 = ~x55 & ~x73 & ~x80 & ~x164 & ~x165 & ~x359 & ~x429 & ~x444 & ~x446 & ~x500 & ~x560 & ~x761;
assign c3288 =  x737 & ~x3 & ~x8 & ~x14 & ~x23 & ~x24 & ~x50 & ~x54 & ~x57 & ~x87 & ~x159 & ~x220 & ~x222 & ~x226 & ~x229 & ~x231 & ~x245 & ~x247 & ~x259 & ~x275 & ~x280 & ~x285 & ~x305 & ~x307 & ~x336 & ~x359 & ~x362 & ~x369 & ~x388 & ~x397 & ~x453 & ~x564 & ~x615 & ~x618 & ~x619 & ~x674 & ~x675 & ~x780;
assign c3290 =  x37 &  x38 &  x45 &  x133 &  x736 &  x738 & ~x27 & ~x55 & ~x112 & ~x141 & ~x167 & ~x225 & ~x248 & ~x256 & ~x276 & ~x280 & ~x310 & ~x361 & ~x362 & ~x392 & ~x504 & ~x506 & ~x557 & ~x560 & ~x614 & ~x781 & ~x782;
assign c3292 = ~x0 & ~x8 & ~x19 & ~x22 & ~x29 & ~x32 & ~x51 & ~x81 & ~x86 & ~x87 & ~x109 & ~x138 & ~x139 & ~x141 & ~x142 & ~x145 & ~x164 & ~x167 & ~x172 & ~x193 & ~x197 & ~x198 & ~x199 & ~x223 & ~x224 & ~x227 & ~x247 & ~x249 & ~x250 & ~x251 & ~x254 & ~x255 & ~x275 & ~x277 & ~x279 & ~x281 & ~x282 & ~x303 & ~x304 & ~x305 & ~x307 & ~x308 & ~x332 & ~x333 & ~x336 & ~x337 & ~x361 & ~x362 & ~x364 & ~x390 & ~x393 & ~x417 & ~x420 & ~x421 & ~x473 & ~x488 & ~x499 & ~x501 & ~x503 & ~x507 & ~x509 & ~x529 & ~x531 & ~x532 & ~x559 & ~x561 & ~x564 & ~x586 & ~x587 & ~x589 & ~x590 & ~x592 & ~x613 & ~x614 & ~x616 & ~x620 & ~x642 & ~x643 & ~x644 & ~x645 & ~x647 & ~x671 & ~x672 & ~x677 & ~x678 & ~x695 & ~x696 & ~x698 & ~x701 & ~x704 & ~x725 & ~x726 & ~x727 & ~x728 & ~x732 & ~x751 & ~x752 & ~x753 & ~x754 & ~x757 & ~x758 & ~x759 & ~x762 & ~x764 & ~x777 & ~x779 & ~x781 & ~x782;
assign c3294 =  x275;
assign c3296 =  x37 &  x47 &  x93 &  x94 &  x95 &  x124 &  x739 &  x742 & ~x58 & ~x87 & ~x113 & ~x139 & ~x249 & ~x256 & ~x310 & ~x388;
assign c3298 =  x742 & ~x3 & ~x4 & ~x6 & ~x19 & ~x26 & ~x29 & ~x32 & ~x53 & ~x59 & ~x80 & ~x81 & ~x110 & ~x111 & ~x112 & ~x139 & ~x144 & ~x170 & ~x171 & ~x194 & ~x196 & ~x198 & ~x199 & ~x200 & ~x220 & ~x222 & ~x223 & ~x229 & ~x243 & ~x244 & ~x252 & ~x255 & ~x260 & ~x272 & ~x276 & ~x302 & ~x305 & ~x307 & ~x309 & ~x314 & ~x330 & ~x331 & ~x334 & ~x336 & ~x340 & ~x343 & ~x363 & ~x370 & ~x371 & ~x388 & ~x390 & ~x395 & ~x398 & ~x399 & ~x418 & ~x425 & ~x426 & ~x441 & ~x444 & ~x447 & ~x450 & ~x455 & ~x469 & ~x472 & ~x478 & ~x479 & ~x480 & ~x482 & ~x500 & ~x510 & ~x527 & ~x531 & ~x532 & ~x534 & ~x555 & ~x558 & ~x564 & ~x587 & ~x612 & ~x613 & ~x614 & ~x615 & ~x620 & ~x638 & ~x643 & ~x649 & ~x673 & ~x696 & ~x697 & ~x729 & ~x731 & ~x732 & ~x760 & ~x761 & ~x779 & ~x781 & ~x782;
assign c3300 = ~x4 & ~x5 & ~x20 & ~x27 & ~x87 & ~x107 & ~x110 & ~x112 & ~x115 & ~x117 & ~x136 & ~x166 & ~x195 & ~x199 & ~x200 & ~x224 & ~x225 & ~x228 & ~x229 & ~x230 & ~x243 & ~x244 & ~x250 & ~x252 & ~x253 & ~x254 & ~x259 & ~x272 & ~x273 & ~x281 & ~x283 & ~x303 & ~x309 & ~x338 & ~x340 & ~x343 & ~x357 & ~x360 & ~x371 & ~x385 & ~x390 & ~x392 & ~x396 & ~x414 & ~x420 & ~x422 & ~x442 & ~x453 & ~x454 & ~x499 & ~x507 & ~x528 & ~x536 & ~x537 & ~x557 & ~x559 & ~x564 & ~x565 & ~x587 & ~x592 & ~x616 & ~x668 & ~x669 & ~x670 & ~x695 & ~x696 & ~x701 & ~x703 & ~x727 & ~x751 & ~x757 & ~x759 & ~x761 & ~x767 & ~x782;
assign c3302 =  x315 &  x548 & ~x52 & ~x55 & ~x58 & ~x62 & ~x108 & ~x109 & ~x110 & ~x117 & ~x118 & ~x162 & ~x198 & ~x202 & ~x220 & ~x226 & ~x257 & ~x310 & ~x366 & ~x418 & ~x446 & ~x449 & ~x504 & ~x563 & ~x581 & ~x609 & ~x610 & ~x617 & ~x618 & ~x669 & ~x705 & ~x723 & ~x727 & ~x752 & ~x756 & ~x758 & ~x782;
assign c3304 = ~x170 & ~x182 & ~x275 & ~x329 & ~x372 & ~x592 & ~x593 & ~x765;
assign c3306 = ~x6 & ~x24 & ~x30 & ~x33 & ~x50 & ~x55 & ~x56 & ~x88 & ~x107 & ~x114 & ~x125 & ~x167 & ~x192 & ~x196 & ~x220 & ~x226 & ~x228 & ~x250 & ~x307 & ~x334 & ~x335 & ~x337 & ~x338 & ~x360 & ~x396 & ~x398 & ~x417 & ~x420 & ~x423 & ~x449 & ~x474 & ~x475 & ~x503 & ~x505 & ~x528 & ~x533 & ~x534 & ~x561 & ~x562 & ~x584 & ~x589 & ~x620 & ~x622 & ~x643 & ~x649 & ~x651 & ~x666 & ~x695 & ~x700 & ~x704 & ~x732 & ~x750 & ~x751 & ~x753 & ~x754 & ~x759 & ~x762 & ~x777 & ~x780;
assign c3308 =  x65 &  x103 &  x128 &  x209 &  x244 &  x272 &  x379 &  x486 &  x604 &  x654 &  x655 &  x685 & ~x28 & ~x82 & ~x117 & ~x172 & ~x256 & ~x303 & ~x341 & ~x364 & ~x418 & ~x559 & ~x642 & ~x672 & ~x675 & ~x727 & ~x777;
assign c3310 =  x541 &  x651 &  x749 & ~x8 & ~x9 & ~x166 & ~x171 & ~x303 & ~x360 & ~x365 & ~x474 & ~x586;
assign c3312 =  x37 & ~x19 & ~x21 & ~x22 & ~x29 & ~x52 & ~x56 & ~x58 & ~x79 & ~x85 & ~x107 & ~x112 & ~x115 & ~x140 & ~x165 & ~x167 & ~x194 & ~x220 & ~x221 & ~x247 & ~x249 & ~x253 & ~x257 & ~x277 & ~x279 & ~x282 & ~x283 & ~x304 & ~x308 & ~x336 & ~x340 & ~x361 & ~x362 & ~x364 & ~x389 & ~x390 & ~x418 & ~x421 & ~x447 & ~x449 & ~x452 & ~x477 & ~x479 & ~x500 & ~x558 & ~x560 & ~x564 & ~x643 & ~x699 & ~x756 & ~x757 & ~x760 & ~x761 & ~x780;
assign c3314 =  x376 &  x682 &  x710 & ~x18 & ~x20 & ~x60 & ~x83 & ~x252 & ~x308 & ~x411 & ~x506 & ~x648 & ~x667 & ~x727;
assign c3316 =  x414 & ~x27 & ~x81 & ~x87 & ~x89 & ~x109 & ~x114 & ~x144 & ~x163 & ~x192 & ~x196 & ~x253 & ~x280 & ~x333 & ~x365 & ~x532 & ~x584 & ~x585 & ~x590 & ~x612 & ~x618 & ~x619 & ~x620 & ~x638 & ~x639 & ~x641 & ~x667 & ~x673 & ~x675 & ~x696 & ~x697 & ~x701 & ~x726 & ~x728 & ~x754 & ~x758 & ~x761 & ~x778;
assign c3318 =  x158 &  x216 &  x405 & ~x5 & ~x33 & ~x87 & ~x89 & ~x106 & ~x109 & ~x114 & ~x143 & ~x197 & ~x221 & ~x222 & ~x228 & ~x248 & ~x255 & ~x277 & ~x279 & ~x305 & ~x310 & ~x419 & ~x420 & ~x503 & ~x530 & ~x556 & ~x590 & ~x592 & ~x595 & ~x613 & ~x615 & ~x643 & ~x668 & ~x676 & ~x696 & ~x729 & ~x733 & ~x751 & ~x755 & ~x759;
assign c3320 = ~x404;
assign c3322 =  x311;
assign c3324 = ~x7 & ~x14 & ~x41 & ~x43 & ~x63 & ~x85 & ~x227 & ~x306 & ~x390 & ~x701 & ~x749 & ~x750 & ~x753 & ~x760 & ~x761 & ~x779;
assign c3326 =  x93 &  x102 &  x152 &  x209 &  x295 &  x297 &  x348 &  x437 &  x461 &  x520 &  x553 &  x579 &  x598 &  x603 &  x653 &  x654 &  x737 & ~x4 & ~x22 & ~x29 & ~x30 & ~x49 & ~x53 & ~x79 & ~x81 & ~x108 & ~x109 & ~x141 & ~x200 & ~x276 & ~x283 & ~x332 & ~x339 & ~x419 & ~x475 & ~x534 & ~x759;
assign c3328 =  x539 & ~x0 & ~x107 & ~x110 & ~x223 & ~x248 & ~x253 & ~x278 & ~x315 & ~x559 & ~x615 & ~x702;
assign c3330 =  x47 & ~x288 & ~x471 & ~x483 & ~x504 & ~x558 & ~x728 & ~x780;
assign c3332 =  x69 &  x70 &  x208 &  x377 &  x405 &  x461 &  x490 &  x546 &  x547 &  x714 &  x739 & ~x86 & ~x88 & ~x141 & ~x162 & ~x166 & ~x219 & ~x221 & ~x307 & ~x313 & ~x385 & ~x416 & ~x443 & ~x472 & ~x480 & ~x499 & ~x505 & ~x557 & ~x561 & ~x611 & ~x636 & ~x639 & ~x693 & ~x726 & ~x727 & ~x752 & ~x780;
assign c3334 = ~x1 & ~x23 & ~x28 & ~x33 & ~x55 & ~x82 & ~x84 & ~x114 & ~x134 & ~x165 & ~x197 & ~x199 & ~x229 & ~x247 & ~x249 & ~x254 & ~x259 & ~x301 & ~x305 & ~x333 & ~x364 & ~x369 & ~x398 & ~x417 & ~x421 & ~x422 & ~x445 & ~x450 & ~x451 & ~x452 & ~x472 & ~x477 & ~x481 & ~x502 & ~x508 & ~x520 & ~x529 & ~x530 & ~x563 & ~x564 & ~x612 & ~x614 & ~x732 & ~x780;
assign c3336 = ~x2 & ~x27 & ~x61 & ~x81 & ~x88 & ~x106 & ~x107 & ~x109 & ~x111 & ~x112 & ~x114 & ~x134 & ~x141 & ~x162 & ~x166 & ~x172 & ~x193 & ~x198 & ~x200 & ~x219 & ~x226 & ~x248 & ~x250 & ~x255 & ~x256 & ~x278 & ~x279 & ~x304 & ~x307 & ~x335 & ~x344 & ~x355 & ~x361 & ~x364 & ~x419 & ~x420 & ~x423 & ~x474 & ~x475 & ~x476 & ~x477 & ~x506 & ~x507 & ~x536 & ~x537 & ~x539 & ~x556 & ~x560 & ~x563 & ~x565 & ~x581 & ~x583 & ~x584 & ~x587 & ~x590 & ~x591 & ~x610 & ~x611 & ~x619 & ~x642 & ~x643 & ~x646 & ~x649 & ~x667 & ~x668 & ~x671 & ~x672 & ~x676 & ~x696 & ~x723 & ~x725 & ~x727 & ~x752 & ~x760 & ~x761 & ~x768 & ~x777;
assign c3338 = ~x55 & ~x144 & ~x249 & ~x310 & ~x325 & ~x334 & ~x390 & ~x473 & ~x522 & ~x556 & ~x642 & ~x676 & ~x703 & ~x747;
assign c3340 =  x397 & ~x30 & ~x56 & ~x84 & ~x109 & ~x136 & ~x167 & ~x171 & ~x193 & ~x195 & ~x281 & ~x334 & ~x336 & ~x392 & ~x533 & ~x559 & ~x590 & ~x670 & ~x676 & ~x701 & ~x723 & ~x726 & ~x757;
assign c3342 =  x95 &  x152 &  x263 &  x598 &  x602 &  x626 & ~x2 & ~x80 & ~x86 & ~x119 & ~x143 & ~x165 & ~x194 & ~x222 & ~x248 & ~x251 & ~x257 & ~x276 & ~x279 & ~x305 & ~x311 & ~x314 & ~x340 & ~x359 & ~x360 & ~x398 & ~x416 & ~x426 & ~x451 & ~x536 & ~x595 & ~x611 & ~x729 & ~x758 & ~x777;
assign c3344 =  x287 &  x385 &  x743 & ~x169 & ~x171 & ~x193 & ~x225 & ~x229 & ~x360 & ~x390 & ~x452 & ~x589 & ~x620 & ~x669 & ~x673 & ~x677 & ~x699 & ~x755 & ~x758 & ~x780;
assign c3346 =  x149 & ~x14 & ~x170 & ~x389 & ~x422 & ~x514 & ~x533 & ~x558 & ~x619 & ~x703 & ~x754;
assign c3348 =  x38 &  x120 &  x350 &  x738 & ~x2 & ~x31 & ~x34 & ~x48 & ~x61 & ~x84 & ~x106 & ~x117 & ~x166 & ~x194 & ~x221 & ~x278 & ~x308 & ~x473 & ~x531 & ~x558 & ~x590 & ~x617 & ~x637 & ~x670 & ~x676 & ~x705 & ~x729;
assign c3350 =  x269 &  x379 &  x438 & ~x2 & ~x24 & ~x25 & ~x26 & ~x28 & ~x31 & ~x50 & ~x54 & ~x55 & ~x58 & ~x60 & ~x79 & ~x80 & ~x81 & ~x82 & ~x83 & ~x107 & ~x112 & ~x136 & ~x138 & ~x139 & ~x140 & ~x141 & ~x144 & ~x163 & ~x170 & ~x192 & ~x193 & ~x196 & ~x197 & ~x199 & ~x221 & ~x222 & ~x224 & ~x247 & ~x249 & ~x251 & ~x253 & ~x254 & ~x276 & ~x278 & ~x279 & ~x280 & ~x281 & ~x303 & ~x304 & ~x305 & ~x310 & ~x311 & ~x312 & ~x327 & ~x333 & ~x336 & ~x338 & ~x362 & ~x363 & ~x364 & ~x367 & ~x390 & ~x392 & ~x417 & ~x418 & ~x420 & ~x422 & ~x444 & ~x447 & ~x451 & ~x476 & ~x504 & ~x505 & ~x506 & ~x532 & ~x556 & ~x561 & ~x562 & ~x587 & ~x590 & ~x615 & ~x618 & ~x641 & ~x642 & ~x645 & ~x669 & ~x671 & ~x673 & ~x701 & ~x702 & ~x703 & ~x723 & ~x729 & ~x757 & ~x758 & ~x762 & ~x781 & ~x783;
assign c3352 =  x132 &  x148 &  x397 &  x440 & ~x112 & ~x279 & ~x363 & ~x616 & ~x648 & ~x675 & ~x676;
assign c3354 =  x179 &  x346 &  x485 & ~x144 & ~x196 & ~x204 & ~x226 & ~x308 & ~x583 & ~x590 & ~x672 & ~x725;
assign c3356 =  x394;
assign c3358 =  x271 &  x288 &  x686 & ~x58 & ~x61 & ~x77 & ~x106 & ~x134 & ~x161 & ~x162 & ~x172 & ~x197 & ~x220 & ~x283 & ~x447 & ~x479 & ~x504 & ~x529 & ~x558 & ~x580 & ~x589 & ~x618 & ~x667 & ~x723 & ~x750;
assign c3360 =  x471 & ~x19 & ~x54 & ~x224;
assign c3362 =  x37 &  x46 &  x47 &  x297 &  x497 & ~x23 & ~x25 & ~x86 & ~x113 & ~x224 & ~x360 & ~x391 & ~x393 & ~x449 & ~x643 & ~x729 & ~x754;
assign c3364 =  x66 &  x67 &  x95 &  x128 &  x401 &  x406 &  x434 &  x461 &  x517 &  x600 & ~x1 & ~x19 & ~x27 & ~x32 & ~x47 & ~x50 & ~x52 & ~x58 & ~x62 & ~x63 & ~x81 & ~x89 & ~x105 & ~x111 & ~x115 & ~x134 & ~x145 & ~x164 & ~x165 & ~x195 & ~x201 & ~x229 & ~x248 & ~x249 & ~x283 & ~x284 & ~x306 & ~x358 & ~x368 & ~x419 & ~x424 & ~x425 & ~x445 & ~x446 & ~x447 & ~x472 & ~x480 & ~x501 & ~x503 & ~x508 & ~x535 & ~x559 & ~x560 & ~x565 & ~x585 & ~x612 & ~x613 & ~x621 & ~x640 & ~x648 & ~x649 & ~x667 & ~x696 & ~x778 & ~x781;
assign c3366 =  x123 &  x124 &  x290 &  x485 &  x653 &  x708 & ~x1 & ~x25 & ~x27 & ~x30 & ~x55 & ~x80 & ~x83 & ~x86 & ~x109 & ~x112 & ~x114 & ~x138 & ~x139 & ~x168 & ~x196 & ~x199 & ~x231 & ~x245 & ~x253 & ~x254 & ~x258 & ~x259 & ~x273 & ~x279 & ~x285 & ~x305 & ~x311 & ~x331 & ~x336 & ~x338 & ~x362 & ~x387 & ~x388 & ~x389 & ~x390 & ~x397 & ~x419 & ~x452 & ~x470 & ~x481 & ~x502 & ~x503 & ~x527 & ~x532 & ~x560 & ~x562 & ~x615 & ~x616 & ~x646 & ~x699 & ~x730 & ~x756 & ~x760 & ~x780 & ~x783;
assign c3368 = ~x5 & ~x9 & ~x31 & ~x62 & ~x78 & ~x84 & ~x115 & ~x116 & ~x136 & ~x138 & ~x144 & ~x145 & ~x168 & ~x197 & ~x219 & ~x252 & ~x257 & ~x281 & ~x285 & ~x308 & ~x392 & ~x450 & ~x477 & ~x509 & ~x531 & ~x592 & ~x615 & ~x619 & ~x683 & ~x695 & ~x704 & ~x721 & ~x729 & ~x749 & ~x750 & ~x755 & ~x781;
assign c3370 = ~x2 & ~x5 & ~x19 & ~x23 & ~x24 & ~x55 & ~x56 & ~x58 & ~x81 & ~x83 & ~x84 & ~x85 & ~x108 & ~x109 & ~x110 & ~x114 & ~x116 & ~x136 & ~x168 & ~x170 & ~x174 & ~x222 & ~x226 & ~x227 & ~x228 & ~x252 & ~x254 & ~x279 & ~x280 & ~x284 & ~x285 & ~x303 & ~x305 & ~x340 & ~x364 & ~x368 & ~x416 & ~x417 & ~x419 & ~x463 & ~x472 & ~x473 & ~x475 & ~x481 & ~x503 & ~x505 & ~x530 & ~x536 & ~x559 & ~x587 & ~x589 & ~x613 & ~x643 & ~x646 & ~x727 & ~x728 & ~x729 & ~x754 & ~x757 & ~x758 & ~x759 & ~x762 & ~x774 & ~x776 & ~x777 & ~x780 & ~x783;
assign c3372 =  x105 &  x133 &  x358 &  x579 & ~x3 & ~x57 & ~x250 & ~x559 & ~x672;
assign c3374 =  x431 &  x436 &  x465 &  x517 &  x598 &  x682 &  x742 & ~x0 & ~x2 & ~x5 & ~x6 & ~x20 & ~x21 & ~x22 & ~x23 & ~x24 & ~x25 & ~x30 & ~x31 & ~x32 & ~x34 & ~x35 & ~x50 & ~x53 & ~x54 & ~x56 & ~x58 & ~x62 & ~x78 & ~x80 & ~x81 & ~x83 & ~x85 & ~x87 & ~x89 & ~x107 & ~x108 & ~x111 & ~x112 & ~x115 & ~x116 & ~x134 & ~x135 & ~x138 & ~x139 & ~x140 & ~x144 & ~x163 & ~x164 & ~x165 & ~x166 & ~x168 & ~x170 & ~x171 & ~x173 & ~x174 & ~x191 & ~x192 & ~x195 & ~x197 & ~x199 & ~x201 & ~x219 & ~x221 & ~x222 & ~x226 & ~x227 & ~x228 & ~x248 & ~x251 & ~x253 & ~x254 & ~x274 & ~x278 & ~x280 & ~x281 & ~x285 & ~x303 & ~x304 & ~x307 & ~x312 & ~x332 & ~x333 & ~x334 & ~x338 & ~x339 & ~x340 & ~x359 & ~x360 & ~x362 & ~x389 & ~x390 & ~x391 & ~x392 & ~x394 & ~x417 & ~x419 & ~x421 & ~x422 & ~x426 & ~x443 & ~x444 & ~x450 & ~x451 & ~x452 & ~x453 & ~x472 & ~x473 & ~x474 & ~x475 & ~x476 & ~x480 & ~x481 & ~x499 & ~x501 & ~x502 & ~x503 & ~x504 & ~x506 & ~x509 & ~x527 & ~x530 & ~x531 & ~x532 & ~x533 & ~x534 & ~x536 & ~x553 & ~x556 & ~x558 & ~x560 & ~x561 & ~x562 & ~x582 & ~x583 & ~x584 & ~x585 & ~x586 & ~x587 & ~x588 & ~x590 & ~x591 & ~x594 & ~x610 & ~x612 & ~x613 & ~x615 & ~x622 & ~x638 & ~x640 & ~x642 & ~x645 & ~x650 & ~x651 & ~x667 & ~x672 & ~x694 & ~x697 & ~x700 & ~x701 & ~x704 & ~x722 & ~x726 & ~x729 & ~x730 & ~x731 & ~x732 & ~x750 & ~x754 & ~x755 & ~x758 & ~x761 & ~x762 & ~x781 & ~x783;
assign c3376 =  x120 &  x629 &  x714 &  x716 &  x738 & ~x6 & ~x19 & ~x20 & ~x23 & ~x24 & ~x27 & ~x30 & ~x59 & ~x60 & ~x90 & ~x107 & ~x117 & ~x136 & ~x253 & ~x257 & ~x278 & ~x330 & ~x335 & ~x341 & ~x387 & ~x390 & ~x391 & ~x451 & ~x453 & ~x478 & ~x479 & ~x502 & ~x530 & ~x532 & ~x535 & ~x587 & ~x650 & ~x651 & ~x678 & ~x699 & ~x700 & ~x702 & ~x754 & ~x763 & ~x781 & ~x782 & ~x783;
assign c3378 =  x37 &  x132 &  x658 & ~x1 & ~x3 & ~x4 & ~x26 & ~x29 & ~x52 & ~x56 & ~x84 & ~x87 & ~x88 & ~x115 & ~x137 & ~x142 & ~x144 & ~x166 & ~x170 & ~x191 & ~x220 & ~x225 & ~x308 & ~x333 & ~x335 & ~x366 & ~x447 & ~x530 & ~x534 & ~x621 & ~x623 & ~x646 & ~x674 & ~x676 & ~x704 & ~x733 & ~x783;
assign c3380 = ~x7 & ~x9 & ~x28 & ~x58 & ~x77 & ~x85 & ~x86 & ~x87 & ~x134 & ~x145 & ~x163 & ~x164 & ~x169 & ~x170 & ~x171 & ~x172 & ~x199 & ~x226 & ~x249 & ~x278 & ~x303 & ~x331 & ~x336 & ~x453 & ~x475 & ~x529 & ~x571 & ~x610 & ~x612 & ~x618 & ~x620 & ~x667 & ~x670 & ~x672 & ~x725 & ~x727 & ~x761 & ~x779 & ~x780 & ~x781;
assign c3382 =  x120 &  x124 &  x125 &  x128 &  x132 &  x160 &  x623 & ~x59 & ~x143 & ~x225 & ~x583 & ~x778;
assign c3384 =  x213 &  x236 &  x265 &  x293 &  x348 &  x467 &  x605 &  x625 &  x629 & ~x30 & ~x57 & ~x81 & ~x253 & ~x272 & ~x282 & ~x365 & ~x501 & ~x530 & ~x559 & ~x618 & ~x730 & ~x754 & ~x759;
assign c3386 =  x97 &  x123 &  x294 &  x318 & ~x27 & ~x53 & ~x140 & ~x232 & ~x259 & ~x281 & ~x336 & ~x505 & ~x530 & ~x561 & ~x728 & ~x755;
assign c3388 = ~x143 & ~x206 & ~x234 & ~x305 & ~x329 & ~x552;
assign c3390 = ~x31 & ~x145 & ~x171 & ~x220 & ~x261 & ~x344 & ~x389 & ~x394 & ~x451 & ~x472 & ~x529 & ~x586 & ~x726 & ~x733 & ~x757 & ~x762 & ~x768 & ~x777;
assign c3392 = ~x8 & ~x19 & ~x53 & ~x54 & ~x58 & ~x61 & ~x106 & ~x138 & ~x139 & ~x145 & ~x168 & ~x196 & ~x201 & ~x223 & ~x248 & ~x281 & ~x306 & ~x331 & ~x333 & ~x360 & ~x365 & ~x379 & ~x418 & ~x471 & ~x474 & ~x550 & ~x561 & ~x589 & ~x590 & ~x614 & ~x648 & ~x672 & ~x728 & ~x733 & ~x752 & ~x759 & ~x761;
assign c3394 = ~x14 & ~x23 & ~x80 & ~x85 & ~x117 & ~x134 & ~x139 & ~x141 & ~x165 & ~x166 & ~x170 & ~x173 & ~x199 & ~x225 & ~x260 & ~x261 & ~x316 & ~x339 & ~x356 & ~x361 & ~x372 & ~x423 & ~x445 & ~x450 & ~x472 & ~x529 & ~x534 & ~x557 & ~x586 & ~x621 & ~x638 & ~x643 & ~x672 & ~x677 & ~x695 & ~x696 & ~x704 & ~x726 & ~x729 & ~x731 & ~x751 & ~x764;
assign c3396 =  x450;
assign c3398 = ~x222 & ~x289 & ~x528 & ~x572;
assign c3400 =  x149 &  x232 &  x319 &  x329 & ~x2 & ~x5 & ~x6 & ~x19 & ~x21 & ~x32 & ~x48 & ~x139 & ~x162 & ~x172 & ~x197 & ~x200 & ~x219 & ~x249 & ~x250 & ~x278 & ~x281 & ~x310 & ~x335 & ~x337 & ~x476 & ~x503 & ~x531 & ~x586 & ~x591 & ~x594 & ~x644 & ~x649 & ~x666 & ~x667 & ~x668 & ~x675 & ~x698 & ~x699 & ~x700 & ~x704 & ~x726 & ~x728 & ~x755;
assign c3402 =  x311;
assign c3404 =  x37 &  x42 &  x205 &  x736 &  x746 & ~x195 & ~x226 & ~x248 & ~x307 & ~x332 & ~x334 & ~x338 & ~x360 & ~x447 & ~x474 & ~x502 & ~x643 & ~x701 & ~x781;
assign c3406 =  x69 &  x70 &  x126 &  x179 &  x182 &  x235 &  x318 &  x629 &  x735 & ~x9 & ~x114 & ~x115 & ~x227 & ~x419 & ~x503 & ~x558 & ~x617;
assign c3408 =  x17 &  x457 &  x485 &  x735 &  x737 & ~x111 & ~x165 & ~x171 & ~x195 & ~x197 & ~x199 & ~x221 & ~x255 & ~x306 & ~x332 & ~x335 & ~x340 & ~x534 & ~x562;
assign c3410 =  x70 &  x125 &  x127 &  x157 &  x209 &  x237 &  x293 &  x375 &  x434 &  x516 &  x547 &  x574 &  x605 &  x633 &  x658 &  x660 &  x714 &  x716 &  x741 &  x743 & ~x3 & ~x7 & ~x35 & ~x54 & ~x60 & ~x63 & ~x82 & ~x106 & ~x108 & ~x112 & ~x117 & ~x138 & ~x144 & ~x171 & ~x228 & ~x229 & ~x250 & ~x251 & ~x280 & ~x305 & ~x338 & ~x339 & ~x341 & ~x360 & ~x390 & ~x425 & ~x475 & ~x478 & ~x482 & ~x504 & ~x506 & ~x508 & ~x555 & ~x581 & ~x587 & ~x594 & ~x612 & ~x642 & ~x644 & ~x650 & ~x674 & ~x726 & ~x762 & ~x778;
assign c3412 =  x745 & ~x1 & ~x2 & ~x3 & ~x5 & ~x7 & ~x12 & ~x24 & ~x27 & ~x28 & ~x31 & ~x32 & ~x34 & ~x49 & ~x50 & ~x56 & ~x57 & ~x58 & ~x60 & ~x61 & ~x78 & ~x85 & ~x86 & ~x89 & ~x108 & ~x110 & ~x111 & ~x114 & ~x117 & ~x136 & ~x139 & ~x141 & ~x142 & ~x164 & ~x165 & ~x169 & ~x170 & ~x194 & ~x196 & ~x197 & ~x200 & ~x222 & ~x223 & ~x224 & ~x227 & ~x228 & ~x229 & ~x247 & ~x248 & ~x249 & ~x253 & ~x254 & ~x255 & ~x256 & ~x276 & ~x278 & ~x279 & ~x282 & ~x284 & ~x304 & ~x306 & ~x307 & ~x309 & ~x310 & ~x311 & ~x312 & ~x331 & ~x334 & ~x336 & ~x337 & ~x339 & ~x359 & ~x360 & ~x362 & ~x363 & ~x366 & ~x368 & ~x387 & ~x388 & ~x389 & ~x391 & ~x395 & ~x416 & ~x419 & ~x424 & ~x443 & ~x447 & ~x449 & ~x450 & ~x451 & ~x471 & ~x472 & ~x474 & ~x476 & ~x480 & ~x481 & ~x501 & ~x502 & ~x505 & ~x506 & ~x507 & ~x532 & ~x534 & ~x535 & ~x557 & ~x558 & ~x562 & ~x584 & ~x586 & ~x588 & ~x589 & ~x590 & ~x591 & ~x612 & ~x613 & ~x614 & ~x618 & ~x644 & ~x646 & ~x647 & ~x651 & ~x666 & ~x673 & ~x674 & ~x679 & ~x693 & ~x694 & ~x696 & ~x698 & ~x699 & ~x700 & ~x701 & ~x702 & ~x703 & ~x704 & ~x705 & ~x707 & ~x722 & ~x724 & ~x729 & ~x730 & ~x731 & ~x733 & ~x734 & ~x750 & ~x755 & ~x758 & ~x762 & ~x778 & ~x779 & ~x780;
assign c3414 =  x711 & ~x2 & ~x8 & ~x17 & ~x21 & ~x22 & ~x23 & ~x28 & ~x35 & ~x50 & ~x51 & ~x56 & ~x59 & ~x61 & ~x62 & ~x78 & ~x80 & ~x86 & ~x87 & ~x90 & ~x110 & ~x111 & ~x112 & ~x135 & ~x144 & ~x163 & ~x165 & ~x192 & ~x195 & ~x200 & ~x201 & ~x202 & ~x219 & ~x222 & ~x225 & ~x249 & ~x250 & ~x251 & ~x253 & ~x256 & ~x257 & ~x278 & ~x280 & ~x303 & ~x304 & ~x309 & ~x331 & ~x333 & ~x335 & ~x340 & ~x360 & ~x361 & ~x363 & ~x364 & ~x392 & ~x394 & ~x395 & ~x397 & ~x401 & ~x416 & ~x420 & ~x422 & ~x445 & ~x446 & ~x447 & ~x449 & ~x451 & ~x452 & ~x472 & ~x474 & ~x478 & ~x500 & ~x501 & ~x507 & ~x508 & ~x528 & ~x530 & ~x537 & ~x559 & ~x563 & ~x586 & ~x591 & ~x592 & ~x593 & ~x613 & ~x621 & ~x638 & ~x639 & ~x641 & ~x642 & ~x646 & ~x649 & ~x675 & ~x676 & ~x678 & ~x679 & ~x694 & ~x702 & ~x704 & ~x705 & ~x728 & ~x729 & ~x731 & ~x734 & ~x752 & ~x753 & ~x763 & ~x778 & ~x783;
assign c3416 = ~x4 & ~x10 & ~x62 & ~x77 & ~x105 & ~x145 & ~x163 & ~x241 & ~x304 & ~x382 & ~x473 & ~x497 & ~x508 & ~x635 & ~x666 & ~x703 & ~x750;
assign c3418 =  x275;
assign c3420 =  x98 &  x99 &  x180 &  x208 &  x601 &  x630 &  x658 & ~x3 & ~x4 & ~x8 & ~x19 & ~x21 & ~x26 & ~x29 & ~x33 & ~x80 & ~x85 & ~x87 & ~x105 & ~x136 & ~x223 & ~x224 & ~x229 & ~x278 & ~x284 & ~x397 & ~x416 & ~x420 & ~x450 & ~x553 & ~x588 & ~x644 & ~x664 & ~x670 & ~x724 & ~x748 & ~x761;
assign c3422 =  x34 &  x46;
assign c3424 =  x124 &  x293 &  x403 &  x663 &  x714 &  x719 & ~x6 & ~x7 & ~x23 & ~x26 & ~x28 & ~x29 & ~x31 & ~x52 & ~x53 & ~x54 & ~x55 & ~x80 & ~x81 & ~x106 & ~x107 & ~x108 & ~x110 & ~x112 & ~x114 & ~x117 & ~x139 & ~x165 & ~x171 & ~x198 & ~x199 & ~x200 & ~x220 & ~x221 & ~x223 & ~x225 & ~x227 & ~x248 & ~x249 & ~x251 & ~x253 & ~x276 & ~x281 & ~x283 & ~x285 & ~x304 & ~x308 & ~x309 & ~x310 & ~x332 & ~x334 & ~x335 & ~x361 & ~x393 & ~x395 & ~x419 & ~x443 & ~x446 & ~x447 & ~x449 & ~x480 & ~x505 & ~x527 & ~x528 & ~x533 & ~x534 & ~x557 & ~x561 & ~x583 & ~x585 & ~x586 & ~x614 & ~x620 & ~x623 & ~x643 & ~x650 & ~x668 & ~x669 & ~x671 & ~x673 & ~x677 & ~x694 & ~x697 & ~x703 & ~x723 & ~x726 & ~x731 & ~x755 & ~x757 & ~x762 & ~x780;
assign c3426 = ~x2 & ~x8 & ~x9 & ~x25 & ~x30 & ~x33 & ~x56 & ~x58 & ~x84 & ~x88 & ~x89 & ~x111 & ~x113 & ~x166 & ~x167 & ~x168 & ~x193 & ~x198 & ~x199 & ~x223 & ~x226 & ~x231 & ~x251 & ~x252 & ~x253 & ~x254 & ~x257 & ~x276 & ~x280 & ~x281 & ~x303 & ~x305 & ~x306 & ~x308 & ~x312 & ~x333 & ~x336 & ~x338 & ~x341 & ~x362 & ~x364 & ~x367 & ~x369 & ~x388 & ~x392 & ~x395 & ~x396 & ~x397 & ~x416 & ~x418 & ~x419 & ~x421 & ~x422 & ~x425 & ~x447 & ~x450 & ~x472 & ~x473 & ~x474 & ~x480 & ~x481 & ~x500 & ~x532 & ~x534 & ~x558 & ~x561 & ~x613 & ~x619 & ~x644 & ~x646 & ~x655 & ~x697 & ~x751 & ~x754 & ~x755 & ~x758 & ~x760 & ~x761 & ~x783;
assign c3428 =  x291 &  x682 &  x710 &  x713 &  x741 & ~x3 & ~x7 & ~x22 & ~x23 & ~x26 & ~x27 & ~x29 & ~x30 & ~x32 & ~x35 & ~x54 & ~x55 & ~x79 & ~x80 & ~x84 & ~x86 & ~x88 & ~x90 & ~x105 & ~x106 & ~x109 & ~x111 & ~x114 & ~x134 & ~x135 & ~x136 & ~x137 & ~x138 & ~x139 & ~x143 & ~x145 & ~x162 & ~x164 & ~x169 & ~x170 & ~x172 & ~x190 & ~x195 & ~x199 & ~x219 & ~x225 & ~x226 & ~x228 & ~x248 & ~x252 & ~x256 & ~x275 & ~x276 & ~x279 & ~x281 & ~x282 & ~x305 & ~x309 & ~x312 & ~x333 & ~x334 & ~x336 & ~x337 & ~x338 & ~x363 & ~x365 & ~x366 & ~x369 & ~x388 & ~x390 & ~x393 & ~x416 & ~x417 & ~x418 & ~x424 & ~x425 & ~x443 & ~x447 & ~x449 & ~x450 & ~x451 & ~x452 & ~x470 & ~x473 & ~x476 & ~x477 & ~x478 & ~x501 & ~x502 & ~x503 & ~x506 & ~x531 & ~x535 & ~x561 & ~x585 & ~x587 & ~x590 & ~x591 & ~x608 & ~x619 & ~x636 & ~x640 & ~x645 & ~x647 & ~x648 & ~x665 & ~x667 & ~x675 & ~x692 & ~x693 & ~x695 & ~x698 & ~x699 & ~x702 & ~x720 & ~x724 & ~x731 & ~x752 & ~x753 & ~x758 & ~x761 & ~x762 & ~x775 & ~x776 & ~x779 & ~x781 & ~x783;
assign c3430 =  x34;
assign c3432 =  x441 &  x624 & ~x35 & ~x113 & ~x194 & ~x257 & ~x331 & ~x337 & ~x674 & ~x705 & ~x727 & ~x754 & ~x763;
assign c3434 =  x678 & ~x231 & ~x259;
assign c3436 =  x123 &  x127 &  x150 &  x211 &  x350 &  x437 &  x463 &  x490 &  x515 &  x517 &  x521 &  x602 & ~x2 & ~x5 & ~x9 & ~x20 & ~x48 & ~x49 & ~x51 & ~x54 & ~x61 & ~x77 & ~x79 & ~x85 & ~x90 & ~x105 & ~x106 & ~x108 & ~x118 & ~x134 & ~x137 & ~x140 & ~x163 & ~x166 & ~x172 & ~x194 & ~x246 & ~x248 & ~x274 & ~x275 & ~x278 & ~x279 & ~x284 & ~x285 & ~x303 & ~x304 & ~x306 & ~x334 & ~x336 & ~x339 & ~x341 & ~x362 & ~x368 & ~x369 & ~x393 & ~x394 & ~x396 & ~x415 & ~x449 & ~x450 & ~x451 & ~x472 & ~x476 & ~x477 & ~x502 & ~x506 & ~x509 & ~x510 & ~x531 & ~x532 & ~x533 & ~x534 & ~x535 & ~x557 & ~x591 & ~x593 & ~x608 & ~x611 & ~x643 & ~x666 & ~x674 & ~x676 & ~x695 & ~x696 & ~x698 & ~x722 & ~x723 & ~x726 & ~x730 & ~x756 & ~x761 & ~x781;
assign c3438 =  x746 & ~x14 & ~x15 & ~x19 & ~x20 & ~x21 & ~x68 & ~x78 & ~x165 & ~x168 & ~x256 & ~x275 & ~x305 & ~x331 & ~x419 & ~x586 & ~x670 & ~x671 & ~x699 & ~x756 & ~x762;
assign c3440 =  x346 &  x513 & ~x24 & ~x289 & ~x363;
assign c3442 = ~x164 & ~x258 & ~x300 & ~x310 & ~x314 & ~x357 & ~x446 & ~x471 & ~x504 & ~x576 & ~x619 & ~x701 & ~x732;
assign c3444 = ~x2 & ~x4 & ~x18 & ~x19 & ~x20 & ~x27 & ~x52 & ~x81 & ~x84 & ~x108 & ~x112 & ~x116 & ~x135 & ~x143 & ~x172 & ~x194 & ~x198 & ~x200 & ~x220 & ~x223 & ~x278 & ~x279 & ~x280 & ~x306 & ~x331 & ~x332 & ~x338 & ~x360 & ~x387 & ~x389 & ~x416 & ~x445 & ~x479 & ~x492 & ~x502 & ~x586 & ~x587 & ~x588 & ~x589 & ~x613 & ~x615 & ~x616 & ~x620 & ~x640 & ~x642 & ~x695 & ~x696 & ~x697 & ~x699 & ~x704 & ~x727 & ~x750 & ~x761 & ~x781;
assign c3446 = ~x10 & ~x25 & ~x29 & ~x31 & ~x32 & ~x48 & ~x49 & ~x56 & ~x58 & ~x78 & ~x82 & ~x89 & ~x90 & ~x105 & ~x109 & ~x134 & ~x136 & ~x142 & ~x143 & ~x145 & ~x172 & ~x199 & ~x202 & ~x203 & ~x219 & ~x222 & ~x226 & ~x230 & ~x251 & ~x255 & ~x257 & ~x280 & ~x286 & ~x303 & ~x307 & ~x331 & ~x334 & ~x336 & ~x340 & ~x353 & ~x361 & ~x362 & ~x387 & ~x395 & ~x397 & ~x419 & ~x445 & ~x448 & ~x453 & ~x472 & ~x477 & ~x498 & ~x509 & ~x560 & ~x613 & ~x615 & ~x620 & ~x635 & ~x643 & ~x649 & ~x669 & ~x676 & ~x692 & ~x694 & ~x702 & ~x727 & ~x749 & ~x750 & ~x757 & ~x775 & ~x776;
assign c3448 =  x100 &  x182 &  x244 &  x545 & ~x6 & ~x14 & ~x35 & ~x90 & ~x168 & ~x249 & ~x363 & ~x446 & ~x504 & ~x562 & ~x589 & ~x753 & ~x755;
assign c3450 =  x37 &  x45 &  x132 &  x246 &  x274 &  x319 & ~x55 & ~x88 & ~x108 & ~x110 & ~x591 & ~x619 & ~x670 & ~x671;
assign c3452 =  x119 &  x120 &  x130 &  x342 &  x483 & ~x53 & ~x89 & ~x140 & ~x170 & ~x308 & ~x668 & ~x675 & ~x701 & ~x703 & ~x730 & ~x779;
assign c3454 =  x577 &  x686 & ~x0 & ~x32 & ~x55 & ~x110 & ~x116 & ~x164 & ~x221 & ~x260 & ~x338 & ~x339 & ~x396 & ~x398 & ~x425 & ~x427 & ~x442 & ~x479 & ~x504 & ~x528 & ~x584 & ~x586 & ~x619 & ~x646 & ~x701 & ~x756 & ~x759;
assign c3456 = ~x25 & ~x55 & ~x80 & ~x84 & ~x146 & ~x167 & ~x171 & ~x245 & ~x258 & ~x259 & ~x273 & ~x363 & ~x381 & ~x398 & ~x415 & ~x443 & ~x472 & ~x481 & ~x550 & ~x558 & ~x584 & ~x616 & ~x751 & ~x755;
assign c3458 =  x538 &  x736 & ~x14 & ~x19 & ~x83 & ~x113 & ~x166 & ~x226 & ~x227 & ~x248 & ~x279 & ~x303 & ~x331 & ~x337 & ~x506 & ~x561 & ~x588 & ~x616;
assign c3460 =  x373 & ~x1 & ~x24 & ~x31 & ~x52 & ~x54 & ~x83 & ~x168 & ~x204 & ~x229 & ~x232 & ~x260 & ~x273 & ~x282 & ~x332 & ~x359 & ~x365 & ~x368 & ~x396 & ~x399 & ~x415 & ~x416 & ~x420 & ~x447 & ~x448 & ~x450 & ~x453 & ~x531 & ~x621 & ~x644 & ~x699 & ~x726 & ~x728 & ~x756 & ~x778;
assign c3462 =  x65 &  x70 &  x148 &  x237 &  x315 &  x519 &  x570 &  x658 &  x688 &  x738 &  x744 & ~x0 & ~x19 & ~x21 & ~x23 & ~x25 & ~x28 & ~x35 & ~x87 & ~x105 & ~x108 & ~x163 & ~x172 & ~x192 & ~x195 & ~x275 & ~x283 & ~x310 & ~x311 & ~x338 & ~x389 & ~x474 & ~x502 & ~x505 & ~x534 & ~x616 & ~x621 & ~x641 & ~x649 & ~x671 & ~x698 & ~x754;
assign c3464 = ~x8 & ~x23 & ~x72 & ~x112 & ~x113 & ~x378 & ~x415 & ~x473 & ~x530;
assign c3466 = ~x74 & ~x318 & ~x330 & ~x505 & ~x506 & ~x513 & ~x586 & ~x680 & ~x704 & ~x709;
assign c3468 =  x350 &  x574 & ~x1 & ~x2 & ~x3 & ~x10 & ~x23 & ~x30 & ~x58 & ~x80 & ~x85 & ~x110 & ~x139 & ~x142 & ~x166 & ~x221 & ~x222 & ~x224 & ~x229 & ~x276 & ~x282 & ~x288 & ~x307 & ~x312 & ~x315 & ~x328 & ~x340 & ~x358 & ~x360 & ~x365 & ~x371 & ~x386 & ~x389 & ~x399 & ~x413 & ~x414 & ~x416 & ~x419 & ~x421 & ~x422 & ~x427 & ~x444 & ~x450 & ~x452 & ~x453 & ~x454 & ~x470 & ~x471 & ~x472 & ~x473 & ~x475 & ~x480 & ~x482 & ~x500 & ~x506 & ~x508 & ~x528 & ~x529 & ~x555 & ~x562 & ~x583 & ~x592 & ~x668 & ~x674 & ~x697 & ~x698 & ~x700 & ~x702 & ~x724 & ~x732 & ~x752 & ~x754 & ~x758 & ~x779;
assign c3470 = ~x57 & ~x71 & ~x85 & ~x87 & ~x114 & ~x199 & ~x282 & ~x307 & ~x363 & ~x407 & ~x472 & ~x500 & ~x530 & ~x532 & ~x586 & ~x640 & ~x697 & ~x700 & ~x705 & ~x725 & ~x779;
assign c3472 =  x538 &  x553 &  x635 & ~x1 & ~x8 & ~x14 & ~x85 & ~x167 & ~x221 & ~x227 & ~x279 & ~x504 & ~x701;
assign c3474 =  x95 &  x104 &  x189 &  x551 &  x739 & ~x32 & ~x87 & ~x166 & ~x228 & ~x365 & ~x392 & ~x476 & ~x477 & ~x700;
assign c3476 = ~x25 & ~x27 & ~x61 & ~x163 & ~x164 & ~x231 & ~x246 & ~x249 & ~x258 & ~x275 & ~x276 & ~x330 & ~x359 & ~x369 & ~x391 & ~x419 & ~x425 & ~x478 & ~x548 & ~x755 & ~x760;
assign c3478 = ~x1 & ~x4 & ~x6 & ~x10 & ~x21 & ~x55 & ~x56 & ~x59 & ~x60 & ~x78 & ~x80 & ~x81 & ~x84 & ~x89 & ~x106 & ~x135 & ~x138 & ~x139 & ~x145 & ~x163 & ~x168 & ~x174 & ~x192 & ~x194 & ~x195 & ~x198 & ~x200 & ~x220 & ~x225 & ~x226 & ~x252 & ~x255 & ~x258 & ~x279 & ~x282 & ~x285 & ~x305 & ~x331 & ~x334 & ~x335 & ~x338 & ~x339 & ~x360 & ~x367 & ~x369 & ~x370 & ~x391 & ~x395 & ~x416 & ~x417 & ~x418 & ~x421 & ~x423 & ~x424 & ~x444 & ~x445 & ~x453 & ~x471 & ~x476 & ~x477 & ~x505 & ~x532 & ~x558 & ~x559 & ~x585 & ~x592 & ~x593 & ~x616 & ~x620 & ~x621 & ~x622 & ~x623 & ~x626 & ~x641 & ~x643 & ~x644 & ~x647 & ~x649 & ~x674 & ~x675 & ~x732 & ~x751 & ~x752 & ~x753 & ~x757 & ~x760 & ~x762 & ~x777 & ~x780;
assign c3480 =  x275;
assign c3482 = ~x181 & ~x249 & ~x255 & ~x317 & ~x359 & ~x428 & ~x450 & ~x453 & ~x528 & ~x529 & ~x530 & ~x561 & ~x639 & ~x764;
assign c3484 =  x36 &  x63 &  x64 &  x742 & ~x26 & ~x82 & ~x110 & ~x224 & ~x363 & ~x364 & ~x392 & ~x503 & ~x586 & ~x756 & ~x777 & ~x783;
assign c3486 =  x34;
assign c3488 =  x148 &  x149 &  x714 &  x738 &  x741 &  x743 & ~x3 & ~x24 & ~x28 & ~x30 & ~x54 & ~x57 & ~x86 & ~x109 & ~x137 & ~x138 & ~x166 & ~x170 & ~x172 & ~x194 & ~x198 & ~x201 & ~x220 & ~x222 & ~x229 & ~x248 & ~x249 & ~x278 & ~x308 & ~x337 & ~x361 & ~x368 & ~x393 & ~x394 & ~x397 & ~x416 & ~x417 & ~x424 & ~x445 & ~x446 & ~x453 & ~x473 & ~x474 & ~x476 & ~x477 & ~x481 & ~x508 & ~x536 & ~x555 & ~x556 & ~x557 & ~x560 & ~x566 & ~x583 & ~x585 & ~x587 & ~x588 & ~x591 & ~x593 & ~x622 & ~x623 & ~x637 & ~x651 & ~x665 & ~x671 & ~x694 & ~x698 & ~x703 & ~x705 & ~x727 & ~x729 & ~x753 & ~x755 & ~x778 & ~x783;
assign c3490 =  x17 &  x70 &  x546 &  x547 &  x658 &  x714 & ~x3 & ~x4 & ~x5 & ~x26 & ~x27 & ~x28 & ~x29 & ~x81 & ~x84 & ~x110 & ~x114 & ~x116 & ~x139 & ~x143 & ~x167 & ~x172 & ~x191 & ~x193 & ~x197 & ~x198 & ~x199 & ~x200 & ~x221 & ~x225 & ~x247 & ~x253 & ~x277 & ~x278 & ~x279 & ~x281 & ~x305 & ~x306 & ~x307 & ~x310 & ~x311 & ~x332 & ~x333 & ~x366 & ~x391 & ~x416 & ~x422 & ~x474 & ~x502 & ~x534 & ~x556 & ~x560 & ~x584 & ~x588 & ~x614 & ~x639 & ~x641 & ~x642 & ~x647 & ~x675 & ~x728 & ~x732 & ~x752 & ~x753 & ~x756 & ~x782;
assign c3492 = ~x2 & ~x30 & ~x84 & ~x89 & ~x116 & ~x121 & ~x133 & ~x144 & ~x164 & ~x167 & ~x205 & ~x224 & ~x246 & ~x260 & ~x273 & ~x287 & ~x299 & ~x312 & ~x329 & ~x333 & ~x336 & ~x337 & ~x340 & ~x343 & ~x356 & ~x363 & ~x370 & ~x384 & ~x385 & ~x394 & ~x398 & ~x412 & ~x426 & ~x427 & ~x445 & ~x468 & ~x475 & ~x478 & ~x481 & ~x508 & ~x528 & ~x529 & ~x534 & ~x536 & ~x537 & ~x552 & ~x554 & ~x562 & ~x563 & ~x566 & ~x588 & ~x591 & ~x615 & ~x616 & ~x646 & ~x668 & ~x704 & ~x726 & ~x730 & ~x750 & ~x763 & ~x777 & ~x783;
assign c3494 =  x124 &  x125 & ~x1 & ~x17 & ~x19 & ~x20 & ~x44 & ~x48 & ~x61 & ~x77 & ~x79 & ~x84 & ~x89 & ~x107 & ~x114 & ~x115 & ~x138 & ~x171 & ~x195 & ~x221 & ~x223 & ~x280 & ~x559 & ~x699 & ~x760 & ~x779;
assign c3496 =  x67 &  x95 &  x129 &  x130 &  x203 &  x375 &  x602 &  x766 & ~x4 & ~x20 & ~x77 & ~x109 & ~x110 & ~x145 & ~x639 & ~x672 & ~x756;
assign c3498 =  x291 & ~x8 & ~x13 & ~x14 & ~x15 & ~x20 & ~x28 & ~x32 & ~x33 & ~x53 & ~x78 & ~x83 & ~x136 & ~x139 & ~x164 & ~x165 & ~x169 & ~x204 & ~x220 & ~x221 & ~x281 & ~x282 & ~x304 & ~x308 & ~x335 & ~x339 & ~x366 & ~x392 & ~x420 & ~x502 & ~x504 & ~x529 & ~x534 & ~x559 & ~x616 & ~x619 & ~x645 & ~x700 & ~x755;
assign c31 = ~x691 & ~x739 & ~x746 & ~x765;
assign c33 =  x334;
assign c35 =  x25;
assign c37 =  x130 &  x213 &  x346 &  x354 &  x373 &  x599 &  x710 & ~x175 & ~x197 & ~x199 & ~x279 & ~x287 & ~x343 & ~x360 & ~x417 & ~x509 & ~x531 & ~x554 & ~x588 & ~x643 & ~x726 & ~x732 & ~x754;
assign c39 =  x275;
assign c311 = ~x574;
assign c313 =  x231 &  x650 & ~x117 & ~x140 & ~x163 & ~x444 & ~x451 & ~x472 & ~x501 & ~x556 & ~x724;
assign c315 =  x41 &  x44 &  x151 &  x152 &  x153 &  x154 &  x155 &  x178 &  x213 &  x235 &  x269 &  x296 &  x375 &  x380 &  x516 &  x544 &  x548 &  x656 &  x683 & ~x9 & ~x27 & ~x32 & ~x55 & ~x57 & ~x79 & ~x86 & ~x110 & ~x113 & ~x139 & ~x194 & ~x199 & ~x221 & ~x249 & ~x334 & ~x336 & ~x362 & ~x365 & ~x417 & ~x443 & ~x473 & ~x476 & ~x506 & ~x532 & ~x535 & ~x559 & ~x564 & ~x590 & ~x623 & ~x637 & ~x638 & ~x641 & ~x647 & ~x672 & ~x679 & ~x729 & ~x734 & ~x748 & ~x752 & ~x762 & ~x764 & ~x776 & ~x779;
assign c317 =  x68 & ~x518 & ~x567 & ~x770;
assign c319 =  x756;
assign c321 = ~x535 & ~x737 & ~x738 & ~x739 & ~x746;
assign c323 =  x11 &  x14 &  x15 &  x122 &  x155 &  x184 &  x211 &  x604 & ~x5 & ~x7 & ~x194 & ~x224 & ~x391 & ~x643 & ~x730;
assign c325 =  x194;
assign c327 =  x615;
assign c329 =  x257;
assign c331 =  x14 &  x15 &  x261 & ~x450;
assign c333 = ~x599 & ~x716;
assign c335 =  x108;
assign c337 =  x219;
assign c339 = ~x291 & ~x516 & ~x743;
assign c341 = ~x551 & ~x601;
assign c343 =  x617;
assign c345 =  x240 &  x269 &  x272 &  x355 &  x373 &  x383 &  x429 &  x513 &  x523 &  x568 & ~x7 & ~x21 & ~x55 & ~x84 & ~x86 & ~x198 & ~x223 & ~x251 & ~x362 & ~x363 & ~x370 & ~x391 & ~x395 & ~x398 & ~x453 & ~x477 & ~x501 & ~x526 & ~x536 & ~x537 & ~x583 & ~x610 & ~x611 & ~x612 & ~x617 & ~x640 & ~x642 & ~x668 & ~x725 & ~x752 & ~x758;
assign c347 =  x154 &  x241 &  x520 & ~x439;
assign c349 =  x344 &  x608 &  x652 & ~x12 & ~x15 & ~x422 & ~x554 & ~x582 & ~x610;
assign c351 = ~x149 & ~x347 & ~x460;
assign c353 =  x17 &  x39 & ~x456;
assign c355 =  x162 &  x230 &  x231 & ~x694;
assign c357 =  x219 &  x258 & ~x750;
assign c359 =  x169;
assign c361 =  x580 & ~x178;
assign c363 =  x148 &  x260 &  x262 &  x288 &  x316 &  x318 &  x323 &  x344 &  x348 &  x374 &  x410 &  x438 &  x465 &  x484 &  x493 &  x576 &  x606 &  x634 & ~x5 & ~x7 & ~x20 & ~x22 & ~x32 & ~x33 & ~x57 & ~x59 & ~x80 & ~x81 & ~x85 & ~x86 & ~x109 & ~x111 & ~x112 & ~x113 & ~x140 & ~x165 & ~x171 & ~x198 & ~x225 & ~x226 & ~x253 & ~x255 & ~x282 & ~x283 & ~x304 & ~x333 & ~x335 & ~x362 & ~x365 & ~x366 & ~x368 & ~x369 & ~x386 & ~x391 & ~x398 & ~x421 & ~x426 & ~x446 & ~x447 & ~x450 & ~x451 & ~x452 & ~x454 & ~x470 & ~x471 & ~x472 & ~x480 & ~x482 & ~x500 & ~x507 & ~x526 & ~x527 & ~x528 & ~x529 & ~x530 & ~x532 & ~x534 & ~x554 & ~x557 & ~x558 & ~x559 & ~x563 & ~x586 & ~x587 & ~x588 & ~x590 & ~x591 & ~x610 & ~x613 & ~x615 & ~x616 & ~x619 & ~x638 & ~x640 & ~x642 & ~x645 & ~x649 & ~x671 & ~x675 & ~x698 & ~x701 & ~x705 & ~x725 & ~x731 & ~x733 & ~x754 & ~x755 & ~x757 & ~x761;
assign c365 =  x152 &  x182 &  x235 &  x352 &  x600 & ~x137 & ~x596;
assign c367 =  x354 &  x566 &  x581 &  x594 &  x682 &  x690 & ~x162 & ~x339;
assign c369 =  x215 &  x261 &  x262 &  x264 &  x265 &  x268 &  x291 &  x292 &  x354 &  x379 &  x401 &  x429 &  x458 &  x521 &  x540 &  x569 &  x596 &  x606 &  x625 &  x662 &  x681 &  x688 &  x709 &  x739 & ~x2 & ~x5 & ~x7 & ~x21 & ~x22 & ~x50 & ~x54 & ~x79 & ~x83 & ~x87 & ~x139 & ~x164 & ~x220 & ~x225 & ~x226 & ~x229 & ~x274 & ~x278 & ~x280 & ~x302 & ~x304 & ~x308 & ~x312 & ~x313 & ~x331 & ~x358 & ~x362 & ~x363 & ~x364 & ~x366 & ~x370 & ~x385 & ~x386 & ~x397 & ~x424 & ~x441 & ~x452 & ~x470 & ~x480 & ~x498 & ~x499 & ~x500 & ~x503 & ~x504 & ~x505 & ~x527 & ~x528 & ~x533 & ~x554 & ~x558 & ~x560 & ~x587 & ~x610 & ~x612 & ~x616 & ~x619 & ~x620 & ~x638 & ~x639 & ~x647 & ~x669 & ~x675 & ~x677 & ~x697 & ~x699 & ~x756 & ~x760 & ~x761 & ~x781 & ~x782;
assign c371 =  x362;
assign c373 =  x86;
assign c375 =  x334;
assign c377 = ~x290 & ~x712;
assign c379 =  x380 & ~x658 & ~x714;
assign c381 =  x62 &  x173 &  x203;
assign c383 = ~x125;
assign c385 =  x305;
assign c387 = ~x94 & ~x744;
assign c389 =  x308;
assign c391 =  x69 &  x125 &  x126 &  x149 &  x153 &  x154 &  x157 &  x176 &  x178 &  x179 &  x180 &  x204 &  x211 &  x214 &  x233 &  x236 &  x237 &  x242 &  x261 &  x265 &  x289 &  x296 &  x299 &  x319 &  x320 &  x327 &  x345 &  x351 &  x355 &  x377 &  x378 &  x380 &  x382 &  x404 &  x407 &  x428 &  x429 &  x430 &  x431 &  x434 &  x457 &  x459 &  x462 &  x463 &  x467 &  x484 &  x485 &  x487 &  x489 &  x491 &  x492 &  x493 &  x515 &  x516 &  x517 &  x519 &  x521 &  x540 &  x541 &  x544 &  x546 &  x547 &  x549 &  x570 &  x573 &  x578 &  x579 &  x602 &  x604 &  x625 &  x626 &  x631 &  x634 &  x655 &  x656 &  x660 &  x683 &  x687 &  x717 &  x718 &  x746 & ~x0 & ~x1 & ~x2 & ~x4 & ~x7 & ~x23 & ~x25 & ~x27 & ~x29 & ~x32 & ~x50 & ~x52 & ~x53 & ~x55 & ~x58 & ~x81 & ~x85 & ~x109 & ~x113 & ~x136 & ~x138 & ~x142 & ~x165 & ~x167 & ~x191 & ~x192 & ~x194 & ~x196 & ~x197 & ~x201 & ~x219 & ~x221 & ~x253 & ~x254 & ~x255 & ~x256 & ~x278 & ~x281 & ~x282 & ~x306 & ~x308 & ~x311 & ~x336 & ~x364 & ~x368 & ~x388 & ~x393 & ~x394 & ~x417 & ~x422 & ~x446 & ~x450 & ~x451 & ~x472 & ~x473 & ~x478 & ~x504 & ~x507 & ~x528 & ~x531 & ~x532 & ~x534 & ~x535 & ~x556 & ~x559 & ~x561 & ~x584 & ~x587 & ~x588 & ~x592 & ~x613 & ~x620 & ~x641 & ~x646 & ~x668 & ~x670 & ~x671 & ~x674 & ~x676 & ~x696 & ~x703 & ~x724 & ~x726 & ~x752 & ~x757 & ~x758 & ~x759 & ~x781;
assign c393 = ~x148 & ~x630 & ~x708;
assign c395 =  x762;
assign c397 =  x334;
assign c399 =  x477;
assign c3101 =  x221;
assign c3103 =  x130 &  x212 &  x234 &  x236 &  x269 &  x270 &  x297 &  x318 &  x326 &  x354 &  x408 &  x410 & ~x62 & ~x80 & ~x116 & ~x118 & ~x163 & ~x167 & ~x218 & ~x257 & ~x315 & ~x359 & ~x365 & ~x469 & ~x528 & ~x538 & ~x554 & ~x557 & ~x609 & ~x637 & ~x750;
assign c3105 =  x672;
assign c3107 =  x364;
assign c3109 =  x24;
assign c3111 =  x45 &  x153 &  x155 &  x176 &  x180 &  x182 &  x186 &  x204 &  x206 &  x209 &  x260 &  x261 &  x262 &  x265 &  x266 &  x271 &  x288 &  x290 &  x293 &  x298 &  x299 &  x317 &  x320 &  x321 &  x323 &  x325 &  x353 &  x355 &  x373 &  x381 &  x401 &  x402 &  x403 &  x411 &  x439 &  x458 &  x463 &  x464 &  x465 &  x467 &  x485 &  x492 &  x493 &  x519 &  x520 &  x540 &  x544 &  x550 &  x551 &  x568 &  x569 &  x571 &  x579 &  x599 &  x603 &  x626 &  x663 &  x688 & ~x2 & ~x6 & ~x21 & ~x27 & ~x29 & ~x53 & ~x55 & ~x58 & ~x60 & ~x81 & ~x83 & ~x86 & ~x110 & ~x138 & ~x143 & ~x166 & ~x170 & ~x196 & ~x222 & ~x226 & ~x229 & ~x253 & ~x254 & ~x279 & ~x307 & ~x336 & ~x362 & ~x364 & ~x366 & ~x417 & ~x418 & ~x419 & ~x445 & ~x447 & ~x449 & ~x450 & ~x473 & ~x501 & ~x503 & ~x505 & ~x506 & ~x508 & ~x534 & ~x557 & ~x558 & ~x564 & ~x590 & ~x591 & ~x611 & ~x613 & ~x615 & ~x620 & ~x640 & ~x644 & ~x647 & ~x668 & ~x672 & ~x696 & ~x700 & ~x702 & ~x704 & ~x726 & ~x728 & ~x758 & ~x760 & ~x780;
assign c3113 =  x611 &  x667;
assign c3115 =  x220;
assign c3117 = ~x177 & ~x233;
assign c3119 =  x106 &  x203 & ~x750;
assign c3121 =  x400 &  x482 &  x566 &  x597 &  x656 &  x662 & ~x10 & ~x18 & ~x36 & ~x84 & ~x173 & ~x615;
assign c3123 =  x583;
assign c3125 = ~x235 & ~x319 & ~x544 & ~x627;
assign c3127 =  x170;
assign c3129 =  x296 & ~x511 & ~x596 & ~x607;
assign c3131 = ~x11 & ~x12 & ~x122 & ~x178 & ~x205;
assign c3133 =  x543 & ~x630 & ~x658;
assign c3135 =  x221;
assign c3137 =  x206 &  x213 &  x239 &  x240 &  x269 &  x320 &  x325 &  x352 &  x380 &  x381 &  x409 &  x515 &  x655 & ~x6 & ~x52 & ~x58 & ~x63 & ~x88 & ~x106 & ~x135 & ~x138 & ~x139 & ~x173 & ~x189 & ~x198 & ~x199 & ~x217 & ~x218 & ~x222 & ~x228 & ~x248 & ~x255 & ~x258 & ~x311 & ~x312 & ~x313 & ~x314 & ~x358 & ~x362 & ~x367 & ~x369 & ~x370 & ~x371 & ~x389 & ~x421 & ~x426 & ~x427 & ~x441 & ~x452 & ~x470 & ~x509 & ~x529 & ~x532 & ~x554 & ~x594 & ~x610 & ~x616 & ~x618 & ~x619 & ~x622 & ~x650 & ~x701 & ~x723 & ~x731 & ~x750 & ~x753 & ~x756;
assign c3139 =  x102 &  x150 &  x158 &  x178 &  x179 &  x206 &  x213 &  x234 &  x236 &  x239 &  x241 &  x262 &  x268 &  x297 &  x325 &  x375 &  x376 &  x515 & ~x6 & ~x22 & ~x49 & ~x80 & ~x83 & ~x90 & ~x108 & ~x109 & ~x110 & ~x114 & ~x141 & ~x146 & ~x170 & ~x173 & ~x191 & ~x217 & ~x250 & ~x255 & ~x258 & ~x310 & ~x315 & ~x331 & ~x341 & ~x398 & ~x415 & ~x417 & ~x418 & ~x426 & ~x478 & ~x480 & ~x497 & ~x507 & ~x508 & ~x537 & ~x556 & ~x582 & ~x586 & ~x612 & ~x621 & ~x669 & ~x674 & ~x695 & ~x703 & ~x752;
assign c3141 = ~x602 & ~x658 & ~x714 & ~x742;
assign c3143 =  x29;
assign c3145 = ~x511 & ~x602 & ~x658 & ~x663;
assign c3147 =  x689 & ~x490 & ~x518 & ~x552 & ~x630;
assign c3149 =  x178 &  x240 &  x268 &  x290 &  x297 &  x318 &  x407 & ~x8 & ~x23 & ~x79 & ~x162 & ~x252 & ~x255 & ~x315 & ~x371 & ~x392 & ~x398 & ~x441 & ~x503 & ~x565 & ~x617 & ~x618 & ~x646 & ~x666 & ~x670 & ~x759 & ~x781;
assign c3151 = ~x16 & ~x181;
assign c3153 = ~x178 & ~x209;
assign c3155 = ~x205 & ~x460;
assign c3157 =  x132 &  x202 &  x230 &  x270 &  x287 &  x327 & ~x10 & ~x422;
assign c3159 =  x213 &  x236 &  x269 &  x324 &  x408 & ~x76 & ~x77 & ~x110 & ~x115 & ~x133 & ~x188 & ~x328 & ~x384 & ~x440 & ~x455 & ~x498 & ~x510 & ~x558 & ~x615 & ~x620 & ~x650 & ~x727 & ~x780;
assign c3161 =  x87;
assign c3163 =  x41 &  x42 &  x45 &  x70 &  x72 &  x94 &  x127 &  x153 &  x177 &  x178 &  x179 &  x182 &  x234 &  x239 &  x261 &  x262 &  x270 &  x289 &  x291 &  x297 &  x348 &  x353 &  x376 &  x401 &  x408 &  x429 &  x431 &  x432 &  x436 &  x438 &  x464 &  x465 &  x466 &  x494 &  x520 &  x522 &  x543 &  x549 &  x578 &  x632 &  x634 &  x655 &  x661 &  x688 &  x710 &  x711 &  x717 &  x718 & ~x21 & ~x22 & ~x23 & ~x24 & ~x25 & ~x26 & ~x50 & ~x54 & ~x56 & ~x85 & ~x86 & ~x110 & ~x112 & ~x136 & ~x140 & ~x145 & ~x170 & ~x191 & ~x198 & ~x219 & ~x246 & ~x281 & ~x285 & ~x303 & ~x306 & ~x313 & ~x367 & ~x392 & ~x393 & ~x419 & ~x423 & ~x451 & ~x506 & ~x527 & ~x529 & ~x583 & ~x584 & ~x588 & ~x592 & ~x611 & ~x615 & ~x618 & ~x620 & ~x668 & ~x696 & ~x703 & ~x704 & ~x725 & ~x750 & ~x753 & ~x763 & ~x778;
assign c3165 =  x257 &  x620;
assign c3167 =  x90 &  x231 & ~x6 & ~x722;
assign c3169 = ~x149 & ~x153 & ~x292 & ~x295;
assign c3171 =  x340;
assign c3173 = ~x126 & ~x130 & ~x187 & ~x265;
assign c3175 =  x220;
assign c3177 =  x424;
assign c3179 =  x136;
assign c3181 =  x222;
assign c3183 =  x224;
assign c3185 =  x700;
assign c3187 =  x177 &  x238 &  x243 &  x268 &  x293 &  x319 &  x327 &  x348 &  x349 &  x354 &  x372 &  x375 &  x377 &  x380 &  x381 &  x402 &  x429 &  x431 &  x457 &  x458 &  x465 &  x484 &  x512 &  x520 &  x540 &  x547 &  x605 &  x663 &  x689 & ~x17 & ~x22 & ~x23 & ~x26 & ~x30 & ~x86 & ~x111 & ~x168 & ~x172 & ~x192 & ~x197 & ~x222 & ~x253 & ~x280 & ~x306 & ~x307 & ~x332 & ~x339 & ~x421 & ~x446 & ~x499 & ~x527 & ~x528 & ~x530 & ~x587 & ~x614 & ~x618 & ~x641 & ~x704 & ~x723 & ~x752 & ~x755;
assign c3189 = ~x75 & ~x153 & ~x160 & ~x205;
assign c3191 = ~x130 & ~x544;
assign c3193 = ~x207 & ~x263;
assign c3197 =  x442 &  x510 &  x594 &  x610 & ~x145;
assign c3199 =  x45 &  x130 &  x182 &  x185 &  x186 &  x210 &  x211 &  x212 &  x237 &  x296 &  x516 & ~x62 & ~x88 & ~x113 & ~x133 & ~x138 & ~x161 & ~x163 & ~x195 & ~x224 & ~x228 & ~x230 & ~x245 & ~x250 & ~x333 & ~x337 & ~x356 & ~x369 & ~x394 & ~x397 & ~x415 & ~x445 & ~x509 & ~x531 & ~x618 & ~x704 & ~x730 & ~x751;
assign c3201 =  x233 &  x271 &  x299 &  x323 &  x383 &  x405 &  x431 &  x436 &  x458 &  x465 &  x487 &  x488 &  x550 &  x633 &  x661 &  x662 &  x709 &  x715 &  x771 & ~x6 & ~x21 & ~x53 & ~x57 & ~x170 & ~x192 & ~x195 & ~x201 & ~x254 & ~x274 & ~x306 & ~x360 & ~x364 & ~x365 & ~x368 & ~x398 & ~x425 & ~x442 & ~x445 & ~x450 & ~x472 & ~x498 & ~x502 & ~x506 & ~x508 & ~x558 & ~x561 & ~x563 & ~x582 & ~x583 & ~x588 & ~x614 & ~x639 & ~x666 & ~x671 & ~x674 & ~x726 & ~x728 & ~x733 & ~x750;
assign c3203 =  x193;
assign c3205 =  x639;
assign c3207 =  x234 & ~x686 & ~x742;
assign c3209 =  x249;
assign c3211 =  x275;
assign c3213 =  x672;
assign c3215 =  x85;
assign c3217 =  x329 &  x386 &  x498 &  x554 &  x610;
assign c3219 = ~x319 & ~x404;
assign c3221 =  x198;
assign c3225 =  x130 &  x149 &  x177 &  x232 &  x234 &  x239 &  x289 &  x292 &  x297 &  x299 &  x324 &  x345 &  x348 &  x353 &  x375 &  x409 &  x520 &  x571 &  x606 &  x655 &  x662 & ~x7 & ~x23 & ~x31 & ~x32 & ~x51 & ~x81 & ~x174 & ~x225 & ~x229 & ~x250 & ~x258 & ~x279 & ~x302 & ~x307 & ~x310 & ~x340 & ~x360 & ~x368 & ~x385 & ~x421 & ~x425 & ~x502 & ~x506 & ~x535 & ~x554 & ~x557 & ~x559 & ~x562 & ~x565 & ~x592 & ~x646 & ~x649 & ~x671 & ~x700 & ~x702 & ~x723 & ~x727 & ~x732 & ~x751 & ~x753;
assign c3227 =  x90 & ~x666;
assign c3229 =  x191;
assign c3231 =  x308;
assign c3233 =  x70 & ~x461 & ~x489;
assign c3235 =  x244 &  x289 &  x406 &  x541 &  x637 & ~x169 & ~x170 & ~x332 & ~x359 & ~x387 & ~x419 & ~x471 & ~x534 & ~x535 & ~x591 & ~x724 & ~x732;
assign c3237 =  x68 &  x101 &  x131 &  x155 &  x156 &  x181 &  x185 &  x243 &  x262 &  x263 &  x271 &  x289 &  x318 &  x327 &  x345 &  x348 &  x351 &  x375 &  x404 &  x429 &  x431 &  x438 &  x439 &  x458 &  x492 &  x514 &  x519 &  x541 &  x542 &  x548 &  x550 &  x597 &  x598 &  x599 &  x661 &  x662 &  x712 &  x717 & ~x28 & ~x31 & ~x32 & ~x54 & ~x85 & ~x138 & ~x142 & ~x198 & ~x221 & ~x225 & ~x249 & ~x282 & ~x306 & ~x307 & ~x334 & ~x363 & ~x366 & ~x367 & ~x385 & ~x387 & ~x388 & ~x392 & ~x393 & ~x416 & ~x421 & ~x424 & ~x425 & ~x442 & ~x446 & ~x451 & ~x452 & ~x477 & ~x480 & ~x527 & ~x530 & ~x531 & ~x533 & ~x535 & ~x554 & ~x556 & ~x557 & ~x560 & ~x561 & ~x584 & ~x588 & ~x592 & ~x610 & ~x613 & ~x614 & ~x617 & ~x642 & ~x643 & ~x649 & ~x671 & ~x674 & ~x677 & ~x700 & ~x703 & ~x750 & ~x752 & ~x755 & ~x757 & ~x759 & ~x782;
assign c3239 =  x309;
assign c3241 =  x129 &  x131 &  x151 &  x153 &  x154 &  x156 &  x158 &  x159 &  x180 &  x181 &  x186 &  x208 &  x236 &  x239 &  x240 &  x261 &  x270 &  x271 &  x296 &  x298 &  x320 &  x324 &  x352 &  x354 &  x374 &  x376 &  x409 &  x432 &  x437 &  x458 &  x464 &  x465 &  x515 &  x543 &  x570 &  x571 &  x577 &  x662 & ~x6 & ~x7 & ~x54 & ~x87 & ~x141 & ~x165 & ~x220 & ~x223 & ~x278 & ~x281 & ~x339 & ~x357 & ~x441 & ~x449 & ~x498 & ~x502 & ~x507 & ~x528 & ~x534 & ~x555 & ~x559 & ~x594 & ~x610 & ~x612 & ~x638 & ~x670 & ~x727 & ~x730 & ~x755 & ~x757 & ~x761 & ~x777;
assign c3243 =  x592;
assign c3245 =  x627 & ~x630 & ~x658;
assign c3247 =  x270 &  x326 &  x465 & ~x658;
assign c3249 = ~x47 & ~x178 & ~x295;
assign c3251 = ~x75 & ~x151 & ~x205 & ~x206;
assign c3253 =  x203 &  x622 & ~x191 & ~x367 & ~x479 & ~x724;
assign c3255 = ~x148 & ~x462 & ~x490 & ~x518 & ~x574 & ~x602;
assign c3257 =  x762;
assign c3259 =  x315 & ~x9 & ~x18 & ~x256 & ~x394 & ~x420 & ~x644 & ~x766 & ~x772 & ~x773 & ~x774;
assign c3261 =  x259 &  x734;
assign c3263 = ~x658 & ~x686 & ~x742 & ~x769;
assign c3265 =  x313 &  x648;
assign c3267 = ~x745;
assign c3269 =  x781;
assign c3271 = ~x12 & ~x75 & ~x178;
assign c3273 = ~x630;
assign c3275 = ~x11 & ~x75 & ~x209;
assign c3277 =  x44 &  x96 &  x152 &  x156 &  x235 &  x297 &  x325 &  x459 &  x515 & ~x4 & ~x9 & ~x36 & ~x64 & ~x76 & ~x80 & ~x222 & ~x312 & ~x336 & ~x417 & ~x449 & ~x474 & ~x533 & ~x646 & ~x702 & ~x727 & ~x736 & ~x765;
assign c3279 =  x645;
assign c3281 =  x118 &  x230 &  x260 &  x274 &  x323 &  x381 & ~x446;
assign c3283 =  x778;
assign c3285 =  x288 &  x345 &  x346 &  x372 &  x374 &  x375 &  x380 &  x400 &  x407 &  x409 &  x429 &  x484 &  x490 &  x522 &  x547 &  x575 &  x577 &  x597 &  x606 &  x653 &  x662 &  x684 &  x688 &  x690 & ~x5 & ~x10 & ~x26 & ~x27 & ~x29 & ~x32 & ~x37 & ~x81 & ~x108 & ~x117 & ~x141 & ~x143 & ~x145 & ~x167 & ~x171 & ~x280 & ~x307 & ~x360 & ~x365 & ~x391 & ~x396 & ~x420 & ~x421 & ~x424 & ~x444 & ~x446 & ~x450 & ~x451 & ~x507 & ~x529 & ~x535 & ~x562 & ~x586 & ~x587 & ~x644 & ~x675 & ~x727;
assign c3287 = ~x130 & ~x215 & ~x235;
assign c3289 =  x639;
assign c3291 =  x0;
assign c3293 =  x717 & ~x518;
assign c3295 =  x257;
assign c3297 =  x212 &  x240 &  x241 &  x267 &  x684 & ~x174 & ~x175 & ~x231 & ~x288 & ~x316 & ~x539;
assign c3299 =  x45 &  x70 &  x101 &  x129 &  x130 &  x152 &  x157 &  x158 &  x180 &  x181 &  x182 &  x183 &  x184 &  x208 &  x211 &  x214 &  x235 &  x236 &  x241 &  x262 &  x264 &  x269 &  x296 &  x318 &  x347 &  x374 &  x380 &  x381 &  x408 &  x431 &  x487 &  x516 &  x543 &  x571 &  x628 & ~x6 & ~x7 & ~x8 & ~x20 & ~x24 & ~x30 & ~x33 & ~x34 & ~x50 & ~x53 & ~x56 & ~x57 & ~x80 & ~x83 & ~x85 & ~x107 & ~x109 & ~x115 & ~x116 & ~x117 & ~x118 & ~x134 & ~x137 & ~x141 & ~x143 & ~x145 & ~x162 & ~x163 & ~x168 & ~x171 & ~x191 & ~x219 & ~x220 & ~x222 & ~x224 & ~x229 & ~x230 & ~x247 & ~x253 & ~x256 & ~x280 & ~x282 & ~x285 & ~x305 & ~x306 & ~x308 & ~x311 & ~x313 & ~x334 & ~x336 & ~x338 & ~x339 & ~x340 & ~x341 & ~x360 & ~x361 & ~x365 & ~x389 & ~x391 & ~x393 & ~x394 & ~x418 & ~x419 & ~x422 & ~x423 & ~x424 & ~x444 & ~x449 & ~x472 & ~x479 & ~x504 & ~x530 & ~x533 & ~x534 & ~x536 & ~x559 & ~x561 & ~x562 & ~x563 & ~x587 & ~x591 & ~x613 & ~x621 & ~x642 & ~x645 & ~x647 & ~x677 & ~x693 & ~x696 & ~x697 & ~x699 & ~x704 & ~x706 & ~x722 & ~x725 & ~x731 & ~x733 & ~x750 & ~x755 & ~x758 & ~x776 & ~x783;
assign c3301 =  x399 &  x489 &  x577 &  x578 & ~x10 & ~x11 & ~x36 & ~x37 & ~x46 & ~x65 & ~x76 & ~x117;
assign c3303 =  x182 & ~x272 & ~x344;
assign c3305 =  x110;
assign c3307 =  x32;
assign c3309 = ~x214 & ~x237 & ~x321;
assign c3311 =  x583;
assign c3313 =  x25;
assign c3315 =  x9;
assign c3317 =  x90 &  x203 &  x272 & ~x471 & ~x510;
assign c3319 =  x203 &  x622 & ~x60 & ~x228 & ~x528;
assign c3321 =  x30;
assign c3323 =  x198;
assign c3325 =  x8;
assign c3327 =  x25;
assign c3329 =  x44 &  x182 &  x684 & ~x512 & ~x720 & ~x724;
assign c3331 =  x303 &  x703;
assign c3333 =  x204 &  x299 &  x345 &  x373 &  x409 &  x429 &  x433 &  x460 &  x608 &  x626 & ~x51 & ~x82 & ~x111 & ~x144 & ~x218 & ~x220 & ~x364 & ~x481 & ~x561 & ~x701 & ~x753;
assign c3335 = ~x75 & ~x181 & ~x293;
assign c3337 =  x639;
assign c3339 =  x727;
assign c3341 = ~x635 & ~x739 & ~x746;
assign c3343 =  x354 &  x547 &  x580 &  x595 &  x597 &  x684 &  x708 & ~x17 & ~x51 & ~x55 & ~x201 & ~x250;
assign c3345 =  x440 &  x608 &  x609 &  x636 &  x637 &  x708 &  x710 & ~x32 & ~x140 & ~x337 & ~x363 & ~x472 & ~x563 & ~x584 & ~x620 & ~x704 & ~x724;
assign c3347 = ~x235 & ~x601;
assign c3349 =  x670;
assign c3351 =  x76 &  x316 &  x428 &  x540 &  x743 & ~x12 & ~x582;
assign c3353 =  x279;
assign c3355 =  x39 &  x40 &  x41 &  x42 &  x96 &  x101 &  x102 &  x126 &  x127 &  x154 &  x157 &  x182 &  x183 &  x206 &  x234 &  x240 &  x241 &  x242 &  x290 &  x297 &  x318 &  x320 &  x323 &  x325 &  x347 &  x351 &  x375 &  x380 &  x403 &  x459 &  x486 &  x543 &  x570 &  x599 &  x627 & ~x27 & ~x28 & ~x30 & ~x79 & ~x80 & ~x85 & ~x109 & ~x110 & ~x111 & ~x143 & ~x164 & ~x171 & ~x196 & ~x224 & ~x227 & ~x248 & ~x249 & ~x252 & ~x253 & ~x276 & ~x389 & ~x390 & ~x474 & ~x526 & ~x560 & ~x561 & ~x581 & ~x588 & ~x614 & ~x616 & ~x637 & ~x647 & ~x665 & ~x693 & ~x697 & ~x707 & ~x725 & ~x728 & ~x729 & ~x754 & ~x758 & ~x760;
assign c3357 =  x355 &  x441 &  x465 & ~x47 & ~x145 & ~x253 & ~x759;
assign c3359 =  x67 &  x157 &  x181 &  x182 &  x206 &  x211 &  x214 &  x234 &  x262 &  x263 &  x264 &  x269 &  x290 &  x291 &  x298 &  x345 &  x346 &  x353 &  x410 &  x431 &  x432 &  x493 &  x548 &  x550 &  x599 & ~x3 & ~x7 & ~x24 & ~x26 & ~x51 & ~x80 & ~x88 & ~x109 & ~x166 & ~x171 & ~x174 & ~x193 & ~x197 & ~x201 & ~x202 & ~x220 & ~x225 & ~x227 & ~x248 & ~x251 & ~x254 & ~x255 & ~x256 & ~x258 & ~x274 & ~x280 & ~x281 & ~x286 & ~x309 & ~x311 & ~x313 & ~x335 & ~x336 & ~x338 & ~x357 & ~x363 & ~x385 & ~x392 & ~x394 & ~x397 & ~x447 & ~x473 & ~x475 & ~x508 & ~x509 & ~x525 & ~x529 & ~x555 & ~x557 & ~x558 & ~x566 & ~x585 & ~x590 & ~x614 & ~x638 & ~x648 & ~x666 & ~x676 & ~x702 & ~x727 & ~x731 & ~x732 & ~x752 & ~x753 & ~x755 & ~x760 & ~x782;
assign c3361 = ~x47 & ~x159 & ~x177 & ~x209 & ~x265;
assign c3365 =  x561;
assign c3367 =  x407 & ~x718 & ~x746 & ~x770;
assign c3369 =  x258 &  x621 & ~x765 & ~x766;
assign c3371 =  x13 &  x97 & ~x742;
assign c3373 =  x562;
assign c3375 = ~x740 & ~x746;
assign c3377 =  x90 &  x259 & ~x553;
assign c3381 =  x40 &  x68 &  x69 &  x125 &  x127 & ~x6 & ~x7 & ~x37 & ~x47 & ~x49 & ~x254 & ~x255 & ~x278 & ~x283 & ~x307 & ~x309 & ~x311 & ~x334 & ~x335 & ~x338 & ~x361 & ~x362 & ~x365 & ~x389 & ~x450 & ~x472 & ~x477 & ~x500 & ~x506 & ~x528 & ~x529 & ~x612 & ~x645 & ~x669 & ~x696 & ~x735 & ~x736 & ~x764 & ~x765 & ~x774 & ~x775;
assign c3383 = ~x37 & ~x159 & ~x209;
assign c3385 =  x84;
assign c3387 =  x700;
assign c3389 =  x66 &  x70 &  x409;
assign c3391 = ~x130 & ~x235 & ~x711;
assign c3393 =  x275;
assign c3395 =  x256;
assign c3397 = ~x148 & ~x178;
assign c3399 = ~x208 & ~x324;
assign c3401 = ~x517 & ~x573 & ~x600;
assign c3403 =  x205 &  x261 &  x271 &  x299 &  x347 &  x348 &  x349 &  x350 &  x354 &  x402 &  x403 &  x407 &  x515 &  x540 &  x568 &  x571 &  x627 &  x635 &  x655 & ~x0 & ~x4 & ~x6 & ~x21 & ~x88 & ~x109 & ~x110 & ~x142 & ~x143 & ~x168 & ~x224 & ~x226 & ~x281 & ~x386 & ~x397 & ~x398 & ~x416 & ~x452 & ~x469 & ~x470 & ~x497 & ~x498 & ~x509 & ~x510 & ~x528 & ~x535 & ~x537 & ~x557 & ~x560 & ~x566 & ~x585 & ~x587 & ~x592 & ~x593 & ~x616 & ~x621 & ~x672 & ~x694 & ~x697 & ~x699 & ~x702 & ~x752 & ~x754;
assign c3405 =  x203 &  x301 &  x329 &  x594 &  x622 & ~x117 & ~x472 & ~x556;
assign c3407 =  x273 & ~x623;
assign c3409 =  x476;
assign c3411 = ~x122 & ~x717 & ~x740;
assign c3413 =  x182 &  x184 &  x186 &  x208 &  x212 &  x213 &  x297 &  x319 &  x324 &  x352 &  x381 &  x432 &  x460 &  x464 &  x544 &  x604 &  x632 &  x688 & ~x21 & ~x52 & ~x88 & ~x109 & ~x111 & ~x175 & ~x259 & ~x307 & ~x313 & ~x314 & ~x330 & ~x335 & ~x369 & ~x371 & ~x393 & ~x419 & ~x443 & ~x531 & ~x535 & ~x565 & ~x582 & ~x590 & ~x591 & ~x617 & ~x618 & ~x620 & ~x639 & ~x641 & ~x642 & ~x650 & ~x675 & ~x698 & ~x699 & ~x727 & ~x728 & ~x734 & ~x760 & ~x781;
assign c3415 =  x695;
assign c3417 =  x176 &  x185 &  x187 &  x204 &  x232 &  x236 &  x240 &  x241 &  x260 &  x290 &  x291 &  x293 &  x296 &  x299 &  x316 &  x321 &  x345 &  x374 &  x379 &  x400 &  x401 &  x407 &  x411 &  x456 &  x468 &  x485 &  x495 &  x496 &  x523 &  x569 &  x574 &  x578 &  x597 &  x602 &  x604 &  x633 &  x683 &  x711 &  x712 &  x744 & ~x25 & ~x30 & ~x33 & ~x51 & ~x53 & ~x56 & ~x79 & ~x86 & ~x117 & ~x136 & ~x138 & ~x144 & ~x165 & ~x193 & ~x197 & ~x225 & ~x226 & ~x229 & ~x252 & ~x253 & ~x256 & ~x281 & ~x282 & ~x311 & ~x312 & ~x332 & ~x338 & ~x341 & ~x359 & ~x369 & ~x416 & ~x474 & ~x475 & ~x476 & ~x501 & ~x502 & ~x505 & ~x507 & ~x529 & ~x531 & ~x532 & ~x591 & ~x612 & ~x619 & ~x643 & ~x648 & ~x669 & ~x672 & ~x698 & ~x704 & ~x728 & ~x754 & ~x757 & ~x758 & ~x760 & ~x781 & ~x782 & ~x783;
assign c3419 = ~x602 & ~x658 & ~x742;
assign c3421 =  x96 &  x98 &  x177 &  x204 &  x232 &  x236 &  x237 &  x238 &  x240 &  x241 &  x261 &  x266 &  x270 &  x271 &  x289 &  x317 &  x322 &  x323 &  x347 &  x382 &  x401 &  x405 &  x430 &  x438 &  x466 &  x494 &  x513 &  x514 &  x519 &  x569 &  x597 &  x599 &  x600 &  x601 &  x603 &  x605 &  x626 &  x634 &  x683 &  x690 &  x745 &  x768 &  x771 & ~x1 & ~x5 & ~x6 & ~x7 & ~x24 & ~x26 & ~x28 & ~x29 & ~x53 & ~x56 & ~x86 & ~x110 & ~x115 & ~x195 & ~x197 & ~x198 & ~x221 & ~x222 & ~x224 & ~x252 & ~x254 & ~x280 & ~x307 & ~x309 & ~x311 & ~x334 & ~x336 & ~x337 & ~x363 & ~x387 & ~x388 & ~x391 & ~x392 & ~x421 & ~x422 & ~x444 & ~x447 & ~x449 & ~x471 & ~x498 & ~x501 & ~x502 & ~x527 & ~x534 & ~x584 & ~x593 & ~x610 & ~x614 & ~x615 & ~x616 & ~x617 & ~x639 & ~x643 & ~x647 & ~x666 & ~x671 & ~x696 & ~x698 & ~x699 & ~x704 & ~x727 & ~x752 & ~x754 & ~x756 & ~x757 & ~x783;
assign c3423 =  x230 & ~x358 & ~x413;
assign c3425 =  x157 &  x159 &  x204 &  x232 &  x243 &  x290 &  x296 &  x319 &  x355 &  x372 &  x407 &  x411 &  x434 &  x464 &  x485 &  x494 &  x512 &  x569 &  x570 &  x575 &  x682 &  x718 & ~x2 & ~x7 & ~x28 & ~x54 & ~x59 & ~x115 & ~x139 & ~x143 & ~x166 & ~x199 & ~x221 & ~x223 & ~x248 & ~x252 & ~x254 & ~x255 & ~x365 & ~x396 & ~x398 & ~x426 & ~x443 & ~x445 & ~x453 & ~x471 & ~x473 & ~x537 & ~x617 & ~x639 & ~x675 & ~x700 & ~x751 & ~x753;
assign c3427 =  x71 &  x184 &  x186 &  x210 &  x232 &  x236 &  x242 &  x243 &  x265 &  x267 &  x271 &  x287 &  x298 &  x315 &  x323 &  x327 &  x343 &  x344 &  x345 &  x355 &  x371 &  x381 &  x405 &  x406 &  x409 &  x427 &  x434 &  x456 &  x461 &  x483 &  x497 &  x514 &  x516 &  x519 &  x550 &  x572 &  x581 &  x599 &  x605 &  x628 &  x655 &  x688 &  x690 &  x711 & ~x22 & ~x55 & ~x60 & ~x87 & ~x109 & ~x113 & ~x135 & ~x168 & ~x169 & ~x197 & ~x200 & ~x223 & ~x275 & ~x279 & ~x284 & ~x366 & ~x395 & ~x419 & ~x449 & ~x500 & ~x504 & ~x507 & ~x528 & ~x529 & ~x560 & ~x563 & ~x585 & ~x588 & ~x670 & ~x671 & ~x701 & ~x724 & ~x726 & ~x730 & ~x755 & ~x756;
assign c3429 =  x171;
assign c3431 =  x219;
assign c3433 =  x40 &  x99 &  x123 &  x152 &  x177 &  x182 &  x204 &  x207 &  x208 &  x214 &  x233 &  x234 &  x236 &  x242 &  x261 &  x263 &  x265 &  x266 &  x269 &  x271 &  x290 &  x291 &  x294 &  x297 &  x298 &  x299 &  x300 &  x317 &  x320 &  x325 &  x327 &  x348 &  x373 &  x403 &  x407 &  x408 &  x437 &  x460 &  x489 &  x513 &  x516 &  x517 &  x518 &  x544 &  x545 &  x547 &  x571 &  x576 &  x598 &  x599 &  x604 &  x627 &  x629 &  x630 &  x684 &  x689 &  x713 & ~x6 & ~x10 & ~x21 & ~x23 & ~x35 & ~x36 & ~x51 & ~x57 & ~x59 & ~x80 & ~x82 & ~x110 & ~x112 & ~x113 & ~x137 & ~x138 & ~x141 & ~x142 & ~x144 & ~x145 & ~x168 & ~x172 & ~x194 & ~x196 & ~x220 & ~x278 & ~x307 & ~x309 & ~x311 & ~x334 & ~x337 & ~x361 & ~x365 & ~x366 & ~x394 & ~x417 & ~x418 & ~x420 & ~x421 & ~x422 & ~x423 & ~x446 & ~x451 & ~x503 & ~x505 & ~x506 & ~x529 & ~x535 & ~x588 & ~x613 & ~x615 & ~x617 & ~x618 & ~x643 & ~x646 & ~x675 & ~x698 & ~x727 & ~x729 & ~x731 & ~x782 & ~x783;
assign c3435 = ~x37 & ~x215 & ~x319 & ~x353;
assign c3437 = ~x206 & ~x233;
assign c3439 =  x454 &  x594 & ~x9 & ~x36 & ~x55 & ~x145 & ~x172 & ~x502 & ~x756;
assign c3441 = ~x549 & ~x550 & ~x772;
assign c3443 =  x604 &  x772 & ~x64 & ~x92 & ~x120 & ~x146 & ~x148 & ~x160 & ~x328 & ~x440 & ~x722;
assign c3445 =  x90 &  x117 &  x118 &  x202 & ~x764;
assign c3447 =  x45 &  x326 &  x345 &  x355 &  x373 &  x375 &  x466 &  x486 &  x488 &  x521 &  x551 &  x552 &  x634 &  x689 &  x745 & ~x18 & ~x22 & ~x90 & ~x112 & ~x115 & ~x168 & ~x198 & ~x225 & ~x251 & ~x255 & ~x277 & ~x280 & ~x304 & ~x333 & ~x334 & ~x389 & ~x420 & ~x422 & ~x450 & ~x500 & ~x530 & ~x560 & ~x646 & ~x696 & ~x730;
assign c3449 = ~x63 & ~x147 & ~x287 & ~x328 & ~x567 & ~x734;
assign c3451 =  x126 &  x182 &  x295 &  x296 &  x297 &  x487 &  x632 & ~x63 & ~x91 & ~x175 & ~x203 & ~x246 & ~x247 & ~x274 & ~x283 & ~x340 & ~x391 & ~x441 & ~x503 & ~x588 & ~x622 & ~x667 & ~x695 & ~x750 & ~x782;
assign c3453 =  x171;
assign c3455 =  x191;
assign c3457 =  x667;
assign c3459 =  x373 & ~x46 & ~x157;
assign c3461 =  x354 &  x373 &  x381 &  x400 &  x461 &  x466 &  x468 &  x485 &  x493 &  x496 &  x522 &  x544 &  x545 &  x550 &  x600 &  x602 &  x603 &  x605 &  x626 &  x627 &  x628 &  x661 &  x662 &  x715 & ~x0 & ~x3 & ~x5 & ~x37 & ~x54 & ~x60 & ~x63 & ~x112 & ~x113 & ~x116 & ~x140 & ~x170 & ~x171 & ~x194 & ~x197 & ~x249 & ~x310 & ~x389 & ~x390 & ~x419 & ~x420 & ~x474 & ~x534 & ~x557 & ~x641 & ~x643 & ~x699 & ~x780 & ~x783;
assign c3463 =  x761;
assign c3465 =  x565 &  x694;
assign c3467 = ~x17 & ~x75 & ~x121 & ~x209;
assign c3469 =  x223;
assign c3471 = ~x518 & ~x574 & ~x595;
assign c3473 =  x561;
assign c3475 =  x778;
assign c3477 =  x159 & ~x133 & ~x273 & ~x384 & ~x412;
assign c3479 =  x173 &  x202 & ~x509 & ~x537 & ~x554;
assign c3481 = ~x518 & ~x574 & ~x743;
assign c3483 =  x14 &  x39 & ~x91;
assign c3485 =  x106 &  x231 & ~x414 & ~x610;
assign c3487 =  x532;
assign c3489 =  x92 &  x201 &  x246 &  x259 & ~x361;
assign c3491 = ~x149 & ~x179;
assign c3493 =  x40 &  x67 &  x152 &  x153 &  x179 &  x319 &  x323 &  x325 &  x346 &  x431 &  x599 & ~x6 & ~x7 & ~x8 & ~x30 & ~x32 & ~x34 & ~x51 & ~x80 & ~x111 & ~x138 & ~x143 & ~x170 & ~x193 & ~x277 & ~x280 & ~x306 & ~x339 & ~x363 & ~x365 & ~x366 & ~x369 & ~x370 & ~x387 & ~x394 & ~x397 & ~x414 & ~x425 & ~x426 & ~x441 & ~x444 & ~x446 & ~x447 & ~x450 & ~x453 & ~x455 & ~x472 & ~x481 & ~x483 & ~x497 & ~x499 & ~x504 & ~x507 & ~x525 & ~x535 & ~x539 & ~x553 & ~x561 & ~x564 & ~x581 & ~x590 & ~x595 & ~x610 & ~x611 & ~x622 & ~x623 & ~x644 & ~x650 & ~x673 & ~x677 & ~x678 & ~x697 & ~x725 & ~x731 & ~x751 & ~x758 & ~x760 & ~x782;
assign c3495 =  x390;
assign c3497 =  x13 &  x40 &  x69 &  x94 &  x97 &  x126 &  x127 &  x152 &  x155 &  x181 &  x240 &  x296 &  x352 &  x488 &  x543 &  x683 & ~x2 & ~x3 & ~x21 & ~x36 & ~x48 & ~x54 & ~x57 & ~x61 & ~x80 & ~x85 & ~x86 & ~x87 & ~x115 & ~x117 & ~x134 & ~x138 & ~x142 & ~x195 & ~x310 & ~x332 & ~x363 & ~x364 & ~x368 & ~x423 & ~x445 & ~x446 & ~x505 & ~x555 & ~x564 & ~x592 & ~x623 & ~x647 & ~x666 & ~x668 & ~x673 & ~x677 & ~x692 & ~x721 & ~x732 & ~x762 & ~x781;
assign c3499 =  x355 &  x383 &  x460 &  x492 &  x512 &  x550 &  x551 &  x578 &  x607 &  x653 &  x655 &  x681 &  x718 &  x745 &  x747 &  x767 & ~x87 & ~x118 & ~x144 & ~x146 & ~x167 & ~x171 & ~x190 & ~x218 & ~x258 & ~x337 & ~x499 & ~x506 & ~x531 & ~x536 & ~x614 & ~x618 & ~x670 & ~x676 & ~x696 & ~x751;
assign c40 =  x368 &  x388 & ~x6 & ~x26 & ~x364;
assign c42 =  x262 &  x298 &  x327 &  x384 &  x412 &  x517 &  x654 & ~x1 & ~x7 & ~x8 & ~x9 & ~x59 & ~x82 & ~x86 & ~x116 & ~x117 & ~x139 & ~x140 & ~x169 & ~x173 & ~x219 & ~x223 & ~x225 & ~x247 & ~x277 & ~x279 & ~x283 & ~x304 & ~x307 & ~x309 & ~x310 & ~x421 & ~x532 & ~x644 & ~x649 & ~x672 & ~x675 & ~x676 & ~x704 & ~x721 & ~x723 & ~x729 & ~x730 & ~x733 & ~x758;
assign c44 =  x41 &  x71 & ~x6 & ~x7 & ~x8 & ~x9 & ~x23 & ~x24 & ~x25 & ~x26 & ~x27 & ~x29 & ~x31 & ~x50 & ~x51 & ~x53 & ~x56 & ~x57 & ~x58 & ~x59 & ~x81 & ~x84 & ~x108 & ~x137 & ~x139 & ~x140 & ~x141 & ~x142 & ~x143 & ~x165 & ~x166 & ~x169 & ~x171 & ~x193 & ~x195 & ~x221 & ~x223 & ~x225 & ~x226 & ~x227 & ~x249 & ~x250 & ~x254 & ~x277 & ~x279 & ~x280 & ~x282 & ~x306 & ~x307 & ~x309 & ~x310 & ~x333 & ~x336 & ~x390 & ~x392 & ~x419 & ~x422 & ~x449 & ~x474 & ~x476 & ~x477 & ~x503 & ~x505 & ~x506 & ~x531 & ~x532 & ~x558 & ~x561 & ~x615 & ~x617 & ~x642 & ~x670 & ~x672 & ~x681 & ~x682 & ~x691 & ~x699 & ~x701 & ~x713 & ~x716 & ~x717 & ~x718 & ~x744 & ~x745 & ~x754 & ~x757 & ~x764 & ~x765 & ~x771 & ~x774 & ~x776;
assign c46 =  x39 &  x185 &  x234 &  x299 &  x323 &  x345 &  x374 &  x482 &  x548 &  x607 &  x684 & ~x4 & ~x111 & ~x112 & ~x118 & ~x170 & ~x256 & ~x277 & ~x312 & ~x361 & ~x448 & ~x615 & ~x616 & ~x699;
assign c48 =  x243 &  x489 & ~x0 & ~x2 & ~x5 & ~x6 & ~x8 & ~x21 & ~x22 & ~x24 & ~x27 & ~x32 & ~x35 & ~x48 & ~x50 & ~x56 & ~x58 & ~x60 & ~x84 & ~x86 & ~x107 & ~x111 & ~x112 & ~x113 & ~x134 & ~x136 & ~x138 & ~x143 & ~x163 & ~x169 & ~x170 & ~x193 & ~x195 & ~x198 & ~x221 & ~x225 & ~x227 & ~x228 & ~x250 & ~x254 & ~x278 & ~x284 & ~x304 & ~x307 & ~x308 & ~x310 & ~x333 & ~x335 & ~x337 & ~x363 & ~x366 & ~x368 & ~x389 & ~x396 & ~x420 & ~x421 & ~x476 & ~x477 & ~x504 & ~x507 & ~x510 & ~x529 & ~x531 & ~x559 & ~x561 & ~x587 & ~x589 & ~x591 & ~x613 & ~x615 & ~x618 & ~x678 & ~x698 & ~x699 & ~x726 & ~x727 & ~x756 & ~x776 & ~x783;
assign c410 = ~x17 & ~x231 & ~x541;
assign c412 =  x41 &  x261 &  x743 & ~x0 & ~x3 & ~x4 & ~x30 & ~x32 & ~x47 & ~x54 & ~x76 & ~x83 & ~x90 & ~x106 & ~x107 & ~x110 & ~x111 & ~x133 & ~x143 & ~x144 & ~x163 & ~x165 & ~x172 & ~x190 & ~x191 & ~x198 & ~x221 & ~x223 & ~x225 & ~x226 & ~x255 & ~x257 & ~x279 & ~x285 & ~x305 & ~x332 & ~x337 & ~x364 & ~x417 & ~x446 & ~x506 & ~x534 & ~x589 & ~x616 & ~x645 & ~x651 & ~x677 & ~x679 & ~x693 & ~x703 & ~x726 & ~x758 & ~x782;
assign c414 =  x38 &  x158 &  x175 &  x187 &  x207 &  x230 &  x261 &  x292 &  x342 &  x369 &  x399 &  x548 &  x654 &  x711 & ~x2 & ~x3 & ~x23 & ~x30 & ~x62 & ~x193 & ~x253 & ~x310 & ~x422 & ~x448 & ~x586 & ~x643 & ~x644 & ~x729 & ~x754 & ~x756;
assign c416 = ~x7 & ~x10 & ~x17 & ~x24 & ~x26 & ~x27 & ~x47 & ~x48 & ~x50 & ~x51 & ~x54 & ~x59 & ~x84 & ~x85 & ~x90 & ~x109 & ~x110 & ~x116 & ~x118 & ~x144 & ~x194 & ~x220 & ~x224 & ~x252 & ~x255 & ~x278 & ~x283 & ~x333 & ~x335 & ~x361 & ~x364 & ~x417 & ~x548 & ~x590 & ~x726 & ~x764;
assign c418 =  x42 &  x443 &  x693 &  x696 & ~x28 & ~x32 & ~x52 & ~x53 & ~x88 & ~x115 & ~x224 & ~x249 & ~x254 & ~x420 & ~x447 & ~x503 & ~x671;
assign c420 = ~x0 & ~x4 & ~x8 & ~x9 & ~x20 & ~x23 & ~x30 & ~x35 & ~x36 & ~x47 & ~x48 & ~x52 & ~x57 & ~x61 & ~x86 & ~x115 & ~x118 & ~x163 & ~x167 & ~x170 & ~x194 & ~x195 & ~x196 & ~x226 & ~x248 & ~x254 & ~x278 & ~x281 & ~x291 & ~x301 & ~x335 & ~x419 & ~x446 & ~x478 & ~x586 & ~x730 & ~x757;
assign c422 =  x210 &  x230 &  x294 &  x378 &  x403 &  x436 &  x486 &  x526 &  x594 &  x704 &  x722 &  x751 & ~x2 & ~x6 & ~x22 & ~x51 & ~x135 & ~x165 & ~x166 & ~x195 & ~x334 & ~x338 & ~x559 & ~x730 & ~x741 & ~x771;
assign c424 =  x156 &  x356 &  x372 &  x384 &  x403 &  x441 &  x457 &  x546 &  x636 & ~x0 & ~x5 & ~x6 & ~x7 & ~x9 & ~x19 & ~x20 & ~x21 & ~x24 & ~x27 & ~x28 & ~x29 & ~x51 & ~x52 & ~x53 & ~x55 & ~x59 & ~x78 & ~x85 & ~x86 & ~x87 & ~x89 & ~x105 & ~x110 & ~x112 & ~x114 & ~x116 & ~x117 & ~x133 & ~x135 & ~x137 & ~x138 & ~x140 & ~x141 & ~x143 & ~x163 & ~x170 & ~x192 & ~x193 & ~x194 & ~x196 & ~x197 & ~x222 & ~x226 & ~x249 & ~x250 & ~x255 & ~x276 & ~x282 & ~x283 & ~x306 & ~x311 & ~x334 & ~x336 & ~x337 & ~x338 & ~x339 & ~x361 & ~x362 & ~x364 & ~x389 & ~x449 & ~x475 & ~x504 & ~x672 & ~x673 & ~x755 & ~x757 & ~x759;
assign c426 =  x44 &  x100 &  x152 &  x244 &  x261 &  x267 &  x291 &  x292 &  x315 &  x324 &  x356 &  x410 &  x411 &  x436 &  x441 &  x442 &  x463 &  x520 &  x596 &  x599 &  x604 &  x708 &  x709 &  x712 &  x719 & ~x2 & ~x23 & ~x28 & ~x33 & ~x57 & ~x80 & ~x135 & ~x140 & ~x165 & ~x169 & ~x192 & ~x193 & ~x224 & ~x226 & ~x277 & ~x305 & ~x306 & ~x307 & ~x309 & ~x334 & ~x336 & ~x420 & ~x532 & ~x535 & ~x557 & ~x587 & ~x588 & ~x754 & ~x758 & ~x783;
assign c428 = ~x1 & ~x9 & ~x19 & ~x23 & ~x32 & ~x59 & ~x61 & ~x81 & ~x116 & ~x140 & ~x169 & ~x251 & ~x269 & ~x277 & ~x282 & ~x307 & ~x389 & ~x420 & ~x478 & ~x728 & ~x737 & ~x738 & ~x740;
assign c430 =  x372 & ~x8 & ~x21 & ~x22 & ~x23 & ~x59 & ~x67 & ~x77 & ~x78 & ~x79 & ~x116 & ~x140 & ~x167 & ~x220 & ~x221 & ~x223 & ~x225 & ~x248 & ~x252 & ~x277 & ~x278 & ~x337 & ~x362 & ~x389 & ~x391 & ~x445 & ~x475 & ~x502 & ~x505 & ~x506 & ~x530 & ~x534 & ~x560 & ~x561 & ~x586 & ~x645 & ~x728;
assign c432 =  x378 &  x430 &  x441 &  x483 &  x708 &  x742 &  x767 & ~x278 & ~x360;
assign c434 =  x171;
assign c436 =  x125 &  x235 &  x239 &  x260 &  x265 &  x266 &  x273 &  x275 &  x348 &  x378 &  x442 &  x443 &  x527 &  x539 &  x565 &  x568 &  x639 &  x668 & ~x53 & ~x54 & ~x56 & ~x80 & ~x110 & ~x114 & ~x278 & ~x476 & ~x783;
assign c438 =  x608 & ~x5 & ~x8 & ~x19 & ~x25 & ~x26 & ~x54 & ~x84 & ~x136 & ~x144 & ~x171 & ~x193 & ~x221 & ~x253 & ~x254 & ~x255 & ~x276 & ~x310 & ~x392 & ~x505 & ~x530 & ~x560 & ~x644 & ~x684 & ~x698 & ~x702 & ~x756 & ~x757;
assign c440 =  x125 &  x203 &  x316 &  x317 &  x371 &  x540 &  x571 &  x572 & ~x5 & ~x6 & ~x30 & ~x53 & ~x56 & ~x57 & ~x58 & ~x61 & ~x62 & ~x86 & ~x90 & ~x109 & ~x111 & ~x113 & ~x115 & ~x118 & ~x135 & ~x138 & ~x141 & ~x162 & ~x172 & ~x194 & ~x225 & ~x226 & ~x227 & ~x253 & ~x254 & ~x276 & ~x279 & ~x281 & ~x310 & ~x333 & ~x367 & ~x394 & ~x395 & ~x419 & ~x422 & ~x446 & ~x448 & ~x474 & ~x501 & ~x507 & ~x531 & ~x590 & ~x616 & ~x644 & ~x698 & ~x699 & ~x702 & ~x728 & ~x755 & ~x756 & ~x758;
assign c442 =  x261 &  x265 &  x267 &  x271 &  x295 &  x320 &  x352 &  x433 &  x491 &  x494 &  x516 &  x547 &  x598 &  x599 &  x629 &  x633 &  x662 &  x682 &  x687 &  x711 & ~x0 & ~x1 & ~x4 & ~x5 & ~x9 & ~x18 & ~x22 & ~x23 & ~x29 & ~x31 & ~x35 & ~x36 & ~x47 & ~x49 & ~x52 & ~x59 & ~x62 & ~x78 & ~x80 & ~x88 & ~x91 & ~x106 & ~x107 & ~x111 & ~x113 & ~x118 & ~x139 & ~x166 & ~x172 & ~x194 & ~x196 & ~x247 & ~x253 & ~x254 & ~x281 & ~x282 & ~x333 & ~x445 & ~x446 & ~x473 & ~x503 & ~x506 & ~x530 & ~x561 & ~x586 & ~x671 & ~x756 & ~x762 & ~x763 & ~x781 & ~x782;
assign c444 =  x345 &  x405 &  x429 & ~x0 & ~x7 & ~x8 & ~x51 & ~x60 & ~x139 & ~x140 & ~x220 & ~x221 & ~x425 & ~x450 & ~x736;
assign c446 =  x259 &  x261 &  x266 &  x299 &  x329 &  x356 &  x375 &  x377 &  x462 &  x493 &  x514 &  x659 &  x662 &  x687 & ~x17 & ~x18 & ~x29 & ~x50 & ~x51 & ~x52 & ~x53 & ~x56 & ~x83 & ~x87 & ~x137 & ~x138 & ~x167 & ~x168 & ~x173 & ~x194 & ~x201 & ~x226 & ~x248 & ~x250 & ~x251 & ~x280 & ~x307 & ~x309 & ~x332 & ~x339 & ~x363 & ~x365 & ~x420 & ~x447 & ~x532 & ~x588 & ~x756 & ~x763 & ~x782;
assign c448 =  x313 &  x623 & ~x49 & ~x56 & ~x80 & ~x227 & ~x334 & ~x335 & ~x362 & ~x534;
assign c450 =  x230 &  x368 &  x452 &  x508 &  x731 & ~x55;
assign c452 =  x602 & ~x20 & ~x35 & ~x48 & ~x78 & ~x137 & ~x164 & ~x193 & ~x336 & ~x432 & ~x476 & ~x699 & ~x702;
assign c454 = ~x0 & ~x1 & ~x2 & ~x4 & ~x6 & ~x7 & ~x8 & ~x10 & ~x17 & ~x20 & ~x21 & ~x22 & ~x23 & ~x25 & ~x27 & ~x28 & ~x29 & ~x30 & ~x31 & ~x34 & ~x35 & ~x36 & ~x48 & ~x50 & ~x53 & ~x54 & ~x55 & ~x56 & ~x57 & ~x59 & ~x61 & ~x78 & ~x79 & ~x80 & ~x81 & ~x82 & ~x83 & ~x85 & ~x87 & ~x88 & ~x89 & ~x90 & ~x107 & ~x108 & ~x110 & ~x112 & ~x116 & ~x136 & ~x140 & ~x143 & ~x144 & ~x164 & ~x167 & ~x168 & ~x169 & ~x172 & ~x190 & ~x193 & ~x195 & ~x197 & ~x198 & ~x222 & ~x223 & ~x225 & ~x226 & ~x227 & ~x248 & ~x250 & ~x251 & ~x254 & ~x277 & ~x278 & ~x280 & ~x281 & ~x283 & ~x304 & ~x305 & ~x306 & ~x307 & ~x308 & ~x310 & ~x331 & ~x333 & ~x334 & ~x335 & ~x336 & ~x337 & ~x338 & ~x361 & ~x362 & ~x363 & ~x364 & ~x365 & ~x366 & ~x367 & ~x389 & ~x390 & ~x391 & ~x392 & ~x393 & ~x394 & ~x417 & ~x418 & ~x423 & ~x444 & ~x445 & ~x446 & ~x447 & ~x448 & ~x450 & ~x451 & ~x473 & ~x475 & ~x477 & ~x500 & ~x501 & ~x502 & ~x506 & ~x507 & ~x532 & ~x535 & ~x558 & ~x560 & ~x561 & ~x585 & ~x586 & ~x613 & ~x616 & ~x643 & ~x644 & ~x646 & ~x670 & ~x671 & ~x673 & ~x675 & ~x698 & ~x699 & ~x702 & ~x725 & ~x726 & ~x727 & ~x728 & ~x729 & ~x731 & ~x736 & ~x747 & ~x755 & ~x756 & ~x759 & ~x765 & ~x772 & ~x775 & ~x776 & ~x781 & ~x783;
assign c456 =  x13 &  x94 &  x121 &  x233 &  x402 &  x463 &  x488 &  x494 & ~x6 & ~x9 & ~x20 & ~x32 & ~x59 & ~x60 & ~x79 & ~x80 & ~x86 & ~x116 & ~x138 & ~x194 & ~x195 & ~x219 & ~x247 & ~x250 & ~x254 & ~x255 & ~x278 & ~x284 & ~x306 & ~x361 & ~x362 & ~x364 & ~x388 & ~x393 & ~x416 & ~x502 & ~x531 & ~x558 & ~x586 & ~x615 & ~x670 & ~x734 & ~x735 & ~x749 & ~x763 & ~x777 & ~x778;
assign c458 =  x39 &  x179 &  x209 &  x210 &  x266 &  x324 &  x357 &  x461 &  x491 &  x566 &  x601 &  x659 &  x712 &  x737 &  x739 & ~x22 & ~x29 & ~x50 & ~x256 & ~x304 & ~x393 & ~x423 & ~x501 & ~x558 & ~x559 & ~x563 & ~x591 & ~x646 & ~x754;
assign c460 =  x245 &  x260 &  x316 &  x351 &  x426 &  x431 &  x554 &  x573 &  x639 &  x693 &  x707 & ~x6 & ~x52 & ~x55 & ~x112 & ~x226 & ~x256 & ~x304 & ~x393 & ~x394 & ~x473 & ~x559 & ~x591 & ~x670 & ~x697;
assign c462 =  x150 &  x178 &  x180 &  x202 &  x208 &  x233 &  x237 &  x261 &  x286 &  x297 &  x302 &  x314 &  x319 &  x325 &  x349 &  x384 &  x386 &  x414 &  x487 &  x554 &  x582 &  x592 &  x654 &  x684 &  x691 &  x732 & ~x55 & ~x62 & ~x79 & ~x107 & ~x112 & ~x165 & ~x168 & ~x475 & ~x671 & ~x757;
assign c464 =  x670;
assign c466 =  x232 &  x239 &  x288 &  x293 &  x356 &  x399 &  x524 &  x581 &  x713 & ~x1 & ~x7 & ~x9 & ~x18 & ~x25 & ~x79 & ~x110 & ~x118 & ~x135 & ~x136 & ~x141 & ~x163 & ~x191 & ~x198 & ~x199 & ~x220 & ~x223 & ~x225 & ~x228 & ~x247 & ~x333 & ~x339 & ~x391 & ~x478 & ~x505 & ~x559 & ~x585 & ~x614 & ~x675 & ~x725 & ~x782 & ~x783;
assign c468 =  x259 &  x511 &  x580 & ~x370;
assign c470 = ~x10 & ~x11 & ~x51 & ~x77 & ~x92 & ~x145 & ~x147 & ~x360 & ~x388 & ~x391 & ~x393 & ~x444 & ~x508 & ~x694 & ~x708 & ~x728;
assign c472 =  x39 &  x566 &  x747 & ~x60 & ~x61 & ~x85 & ~x170 & ~x194 & ~x283 & ~x284 & ~x312 & ~x363 & ~x367 & ~x423 & ~x478 & ~x535 & ~x644 & ~x702 & ~x781;
assign c474 = ~x222 & ~x241 & ~x272 & ~x318;
assign c476 =  x506;
assign c478 =  x331 & ~x3 & ~x32 & ~x49 & ~x52 & ~x58 & ~x60 & ~x85 & ~x166 & ~x195 & ~x197 & ~x225 & ~x249 & ~x448 & ~x504 & ~x560 & ~x587 & ~x617 & ~x715 & ~x743 & ~x747;
assign c480 =  x375 &  x387 &  x413 & ~x0 & ~x10 & ~x19 & ~x26 & ~x30 & ~x34 & ~x52 & ~x254 & ~x309 & ~x363 & ~x450 & ~x530 & ~x533 & ~x585 & ~x617 & ~x669 & ~x743 & ~x753;
assign c482 =  x715 & ~x0 & ~x7 & ~x10 & ~x18 & ~x23 & ~x28 & ~x29 & ~x30 & ~x31 & ~x35 & ~x36 & ~x50 & ~x56 & ~x61 & ~x63 & ~x77 & ~x78 & ~x84 & ~x86 & ~x88 & ~x92 & ~x116 & ~x133 & ~x138 & ~x139 & ~x140 & ~x141 & ~x162 & ~x163 & ~x169 & ~x171 & ~x172 & ~x174 & ~x190 & ~x192 & ~x193 & ~x194 & ~x197 & ~x223 & ~x225 & ~x226 & ~x227 & ~x246 & ~x248 & ~x252 & ~x257 & ~x276 & ~x277 & ~x282 & ~x283 & ~x285 & ~x306 & ~x308 & ~x312 & ~x331 & ~x338 & ~x340 & ~x361 & ~x364 & ~x368 & ~x388 & ~x419 & ~x423 & ~x446 & ~x452 & ~x474 & ~x501 & ~x530 & ~x562 & ~x563 & ~x587 & ~x613 & ~x618 & ~x619 & ~x642 & ~x644 & ~x672 & ~x698 & ~x699 & ~x700 & ~x702 & ~x731 & ~x754 & ~x775 & ~x780;
assign c484 =  x602 & ~x20 & ~x78 & ~x79 & ~x87 & ~x116 & ~x137 & ~x250 & ~x364 & ~x379 & ~x764;
assign c486 =  x291 &  x294 &  x328 &  x427 &  x431 &  x538 &  x541 &  x543 &  x572 &  x579 &  x651 &  x656 &  x690 &  x743 & ~x1 & ~x24 & ~x32 & ~x78 & ~x82 & ~x83 & ~x110 & ~x111 & ~x166 & ~x167 & ~x170 & ~x197 & ~x222 & ~x334 & ~x336 & ~x339 & ~x365 & ~x418 & ~x420 & ~x421 & ~x447 & ~x503 & ~x504 & ~x725 & ~x754 & ~x781;
assign c488 =  x71 &  x731 & ~x29 & ~x50 & ~x51 & ~x165 & ~x168 & ~x280;
assign c490 =  x523 & ~x9 & ~x10 & ~x28 & ~x51 & ~x110 & ~x137 & ~x146 & ~x162 & ~x166 & ~x191 & ~x198 & ~x247 & ~x277 & ~x283 & ~x337 & ~x340 & ~x361 & ~x422 & ~x507 & ~x557 & ~x559 & ~x560 & ~x619 & ~x646 & ~x700 & ~x736 & ~x754 & ~x768 & ~x775 & ~x780;
assign c492 =  x14 &  x156 &  x240 &  x270 &  x320 &  x356 &  x460 &  x603 &  x740 & ~x4 & ~x83 & ~x137 & ~x144 & ~x166 & ~x190 & ~x191 & ~x196 & ~x218 & ~x227 & ~x281 & ~x335 & ~x362 & ~x363 & ~x533 & ~x642 & ~x755 & ~x763;
assign c494 =  x238 &  x262 &  x265 &  x295 &  x372 &  x469 &  x497 &  x516 &  x543 &  x545 &  x568 &  x579 &  x598 &  x681 & ~x3 & ~x8 & ~x19 & ~x27 & ~x50 & ~x56 & ~x59 & ~x112 & ~x164 & ~x166 & ~x168 & ~x169 & ~x171 & ~x190 & ~x223 & ~x224 & ~x251 & ~x255 & ~x256 & ~x281 & ~x308 & ~x309 & ~x311 & ~x335 & ~x336 & ~x339 & ~x340 & ~x360 & ~x364 & ~x367 & ~x389 & ~x390 & ~x393 & ~x395 & ~x419 & ~x450 & ~x474 & ~x477 & ~x478 & ~x502 & ~x504 & ~x505 & ~x532 & ~x560 & ~x561 & ~x613 & ~x615 & ~x616 & ~x671 & ~x673 & ~x727 & ~x730 & ~x755 & ~x756 & ~x757 & ~x758;
assign c496 =  x98 &  x484 &  x553 &  x567 &  x745 & ~x1 & ~x5 & ~x18 & ~x20 & ~x25 & ~x26 & ~x28 & ~x47 & ~x49 & ~x50 & ~x51 & ~x53 & ~x76 & ~x77 & ~x78 & ~x79 & ~x82 & ~x88 & ~x107 & ~x108 & ~x110 & ~x114 & ~x140 & ~x164 & ~x165 & ~x166 & ~x193 & ~x196 & ~x197 & ~x225 & ~x251 & ~x255 & ~x277 & ~x278 & ~x307 & ~x310 & ~x364 & ~x420 & ~x421 & ~x445 & ~x447 & ~x450 & ~x477 & ~x478 & ~x504 & ~x505 & ~x532 & ~x533 & ~x587 & ~x588 & ~x590 & ~x617 & ~x645 & ~x646 & ~x701 & ~x702 & ~x726 & ~x757 & ~x781;
assign c498 =  x372 & ~x0 & ~x8 & ~x9 & ~x10 & ~x21 & ~x54 & ~x60 & ~x62 & ~x77 & ~x85 & ~x111 & ~x140 & ~x162 & ~x164 & ~x171 & ~x199 & ~x225 & ~x251 & ~x276 & ~x278 & ~x304 & ~x305 & ~x306 & ~x308 & ~x331 & ~x334 & ~x393 & ~x448 & ~x501 & ~x527 & ~x531 & ~x563 & ~x564 & ~x615 & ~x667 & ~x674 & ~x678 & ~x697 & ~x698 & ~x701 & ~x757 & ~x764 & ~x774;
assign c4100 =  x238 &  x378 &  x433 &  x568 &  x582 &  x596 &  x662 &  x683 &  x709 &  x737 & ~x5 & ~x21 & ~x51 & ~x56 & ~x85 & ~x110 & ~x138 & ~x224 & ~x275 & ~x360 & ~x363 & ~x475 & ~x477 & ~x500 & ~x503 & ~x528 & ~x585 & ~x614 & ~x645 & ~x671 & ~x759;
assign c4102 =  x533;
assign c4104 = ~x2 & ~x3 & ~x8 & ~x20 & ~x48 & ~x54 & ~x55 & ~x59 & ~x78 & ~x81 & ~x85 & ~x109 & ~x112 & ~x135 & ~x140 & ~x169 & ~x171 & ~x196 & ~x200 & ~x225 & ~x248 & ~x249 & ~x252 & ~x253 & ~x254 & ~x255 & ~x276 & ~x282 & ~x305 & ~x306 & ~x307 & ~x310 & ~x333 & ~x334 & ~x336 & ~x338 & ~x363 & ~x364 & ~x365 & ~x380 & ~x391 & ~x392 & ~x394 & ~x419 & ~x420 & ~x421 & ~x474 & ~x476 & ~x505 & ~x506 & ~x534 & ~x558 & ~x559 & ~x562 & ~x587 & ~x616 & ~x645 & ~x646 & ~x699 & ~x701 & ~x755 & ~x757 & ~x782 & ~x783;
assign c4106 = ~x3 & ~x5 & ~x6 & ~x7 & ~x22 & ~x25 & ~x26 & ~x27 & ~x28 & ~x31 & ~x34 & ~x49 & ~x56 & ~x57 & ~x61 & ~x78 & ~x79 & ~x80 & ~x83 & ~x88 & ~x106 & ~x109 & ~x111 & ~x115 & ~x116 & ~x137 & ~x166 & ~x194 & ~x196 & ~x199 & ~x221 & ~x222 & ~x223 & ~x249 & ~x250 & ~x254 & ~x255 & ~x277 & ~x278 & ~x279 & ~x280 & ~x282 & ~x307 & ~x334 & ~x337 & ~x348 & ~x361 & ~x366 & ~x382 & ~x390 & ~x392 & ~x418 & ~x421 & ~x450 & ~x474 & ~x477 & ~x505 & ~x532 & ~x561 & ~x587 & ~x671 & ~x672 & ~x673 & ~x699 & ~x702 & ~x729 & ~x755 & ~x781;
assign c4108 =  x100 &  x523 &  x695 &  x706 &  x721 &  x752 & ~x26 & ~x165;
assign c4110 =  x357 &  x455 &  x483 &  x553 &  x609 & ~x0 & ~x2 & ~x6 & ~x33 & ~x59 & ~x84 & ~x86 & ~x107 & ~x115 & ~x141 & ~x169 & ~x222 & ~x226 & ~x254 & ~x338 & ~x363 & ~x392 & ~x446 & ~x534 & ~x558 & ~x645 & ~x734 & ~x750 & ~x753 & ~x755 & ~x781;
assign c4112 =  x184 &  x316 &  x408 &  x424 &  x452 &  x536 &  x545 &  x648 &  x704 & ~x1 & ~x2 & ~x28 & ~x32 & ~x48 & ~x55 & ~x61 & ~x78 & ~x87 & ~x165 & ~x171 & ~x194 & ~x280 & ~x310 & ~x333 & ~x394 & ~x477 & ~x529 & ~x617 & ~x642 & ~x644 & ~x754 & ~x771 & ~x781;
assign c4114 =  x204 &  x211 &  x234 &  x240 &  x242 &  x261 &  x270 &  x293 &  x299 &  x344 &  x384 &  x434 &  x435 &  x462 &  x464 &  x548 & ~x1 & ~x4 & ~x5 & ~x7 & ~x20 & ~x23 & ~x25 & ~x28 & ~x32 & ~x33 & ~x59 & ~x78 & ~x83 & ~x87 & ~x112 & ~x113 & ~x114 & ~x116 & ~x163 & ~x166 & ~x172 & ~x191 & ~x196 & ~x198 & ~x220 & ~x223 & ~x226 & ~x256 & ~x275 & ~x281 & ~x282 & ~x283 & ~x305 & ~x310 & ~x335 & ~x336 & ~x361 & ~x363 & ~x390 & ~x395 & ~x421 & ~x445 & ~x446 & ~x447 & ~x476 & ~x501 & ~x502 & ~x503 & ~x506 & ~x529 & ~x532 & ~x533 & ~x534 & ~x535 & ~x563 & ~x584 & ~x588 & ~x590 & ~x613 & ~x615 & ~x616 & ~x618 & ~x644 & ~x648 & ~x669 & ~x671 & ~x696 & ~x700 & ~x705 & ~x706 & ~x751 & ~x755 & ~x757 & ~x776 & ~x781;
assign c4116 =  x38 &  x39 &  x41 &  x43 &  x120 &  x291 &  x319 &  x321 &  x347 &  x352 &  x355 &  x403 &  x426 &  x495 &  x523 &  x545 &  x575 &  x578 &  x684 &  x746 & ~x51 & ~x53 & ~x85 & ~x108 & ~x111 & ~x135 & ~x167 & ~x168 & ~x196 & ~x198 & ~x223 & ~x228 & ~x283 & ~x304 & ~x311 & ~x333 & ~x336 & ~x447 & ~x450 & ~x533 & ~x700 & ~x728 & ~x758;
assign c4118 =  x40 &  x42 &  x152 &  x207 &  x233 &  x296 &  x321 &  x323 &  x354 &  x372 &  x379 &  x382 &  x439 &  x461 &  x488 &  x514 &  x515 &  x576 & ~x5 & ~x21 & ~x30 & ~x53 & ~x54 & ~x60 & ~x85 & ~x113 & ~x119 & ~x137 & ~x138 & ~x140 & ~x199 & ~x220 & ~x282 & ~x284 & ~x333 & ~x334 & ~x338 & ~x364 & ~x389 & ~x391 & ~x420 & ~x446 & ~x448 & ~x450 & ~x474 & ~x476 & ~x503 & ~x585 & ~x587 & ~x614 & ~x615 & ~x642 & ~x644 & ~x645 & ~x700 & ~x757;
assign c4120 =  x121 &  x129 &  x205 &  x329 &  x457 &  x592 &  x647 & ~x30 & ~x49 & ~x140 & ~x503;
assign c4122 = ~x0 & ~x10 & ~x25 & ~x34 & ~x46 & ~x56 & ~x117 & ~x136 & ~x141 & ~x166 & ~x195 & ~x198 & ~x200 & ~x201 & ~x228 & ~x255 & ~x256 & ~x285 & ~x332 & ~x334 & ~x390 & ~x450 & ~x501 & ~x535 & ~x585 & ~x624 & ~x666 & ~x668 & ~x693 & ~x706 & ~x734 & ~x750 & ~x756 & ~x757 & ~x759 & ~x764 & ~x783;
assign c4124 =  x42 &  x317 &  x411 &  x434 & ~x10 & ~x18 & ~x49 & ~x117 & ~x141 & ~x145 & ~x168 & ~x192 & ~x193 & ~x222 & ~x226 & ~x248 & ~x251 & ~x304 & ~x309 & ~x310 & ~x333 & ~x421 & ~x531 & ~x585 & ~x590 & ~x616 & ~x678 & ~x775;
assign c4126 =  x261 &  x289 &  x327 & ~x253 & ~x418 & ~x622 & ~x652 & ~x764 & ~x775;
assign c4128 =  x289 & ~x10 & ~x56 & ~x61 & ~x75 & ~x118 & ~x135 & ~x147 & ~x173 & ~x174 & ~x190 & ~x195 & ~x249 & ~x253 & ~x257 & ~x313 & ~x333 & ~x365 & ~x388 & ~x396 & ~x450 & ~x451 & ~x475 & ~x501 & ~x504 & ~x587 & ~x615 & ~x782 & ~x783;
assign c4130 =  x258 &  x300 &  x313 &  x340 &  x350 &  x377 &  x519 &  x526 &  x547 & ~x20 & ~x25 & ~x28 & ~x35 & ~x61 & ~x77 & ~x169 & ~x252 & ~x308 & ~x337 & ~x363 & ~x390 & ~x532 & ~x588 & ~x642 & ~x643 & ~x726 & ~x763 & ~x769;
assign c4132 =  x270 &  x516 &  x546 & ~x2 & ~x4 & ~x5 & ~x21 & ~x27 & ~x55 & ~x82 & ~x140 & ~x226 & ~x229 & ~x248 & ~x249 & ~x275 & ~x279 & ~x283 & ~x304 & ~x359 & ~x390 & ~x392 & ~x419 & ~x589 & ~x616 & ~x620 & ~x621 & ~x666 & ~x674 & ~x678 & ~x679 & ~x696 & ~x703 & ~x726 & ~x729 & ~x732 & ~x775 & ~x780;
assign c4134 =  x285 &  x287 &  x374 &  x380 &  x397 &  x410 &  x431 &  x465 &  x466 &  x485 &  x494 &  x513 &  x542 & ~x5 & ~x7 & ~x24 & ~x26 & ~x33 & ~x61 & ~x84 & ~x85 & ~x87 & ~x88 & ~x106 & ~x144 & ~x167 & ~x195 & ~x199 & ~x250 & ~x310 & ~x334 & ~x338 & ~x363 & ~x394 & ~x506 & ~x530 & ~x532 & ~x561 & ~x562 & ~x585 & ~x613 & ~x645 & ~x669 & ~x674 & ~x698 & ~x726 & ~x746 & ~x765 & ~x782;
assign c4136 = ~x50 & ~x208 & ~x241 & ~x290 & ~x446 & ~x770;
assign c4138 =  x312 & ~x721 & ~x742;
assign c4140 =  x117 &  x567;
assign c4142 =  x286 &  x302 &  x325 &  x374 &  x380 &  x481 &  x733 &  x751 & ~x4 & ~x20 & ~x21 & ~x30 & ~x63 & ~x76 & ~x77 & ~x106 & ~x141 & ~x222 & ~x225 & ~x254 & ~x278 & ~x365 & ~x390 & ~x420 & ~x421 & ~x447 & ~x534 & ~x587 & ~x615 & ~x642 & ~x644 & ~x699 & ~x772;
assign c4144 =  x125 & ~x3 & ~x7 & ~x22 & ~x24 & ~x30 & ~x33 & ~x35 & ~x48 & ~x51 & ~x54 & ~x56 & ~x58 & ~x63 & ~x78 & ~x79 & ~x105 & ~x110 & ~x115 & ~x134 & ~x136 & ~x140 & ~x143 & ~x144 & ~x163 & ~x191 & ~x193 & ~x194 & ~x199 & ~x219 & ~x220 & ~x223 & ~x249 & ~x251 & ~x256 & ~x284 & ~x304 & ~x305 & ~x309 & ~x310 & ~x360 & ~x363 & ~x365 & ~x388 & ~x389 & ~x393 & ~x418 & ~x419 & ~x446 & ~x448 & ~x475 & ~x531 & ~x560 & ~x588 & ~x644 & ~x646 & ~x670 & ~x675 & ~x678 & ~x699 & ~x726 & ~x727 & ~x756 & ~x764 & ~x773 & ~x774;
assign c4146 = ~x231 & ~x362 & ~x363 & ~x375 & ~x505;
assign c4148 =  x206 &  x207 &  x243 &  x270 &  x271 &  x345 &  x377 &  x381 &  x438 &  x461 &  x630 &  x654 &  x683 & ~x4 & ~x28 & ~x30 & ~x50 & ~x55 & ~x79 & ~x82 & ~x115 & ~x141 & ~x163 & ~x165 & ~x167 & ~x226 & ~x228 & ~x255 & ~x280 & ~x284 & ~x309 & ~x365 & ~x389 & ~x390 & ~x445 & ~x530 & ~x560 & ~x618 & ~x646 & ~x674 & ~x675 & ~x697 & ~x725 & ~x734 & ~x780;
assign c4150 =  x345 & ~x7 & ~x561 & ~x653 & ~x716;
assign c4152 = ~x17 & ~x33 & ~x47 & ~x49 & ~x78 & ~x109 & ~x114 & ~x118 & ~x133 & ~x169 & ~x196 & ~x200 & ~x220 & ~x225 & ~x226 & ~x280 & ~x376 & ~x389 & ~x390 & ~x473 & ~x500 & ~x504 & ~x506 & ~x532 & ~x669;
assign c4154 =  x13 &  x210 &  x303 &  x331 &  x342 &  x343 &  x432 &  x676 & ~x22 & ~x86 & ~x108 & ~x112 & ~x139 & ~x475 & ~x756;
assign c4156 =  x72 &  x357 &  x406 &  x427 &  x563 &  x619 & ~x1 & ~x26 & ~x33;
assign c4158 =  x43 &  x70 &  x98 &  x315 &  x343 &  x356 &  x413 &  x441 &  x593 &  x694 & ~x3 & ~x5 & ~x6 & ~x7 & ~x8 & ~x17 & ~x18 & ~x19 & ~x20 & ~x21 & ~x23 & ~x25 & ~x27 & ~x28 & ~x31 & ~x33 & ~x34 & ~x35 & ~x47 & ~x48 & ~x49 & ~x50 & ~x51 & ~x54 & ~x55 & ~x57 & ~x60 & ~x62 & ~x63 & ~x76 & ~x78 & ~x79 & ~x81 & ~x83 & ~x84 & ~x86 & ~x89 & ~x106 & ~x109 & ~x113 & ~x115 & ~x135 & ~x137 & ~x138 & ~x139 & ~x140 & ~x141 & ~x143 & ~x144 & ~x168 & ~x169 & ~x170 & ~x192 & ~x193 & ~x195 & ~x197 & ~x198 & ~x199 & ~x223 & ~x224 & ~x226 & ~x227 & ~x249 & ~x251 & ~x252 & ~x253 & ~x279 & ~x280 & ~x281 & ~x282 & ~x283 & ~x304 & ~x305 & ~x306 & ~x307 & ~x309 & ~x332 & ~x333 & ~x335 & ~x337 & ~x338 & ~x361 & ~x363 & ~x365 & ~x391 & ~x392 & ~x393 & ~x419 & ~x421 & ~x422 & ~x446 & ~x447 & ~x450 & ~x473 & ~x474 & ~x475 & ~x476 & ~x501 & ~x502 & ~x504 & ~x505 & ~x532 & ~x557 & ~x560 & ~x561 & ~x562 & ~x586 & ~x588 & ~x590 & ~x614 & ~x615 & ~x617 & ~x641 & ~x643 & ~x644 & ~x645 & ~x671 & ~x672 & ~x698 & ~x699 & ~x700 & ~x701 & ~x726 & ~x728 & ~x729 & ~x730 & ~x755 & ~x756 & ~x757 & ~x765 & ~x767 & ~x769 & ~x770 & ~x772 & ~x773 & ~x774 & ~x775 & ~x776 & ~x781 & ~x782;
assign c4160 =  x329 &  x428 &  x459 &  x490 &  x554 &  x566 &  x573 &  x623 &  x628 &  x653 &  x683 &  x690 &  x743 &  x745 & ~x27 & ~x54 & ~x55 & ~x59 & ~x89 & ~x168 & ~x171 & ~x192 & ~x249 & ~x307 & ~x334 & ~x419 & ~x504 & ~x647 & ~x699 & ~x729;
assign c4162 =  x294 &  x434 &  x462 &  x574 &  x602 & ~x4 & ~x19 & ~x23 & ~x24 & ~x36 & ~x56 & ~x57 & ~x59 & ~x61 & ~x80 & ~x83 & ~x107 & ~x108 & ~x148 & ~x192 & ~x219 & ~x223 & ~x227 & ~x248 & ~x251 & ~x252 & ~x277 & ~x279 & ~x282 & ~x304 & ~x305 & ~x307 & ~x308 & ~x362 & ~x364 & ~x367 & ~x389 & ~x392 & ~x417 & ~x473 & ~x474 & ~x475 & ~x478 & ~x502 & ~x533 & ~x534 & ~x558 & ~x588 & ~x589 & ~x615 & ~x616 & ~x617 & ~x645 & ~x673 & ~x700 & ~x701 & ~x728 & ~x759;
assign c4164 =  x176 &  x185 &  x236 &  x262 &  x267 &  x275 &  x567 &  x592 & ~x165;
assign c4166 =  x45 &  x100 &  x268 &  x483 &  x540 &  x599 &  x653 &  x691 &  x715 & ~x48 & ~x62 & ~x82 & ~x86 & ~x89 & ~x135 & ~x279 & ~x310 & ~x334 & ~x338 & ~x447 & ~x479 & ~x535 & ~x589 & ~x617 & ~x675 & ~x777 & ~x783;
assign c4168 =  x236 &  x241 &  x261 &  x294 &  x459 &  x517 &  x547 &  x603 &  x631 &  x657 &  x659 &  x660 & ~x3 & ~x7 & ~x8 & ~x17 & ~x26 & ~x58 & ~x111 & ~x118 & ~x132 & ~x136 & ~x139 & ~x169 & ~x250 & ~x252 & ~x253 & ~x277 & ~x280 & ~x332 & ~x338 & ~x394 & ~x417 & ~x447 & ~x590 & ~x614 & ~x615 & ~x645 & ~x673;
assign c4170 = ~x2 & ~x18 & ~x19 & ~x49 & ~x50 & ~x53 & ~x61 & ~x84 & ~x87 & ~x115 & ~x139 & ~x141 & ~x166 & ~x170 & ~x193 & ~x198 & ~x230 & ~x258 & ~x283 & ~x308 & ~x333 & ~x358 & ~x419 & ~x477 & ~x529 & ~x531 & ~x534 & ~x557 & ~x558 & ~x559 & ~x560 & ~x674 & ~x697 & ~x729 & ~x737 & ~x768 & ~x774;
assign c4172 =  x585;
assign c4174 =  x751 &  x760 & ~x62 & ~x85 & ~x309 & ~x334 & ~x504 & ~x642;
assign c4176 =  x40 &  x41 &  x211 &  x269 &  x293 &  x320 &  x327 &  x344 &  x351 &  x403 &  x405 &  x433 &  x459 &  x460 &  x491 &  x493 &  x514 &  x516 &  x521 &  x570 &  x571 &  x629 &  x632 &  x654 &  x656 &  x682 &  x687 &  x688 & ~x3 & ~x6 & ~x9 & ~x10 & ~x25 & ~x31 & ~x54 & ~x55 & ~x61 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x108 & ~x110 & ~x117 & ~x136 & ~x138 & ~x140 & ~x143 & ~x144 & ~x163 & ~x164 & ~x190 & ~x197 & ~x218 & ~x219 & ~x224 & ~x225 & ~x226 & ~x249 & ~x255 & ~x256 & ~x277 & ~x283 & ~x305 & ~x308 & ~x310 & ~x334 & ~x363 & ~x364 & ~x365 & ~x368 & ~x390 & ~x392 & ~x395 & ~x396 & ~x420 & ~x444 & ~x476 & ~x501 & ~x503 & ~x504 & ~x508 & ~x531 & ~x533 & ~x561 & ~x611 & ~x615 & ~x619 & ~x641 & ~x643 & ~x645 & ~x646 & ~x670 & ~x671 & ~x672 & ~x702 & ~x726 & ~x757 & ~x776 & ~x783;
assign c4178 =  x100 &  x124 &  x153 &  x156 &  x158 &  x181 &  x184 &  x217 &  x230 &  x237 &  x259 &  x290 &  x291 &  x296 &  x315 &  x317 &  x321 &  x327 &  x342 &  x346 &  x351 &  x353 &  x371 &  x399 &  x425 &  x427 &  x434 &  x437 &  x461 &  x487 &  x497 &  x498 &  x512 &  x517 &  x547 &  x568 &  x570 &  x571 &  x578 &  x593 &  x605 &  x610 &  x666 &  x676 &  x693 &  x705 & ~x1 & ~x2 & ~x29 & ~x32 & ~x79 & ~x81 & ~x82 & ~x85 & ~x87 & ~x107 & ~x115 & ~x140 & ~x165 & ~x166 & ~x194 & ~x195 & ~x221 & ~x279 & ~x304 & ~x335 & ~x336 & ~x388 & ~x389 & ~x391 & ~x417 & ~x447 & ~x448 & ~x450 & ~x473 & ~x475 & ~x476 & ~x477 & ~x504 & ~x505 & ~x530 & ~x533 & ~x559 & ~x585 & ~x589 & ~x613 & ~x669 & ~x670 & ~x674 & ~x699 & ~x702 & ~x755;
assign c4180 =  x236 &  x243 &  x262 &  x263 &  x272 &  x291 &  x298 &  x329 &  x375 &  x384 &  x407 &  x441 &  x458 &  x463 &  x498 &  x520 &  x582 &  x603 &  x606 &  x607 &  x608 &  x621 &  x634 &  x638 &  x653 &  x667 &  x695 &  x706 & ~x1 & ~x20 & ~x82 & ~x137 & ~x163 & ~x165 & ~x167 & ~x305 & ~x310 & ~x337 & ~x501 & ~x618 & ~x674 & ~x702 & ~x727 & ~x755 & ~x781;
assign c4182 =  x43 &  x206 &  x261 &  x265 &  x271 &  x322 &  x345 &  x349 &  x432 &  x460 &  x489 &  x494 &  x515 &  x548 &  x598 &  x627 &  x690 & ~x1 & ~x20 & ~x28 & ~x62 & ~x108 & ~x169 & ~x225 & ~x252 & ~x303 & ~x304 & ~x305 & ~x307 & ~x331 & ~x367 & ~x419 & ~x421 & ~x473 & ~x502 & ~x668 & ~x672 & ~x706 & ~x734 & ~x778;
assign c4184 =  x97 &  x358 &  x488 & ~x3 & ~x9 & ~x22 & ~x25 & ~x26 & ~x27 & ~x31 & ~x33 & ~x49 & ~x52 & ~x54 & ~x55 & ~x57 & ~x78 & ~x79 & ~x81 & ~x82 & ~x92 & ~x106 & ~x135 & ~x163 & ~x165 & ~x169 & ~x171 & ~x223 & ~x224 & ~x226 & ~x281 & ~x306 & ~x334 & ~x360 & ~x362 & ~x363 & ~x389 & ~x392 & ~x393 & ~x394 & ~x417 & ~x447 & ~x448 & ~x449 & ~x474 & ~x475 & ~x477 & ~x502 & ~x532 & ~x533 & ~x558 & ~x587 & ~x615 & ~x643 & ~x756 & ~x763;
assign c4186 =  x126 &  x268 &  x315 &  x355 &  x412 &  x424 &  x434 &  x458 &  x488 &  x520 &  x538 &  x541 &  x549 &  x571 &  x575 &  x578 &  x650 & ~x1 & ~x3 & ~x23 & ~x30 & ~x52 & ~x60 & ~x61 & ~x62 & ~x85 & ~x88 & ~x560 & ~x698;
assign c4188 =  x98 &  x384 &  x385 &  x441 &  x497 & ~x0 & ~x1 & ~x3 & ~x4 & ~x6 & ~x7 & ~x8 & ~x19 & ~x25 & ~x26 & ~x29 & ~x30 & ~x35 & ~x48 & ~x51 & ~x52 & ~x53 & ~x54 & ~x57 & ~x59 & ~x81 & ~x83 & ~x84 & ~x85 & ~x86 & ~x88 & ~x90 & ~x106 & ~x107 & ~x108 & ~x109 & ~x111 & ~x114 & ~x115 & ~x116 & ~x117 & ~x135 & ~x136 & ~x137 & ~x139 & ~x140 & ~x144 & ~x145 & ~x164 & ~x165 & ~x166 & ~x168 & ~x169 & ~x171 & ~x193 & ~x198 & ~x221 & ~x222 & ~x223 & ~x224 & ~x225 & ~x226 & ~x228 & ~x249 & ~x250 & ~x251 & ~x253 & ~x255 & ~x276 & ~x277 & ~x279 & ~x283 & ~x307 & ~x310 & ~x333 & ~x335 & ~x338 & ~x363 & ~x367 & ~x389 & ~x390 & ~x391 & ~x392 & ~x395 & ~x423 & ~x447 & ~x449 & ~x451 & ~x473 & ~x474 & ~x475 & ~x476 & ~x501 & ~x530 & ~x533 & ~x559 & ~x560 & ~x586 & ~x613 & ~x615 & ~x616 & ~x617 & ~x641 & ~x642 & ~x643 & ~x645 & ~x673 & ~x674 & ~x702 & ~x728 & ~x729 & ~x736 & ~x737 & ~x738 & ~x740 & ~x742 & ~x743 & ~x745 & ~x746 & ~x755 & ~x757 & ~x759 & ~x765 & ~x767 & ~x769 & ~x772 & ~x773 & ~x774 & ~x775 & ~x776 & ~x782 & ~x783;
assign c4190 =  x261 &  x405 &  x462 & ~x4 & ~x85 & ~x172 & ~x195 & ~x201 & ~x282 & ~x304 & ~x332 & ~x447 & ~x648 & ~x650 & ~x679 & ~x735 & ~x774;
assign c4192 = ~x1 & ~x6 & ~x8 & ~x9 & ~x10 & ~x17 & ~x20 & ~x24 & ~x25 & ~x27 & ~x30 & ~x32 & ~x49 & ~x50 & ~x56 & ~x59 & ~x63 & ~x77 & ~x78 & ~x89 & ~x106 & ~x107 & ~x114 & ~x116 & ~x138 & ~x140 & ~x142 & ~x143 & ~x163 & ~x164 & ~x166 & ~x167 & ~x192 & ~x219 & ~x220 & ~x228 & ~x255 & ~x309 & ~x311 & ~x332 & ~x362 & ~x365 & ~x366 & ~x389 & ~x392 & ~x393 & ~x395 & ~x420 & ~x449 & ~x507 & ~x530 & ~x531 & ~x557 & ~x559 & ~x563 & ~x585 & ~x588 & ~x590 & ~x614 & ~x615 & ~x618 & ~x643 & ~x672 & ~x674 & ~x675 & ~x690 & ~x691 & ~x701 & ~x702 & ~x727 & ~x729 & ~x736 & ~x739 & ~x741 & ~x745 & ~x746 & ~x757 & ~x766 & ~x772 & ~x774 & ~x780 & ~x782;
assign c4194 =  x43 &  x98 & ~x6 & ~x8 & ~x24 & ~x48 & ~x59 & ~x144 & ~x196 & ~x199 & ~x200 & ~x221 & ~x248 & ~x250 & ~x308 & ~x311 & ~x392 & ~x395 & ~x419 & ~x448 & ~x475 & ~x476 & ~x479 & ~x504 & ~x532 & ~x535 & ~x585 & ~x646 & ~x674 & ~x702 & ~x746 & ~x754 & ~x759 & ~x774 & ~x776;
assign c4196 =  x376 &  x463 &  x487 &  x547 & ~x1 & ~x2 & ~x5 & ~x9 & ~x22 & ~x23 & ~x24 & ~x25 & ~x27 & ~x28 & ~x30 & ~x31 & ~x35 & ~x36 & ~x53 & ~x56 & ~x57 & ~x60 & ~x79 & ~x80 & ~x81 & ~x90 & ~x106 & ~x107 & ~x113 & ~x133 & ~x143 & ~x145 & ~x162 & ~x163 & ~x165 & ~x169 & ~x170 & ~x192 & ~x195 & ~x197 & ~x198 & ~x219 & ~x222 & ~x224 & ~x225 & ~x254 & ~x255 & ~x276 & ~x277 & ~x280 & ~x281 & ~x283 & ~x305 & ~x308 & ~x311 & ~x335 & ~x338 & ~x361 & ~x362 & ~x363 & ~x366 & ~x391 & ~x392 & ~x394 & ~x419 & ~x421 & ~x450 & ~x474 & ~x475 & ~x535 & ~x559 & ~x560 & ~x561 & ~x616 & ~x644 & ~x646 & ~x700 & ~x728 & ~x748 & ~x754 & ~x765 & ~x766 & ~x767 & ~x774 & ~x776 & ~x781;
assign c4198 =  x209 &  x780 & ~x49;
assign c4200 =  x375 &  x430 &  x492 &  x650 & ~x5 & ~x37 & ~x51 & ~x52 & ~x53 & ~x62 & ~x63 & ~x88 & ~x143 & ~x166 & ~x193 & ~x196 & ~x252 & ~x278 & ~x283 & ~x306 & ~x334 & ~x363 & ~x422 & ~x502 & ~x504 & ~x561 & ~x616 & ~x617 & ~x642 & ~x643 & ~x644 & ~x673 & ~x698 & ~x754 & ~x772;
assign c4202 =  x41 &  x45 &  x158 &  x207 &  x238 &  x528 &  x567 &  x665 & ~x6 & ~x137 & ~x279 & ~x307 & ~x308 & ~x446 & ~x448 & ~x756;
assign c4204 =  x203 &  x237 &  x315 &  x371 &  x376 &  x385 &  x442 &  x486 &  x515 &  x542 &  x569 &  x600 &  x724 & ~x0 & ~x5 & ~x33 & ~x51 & ~x52 & ~x55 & ~x61 & ~x77 & ~x89 & ~x144 & ~x171 & ~x195 & ~x220 & ~x224 & ~x251 & ~x280 & ~x394 & ~x421 & ~x446 & ~x448 & ~x504 & ~x532 & ~x617;
assign c4206 =  x416 & ~x113 & ~x142 & ~x721;
assign c4208 =  x489 & ~x6 & ~x9 & ~x18 & ~x26 & ~x37 & ~x83 & ~x144 & ~x194 & ~x196 & ~x281 & ~x333 & ~x395 & ~x476 & ~x506 & ~x531 & ~x534 & ~x562 & ~x587 & ~x589 & ~x613 & ~x643 & ~x671 & ~x700 & ~x702 & ~x709 & ~x737 & ~x739 & ~x741 & ~x755 & ~x768;
assign c4210 =  x43 &  x94 &  x209 &  x261 &  x271 &  x289 &  x296 &  x298 &  x299 &  x320 &  x375 &  x376 &  x402 &  x405 &  x409 &  x433 &  x461 &  x486 &  x488 &  x489 &  x517 &  x545 &  x599 &  x600 &  x601 &  x626 &  x632 &  x654 &  x655 &  x658 &  x683 &  x686 & ~x4 & ~x20 & ~x29 & ~x34 & ~x50 & ~x60 & ~x111 & ~x113 & ~x116 & ~x138 & ~x142 & ~x144 & ~x163 & ~x171 & ~x220 & ~x222 & ~x224 & ~x226 & ~x248 & ~x249 & ~x250 & ~x276 & ~x281 & ~x282 & ~x283 & ~x304 & ~x305 & ~x307 & ~x333 & ~x337 & ~x338 & ~x340 & ~x365 & ~x388 & ~x389 & ~x392 & ~x446 & ~x449 & ~x472 & ~x473 & ~x475 & ~x476 & ~x478 & ~x479 & ~x503 & ~x529 & ~x533 & ~x560 & ~x561 & ~x585 & ~x587 & ~x588 & ~x589 & ~x618 & ~x671 & ~x673 & ~x675 & ~x699 & ~x700 & ~x728 & ~x729 & ~x730 & ~x750 & ~x752 & ~x754 & ~x757 & ~x777 & ~x779 & ~x780 & ~x781;
assign c4212 =  x197;
assign c4214 =  x261 &  x289 &  x356 &  x546 & ~x0 & ~x20 & ~x27 & ~x50 & ~x51 & ~x59 & ~x79 & ~x84 & ~x85 & ~x195 & ~x197 & ~x225 & ~x253 & ~x279 & ~x280 & ~x284 & ~x306 & ~x332 & ~x338 & ~x361 & ~x417 & ~x445 & ~x700 & ~x701 & ~x705 & ~x727 & ~x733 & ~x734 & ~x750 & ~x751 & ~x755 & ~x782 & ~x783;
assign c4216 =  x242 &  x270 &  x345 &  x461 &  x546 & ~x48 & ~x111 & ~x197 & ~x225 & ~x247 & ~x283 & ~x331 & ~x332 & ~x336 & ~x339 & ~x366 & ~x391 & ~x416 & ~x651 & ~x652;
assign c4218 = ~x2 & ~x6 & ~x7 & ~x8 & ~x9 & ~x10 & ~x20 & ~x22 & ~x24 & ~x25 & ~x28 & ~x31 & ~x56 & ~x57 & ~x84 & ~x109 & ~x111 & ~x115 & ~x135 & ~x138 & ~x141 & ~x165 & ~x193 & ~x198 & ~x227 & ~x249 & ~x255 & ~x309 & ~x365 & ~x419 & ~x447 & ~x476 & ~x503 & ~x531 & ~x559 & ~x572 & ~x587 & ~x671 & ~x698 & ~x728 & ~x756 & ~x757 & ~x764;
assign c4220 =  x12 &  x269 &  x320 &  x327 &  x345 &  x378 &  x424 &  x457 &  x492 &  x676 & ~x88 & ~x114 & ~x135 & ~x193 & ~x196 & ~x277 & ~x308 & ~x365 & ~x476 & ~x532 & ~x699;
assign c4222 =  x13 &  x323 &  x443 &  x471 &  x523 &  x608 &  x650 & ~x56 & ~x422 & ~x506 & ~x558 & ~x700 & ~x782;
assign c4224 =  x42 &  x230 &  x415 &  x428 &  x513 &  x581 &  x596 &  x637 &  x665 &  x744 & ~x24 & ~x31 & ~x81 & ~x674 & ~x758;
assign c4226 = ~x0 & ~x2 & ~x3 & ~x9 & ~x10 & ~x18 & ~x19 & ~x22 & ~x23 & ~x25 & ~x31 & ~x32 & ~x36 & ~x37 & ~x48 & ~x51 & ~x53 & ~x54 & ~x55 & ~x57 & ~x58 & ~x59 & ~x61 & ~x79 & ~x80 & ~x83 & ~x106 & ~x109 & ~x110 & ~x114 & ~x115 & ~x137 & ~x139 & ~x142 & ~x164 & ~x166 & ~x167 & ~x168 & ~x170 & ~x171 & ~x195 & ~x221 & ~x222 & ~x227 & ~x250 & ~x278 & ~x279 & ~x280 & ~x281 & ~x304 & ~x305 & ~x307 & ~x309 & ~x335 & ~x336 & ~x366 & ~x389 & ~x390 & ~x391 & ~x392 & ~x394 & ~x395 & ~x417 & ~x418 & ~x422 & ~x445 & ~x447 & ~x450 & ~x451 & ~x476 & ~x503 & ~x529 & ~x530 & ~x535 & ~x559 & ~x561 & ~x614 & ~x618 & ~x643 & ~x645 & ~x670 & ~x673 & ~x708 & ~x709 & ~x712 & ~x718 & ~x728 & ~x729 & ~x738 & ~x739 & ~x740 & ~x741 & ~x742 & ~x746 & ~x747 & ~x748 & ~x754 & ~x756 & ~x758 & ~x764 & ~x769 & ~x770 & ~x774 & ~x776 & ~x781 & ~x782;
assign c4228 =  x701;
assign c4230 =  x602 & ~x4 & ~x114 & ~x129 & ~x255 & ~x474 & ~x534 & ~x736 & ~x766;
assign c4232 =  x317 &  x434 &  x461 & ~x7 & ~x21 & ~x23 & ~x46 & ~x55 & ~x57 & ~x77 & ~x80 & ~x117 & ~x132 & ~x135 & ~x139 & ~x144 & ~x146 & ~x172 & ~x173 & ~x197 & ~x199 & ~x251 & ~x309 & ~x367 & ~x390 & ~x418 & ~x419 & ~x423 & ~x448 & ~x479 & ~x501 & ~x557 & ~x563 & ~x585 & ~x591 & ~x728 & ~x729 & ~x782;
assign c4234 =  x42 &  x43 &  x70 &  x71 &  x378 & ~x1 & ~x2 & ~x3 & ~x5 & ~x7 & ~x8 & ~x21 & ~x24 & ~x26 & ~x29 & ~x31 & ~x32 & ~x33 & ~x34 & ~x51 & ~x52 & ~x60 & ~x85 & ~x86 & ~x87 & ~x107 & ~x108 & ~x110 & ~x111 & ~x112 & ~x116 & ~x139 & ~x140 & ~x141 & ~x142 & ~x143 & ~x167 & ~x169 & ~x171 & ~x193 & ~x194 & ~x195 & ~x198 & ~x221 & ~x222 & ~x226 & ~x250 & ~x251 & ~x252 & ~x254 & ~x276 & ~x279 & ~x282 & ~x306 & ~x309 & ~x310 & ~x332 & ~x334 & ~x338 & ~x366 & ~x390 & ~x421 & ~x422 & ~x445 & ~x448 & ~x449 & ~x450 & ~x474 & ~x475 & ~x476 & ~x503 & ~x504 & ~x531 & ~x557 & ~x558 & ~x559 & ~x560 & ~x585 & ~x588 & ~x616 & ~x617 & ~x618 & ~x641 & ~x645 & ~x670 & ~x672 & ~x698 & ~x701 & ~x713 & ~x737 & ~x738 & ~x739 & ~x765 & ~x767 & ~x768 & ~x771 & ~x775 & ~x782 & ~x783;
assign c4236 =  x262 &  x271 &  x289 &  x292 &  x298 &  x319 &  x326 &  x354 &  x384 &  x515 &  x548 & ~x10 & ~x21 & ~x50 & ~x57 & ~x61 & ~x86 & ~x145 & ~x168 & ~x194 & ~x225 & ~x256 & ~x280 & ~x308 & ~x362 & ~x366 & ~x390 & ~x395 & ~x450 & ~x478 & ~x533 & ~x534 & ~x558 & ~x561 & ~x616 & ~x645 & ~x734 & ~x751 & ~x756 & ~x779;
assign c4238 =  x232 &  x267 &  x295 &  x301 &  x372 &  x403 &  x494 &  x553 &  x580 &  x581 &  x603 &  x720 & ~x1 & ~x27 & ~x50 & ~x53 & ~x110 & ~x140 & ~x141 & ~x165 & ~x193 & ~x280 & ~x304 & ~x305 & ~x310 & ~x332 & ~x393 & ~x418 & ~x445 & ~x451 & ~x473 & ~x503 & ~x562 & ~x675 & ~x726 & ~x780 & ~x783;
assign c4240 =  x247 &  x286 &  x638 & ~x59 & ~x165 & ~x225 & ~x306;
assign c4242 =  x399 &  x461 & ~x1 & ~x2 & ~x5 & ~x8 & ~x22 & ~x23 & ~x26 & ~x28 & ~x32 & ~x37 & ~x46 & ~x53 & ~x56 & ~x60 & ~x63 & ~x78 & ~x79 & ~x84 & ~x87 & ~x113 & ~x136 & ~x142 & ~x166 & ~x192 & ~x194 & ~x196 & ~x198 & ~x199 & ~x249 & ~x252 & ~x276 & ~x283 & ~x305 & ~x308 & ~x310 & ~x336 & ~x337 & ~x362 & ~x363 & ~x364 & ~x365 & ~x390 & ~x476 & ~x559 & ~x587 & ~x615 & ~x643 & ~x644 & ~x671 & ~x699 & ~x737 & ~x743 & ~x744 & ~x745 & ~x757 & ~x759 & ~x768 & ~x769 & ~x774;
assign c4244 =  x295 &  x527 &  x662 &  x748 & ~x27 & ~x31 & ~x81 & ~x111 & ~x166 & ~x196 & ~x224 & ~x251 & ~x276 & ~x283 & ~x335 & ~x336 & ~x339 & ~x417 & ~x447 & ~x530 & ~x531 & ~x560 & ~x617 & ~x700;
assign c4246 =  x154 &  x459 &  x517 &  x766 & ~x10 & ~x60 & ~x87 & ~x105 & ~x139 & ~x170 & ~x250 & ~x360 & ~x362 & ~x645 & ~x727 & ~x754;
assign c4248 =  x725;
assign c4250 =  x377 &  x551 &  x581 &  x599 & ~x28 & ~x32 & ~x56 & ~x60 & ~x82 & ~x107 & ~x168 & ~x170 & ~x195 & ~x198 & ~x250 & ~x251 & ~x254 & ~x309 & ~x335 & ~x336 & ~x559 & ~x588 & ~x615 & ~x671 & ~x700 & ~x725 & ~x733 & ~x734 & ~x750 & ~x758 & ~x778 & ~x782 & ~x783;
assign c4252 =  x70 & ~x10 & ~x18 & ~x36 & ~x198 & ~x255 & ~x300 & ~x446 & ~x478 & ~x558 & ~x614;
assign c4254 =  x355 &  x459 &  x462 &  x495 & ~x1 & ~x4 & ~x9 & ~x21 & ~x23 & ~x29 & ~x52 & ~x53 & ~x57 & ~x61 & ~x81 & ~x107 & ~x163 & ~x165 & ~x166 & ~x169 & ~x171 & ~x192 & ~x193 & ~x198 & ~x221 & ~x227 & ~x249 & ~x250 & ~x252 & ~x276 & ~x332 & ~x336 & ~x339 & ~x360 & ~x362 & ~x365 & ~x388 & ~x391 & ~x392 & ~x393 & ~x416 & ~x447 & ~x448 & ~x450 & ~x502 & ~x503 & ~x504 & ~x529 & ~x530 & ~x533 & ~x563 & ~x585 & ~x586 & ~x591 & ~x645 & ~x646 & ~x671 & ~x673 & ~x674 & ~x701 & ~x730 & ~x741 & ~x754 & ~x774;
assign c4256 =  x98 & ~x7 & ~x18 & ~x19 & ~x26 & ~x27 & ~x50 & ~x51 & ~x53 & ~x81 & ~x84 & ~x87 & ~x137 & ~x143 & ~x144 & ~x193 & ~x194 & ~x195 & ~x196 & ~x239 & ~x252 & ~x254 & ~x278 & ~x305 & ~x307 & ~x333 & ~x335 & ~x361 & ~x364 & ~x365 & ~x390 & ~x392 & ~x419 & ~x423 & ~x447 & ~x450 & ~x503 & ~x530 & ~x533 & ~x557 & ~x559 & ~x617 & ~x643 & ~x644 & ~x669 & ~x756;
assign c4258 =  x289 &  x317 &  x345 & ~x1 & ~x4 & ~x10 & ~x21 & ~x23 & ~x36 & ~x37 & ~x64 & ~x86 & ~x107 & ~x108 & ~x116 & ~x133 & ~x139 & ~x144 & ~x145 & ~x162 & ~x167 & ~x190 & ~x191 & ~x218 & ~x222 & ~x224 & ~x226 & ~x247 & ~x248 & ~x257 & ~x277 & ~x280 & ~x283 & ~x285 & ~x331 & ~x333 & ~x338 & ~x361 & ~x362 & ~x366 & ~x396 & ~x415 & ~x422 & ~x450 & ~x451 & ~x471 & ~x472 & ~x477 & ~x479 & ~x501 & ~x504 & ~x505 & ~x529 & ~x646 & ~x675 & ~x701 & ~x729 & ~x753 & ~x754 & ~x765 & ~x781;
assign c4260 =  x219 &  x638 &  x696 &  x750 & ~x6 & ~x448 & ~x769;
assign c4262 =  x754;
assign c4264 =  x270 & ~x2 & ~x4 & ~x8 & ~x10 & ~x17 & ~x18 & ~x19 & ~x25 & ~x26 & ~x30 & ~x34 & ~x36 & ~x47 & ~x48 & ~x63 & ~x85 & ~x86 & ~x87 & ~x90 & ~x91 & ~x109 & ~x116 & ~x133 & ~x138 & ~x140 & ~x141 & ~x146 & ~x161 & ~x163 & ~x164 & ~x169 & ~x173 & ~x190 & ~x197 & ~x198 & ~x219 & ~x225 & ~x227 & ~x248 & ~x249 & ~x251 & ~x277 & ~x280 & ~x304 & ~x306 & ~x308 & ~x334 & ~x339 & ~x363 & ~x364 & ~x365 & ~x389 & ~x390 & ~x418 & ~x445 & ~x448 & ~x505 & ~x587 & ~x589 & ~x673 & ~x703 & ~x730 & ~x750 & ~x752 & ~x754 & ~x762 & ~x777;
assign c4266 =  x235 &  x346 &  x412 &  x497 &  x551 &  x569 &  x598 &  x609 &  x621 &  x624 &  x628 &  x665 &  x684 &  x711 & ~x3 & ~x19 & ~x26 & ~x28 & ~x52 & ~x169 & ~x277 & ~x336 & ~x361 & ~x388 & ~x476 & ~x502 & ~x503 & ~x506 & ~x530 & ~x617 & ~x647 & ~x702 & ~x754;
assign c4268 =  x14 &  x40 &  x44 &  x45 &  x99 &  x180 &  x213 &  x235 &  x267 &  x329 &  x405 &  x481 &  x551 &  x565 &  x566 & ~x2 & ~x52 & ~x62 & ~x254 & ~x307 & ~x420 & ~x533;
assign c4270 =  x42 &  x70 &  x286 &  x314 &  x431 &  x433 &  x440 &  x454 &  x483 &  x484 &  x572 &  x621 &  x622 &  x625 &  x628 &  x637 & ~x4 & ~x23 & ~x141 & ~x144 & ~x169 & ~x192 & ~x222 & ~x224 & ~x278 & ~x338 & ~x534 & ~x559 & ~x560 & ~x586 & ~x615 & ~x616 & ~x643 & ~x783;
assign c4272 =  x322 &  x343 &  x592 & ~x26 & ~x27 & ~x28 & ~x49 & ~x57 & ~x63 & ~x76 & ~x77 & ~x78 & ~x107 & ~x115 & ~x136 & ~x172 & ~x192 & ~x194 & ~x197 & ~x221 & ~x253 & ~x278 & ~x281 & ~x282 & ~x283 & ~x445 & ~x474 & ~x503 & ~x778;
assign c4274 =  x322 &  x384 &  x541 &  x551 &  x610 &  x634 &  x704 &  x733 & ~x6 & ~x9 & ~x20 & ~x48 & ~x49 & ~x56 & ~x58 & ~x59 & ~x63 & ~x82 & ~x114 & ~x140 & ~x165 & ~x167 & ~x169 & ~x170 & ~x171 & ~x194 & ~x222 & ~x226 & ~x253 & ~x389 & ~x390 & ~x419 & ~x449 & ~x478 & ~x502 & ~x530 & ~x561 & ~x645 & ~x646 & ~x672 & ~x673 & ~x698 & ~x700 & ~x766 & ~x768 & ~x770;
assign c4276 = ~x10 & ~x18 & ~x20 & ~x61 & ~x85 & ~x115 & ~x136 & ~x164 & ~x171 & ~x196 & ~x231 & ~x364 & ~x419 & ~x459 & ~x533 & ~x587 & ~x644;
assign c4278 =  x321 &  x350 &  x400 &  x462 &  x467 &  x599 &  x660 &  x689 &  x736 & ~x59 & ~x107 & ~x108 & ~x191 & ~x251 & ~x256 & ~x282 & ~x476 & ~x560 & ~x562 & ~x614 & ~x615 & ~x675 & ~x728;
assign c4280 =  x359 &  x623 &  x680 & ~x3 & ~x62 & ~x278;
assign c4282 =  x43 &  x124 &  x154 &  x177 &  x181 &  x186 &  x206 &  x208 &  x211 &  x212 &  x214 &  x215 &  x233 &  x234 &  x235 &  x239 &  x261 &  x262 &  x264 &  x265 &  x269 &  x270 &  x271 &  x291 &  x294 &  x295 &  x297 &  x317 &  x319 &  x323 &  x344 &  x345 &  x347 &  x352 &  x353 &  x356 &  x372 &  x373 &  x375 &  x381 &  x400 &  x401 &  x402 &  x404 &  x405 &  x408 &  x409 &  x411 &  x429 &  x432 &  x433 &  x435 &  x437 &  x439 &  x458 &  x461 &  x462 &  x465 &  x466 &  x467 &  x489 &  x491 &  x492 &  x493 &  x494 &  x513 &  x514 &  x516 &  x517 &  x519 &  x521 &  x546 &  x549 &  x571 &  x572 &  x577 & ~x1 & ~x2 & ~x4 & ~x7 & ~x20 & ~x26 & ~x27 & ~x28 & ~x30 & ~x32 & ~x33 & ~x50 & ~x51 & ~x53 & ~x54 & ~x55 & ~x56 & ~x60 & ~x78 & ~x79 & ~x81 & ~x83 & ~x84 & ~x85 & ~x110 & ~x111 & ~x118 & ~x139 & ~x142 & ~x143 & ~x165 & ~x169 & ~x170 & ~x191 & ~x195 & ~x196 & ~x220 & ~x222 & ~x225 & ~x247 & ~x248 & ~x250 & ~x252 & ~x254 & ~x256 & ~x276 & ~x277 & ~x278 & ~x279 & ~x281 & ~x282 & ~x283 & ~x284 & ~x304 & ~x305 & ~x310 & ~x311 & ~x332 & ~x340 & ~x360 & ~x362 & ~x363 & ~x392 & ~x393 & ~x394 & ~x418 & ~x419 & ~x421 & ~x422 & ~x423 & ~x446 & ~x448 & ~x449 & ~x472 & ~x476 & ~x479 & ~x501 & ~x505 & ~x531 & ~x558 & ~x559 & ~x560 & ~x585 & ~x590 & ~x591 & ~x613 & ~x617 & ~x640 & ~x641 & ~x642 & ~x672 & ~x673 & ~x674 & ~x700 & ~x701 & ~x703 & ~x727 & ~x728 & ~x729 & ~x753 & ~x757 & ~x758 & ~x759 & ~x764;
assign c4284 = ~x1 & ~x7 & ~x8 & ~x25 & ~x28 & ~x32 & ~x52 & ~x78 & ~x83 & ~x84 & ~x115 & ~x164 & ~x192 & ~x197 & ~x249 & ~x253 & ~x269 & ~x297 & ~x298 & ~x305 & ~x309 & ~x333 & ~x364 & ~x390 & ~x418 & ~x450 & ~x559 & ~x561 & ~x586 & ~x587 & ~x670 & ~x765 & ~x768 & ~x769 & ~x771;
assign c4286 =  x151 &  x184 &  x202 &  x211 &  x319 &  x370 &  x413 &  x438 &  x439 &  x471 &  x491 &  x495 &  x554 & ~x6 & ~x77 & ~x80 & ~x81 & ~x82 & ~x250 & ~x533 & ~x728;
assign c4288 =  x380 &  x408 &  x639 &  x733 & ~x2 & ~x3 & ~x20 & ~x29 & ~x30 & ~x31 & ~x37 & ~x51 & ~x53 & ~x56 & ~x59 & ~x61 & ~x113 & ~x143 & ~x167 & ~x221 & ~x251 & ~x255 & ~x280 & ~x306 & ~x309 & ~x310 & ~x334 & ~x394 & ~x475 & ~x476 & ~x530 & ~x558 & ~x559 & ~x588 & ~x617 & ~x644 & ~x700 & ~x701 & ~x702 & ~x727 & ~x744 & ~x745 & ~x755 & ~x766 & ~x770 & ~x774 & ~x775 & ~x781;
assign c4290 =  x489 &  x566 &  x658 & ~x1 & ~x5 & ~x30 & ~x58 & ~x85 & ~x110 & ~x171 & ~x192 & ~x193 & ~x198 & ~x249 & ~x281 & ~x282 & ~x283 & ~x310 & ~x390 & ~x392 & ~x420 & ~x446 & ~x447 & ~x477 & ~x588 & ~x722 & ~x724 & ~x780;
assign c4292 = ~x3 & ~x7 & ~x8 & ~x19 & ~x21 & ~x30 & ~x31 & ~x33 & ~x36 & ~x50 & ~x54 & ~x55 & ~x58 & ~x79 & ~x80 & ~x82 & ~x85 & ~x86 & ~x87 & ~x88 & ~x107 & ~x108 & ~x110 & ~x113 & ~x162 & ~x165 & ~x166 & ~x169 & ~x191 & ~x193 & ~x196 & ~x197 & ~x198 & ~x199 & ~x200 & ~x208 & ~x222 & ~x226 & ~x250 & ~x251 & ~x277 & ~x278 & ~x308 & ~x309 & ~x332 & ~x339 & ~x363 & ~x367 & ~x390 & ~x395 & ~x423 & ~x445 & ~x447 & ~x449 & ~x475 & ~x478 & ~x479 & ~x505 & ~x529 & ~x530 & ~x531 & ~x533 & ~x534 & ~x560 & ~x561 & ~x616 & ~x644 & ~x646 & ~x670 & ~x671 & ~x672 & ~x702 & ~x725 & ~x726 & ~x754 & ~x756 & ~x759 & ~x764 & ~x765 & ~x775 & ~x776 & ~x783;
assign c4294 = ~x2 & ~x7 & ~x8 & ~x19 & ~x30 & ~x54 & ~x88 & ~x108 & ~x115 & ~x134 & ~x138 & ~x163 & ~x197 & ~x200 & ~x249 & ~x264 & ~x282 & ~x297 & ~x307 & ~x308 & ~x309 & ~x334 & ~x361 & ~x394 & ~x479 & ~x502 & ~x530 & ~x534 & ~x562 & ~x586 & ~x616 & ~x765 & ~x771;
assign c4296 =  x15 &  x327 & ~x0 & ~x2 & ~x22 & ~x29 & ~x53 & ~x58 & ~x59 & ~x79 & ~x81 & ~x83 & ~x114 & ~x140 & ~x141 & ~x142 & ~x166 & ~x167 & ~x193 & ~x196 & ~x224 & ~x249 & ~x280 & ~x282 & ~x306 & ~x363 & ~x390 & ~x559 & ~x587 & ~x615 & ~x643 & ~x711 & ~x755 & ~x768 & ~x769;
assign c4298 = ~x1 & ~x9 & ~x10 & ~x18 & ~x19 & ~x23 & ~x25 & ~x27 & ~x30 & ~x31 & ~x35 & ~x36 & ~x51 & ~x52 & ~x54 & ~x55 & ~x60 & ~x62 & ~x81 & ~x84 & ~x88 & ~x106 & ~x107 & ~x108 & ~x109 & ~x110 & ~x112 & ~x114 & ~x116 & ~x135 & ~x137 & ~x144 & ~x169 & ~x170 & ~x192 & ~x194 & ~x195 & ~x196 & ~x197 & ~x199 & ~x200 & ~x222 & ~x223 & ~x224 & ~x226 & ~x227 & ~x249 & ~x251 & ~x253 & ~x254 & ~x256 & ~x277 & ~x279 & ~x280 & ~x282 & ~x283 & ~x284 & ~x305 & ~x307 & ~x333 & ~x334 & ~x336 & ~x337 & ~x362 & ~x365 & ~x367 & ~x378 & ~x392 & ~x393 & ~x394 & ~x395 & ~x419 & ~x420 & ~x423 & ~x446 & ~x450 & ~x451 & ~x475 & ~x476 & ~x503 & ~x531 & ~x533 & ~x559 & ~x562 & ~x587 & ~x588 & ~x589 & ~x590 & ~x614 & ~x616 & ~x617 & ~x618 & ~x642 & ~x672 & ~x673 & ~x728 & ~x754 & ~x757 & ~x776;
assign c4300 =  x70 & ~x2 & ~x4 & ~x5 & ~x6 & ~x19 & ~x22 & ~x25 & ~x28 & ~x32 & ~x81 & ~x109 & ~x113 & ~x114 & ~x141 & ~x166 & ~x193 & ~x197 & ~x223 & ~x281 & ~x307 & ~x335 & ~x337 & ~x390 & ~x447 & ~x448 & ~x475 & ~x476 & ~x502 & ~x504 & ~x587 & ~x615 & ~x700 & ~x721 & ~x736 & ~x737 & ~x738 & ~x740 & ~x741 & ~x744 & ~x746 & ~x748 & ~x769 & ~x771 & ~x774;
assign c4302 =  x40 &  x173 &  x340 &  x552 &  x648 & ~x475;
assign c4304 =  x40 &  x43 &  x70 &  x98 &  x733 &  x750 & ~x0 & ~x2 & ~x3 & ~x5 & ~x6 & ~x7 & ~x19 & ~x20 & ~x26 & ~x30 & ~x31 & ~x48 & ~x49 & ~x50 & ~x51 & ~x52 & ~x53 & ~x54 & ~x55 & ~x56 & ~x57 & ~x58 & ~x59 & ~x60 & ~x62 & ~x84 & ~x85 & ~x88 & ~x106 & ~x111 & ~x115 & ~x140 & ~x141 & ~x142 & ~x143 & ~x167 & ~x170 & ~x172 & ~x192 & ~x195 & ~x196 & ~x199 & ~x221 & ~x223 & ~x255 & ~x279 & ~x280 & ~x282 & ~x304 & ~x308 & ~x311 & ~x334 & ~x336 & ~x338 & ~x360 & ~x361 & ~x388 & ~x390 & ~x392 & ~x393 & ~x394 & ~x418 & ~x420 & ~x422 & ~x445 & ~x446 & ~x448 & ~x449 & ~x450 & ~x451 & ~x476 & ~x479 & ~x505 & ~x506 & ~x507 & ~x530 & ~x534 & ~x558 & ~x559 & ~x560 & ~x562 & ~x563 & ~x587 & ~x588 & ~x589 & ~x613 & ~x617 & ~x641 & ~x643 & ~x644 & ~x645 & ~x646 & ~x647 & ~x669 & ~x673 & ~x698 & ~x699 & ~x700 & ~x701 & ~x725 & ~x728 & ~x730 & ~x737 & ~x738 & ~x739 & ~x742 & ~x744 & ~x745 & ~x746 & ~x747 & ~x753 & ~x756 & ~x757 & ~x758 & ~x765 & ~x767 & ~x769 & ~x770 & ~x773 & ~x774 & ~x782;
assign c4306 =  x154 &  x229 &  x406 &  x440 &  x455 &  x489 &  x539 & ~x2 & ~x51 & ~x86 & ~x307 & ~x337 & ~x363 & ~x761 & ~x782;
assign c4308 =  x42 &  x152 &  x179 &  x289 &  x415 &  x435 &  x453 &  x482 &  x567 &  x595 &  x597 &  x665 &  x666 & ~x5 & ~x137 & ~x138 & ~x278 & ~x420 & ~x532 & ~x589 & ~x615;
assign c4310 =  x126 & ~x435;
assign c4312 =  x154 &  x300 &  x356 & ~x6 & ~x9 & ~x18 & ~x19 & ~x27 & ~x31 & ~x32 & ~x36 & ~x48 & ~x51 & ~x58 & ~x59 & ~x79 & ~x81 & ~x82 & ~x83 & ~x87 & ~x105 & ~x106 & ~x110 & ~x111 & ~x113 & ~x115 & ~x116 & ~x132 & ~x133 & ~x134 & ~x138 & ~x139 & ~x146 & ~x164 & ~x165 & ~x166 & ~x167 & ~x168 & ~x170 & ~x171 & ~x192 & ~x194 & ~x198 & ~x219 & ~x220 & ~x223 & ~x225 & ~x226 & ~x228 & ~x248 & ~x249 & ~x250 & ~x253 & ~x255 & ~x278 & ~x280 & ~x281 & ~x282 & ~x283 & ~x304 & ~x306 & ~x308 & ~x311 & ~x312 & ~x332 & ~x336 & ~x337 & ~x338 & ~x339 & ~x363 & ~x391 & ~x393 & ~x394 & ~x417 & ~x418 & ~x420 & ~x423 & ~x446 & ~x447 & ~x474 & ~x479 & ~x502 & ~x503 & ~x504 & ~x505 & ~x507 & ~x530 & ~x557 & ~x561 & ~x590 & ~x616 & ~x618 & ~x643 & ~x644 & ~x646 & ~x701 & ~x728 & ~x729 & ~x730 & ~x753 & ~x756 & ~x758;
assign c4314 =  x42 &  x70 &  x428 & ~x0 & ~x1 & ~x2 & ~x3 & ~x4 & ~x5 & ~x6 & ~x7 & ~x9 & ~x10 & ~x17 & ~x18 & ~x19 & ~x20 & ~x23 & ~x24 & ~x25 & ~x26 & ~x27 & ~x29 & ~x30 & ~x31 & ~x33 & ~x35 & ~x36 & ~x48 & ~x49 & ~x50 & ~x51 & ~x52 & ~x55 & ~x56 & ~x57 & ~x58 & ~x60 & ~x61 & ~x62 & ~x76 & ~x78 & ~x79 & ~x80 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x86 & ~x87 & ~x88 & ~x89 & ~x90 & ~x105 & ~x106 & ~x107 & ~x108 & ~x109 & ~x112 & ~x114 & ~x115 & ~x116 & ~x117 & ~x118 & ~x134 & ~x135 & ~x136 & ~x137 & ~x138 & ~x139 & ~x140 & ~x141 & ~x142 & ~x143 & ~x144 & ~x145 & ~x163 & ~x164 & ~x165 & ~x166 & ~x167 & ~x168 & ~x169 & ~x171 & ~x172 & ~x189 & ~x191 & ~x192 & ~x193 & ~x194 & ~x195 & ~x196 & ~x197 & ~x198 & ~x199 & ~x201 & ~x220 & ~x223 & ~x225 & ~x227 & ~x228 & ~x229 & ~x248 & ~x249 & ~x250 & ~x251 & ~x252 & ~x254 & ~x255 & ~x276 & ~x277 & ~x278 & ~x279 & ~x280 & ~x281 & ~x282 & ~x284 & ~x304 & ~x305 & ~x306 & ~x307 & ~x308 & ~x310 & ~x332 & ~x333 & ~x335 & ~x336 & ~x337 & ~x338 & ~x339 & ~x360 & ~x361 & ~x362 & ~x363 & ~x364 & ~x365 & ~x366 & ~x367 & ~x389 & ~x390 & ~x391 & ~x392 & ~x393 & ~x394 & ~x395 & ~x417 & ~x418 & ~x419 & ~x420 & ~x421 & ~x422 & ~x423 & ~x444 & ~x445 & ~x446 & ~x447 & ~x448 & ~x450 & ~x472 & ~x473 & ~x474 & ~x475 & ~x476 & ~x477 & ~x502 & ~x503 & ~x504 & ~x505 & ~x506 & ~x508 & ~x528 & ~x529 & ~x530 & ~x531 & ~x532 & ~x533 & ~x534 & ~x535 & ~x556 & ~x557 & ~x559 & ~x560 & ~x561 & ~x562 & ~x585 & ~x586 & ~x587 & ~x588 & ~x590 & ~x613 & ~x615 & ~x616 & ~x617 & ~x618 & ~x619 & ~x644 & ~x646 & ~x647 & ~x669 & ~x670 & ~x671 & ~x673 & ~x674 & ~x675 & ~x697 & ~x699 & ~x701 & ~x703 & ~x726 & ~x728 & ~x729 & ~x730 & ~x731 & ~x752 & ~x753 & ~x755 & ~x756 & ~x757 & ~x758 & ~x759 & ~x775 & ~x776 & ~x781 & ~x782 & ~x783;
assign c4316 =  x286 &  x288 &  x321 &  x352 &  x460 &  x487 &  x620 &  x676 & ~x2 & ~x5 & ~x19 & ~x109 & ~x196 & ~x223 & ~x250 & ~x393 & ~x709;
assign c4318 =  x230 &  x312 &  x340 &  x424 &  x647 & ~x32 & ~x57 & ~x80 & ~x282 & ~x337 & ~x363 & ~x447 & ~x476 & ~x561 & ~x645;
assign c4320 = ~x232 & ~x292 & ~x393 & ~x474 & ~x765;
assign c4322 =  x203 &  x260 &  x267 &  x271 &  x298 &  x328 &  x358 &  x380 &  x399 &  x403 &  x407 &  x408 &  x440 &  x470 &  x519 &  x566 &  x576 &  x580 &  x596 &  x632 &  x636 &  x650 & ~x4 & ~x33 & ~x141 & ~x252 & ~x276 & ~x310 & ~x334 & ~x335 & ~x364 & ~x417 & ~x448 & ~x616 & ~x702 & ~x731 & ~x752;
assign c4324 =  x764 &  x773;
assign c4326 =  x275 &  x387 &  x552 &  x582 &  x694 &  x750 & ~x86 & ~x311 & ~x365 & ~x533 & ~x772 & ~x783;
assign c4328 =  x238 &  x344 &  x355 &  x357 &  x412 &  x465 &  x518 &  x539 &  x542 &  x545 &  x550 &  x567 &  x580 &  x606 &  x624 &  x660 & ~x8 & ~x9 & ~x33 & ~x56 & ~x57 & ~x133 & ~x143 & ~x163 & ~x168 & ~x197 & ~x224 & ~x227 & ~x255 & ~x279 & ~x305 & ~x306 & ~x308 & ~x389 & ~x446 & ~x448 & ~x504 & ~x531 & ~x560 & ~x673 & ~x675 & ~x700 & ~x702 & ~x728 & ~x755 & ~x758 & ~x759 & ~x781 & ~x782;
assign c4330 =  x208 &  x209 &  x235 &  x245 &  x321 &  x325 &  x327 &  x429 &  x438 &  x442 &  x466 &  x526 &  x542 &  x569 &  x605 &  x610 &  x631 &  x751 & ~x5 & ~x6 & ~x8 & ~x28 & ~x51 & ~x55 & ~x56 & ~x77 & ~x83 & ~x85 & ~x113 & ~x165 & ~x166 & ~x194 & ~x223 & ~x255 & ~x281 & ~x308 & ~x362 & ~x363 & ~x365 & ~x391 & ~x394 & ~x421 & ~x447 & ~x534 & ~x561 & ~x589 & ~x642 & ~x643 & ~x699 & ~x748 & ~x771;
assign c4332 =  x43 &  x270 &  x380 &  x434 &  x462 &  x543 & ~x6 & ~x18 & ~x56 & ~x77 & ~x173 & ~x219 & ~x451 & ~x623 & ~x650 & ~x763;
assign c4334 =  x228 &  x696 & ~x30 & ~x194 & ~x224 & ~x225 & ~x448 & ~x532;
assign c4336 =  x573 & ~x598;
assign c4338 =  x38 &  x180 &  x210 &  x231 &  x238 &  x267 &  x287 &  x293 &  x324 &  x341 &  x353 &  x369 &  x381 &  x406 &  x434 &  x436 &  x509 &  x570 &  x685 & ~x51 & ~x62 & ~x78 & ~x110 & ~x254 & ~x478 & ~x754;
assign c4340 =  x289 &  x327 & ~x22 & ~x33 & ~x54 & ~x80 & ~x113 & ~x116 & ~x143 & ~x201 & ~x279 & ~x333 & ~x389 & ~x479 & ~x501 & ~x562 & ~x563 & ~x623 & ~x652 & ~x673 & ~x700 & ~x705 & ~x731 & ~x734 & ~x759 & ~x776;
assign c4342 =  x126 & ~x9 & ~x60 & ~x78 & ~x83 & ~x140 & ~x167 & ~x194 & ~x306 & ~x360 & ~x361 & ~x432 & ~x584;
assign c4344 =  x43 &  x647 & ~x7 & ~x61 & ~x114 & ~x279;
assign c4346 =  x230 &  x570 &  x679 &  x733 & ~x61 & ~x87 & ~x114 & ~x169 & ~x198 & ~x249 & ~x253 & ~x310 & ~x422 & ~x479 & ~x700 & ~x768 & ~x775 & ~x781;
assign c4348 =  x259 &  x551 &  x593 &  x596 &  x604 &  x608 &  x707 & ~x28 & ~x60 & ~x79 & ~x83 & ~x138 & ~x144 & ~x169 & ~x172 & ~x193 & ~x196 & ~x200 & ~x364 & ~x418 & ~x419 & ~x449 & ~x502 & ~x505 & ~x530 & ~x558 & ~x644 & ~x674 & ~x675 & ~x703 & ~x757;
assign c4350 =  x174 &  x300 &  x407 &  x431 &  x549 &  x638 &  x732 & ~x9 & ~x20 & ~x84 & ~x139 & ~x167 & ~x389 & ~x391 & ~x417 & ~x505 & ~x533 & ~x728 & ~x738 & ~x746 & ~x766;
assign c4352 =  x43 &  x241 &  x378 &  x490 &  x518 &  x546 &  x602 &  x630 & ~x9 & ~x26 & ~x162 & ~x166 & ~x169 & ~x225 & ~x309 & ~x335 & ~x419 & ~x451 & ~x475 & ~x534 & ~x536 & ~x644 & ~x651 & ~x670 & ~x679 & ~x775;
assign c4354 =  x658 & ~x7 & ~x466 & ~x503 & ~x769;
assign c4356 = ~x4 & ~x10 & ~x18 & ~x30 & ~x33 & ~x46 & ~x58 & ~x64 & ~x75 & ~x85 & ~x87 & ~x112 & ~x114 & ~x139 & ~x144 & ~x168 & ~x192 & ~x195 & ~x221 & ~x223 & ~x227 & ~x283 & ~x304 & ~x310 & ~x335 & ~x336 & ~x337 & ~x361 & ~x391 & ~x423 & ~x447 & ~x477 & ~x478 & ~x534 & ~x557 & ~x559 & ~x587 & ~x618 & ~x672 & ~x697 & ~x698 & ~x699 & ~x701 & ~x726 & ~x728 & ~x729 & ~x740 & ~x746 & ~x769 & ~x783;
assign c4358 = ~x21 & ~x32 & ~x62 & ~x80 & ~x85 & ~x223 & ~x264 & ~x333 & ~x348 & ~x381 & ~x389 & ~x394 & ~x420 & ~x474 & ~x700;
assign c4360 =  x457 &  x577 &  x596 &  x600 & ~x2 & ~x5 & ~x6 & ~x8 & ~x9 & ~x18 & ~x19 & ~x21 & ~x26 & ~x28 & ~x29 & ~x30 & ~x32 & ~x49 & ~x50 & ~x51 & ~x52 & ~x53 & ~x57 & ~x58 & ~x60 & ~x61 & ~x63 & ~x78 & ~x81 & ~x83 & ~x84 & ~x85 & ~x87 & ~x108 & ~x111 & ~x114 & ~x116 & ~x135 & ~x137 & ~x141 & ~x163 & ~x164 & ~x168 & ~x169 & ~x170 & ~x171 & ~x172 & ~x196 & ~x197 & ~x220 & ~x222 & ~x224 & ~x227 & ~x248 & ~x252 & ~x253 & ~x276 & ~x277 & ~x278 & ~x281 & ~x282 & ~x304 & ~x307 & ~x334 & ~x362 & ~x363 & ~x364 & ~x366 & ~x389 & ~x392 & ~x394 & ~x421 & ~x444 & ~x447 & ~x448 & ~x450 & ~x451 & ~x502 & ~x503 & ~x504 & ~x528 & ~x530 & ~x532 & ~x557 & ~x558 & ~x559 & ~x561 & ~x587 & ~x588 & ~x613 & ~x616 & ~x642 & ~x644 & ~x645 & ~x669 & ~x670 & ~x674 & ~x702 & ~x727 & ~x729 & ~x754 & ~x755 & ~x758 & ~x759 & ~x764 & ~x766 & ~x769 & ~x770 & ~x772 & ~x773;
assign c4362 =  x40 &  x42 &  x630 & ~x7 & ~x24 & ~x26 & ~x36 & ~x51 & ~x55 & ~x79 & ~x82 & ~x86 & ~x106 & ~x115 & ~x137 & ~x166 & ~x168 & ~x196 & ~x199 & ~x250 & ~x252 & ~x363 & ~x364 & ~x365 & ~x448 & ~x477 & ~x502 & ~x504 & ~x588 & ~x720 & ~x739 & ~x740 & ~x745 & ~x747 & ~x757 & ~x775;
assign c4364 =  x43 &  x45 &  x180 &  x233 &  x272 &  x287 &  x327 &  x347 &  x351 &  x371 &  x375 &  x413 &  x519 &  x571 &  x576 &  x601 &  x635 &  x655 & ~x1 & ~x3 & ~x20 & ~x21 & ~x51 & ~x56 & ~x57 & ~x60 & ~x61 & ~x78 & ~x85 & ~x109 & ~x138 & ~x194 & ~x224 & ~x227 & ~x335 & ~x418 & ~x422 & ~x449 & ~x474 & ~x502 & ~x701 & ~x729 & ~x777 & ~x778;
assign c4366 = ~x0 & ~x4 & ~x7 & ~x8 & ~x19 & ~x21 & ~x23 & ~x28 & ~x29 & ~x30 & ~x31 & ~x32 & ~x51 & ~x54 & ~x55 & ~x56 & ~x78 & ~x109 & ~x111 & ~x115 & ~x116 & ~x135 & ~x138 & ~x140 & ~x141 & ~x143 & ~x166 & ~x194 & ~x220 & ~x227 & ~x249 & ~x252 & ~x253 & ~x255 & ~x264 & ~x281 & ~x304 & ~x309 & ~x335 & ~x338 & ~x366 & ~x389 & ~x422 & ~x445 & ~x448 & ~x449 & ~x473 & ~x488 & ~x505 & ~x506 & ~x529 & ~x531 & ~x532 & ~x533 & ~x534 & ~x557 & ~x559 & ~x562 & ~x614 & ~x671 & ~x698 & ~x700 & ~x725 & ~x727 & ~x728 & ~x756 & ~x765 & ~x783;
assign c4368 = ~x0 & ~x18 & ~x49 & ~x57 & ~x84 & ~x135 & ~x138 & ~x139 & ~x140 & ~x142 & ~x165 & ~x220 & ~x249 & ~x251 & ~x336 & ~x365 & ~x367 & ~x391 & ~x393 & ~x418 & ~x475 & ~x503 & ~x529 & ~x558 & ~x599 & ~x741 & ~x768;
assign c4370 =  x266 &  x323 &  x343 &  x441 &  x565 &  x610 &  x748 & ~x2 & ~x135 & ~x164 & ~x193 & ~x197 & ~x306 & ~x336 & ~x503 & ~x727;
assign c4372 =  x540 & ~x1 & ~x3 & ~x4 & ~x5 & ~x6 & ~x18 & ~x19 & ~x20 & ~x21 & ~x22 & ~x24 & ~x25 & ~x29 & ~x30 & ~x31 & ~x33 & ~x34 & ~x35 & ~x36 & ~x37 & ~x47 & ~x48 & ~x51 & ~x52 & ~x59 & ~x78 & ~x80 & ~x82 & ~x84 & ~x108 & ~x109 & ~x110 & ~x112 & ~x113 & ~x114 & ~x136 & ~x137 & ~x138 & ~x139 & ~x140 & ~x142 & ~x164 & ~x166 & ~x167 & ~x168 & ~x170 & ~x171 & ~x172 & ~x192 & ~x197 & ~x220 & ~x223 & ~x224 & ~x225 & ~x227 & ~x249 & ~x251 & ~x253 & ~x254 & ~x278 & ~x280 & ~x281 & ~x283 & ~x305 & ~x309 & ~x333 & ~x334 & ~x335 & ~x336 & ~x362 & ~x363 & ~x364 & ~x365 & ~x367 & ~x389 & ~x392 & ~x394 & ~x395 & ~x417 & ~x418 & ~x419 & ~x420 & ~x421 & ~x446 & ~x447 & ~x448 & ~x449 & ~x450 & ~x474 & ~x475 & ~x477 & ~x478 & ~x501 & ~x502 & ~x504 & ~x505 & ~x506 & ~x529 & ~x530 & ~x532 & ~x533 & ~x534 & ~x558 & ~x560 & ~x562 & ~x588 & ~x590 & ~x615 & ~x617 & ~x618 & ~x643 & ~x645 & ~x646 & ~x669 & ~x672 & ~x674 & ~x698 & ~x700 & ~x701 & ~x725 & ~x727 & ~x729 & ~x730 & ~x736 & ~x754 & ~x758 & ~x764 & ~x765 & ~x766 & ~x767 & ~x768 & ~x769 & ~x770 & ~x782 & ~x783;
assign c4374 =  x97 &  x287 &  x315 &  x384 &  x456 &  x468 &  x512 &  x538 &  x539 &  x552 &  x595 &  x651 & ~x1 & ~x6 & ~x9 & ~x23 & ~x33 & ~x52 & ~x57 & ~x61 & ~x77 & ~x81 & ~x82 & ~x90 & ~x107 & ~x113 & ~x114 & ~x135 & ~x136 & ~x137 & ~x138 & ~x143 & ~x168 & ~x169 & ~x192 & ~x194 & ~x195 & ~x196 & ~x225 & ~x226 & ~x249 & ~x250 & ~x253 & ~x276 & ~x277 & ~x278 & ~x280 & ~x281 & ~x334 & ~x339 & ~x363 & ~x388 & ~x390 & ~x392 & ~x418 & ~x419 & ~x448 & ~x474 & ~x529 & ~x615 & ~x644 & ~x697 & ~x702 & ~x726 & ~x727 & ~x764;
assign c4376 =  x15 &  x45 &  x127 &  x244 &  x269 &  x300 &  x348 &  x401 &  x465 &  x565 &  x622 &  x639 & ~x25 & ~x33 & ~x35 & ~x56 & ~x81 & ~x85 & ~x167 & ~x192 & ~x222 & ~x278 & ~x364 & ~x532 & ~x588 & ~x589 & ~x672 & ~x755;
assign c4378 =  x218 &  x413 &  x582 & ~x0 & ~x9 & ~x20 & ~x31 & ~x35 & ~x53 & ~x57 & ~x59 & ~x60 & ~x62 & ~x77 & ~x78 & ~x84 & ~x85 & ~x106 & ~x109 & ~x110 & ~x112 & ~x113 & ~x138 & ~x143 & ~x167 & ~x169 & ~x193 & ~x197 & ~x198 & ~x199 & ~x226 & ~x249 & ~x251 & ~x254 & ~x277 & ~x280 & ~x283 & ~x307 & ~x309 & ~x337 & ~x390 & ~x391 & ~x393 & ~x448 & ~x450 & ~x474 & ~x475 & ~x476 & ~x531 & ~x532 & ~x533 & ~x558 & ~x588 & ~x589 & ~x613 & ~x616 & ~x669 & ~x670 & ~x672 & ~x700 & ~x702 & ~x728 & ~x738 & ~x740 & ~x746 & ~x757 & ~x769 & ~x773;
assign c4380 =  x124 &  x185 &  x263 &  x299 &  x325 &  x353 &  x376 &  x402 &  x403 &  x409 &  x434 &  x489 &  x514 &  x546 &  x575 &  x632 &  x686 &  x688 &  x709 &  x717 & ~x3 & ~x7 & ~x8 & ~x10 & ~x30 & ~x31 & ~x48 & ~x50 & ~x51 & ~x54 & ~x62 & ~x220 & ~x224 & ~x248 & ~x254 & ~x277 & ~x281 & ~x284 & ~x310 & ~x340 & ~x366 & ~x368 & ~x395 & ~x452 & ~x476 & ~x591 & ~x642 & ~x670 & ~x727 & ~x728 & ~x734;
assign c4382 = ~x5 & ~x8 & ~x9 & ~x11 & ~x18 & ~x20 & ~x35 & ~x47 & ~x52 & ~x53 & ~x80 & ~x83 & ~x106 & ~x109 & ~x110 & ~x114 & ~x136 & ~x137 & ~x138 & ~x141 & ~x144 & ~x145 & ~x165 & ~x170 & ~x174 & ~x191 & ~x192 & ~x197 & ~x200 & ~x221 & ~x225 & ~x227 & ~x244 & ~x248 & ~x251 & ~x253 & ~x276 & ~x278 & ~x281 & ~x304 & ~x311 & ~x332 & ~x335 & ~x360 & ~x362 & ~x367 & ~x389 & ~x393 & ~x397 & ~x422 & ~x445 & ~x474 & ~x476 & ~x477 & ~x504 & ~x506 & ~x533 & ~x560 & ~x562 & ~x615 & ~x616 & ~x617 & ~x618 & ~x700 & ~x702 & ~x725 & ~x729 & ~x747 & ~x756 & ~x759 & ~x783;
assign c4384 =  x69 &  x591 & ~x30 & ~x78 & ~x86 & ~x106 & ~x194 & ~x249 & ~x336 & ~x560 & ~x615;
assign c4386 =  x455 &  x658 & ~x7 & ~x8 & ~x20 & ~x22 & ~x55 & ~x60 & ~x61 & ~x80 & ~x81 & ~x88 & ~x111 & ~x115 & ~x142 & ~x144 & ~x164 & ~x192 & ~x193 & ~x197 & ~x199 & ~x251 & ~x253 & ~x276 & ~x306 & ~x318 & ~x333 & ~x417 & ~x418 & ~x446 & ~x450 & ~x474 & ~x506 & ~x529 & ~x534 & ~x559 & ~x561 & ~x587 & ~x619 & ~x674 & ~x701 & ~x726 & ~x730 & ~x755 & ~x782;
assign c4388 =  x158 &  x245 &  x291 &  x500 &  x608 &  x629 & ~x165 & ~x252 & ~x336 & ~x392;
assign c4390 = ~x17 & ~x46 & ~x48 & ~x54 & ~x62 & ~x65 & ~x81 & ~x92 & ~x106 & ~x118 & ~x141 & ~x169 & ~x174 & ~x221 & ~x222 & ~x249 & ~x332 & ~x666 & ~x694 & ~x722;
assign c4392 =  x44 &  x185 &  x242 &  x261 &  x267 &  x345 &  x436 &  x462 &  x463 &  x466 &  x491 &  x493 &  x517 &  x547 &  x548 &  x575 &  x576 & ~x9 & ~x20 & ~x21 & ~x23 & ~x25 & ~x29 & ~x31 & ~x52 & ~x56 & ~x78 & ~x80 & ~x81 & ~x83 & ~x86 & ~x115 & ~x145 & ~x166 & ~x191 & ~x193 & ~x195 & ~x253 & ~x276 & ~x279 & ~x284 & ~x304 & ~x305 & ~x306 & ~x310 & ~x311 & ~x312 & ~x337 & ~x339 & ~x388 & ~x393 & ~x418 & ~x420 & ~x445 & ~x446 & ~x449 & ~x450 & ~x477 & ~x505 & ~x530 & ~x589 & ~x669 & ~x700 & ~x722 & ~x729 & ~x733 & ~x750 & ~x759 & ~x762 & ~x763 & ~x776;
assign c4394 =  x98 & ~x0 & ~x2 & ~x5 & ~x6 & ~x7 & ~x8 & ~x19 & ~x21 & ~x25 & ~x26 & ~x27 & ~x28 & ~x30 & ~x31 & ~x34 & ~x48 & ~x49 & ~x53 & ~x54 & ~x56 & ~x59 & ~x61 & ~x62 & ~x79 & ~x80 & ~x83 & ~x85 & ~x87 & ~x108 & ~x111 & ~x112 & ~x113 & ~x114 & ~x115 & ~x136 & ~x137 & ~x164 & ~x165 & ~x167 & ~x168 & ~x170 & ~x171 & ~x192 & ~x193 & ~x194 & ~x195 & ~x196 & ~x221 & ~x227 & ~x249 & ~x250 & ~x251 & ~x252 & ~x278 & ~x279 & ~x281 & ~x283 & ~x304 & ~x305 & ~x306 & ~x307 & ~x309 & ~x310 & ~x311 & ~x333 & ~x334 & ~x335 & ~x337 & ~x352 & ~x362 & ~x365 & ~x367 & ~x390 & ~x391 & ~x392 & ~x393 & ~x394 & ~x420 & ~x421 & ~x422 & ~x445 & ~x446 & ~x448 & ~x475 & ~x476 & ~x477 & ~x503 & ~x504 & ~x505 & ~x530 & ~x531 & ~x532 & ~x534 & ~x558 & ~x559 & ~x560 & ~x561 & ~x589 & ~x614 & ~x616 & ~x617 & ~x643 & ~x644 & ~x645 & ~x646 & ~x671 & ~x672 & ~x698 & ~x728 & ~x729 & ~x753 & ~x755 & ~x759 & ~x763 & ~x783;
assign c4396 = ~x25 & ~x27 & ~x49 & ~x51 & ~x90 & ~x133 & ~x145 & ~x146 & ~x198 & ~x253 & ~x308 & ~x394 & ~x419 & ~x477 & ~x493;
assign c4398 =  x333;
assign c4400 = ~x1 & ~x2 & ~x3 & ~x4 & ~x5 & ~x6 & ~x7 & ~x8 & ~x9 & ~x19 & ~x20 & ~x21 & ~x23 & ~x24 & ~x25 & ~x26 & ~x27 & ~x28 & ~x30 & ~x31 & ~x32 & ~x35 & ~x36 & ~x48 & ~x49 & ~x50 & ~x51 & ~x52 & ~x53 & ~x54 & ~x55 & ~x56 & ~x57 & ~x58 & ~x59 & ~x61 & ~x62 & ~x63 & ~x77 & ~x78 & ~x79 & ~x80 & ~x81 & ~x82 & ~x83 & ~x85 & ~x87 & ~x89 & ~x106 & ~x107 & ~x108 & ~x110 & ~x111 & ~x113 & ~x114 & ~x115 & ~x117 & ~x134 & ~x135 & ~x136 & ~x138 & ~x139 & ~x140 & ~x141 & ~x142 & ~x144 & ~x163 & ~x164 & ~x165 & ~x166 & ~x167 & ~x169 & ~x170 & ~x171 & ~x172 & ~x191 & ~x193 & ~x194 & ~x195 & ~x196 & ~x198 & ~x200 & ~x219 & ~x222 & ~x223 & ~x224 & ~x225 & ~x226 & ~x227 & ~x248 & ~x249 & ~x251 & ~x252 & ~x253 & ~x254 & ~x255 & ~x276 & ~x277 & ~x278 & ~x279 & ~x280 & ~x281 & ~x282 & ~x284 & ~x304 & ~x305 & ~x306 & ~x307 & ~x308 & ~x309 & ~x310 & ~x311 & ~x334 & ~x335 & ~x337 & ~x338 & ~x339 & ~x360 & ~x361 & ~x362 & ~x363 & ~x364 & ~x366 & ~x367 & ~x391 & ~x392 & ~x393 & ~x394 & ~x395 & ~x417 & ~x418 & ~x419 & ~x420 & ~x421 & ~x422 & ~x423 & ~x444 & ~x445 & ~x447 & ~x448 & ~x449 & ~x450 & ~x451 & ~x472 & ~x473 & ~x475 & ~x478 & ~x479 & ~x501 & ~x502 & ~x503 & ~x504 & ~x505 & ~x507 & ~x529 & ~x531 & ~x532 & ~x533 & ~x534 & ~x535 & ~x556 & ~x557 & ~x558 & ~x560 & ~x563 & ~x584 & ~x585 & ~x586 & ~x587 & ~x590 & ~x591 & ~x612 & ~x613 & ~x617 & ~x619 & ~x640 & ~x644 & ~x645 & ~x646 & ~x647 & ~x668 & ~x669 & ~x670 & ~x673 & ~x674 & ~x675 & ~x697 & ~x698 & ~x699 & ~x700 & ~x701 & ~x702 & ~x703 & ~x708 & ~x724 & ~x725 & ~x727 & ~x728 & ~x729 & ~x737 & ~x738 & ~x739 & ~x740 & ~x741 & ~x742 & ~x743 & ~x744 & ~x745 & ~x747 & ~x752 & ~x753 & ~x755 & ~x756 & ~x759 & ~x760 & ~x764 & ~x765 & ~x766 & ~x767 & ~x768 & ~x769 & ~x770 & ~x772 & ~x773 & ~x775 & ~x776 & ~x781 & ~x783;
assign c4402 = ~x6 & ~x7 & ~x10 & ~x20 & ~x21 & ~x23 & ~x30 & ~x32 & ~x34 & ~x48 & ~x49 & ~x52 & ~x53 & ~x55 & ~x79 & ~x81 & ~x86 & ~x87 & ~x107 & ~x109 & ~x115 & ~x137 & ~x144 & ~x169 & ~x170 & ~x192 & ~x193 & ~x195 & ~x199 & ~x248 & ~x250 & ~x251 & ~x254 & ~x277 & ~x282 & ~x308 & ~x334 & ~x338 & ~x339 & ~x361 & ~x362 & ~x364 & ~x389 & ~x393 & ~x418 & ~x419 & ~x422 & ~x448 & ~x474 & ~x505 & ~x529 & ~x534 & ~x561 & ~x597 & ~x615 & ~x671 & ~x674 & ~x728 & ~x755 & ~x757 & ~x764 & ~x765 & ~x767 & ~x769 & ~x770;
assign c4404 = ~x20 & ~x334 & ~x529 & ~x586 & ~x605 & ~x719 & ~x737 & ~x738 & ~x741;
assign c4406 =  x574 & ~x460;
assign c4408 =  x248;
assign c4410 =  x145 &  x490 &  x623 & ~x27 & ~x55 & ~x59 & ~x391 & ~x671;
assign c4412 =  x327 &  x355 & ~x4 & ~x6 & ~x10 & ~x20 & ~x46 & ~x54 & ~x55 & ~x80 & ~x85 & ~x163 & ~x166 & ~x254 & ~x274 & ~x303 & ~x306 & ~x420 & ~x448 & ~x559 & ~x585 & ~x586 & ~x588 & ~x615 & ~x666 & ~x672 & ~x677 & ~x693 & ~x695;
assign c4414 =  x385 &  x542 &  x577 &  x692 & ~x8 & ~x23 & ~x24 & ~x59 & ~x60 & ~x107 & ~x135 & ~x169 & ~x220 & ~x338 & ~x444 & ~x451 & ~x507 & ~x534 & ~x618 & ~x644 & ~x702 & ~x726 & ~x753;
assign c4416 =  x261 &  x262 &  x345 &  x411 &  x489 &  x629 &  x633 &  x687 & ~x5 & ~x7 & ~x18 & ~x80 & ~x112 & ~x142 & ~x164 & ~x192 & ~x219 & ~x222 & ~x224 & ~x275 & ~x283 & ~x304 & ~x364 & ~x446 & ~x448 & ~x500 & ~x501 & ~x560 & ~x587 & ~x615 & ~x644 & ~x645 & ~x697 & ~x721 & ~x776;
assign c4418 =  x69 &  x296 &  x355 &  x380 &  x384 &  x403 &  x412 &  x440 &  x466 &  x493 &  x517 &  x547 &  x573 & ~x7 & ~x19 & ~x25 & ~x26 & ~x53 & ~x57 & ~x80 & ~x86 & ~x87 & ~x111 & ~x112 & ~x113 & ~x115 & ~x116 & ~x140 & ~x142 & ~x171 & ~x198 & ~x222 & ~x247 & ~x248 & ~x253 & ~x256 & ~x282 & ~x305 & ~x310 & ~x312 & ~x340 & ~x360 & ~x367 & ~x388 & ~x389 & ~x393 & ~x418 & ~x420 & ~x476 & ~x500 & ~x505 & ~x590 & ~x614 & ~x671 & ~x674 & ~x700 & ~x704 & ~x729 & ~x734 & ~x749 & ~x750 & ~x757 & ~x760 & ~x762 & ~x778 & ~x779 & ~x780;
assign c4420 =  x596 & ~x0 & ~x1 & ~x3 & ~x6 & ~x25 & ~x31 & ~x52 & ~x58 & ~x59 & ~x80 & ~x82 & ~x85 & ~x86 & ~x111 & ~x112 & ~x137 & ~x141 & ~x163 & ~x166 & ~x169 & ~x171 & ~x194 & ~x221 & ~x251 & ~x277 & ~x279 & ~x282 & ~x283 & ~x305 & ~x309 & ~x335 & ~x367 & ~x420 & ~x421 & ~x445 & ~x446 & ~x473 & ~x474 & ~x475 & ~x477 & ~x521 & ~x560 & ~x642 & ~x644 & ~x645 & ~x670 & ~x698 & ~x700 & ~x702 & ~x729 & ~x782;
assign c4422 =  x289 &  x619 &  x675 &  x703 & ~x277;
assign c4424 =  x218 &  x257 &  x459 & ~x29 & ~x34 & ~x76 & ~x196 & ~x308 & ~x769;
assign c4426 = ~x1 & ~x2 & ~x3 & ~x5 & ~x6 & ~x7 & ~x8 & ~x19 & ~x20 & ~x23 & ~x25 & ~x26 & ~x27 & ~x29 & ~x30 & ~x31 & ~x32 & ~x33 & ~x34 & ~x49 & ~x50 & ~x52 & ~x53 & ~x55 & ~x57 & ~x58 & ~x59 & ~x60 & ~x61 & ~x78 & ~x79 & ~x81 & ~x82 & ~x84 & ~x85 & ~x87 & ~x88 & ~x106 & ~x107 & ~x108 & ~x109 & ~x110 & ~x112 & ~x115 & ~x135 & ~x137 & ~x138 & ~x139 & ~x141 & ~x142 & ~x144 & ~x164 & ~x165 & ~x166 & ~x167 & ~x169 & ~x170 & ~x171 & ~x193 & ~x194 & ~x195 & ~x196 & ~x197 & ~x198 & ~x199 & ~x220 & ~x222 & ~x223 & ~x224 & ~x225 & ~x249 & ~x250 & ~x251 & ~x252 & ~x253 & ~x254 & ~x267 & ~x277 & ~x278 & ~x279 & ~x280 & ~x281 & ~x282 & ~x283 & ~x305 & ~x307 & ~x308 & ~x309 & ~x334 & ~x335 & ~x336 & ~x337 & ~x338 & ~x339 & ~x362 & ~x363 & ~x364 & ~x365 & ~x366 & ~x367 & ~x389 & ~x390 & ~x392 & ~x394 & ~x418 & ~x419 & ~x420 & ~x421 & ~x422 & ~x445 & ~x448 & ~x449 & ~x450 & ~x474 & ~x475 & ~x476 & ~x477 & ~x478 & ~x502 & ~x503 & ~x504 & ~x505 & ~x530 & ~x531 & ~x532 & ~x559 & ~x561 & ~x586 & ~x587 & ~x588 & ~x590 & ~x615 & ~x617 & ~x618 & ~x642 & ~x643 & ~x644 & ~x645 & ~x646 & ~x670 & ~x672 & ~x698 & ~x699 & ~x701 & ~x702 & ~x726 & ~x727 & ~x728 & ~x729 & ~x741 & ~x755 & ~x757 & ~x758 & ~x764 & ~x765 & ~x769 & ~x773 & ~x774 & ~x775 & ~x776 & ~x782 & ~x783;
assign c4428 =  x697;
assign c4430 =  x270 &  x289 & ~x10 & ~x17 & ~x28 & ~x54 & ~x60 & ~x77 & ~x105 & ~x135 & ~x162 & ~x163 & ~x190 & ~x310 & ~x619 & ~x640 & ~x644 & ~x666 & ~x668 & ~x700 & ~x729 & ~x753 & ~x765 & ~x775;
assign c4432 =  x262 &  x270 &  x373 &  x411 &  x462 & ~x171 & ~x255 & ~x257 & ~x416 & ~x424 & ~x508 & ~x641 & ~x651 & ~x733 & ~x781;
assign c4434 =  x298 & ~x6 & ~x8 & ~x10 & ~x17 & ~x19 & ~x26 & ~x31 & ~x50 & ~x84 & ~x108 & ~x115 & ~x117 & ~x143 & ~x170 & ~x190 & ~x247 & ~x249 & ~x303 & ~x304 & ~x390 & ~x416 & ~x423 & ~x451 & ~x503 & ~x527 & ~x529 & ~x589 & ~x670 & ~x671 & ~x675 & ~x698 & ~x702 & ~x708 & ~x752 & ~x759 & ~x760 & ~x765;
assign c4436 =  x230 &  x424 &  x647 &  x675 & ~x27 & ~x29 & ~x31 & ~x32 & ~x49 & ~x53 & ~x56 & ~x60 & ~x62 & ~x78 & ~x109 & ~x111 & ~x113 & ~x136 & ~x168 & ~x193 & ~x222 & ~x223 & ~x250 & ~x251 & ~x279 & ~x280 & ~x337 & ~x419;
assign c4438 =  x557;
assign c4440 =  x103 &  x372 &  x408 &  x485 & ~x7 & ~x9 & ~x20 & ~x26 & ~x30 & ~x36 & ~x48 & ~x50 & ~x54 & ~x62 & ~x78 & ~x79 & ~x84 & ~x108 & ~x115 & ~x138 & ~x142 & ~x167 & ~x195 & ~x225 & ~x252 & ~x335 & ~x391 & ~x393 & ~x418 & ~x420 & ~x445 & ~x449 & ~x450 & ~x501 & ~x529 & ~x533 & ~x557 & ~x559 & ~x560 & ~x642 & ~x670 & ~x672 & ~x738 & ~x768 & ~x774;
assign c4442 =  x602 & ~x6 & ~x26 & ~x36 & ~x62 & ~x89 & ~x140 & ~x141 & ~x278 & ~x395 & ~x457 & ~x502 & ~x533 & ~x644 & ~x701;
assign c4444 =  x70 &  x71 &  x126 & ~x1 & ~x2 & ~x3 & ~x4 & ~x9 & ~x21 & ~x23 & ~x24 & ~x49 & ~x50 & ~x52 & ~x53 & ~x54 & ~x56 & ~x57 & ~x58 & ~x60 & ~x80 & ~x82 & ~x84 & ~x87 & ~x109 & ~x110 & ~x111 & ~x112 & ~x116 & ~x135 & ~x136 & ~x137 & ~x139 & ~x140 & ~x165 & ~x167 & ~x194 & ~x195 & ~x220 & ~x221 & ~x222 & ~x227 & ~x249 & ~x250 & ~x252 & ~x253 & ~x278 & ~x280 & ~x281 & ~x283 & ~x305 & ~x306 & ~x307 & ~x309 & ~x310 & ~x311 & ~x337 & ~x338 & ~x363 & ~x390 & ~x393 & ~x394 & ~x445 & ~x447 & ~x449 & ~x450 & ~x474 & ~x475 & ~x478 & ~x501 & ~x503 & ~x504 & ~x506 & ~x532 & ~x558 & ~x559 & ~x586 & ~x587 & ~x588 & ~x590 & ~x670 & ~x672 & ~x673 & ~x674 & ~x702 & ~x709 & ~x711 & ~x716 & ~x719 & ~x726 & ~x727 & ~x728 & ~x738 & ~x739 & ~x745 & ~x746 & ~x756 & ~x766 & ~x768 & ~x771 & ~x774 & ~x780;
assign c4446 =  x45 &  x180 &  x261 &  x272 &  x292 &  x295 &  x317 &  x321 &  x348 &  x464 &  x522 &  x547 &  x548 &  x599 &  x607 &  x632 &  x687 & ~x2 & ~x3 & ~x9 & ~x24 & ~x52 & ~x88 & ~x113 & ~x166 & ~x194 & ~x199 & ~x227 & ~x311 & ~x388 & ~x420 & ~x447 & ~x503 & ~x558 & ~x700 & ~x727 & ~x762 & ~x782;
assign c4448 = ~x3 & ~x4 & ~x6 & ~x8 & ~x9 & ~x10 & ~x18 & ~x19 & ~x20 & ~x21 & ~x22 & ~x23 & ~x24 & ~x25 & ~x26 & ~x27 & ~x28 & ~x29 & ~x30 & ~x31 & ~x32 & ~x33 & ~x34 & ~x48 & ~x49 & ~x50 & ~x51 & ~x52 & ~x53 & ~x56 & ~x58 & ~x59 & ~x61 & ~x77 & ~x78 & ~x79 & ~x80 & ~x81 & ~x84 & ~x85 & ~x87 & ~x88 & ~x107 & ~x108 & ~x110 & ~x113 & ~x114 & ~x116 & ~x117 & ~x138 & ~x139 & ~x140 & ~x142 & ~x143 & ~x144 & ~x163 & ~x164 & ~x167 & ~x168 & ~x169 & ~x170 & ~x171 & ~x172 & ~x193 & ~x195 & ~x196 & ~x200 & ~x220 & ~x222 & ~x223 & ~x224 & ~x227 & ~x228 & ~x248 & ~x250 & ~x251 & ~x252 & ~x276 & ~x277 & ~x278 & ~x280 & ~x281 & ~x283 & ~x304 & ~x305 & ~x306 & ~x307 & ~x308 & ~x309 & ~x311 & ~x333 & ~x334 & ~x336 & ~x338 & ~x339 & ~x361 & ~x362 & ~x364 & ~x389 & ~x390 & ~x391 & ~x392 & ~x393 & ~x394 & ~x395 & ~x418 & ~x422 & ~x423 & ~x446 & ~x447 & ~x448 & ~x449 & ~x450 & ~x451 & ~x473 & ~x474 & ~x478 & ~x486 & ~x503 & ~x507 & ~x529 & ~x530 & ~x531 & ~x533 & ~x534 & ~x535 & ~x558 & ~x559 & ~x560 & ~x561 & ~x562 & ~x586 & ~x588 & ~x589 & ~x614 & ~x615 & ~x642 & ~x643 & ~x644 & ~x645 & ~x646 & ~x670 & ~x673 & ~x698 & ~x699 & ~x700 & ~x702 & ~x727 & ~x728 & ~x729 & ~x755 & ~x756 & ~x758 & ~x760 & ~x783;
assign c4450 =  x484 & ~x1 & ~x115 & ~x390 & ~x392 & ~x627;
assign c4452 =  x180 &  x212 &  x275 &  x452 & ~x8 & ~x77;
assign c4454 =  x248;
assign c4456 =  x270 &  x317 &  x436 &  x459 &  x514 &  x518 &  x577 & ~x1 & ~x9 & ~x20 & ~x24 & ~x30 & ~x32 & ~x36 & ~x50 & ~x51 & ~x57 & ~x60 & ~x79 & ~x87 & ~x89 & ~x110 & ~x111 & ~x113 & ~x117 & ~x169 & ~x173 & ~x191 & ~x192 & ~x193 & ~x199 & ~x201 & ~x219 & ~x223 & ~x224 & ~x225 & ~x227 & ~x248 & ~x254 & ~x280 & ~x335 & ~x366 & ~x448 & ~x532 & ~x560 & ~x586 & ~x587 & ~x591 & ~x615 & ~x617 & ~x672 & ~x705 & ~x722 & ~x727 & ~x735 & ~x749 & ~x757 & ~x763 & ~x781;
assign c4458 =  x618;
assign c4460 =  x236 &  x240 &  x269 &  x289 &  x295 &  x344 &  x353 &  x376 &  x408 &  x437 &  x460 &  x482 &  x485 &  x493 &  x520 &  x538 &  x545 &  x549 &  x567 &  x569 &  x595 &  x596 &  x624 & ~x18 & ~x32 & ~x56 & ~x107 & ~x114 & ~x134 & ~x199 & ~x253 & ~x256 & ~x279 & ~x333 & ~x340 & ~x418 & ~x419 & ~x503 & ~x506 & ~x535 & ~x558 & ~x589 & ~x616 & ~x643 & ~x701 & ~x726 & ~x754 & ~x758 & ~x759;
assign c4462 =  x129 &  x318 &  x547 &  x575 & ~x84 & ~x142 & ~x311 & ~x389 & ~x446 & ~x449 & ~x642 & ~x711;
assign c4464 =  x45 &  x234 &  x292 &  x443 &  x466 &  x518 & ~x2 & ~x20 & ~x52 & ~x63 & ~x79 & ~x137 & ~x144 & ~x220 & ~x226 & ~x281 & ~x306 & ~x311 & ~x336 & ~x366 & ~x503 & ~x587;
assign c4466 =  x70 & ~x2 & ~x3 & ~x6 & ~x17 & ~x18 & ~x20 & ~x23 & ~x25 & ~x28 & ~x29 & ~x33 & ~x34 & ~x35 & ~x51 & ~x52 & ~x59 & ~x79 & ~x82 & ~x84 & ~x87 & ~x107 & ~x111 & ~x113 & ~x114 & ~x115 & ~x116 & ~x137 & ~x143 & ~x163 & ~x169 & ~x219 & ~x221 & ~x223 & ~x225 & ~x251 & ~x253 & ~x276 & ~x277 & ~x278 & ~x280 & ~x281 & ~x283 & ~x334 & ~x367 & ~x390 & ~x391 & ~x394 & ~x421 & ~x448 & ~x475 & ~x476 & ~x477 & ~x502 & ~x503 & ~x534 & ~x561 & ~x562 & ~x586 & ~x587 & ~x588 & ~x589 & ~x590 & ~x614 & ~x617 & ~x642 & ~x645 & ~x646 & ~x671 & ~x690 & ~x700 & ~x709 & ~x711 & ~x719 & ~x727 & ~x729 & ~x737 & ~x738 & ~x741 & ~x746 & ~x754 & ~x756 & ~x758 & ~x776 & ~x782;
assign c4468 =  x72 &  x285 &  x341 &  x539 & ~x0 & ~x58 & ~x167 & ~x199 & ~x249 & ~x250 & ~x418 & ~x445 & ~x618 & ~x672 & ~x674;
assign c4470 = ~x4 & ~x5 & ~x23 & ~x62 & ~x81 & ~x87 & ~x108 & ~x138 & ~x140 & ~x142 & ~x168 & ~x192 & ~x194 & ~x195 & ~x222 & ~x262 & ~x264 & ~x282 & ~x308 & ~x339 & ~x348 & ~x365 & ~x421 & ~x493 & ~x502 & ~x530;
assign c4472 = ~x2 & ~x3 & ~x8 & ~x9 & ~x10 & ~x17 & ~x18 & ~x20 & ~x21 & ~x23 & ~x24 & ~x26 & ~x34 & ~x35 & ~x49 & ~x51 & ~x52 & ~x53 & ~x54 & ~x56 & ~x60 & ~x79 & ~x80 & ~x81 & ~x82 & ~x83 & ~x85 & ~x86 & ~x87 & ~x107 & ~x110 & ~x111 & ~x112 & ~x113 & ~x114 & ~x115 & ~x139 & ~x141 & ~x142 & ~x168 & ~x193 & ~x194 & ~x195 & ~x196 & ~x200 & ~x225 & ~x250 & ~x277 & ~x280 & ~x282 & ~x283 & ~x305 & ~x310 & ~x335 & ~x337 & ~x362 & ~x363 & ~x418 & ~x420 & ~x421 & ~x448 & ~x474 & ~x477 & ~x530 & ~x531 & ~x557 & ~x559 & ~x561 & ~x576 & ~x616 & ~x617 & ~x643 & ~x645 & ~x669 & ~x670 & ~x674 & ~x700 & ~x702 & ~x725 & ~x728 & ~x729 & ~x759;
assign c4474 = ~x575;
assign c4476 =  x41 &  x45 &  x67 &  x95 &  x536 & ~x25 & ~x32 & ~x54 & ~x86 & ~x88 & ~x108 & ~x111 & ~x113 & ~x136 & ~x171 & ~x224 & ~x250 & ~x252 & ~x278 & ~x281 & ~x363 & ~x366 & ~x420 & ~x587 & ~x778;
assign c4478 =  x70 & ~x3 & ~x6 & ~x8 & ~x52 & ~x100 & ~x115 & ~x136 & ~x137 & ~x163 & ~x167 & ~x169 & ~x171 & ~x193 & ~x197 & ~x199 & ~x223 & ~x248 & ~x251 & ~x254 & ~x283 & ~x307 & ~x336 & ~x393 & ~x394 & ~x418 & ~x451 & ~x478 & ~x502 & ~x531 & ~x562 & ~x589 & ~x590 & ~x616 & ~x645 & ~x646 & ~x700 & ~x702 & ~x703;
assign c4480 =  x551 & ~x27 & ~x30 & ~x48 & ~x53 & ~x56 & ~x85 & ~x106 & ~x112 & ~x139 & ~x143 & ~x164 & ~x165 & ~x167 & ~x168 & ~x220 & ~x248 & ~x249 & ~x252 & ~x276 & ~x309 & ~x336 & ~x365 & ~x503 & ~x606 & ~x643 & ~x758;
assign c4482 =  x12 &  x41 &  x585;
assign c4484 =  x423;
assign c4486 = ~x3 & ~x6 & ~x8 & ~x9 & ~x18 & ~x20 & ~x21 & ~x22 & ~x24 & ~x26 & ~x27 & ~x29 & ~x30 & ~x31 & ~x32 & ~x36 & ~x49 & ~x50 & ~x55 & ~x57 & ~x59 & ~x60 & ~x75 & ~x81 & ~x82 & ~x86 & ~x106 & ~x108 & ~x109 & ~x113 & ~x115 & ~x116 & ~x117 & ~x137 & ~x138 & ~x139 & ~x143 & ~x165 & ~x166 & ~x167 & ~x168 & ~x169 & ~x171 & ~x172 & ~x191 & ~x192 & ~x193 & ~x194 & ~x200 & ~x222 & ~x225 & ~x226 & ~x227 & ~x249 & ~x250 & ~x251 & ~x252 & ~x276 & ~x277 & ~x278 & ~x282 & ~x304 & ~x307 & ~x308 & ~x309 & ~x311 & ~x332 & ~x333 & ~x336 & ~x338 & ~x339 & ~x361 & ~x362 & ~x363 & ~x364 & ~x366 & ~x367 & ~x389 & ~x395 & ~x417 & ~x418 & ~x421 & ~x423 & ~x446 & ~x449 & ~x451 & ~x473 & ~x474 & ~x475 & ~x502 & ~x503 & ~x506 & ~x530 & ~x531 & ~x534 & ~x558 & ~x560 & ~x561 & ~x562 & ~x585 & ~x586 & ~x587 & ~x588 & ~x589 & ~x613 & ~x617 & ~x642 & ~x670 & ~x671 & ~x672 & ~x698 & ~x702 & ~x703 & ~x709 & ~x725 & ~x726 & ~x728 & ~x729 & ~x730 & ~x738 & ~x741 & ~x754 & ~x755 & ~x757 & ~x764 & ~x765 & ~x766 & ~x768 & ~x773 & ~x775 & ~x776;
assign c4488 =  x219 &  x258 &  x582 & ~x30 & ~x107 & ~x141 & ~x199 & ~x250 & ~x253 & ~x309 & ~x391 & ~x392 & ~x475 & ~x558 & ~x699 & ~x728 & ~x755 & ~x770;
assign c4490 =  x236 &  x287 &  x288 &  x315 &  x321 &  x346 &  x384 &  x430 &  x433 &  x435 &  x498 &  x540 &  x544 &  x573 &  x578 &  x604 &  x628 &  x639 &  x650 &  x651 &  x652 &  x653 &  x688 & ~x1 & ~x31 & ~x51 & ~x53 & ~x112 & ~x117 & ~x142 & ~x169 & ~x248 & ~x251 & ~x304 & ~x309 & ~x337 & ~x338 & ~x366 & ~x393 & ~x419 & ~x447 & ~x476 & ~x531 & ~x701;
assign c4492 = ~x231 & ~x320;
assign c4494 =  x126 &  x353 &  x359 &  x469 & ~x0 & ~x3 & ~x4 & ~x7 & ~x19 & ~x20 & ~x24 & ~x26 & ~x33 & ~x53 & ~x55 & ~x59 & ~x83 & ~x107 & ~x108 & ~x111 & ~x137 & ~x143 & ~x170 & ~x199 & ~x221 & ~x225 & ~x227 & ~x249 & ~x252 & ~x254 & ~x278 & ~x282 & ~x306 & ~x307 & ~x310 & ~x335 & ~x337 & ~x338 & ~x365 & ~x446 & ~x448 & ~x502 & ~x504 & ~x533 & ~x558 & ~x559 & ~x560 & ~x586 & ~x588 & ~x615 & ~x616 & ~x617 & ~x642 & ~x645 & ~x672 & ~x687 & ~x700 & ~x727 & ~x756 & ~x757 & ~x767 & ~x783;
assign c4496 =  x413 & ~x34 & ~x351 & ~x726;
assign c4498 =  x177 &  x214 &  x359 &  x639 & ~x10 & ~x63 & ~x78 & ~x197 & ~x220 & ~x221 & ~x223 & ~x225 & ~x252 & ~x335 & ~x392 & ~x753;
assign c41 =  x86;
assign c43 =  x249;
assign c45 = ~x544 & ~x688;
assign c47 =  x95 &  x97 &  x98 &  x101 &  x130 &  x149 &  x150 &  x158 &  x159 &  x177 &  x178 &  x184 &  x212 &  x214 &  x319 &  x324 &  x325 &  x351 &  x377 &  x378 &  x382 &  x406 &  x430 &  x464 &  x494 &  x495 &  x518 &  x541 &  x597 &  x600 &  x602 &  x604 &  x606 &  x630 & ~x14 & ~x24 & ~x31 & ~x51 & ~x61 & ~x78 & ~x87 & ~x88 & ~x109 & ~x111 & ~x113 & ~x139 & ~x140 & ~x165 & ~x166 & ~x168 & ~x171 & ~x193 & ~x199 & ~x226 & ~x248 & ~x256 & ~x304 & ~x306 & ~x307 & ~x333 & ~x335 & ~x360 & ~x361 & ~x366 & ~x367 & ~x389 & ~x420 & ~x423 & ~x445 & ~x446 & ~x450 & ~x477 & ~x557 & ~x558 & ~x618 & ~x642 & ~x670 & ~x673 & ~x729 & ~x757 & ~x781 & ~x782;
assign c49 =  x54;
assign c411 =  x44 &  x45 &  x207 & ~x136 & ~x193 & ~x366 & ~x369 & ~x425 & ~x443 & ~x565 & ~x649 & ~x761;
assign c415 = ~x66 & ~x176;
assign c417 =  x46 &  x74 &  x94 &  x121 &  x126 &  x156 &  x158 &  x208 &  x239 &  x263 &  x292 &  x294 &  x376 &  x430 &  x432 & ~x13 & ~x778;
assign c419 =  x502;
assign c421 =  x419;
assign c423 =  x390;
assign c425 =  x1;
assign c429 =  x774 & ~x565;
assign c431 = ~x126 & ~x240;
assign c433 = ~x125 & ~x126;
assign c435 = ~x355 & ~x411 & ~x696 & ~x751;
assign c437 =  x212 & ~x525;
assign c439 =  x77;
assign c441 = ~x125;
assign c443 =  x57;
assign c445 =  x153 &  x180 &  x348 & ~x217 & ~x454 & ~x704;
assign c447 =  x101 &  x132 &  x182 &  x320 &  x522 &  x573 &  x600 &  x626 & ~x4 & ~x13 & ~x22 & ~x50 & ~x51 & ~x80 & ~x116 & ~x193 & ~x197 & ~x223 & ~x227 & ~x305 & ~x366 & ~x417 & ~x450 & ~x504 & ~x505 & ~x531 & ~x586 & ~x703 & ~x731 & ~x757 & ~x780;
assign c449 =  x135;
assign c451 =  x114;
assign c453 =  x24;
assign c455 =  x309;
assign c457 =  x125 &  x177 &  x183 &  x235 &  x240 &  x291 &  x325 &  x438 &  x520 &  x578 &  x653 &  x710 &  x738 &  x742 & ~x2 & ~x53 & ~x140 & ~x248 & ~x256 & ~x278 & ~x531 & ~x533 & ~x536 & ~x556 & ~x564 & ~x583 & ~x613 & ~x616 & ~x701 & ~x751;
assign c459 = ~x398 & ~x428;
assign c461 =  x46 &  x208 &  x210 &  x212 &  x264 & ~x369;
assign c463 =  x7;
assign c465 =  x109;
assign c467 =  x250;
assign c469 =  x475;
assign c471 = ~x129 & ~x607;
assign c473 =  x196;
assign c475 = ~x572;
assign c477 =  x111;
assign c479 =  x1;
assign c481 =  x67 &  x73 &  x74 &  x92 &  x98 &  x104 &  x120 &  x129 &  x148 &  x154 &  x157 &  x182 &  x186 &  x188 &  x233 &  x259 &  x296 &  x301 &  x315 &  x323 &  x352 &  x369 &  x373 &  x381 &  x397 &  x407 &  x438 &  x457 &  x459 &  x489 &  x492 &  x493 &  x495 &  x510 &  x526 &  x542 &  x546 &  x571 &  x573 &  x574 &  x579 &  x593 &  x598 &  x599 &  x601 &  x621 &  x625 &  x627 &  x628 &  x630 &  x631 &  x639 &  x658 &  x660 &  x662 &  x676 &  x695 & ~x19 & ~x21 & ~x34 & ~x35 & ~x50 & ~x56 & ~x58 & ~x88 & ~x112 & ~x116 & ~x137 & ~x139 & ~x165 & ~x197 & ~x250 & ~x277 & ~x281 & ~x305 & ~x307 & ~x311 & ~x360 & ~x366 & ~x417 & ~x420 & ~x587 & ~x589 & ~x617 & ~x701 & ~x729 & ~x757 & ~x758 & ~x776;
assign c483 =  x62;
assign c485 = ~x95;
assign c487 =  x105 &  x118 &  x155 &  x230 &  x244 &  x549 &  x649 & ~x13 & ~x249;
assign c489 =  x531;
assign c491 =  x77 & ~x749;
assign c495 = ~x513 & ~x636;
assign c497 = ~x153 & ~x154 & ~x182;
assign c499 =  x118 &  x243 &  x627 &  x631 &  x653 &  x677 & ~x3 & ~x110 & ~x361 & ~x367 & ~x478 & ~x507 & ~x563 & ~x735;
assign c4101 = ~x327 & ~x411 & ~x664;
assign c4103 =  x195 &  x476;
assign c4105 =  x118 &  x201 &  x625 & ~x224 & ~x361 & ~x366 & ~x417 & ~x445 & ~x449 & ~x567 & ~x589;
assign c4107 = ~x544 & ~x602;
assign c4109 =  x70 &  x91 &  x100 &  x101 &  x104 &  x125 &  x126 &  x133 &  x146 &  x178 &  x188 &  x230 &  x234 &  x274 &  x287 &  x289 &  x348 &  x374 &  x376 &  x378 &  x487 &  x497 &  x601 &  x633 &  x635 &  x657 &  x711 &  x714 & ~x7 & ~x51 & ~x112 & ~x417 & ~x531 & ~x532 & ~x560 & ~x586 & ~x757 & ~x758 & ~x775 & ~x777;
assign c4111 =  x251;
assign c4113 =  x20;
assign c4115 =  x90 &  x106 &  x133 &  x498;
assign c4117 = ~x400 & ~x454;
assign c4119 =  x86;
assign c4121 =  x53;
assign c4123 =  x672;
assign c4125 = ~x343 & ~x398;
assign c4127 =  x21;
assign c4129 =  x142;
assign c4131 =  x504;
assign c4135 = ~x372 & ~x440;
assign c4137 = ~x153;
assign c4139 = ~x66 & ~x98 & ~x153;
assign c4141 =  x737 & ~x565;
assign c4143 = ~x65 & ~x239;
assign c4145 =  x165;
assign c4147 = ~x342 & ~x483 & ~x511 & ~x762;
assign c4149 =  x46 &  x95 &  x102 &  x156 & ~x6 & ~x14 & ~x15 & ~x116 & ~x283 & ~x417 & ~x702;
assign c4151 =  x447;
assign c4153 = ~x440 & ~x650;
assign c4155 =  x102 &  x103 &  x203 &  x244 &  x245 &  x601 &  x657 & ~x38 & ~x46 & ~x109 & ~x366 & ~x389 & ~x702 & ~x748 & ~x764;
assign c4157 =  x587;
assign c4159 =  x337;
assign c4161 =  x166;
assign c4163 =  x532;
assign c4167 =  x142;
assign c4169 =  x225;
assign c4173 =  x291 &  x464 &  x711 & ~x231 & ~x413;
assign c4175 =  x70 &  x101 & ~x484 & ~x512 & ~x556 & ~x640 & ~x724;
assign c4177 =  x67 &  x103 &  x129 &  x148 &  x160 &  x211 &  x244 &  x291 &  x346 &  x569 &  x625 &  x681 & ~x38 & ~x643 & ~x757 & ~x775;
assign c4179 =  x164;
assign c4181 =  x522 &  x747 & ~x245 & ~x274;
assign c4183 =  x65 &  x68 &  x69 &  x71 &  x91 &  x92 &  x97 &  x101 &  x103 &  x120 &  x124 &  x126 &  x127 &  x133 &  x146 &  x152 &  x158 &  x159 &  x174 &  x177 &  x187 &  x205 &  x210 &  x214 &  x216 &  x218 &  x236 &  x246 &  x266 &  x270 &  x274 &  x294 &  x299 &  x300 &  x302 &  x315 &  x322 &  x323 &  x324 &  x325 &  x342 &  x343 &  x345 &  x346 &  x347 &  x348 &  x376 &  x377 &  x382 &  x386 &  x405 &  x406 &  x407 &  x410 &  x411 &  x413 &  x414 &  x430 &  x438 &  x441 &  x458 &  x460 &  x463 &  x466 &  x471 &  x481 &  x492 &  x493 &  x494 &  x514 &  x515 &  x516 &  x525 &  x527 &  x541 &  x548 &  x565 &  x566 &  x569 &  x571 &  x573 &  x638 &  x660 &  x661 &  x666 & ~x3 & ~x5 & ~x8 & ~x22 & ~x24 & ~x28 & ~x33 & ~x34 & ~x49 & ~x57 & ~x59 & ~x61 & ~x83 & ~x84 & ~x108 & ~x138 & ~x139 & ~x143 & ~x164 & ~x171 & ~x195 & ~x197 & ~x223 & ~x225 & ~x249 & ~x252 & ~x283 & ~x305 & ~x309 & ~x334 & ~x336 & ~x361 & ~x363 & ~x364 & ~x390 & ~x420 & ~x422 & ~x445 & ~x447 & ~x477 & ~x501 & ~x530 & ~x531 & ~x534 & ~x588 & ~x669 & ~x672 & ~x702 & ~x755 & ~x758 & ~x776;
assign c4185 =  x107;
assign c4189 =  x166;
assign c4191 =  x67 &  x69 &  x92 &  x96 &  x101 &  x119 &  x120 &  x122 &  x124 &  x128 &  x129 &  x131 &  x146 &  x149 &  x151 &  x161 &  x174 &  x186 &  x209 &  x213 &  x216 &  x231 &  x236 &  x242 &  x244 &  x259 &  x266 &  x267 &  x270 &  x272 &  x285 &  x286 &  x293 &  x300 &  x314 &  x315 &  x320 &  x324 &  x342 &  x347 &  x352 &  x354 &  x369 &  x373 &  x382 &  x397 &  x402 &  x406 &  x409 &  x426 &  x429 &  x454 &  x461 &  x467 &  x498 &  x515 &  x516 &  x527 &  x536 &  x555 &  x564 &  x594 &  x603 &  x622 &  x627 &  x628 &  x631 &  x649 &  x652 &  x656 &  x661 &  x677 & ~x1 & ~x21 & ~x29 & ~x30 & ~x32 & ~x33 & ~x54 & ~x60 & ~x81 & ~x82 & ~x109 & ~x110 & ~x111 & ~x112 & ~x114 & ~x137 & ~x140 & ~x141 & ~x167 & ~x171 & ~x195 & ~x198 & ~x220 & ~x221 & ~x249 & ~x254 & ~x277 & ~x333 & ~x335 & ~x360 & ~x390 & ~x392 & ~x395 & ~x473 & ~x501 & ~x503 & ~x586 & ~x618 & ~x670 & ~x726 & ~x729 & ~x730 & ~x754 & ~x757 & ~x763;
assign c4193 = ~x97 & ~x98 & ~x99;
assign c4195 = ~x495 & ~x572;
assign c4197 = ~x65 & ~x149;
assign c4199 =  x222;
assign c4201 =  x30;
assign c4203 =  x10 &  x97 &  x150 &  x183 & ~x556 & ~x613 & ~x641 & ~x780;
assign c4205 = ~x12 & ~x42;
assign c4207 =  x79;
assign c4209 =  x109;
assign c4211 =  x69 &  x73 &  x75 &  x91 &  x93 &  x97 &  x105 &  x151 &  x154 &  x174 &  x175 & ~x13 & ~x82 & ~x168 & ~x249 & ~x333 & ~x757;
assign c4213 =  x65 &  x66 &  x73 &  x75 &  x94 &  x95 &  x100 &  x103 &  x126 &  x127 &  x131 &  x152 &  x158 &  x179 &  x183 &  x186 &  x213 &  x267 &  x322 &  x325 &  x350 &  x430 &  x432 &  x493 &  x519 &  x521 &  x598 &  x604 &  x628 &  x631 & ~x14 & ~x21 & ~x27 & ~x30 & ~x57 & ~x60 & ~x61 & ~x80 & ~x86 & ~x135 & ~x137 & ~x140 & ~x170 & ~x197 & ~x226 & ~x255 & ~x306 & ~x334 & ~x338 & ~x361 & ~x363 & ~x364 & ~x389 & ~x393 & ~x394 & ~x418 & ~x446 & ~x502 & ~x532 & ~x560 & ~x618 & ~x645 & ~x671 & ~x728 & ~x754 & ~x755 & ~x756 & ~x757 & ~x781;
assign c4215 = ~x70 & ~x99;
assign c4217 =  x23;
assign c4219 =  x73 &  x97 &  x102 &  x105 &  x121 &  x128 &  x134 &  x146 &  x162 &  x174 &  x240 &  x247 &  x289 &  x346 &  x377 &  x407 &  x523 &  x547 &  x549 &  x579 &  x603 &  x604 &  x626 &  x630 &  x632 &  x657 &  x683 &  x713 &  x715 &  x716 &  x718 & ~x50 & ~x51 & ~x170 & ~x221 & ~x253 & ~x277 & ~x278 & ~x282 & ~x306 & ~x365 & ~x392 & ~x615;
assign c4221 =  x78;
assign c4223 =  x69 &  x73 &  x74 &  x75 &  x92 &  x103 &  x120 &  x130 &  x176 &  x382 &  x466 &  x521 & ~x5 & ~x12 & ~x13 & ~x14 & ~x15 & ~x30 & ~x58 & ~x108 & ~x138 & ~x277 & ~x282 & ~x390 & ~x393 & ~x421;
assign c4225 = ~x356 & ~x440 & ~x511;
assign c4227 =  x134 &  x190 &  x740 &  x741 & ~x731;
assign c4229 =  x291 & ~x358;
assign c4231 =  x362;
assign c4233 =  x336;
assign c4235 =  x193;
assign c4237 = ~x74 & ~x154;
assign c4239 =  x417;
assign c4241 =  x153 &  x295 &  x541 & ~x23 & ~x114 & ~x305 & ~x308 & ~x609 & ~x731;
assign c4243 =  x107;
assign c4245 =  x165;
assign c4247 =  x108;
assign c4249 =  x252;
assign c4251 = ~x126 & ~x151 & ~x182;
assign c4253 =  x65 &  x73 &  x103 &  x119 &  x126 &  x150 &  x159 &  x160 &  x177 &  x179 &  x203 &  x206 &  x213 &  x214 &  x217 &  x261 &  x268 &  x270 &  x273 &  x293 &  x297 &  x298 &  x320 &  x342 &  x351 &  x353 &  x377 &  x516 &  x540 &  x598 &  x603 &  x605 &  x629 &  x653 &  x660 &  x661 & ~x24 & ~x26 & ~x27 & ~x30 & ~x50 & ~x52 & ~x58 & ~x61 & ~x112 & ~x135 & ~x137 & ~x163 & ~x168 & ~x221 & ~x223 & ~x252 & ~x335 & ~x339 & ~x367 & ~x392 & ~x393 & ~x418 & ~x421 & ~x422 & ~x448 & ~x449 & ~x477 & ~x530 & ~x586 & ~x589 & ~x615 & ~x618 & ~x643 & ~x729 & ~x748 & ~x756 & ~x763 & ~x776 & ~x783;
assign c4255 = ~x489;
assign c4257 = ~x440 & ~x468 & ~x469;
assign c4259 =  x475;
assign c4261 =  x249;
assign c4263 =  x588;
assign c4265 =  x250;
assign c4267 =  x81;
assign c4269 =  x28;
assign c4271 =  x112;
assign c4273 =  x24;
assign c4275 =  x281;
assign c4277 =  x20;
assign c4279 =  x84;
assign c4281 =  x44 &  x68 &  x74 &  x92 &  x94 &  x95 &  x96 &  x98 &  x104 &  x127 &  x133 &  x157 &  x178 &  x181 &  x182 &  x218 &  x232 &  x266 &  x273 &  x352 &  x382 &  x386 &  x431 &  x437 &  x442 &  x443 &  x461 &  x471 &  x498 &  x499 &  x523 &  x549 &  x555 &  x565 &  x632 &  x658 &  x663 & ~x22 & ~x25 & ~x32 & ~x51 & ~x55 & ~x59 & ~x82 & ~x108 & ~x139 & ~x171 & ~x199 & ~x223 & ~x224 & ~x255 & ~x279 & ~x333 & ~x361 & ~x476 & ~x531 & ~x728 & ~x757 & ~x762 & ~x775;
assign c4283 = ~x120 & ~x126;
assign c4285 = ~x546;
assign c4287 =  x80;
assign c4289 =  x281;
assign c4291 =  x617;
assign c4293 =  x365;
assign c4295 =  x66 &  x73 &  x74 &  x91 &  x97 &  x98 &  x104 &  x123 &  x157 &  x162 &  x183 &  x188 &  x203 &  x206 &  x211 &  x212 &  x213 &  x218 &  x238 &  x239 &  x245 &  x260 &  x315 &  x323 &  x329 &  x397 &  x406 &  x408 &  x425 &  x436 &  x453 &  x463 &  x469 &  x480 &  x495 &  x499 &  x508 &  x538 &  x544 &  x553 &  x554 &  x572 &  x577 &  x597 &  x604 &  x630 &  x658 &  x662 &  x691 & ~x29 & ~x32 & ~x53 & ~x87 & ~x111 & ~x113 & ~x114 & ~x139 & ~x223 & ~x225 & ~x249 & ~x251 & ~x307 & ~x334 & ~x363 & ~x366 & ~x390 & ~x445 & ~x476 & ~x560 & ~x588 & ~x589 & ~x644 & ~x672 & ~x727 & ~x755;
assign c4297 =  x783;
assign c4299 =  x66 &  x105 &  x119 &  x161 &  x354 &  x481 &  x490 & ~x13 & ~x227;
assign c4301 =  x64 &  x69 &  x76 &  x102 &  x105 &  x123 &  x126 &  x216 &  x236 &  x246 &  x350 &  x379 &  x414 &  x426 &  x628 &  x635 & ~x3 & ~x4 & ~x84 & ~x361 & ~x772 & ~x774;
assign c4303 =  x419;
assign c4305 =  x110 &  x163;
assign c4307 =  x364;
assign c4309 =  x62;
assign c4311 = ~x440 & ~x733;
assign c4313 =  x334;
assign c4315 =  x197;
assign c4317 =  x122 &  x129 &  x158 &  x541 &  x599 &  x740 &  x743 & ~x49 & ~x558 & ~x583 & ~x638;
assign c4319 = ~x126 & ~x182 & ~x214;
assign c4321 =  x39 &  x64 &  x90 &  x102 &  x104 &  x105 &  x119 &  x120 &  x132 &  x133 &  x204 &  x218 &  x232 &  x321 &  x374 &  x426 &  x488 &  x625 &  x631 &  x635 &  x655 &  x656 &  x658 & ~x2 & ~x4 & ~x87 & ~x111 & ~x195 & ~x220 & ~x282 & ~x333 & ~x449 & ~x477 & ~x534 & ~x559 & ~x586 & ~x727 & ~x763;
assign c4323 =  x587;
assign c4325 =  x67 &  x147 &  x177 &  x185 &  x186 &  x203 &  x214 &  x237 &  x260 &  x264 &  x270 &  x316 &  x351 &  x404 &  x407 &  x430 &  x455 &  x457 &  x483 &  x492 &  x494 &  x511 &  x525 &  x539 &  x594 &  x638 &  x710 &  x750 & ~x77 & ~x250 & ~x252 & ~x563 & ~x754 & ~x760;
assign c4327 =  x20;
assign c4329 =  x197;
assign c4331 =  x95 &  x155 &  x184 &  x208 & ~x538 & ~x583 & ~x704 & ~x754 & ~x762;
assign c4333 = ~x426 & ~x455;
assign c4337 =  x47 &  x117;
assign c4339 =  x727;
assign c4341 =  x59;
assign c4343 =  x135;
assign c4345 =  x57;
assign c4349 = ~x497;
assign c4351 =  x56;
assign c4353 = ~x343 & ~x356;
assign c4355 =  x116;
assign c4357 =  x138;
assign c4359 =  x25;
assign c4361 =  x305;
assign c4363 =  x79;
assign c4365 =  x587;
assign c4367 = ~x98;
assign c4369 =  x34;
assign c4371 =  x75 &  x95 &  x96 &  x97 &  x101 &  x102 &  x105 &  x122 &  x126 &  x146 &  x147 &  x152 &  x154 &  x158 &  x160 &  x176 &  x179 &  x186 &  x187 &  x189 &  x203 &  x204 &  x205 &  x206 &  x208 &  x211 &  x213 &  x217 &  x237 &  x243 &  x285 &  x296 &  x297 &  x298 &  x315 &  x318 &  x326 &  x348 &  x382 &  x425 &  x453 &  x463 &  x469 &  x481 &  x492 &  x493 &  x509 &  x525 &  x544 &  x565 &  x593 &  x598 &  x601 &  x604 &  x628 &  x630 &  x634 &  x635 &  x677 & ~x1 & ~x20 & ~x31 & ~x33 & ~x34 & ~x50 & ~x79 & ~x84 & ~x85 & ~x108 & ~x113 & ~x139 & ~x143 & ~x164 & ~x167 & ~x192 & ~x194 & ~x199 & ~x250 & ~x276 & ~x304 & ~x305 & ~x336 & ~x389 & ~x419 & ~x422 & ~x474 & ~x504 & ~x589 & ~x615 & ~x644 & ~x645 & ~x699 & ~x755 & ~x763 & ~x781;
assign c4373 =  x92 &  x101 &  x103 &  x123 &  x130 &  x159 &  x183 &  x234 &  x259 &  x268 &  x322 &  x486 &  x493 &  x625 &  x689 &  x745 & ~x46 & ~x52 & ~x59 & ~x89 & ~x106 & ~x107 & ~x165 & ~x534 & ~x557 & ~x588 & ~x646 & ~x672 & ~x725 & ~x763 & ~x764 & ~x775;
assign c4375 = ~x327 & ~x383 & ~x411 & ~x607;
assign c4377 = ~x434 & ~x547 & ~x572;
assign c4379 =  x66 &  x68 &  x69 &  x73 &  x96 &  x98 &  x99 &  x101 &  x102 &  x121 &  x126 &  x130 &  x147 &  x149 &  x150 &  x157 &  x158 &  x176 &  x177 &  x183 &  x210 &  x234 &  x235 &  x239 &  x244 &  x271 &  x288 &  x319 &  x328 &  x348 &  x373 &  x381 &  x385 &  x406 &  x432 &  x434 &  x457 &  x458 &  x460 &  x465 &  x486 &  x525 &  x543 &  x544 &  x553 &  x565 &  x570 &  x574 &  x575 &  x598 &  x621 &  x627 &  x658 &  x662 &  x678 & ~x3 & ~x20 & ~x24 & ~x30 & ~x54 & ~x55 & ~x78 & ~x80 & ~x109 & ~x116 & ~x142 & ~x143 & ~x170 & ~x221 & ~x222 & ~x223 & ~x254 & ~x278 & ~x280 & ~x306 & ~x309 & ~x310 & ~x334 & ~x362 & ~x392 & ~x394 & ~x395 & ~x445 & ~x448 & ~x450 & ~x451 & ~x532 & ~x563 & ~x590 & ~x615 & ~x616 & ~x645 & ~x669 & ~x731 & ~x748 & ~x759 & ~x764;
assign c4381 =  x112;
assign c4383 =  x63 &  x76 &  x90 &  x97 &  x285 &  x330 &  x380 & ~x5 & ~x22 & ~x34 & ~x616;
assign c4385 = ~x372;
assign c4389 =  x141;
assign c4391 =  x617;
assign c4393 =  x40 &  x41 &  x73 &  x92 &  x93 &  x94 &  x95 &  x97 &  x99 &  x120 &  x124 &  x126 &  x127 &  x129 &  x132 &  x148 &  x150 &  x152 &  x154 &  x156 &  x158 &  x160 &  x176 &  x178 &  x179 &  x184 &  x186 &  x188 &  x204 &  x215 &  x233 &  x234 &  x235 &  x239 &  x241 &  x244 &  x259 &  x264 &  x265 &  x267 &  x271 &  x287 &  x290 &  x293 &  x294 &  x295 &  x296 &  x297 &  x318 &  x320 &  x321 &  x322 &  x323 &  x324 &  x325 &  x343 &  x346 &  x348 &  x350 &  x351 &  x375 &  x376 &  x378 &  x380 &  x404 &  x406 &  x408 &  x409 &  x410 &  x430 &  x431 &  x432 &  x433 &  x434 &  x458 &  x462 &  x463 &  x485 &  x487 &  x513 &  x515 &  x519 &  x520 &  x521 &  x541 &  x575 &  x597 &  x602 &  x605 &  x633 &  x654 &  x656 &  x682 &  x683 &  x713 &  x716 &  x740 &  x741 &  x744 &  x745 &  x746 & ~x0 & ~x4 & ~x19 & ~x20 & ~x24 & ~x26 & ~x27 & ~x31 & ~x34 & ~x48 & ~x49 & ~x52 & ~x57 & ~x58 & ~x61 & ~x79 & ~x81 & ~x83 & ~x84 & ~x85 & ~x86 & ~x88 & ~x107 & ~x109 & ~x115 & ~x138 & ~x141 & ~x164 & ~x167 & ~x168 & ~x169 & ~x170 & ~x193 & ~x195 & ~x197 & ~x199 & ~x221 & ~x222 & ~x223 & ~x224 & ~x225 & ~x249 & ~x250 & ~x280 & ~x281 & ~x305 & ~x306 & ~x307 & ~x333 & ~x335 & ~x336 & ~x337 & ~x338 & ~x364 & ~x365 & ~x367 & ~x390 & ~x474 & ~x477 & ~x501 & ~x504 & ~x505 & ~x506 & ~x530 & ~x533 & ~x534 & ~x558 & ~x562 & ~x585 & ~x587 & ~x588 & ~x590 & ~x615 & ~x618 & ~x642 & ~x643 & ~x646 & ~x670 & ~x697 & ~x701 & ~x703 & ~x726 & ~x730 & ~x755 & ~x756 & ~x758 & ~x763;
assign c4395 = ~x98;
assign c4397 = ~x71;
assign c4399 =  x67 &  x68 &  x70 &  x94 &  x123 &  x127 &  x132 &  x150 &  x176 &  x182 &  x183 &  x245 &  x274 &  x286 &  x295 &  x314 &  x325 &  x343 &  x357 &  x374 &  x380 &  x403 &  x410 &  x453 &  x455 &  x460 &  x487 &  x489 &  x490 &  x491 &  x496 &  x515 &  x539 &  x543 &  x549 &  x565 &  x570 &  x576 &  x578 &  x605 &  x611 &  x621 &  x622 &  x630 &  x634 &  x661 & ~x2 & ~x22 & ~x51 & ~x52 & ~x54 & ~x82 & ~x109 & ~x137 & ~x167 & ~x170 & ~x249 & ~x252 & ~x306 & ~x307 & ~x309 & ~x365 & ~x366 & ~x394 & ~x473 & ~x478 & ~x479 & ~x505 & ~x561 & ~x585 & ~x616 & ~x647 & ~x671 & ~x701 & ~x728 & ~x729 & ~x756 & ~x763;
assign c4401 =  x10 &  x44 &  x130 &  x152 &  x297 &  x353 &  x408 &  x428 &  x487 &  x605 & ~x5 & ~x32 & ~x420 & ~x475 & ~x781;
assign c4403 = ~x412 & ~x510 & ~x539;
assign c4405 =  x89;
assign c4407 =  x196;
assign c4409 =  x304;
assign c4413 =  x58;
assign c4415 = ~x98;
assign c4417 =  x63 &  x90 &  x119 &  x162 &  x425 &  x634 &  x655 & ~x25 & ~x333;
assign c4419 = ~x664 & ~x686 & ~x688;
assign c4421 =  x337;
assign c4423 =  x69 &  x96 &  x101 &  x121 &  x126 &  x132 &  x154 &  x185 &  x204 &  x213 &  x232 &  x242 &  x244 &  x293 &  x314 &  x323 &  x330 &  x378 &  x433 &  x464 &  x493 &  x514 &  x522 &  x544 &  x627 &  x629 &  x654 & ~x3 & ~x26 & ~x28 & ~x29 & ~x36 & ~x37 & ~x47 & ~x81 & ~x82 & ~x83 & ~x106 & ~x109 & ~x138 & ~x143 & ~x167 & ~x171 & ~x194 & ~x336 & ~x338 & ~x396 & ~x417 & ~x420 & ~x446 & ~x475 & ~x530;
assign c4425 =  x419;
assign c4429 =  x587;
assign c4431 =  x15 &  x41 &  x42 &  x68 &  x69 &  x73 &  x95 &  x98 &  x126 &  x131 &  x149 &  x160 &  x176 &  x177 &  x213 &  x217 &  x241 &  x244 &  x260 &  x295 &  x300 &  x301 &  x344 &  x345 &  x375 &  x405 &  x407 &  x410 &  x442 &  x457 &  x459 &  x462 &  x517 &  x521 &  x570 &  x574 &  x626 &  x632 &  x685 &  x710 & ~x1 & ~x4 & ~x25 & ~x32 & ~x47 & ~x57 & ~x61 & ~x84 & ~x88 & ~x89 & ~x110 & ~x113 & ~x138 & ~x163 & ~x172 & ~x192 & ~x199 & ~x248 & ~x249 & ~x251 & ~x307 & ~x308 & ~x309 & ~x332 & ~x365 & ~x393 & ~x420 & ~x423 & ~x451 & ~x474 & ~x475 & ~x504 & ~x531 & ~x560 & ~x561 & ~x588 & ~x729 & ~x764 & ~x765;
assign c4433 =  x282;
assign c4435 =  x85;
assign c4437 = ~x98 & ~x181;
assign c4439 =  x87;
assign c4441 =  x69 &  x96 &  x119 &  x121 &  x122 &  x124 &  x125 &  x129 &  x146 &  x147 &  x154 &  x157 &  x158 &  x161 &  x174 &  x179 &  x209 &  x216 &  x217 &  x232 &  x241 &  x267 &  x293 &  x295 &  x301 &  x314 &  x317 &  x319 &  x321 &  x342 &  x348 &  x349 &  x409 &  x413 &  x427 &  x433 &  x435 &  x463 &  x491 &  x493 &  x497 &  x513 &  x517 &  x518 &  x519 &  x594 &  x597 &  x599 &  x627 &  x631 &  x649 &  x666 &  x706 &  x722 & ~x9 & ~x18 & ~x34 & ~x49 & ~x78 & ~x107 & ~x108 & ~x135 & ~x137 & ~x138 & ~x139 & ~x142 & ~x144 & ~x165 & ~x168 & ~x172 & ~x195 & ~x250 & ~x254 & ~x277 & ~x311 & ~x361 & ~x365 & ~x367 & ~x393 & ~x417 & ~x421 & ~x449 & ~x476 & ~x479 & ~x534 & ~x535 & ~x557 & ~x587 & ~x619 & ~x647 & ~x673 & ~x697 & ~x783;
assign c4443 =  x165;
assign c4445 = ~x210 & ~x571 & ~x660;
assign c4447 =  x77 &  x146 &  x218 & ~x333;
assign c4449 =  x66 &  x73 &  x75 &  x96 &  x97 &  x98 &  x99 &  x103 &  x125 &  x126 &  x130 &  x177 &  x186 &  x210 &  x265 &  x348 &  x352 &  x380 &  x405 &  x516 &  x542 &  x576 &  x629 &  x633 &  x655 &  x689 & ~x0 & ~x13 & ~x32 & ~x60 & ~x61 & ~x85 & ~x107 & ~x110 & ~x223 & ~x254 & ~x283 & ~x333 & ~x448 & ~x589 & ~x757;
assign c4451 =  x309;
assign c4455 =  x30;
assign c4457 =  x140;
assign c4459 =  x212 &  x716 & ~x369 & ~x510 & ~x526;
assign c4461 = ~x177 & ~x266;
assign c4463 =  x76 &  x104 &  x120 &  x121 &  x294 &  x462 &  x514 & ~x13 & ~x29 & ~x52 & ~x53 & ~x171 & ~x220 & ~x362 & ~x446 & ~x449;
assign c4465 =  x127 &  x182 & ~x199 & ~x443 & ~x453 & ~x529 & ~x554 & ~x566;
assign c4467 =  x77;
assign c4469 =  x108;
assign c4471 = ~x122 & ~x125;
assign c4473 =  x167;
assign c4475 =  x140;
assign c4477 =  x21;
assign c4479 =  x137;
assign c4481 = ~x518;
assign c4483 = ~x129 & ~x238;
assign c4485 = ~x384 & ~x496;
assign c4487 =  x54;
assign c4489 = ~x150 & ~x512 & ~x676;
assign c4491 =  x108;
assign c4493 =  x62 &  x117 &  x711;
assign c4495 =  x80;
assign c4497 =  x307;
assign c4499 =  x59;
assign c50 =  x484 & ~x268 & ~x297 & ~x578 & ~x687 & ~x765 & ~x775;
assign c52 = ~x0 & ~x5 & ~x7 & ~x8 & ~x13 & ~x15 & ~x33 & ~x34 & ~x36 & ~x41 & ~x59 & ~x69 & ~x84 & ~x91 & ~x94 & ~x97 & ~x111 & ~x121 & ~x139 & ~x140 & ~x142 & ~x146 & ~x148 & ~x170 & ~x174 & ~x177 & ~x178 & ~x198 & ~x199 & ~x201 & ~x202 & ~x205 & ~x225 & ~x228 & ~x229 & ~x230 & ~x232 & ~x252 & ~x258 & ~x281 & ~x285 & ~x286 & ~x287 & ~x288 & ~x313 & ~x338 & ~x364 & ~x365 & ~x378 & ~x392 & ~x393 & ~x407 & ~x422 & ~x435 & ~x734 & ~x758 & ~x761 & ~x764 & ~x781;
assign c54 =  x595 & ~x4 & ~x6 & ~x8 & ~x16 & ~x17 & ~x19 & ~x21 & ~x28 & ~x29 & ~x32 & ~x38 & ~x39 & ~x41 & ~x45 & ~x47 & ~x53 & ~x55 & ~x59 & ~x72 & ~x84 & ~x86 & ~x87 & ~x97 & ~x113 & ~x114 & ~x115 & ~x120 & ~x139 & ~x140 & ~x143 & ~x144 & ~x145 & ~x147 & ~x148 & ~x149 & ~x152 & ~x168 & ~x174 & ~x179 & ~x202 & ~x203 & ~x204 & ~x205 & ~x232 & ~x252 & ~x255 & ~x256 & ~x276 & ~x281 & ~x282 & ~x283 & ~x303 & ~x311 & ~x338 & ~x734 & ~x760 & ~x762 & ~x764 & ~x772 & ~x773 & ~x774 & ~x777;
assign c56 = ~x1 & ~x4 & ~x12 & ~x24 & ~x26 & ~x29 & ~x36 & ~x39 & ~x40 & ~x43 & ~x44 & ~x56 & ~x58 & ~x59 & ~x61 & ~x71 & ~x72 & ~x73 & ~x84 & ~x86 & ~x88 & ~x92 & ~x93 & ~x98 & ~x101 & ~x104 & ~x106 & ~x109 & ~x115 & ~x118 & ~x125 & ~x126 & ~x130 & ~x137 & ~x138 & ~x147 & ~x149 & ~x152 & ~x164 & ~x178 & ~x181 & ~x184 & ~x185 & ~x192 & ~x193 & ~x194 & ~x204 & ~x205 & ~x216 & ~x218 & ~x225 & ~x240 & ~x242 & ~x243 & ~x252 & ~x270 & ~x278 & ~x279 & ~x308 & ~x335 & ~x390 & ~x391 & ~x561 & ~x572 & ~x575 & ~x576 & ~x586 & ~x593 & ~x596 & ~x599 & ~x601 & ~x602 & ~x603 & ~x604 & ~x609 & ~x613 & ~x616 & ~x621 & ~x622 & ~x624 & ~x627 & ~x631 & ~x639 & ~x644 & ~x652 & ~x656 & ~x658 & ~x665 & ~x667 & ~x675 & ~x677 & ~x678 & ~x686 & ~x699 & ~x702 & ~x708 & ~x712 & ~x717 & ~x718 & ~x720 & ~x729 & ~x734 & ~x736 & ~x742 & ~x747 & ~x751 & ~x755 & ~x758 & ~x759 & ~x769 & ~x772 & ~x774;
assign c58 =  x549 & ~x2 & ~x3 & ~x11 & ~x15 & ~x18 & ~x21 & ~x22 & ~x25 & ~x30 & ~x32 & ~x33 & ~x35 & ~x36 & ~x37 & ~x42 & ~x53 & ~x59 & ~x60 & ~x61 & ~x62 & ~x72 & ~x83 & ~x88 & ~x89 & ~x90 & ~x93 & ~x111 & ~x113 & ~x117 & ~x118 & ~x120 & ~x142 & ~x143 & ~x144 & ~x145 & ~x148 & ~x166 & ~x168 & ~x174 & ~x176 & ~x198 & ~x200 & ~x202 & ~x203 & ~x204 & ~x205 & ~x227 & ~x229 & ~x230 & ~x252 & ~x255 & ~x259 & ~x260 & ~x280 & ~x282 & ~x289 & ~x308 & ~x311 & ~x336 & ~x340 & ~x391 & ~x419 & ~x448 & ~x503 & ~x614 & ~x615 & ~x699 & ~x756 & ~x758 & ~x762 & ~x772;
assign c510 =  x235 &  x266;
assign c512 =  x362 &  x593 & ~x10 & ~x31 & ~x35 & ~x43 & ~x55 & ~x69 & ~x71 & ~x95 & ~x149 & ~x168 & ~x173 & ~x197 & ~x252 & ~x256 & ~x259 & ~x260 & ~x283 & ~x339 & ~x341 & ~x364 & ~x366 & ~x392 & ~x759 & ~x769 & ~x770;
assign c514 = ~x0 & ~x3 & ~x7 & ~x11 & ~x31 & ~x35 & ~x37 & ~x42 & ~x58 & ~x66 & ~x112 & ~x114 & ~x116 & ~x121 & ~x175 & ~x196 & ~x203 & ~x204 & ~x223 & ~x225 & ~x228 & ~x230 & ~x232 & ~x233 & ~x256 & ~x258 & ~x280 & ~x284 & ~x286 & ~x311 & ~x336 & ~x338 & ~x340 & ~x341 & ~x394 & ~x421 & ~x423 & ~x435 & ~x476 & ~x477 & ~x580 & ~x608 & ~x636 & ~x663 & ~x689 & ~x746 & ~x748 & ~x755 & ~x770 & ~x773 & ~x774;
assign c516 =  x454 & ~x0 & ~x6 & ~x10 & ~x16 & ~x25 & ~x29 & ~x37 & ~x41 & ~x42 & ~x44 & ~x47 & ~x52 & ~x53 & ~x54 & ~x55 & ~x59 & ~x60 & ~x61 & ~x62 & ~x64 & ~x69 & ~x72 & ~x73 & ~x79 & ~x81 & ~x82 & ~x84 & ~x88 & ~x90 & ~x91 & ~x96 & ~x97 & ~x98 & ~x101 & ~x108 & ~x111 & ~x113 & ~x115 & ~x117 & ~x132 & ~x133 & ~x134 & ~x137 & ~x142 & ~x145 & ~x148 & ~x151 & ~x158 & ~x159 & ~x167 & ~x178 & ~x179 & ~x182 & ~x184 & ~x202 & ~x203 & ~x204 & ~x208 & ~x222 & ~x228 & ~x230 & ~x231 & ~x257 & ~x283 & ~x284 & ~x310 & ~x348 & ~x394 & ~x615 & ~x637 & ~x657 & ~x658 & ~x663 & ~x672 & ~x673 & ~x674 & ~x678 & ~x686 & ~x689 & ~x690 & ~x693 & ~x697 & ~x701 & ~x705 & ~x710 & ~x715 & ~x716 & ~x719 & ~x721 & ~x738 & ~x739 & ~x746 & ~x747 & ~x748 & ~x751 & ~x761 & ~x762 & ~x763 & ~x764 & ~x771 & ~x779;
assign c518 =  x481 & ~x9 & ~x42 & ~x68 & ~x111 & ~x123 & ~x150 & ~x228 & ~x232 & ~x310 & ~x337 & ~x377 & ~x657 & ~x677 & ~x717 & ~x722;
assign c520 =  x78 & ~x21 & ~x62 & ~x115 & ~x197 & ~x368 & ~x371;
assign c522 =  x457 & ~x91 & ~x298 & ~x506 & ~x507 & ~x531 & ~x652;
assign c524 = ~x0 & ~x1 & ~x3 & ~x7 & ~x13 & ~x22 & ~x55 & ~x62 & ~x64 & ~x67 & ~x83 & ~x89 & ~x120 & ~x139 & ~x143 & ~x144 & ~x145 & ~x146 & ~x169 & ~x177 & ~x178 & ~x198 & ~x199 & ~x200 & ~x202 & ~x203 & ~x225 & ~x226 & ~x231 & ~x252 & ~x281 & ~x287 & ~x288 & ~x312 & ~x314 & ~x367 & ~x414 & ~x420 & ~x423 & ~x448 & ~x451 & ~x478 & ~x504 & ~x532 & ~x643 & ~x671 & ~x672 & ~x727 & ~x743 & ~x755 & ~x759 & ~x772;
assign c526 =  x428 &  x429 &  x455 & ~x7 & ~x88 & ~x98 & ~x140 & ~x166 & ~x214 & ~x334 & ~x491 & ~x657 & ~x750 & ~x751;
assign c528 = ~x5 & ~x9 & ~x12 & ~x16 & ~x18 & ~x26 & ~x28 & ~x29 & ~x30 & ~x31 & ~x34 & ~x36 & ~x38 & ~x39 & ~x54 & ~x59 & ~x60 & ~x61 & ~x63 & ~x64 & ~x82 & ~x84 & ~x86 & ~x89 & ~x91 & ~x92 & ~x113 & ~x116 & ~x117 & ~x118 & ~x119 & ~x121 & ~x138 & ~x140 & ~x142 & ~x143 & ~x144 & ~x145 & ~x146 & ~x169 & ~x170 & ~x173 & ~x174 & ~x197 & ~x200 & ~x203 & ~x205 & ~x206 & ~x222 & ~x226 & ~x227 & ~x229 & ~x231 & ~x252 & ~x254 & ~x256 & ~x257 & ~x283 & ~x286 & ~x288 & ~x311 & ~x314 & ~x337 & ~x364 & ~x365 & ~x368 & ~x448 & ~x475 & ~x476 & ~x478 & ~x504 & ~x507 & ~x532 & ~x552 & ~x563 & ~x579 & ~x580 & ~x590 & ~x607 & ~x616 & ~x617 & ~x700 & ~x744 & ~x755 & ~x771 & ~x772;
assign c530 =  x75 & ~x61 & ~x140 & ~x147 & ~x203 & ~x230 & ~x255 & ~x256 & ~x309 & ~x341 & ~x370 & ~x478;
assign c532 =  x427 &  x543 &  x567 & ~x13 & ~x110 & ~x202 & ~x232 & ~x279 & ~x287 & ~x288 & ~x311 & ~x312 & ~x616 & ~x717 & ~x719 & ~x745 & ~x756 & ~x764;
assign c534 = ~x4 & ~x6 & ~x7 & ~x14 & ~x18 & ~x19 & ~x21 & ~x27 & ~x36 & ~x40 & ~x49 & ~x57 & ~x60 & ~x63 & ~x69 & ~x70 & ~x86 & ~x90 & ~x97 & ~x115 & ~x116 & ~x119 & ~x121 & ~x123 & ~x140 & ~x141 & ~x149 & ~x169 & ~x173 & ~x175 & ~x181 & ~x201 & ~x202 & ~x203 & ~x224 & ~x226 & ~x227 & ~x228 & ~x252 & ~x253 & ~x257 & ~x258 & ~x261 & ~x281 & ~x283 & ~x284 & ~x286 & ~x288 & ~x289 & ~x308 & ~x312 & ~x313 & ~x339 & ~x361 & ~x364 & ~x367 & ~x394 & ~x395 & ~x531 & ~x560 & ~x579 & ~x580 & ~x661 & ~x662 & ~x672 & ~x700 & ~x715 & ~x729 & ~x747 & ~x748 & ~x767 & ~x777 & ~x781 & ~x782;
assign c536 =  x425 & ~x93 & ~x269 & ~x297 & ~x692 & ~x693 & ~x736 & ~x750;
assign c538 =  x131 &  x132 & ~x10 & ~x11 & ~x21 & ~x30 & ~x33 & ~x34 & ~x58 & ~x60 & ~x61 & ~x62 & ~x84 & ~x85 & ~x86 & ~x87 & ~x88 & ~x89 & ~x112 & ~x116 & ~x119 & ~x140 & ~x143 & ~x167 & ~x173 & ~x174 & ~x197 & ~x199 & ~x223 & ~x224 & ~x225 & ~x227 & ~x230 & ~x231 & ~x256 & ~x258 & ~x259 & ~x286 & ~x288 & ~x312 & ~x313 & ~x316 & ~x336 & ~x337 & ~x338 & ~x341 & ~x342 & ~x364 & ~x369 & ~x393 & ~x395 & ~x421 & ~x423 & ~x448 & ~x450 & ~x451 & ~x671;
assign c540 =  x444 &  x472 &  x473 & ~x3 & ~x5 & ~x6 & ~x15 & ~x17 & ~x19 & ~x25 & ~x34 & ~x35 & ~x37 & ~x85 & ~x87 & ~x117 & ~x118 & ~x140 & ~x142 & ~x146 & ~x148 & ~x149 & ~x173 & ~x177 & ~x200 & ~x201 & ~x203 & ~x204 & ~x230 & ~x233 & ~x256 & ~x257 & ~x260 & ~x261 & ~x284 & ~x308 & ~x309 & ~x310 & ~x313 & ~x350 & ~x379 & ~x420 & ~x730 & ~x757 & ~x758 & ~x762 & ~x771 & ~x772 & ~x773 & ~x778;
assign c542 =  x351 &  x482 &  x483 &  x486 & ~x2 & ~x10 & ~x16 & ~x21 & ~x24 & ~x37 & ~x50 & ~x56 & ~x61 & ~x64 & ~x67 & ~x73 & ~x74 & ~x79 & ~x83 & ~x86 & ~x99 & ~x101 & ~x118 & ~x126 & ~x131 & ~x135 & ~x144 & ~x146 & ~x152 & ~x154 & ~x155 & ~x166 & ~x169 & ~x170 & ~x174 & ~x176 & ~x177 & ~x188 & ~x209 & ~x211 & ~x214 & ~x226 & ~x229 & ~x230 & ~x240 & ~x243 & ~x252 & ~x257 & ~x259 & ~x269 & ~x270 & ~x310 & ~x504 & ~x573 & ~x574 & ~x576 & ~x591 & ~x593 & ~x600 & ~x606 & ~x616 & ~x617 & ~x618 & ~x630 & ~x644 & ~x649 & ~x650 & ~x675 & ~x679 & ~x683 & ~x688 & ~x690 & ~x692 & ~x699 & ~x703 & ~x714 & ~x721 & ~x723 & ~x737 & ~x748 & ~x751 & ~x756 & ~x777;
assign c544 = ~x1 & ~x2 & ~x3 & ~x5 & ~x6 & ~x7 & ~x10 & ~x11 & ~x12 & ~x13 & ~x14 & ~x16 & ~x20 & ~x21 & ~x28 & ~x29 & ~x31 & ~x32 & ~x33 & ~x35 & ~x36 & ~x37 & ~x39 & ~x40 & ~x55 & ~x57 & ~x61 & ~x64 & ~x67 & ~x83 & ~x84 & ~x85 & ~x89 & ~x90 & ~x91 & ~x92 & ~x111 & ~x113 & ~x116 & ~x117 & ~x119 & ~x120 & ~x122 & ~x123 & ~x124 & ~x140 & ~x142 & ~x143 & ~x144 & ~x145 & ~x146 & ~x148 & ~x149 & ~x150 & ~x151 & ~x152 & ~x168 & ~x172 & ~x173 & ~x177 & ~x178 & ~x195 & ~x196 & ~x199 & ~x201 & ~x202 & ~x203 & ~x207 & ~x208 & ~x223 & ~x224 & ~x227 & ~x229 & ~x231 & ~x233 & ~x253 & ~x254 & ~x256 & ~x257 & ~x258 & ~x259 & ~x260 & ~x261 & ~x264 & ~x280 & ~x283 & ~x284 & ~x308 & ~x309 & ~x310 & ~x311 & ~x353 & ~x354 & ~x365 & ~x366 & ~x420 & ~x476 & ~x587 & ~x588 & ~x616 & ~x643 & ~x672 & ~x728 & ~x729 & ~x758 & ~x773 & ~x782;
assign c546 = ~x0 & ~x11 & ~x12 & ~x14 & ~x27 & ~x30 & ~x35 & ~x57 & ~x60 & ~x63 & ~x84 & ~x86 & ~x111 & ~x113 & ~x114 & ~x116 & ~x170 & ~x171 & ~x173 & ~x175 & ~x200 & ~x201 & ~x204 & ~x225 & ~x226 & ~x230 & ~x286 & ~x288 & ~x308 & ~x312 & ~x314 & ~x336 & ~x342 & ~x344 & ~x368 & ~x395 & ~x396 & ~x398 & ~x420 & ~x421 & ~x432 & ~x433 & ~x449 & ~x451 & ~x461 & ~x700 & ~x782;
assign c548 =  x485 & ~x12 & ~x38 & ~x40 & ~x45 & ~x64 & ~x69 & ~x92 & ~x95 & ~x112 & ~x113 & ~x115 & ~x141 & ~x145 & ~x152 & ~x202 & ~x225 & ~x446 & ~x737 & ~x744 & ~x771 & ~x772 & ~x774 & ~x780;
assign c550 =  x331 &  x358 &  x359 & ~x42 & ~x109 & ~x318 & ~x731;
assign c552 =  x428 & ~x3 & ~x5 & ~x7 & ~x11 & ~x13 & ~x20 & ~x21 & ~x23 & ~x28 & ~x35 & ~x38 & ~x39 & ~x56 & ~x59 & ~x62 & ~x71 & ~x72 & ~x86 & ~x90 & ~x112 & ~x117 & ~x118 & ~x119 & ~x120 & ~x142 & ~x172 & ~x173 & ~x174 & ~x197 & ~x199 & ~x224 & ~x227 & ~x252 & ~x254 & ~x259 & ~x284 & ~x286 & ~x313 & ~x314 & ~x340 & ~x449 & ~x559 & ~x728 & ~x756 & ~x761 & ~x764 & ~x765 & ~x770 & ~x774 & ~x781;
assign c554 =  x301 & ~x64 & ~x146 & ~x338 & ~x410;
assign c556 =  x621 & ~x10 & ~x13 & ~x14 & ~x19 & ~x36 & ~x113 & ~x144 & ~x202 & ~x225 & ~x227 & ~x281 & ~x285 & ~x308 & ~x312 & ~x313 & ~x316 & ~x396 & ~x421 & ~x448 & ~x763;
assign c558 =  x466 & ~x64 & ~x230 & ~x286 & ~x333 & ~x359 & ~x360 & ~x367 & ~x718;
assign c560 =  x595 &  x697 & ~x10 & ~x225 & ~x258 & ~x422;
assign c562 =  x248 & ~x16 & ~x35 & ~x55 & ~x58 & ~x64 & ~x93 & ~x118 & ~x119 & ~x141 & ~x174 & ~x176 & ~x223 & ~x226 & ~x228 & ~x337 & ~x561 & ~x615 & ~x618 & ~x633 & ~x635 & ~x692 & ~x745 & ~x779;
assign c564 =  x397 &  x426 & ~x8 & ~x60 & ~x92 & ~x371 & ~x559 & ~x765;
assign c566 =  x438 & ~x13 & ~x41 & ~x94 & ~x118 & ~x180 & ~x295 & ~x333 & ~x560;
assign c568 =  x377 & ~x5 & ~x6 & ~x7 & ~x24 & ~x31 & ~x39 & ~x43 & ~x64 & ~x67 & ~x89 & ~x92 & ~x120 & ~x140 & ~x144 & ~x175 & ~x201 & ~x205 & ~x226 & ~x231 & ~x259 & ~x262 & ~x283 & ~x285 & ~x286 & ~x309 & ~x312 & ~x367 & ~x381 & ~x643 & ~x671 & ~x761 & ~x771 & ~x772;
assign c570 =  x399 &  x499 & ~x3 & ~x11 & ~x13 & ~x18 & ~x23 & ~x39 & ~x42 & ~x63 & ~x84 & ~x101 & ~x103 & ~x105 & ~x110 & ~x112 & ~x116 & ~x117 & ~x118 & ~x144 & ~x172 & ~x319 & ~x335 & ~x632 & ~x647 & ~x652 & ~x659 & ~x663 & ~x665 & ~x666 & ~x677 & ~x678 & ~x686 & ~x712 & ~x714 & ~x727 & ~x756 & ~x761 & ~x770;
assign c572 =  x165 & ~x31 & ~x81 & ~x171;
assign c574 =  x736 &  x738 &  x739 & ~x3 & ~x7 & ~x12 & ~x33 & ~x34 & ~x56 & ~x57 & ~x86 & ~x115 & ~x117 & ~x170 & ~x197 & ~x230 & ~x233 & ~x253 & ~x256 & ~x284 & ~x287 & ~x314 & ~x341 & ~x344 & ~x369 & ~x370 & ~x392 & ~x395 & ~x398 & ~x399 & ~x400 & ~x420 & ~x421 & ~x426 & ~x427 & ~x452 & ~x477 & ~x478 & ~x504 & ~x505 & ~x560 & ~x587;
assign c576 =  x549 & ~x55 & ~x87 & ~x113 & ~x141 & ~x216 & ~x224 & ~x285 & ~x312 & ~x316 & ~x339 & ~x344 & ~x365 & ~x373 & ~x449 & ~x478 & ~x771;
assign c578 = ~x4 & ~x6 & ~x7 & ~x10 & ~x13 & ~x16 & ~x17 & ~x24 & ~x32 & ~x33 & ~x37 & ~x39 & ~x45 & ~x53 & ~x58 & ~x63 & ~x65 & ~x70 & ~x75 & ~x77 & ~x81 & ~x83 & ~x84 & ~x88 & ~x89 & ~x91 & ~x100 & ~x104 & ~x112 & ~x116 & ~x117 & ~x127 & ~x128 & ~x139 & ~x142 & ~x150 & ~x167 & ~x171 & ~x172 & ~x173 & ~x195 & ~x197 & ~x198 & ~x202 & ~x206 & ~x225 & ~x226 & ~x228 & ~x255 & ~x257 & ~x258 & ~x259 & ~x260 & ~x281 & ~x283 & ~x308 & ~x314 & ~x337 & ~x341 & ~x365 & ~x368 & ~x392 & ~x393 & ~x532 & ~x534 & ~x702 & ~x713 & ~x716 & ~x727 & ~x728 & ~x731 & ~x736 & ~x737 & ~x741 & ~x745 & ~x746 & ~x747 & ~x749 & ~x750 & ~x767 & ~x769 & ~x770 & ~x773 & ~x776 & ~x778 & ~x782;
assign c580 =  x482 & ~x4 & ~x12 & ~x15 & ~x19 & ~x28 & ~x35 & ~x38 & ~x39 & ~x40 & ~x41 & ~x44 & ~x52 & ~x61 & ~x62 & ~x64 & ~x68 & ~x70 & ~x72 & ~x92 & ~x94 & ~x95 & ~x98 & ~x114 & ~x121 & ~x128 & ~x148 & ~x149 & ~x151 & ~x173 & ~x174 & ~x176 & ~x179 & ~x200 & ~x201 & ~x225 & ~x256 & ~x270 & ~x308 & ~x310 & ~x311 & ~x338 & ~x419 & ~x445 & ~x560 & ~x631 & ~x716 & ~x721 & ~x730 & ~x734 & ~x746 & ~x748 & ~x751 & ~x760 & ~x764 & ~x767 & ~x769 & ~x773 & ~x777 & ~x778 & ~x779 & ~x781;
assign c582 = ~x12 & ~x27 & ~x38 & ~x44 & ~x56 & ~x63 & ~x64 & ~x66 & ~x68 & ~x71 & ~x94 & ~x96 & ~x113 & ~x116 & ~x139 & ~x141 & ~x145 & ~x149 & ~x151 & ~x172 & ~x173 & ~x177 & ~x195 & ~x198 & ~x206 & ~x226 & ~x227 & ~x334 & ~x336 & ~x448 & ~x469 & ~x603 & ~x606 & ~x607 & ~x635 & ~x663 & ~x716 & ~x727 & ~x757 & ~x759 & ~x774;
assign c584 =  x400 &  x427 &  x537 &  x547 & ~x0 & ~x3 & ~x9 & ~x15 & ~x21 & ~x30 & ~x32 & ~x36 & ~x52 & ~x53 & ~x69 & ~x71 & ~x75 & ~x90 & ~x91 & ~x93 & ~x103 & ~x110 & ~x114 & ~x121 & ~x126 & ~x133 & ~x172 & ~x178 & ~x196 & ~x197 & ~x199 & ~x280 & ~x281 & ~x308 & ~x309 & ~x649 & ~x673 & ~x676 & ~x692 & ~x699 & ~x717 & ~x733 & ~x744 & ~x746 & ~x748 & ~x765 & ~x769 & ~x771 & ~x774;
assign c586 = ~x55 & ~x170 & ~x233 & ~x287 & ~x297 & ~x343 & ~x344 & ~x378;
assign c588 = ~x1 & ~x2 & ~x3 & ~x4 & ~x11 & ~x15 & ~x21 & ~x24 & ~x32 & ~x33 & ~x40 & ~x42 & ~x51 & ~x54 & ~x55 & ~x57 & ~x59 & ~x63 & ~x67 & ~x84 & ~x114 & ~x119 & ~x123 & ~x141 & ~x143 & ~x147 & ~x149 & ~x170 & ~x171 & ~x172 & ~x173 & ~x176 & ~x177 & ~x196 & ~x201 & ~x207 & ~x223 & ~x224 & ~x226 & ~x227 & ~x228 & ~x231 & ~x232 & ~x233 & ~x253 & ~x254 & ~x255 & ~x257 & ~x260 & ~x281 & ~x284 & ~x286 & ~x288 & ~x308 & ~x309 & ~x311 & ~x313 & ~x314 & ~x315 & ~x316 & ~x337 & ~x345 & ~x364 & ~x370 & ~x421 & ~x435 & ~x448 & ~x451 & ~x463 & ~x616 & ~x757 & ~x758 & ~x781;
assign c590 =  x267 &  x481 &  x545 & ~x16 & ~x29 & ~x102 & ~x158 & ~x290 & ~x767 & ~x781;
assign c592 =  x357 &  x360 &  x399 &  x412 &  x466 & ~x42 & ~x46 & ~x77 & ~x116 & ~x197 & ~x311 & ~x318 & ~x319 & ~x700 & ~x775;
assign c594 =  x265 &  x438 & ~x71 & ~x281 & ~x311 & ~x636 & ~x647 & ~x669 & ~x728 & ~x778;
assign c596 =  x359 &  x362 &  x427 &  x466 &  x482 & ~x11 & ~x13 & ~x36 & ~x69 & ~x96 & ~x121 & ~x140 & ~x141 & ~x167 & ~x204 & ~x226 & ~x257 & ~x281 & ~x286 & ~x364 & ~x531 & ~x559 & ~x671 & ~x776;
assign c598 =  x217 & ~x27 & ~x203 & ~x249 & ~x392 & ~x450 & ~x752;
assign c5100 =  x370 &  x480 &  x494 &  x502 & ~x13 & ~x36 & ~x40 & ~x44 & ~x60 & ~x74 & ~x97 & ~x114 & ~x169 & ~x228 & ~x242 & ~x627 & ~x631 & ~x654 & ~x678 & ~x687 & ~x689 & ~x704 & ~x760 & ~x769;
assign c5102 =  x266 &  x425 &  x511 &  x520 &  x542 & ~x5 & ~x27 & ~x63 & ~x88 & ~x97 & ~x145 & ~x146 & ~x157 & ~x176 & ~x178 & ~x185 & ~x198 & ~x255 & ~x258 & ~x660 & ~x702 & ~x740 & ~x747 & ~x771;
assign c5104 =  x106 & ~x0 & ~x5 & ~x8 & ~x9 & ~x12 & ~x20 & ~x30 & ~x59 & ~x84 & ~x115 & ~x116 & ~x139 & ~x143 & ~x199 & ~x225 & ~x228 & ~x283 & ~x284 & ~x340 & ~x341 & ~x342 & ~x365 & ~x366 & ~x644 & ~x728 & ~x755 & ~x756 & ~x783;
assign c5106 =  x451 &  x456 & ~x53 & ~x57 & ~x70 & ~x94 & ~x120 & ~x126 & ~x132 & ~x139 & ~x144 & ~x181 & ~x211 & ~x226 & ~x268 & ~x269 & ~x311 & ~x614 & ~x616 & ~x643 & ~x648 & ~x649 & ~x658 & ~x659 & ~x717 & ~x720 & ~x722 & ~x724 & ~x743 & ~x750;
assign c5108 =  x453 & ~x55 & ~x64 & ~x70 & ~x71 & ~x75 & ~x145 & ~x199 & ~x208 & ~x211 & ~x214 & ~x240 & ~x268 & ~x269 & ~x270 & ~x572 & ~x575 & ~x583 & ~x695 & ~x713 & ~x718 & ~x742 & ~x744 & ~x752 & ~x760;
assign c5110 =  x565 &  x567 & ~x0 & ~x1 & ~x9 & ~x13 & ~x14 & ~x18 & ~x20 & ~x27 & ~x33 & ~x36 & ~x39 & ~x40 & ~x41 & ~x44 & ~x45 & ~x55 & ~x60 & ~x61 & ~x66 & ~x86 & ~x94 & ~x95 & ~x113 & ~x116 & ~x120 & ~x140 & ~x141 & ~x143 & ~x144 & ~x168 & ~x170 & ~x171 & ~x172 & ~x202 & ~x204 & ~x226 & ~x227 & ~x228 & ~x230 & ~x232 & ~x253 & ~x254 & ~x259 & ~x281 & ~x286 & ~x312 & ~x313 & ~x314 & ~x342 & ~x366 & ~x368 & ~x392 & ~x395 & ~x421 & ~x422 & ~x449 & ~x506 & ~x700 & ~x730 & ~x732 & ~x762 & ~x766 & ~x769 & ~x777 & ~x780 & ~x783;
assign c5112 =  x267 &  x295 &  x325 &  x326 &  x483 &  x526 & ~x7 & ~x11 & ~x18 & ~x21 & ~x37 & ~x57 & ~x59 & ~x68 & ~x69 & ~x70 & ~x72 & ~x79 & ~x87 & ~x91 & ~x100 & ~x116 & ~x120 & ~x127 & ~x130 & ~x137 & ~x140 & ~x150 & ~x154 & ~x155 & ~x158 & ~x179 & ~x194 & ~x203 & ~x225 & ~x229 & ~x232 & ~x252 & ~x259 & ~x282 & ~x286 & ~x309 & ~x339 & ~x364 & ~x365 & ~x532 & ~x590 & ~x607 & ~x614 & ~x615 & ~x636 & ~x671 & ~x672 & ~x674 & ~x700 & ~x706 & ~x735 & ~x744 & ~x745 & ~x747 & ~x748 & ~x750 & ~x782 & ~x783;
assign c5114 =  x412 & ~x2 & ~x10 & ~x12 & ~x15 & ~x21 & ~x26 & ~x31 & ~x32 & ~x36 & ~x37 & ~x43 & ~x46 & ~x52 & ~x59 & ~x62 & ~x66 & ~x67 & ~x71 & ~x75 & ~x78 & ~x82 & ~x83 & ~x85 & ~x97 & ~x98 & ~x99 & ~x102 & ~x124 & ~x170 & ~x173 & ~x176 & ~x195 & ~x197 & ~x201 & ~x202 & ~x207 & ~x208 & ~x227 & ~x285 & ~x287 & ~x289 & ~x309 & ~x310 & ~x337 & ~x406 & ~x672 & ~x703 & ~x742 & ~x743 & ~x744 & ~x745 & ~x754 & ~x757 & ~x759 & ~x761 & ~x769 & ~x773 & ~x774 & ~x783;
assign c5116 =  x490 &  x500 & ~x0 & ~x30 & ~x39 & ~x117 & ~x202 & ~x213 & ~x241 & ~x242 & ~x270 & ~x551 & ~x554 & ~x587 & ~x653 & ~x689 & ~x724 & ~x726 & ~x760 & ~x769;
assign c5118 =  x399 &  x453 &  x508 &  x523 &  x543 & ~x1 & ~x18 & ~x32 & ~x33 & ~x64 & ~x83 & ~x91 & ~x93 & ~x130 & ~x140 & ~x145 & ~x150 & ~x232 & ~x616 & ~x679 & ~x681 & ~x686 & ~x695 & ~x700 & ~x705 & ~x731 & ~x741 & ~x745 & ~x749 & ~x761;
assign c5120 =  x334 &  x359 &  x622 &  x624 & ~x0 & ~x11 & ~x12 & ~x20 & ~x26 & ~x30 & ~x31 & ~x84 & ~x111 & ~x115 & ~x141 & ~x170 & ~x197 & ~x254 & ~x259 & ~x282 & ~x314 & ~x338 & ~x340 & ~x342 & ~x364 & ~x559 & ~x783;
assign c5122 =  x326 &  x535 &  x545 &  x557 & ~x39 & ~x213;
assign c5124 =  x585 & ~x6 & ~x13 & ~x27 & ~x32 & ~x33 & ~x57 & ~x61 & ~x87 & ~x199 & ~x200 & ~x201 & ~x280 & ~x284 & ~x534 & ~x579 & ~x607 & ~x718 & ~x719 & ~x757 & ~x775;
assign c5126 =  x708 &  x711 & ~x4 & ~x9 & ~x13 & ~x25 & ~x26 & ~x29 & ~x36 & ~x57 & ~x58 & ~x59 & ~x63 & ~x64 & ~x88 & ~x89 & ~x170 & ~x253 & ~x285 & ~x308 & ~x313 & ~x338 & ~x340 & ~x344 & ~x369 & ~x371 & ~x372 & ~x392 & ~x393 & ~x395 & ~x396 & ~x398 & ~x400 & ~x421 & ~x478 & ~x503 & ~x507 & ~x587 & ~x644 & ~x671;
assign c5128 =  x412 &  x427 & ~x16 & ~x57 & ~x58 & ~x64 & ~x77 & ~x86 & ~x89 & ~x97 & ~x101 & ~x104 & ~x118 & ~x146 & ~x180 & ~x197 & ~x209 & ~x214 & ~x225 & ~x241 & ~x256 & ~x286 & ~x306 & ~x334 & ~x335 & ~x560 & ~x575 & ~x635 & ~x676 & ~x692 & ~x705 & ~x707 & ~x713 & ~x716 & ~x718 & ~x730 & ~x731 & ~x744 & ~x761 & ~x775 & ~x781;
assign c5130 =  x714 & ~x37 & ~x83 & ~x90 & ~x144 & ~x145 & ~x230 & ~x284 & ~x309 & ~x343 & ~x370 & ~x391 & ~x392 & ~x397 & ~x398 & ~x400 & ~x451 & ~x478 & ~x643 & ~x671 & ~x672;
assign c5132 =  x439 & ~x0 & ~x1 & ~x3 & ~x4 & ~x5 & ~x6 & ~x8 & ~x9 & ~x10 & ~x11 & ~x13 & ~x14 & ~x20 & ~x21 & ~x24 & ~x28 & ~x30 & ~x31 & ~x32 & ~x33 & ~x40 & ~x53 & ~x55 & ~x56 & ~x57 & ~x58 & ~x59 & ~x60 & ~x61 & ~x62 & ~x63 & ~x84 & ~x86 & ~x87 & ~x88 & ~x89 & ~x91 & ~x113 & ~x115 & ~x116 & ~x117 & ~x119 & ~x143 & ~x145 & ~x149 & ~x150 & ~x167 & ~x168 & ~x169 & ~x170 & ~x173 & ~x174 & ~x175 & ~x177 & ~x197 & ~x199 & ~x200 & ~x202 & ~x204 & ~x205 & ~x224 & ~x225 & ~x228 & ~x230 & ~x232 & ~x233 & ~x252 & ~x253 & ~x254 & ~x255 & ~x256 & ~x259 & ~x261 & ~x280 & ~x281 & ~x282 & ~x283 & ~x286 & ~x287 & ~x309 & ~x310 & ~x312 & ~x314 & ~x338 & ~x339 & ~x340 & ~x364 & ~x366 & ~x372 & ~x391 & ~x448 & ~x476 & ~x477 & ~x478 & ~x479 & ~x504 & ~x505 & ~x506 & ~x507 & ~x532 & ~x559 & ~x560 & ~x616 & ~x699 & ~x728 & ~x755 & ~x756 & ~x757 & ~x758 & ~x759 & ~x783;
assign c5134 =  x539 & ~x1 & ~x3 & ~x4 & ~x5 & ~x7 & ~x9 & ~x10 & ~x12 & ~x14 & ~x15 & ~x17 & ~x20 & ~x22 & ~x25 & ~x26 & ~x27 & ~x28 & ~x29 & ~x30 & ~x32 & ~x38 & ~x39 & ~x40 & ~x41 & ~x42 & ~x43 & ~x44 & ~x45 & ~x46 & ~x52 & ~x53 & ~x54 & ~x56 & ~x58 & ~x59 & ~x60 & ~x61 & ~x62 & ~x63 & ~x64 & ~x65 & ~x66 & ~x68 & ~x69 & ~x70 & ~x71 & ~x73 & ~x74 & ~x77 & ~x79 & ~x82 & ~x83 & ~x84 & ~x85 & ~x87 & ~x89 & ~x92 & ~x94 & ~x110 & ~x111 & ~x112 & ~x113 & ~x114 & ~x115 & ~x117 & ~x118 & ~x120 & ~x122 & ~x123 & ~x125 & ~x126 & ~x138 & ~x140 & ~x141 & ~x142 & ~x143 & ~x146 & ~x147 & ~x148 & ~x149 & ~x150 & ~x167 & ~x168 & ~x169 & ~x170 & ~x171 & ~x173 & ~x174 & ~x177 & ~x178 & ~x179 & ~x180 & ~x195 & ~x197 & ~x198 & ~x199 & ~x201 & ~x203 & ~x204 & ~x223 & ~x224 & ~x226 & ~x229 & ~x230 & ~x231 & ~x232 & ~x233 & ~x252 & ~x253 & ~x254 & ~x256 & ~x257 & ~x259 & ~x283 & ~x284 & ~x285 & ~x289 & ~x308 & ~x310 & ~x312 & ~x337 & ~x338 & ~x340 & ~x364 & ~x365 & ~x392 & ~x393 & ~x395 & ~x420 & ~x421 & ~x422 & ~x450 & ~x477 & ~x478 & ~x700 & ~x703 & ~x704 & ~x706 & ~x711 & ~x718 & ~x727 & ~x730 & ~x732 & ~x733 & ~x735 & ~x737 & ~x738 & ~x739 & ~x740 & ~x741 & ~x742 & ~x743 & ~x745 & ~x746 & ~x747 & ~x748 & ~x749 & ~x750 & ~x754 & ~x755 & ~x756 & ~x757 & ~x758 & ~x759 & ~x760 & ~x761 & ~x763 & ~x764 & ~x766 & ~x767 & ~x771 & ~x773 & ~x775 & ~x776 & ~x778 & ~x780 & ~x781 & ~x782 & ~x783;
assign c5136 =  x652 & ~x9 & ~x11 & ~x59 & ~x141 & ~x148 & ~x195 & ~x254 & ~x255 & ~x280 & ~x310 & ~x314 & ~x315 & ~x341 & ~x369 & ~x398 & ~x423 & ~x449 & ~x591 & ~x692;
assign c5138 = ~x5 & ~x37 & ~x39 & ~x43 & ~x71 & ~x82 & ~x85 & ~x93 & ~x95 & ~x111 & ~x168 & ~x172 & ~x178 & ~x203 & ~x205 & ~x226 & ~x230 & ~x260 & ~x284 & ~x287 & ~x288 & ~x310 & ~x314 & ~x316 & ~x339 & ~x368 & ~x394 & ~x395 & ~x410 & ~x421 & ~x437 & ~x699 & ~x702 & ~x716 & ~x723 & ~x777 & ~x783;
assign c5140 =  x191 & ~x2 & ~x29 & ~x36 & ~x56 & ~x61 & ~x89 & ~x114 & ~x115 & ~x117 & ~x118 & ~x119 & ~x139 & ~x145 & ~x167 & ~x168 & ~x199 & ~x200 & ~x224 & ~x225 & ~x230 & ~x309 & ~x560 & ~x617 & ~x618 & ~x661 & ~x716 & ~x717 & ~x720 & ~x773 & ~x777;
assign c5142 =  x512 & ~x1 & ~x35 & ~x43 & ~x113 & ~x195 & ~x422 & ~x451 & ~x462 & ~x671 & ~x700 & ~x728 & ~x783;
assign c5144 =  x265 &  x466 & ~x0 & ~x1 & ~x4 & ~x24 & ~x27 & ~x32 & ~x33 & ~x37 & ~x56 & ~x60 & ~x63 & ~x64 & ~x82 & ~x89 & ~x94 & ~x110 & ~x111 & ~x117 & ~x118 & ~x120 & ~x121 & ~x140 & ~x146 & ~x167 & ~x169 & ~x176 & ~x197 & ~x200 & ~x203 & ~x223 & ~x226 & ~x227 & ~x228 & ~x230 & ~x255 & ~x256 & ~x283 & ~x312 & ~x337 & ~x338 & ~x365 & ~x587 & ~x616 & ~x617 & ~x618 & ~x634 & ~x635 & ~x644 & ~x662 & ~x672 & ~x674 & ~x716 & ~x743 & ~x746 & ~x770 & ~x772 & ~x775;
assign c5146 =  x537 & ~x1 & ~x17 & ~x18 & ~x20 & ~x23 & ~x27 & ~x30 & ~x31 & ~x35 & ~x36 & ~x39 & ~x40 & ~x41 & ~x42 & ~x44 & ~x45 & ~x57 & ~x59 & ~x60 & ~x61 & ~x65 & ~x84 & ~x113 & ~x115 & ~x116 & ~x118 & ~x139 & ~x144 & ~x149 & ~x152 & ~x153 & ~x167 & ~x173 & ~x174 & ~x176 & ~x177 & ~x180 & ~x201 & ~x202 & ~x203 & ~x224 & ~x235 & ~x260 & ~x261 & ~x281 & ~x282 & ~x283 & ~x286 & ~x287 & ~x288 & ~x308 & ~x311 & ~x337 & ~x342 & ~x343 & ~x364 & ~x369 & ~x423 & ~x450 & ~x478 & ~x671 & ~x732 & ~x733 & ~x734 & ~x741 & ~x743 & ~x745 & ~x748 & ~x756 & ~x760 & ~x769 & ~x771 & ~x774 & ~x775 & ~x781 & ~x783;
assign c5148 =  x220 & ~x0 & ~x2 & ~x10 & ~x18 & ~x22 & ~x27 & ~x28 & ~x29 & ~x30 & ~x31 & ~x32 & ~x34 & ~x35 & ~x41 & ~x53 & ~x54 & ~x56 & ~x57 & ~x61 & ~x62 & ~x83 & ~x85 & ~x86 & ~x87 & ~x89 & ~x91 & ~x92 & ~x93 & ~x112 & ~x115 & ~x118 & ~x119 & ~x121 & ~x131 & ~x138 & ~x139 & ~x144 & ~x146 & ~x167 & ~x170 & ~x172 & ~x175 & ~x196 & ~x197 & ~x199 & ~x200 & ~x202 & ~x204 & ~x223 & ~x224 & ~x227 & ~x229 & ~x231 & ~x252 & ~x253 & ~x255 & ~x281 & ~x283 & ~x308 & ~x336 & ~x337 & ~x365 & ~x532 & ~x560 & ~x616 & ~x619 & ~x727 & ~x744 & ~x745 & ~x746 & ~x756 & ~x769 & ~x774 & ~x775 & ~x777 & ~x778 & ~x779 & ~x783;
assign c5150 = ~x3 & ~x4 & ~x6 & ~x8 & ~x9 & ~x11 & ~x12 & ~x14 & ~x21 & ~x24 & ~x29 & ~x30 & ~x33 & ~x34 & ~x36 & ~x37 & ~x39 & ~x40 & ~x41 & ~x42 & ~x43 & ~x44 & ~x45 & ~x48 & ~x49 & ~x54 & ~x55 & ~x58 & ~x59 & ~x60 & ~x62 & ~x64 & ~x65 & ~x66 & ~x67 & ~x68 & ~x69 & ~x71 & ~x72 & ~x81 & ~x84 & ~x86 & ~x88 & ~x89 & ~x91 & ~x92 & ~x93 & ~x97 & ~x100 & ~x102 & ~x108 & ~x111 & ~x112 & ~x115 & ~x118 & ~x119 & ~x124 & ~x125 & ~x129 & ~x137 & ~x143 & ~x146 & ~x147 & ~x158 & ~x165 & ~x168 & ~x169 & ~x171 & ~x172 & ~x173 & ~x178 & ~x180 & ~x182 & ~x183 & ~x185 & ~x187 & ~x188 & ~x192 & ~x197 & ~x198 & ~x203 & ~x204 & ~x205 & ~x206 & ~x224 & ~x232 & ~x252 & ~x253 & ~x255 & ~x256 & ~x257 & ~x280 & ~x281 & ~x309 & ~x311 & ~x312 & ~x338 & ~x391 & ~x418 & ~x444 & ~x447 & ~x559 & ~x615 & ~x617 & ~x644 & ~x646 & ~x656 & ~x658 & ~x664 & ~x667 & ~x672 & ~x682 & ~x684 & ~x685 & ~x692 & ~x693 & ~x694 & ~x699 & ~x700 & ~x701 & ~x706 & ~x707 & ~x708 & ~x711 & ~x715 & ~x716 & ~x718 & ~x719 & ~x721 & ~x723 & ~x724 & ~x730 & ~x731 & ~x734 & ~x735 & ~x741 & ~x747 & ~x748 & ~x749 & ~x750 & ~x751 & ~x753 & ~x755 & ~x756 & ~x757 & ~x758 & ~x761 & ~x768 & ~x771 & ~x774 & ~x778 & ~x782;
assign c5152 =  x455 &  x537 & ~x4 & ~x20 & ~x27 & ~x38 & ~x39 & ~x40 & ~x44 & ~x51 & ~x55 & ~x72 & ~x85 & ~x97 & ~x103 & ~x116 & ~x119 & ~x121 & ~x127 & ~x136 & ~x145 & ~x147 & ~x154 & ~x177 & ~x180 & ~x196 & ~x197 & ~x203 & ~x253 & ~x263 & ~x283 & ~x336 & ~x365 & ~x478 & ~x645 & ~x700 & ~x704 & ~x709 & ~x710 & ~x712 & ~x729 & ~x732 & ~x734 & ~x751 & ~x753 & ~x776 & ~x782;
assign c5154 =  x452 &  x454 & ~x35 & ~x250 & ~x270 & ~x277 & ~x556;
assign c5156 =  x326 &  x544 &  x569 & ~x32 & ~x56 & ~x68 & ~x214 & ~x230 & ~x281 & ~x282 & ~x336 & ~x728 & ~x732 & ~x773;
assign c5158 =  x160 & ~x300;
assign c5160 =  x510 & ~x13 & ~x24 & ~x37 & ~x43 & ~x56 & ~x71 & ~x83 & ~x91 & ~x99 & ~x128 & ~x207 & ~x253 & ~x286 & ~x313 & ~x314 & ~x338 & ~x345 & ~x435 & ~x704 & ~x750 & ~x761 & ~x772;
assign c5162 =  x541 & ~x27 & ~x30 & ~x40 & ~x45 & ~x90 & ~x113 & ~x121 & ~x141 & ~x168 & ~x170 & ~x172 & ~x175 & ~x194 & ~x202 & ~x338 & ~x432 & ~x672 & ~x715 & ~x730 & ~x743 & ~x747 & ~x757 & ~x769 & ~x783;
assign c5164 =  x329 &  x332 & ~x2 & ~x5 & ~x6 & ~x9 & ~x13 & ~x14 & ~x17 & ~x18 & ~x20 & ~x22 & ~x26 & ~x27 & ~x29 & ~x30 & ~x34 & ~x35 & ~x40 & ~x44 & ~x47 & ~x50 & ~x51 & ~x53 & ~x56 & ~x73 & ~x74 & ~x79 & ~x85 & ~x89 & ~x90 & ~x95 & ~x98 & ~x100 & ~x102 & ~x103 & ~x105 & ~x109 & ~x115 & ~x126 & ~x130 & ~x137 & ~x138 & ~x139 & ~x142 & ~x145 & ~x151 & ~x156 & ~x158 & ~x164 & ~x167 & ~x169 & ~x175 & ~x177 & ~x181 & ~x182 & ~x183 & ~x184 & ~x185 & ~x190 & ~x191 & ~x204 & ~x213 & ~x214 & ~x217 & ~x227 & ~x229 & ~x241 & ~x242 & ~x244 & ~x253 & ~x255 & ~x283 & ~x308 & ~x336 & ~x363 & ~x504 & ~x559 & ~x575 & ~x587 & ~x589 & ~x593 & ~x602 & ~x608 & ~x615 & ~x620 & ~x626 & ~x629 & ~x633 & ~x636 & ~x637 & ~x638 & ~x642 & ~x648 & ~x652 & ~x660 & ~x661 & ~x663 & ~x667 & ~x668 & ~x669 & ~x670 & ~x679 & ~x680 & ~x682 & ~x686 & ~x687 & ~x693 & ~x694 & ~x702 & ~x703 & ~x707 & ~x709 & ~x710 & ~x718 & ~x720 & ~x721 & ~x722 & ~x723 & ~x724 & ~x727 & ~x735 & ~x740 & ~x742 & ~x749 & ~x751 & ~x752 & ~x756 & ~x757 & ~x766 & ~x769 & ~x770 & ~x778 & ~x780 & ~x783;
assign c5166 =  x135 & ~x13 & ~x14 & ~x19 & ~x20 & ~x32 & ~x35 & ~x57 & ~x58 & ~x61 & ~x83 & ~x85 & ~x87 & ~x90 & ~x91 & ~x112 & ~x113 & ~x114 & ~x116 & ~x117 & ~x144 & ~x167 & ~x168 & ~x169 & ~x170 & ~x172 & ~x174 & ~x195 & ~x196 & ~x201 & ~x228 & ~x229 & ~x230 & ~x231 & ~x255 & ~x256 & ~x257 & ~x310 & ~x336 & ~x337 & ~x338 & ~x364 & ~x394 & ~x395 & ~x421 & ~x450 & ~x478 & ~x616 & ~x700 & ~x756 & ~x759;
assign c5168 =  x741 &  x766 & ~x174 & ~x228 & ~x365 & ~x399 & ~x426 & ~x455;
assign c5170 = ~x6 & ~x18 & ~x65 & ~x69 & ~x91 & ~x145 & ~x152 & ~x173 & ~x205 & ~x206 & ~x228 & ~x253 & ~x255 & ~x257 & ~x261 & ~x289 & ~x380 & ~x409 & ~x422 & ~x563 & ~x582 & ~x633 & ~x635 & ~x663 & ~x688 & ~x690 & ~x693 & ~x729 & ~x742 & ~x743 & ~x759 & ~x772 & ~x782;
assign c5172 =  x397 & ~x24 & ~x42 & ~x66 & ~x69 & ~x72 & ~x84 & ~x97 & ~x104 & ~x151 & ~x177 & ~x308 & ~x390 & ~x577 & ~x641 & ~x653 & ~x696 & ~x701 & ~x737 & ~x740 & ~x773 & ~x782;
assign c5174 =  x397 &  x542 & ~x2 & ~x9 & ~x10 & ~x24 & ~x30 & ~x36 & ~x58 & ~x67 & ~x87 & ~x96 & ~x147 & ~x308 & ~x317 & ~x336 & ~x644 & ~x645 & ~x656 & ~x661 & ~x675 & ~x690 & ~x700 & ~x703 & ~x716 & ~x747 & ~x749 & ~x769 & ~x772 & ~x779;
assign c5176 = ~x1 & ~x2 & ~x8 & ~x10 & ~x11 & ~x12 & ~x13 & ~x14 & ~x15 & ~x21 & ~x25 & ~x26 & ~x32 & ~x33 & ~x35 & ~x36 & ~x38 & ~x54 & ~x55 & ~x57 & ~x59 & ~x60 & ~x62 & ~x63 & ~x84 & ~x87 & ~x89 & ~x90 & ~x91 & ~x110 & ~x112 & ~x118 & ~x140 & ~x141 & ~x142 & ~x144 & ~x145 & ~x146 & ~x147 & ~x148 & ~x151 & ~x168 & ~x169 & ~x171 & ~x174 & ~x175 & ~x176 & ~x177 & ~x196 & ~x198 & ~x199 & ~x200 & ~x201 & ~x204 & ~x205 & ~x225 & ~x226 & ~x227 & ~x228 & ~x229 & ~x230 & ~x231 & ~x232 & ~x233 & ~x234 & ~x252 & ~x253 & ~x254 & ~x256 & ~x257 & ~x258 & ~x259 & ~x261 & ~x281 & ~x282 & ~x283 & ~x285 & ~x286 & ~x287 & ~x288 & ~x289 & ~x309 & ~x313 & ~x315 & ~x316 & ~x336 & ~x338 & ~x339 & ~x342 & ~x343 & ~x344 & ~x364 & ~x366 & ~x367 & ~x368 & ~x369 & ~x392 & ~x393 & ~x394 & ~x395 & ~x404 & ~x420 & ~x421 & ~x422 & ~x424 & ~x433 & ~x449 & ~x450 & ~x728 & ~x755 & ~x756 & ~x759 & ~x771 & ~x776;
assign c5178 =  x397 &  x481 & ~x7 & ~x11 & ~x48 & ~x86 & ~x87 & ~x116 & ~x127 & ~x222 & ~x318 & ~x660 & ~x700 & ~x713 & ~x728 & ~x777;
assign c5180 =  x107 &  x134 &  x623 &  x677;
assign c5182 =  x329 &  x330 &  x331 &  x358 & ~x9 & ~x43 & ~x90 & ~x212 & ~x244 & ~x270 & ~x271 & ~x615 & ~x621 & ~x646 & ~x661 & ~x665 & ~x744;
assign c5184 =  x529 & ~x1 & ~x2 & ~x9 & ~x10 & ~x11 & ~x21 & ~x29 & ~x30 & ~x39 & ~x54 & ~x64 & ~x65 & ~x85 & ~x86 & ~x91 & ~x109 & ~x114 & ~x116 & ~x120 & ~x150 & ~x151 & ~x173 & ~x174 & ~x175 & ~x176 & ~x179 & ~x200 & ~x201 & ~x226 & ~x227 & ~x229 & ~x234 & ~x253 & ~x259 & ~x260 & ~x280 & ~x336 & ~x465 & ~x717 & ~x744 & ~x745 & ~x746 & ~x774;
assign c5186 = ~x5 & ~x13 & ~x20 & ~x30 & ~x43 & ~x69 & ~x78 & ~x87 & ~x94 & ~x113 & ~x123 & ~x126 & ~x150 & ~x200 & ~x234 & ~x259 & ~x262 & ~x364 & ~x390 & ~x417 & ~x419 & ~x559 & ~x623 & ~x627 & ~x630 & ~x635 & ~x646 & ~x676 & ~x694 & ~x700 & ~x719 & ~x727 & ~x728 & ~x739 & ~x744 & ~x746 & ~x749 & ~x774 & ~x776 & ~x782;
assign c5188 =  x443 & ~x4 & ~x6 & ~x39 & ~x42 & ~x54 & ~x56 & ~x62 & ~x70 & ~x74 & ~x87 & ~x91 & ~x97 & ~x120 & ~x196 & ~x197 & ~x203 & ~x235 & ~x281 & ~x312 & ~x340 & ~x356 & ~x450 & ~x746 & ~x747;
assign c5190 =  x218 & ~x15 & ~x17 & ~x39 & ~x62 & ~x99 & ~x128 & ~x278 & ~x705;
assign c5192 =  x523 &  x538 & ~x148 & ~x212 & ~x577 & ~x590;
assign c5194 = ~x2 & ~x5 & ~x9 & ~x25 & ~x33 & ~x41 & ~x42 & ~x54 & ~x56 & ~x60 & ~x70 & ~x72 & ~x83 & ~x118 & ~x143 & ~x145 & ~x169 & ~x201 & ~x202 & ~x205 & ~x230 & ~x232 & ~x233 & ~x259 & ~x285 & ~x354 & ~x355 & ~x504 & ~x505 & ~x508 & ~x560 & ~x634 & ~x636 & ~x689 & ~x717 & ~x770 & ~x772;
assign c5196 =  x501 & ~x1 & ~x4 & ~x7 & ~x19 & ~x26 & ~x34 & ~x35 & ~x56 & ~x60 & ~x63 & ~x84 & ~x86 & ~x87 & ~x90 & ~x92 & ~x111 & ~x117 & ~x118 & ~x140 & ~x141 & ~x143 & ~x147 & ~x169 & ~x174 & ~x228 & ~x230 & ~x231 & ~x233 & ~x252 & ~x253 & ~x256 & ~x259 & ~x281 & ~x282 & ~x283 & ~x286 & ~x289 & ~x309 & ~x312 & ~x324 & ~x337 & ~x339 & ~x340 & ~x342 & ~x368 & ~x395 & ~x559 & ~x615 & ~x643 & ~x700 & ~x755 & ~x758 & ~x760 & ~x772 & ~x783;
assign c5198 = ~x4 & ~x6 & ~x20 & ~x23 & ~x29 & ~x90 & ~x114 & ~x118 & ~x281 & ~x302 & ~x303 & ~x367 & ~x701;
assign c5200 = ~x1 & ~x2 & ~x13 & ~x28 & ~x35 & ~x37 & ~x56 & ~x60 & ~x63 & ~x85 & ~x178 & ~x226 & ~x233 & ~x256 & ~x258 & ~x259 & ~x288 & ~x312 & ~x338 & ~x394 & ~x398 & ~x448 & ~x478 & ~x489 & ~x672 & ~x759;
assign c5202 =  x454 & ~x96 & ~x350 & ~x716;
assign c5204 =  x386 & ~x0 & ~x4 & ~x12 & ~x16 & ~x17 & ~x22 & ~x28 & ~x38 & ~x57 & ~x65 & ~x66 & ~x84 & ~x166 & ~x167 & ~x170 & ~x171 & ~x195 & ~x224 & ~x225 & ~x226 & ~x228 & ~x252 & ~x285 & ~x313 & ~x337 & ~x338 & ~x365 & ~x379 & ~x393 & ~x419 & ~x420 & ~x729 & ~x755 & ~x758 & ~x760 & ~x770 & ~x772 & ~x774;
assign c5206 = ~x0 & ~x4 & ~x5 & ~x9 & ~x11 & ~x12 & ~x26 & ~x29 & ~x30 & ~x32 & ~x36 & ~x38 & ~x39 & ~x54 & ~x57 & ~x58 & ~x61 & ~x84 & ~x88 & ~x114 & ~x116 & ~x117 & ~x118 & ~x140 & ~x141 & ~x143 & ~x144 & ~x167 & ~x168 & ~x169 & ~x172 & ~x174 & ~x175 & ~x177 & ~x195 & ~x198 & ~x199 & ~x201 & ~x202 & ~x204 & ~x225 & ~x226 & ~x231 & ~x233 & ~x252 & ~x253 & ~x255 & ~x256 & ~x259 & ~x260 & ~x280 & ~x281 & ~x283 & ~x284 & ~x285 & ~x286 & ~x287 & ~x289 & ~x309 & ~x310 & ~x311 & ~x313 & ~x314 & ~x315 & ~x316 & ~x317 & ~x339 & ~x340 & ~x341 & ~x364 & ~x365 & ~x366 & ~x368 & ~x369 & ~x392 & ~x393 & ~x420 & ~x422 & ~x423 & ~x427 & ~x448 & ~x475 & ~x476 & ~x477 & ~x478 & ~x505 & ~x506 & ~x531 & ~x535 & ~x559 & ~x560 & ~x561 & ~x563 & ~x587 & ~x589 & ~x615 & ~x617 & ~x618 & ~x671 & ~x727 & ~x756 & ~x757;
assign c5208 = ~x3 & ~x10 & ~x14 & ~x21 & ~x44 & ~x49 & ~x69 & ~x70 & ~x72 & ~x73 & ~x82 & ~x96 & ~x129 & ~x146 & ~x178 & ~x200 & ~x204 & ~x207 & ~x214 & ~x227 & ~x230 & ~x233 & ~x234 & ~x308 & ~x334 & ~x362 & ~x546 & ~x553 & ~x564 & ~x570 & ~x574 & ~x578 & ~x579 & ~x602 & ~x606 & ~x608 & ~x649 & ~x684 & ~x689 & ~x713 & ~x717 & ~x718 & ~x719 & ~x732 & ~x734 & ~x736 & ~x750 & ~x763 & ~x764 & ~x769 & ~x782;
assign c5210 =  x358 &  x412 &  x482 & ~x3 & ~x5 & ~x6 & ~x7 & ~x11 & ~x12 & ~x14 & ~x15 & ~x19 & ~x28 & ~x37 & ~x38 & ~x39 & ~x41 & ~x42 & ~x43 & ~x47 & ~x50 & ~x51 & ~x55 & ~x61 & ~x62 & ~x68 & ~x73 & ~x75 & ~x80 & ~x85 & ~x89 & ~x91 & ~x92 & ~x93 & ~x94 & ~x95 & ~x96 & ~x98 & ~x99 & ~x101 & ~x103 & ~x108 & ~x111 & ~x112 & ~x120 & ~x122 & ~x123 & ~x125 & ~x130 & ~x132 & ~x133 & ~x134 & ~x135 & ~x137 & ~x141 & ~x144 & ~x145 & ~x146 & ~x154 & ~x167 & ~x175 & ~x177 & ~x178 & ~x182 & ~x184 & ~x185 & ~x186 & ~x187 & ~x189 & ~x194 & ~x195 & ~x197 & ~x200 & ~x205 & ~x209 & ~x210 & ~x214 & ~x215 & ~x230 & ~x240 & ~x241 & ~x242 & ~x250 & ~x251 & ~x280 & ~x282 & ~x284 & ~x285 & ~x286 & ~x307 & ~x310 & ~x504 & ~x574 & ~x577 & ~x578 & ~x587 & ~x588 & ~x596 & ~x598 & ~x599 & ~x602 & ~x605 & ~x606 & ~x609 & ~x610 & ~x612 & ~x613 & ~x614 & ~x615 & ~x617 & ~x620 & ~x623 & ~x628 & ~x629 & ~x639 & ~x640 & ~x641 & ~x645 & ~x650 & ~x651 & ~x653 & ~x666 & ~x672 & ~x676 & ~x679 & ~x682 & ~x684 & ~x685 & ~x687 & ~x690 & ~x697 & ~x702 & ~x704 & ~x710 & ~x714 & ~x719 & ~x723 & ~x730 & ~x734 & ~x736 & ~x737 & ~x744 & ~x752 & ~x754 & ~x757 & ~x761 & ~x762 & ~x764 & ~x765 & ~x769 & ~x771 & ~x772 & ~x774 & ~x778;
assign c5212 =  x425 & ~x43 & ~x46 & ~x47 & ~x70 & ~x74 & ~x166 & ~x169 & ~x173 & ~x283 & ~x348 & ~x660 & ~x690 & ~x704;
assign c5214 =  x427 &  x564 & ~x13 & ~x201 & ~x759;
assign c5216 =  x594 &  x595 & ~x3 & ~x13 & ~x14 & ~x21 & ~x35 & ~x60 & ~x84 & ~x118 & ~x141 & ~x142 & ~x168 & ~x172 & ~x173 & ~x195 & ~x201 & ~x226 & ~x228 & ~x252 & ~x256 & ~x257 & ~x259 & ~x260 & ~x281 & ~x284 & ~x337 & ~x338 & ~x341 & ~x342 & ~x364 & ~x368 & ~x394 & ~x420 & ~x605 & ~x671 & ~x729 & ~x774;
assign c5218 =  x679 &  x683 & ~x112 & ~x118 & ~x174 & ~x197 & ~x337 & ~x340 & ~x395 & ~x419 & ~x758;
assign c5220 =  x428 &  x566 & ~x2 & ~x7 & ~x10 & ~x16 & ~x21 & ~x37 & ~x46 & ~x58 & ~x59 & ~x89 & ~x113 & ~x121 & ~x141 & ~x168 & ~x171 & ~x176 & ~x196 & ~x199 & ~x223 & ~x228 & ~x231 & ~x252 & ~x254 & ~x259 & ~x280 & ~x281 & ~x282 & ~x283 & ~x309 & ~x313 & ~x340 & ~x365 & ~x559 & ~x701 & ~x733 & ~x734 & ~x735 & ~x743 & ~x745 & ~x747 & ~x757 & ~x763 & ~x764 & ~x767 & ~x773 & ~x779 & ~x780;
assign c5222 =  x291 & ~x10 & ~x47 & ~x72 & ~x227 & ~x229 & ~x280 & ~x337;
assign c5224 =  x331 & ~x4 & ~x32 & ~x37 & ~x40 & ~x65 & ~x91 & ~x92 & ~x96 & ~x113 & ~x147 & ~x168 & ~x197 & ~x252 & ~x255 & ~x259 & ~x281 & ~x391 & ~x416 & ~x417 & ~x702 & ~x718 & ~x719 & ~x727 & ~x744 & ~x747 & ~x770 & ~x771;
assign c5226 =  x219 & ~x13 & ~x86 & ~x140 & ~x146 & ~x169 & ~x203 & ~x225 & ~x277 & ~x281 & ~x727 & ~x774;
assign c5228 =  x697 & ~x88 & ~x197 & ~x198 & ~x200 & ~x203 & ~x225 & ~x227 & ~x312 & ~x337 & ~x341 & ~x392 & ~x394 & ~x395 & ~x421 & ~x448 & ~x776 & ~x782;
assign c5230 = ~x11 & ~x88 & ~x90 & ~x197 & ~x200 & ~x230 & ~x233 & ~x260 & ~x325 & ~x326 & ~x340 & ~x344 & ~x368 & ~x371 & ~x396 & ~x400 & ~x401 & ~x449 & ~x450 & ~x451 & ~x507 & ~x560;
assign c5232 =  x481 & ~x9 & ~x10 & ~x13 & ~x14 & ~x28 & ~x45 & ~x54 & ~x74 & ~x96 & ~x129 & ~x143 & ~x173 & ~x179 & ~x196 & ~x199 & ~x231 & ~x251 & ~x284 & ~x393 & ~x394 & ~x420 & ~x451 & ~x699 & ~x723 & ~x764 & ~x780;
assign c5234 =  x216 & ~x0 & ~x4 & ~x6 & ~x7 & ~x27 & ~x31 & ~x60 & ~x90 & ~x145 & ~x146 & ~x150 & ~x202 & ~x224 & ~x283 & ~x302 & ~x308;
assign c5236 = ~x8 & ~x15 & ~x28 & ~x30 & ~x31 & ~x38 & ~x43 & ~x167 & ~x172 & ~x204 & ~x257 & ~x259 & ~x341 & ~x349 & ~x377 & ~x393 & ~x421 & ~x642 & ~x671 & ~x762;
assign c5238 = ~x1 & ~x2 & ~x5 & ~x8 & ~x9 & ~x10 & ~x11 & ~x14 & ~x19 & ~x26 & ~x33 & ~x34 & ~x35 & ~x43 & ~x55 & ~x59 & ~x63 & ~x65 & ~x68 & ~x85 & ~x86 & ~x87 & ~x89 & ~x90 & ~x92 & ~x93 & ~x94 & ~x95 & ~x96 & ~x112 & ~x114 & ~x117 & ~x142 & ~x144 & ~x145 & ~x147 & ~x148 & ~x150 & ~x168 & ~x171 & ~x172 & ~x173 & ~x175 & ~x177 & ~x178 & ~x198 & ~x200 & ~x201 & ~x204 & ~x205 & ~x224 & ~x225 & ~x226 & ~x227 & ~x229 & ~x230 & ~x231 & ~x232 & ~x233 & ~x252 & ~x255 & ~x256 & ~x259 & ~x271 & ~x281 & ~x283 & ~x308 & ~x310 & ~x313 & ~x336 & ~x338 & ~x339 & ~x370 & ~x371 & ~x372 & ~x392 & ~x393 & ~x394 & ~x395 & ~x420 & ~x424 & ~x478 & ~x503 & ~x531 & ~x560 & ~x587 & ~x615 & ~x616 & ~x699 & ~x700 & ~x727 & ~x755 & ~x757 & ~x758;
assign c5240 =  x441 &  x584 & ~x3 & ~x6 & ~x10 & ~x27 & ~x37 & ~x62 & ~x63 & ~x64 & ~x68 & ~x94 & ~x112 & ~x117 & ~x139 & ~x141 & ~x146 & ~x175 & ~x177 & ~x202 & ~x224 & ~x280 & ~x309 & ~x310 & ~x337 & ~x378 & ~x671;
assign c5242 =  x273 & ~x1 & ~x3 & ~x4 & ~x7 & ~x14 & ~x16 & ~x20 & ~x25 & ~x30 & ~x32 & ~x34 & ~x37 & ~x42 & ~x44 & ~x55 & ~x60 & ~x63 & ~x64 & ~x66 & ~x71 & ~x81 & ~x83 & ~x84 & ~x88 & ~x97 & ~x122 & ~x142 & ~x144 & ~x147 & ~x173 & ~x175 & ~x179 & ~x198 & ~x203 & ~x226 & ~x228 & ~x254 & ~x255 & ~x256 & ~x257 & ~x281 & ~x308 & ~x309 & ~x310 & ~x311 & ~x336 & ~x337 & ~x357 & ~x691 & ~x702 & ~x719 & ~x730 & ~x743 & ~x744 & ~x749 & ~x750 & ~x752 & ~x760 & ~x766 & ~x768 & ~x776 & ~x781 & ~x783;
assign c5244 =  x538 & ~x7 & ~x14 & ~x32 & ~x39 & ~x40 & ~x43 & ~x44 & ~x45 & ~x46 & ~x47 & ~x49 & ~x55 & ~x58 & ~x66 & ~x68 & ~x70 & ~x71 & ~x87 & ~x90 & ~x99 & ~x104 & ~x114 & ~x116 & ~x124 & ~x125 & ~x126 & ~x128 & ~x139 & ~x140 & ~x146 & ~x148 & ~x173 & ~x175 & ~x180 & ~x197 & ~x199 & ~x203 & ~x223 & ~x225 & ~x229 & ~x254 & ~x257 & ~x258 & ~x259 & ~x260 & ~x280 & ~x308 & ~x310 & ~x311 & ~x316 & ~x342 & ~x343 & ~x344 & ~x394 & ~x395 & ~x396 & ~x420 & ~x421 & ~x422 & ~x478 & ~x671 & ~x717 & ~x728 & ~x729 & ~x742 & ~x744 & ~x746 & ~x770 & ~x779;
assign c5246 =  x567 & ~x0 & ~x2 & ~x3 & ~x9 & ~x13 & ~x15 & ~x25 & ~x28 & ~x30 & ~x37 & ~x40 & ~x56 & ~x64 & ~x66 & ~x67 & ~x71 & ~x84 & ~x90 & ~x92 & ~x112 & ~x118 & ~x120 & ~x125 & ~x142 & ~x145 & ~x171 & ~x176 & ~x180 & ~x202 & ~x207 & ~x209 & ~x230 & ~x255 & ~x259 & ~x287 & ~x395 & ~x449 & ~x507 & ~x531 & ~x699 & ~x759 & ~x768 & ~x777 & ~x780;
assign c5248 = ~x2 & ~x6 & ~x8 & ~x16 & ~x17 & ~x19 & ~x21 & ~x29 & ~x30 & ~x31 & ~x34 & ~x36 & ~x37 & ~x38 & ~x45 & ~x49 & ~x50 & ~x58 & ~x60 & ~x61 & ~x62 & ~x65 & ~x66 & ~x67 & ~x69 & ~x72 & ~x73 & ~x75 & ~x76 & ~x78 & ~x79 & ~x81 & ~x82 & ~x85 & ~x88 & ~x89 & ~x90 & ~x92 & ~x93 & ~x94 & ~x95 & ~x96 & ~x99 & ~x102 & ~x104 & ~x106 & ~x107 & ~x108 & ~x110 & ~x118 & ~x122 & ~x124 & ~x126 & ~x127 & ~x130 & ~x133 & ~x134 & ~x136 & ~x137 & ~x138 & ~x139 & ~x141 & ~x142 & ~x143 & ~x144 & ~x145 & ~x146 & ~x149 & ~x155 & ~x156 & ~x157 & ~x169 & ~x170 & ~x172 & ~x173 & ~x177 & ~x178 & ~x180 & ~x181 & ~x183 & ~x184 & ~x190 & ~x192 & ~x194 & ~x195 & ~x198 & ~x200 & ~x201 & ~x202 & ~x203 & ~x205 & ~x208 & ~x210 & ~x211 & ~x212 & ~x214 & ~x218 & ~x227 & ~x231 & ~x235 & ~x236 & ~x241 & ~x242 & ~x243 & ~x248 & ~x250 & ~x252 & ~x254 & ~x255 & ~x258 & ~x279 & ~x280 & ~x281 & ~x283 & ~x307 & ~x308 & ~x334 & ~x336 & ~x362 & ~x363 & ~x391 & ~x532 & ~x562 & ~x568 & ~x572 & ~x573 & ~x578 & ~x582 & ~x583 & ~x586 & ~x590 & ~x593 & ~x594 & ~x595 & ~x596 & ~x598 & ~x599 & ~x600 & ~x602 & ~x603 & ~x610 & ~x615 & ~x621 & ~x622 & ~x623 & ~x624 & ~x627 & ~x629 & ~x635 & ~x637 & ~x642 & ~x643 & ~x644 & ~x648 & ~x651 & ~x655 & ~x656 & ~x660 & ~x664 & ~x666 & ~x670 & ~x674 & ~x676 & ~x679 & ~x682 & ~x684 & ~x687 & ~x688 & ~x689 & ~x690 & ~x691 & ~x693 & ~x695 & ~x707 & ~x708 & ~x709 & ~x713 & ~x716 & ~x717 & ~x718 & ~x719 & ~x722 & ~x723 & ~x725 & ~x727 & ~x728 & ~x732 & ~x733 & ~x734 & ~x737 & ~x739 & ~x741 & ~x743 & ~x746 & ~x747 & ~x749 & ~x752 & ~x760 & ~x764 & ~x766 & ~x767 & ~x771 & ~x773 & ~x774 & ~x777 & ~x780 & ~x781 & ~x782;
assign c5250 =  x327 &  x484 &  x498 & ~x11 & ~x29 & ~x31 & ~x44 & ~x49 & ~x55 & ~x64 & ~x71 & ~x112 & ~x122 & ~x123 & ~x137 & ~x139 & ~x147 & ~x179 & ~x186 & ~x198 & ~x199 & ~x215 & ~x339 & ~x590 & ~x633 & ~x635 & ~x646 & ~x652 & ~x684 & ~x708 & ~x729 & ~x734 & ~x752 & ~x758 & ~x760 & ~x776;
assign c5252 =  x738 & ~x0 & ~x2 & ~x8 & ~x31 & ~x33 & ~x34 & ~x55 & ~x58 & ~x64 & ~x84 & ~x87 & ~x88 & ~x116 & ~x140 & ~x141 & ~x146 & ~x171 & ~x198 & ~x201 & ~x202 & ~x227 & ~x229 & ~x253 & ~x255 & ~x257 & ~x259 & ~x281 & ~x283 & ~x284 & ~x286 & ~x287 & ~x288 & ~x310 & ~x311 & ~x341 & ~x342 & ~x343 & ~x344 & ~x364 & ~x366 & ~x367 & ~x369 & ~x371 & ~x397 & ~x398 & ~x424 & ~x450 & ~x452 & ~x454 & ~x478 & ~x479 & ~x559 & ~x615 & ~x644 & ~x672 & ~x699 & ~x728;
assign c5254 =  x733 &  x734 &  x737 & ~x63 & ~x313 & ~x372 & ~x396 & ~x424 & ~x453 & ~x644;
assign c5256 = ~x3 & ~x4 & ~x6 & ~x9 & ~x14 & ~x26 & ~x28 & ~x31 & ~x36 & ~x37 & ~x38 & ~x39 & ~x40 & ~x44 & ~x55 & ~x57 & ~x60 & ~x63 & ~x65 & ~x66 & ~x67 & ~x68 & ~x87 & ~x94 & ~x96 & ~x110 & ~x123 & ~x139 & ~x173 & ~x175 & ~x176 & ~x177 & ~x195 & ~x202 & ~x203 & ~x204 & ~x205 & ~x206 & ~x230 & ~x231 & ~x234 & ~x251 & ~x261 & ~x262 & ~x305 & ~x313 & ~x336 & ~x402 & ~x404 & ~x430 & ~x504 & ~x728 & ~x757 & ~x782;
assign c5258 =  x162 &  x595 & ~x38 & ~x58 & ~x98 & ~x110 & ~x112 & ~x115 & ~x203 & ~x762 & ~x774;
assign c5260 = ~x9 & ~x37 & ~x38 & ~x39 & ~x42 & ~x89 & ~x90 & ~x93 & ~x94 & ~x113 & ~x119 & ~x139 & ~x177 & ~x202 & ~x206 & ~x224 & ~x230 & ~x256 & ~x285 & ~x313 & ~x315 & ~x317 & ~x346 & ~x424 & ~x435 & ~x449 & ~x451 & ~x463 & ~x559 & ~x756;
assign c5262 = ~x3 & ~x4 & ~x5 & ~x7 & ~x8 & ~x10 & ~x11 & ~x13 & ~x15 & ~x17 & ~x20 & ~x27 & ~x35 & ~x40 & ~x41 & ~x45 & ~x51 & ~x62 & ~x71 & ~x72 & ~x74 & ~x81 & ~x84 & ~x95 & ~x98 & ~x114 & ~x115 & ~x117 & ~x119 & ~x122 & ~x124 & ~x125 & ~x126 & ~x138 & ~x146 & ~x151 & ~x155 & ~x157 & ~x159 & ~x177 & ~x183 & ~x194 & ~x197 & ~x202 & ~x203 & ~x204 & ~x205 & ~x206 & ~x207 & ~x208 & ~x230 & ~x254 & ~x269 & ~x280 & ~x281 & ~x308 & ~x337 & ~x390 & ~x391 & ~x577 & ~x611 & ~x630 & ~x636 & ~x637 & ~x638 & ~x639 & ~x650 & ~x654 & ~x662 & ~x667 & ~x672 & ~x673 & ~x678 & ~x690 & ~x691 & ~x692 & ~x694 & ~x696 & ~x697 & ~x700 & ~x706 & ~x716 & ~x719 & ~x720 & ~x721 & ~x723 & ~x727 & ~x730 & ~x740 & ~x744 & ~x747 & ~x748 & ~x750 & ~x752 & ~x755 & ~x757 & ~x765 & ~x767 & ~x768 & ~x770 & ~x776 & ~x778 & ~x783;
assign c5264 =  x545 &  x569 & ~x5 & ~x9 & ~x11 & ~x15 & ~x19 & ~x21 & ~x23 & ~x26 & ~x28 & ~x35 & ~x40 & ~x46 & ~x47 & ~x53 & ~x62 & ~x73 & ~x76 & ~x81 & ~x83 & ~x85 & ~x86 & ~x90 & ~x92 & ~x95 & ~x96 & ~x98 & ~x99 & ~x102 & ~x104 & ~x111 & ~x113 & ~x114 & ~x116 & ~x118 & ~x121 & ~x129 & ~x131 & ~x137 & ~x142 & ~x143 & ~x146 & ~x147 & ~x149 & ~x153 & ~x205 & ~x215 & ~x227 & ~x252 & ~x254 & ~x257 & ~x258 & ~x280 & ~x282 & ~x285 & ~x286 & ~x287 & ~x313 & ~x315 & ~x340 & ~x607 & ~x616 & ~x663 & ~x666 & ~x676 & ~x689 & ~x714 & ~x715 & ~x721 & ~x727 & ~x728 & ~x733 & ~x737 & ~x742 & ~x745 & ~x747 & ~x756 & ~x763 & ~x769 & ~x770 & ~x773 & ~x774 & ~x775 & ~x781 & ~x782;
assign c5266 =  x239 &  x510 & ~x55 & ~x57 & ~x62 & ~x85 & ~x93 & ~x187 & ~x257 & ~x335 & ~x532 & ~x683 & ~x690 & ~x696 & ~x713 & ~x728 & ~x736 & ~x742 & ~x781;
assign c5268 =  x274 & ~x230 & ~x357 & ~x717;
assign c5270 = ~x0 & ~x5 & ~x6 & ~x8 & ~x16 & ~x21 & ~x22 & ~x26 & ~x31 & ~x38 & ~x39 & ~x42 & ~x44 & ~x53 & ~x54 & ~x61 & ~x64 & ~x65 & ~x67 & ~x71 & ~x84 & ~x85 & ~x91 & ~x95 & ~x96 & ~x101 & ~x110 & ~x121 & ~x124 & ~x125 & ~x126 & ~x127 & ~x135 & ~x142 & ~x143 & ~x145 & ~x146 & ~x169 & ~x173 & ~x181 & ~x185 & ~x194 & ~x196 & ~x200 & ~x212 & ~x225 & ~x228 & ~x230 & ~x233 & ~x234 & ~x237 & ~x253 & ~x259 & ~x261 & ~x336 & ~x418 & ~x419 & ~x420 & ~x632 & ~x661 & ~x664 & ~x688 & ~x700 & ~x704 & ~x706 & ~x712 & ~x716 & ~x717 & ~x720 & ~x741 & ~x747 & ~x748 & ~x751 & ~x759 & ~x773 & ~x783;
assign c5272 = ~x8 & ~x9 & ~x10 & ~x11 & ~x14 & ~x24 & ~x28 & ~x35 & ~x40 & ~x41 & ~x42 & ~x56 & ~x62 & ~x63 & ~x64 & ~x87 & ~x89 & ~x93 & ~x94 & ~x95 & ~x112 & ~x116 & ~x120 & ~x141 & ~x145 & ~x146 & ~x147 & ~x148 & ~x149 & ~x169 & ~x177 & ~x178 & ~x197 & ~x198 & ~x199 & ~x203 & ~x206 & ~x229 & ~x232 & ~x234 & ~x252 & ~x254 & ~x255 & ~x258 & ~x259 & ~x260 & ~x261 & ~x262 & ~x281 & ~x282 & ~x287 & ~x288 & ~x290 & ~x310 & ~x311 & ~x313 & ~x315 & ~x338 & ~x340 & ~x375 & ~x394 & ~x422 & ~x423 & ~x435 & ~x476 & ~x587 & ~x615 & ~x643 & ~x699 & ~x783;
assign c5274 = ~x2 & ~x6 & ~x8 & ~x9 & ~x20 & ~x26 & ~x34 & ~x35 & ~x41 & ~x44 & ~x46 & ~x52 & ~x54 & ~x56 & ~x59 & ~x62 & ~x64 & ~x66 & ~x68 & ~x73 & ~x81 & ~x82 & ~x83 & ~x85 & ~x87 & ~x88 & ~x89 & ~x111 & ~x112 & ~x114 & ~x117 & ~x118 & ~x121 & ~x141 & ~x144 & ~x145 & ~x169 & ~x197 & ~x199 & ~x201 & ~x202 & ~x206 & ~x223 & ~x225 & ~x228 & ~x229 & ~x230 & ~x233 & ~x252 & ~x253 & ~x254 & ~x256 & ~x257 & ~x258 & ~x280 & ~x282 & ~x285 & ~x286 & ~x288 & ~x311 & ~x366 & ~x394 & ~x395 & ~x475 & ~x507 & ~x525 & ~x531 & ~x552 & ~x579 & ~x580 & ~x581 & ~x588 & ~x589 & ~x591 & ~x609 & ~x644 & ~x661 & ~x663 & ~x665 & ~x690 & ~x699 & ~x716 & ~x719 & ~x720 & ~x723 & ~x727 & ~x745 & ~x747 & ~x748 & ~x749 & ~x754 & ~x759 & ~x770 & ~x771 & ~x772 & ~x774 & ~x775 & ~x776 & ~x778 & ~x781 & ~x783;
assign c5276 = ~x10 & ~x13 & ~x39 & ~x42 & ~x60 & ~x117 & ~x174 & ~x196 & ~x202 & ~x226 & ~x257 & ~x260 & ~x285 & ~x288 & ~x315 & ~x316 & ~x343 & ~x345 & ~x347 & ~x366 & ~x395 & ~x420 & ~x421 & ~x424 & ~x449 & ~x558 & ~x586 & ~x614 & ~x643;
assign c5278 =  x246 &  x539 & ~x9 & ~x13 & ~x38 & ~x76 & ~x104 & ~x106 & ~x112 & ~x122 & ~x151 & ~x171 & ~x196 & ~x199 & ~x256 & ~x278;
assign c5280 = ~x0 & ~x2 & ~x3 & ~x7 & ~x13 & ~x14 & ~x19 & ~x21 & ~x24 & ~x28 & ~x34 & ~x35 & ~x36 & ~x37 & ~x38 & ~x42 & ~x43 & ~x51 & ~x55 & ~x58 & ~x62 & ~x63 & ~x65 & ~x66 & ~x67 & ~x87 & ~x88 & ~x89 & ~x90 & ~x91 & ~x94 & ~x96 & ~x111 & ~x113 & ~x119 & ~x121 & ~x123 & ~x138 & ~x139 & ~x143 & ~x146 & ~x147 & ~x148 & ~x149 & ~x167 & ~x168 & ~x169 & ~x170 & ~x174 & ~x179 & ~x195 & ~x198 & ~x199 & ~x200 & ~x205 & ~x206 & ~x207 & ~x224 & ~x225 & ~x230 & ~x231 & ~x234 & ~x235 & ~x252 & ~x255 & ~x257 & ~x259 & ~x260 & ~x264 & ~x280 & ~x281 & ~x287 & ~x288 & ~x292 & ~x308 & ~x312 & ~x313 & ~x315 & ~x316 & ~x320 & ~x321 & ~x336 & ~x337 & ~x339 & ~x367 & ~x393 & ~x406 & ~x531 & ~x560 & ~x587 & ~x671 & ~x700 & ~x729 & ~x755 & ~x756 & ~x757 & ~x772;
assign c5282 =  x210 & ~x26 & ~x88 & ~x91 & ~x113 & ~x170 & ~x178 & ~x311 & ~x338 & ~x744 & ~x751;
assign c5284 =  x731 & ~x399;
assign c5286 =  x299 &  x300 &  x326 & ~x1 & ~x2 & ~x22 & ~x29 & ~x48 & ~x68 & ~x70 & ~x92 & ~x127 & ~x128 & ~x139 & ~x140 & ~x166 & ~x173 & ~x224 & ~x242 & ~x308 & ~x337 & ~x560 & ~x588 & ~x608 & ~x633 & ~x678 & ~x693 & ~x704 & ~x706 & ~x715 & ~x719;
assign c5288 =  x442 & ~x3 & ~x11 & ~x19 & ~x25 & ~x33 & ~x86 & ~x88 & ~x112 & ~x118 & ~x145 & ~x196 & ~x203 & ~x231 & ~x255 & ~x282 & ~x288 & ~x314 & ~x372 & ~x373 & ~x477 & ~x532 & ~x534 & ~x616 & ~x636 & ~x719 & ~x720 & ~x757;
assign c5290 =  x511 & ~x5 & ~x15 & ~x19 & ~x29 & ~x38 & ~x48 & ~x53 & ~x58 & ~x63 & ~x74 & ~x80 & ~x98 & ~x99 & ~x100 & ~x110 & ~x114 & ~x115 & ~x122 & ~x130 & ~x131 & ~x140 & ~x141 & ~x142 & ~x146 & ~x147 & ~x149 & ~x150 & ~x156 & ~x170 & ~x171 & ~x174 & ~x195 & ~x201 & ~x203 & ~x206 & ~x222 & ~x227 & ~x229 & ~x232 & ~x254 & ~x261 & ~x282 & ~x283 & ~x288 & ~x309 & ~x310 & ~x311 & ~x366 & ~x392 & ~x420 & ~x478 & ~x672 & ~x714 & ~x720 & ~x724 & ~x727 & ~x728 & ~x733 & ~x734 & ~x747 & ~x750 & ~x751 & ~x752 & ~x760 & ~x762 & ~x764 & ~x766 & ~x770 & ~x773;
assign c5292 =  x454 & ~x33 & ~x43 & ~x149 & ~x161 & ~x179 & ~x201 & ~x394 & ~x403 & ~x644 & ~x726 & ~x738 & ~x758 & ~x759 & ~x778;
assign c5294 =  x482 &  x601 & ~x32 & ~x50 & ~x57 & ~x65 & ~x73 & ~x168 & ~x170 & ~x174 & ~x196 & ~x197 & ~x256 & ~x258 & ~x285 & ~x364 & ~x368 & ~x700 & ~x743 & ~x764 & ~x780 & ~x783;
assign c5296 =  x160 & ~x2 & ~x21 & ~x62 & ~x122 & ~x175 & ~x310 & ~x315 & ~x778;
assign c5298 =  x264 & ~x4 & ~x28 & ~x29 & ~x37 & ~x40 & ~x48 & ~x52 & ~x115 & ~x142 & ~x149 & ~x175 & ~x199 & ~x201 & ~x233 & ~x587 & ~x671 & ~x730 & ~x736 & ~x765;
assign c5300 =  x455 & ~x23 & ~x37 & ~x38 & ~x41 & ~x42 & ~x47 & ~x54 & ~x70 & ~x71 & ~x82 & ~x86 & ~x223 & ~x226 & ~x281 & ~x297 & ~x334 & ~x476 & ~x691 & ~x709 & ~x758 & ~x772;
assign c5302 =  x529 & ~x7 & ~x12 & ~x26 & ~x30 & ~x31 & ~x36 & ~x56 & ~x63 & ~x91 & ~x114 & ~x145 & ~x150 & ~x175 & ~x178 & ~x203 & ~x225 & ~x254 & ~x309 & ~x312 & ~x336 & ~x465 & ~x504 & ~x767 & ~x768 & ~x773;
assign c5304 = ~x2 & ~x3 & ~x5 & ~x8 & ~x14 & ~x27 & ~x36 & ~x38 & ~x39 & ~x53 & ~x55 & ~x57 & ~x58 & ~x61 & ~x62 & ~x83 & ~x84 & ~x87 & ~x89 & ~x113 & ~x116 & ~x119 & ~x120 & ~x139 & ~x148 & ~x168 & ~x171 & ~x177 & ~x200 & ~x203 & ~x229 & ~x232 & ~x252 & ~x254 & ~x258 & ~x259 & ~x280 & ~x282 & ~x288 & ~x314 & ~x340 & ~x342 & ~x368 & ~x370 & ~x393 & ~x394 & ~x395 & ~x421 & ~x449 & ~x451 & ~x478 & ~x504 & ~x552 & ~x560 & ~x561 & ~x562 & ~x579 & ~x606 & ~x607 & ~x662 & ~x671 & ~x719 & ~x727 & ~x743 & ~x746 & ~x770 & ~x772 & ~x774;
assign c5306 =  x399 & ~x1 & ~x6 & ~x15 & ~x30 & ~x38 & ~x40 & ~x41 & ~x43 & ~x44 & ~x47 & ~x71 & ~x96 & ~x99 & ~x101 & ~x103 & ~x117 & ~x143 & ~x148 & ~x171 & ~x172 & ~x228 & ~x245 & ~x269 & ~x270 & ~x272 & ~x275 & ~x391 & ~x504 & ~x563 & ~x564 & ~x565 & ~x567 & ~x575 & ~x587 & ~x589 & ~x596 & ~x602 & ~x649 & ~x650 & ~x654 & ~x658 & ~x668 & ~x720 & ~x721 & ~x738 & ~x739 & ~x760 & ~x769;
assign c5308 =  x329 &  x489 & ~x149 & ~x203 & ~x242 & ~x270 & ~x318 & ~x717;
assign c5310 = ~x0 & ~x1 & ~x3 & ~x32 & ~x33 & ~x34 & ~x35 & ~x36 & ~x40 & ~x41 & ~x42 & ~x43 & ~x46 & ~x49 & ~x50 & ~x56 & ~x65 & ~x66 & ~x68 & ~x69 & ~x71 & ~x78 & ~x84 & ~x89 & ~x91 & ~x93 & ~x95 & ~x96 & ~x97 & ~x98 & ~x100 & ~x104 & ~x111 & ~x112 & ~x119 & ~x121 & ~x124 & ~x126 & ~x151 & ~x163 & ~x168 & ~x174 & ~x180 & ~x197 & ~x216 & ~x223 & ~x228 & ~x230 & ~x233 & ~x261 & ~x280 & ~x336 & ~x362 & ~x389 & ~x390 & ~x391 & ~x504 & ~x532 & ~x573 & ~x579 & ~x583 & ~x584 & ~x587 & ~x588 & ~x620 & ~x623 & ~x626 & ~x629 & ~x647 & ~x653 & ~x666 & ~x667 & ~x671 & ~x701 & ~x707 & ~x716 & ~x720 & ~x725 & ~x735 & ~x742 & ~x744 & ~x749 & ~x768 & ~x771 & ~x783;
assign c5312 =  x237 &  x443 & ~x1 & ~x38 & ~x65 & ~x144 & ~x308 & ~x448 & ~x775;
assign c5314 =  x537 &  x581 &  x584 & ~x14 & ~x66 & ~x112 & ~x183 & ~x195 & ~x210 & ~x236 & ~x261 & ~x281 & ~x309 & ~x649 & ~x679 & ~x762 & ~x776;
assign c5316 = ~x2 & ~x3 & ~x5 & ~x6 & ~x10 & ~x59 & ~x61 & ~x62 & ~x112 & ~x116 & ~x119 & ~x141 & ~x145 & ~x168 & ~x172 & ~x174 & ~x175 & ~x196 & ~x199 & ~x200 & ~x202 & ~x225 & ~x226 & ~x229 & ~x230 & ~x231 & ~x255 & ~x257 & ~x258 & ~x260 & ~x281 & ~x282 & ~x284 & ~x286 & ~x287 & ~x288 & ~x314 & ~x316 & ~x336 & ~x338 & ~x339 & ~x341 & ~x365 & ~x366 & ~x367 & ~x392 & ~x394 & ~x395 & ~x396 & ~x421 & ~x423 & ~x426 & ~x505 & ~x506 & ~x562 & ~x607 & ~x635 & ~x662 & ~x663 & ~x689 & ~x690 & ~x692 & ~x744 & ~x745 & ~x755 & ~x772 & ~x776 & ~x778;
assign c5318 =  x211 & ~x12 & ~x38 & ~x51 & ~x94 & ~x116 & ~x122 & ~x197 & ~x224 & ~x253 & ~x254 & ~x259 & ~x311 & ~x316 & ~x534 & ~x559 & ~x560 & ~x617 & ~x643;
assign c5320 = ~x1 & ~x8 & ~x13 & ~x26 & ~x32 & ~x39 & ~x40 & ~x41 & ~x43 & ~x47 & ~x59 & ~x70 & ~x72 & ~x94 & ~x95 & ~x96 & ~x102 & ~x121 & ~x122 & ~x123 & ~x134 & ~x145 & ~x146 & ~x155 & ~x169 & ~x173 & ~x177 & ~x179 & ~x205 & ~x207 & ~x208 & ~x280 & ~x307 & ~x333 & ~x334 & ~x335 & ~x362 & ~x387 & ~x388 & ~x617 & ~x664 & ~x666 & ~x671 & ~x756 & ~x777;
assign c5322 =  x511 & ~x6 & ~x11 & ~x13 & ~x22 & ~x23 & ~x34 & ~x35 & ~x46 & ~x57 & ~x59 & ~x60 & ~x66 & ~x67 & ~x70 & ~x81 & ~x115 & ~x116 & ~x139 & ~x174 & ~x197 & ~x202 & ~x423 & ~x460 & ~x743 & ~x756 & ~x760 & ~x764 & ~x771 & ~x775 & ~x778;
assign c5324 =  x271 & ~x7 & ~x10 & ~x12 & ~x58 & ~x63 & ~x82 & ~x84 & ~x91 & ~x95 & ~x111 & ~x116 & ~x120 & ~x144 & ~x145 & ~x147 & ~x148 & ~x176 & ~x196 & ~x199 & ~x224 & ~x254 & ~x256 & ~x357 & ~x782;
assign c5326 =  x361 & ~x110 & ~x150 & ~x319 & ~x445 & ~x649 & ~x755;
assign c5328 =  x470 &  x526 & ~x0 & ~x3 & ~x5 & ~x6 & ~x14 & ~x30 & ~x42 & ~x45 & ~x84 & ~x97 & ~x112 & ~x118 & ~x124 & ~x139 & ~x142 & ~x206 & ~x230 & ~x231 & ~x288 & ~x291 & ~x315 & ~x672 & ~x703 & ~x719 & ~x742 & ~x764;
assign c5330 =  x453 &  x537 &  x539 & ~x8 & ~x12 & ~x31 & ~x32 & ~x68 & ~x81 & ~x82 & ~x85 & ~x118 & ~x125 & ~x144 & ~x145 & ~x154 & ~x167 & ~x205 & ~x227 & ~x259 & ~x262 & ~x364 & ~x365 & ~x709 & ~x711 & ~x714 & ~x723 & ~x728 & ~x743 & ~x753 & ~x779 & ~x782;
assign c5332 =  x686 & ~x7 & ~x8 & ~x28 & ~x84 & ~x284 & ~x288 & ~x344 & ~x371 & ~x372 & ~x397 & ~x399 & ~x424 & ~x428 & ~x452 & ~x477 & ~x479 & ~x563 & ~x590 & ~x619 & ~x644 & ~x646 & ~x772;
assign c5334 = ~x2 & ~x7 & ~x10 & ~x16 & ~x22 & ~x27 & ~x28 & ~x31 & ~x34 & ~x36 & ~x37 & ~x40 & ~x42 & ~x43 & ~x44 & ~x84 & ~x90 & ~x111 & ~x117 & ~x120 & ~x146 & ~x148 & ~x171 & ~x175 & ~x176 & ~x196 & ~x200 & ~x227 & ~x230 & ~x231 & ~x233 & ~x254 & ~x258 & ~x259 & ~x280 & ~x353 & ~x476 & ~x504 & ~x523 & ~x524 & ~x525 & ~x552 & ~x553 & ~x580 & ~x688 & ~x689 & ~x690 & ~x743 & ~x761 & ~x769 & ~x770;
assign c5336 =  x435 & ~x30 & ~x36 & ~x89 & ~x233 & ~x258 & ~x306 & ~x332 & ~x333 & ~x551 & ~x588 & ~x716;
assign c5338 =  x732 & ~x231 & ~x281 & ~x342 & ~x344 & ~x396 & ~x426 & ~x427 & ~x534;
assign c5340 = ~x9 & ~x13 & ~x89 & ~x112 & ~x118 & ~x145 & ~x146 & ~x167 & ~x177 & ~x205 & ~x223 & ~x259 & ~x260 & ~x280 & ~x288 & ~x319 & ~x321 & ~x322 & ~x336 & ~x348 & ~x373 & ~x375 & ~x398 & ~x434 & ~x435 & ~x452 & ~x700;
assign c5342 =  x105 & ~x3 & ~x90 & ~x174 & ~x199 & ~x200 & ~x202 & ~x252 & ~x342 & ~x365 & ~x371 & ~x534 & ~x616 & ~x617;
assign c5344 = ~x4 & ~x10 & ~x13 & ~x14 & ~x16 & ~x28 & ~x30 & ~x42 & ~x43 & ~x55 & ~x61 & ~x67 & ~x69 & ~x85 & ~x89 & ~x109 & ~x110 & ~x113 & ~x114 & ~x115 & ~x116 & ~x117 & ~x139 & ~x145 & ~x147 & ~x150 & ~x152 & ~x173 & ~x174 & ~x176 & ~x178 & ~x179 & ~x185 & ~x202 & ~x209 & ~x225 & ~x282 & ~x287 & ~x288 & ~x338 & ~x364 & ~x365 & ~x367 & ~x393 & ~x394 & ~x422 & ~x448 & ~x451 & ~x478 & ~x479 & ~x506 & ~x507 & ~x699 & ~x700 & ~x727 & ~x755 & ~x770 & ~x783;
assign c5346 =  x679 & ~x8 & ~x26 & ~x82 & ~x115 & ~x116 & ~x170 & ~x196 & ~x258 & ~x311 & ~x336 & ~x341 & ~x343 & ~x606 & ~x634 & ~x635 & ~x716 & ~x718 & ~x770;
assign c5348 =  x362 &  x622 & ~x69 & ~x144 & ~x254 & ~x342;
assign c5350 =  x328 & ~x12 & ~x20 & ~x21 & ~x24 & ~x33 & ~x34 & ~x35 & ~x53 & ~x64 & ~x70 & ~x74 & ~x91 & ~x92 & ~x103 & ~x112 & ~x113 & ~x161 & ~x170 & ~x172 & ~x173 & ~x177 & ~x179 & ~x185 & ~x188 & ~x201 & ~x208 & ~x213 & ~x216 & ~x224 & ~x226 & ~x261 & ~x283 & ~x290 & ~x318 & ~x366 & ~x367 & ~x448 & ~x587 & ~x588 & ~x614 & ~x618 & ~x635 & ~x644 & ~x653 & ~x665 & ~x672 & ~x674 & ~x684 & ~x686 & ~x687 & ~x717 & ~x718 & ~x730 & ~x737 & ~x743 & ~x755 & ~x757 & ~x761 & ~x762 & ~x771 & ~x773 & ~x776 & ~x778;
assign c5352 =  x444 & ~x9 & ~x11 & ~x35 & ~x86 & ~x110 & ~x112 & ~x116 & ~x147 & ~x148 & ~x150 & ~x177 & ~x198 & ~x228 & ~x252 & ~x282 & ~x285 & ~x312 & ~x314 & ~x351 & ~x366 & ~x380 & ~x773 & ~x776;
assign c5354 =  x764;
assign c5356 = ~x1 & ~x4 & ~x12 & ~x14 & ~x15 & ~x16 & ~x18 & ~x24 & ~x29 & ~x39 & ~x40 & ~x41 & ~x42 & ~x43 & ~x45 & ~x46 & ~x49 & ~x50 & ~x52 & ~x55 & ~x65 & ~x66 & ~x67 & ~x68 & ~x69 & ~x70 & ~x71 & ~x72 & ~x74 & ~x75 & ~x82 & ~x89 & ~x91 & ~x92 & ~x94 & ~x95 & ~x97 & ~x98 & ~x99 & ~x101 & ~x102 & ~x104 & ~x105 & ~x114 & ~x121 & ~x122 & ~x125 & ~x128 & ~x130 & ~x131 & ~x133 & ~x134 & ~x139 & ~x140 & ~x142 & ~x144 & ~x145 & ~x146 & ~x149 & ~x150 & ~x152 & ~x159 & ~x166 & ~x169 & ~x172 & ~x176 & ~x184 & ~x185 & ~x194 & ~x196 & ~x197 & ~x200 & ~x201 & ~x203 & ~x207 & ~x209 & ~x216 & ~x224 & ~x227 & ~x229 & ~x230 & ~x234 & ~x253 & ~x255 & ~x257 & ~x259 & ~x281 & ~x283 & ~x284 & ~x308 & ~x309 & ~x336 & ~x337 & ~x390 & ~x417 & ~x418 & ~x419 & ~x504 & ~x532 & ~x560 & ~x604 & ~x628 & ~x633 & ~x645 & ~x658 & ~x662 & ~x664 & ~x669 & ~x676 & ~x684 & ~x686 & ~x690 & ~x691 & ~x692 & ~x700 & ~x702 & ~x703 & ~x704 & ~x706 & ~x707 & ~x708 & ~x710 & ~x711 & ~x713 & ~x714 & ~x716 & ~x717 & ~x719 & ~x728 & ~x730 & ~x733 & ~x738 & ~x747 & ~x751 & ~x754 & ~x759 & ~x761 & ~x763 & ~x770 & ~x771 & ~x774 & ~x776 & ~x777 & ~x780 & ~x782;
assign c5358 = ~x0 & ~x2 & ~x3 & ~x4 & ~x5 & ~x6 & ~x7 & ~x8 & ~x9 & ~x10 & ~x11 & ~x12 & ~x13 & ~x14 & ~x17 & ~x21 & ~x23 & ~x24 & ~x25 & ~x26 & ~x29 & ~x30 & ~x31 & ~x32 & ~x33 & ~x34 & ~x36 & ~x37 & ~x38 & ~x39 & ~x40 & ~x41 & ~x51 & ~x54 & ~x55 & ~x56 & ~x58 & ~x60 & ~x61 & ~x62 & ~x63 & ~x64 & ~x83 & ~x84 & ~x85 & ~x86 & ~x87 & ~x88 & ~x89 & ~x93 & ~x112 & ~x113 & ~x114 & ~x115 & ~x116 & ~x117 & ~x118 & ~x120 & ~x142 & ~x143 & ~x144 & ~x145 & ~x146 & ~x147 & ~x149 & ~x168 & ~x169 & ~x170 & ~x172 & ~x173 & ~x175 & ~x176 & ~x177 & ~x194 & ~x195 & ~x197 & ~x198 & ~x202 & ~x204 & ~x205 & ~x224 & ~x225 & ~x226 & ~x227 & ~x228 & ~x229 & ~x230 & ~x231 & ~x232 & ~x253 & ~x255 & ~x256 & ~x258 & ~x260 & ~x280 & ~x281 & ~x282 & ~x283 & ~x286 & ~x287 & ~x288 & ~x308 & ~x309 & ~x310 & ~x313 & ~x323 & ~x336 & ~x337 & ~x340 & ~x364 & ~x365 & ~x366 & ~x367 & ~x368 & ~x369 & ~x392 & ~x393 & ~x394 & ~x395 & ~x448 & ~x475 & ~x503 & ~x615 & ~x643 & ~x699 & ~x727 & ~x729 & ~x755 & ~x756 & ~x757 & ~x759 & ~x771 & ~x772 & ~x782 & ~x783;
assign c5360 = ~x2 & ~x6 & ~x12 & ~x14 & ~x16 & ~x19 & ~x20 & ~x21 & ~x24 & ~x26 & ~x27 & ~x29 & ~x31 & ~x37 & ~x38 & ~x42 & ~x43 & ~x46 & ~x56 & ~x63 & ~x64 & ~x65 & ~x67 & ~x74 & ~x76 & ~x78 & ~x82 & ~x88 & ~x89 & ~x91 & ~x92 & ~x99 & ~x100 & ~x101 & ~x110 & ~x111 & ~x113 & ~x118 & ~x120 & ~x122 & ~x126 & ~x132 & ~x133 & ~x134 & ~x135 & ~x140 & ~x143 & ~x144 & ~x149 & ~x151 & ~x155 & ~x166 & ~x171 & ~x174 & ~x175 & ~x178 & ~x187 & ~x188 & ~x190 & ~x196 & ~x197 & ~x198 & ~x199 & ~x200 & ~x201 & ~x204 & ~x205 & ~x207 & ~x209 & ~x211 & ~x212 & ~x213 & ~x214 & ~x215 & ~x220 & ~x223 & ~x224 & ~x226 & ~x231 & ~x234 & ~x241 & ~x242 & ~x243 & ~x252 & ~x254 & ~x260 & ~x270 & ~x278 & ~x280 & ~x282 & ~x283 & ~x308 & ~x309 & ~x362 & ~x391 & ~x532 & ~x559 & ~x560 & ~x562 & ~x566 & ~x574 & ~x575 & ~x578 & ~x579 & ~x587 & ~x592 & ~x608 & ~x616 & ~x628 & ~x629 & ~x631 & ~x637 & ~x638 & ~x641 & ~x652 & ~x654 & ~x660 & ~x661 & ~x662 & ~x663 & ~x666 & ~x669 & ~x671 & ~x672 & ~x674 & ~x676 & ~x678 & ~x682 & ~x683 & ~x686 & ~x688 & ~x692 & ~x699 & ~x700 & ~x702 & ~x703 & ~x709 & ~x711 & ~x712 & ~x714 & ~x723 & ~x728 & ~x729 & ~x733 & ~x737 & ~x738 & ~x740 & ~x746 & ~x747 & ~x750 & ~x761 & ~x763 & ~x767 & ~x768 & ~x769 & ~x771 & ~x772 & ~x775 & ~x777 & ~x781;
assign c5362 =  x483 &  x537 &  x566 & ~x1 & ~x5 & ~x9 & ~x14 & ~x30 & ~x38 & ~x43 & ~x45 & ~x60 & ~x61 & ~x71 & ~x83 & ~x89 & ~x97 & ~x99 & ~x101 & ~x126 & ~x128 & ~x146 & ~x167 & ~x172 & ~x173 & ~x175 & ~x198 & ~x202 & ~x282 & ~x286 & ~x309 & ~x312 & ~x337 & ~x730 & ~x739 & ~x741 & ~x742 & ~x750 & ~x757 & ~x760 & ~x763 & ~x768 & ~x772;
assign c5364 =  x332 &  x357 &  x358 &  x359 &  x360 &  x453 & ~x2 & ~x17 & ~x19 & ~x21 & ~x30 & ~x34 & ~x36 & ~x51 & ~x72 & ~x79 & ~x89 & ~x111 & ~x134 & ~x141 & ~x150 & ~x163 & ~x169 & ~x173 & ~x198 & ~x208 & ~x224 & ~x230 & ~x234 & ~x241 & ~x242 & ~x243 & ~x248 & ~x254 & ~x289 & ~x290 & ~x310 & ~x313 & ~x318 & ~x575 & ~x577 & ~x596 & ~x599 & ~x631 & ~x633 & ~x641 & ~x646 & ~x692 & ~x704 & ~x718 & ~x722 & ~x728 & ~x748 & ~x757 & ~x763 & ~x768 & ~x770;
assign c5366 = ~x13 & ~x14 & ~x17 & ~x27 & ~x30 & ~x33 & ~x35 & ~x38 & ~x42 & ~x43 & ~x58 & ~x66 & ~x68 & ~x69 & ~x71 & ~x84 & ~x87 & ~x89 & ~x90 & ~x93 & ~x95 & ~x98 & ~x118 & ~x120 & ~x140 & ~x141 & ~x144 & ~x172 & ~x174 & ~x197 & ~x198 & ~x226 & ~x227 & ~x229 & ~x231 & ~x232 & ~x258 & ~x280 & ~x281 & ~x284 & ~x285 & ~x286 & ~x312 & ~x326 & ~x337 & ~x354 & ~x355 & ~x365 & ~x367 & ~x476 & ~x504 & ~x505 & ~x506 & ~x643 & ~x700 & ~x744 & ~x745 & ~x761 & ~x770;
assign c5368 =  x639 & ~x15 & ~x29 & ~x31 & ~x33 & ~x35 & ~x56 & ~x83 & ~x91 & ~x146 & ~x173 & ~x175 & ~x196 & ~x226 & ~x232 & ~x260 & ~x262 & ~x280 & ~x296 & ~x314 & ~x345 & ~x367 & ~x392 & ~x398 & ~x756 & ~x758;
assign c5370 =  x382 &  x440 &  x481 &  x494 &  x495 &  x512 & ~x2 & ~x8 & ~x11 & ~x12 & ~x14 & ~x15 & ~x22 & ~x23 & ~x34 & ~x37 & ~x40 & ~x55 & ~x56 & ~x57 & ~x59 & ~x70 & ~x85 & ~x90 & ~x91 & ~x101 & ~x108 & ~x112 & ~x114 & ~x116 & ~x121 & ~x123 & ~x125 & ~x144 & ~x146 & ~x157 & ~x174 & ~x176 & ~x195 & ~x200 & ~x206 & ~x214 & ~x223 & ~x232 & ~x256 & ~x281 & ~x335 & ~x587 & ~x638 & ~x644 & ~x647 & ~x671 & ~x672 & ~x685 & ~x691 & ~x692 & ~x694 & ~x700 & ~x701 & ~x702 & ~x706 & ~x716 & ~x719 & ~x724 & ~x727 & ~x732 & ~x734 & ~x738 & ~x742 & ~x743 & ~x746 & ~x751 & ~x753 & ~x756 & ~x771 & ~x777 & ~x782;
assign c5372 =  x398 &  x483 &  x525 & ~x5 & ~x19 & ~x69 & ~x93 & ~x101 & ~x213 & ~x241 & ~x391 & ~x615 & ~x711 & ~x747;
assign c5374 =  x426 & ~x15 & ~x26 & ~x58 & ~x67 & ~x77 & ~x104 & ~x146 & ~x147 & ~x176 & ~x319 & ~x349 & ~x587 & ~x670 & ~x686 & ~x769;
assign c5376 = ~x7 & ~x8 & ~x13 & ~x39 & ~x47 & ~x48 & ~x55 & ~x69 & ~x84 & ~x91 & ~x93 & ~x95 & ~x108 & ~x118 & ~x124 & ~x140 & ~x142 & ~x174 & ~x175 & ~x182 & ~x183 & ~x201 & ~x234 & ~x253 & ~x268 & ~x271 & ~x281 & ~x297 & ~x298 & ~x309 & ~x310 & ~x547 & ~x563 & ~x564 & ~x566 & ~x568 & ~x571 & ~x582 & ~x588 & ~x591 & ~x593 & ~x610 & ~x633 & ~x634 & ~x643 & ~x657 & ~x671 & ~x699 & ~x717 & ~x722 & ~x728 & ~x742 & ~x782;
assign c5378 =  x593 &  x598 & ~x19 & ~x39 & ~x55 & ~x127 & ~x252 & ~x280 & ~x312 & ~x340 & ~x341 & ~x759;
assign c5380 =  x557 & ~x3 & ~x5 & ~x8 & ~x10 & ~x11 & ~x115 & ~x116 & ~x144 & ~x168 & ~x172 & ~x200 & ~x201 & ~x202 & ~x256 & ~x364 & ~x368 & ~x394 & ~x476 & ~x478 & ~x497 & ~x506 & ~x757 & ~x782;
assign c5382 =  x423 &  x432 &  x438 & ~x43 & ~x242 & ~x269 & ~x713;
assign c5384 = ~x0 & ~x2 & ~x13 & ~x29 & ~x31 & ~x41 & ~x57 & ~x65 & ~x71 & ~x88 & ~x90 & ~x124 & ~x126 & ~x137 & ~x142 & ~x143 & ~x145 & ~x150 & ~x151 & ~x157 & ~x169 & ~x171 & ~x175 & ~x177 & ~x179 & ~x182 & ~x199 & ~x203 & ~x206 & ~x208 & ~x215 & ~x224 & ~x230 & ~x231 & ~x232 & ~x233 & ~x250 & ~x254 & ~x279 & ~x390 & ~x391 & ~x417 & ~x418 & ~x419 & ~x532 & ~x583 & ~x608 & ~x688 & ~x711 & ~x722 & ~x724 & ~x725 & ~x749 & ~x753 & ~x757 & ~x761 & ~x764;
assign c5386 =  x400 &  x534 &  x546 & ~x61 & ~x67 & ~x83 & ~x206 & ~x750 & ~x782;
assign c5388 = ~x44 & ~x69 & ~x99 & ~x102 & ~x282 & ~x309 & ~x665 & ~x690;
assign c5390 =  x738 & ~x552;
assign c5392 =  x266 &  x495 & ~x14 & ~x17 & ~x19 & ~x24 & ~x38 & ~x45 & ~x52 & ~x54 & ~x58 & ~x63 & ~x65 & ~x67 & ~x70 & ~x77 & ~x97 & ~x99 & ~x106 & ~x110 & ~x112 & ~x115 & ~x124 & ~x128 & ~x132 & ~x133 & ~x156 & ~x158 & ~x176 & ~x179 & ~x191 & ~x197 & ~x214 & ~x215 & ~x229 & ~x232 & ~x253 & ~x256 & ~x257 & ~x259 & ~x260 & ~x290 & ~x291 & ~x532 & ~x615 & ~x655 & ~x664 & ~x681 & ~x685 & ~x687 & ~x703 & ~x713 & ~x718 & ~x731 & ~x732 & ~x737 & ~x738 & ~x741 & ~x745 & ~x748 & ~x755 & ~x758 & ~x767 & ~x773 & ~x775 & ~x782;
assign c5394 = ~x8 & ~x21 & ~x29 & ~x33 & ~x41 & ~x45 & ~x56 & ~x57 & ~x58 & ~x60 & ~x64 & ~x68 & ~x84 & ~x88 & ~x94 & ~x97 & ~x98 & ~x105 & ~x116 & ~x146 & ~x148 & ~x151 & ~x178 & ~x200 & ~x209 & ~x223 & ~x226 & ~x233 & ~x279 & ~x280 & ~x418 & ~x445 & ~x564 & ~x575 & ~x616 & ~x623 & ~x625 & ~x636 & ~x646 & ~x649 & ~x650 & ~x665 & ~x666 & ~x669 & ~x681 & ~x690 & ~x694 & ~x700 & ~x706 & ~x714 & ~x781;
assign c5396 =  x237 & ~x8 & ~x14 & ~x22 & ~x24 & ~x72 & ~x81 & ~x111 & ~x141 & ~x147 & ~x148 & ~x172 & ~x196 & ~x225 & ~x226 & ~x282 & ~x364 & ~x689 & ~x730 & ~x747 & ~x770 & ~x775;
assign c5398 =  x481 & ~x7 & ~x20 & ~x84 & ~x104 & ~x123 & ~x149 & ~x196 & ~x202 & ~x444 & ~x615 & ~x649 & ~x695 & ~x702 & ~x744 & ~x750 & ~x761;
assign c5400 =  x510 & ~x9 & ~x16 & ~x25 & ~x43 & ~x65 & ~x82 & ~x83 & ~x87 & ~x120 & ~x145 & ~x148 & ~x197 & ~x198 & ~x224 & ~x226 & ~x252 & ~x256 & ~x257 & ~x280 & ~x283 & ~x284 & ~x309 & ~x337 & ~x394 & ~x423 & ~x477 & ~x691 & ~x692 & ~x717 & ~x721 & ~x722 & ~x734 & ~x747 & ~x751 & ~x758 & ~x774;
assign c5402 = ~x2 & ~x4 & ~x8 & ~x10 & ~x11 & ~x12 & ~x13 & ~x31 & ~x33 & ~x35 & ~x63 & ~x86 & ~x87 & ~x89 & ~x112 & ~x117 & ~x140 & ~x142 & ~x143 & ~x147 & ~x150 & ~x169 & ~x173 & ~x175 & ~x176 & ~x200 & ~x204 & ~x205 & ~x206 & ~x227 & ~x228 & ~x231 & ~x232 & ~x260 & ~x280 & ~x281 & ~x283 & ~x287 & ~x288 & ~x295 & ~x296 & ~x297 & ~x309 & ~x310 & ~x311 & ~x313 & ~x314 & ~x324 & ~x325 & ~x336 & ~x339 & ~x340 & ~x448 & ~x477 & ~x478 & ~x503 & ~x643 & ~x671 & ~x699 & ~x744 & ~x772 & ~x775;
assign c5404 =  x300 & ~x0 & ~x3 & ~x4 & ~x5 & ~x6 & ~x8 & ~x9 & ~x10 & ~x11 & ~x12 & ~x13 & ~x15 & ~x16 & ~x17 & ~x18 & ~x21 & ~x23 & ~x24 & ~x25 & ~x26 & ~x28 & ~x29 & ~x32 & ~x33 & ~x34 & ~x35 & ~x37 & ~x38 & ~x41 & ~x42 & ~x43 & ~x45 & ~x46 & ~x50 & ~x51 & ~x52 & ~x53 & ~x55 & ~x56 & ~x57 & ~x61 & ~x64 & ~x68 & ~x69 & ~x70 & ~x75 & ~x80 & ~x82 & ~x83 & ~x88 & ~x89 & ~x90 & ~x91 & ~x92 & ~x93 & ~x94 & ~x95 & ~x96 & ~x98 & ~x100 & ~x105 & ~x110 & ~x112 & ~x115 & ~x116 & ~x117 & ~x119 & ~x120 & ~x123 & ~x124 & ~x125 & ~x128 & ~x129 & ~x138 & ~x139 & ~x140 & ~x143 & ~x144 & ~x145 & ~x147 & ~x150 & ~x151 & ~x157 & ~x158 & ~x159 & ~x170 & ~x171 & ~x173 & ~x175 & ~x177 & ~x178 & ~x179 & ~x187 & ~x194 & ~x196 & ~x197 & ~x199 & ~x201 & ~x203 & ~x204 & ~x206 & ~x214 & ~x215 & ~x222 & ~x224 & ~x225 & ~x228 & ~x229 & ~x232 & ~x233 & ~x234 & ~x253 & ~x255 & ~x256 & ~x257 & ~x259 & ~x262 & ~x280 & ~x281 & ~x282 & ~x283 & ~x284 & ~x287 & ~x309 & ~x310 & ~x311 & ~x312 & ~x336 & ~x338 & ~x340 & ~x367 & ~x392 & ~x393 & ~x588 & ~x626 & ~x642 & ~x643 & ~x670 & ~x671 & ~x683 & ~x702 & ~x716 & ~x718 & ~x721 & ~x727 & ~x729 & ~x734 & ~x736 & ~x737 & ~x738 & ~x739 & ~x742 & ~x743 & ~x744 & ~x746 & ~x747 & ~x748 & ~x751 & ~x752 & ~x754 & ~x755 & ~x756 & ~x757 & ~x758 & ~x759 & ~x761 & ~x763 & ~x765 & ~x766 & ~x768 & ~x769 & ~x770 & ~x771 & ~x772 & ~x774 & ~x775 & ~x778 & ~x779 & ~x781 & ~x782 & ~x783;
assign c5406 =  x686 & ~x4 & ~x7 & ~x10 & ~x11 & ~x33 & ~x84 & ~x89 & ~x115 & ~x142 & ~x145 & ~x168 & ~x170 & ~x255 & ~x256 & ~x257 & ~x258 & ~x282 & ~x287 & ~x288 & ~x309 & ~x315 & ~x338 & ~x342 & ~x343 & ~x344 & ~x364 & ~x369 & ~x371 & ~x395 & ~x396 & ~x398 & ~x400 & ~x422 & ~x424 & ~x425 & ~x426 & ~x447 & ~x450 & ~x451 & ~x452 & ~x506 & ~x534 & ~x559 & ~x644 & ~x671 & ~x759;
assign c5408 = ~x0 & ~x14 & ~x17 & ~x26 & ~x29 & ~x42 & ~x50 & ~x56 & ~x67 & ~x68 & ~x69 & ~x82 & ~x94 & ~x95 & ~x96 & ~x98 & ~x113 & ~x117 & ~x121 & ~x123 & ~x125 & ~x135 & ~x146 & ~x151 & ~x163 & ~x165 & ~x170 & ~x177 & ~x179 & ~x185 & ~x195 & ~x230 & ~x250 & ~x283 & ~x390 & ~x417 & ~x418 & ~x607 & ~x609 & ~x627 & ~x628 & ~x629 & ~x633 & ~x640 & ~x646 & ~x654 & ~x663 & ~x690 & ~x694 & ~x697 & ~x702 & ~x707 & ~x708 & ~x711 & ~x717 & ~x719 & ~x721 & ~x723 & ~x724 & ~x730 & ~x733 & ~x734 & ~x760 & ~x764 & ~x771;
assign c5410 =  x708 & ~x2 & ~x4 & ~x54 & ~x62 & ~x84 & ~x114 & ~x117 & ~x140 & ~x143 & ~x230 & ~x255 & ~x280 & ~x284 & ~x286 & ~x315 & ~x316 & ~x367 & ~x661 & ~x664 & ~x757;
assign c5412 =  x75 & ~x288 & ~x315 & ~x371 & ~x399 & ~x424 & ~x505;
assign c5414 =  x358 &  x425 & ~x4 & ~x10 & ~x21 & ~x27 & ~x29 & ~x41 & ~x43 & ~x46 & ~x48 & ~x50 & ~x60 & ~x77 & ~x79 & ~x82 & ~x92 & ~x94 & ~x97 & ~x131 & ~x132 & ~x146 & ~x159 & ~x163 & ~x185 & ~x186 & ~x200 & ~x204 & ~x223 & ~x225 & ~x257 & ~x319 & ~x391 & ~x560 & ~x586 & ~x613 & ~x638 & ~x639 & ~x650 & ~x652 & ~x654 & ~x663 & ~x671 & ~x715 & ~x722 & ~x726 & ~x733 & ~x737 & ~x742 & ~x756 & ~x771;
assign c5416 =  x426 &  x542 & ~x15 & ~x54 & ~x117 & ~x151 & ~x195 & ~x253 & ~x255 & ~x319 & ~x616 & ~x733 & ~x770;
assign c5418 =  x489 & ~x2 & ~x7 & ~x8 & ~x10 & ~x11 & ~x13 & ~x23 & ~x29 & ~x33 & ~x34 & ~x38 & ~x59 & ~x65 & ~x88 & ~x154 & ~x166 & ~x175 & ~x176 & ~x203 & ~x226 & ~x241 & ~x243 & ~x251 & ~x252 & ~x310 & ~x336 & ~x338 & ~x393 & ~x395 & ~x552 & ~x554 & ~x562 & ~x579 & ~x580 & ~x581 & ~x582 & ~x671 & ~x718 & ~x720 & ~x749 & ~x775 & ~x776;
assign c5420 =  x296 &  x484 & ~x4 & ~x215 & ~x348;
assign c5422 =  x440 & ~x3 & ~x11 & ~x17 & ~x21 & ~x27 & ~x32 & ~x35 & ~x41 & ~x43 & ~x50 & ~x55 & ~x56 & ~x59 & ~x60 & ~x61 & ~x67 & ~x68 & ~x85 & ~x86 & ~x99 & ~x114 & ~x120 & ~x141 & ~x142 & ~x145 & ~x150 & ~x170 & ~x172 & ~x175 & ~x200 & ~x201 & ~x226 & ~x230 & ~x254 & ~x255 & ~x257 & ~x280 & ~x282 & ~x379 & ~x475 & ~x560 & ~x587 & ~x588 & ~x615 & ~x616 & ~x718 & ~x729 & ~x742 & ~x744 & ~x746 & ~x749 & ~x758 & ~x761 & ~x767 & ~x768 & ~x769 & ~x771 & ~x775 & ~x777 & ~x780;
assign c5424 =  x613 & ~x49 & ~x126 & ~x139 & ~x339 & ~x340 & ~x507 & ~x643 & ~x714 & ~x745;
assign c5426 =  x529 &  x585 & ~x0 & ~x18 & ~x31 & ~x33 & ~x35 & ~x51 & ~x91 & ~x167 & ~x201 & ~x230 & ~x253 & ~x256 & ~x283 & ~x284 & ~x310 & ~x342 & ~x477 & ~x506 & ~x507 & ~x756 & ~x759;
assign c5428 =  x481 & ~x43 & ~x44 & ~x58 & ~x68 & ~x70 & ~x87 & ~x91 & ~x119 & ~x128 & ~x136 & ~x142 & ~x147 & ~x155 & ~x160 & ~x172 & ~x186 & ~x199 & ~x204 & ~x212 & ~x213 & ~x214 & ~x215 & ~x224 & ~x227 & ~x229 & ~x254 & ~x337 & ~x365 & ~x423 & ~x531 & ~x575 & ~x602 & ~x603 & ~x615 & ~x631 & ~x644 & ~x646 & ~x663 & ~x677 & ~x712 & ~x732 & ~x744 & ~x778 & ~x779;
assign c5430 =  x103 & ~x140 & ~x314 & ~x344 & ~x364 & ~x368 & ~x399 & ~x536 & ~x643;
assign c5432 = ~x0 & ~x2 & ~x3 & ~x5 & ~x9 & ~x10 & ~x11 & ~x13 & ~x14 & ~x15 & ~x16 & ~x18 & ~x20 & ~x21 & ~x23 & ~x25 & ~x26 & ~x28 & ~x31 & ~x32 & ~x35 & ~x36 & ~x37 & ~x38 & ~x39 & ~x40 & ~x41 & ~x42 & ~x43 & ~x44 & ~x45 & ~x46 & ~x47 & ~x49 & ~x50 & ~x54 & ~x55 & ~x56 & ~x58 & ~x62 & ~x63 & ~x70 & ~x71 & ~x73 & ~x74 & ~x83 & ~x91 & ~x94 & ~x95 & ~x97 & ~x100 & ~x114 & ~x116 & ~x117 & ~x118 & ~x120 & ~x122 & ~x125 & ~x140 & ~x143 & ~x146 & ~x147 & ~x150 & ~x169 & ~x170 & ~x171 & ~x174 & ~x176 & ~x177 & ~x179 & ~x196 & ~x197 & ~x200 & ~x203 & ~x204 & ~x205 & ~x226 & ~x227 & ~x228 & ~x231 & ~x254 & ~x257 & ~x280 & ~x281 & ~x282 & ~x283 & ~x284 & ~x285 & ~x309 & ~x337 & ~x340 & ~x367 & ~x381 & ~x392 & ~x395 & ~x448 & ~x560 & ~x616 & ~x672 & ~x727 & ~x728 & ~x729 & ~x730 & ~x732 & ~x741 & ~x744 & ~x747 & ~x757 & ~x758 & ~x762 & ~x765 & ~x767 & ~x770 & ~x771 & ~x774 & ~x775 & ~x781 & ~x783;
assign c5434 =  x439 & ~x2 & ~x15 & ~x22 & ~x23 & ~x32 & ~x38 & ~x50 & ~x52 & ~x55 & ~x68 & ~x70 & ~x74 & ~x84 & ~x86 & ~x91 & ~x92 & ~x97 & ~x98 & ~x112 & ~x120 & ~x124 & ~x151 & ~x171 & ~x173 & ~x175 & ~x179 & ~x180 & ~x182 & ~x197 & ~x202 & ~x206 & ~x230 & ~x238 & ~x252 & ~x255 & ~x257 & ~x259 & ~x268 & ~x269 & ~x282 & ~x309 & ~x336 & ~x447 & ~x560 & ~x615 & ~x644 & ~x671 & ~x704 & ~x705 & ~x763 & ~x771 & ~x781;
assign c5436 = ~x41 & ~x48 & ~x68 & ~x69 & ~x80 & ~x100 & ~x114 & ~x161 & ~x174 & ~x184 & ~x186 & ~x195 & ~x214 & ~x217 & ~x223 & ~x226 & ~x228 & ~x242 & ~x308 & ~x390 & ~x417 & ~x575 & ~x577 & ~x587 & ~x601 & ~x608 & ~x644 & ~x676 & ~x682 & ~x686 & ~x692 & ~x698 & ~x713 & ~x719 & ~x722 & ~x724 & ~x725 & ~x731 & ~x750 & ~x758 & ~x764 & ~x772 & ~x774;
assign c5438 =  x408 & ~x1 & ~x2 & ~x3 & ~x6 & ~x7 & ~x8 & ~x13 & ~x14 & ~x15 & ~x16 & ~x18 & ~x21 & ~x22 & ~x23 & ~x24 & ~x25 & ~x28 & ~x30 & ~x31 & ~x32 & ~x34 & ~x35 & ~x36 & ~x37 & ~x38 & ~x40 & ~x42 & ~x43 & ~x44 & ~x46 & ~x47 & ~x48 & ~x51 & ~x54 & ~x55 & ~x56 & ~x58 & ~x59 & ~x60 & ~x63 & ~x65 & ~x66 & ~x67 & ~x68 & ~x69 & ~x70 & ~x71 & ~x72 & ~x73 & ~x76 & ~x77 & ~x80 & ~x82 & ~x84 & ~x87 & ~x88 & ~x89 & ~x91 & ~x92 & ~x94 & ~x96 & ~x97 & ~x98 & ~x99 & ~x100 & ~x101 & ~x102 & ~x106 & ~x108 & ~x110 & ~x111 & ~x114 & ~x115 & ~x116 & ~x121 & ~x123 & ~x124 & ~x125 & ~x126 & ~x127 & ~x130 & ~x131 & ~x132 & ~x135 & ~x136 & ~x138 & ~x139 & ~x140 & ~x143 & ~x145 & ~x146 & ~x148 & ~x149 & ~x150 & ~x151 & ~x153 & ~x155 & ~x156 & ~x157 & ~x158 & ~x160 & ~x165 & ~x166 & ~x168 & ~x170 & ~x173 & ~x176 & ~x178 & ~x179 & ~x180 & ~x182 & ~x185 & ~x186 & ~x187 & ~x189 & ~x190 & ~x191 & ~x199 & ~x200 & ~x205 & ~x206 & ~x211 & ~x213 & ~x214 & ~x215 & ~x218 & ~x224 & ~x225 & ~x226 & ~x227 & ~x228 & ~x229 & ~x231 & ~x232 & ~x233 & ~x234 & ~x235 & ~x238 & ~x239 & ~x240 & ~x241 & ~x250 & ~x251 & ~x255 & ~x256 & ~x257 & ~x259 & ~x261 & ~x263 & ~x269 & ~x270 & ~x279 & ~x281 & ~x282 & ~x285 & ~x286 & ~x287 & ~x288 & ~x307 & ~x308 & ~x309 & ~x311 & ~x312 & ~x334 & ~x336 & ~x337 & ~x340 & ~x560 & ~x564 & ~x565 & ~x575 & ~x576 & ~x577 & ~x587 & ~x588 & ~x589 & ~x590 & ~x591 & ~x592 & ~x593 & ~x594 & ~x595 & ~x596 & ~x600 & ~x601 & ~x606 & ~x609 & ~x612 & ~x613 & ~x615 & ~x617 & ~x618 & ~x623 & ~x625 & ~x627 & ~x628 & ~x629 & ~x633 & ~x634 & ~x635 & ~x638 & ~x639 & ~x641 & ~x643 & ~x645 & ~x646 & ~x649 & ~x652 & ~x653 & ~x656 & ~x657 & ~x658 & ~x659 & ~x662 & ~x664 & ~x665 & ~x666 & ~x671 & ~x673 & ~x674 & ~x676 & ~x677 & ~x679 & ~x680 & ~x681 & ~x682 & ~x683 & ~x686 & ~x687 & ~x688 & ~x689 & ~x690 & ~x695 & ~x697 & ~x699 & ~x700 & ~x701 & ~x702 & ~x703 & ~x706 & ~x708 & ~x710 & ~x711 & ~x712 & ~x716 & ~x717 & ~x719 & ~x720 & ~x723 & ~x724 & ~x727 & ~x728 & ~x730 & ~x731 & ~x732 & ~x735 & ~x736 & ~x739 & ~x741 & ~x742 & ~x743 & ~x744 & ~x746 & ~x747 & ~x748 & ~x749 & ~x750 & ~x751 & ~x754 & ~x755 & ~x756 & ~x758 & ~x760 & ~x765 & ~x767 & ~x769 & ~x774 & ~x776 & ~x777 & ~x778 & ~x782 & ~x783;
assign c5440 =  x317;
assign c5442 = ~x9 & ~x11 & ~x27 & ~x28 & ~x38 & ~x41 & ~x57 & ~x66 & ~x68 & ~x92 & ~x97 & ~x114 & ~x115 & ~x122 & ~x145 & ~x148 & ~x152 & ~x169 & ~x171 & ~x177 & ~x204 & ~x206 & ~x253 & ~x268 & ~x277 & ~x335 & ~x418 & ~x419 & ~x447 & ~x503 & ~x504 & ~x692 & ~x773;
assign c5444 =  x302 & ~x0 & ~x2 & ~x12 & ~x15 & ~x19 & ~x27 & ~x32 & ~x33 & ~x88 & ~x145 & ~x166 & ~x201 & ~x224 & ~x225 & ~x255 & ~x257 & ~x310 & ~x364 & ~x379 & ~x672 & ~x700 & ~x771 & ~x783;
assign c5446 = ~x0 & ~x2 & ~x3 & ~x6 & ~x11 & ~x25 & ~x26 & ~x62 & ~x114 & ~x166 & ~x172 & ~x232 & ~x234 & ~x256 & ~x258 & ~x259 & ~x261 & ~x309 & ~x316 & ~x337 & ~x341 & ~x373 & ~x375 & ~x394 & ~x395 & ~x401 & ~x454 & ~x474 & ~x506 & ~x531 & ~x642 & ~x671 & ~x700 & ~x756 & ~x759 & ~x783;
assign c5448 =  x732 & ~x7 & ~x340 & ~x368 & ~x533 & ~x534;
assign c5450 =  x400 &  x537 &  x547 & ~x76 & ~x719 & ~x744;
assign c5452 =  x511 & ~x0 & ~x1 & ~x5 & ~x7 & ~x8 & ~x12 & ~x14 & ~x26 & ~x28 & ~x29 & ~x32 & ~x33 & ~x38 & ~x41 & ~x46 & ~x48 & ~x51 & ~x54 & ~x55 & ~x58 & ~x60 & ~x67 & ~x74 & ~x75 & ~x82 & ~x83 & ~x84 & ~x91 & ~x97 & ~x104 & ~x105 & ~x106 & ~x115 & ~x116 & ~x117 & ~x121 & ~x122 & ~x141 & ~x144 & ~x147 & ~x148 & ~x154 & ~x195 & ~x198 & ~x200 & ~x201 & ~x202 & ~x204 & ~x223 & ~x224 & ~x226 & ~x229 & ~x235 & ~x256 & ~x259 & ~x260 & ~x282 & ~x287 & ~x288 & ~x289 & ~x290 & ~x308 & ~x309 & ~x312 & ~x340 & ~x341 & ~x366 & ~x479 & ~x559 & ~x588 & ~x644 & ~x671 & ~x672 & ~x674 & ~x678 & ~x703 & ~x705 & ~x710 & ~x714 & ~x715 & ~x716 & ~x719 & ~x723 & ~x724 & ~x727 & ~x730 & ~x733 & ~x737 & ~x741 & ~x747 & ~x751 & ~x752 & ~x753 & ~x754 & ~x758 & ~x761 & ~x763 & ~x764 & ~x765 & ~x767 & ~x768 & ~x773 & ~x774 & ~x776 & ~x779 & ~x780 & ~x782;
assign c5454 =  x299 &  x301 & ~x57 & ~x59 & ~x97 & ~x123 & ~x198 & ~x201 & ~x227 & ~x308 & ~x385;
assign c5456 = ~x2 & ~x7 & ~x12 & ~x16 & ~x26 & ~x42 & ~x46 & ~x50 & ~x53 & ~x54 & ~x60 & ~x70 & ~x75 & ~x81 & ~x90 & ~x95 & ~x98 & ~x100 & ~x114 & ~x120 & ~x124 & ~x125 & ~x132 & ~x142 & ~x148 & ~x163 & ~x167 & ~x225 & ~x228 & ~x250 & ~x273 & ~x281 & ~x306 & ~x336 & ~x337 & ~x419 & ~x445 & ~x446 & ~x628 & ~x659 & ~x663 & ~x671 & ~x681 & ~x684 & ~x690 & ~x699 & ~x715 & ~x716 & ~x717 & ~x718 & ~x723 & ~x725 & ~x726 & ~x728 & ~x729 & ~x730 & ~x734 & ~x742 & ~x745 & ~x748 & ~x760 & ~x766 & ~x768 & ~x777;
assign c5458 =  x301 &  x482 &  x484 &  x510 & ~x1 & ~x10 & ~x17 & ~x19 & ~x20 & ~x22 & ~x24 & ~x26 & ~x31 & ~x32 & ~x33 & ~x38 & ~x39 & ~x41 & ~x42 & ~x44 & ~x52 & ~x71 & ~x74 & ~x75 & ~x85 & ~x88 & ~x96 & ~x112 & ~x117 & ~x125 & ~x144 & ~x149 & ~x151 & ~x152 & ~x167 & ~x171 & ~x172 & ~x173 & ~x174 & ~x180 & ~x200 & ~x201 & ~x202 & ~x204 & ~x229 & ~x252 & ~x253 & ~x254 & ~x308 & ~x309 & ~x310 & ~x364 & ~x559 & ~x587 & ~x616 & ~x671 & ~x734 & ~x739 & ~x741 & ~x742 & ~x747 & ~x754 & ~x758 & ~x768 & ~x770 & ~x771 & ~x773 & ~x774 & ~x775 & ~x778 & ~x779 & ~x781 & ~x782;
assign c5460 = ~x0 & ~x1 & ~x3 & ~x4 & ~x6 & ~x10 & ~x11 & ~x13 & ~x15 & ~x24 & ~x28 & ~x29 & ~x30 & ~x31 & ~x32 & ~x37 & ~x38 & ~x54 & ~x59 & ~x62 & ~x64 & ~x66 & ~x83 & ~x89 & ~x92 & ~x116 & ~x119 & ~x120 & ~x139 & ~x141 & ~x142 & ~x143 & ~x146 & ~x147 & ~x149 & ~x151 & ~x167 & ~x171 & ~x173 & ~x174 & ~x177 & ~x178 & ~x195 & ~x196 & ~x197 & ~x198 & ~x202 & ~x203 & ~x206 & ~x228 & ~x233 & ~x252 & ~x255 & ~x257 & ~x259 & ~x260 & ~x281 & ~x282 & ~x288 & ~x289 & ~x290 & ~x312 & ~x336 & ~x339 & ~x341 & ~x342 & ~x343 & ~x344 & ~x365 & ~x367 & ~x369 & ~x370 & ~x394 & ~x395 & ~x421 & ~x423 & ~x424 & ~x433 & ~x448 & ~x451 & ~x461 & ~x476 & ~x478 & ~x504 & ~x505 & ~x700 & ~x728 & ~x756;
assign c5462 =  x237 & ~x1 & ~x32 & ~x54 & ~x80 & ~x91 & ~x108 & ~x144 & ~x175 & ~x176;
assign c5464 =  x134 & ~x58 & ~x168 & ~x196 & ~x201 & ~x228 & ~x367 & ~x449 & ~x476 & ~x698;
assign c5466 = ~x4 & ~x23 & ~x39 & ~x40 & ~x43 & ~x65 & ~x69 & ~x70 & ~x97 & ~x150 & ~x151 & ~x153 & ~x173 & ~x178 & ~x180 & ~x203 & ~x232 & ~x361 & ~x362 & ~x555 & ~x560 & ~x567 & ~x568 & ~x569 & ~x572 & ~x574 & ~x580 & ~x581 & ~x583 & ~x584 & ~x694 & ~x697 & ~x720 & ~x743;
assign c5468 = ~x9 & ~x13 & ~x20 & ~x30 & ~x41 & ~x66 & ~x69 & ~x71 & ~x82 & ~x97 & ~x104 & ~x143 & ~x171 & ~x173 & ~x179 & ~x232 & ~x233 & ~x242 & ~x362 & ~x363 & ~x388 & ~x389 & ~x390 & ~x607 & ~x615 & ~x619 & ~x624 & ~x669 & ~x686 & ~x688 & ~x695 & ~x716 & ~x719 & ~x726 & ~x733 & ~x734 & ~x747 & ~x752 & ~x770 & ~x778 & ~x780;
assign c5470 = ~x6 & ~x11 & ~x13 & ~x22 & ~x25 & ~x26 & ~x39 & ~x40 & ~x43 & ~x46 & ~x59 & ~x60 & ~x67 & ~x68 & ~x87 & ~x94 & ~x95 & ~x96 & ~x97 & ~x114 & ~x117 & ~x118 & ~x120 & ~x143 & ~x145 & ~x167 & ~x171 & ~x173 & ~x174 & ~x176 & ~x180 & ~x181 & ~x196 & ~x202 & ~x203 & ~x207 & ~x226 & ~x230 & ~x232 & ~x235 & ~x236 & ~x238 & ~x259 & ~x266 & ~x336 & ~x361 & ~x362 & ~x388 & ~x390 & ~x391 & ~x504 & ~x560 & ~x587 & ~x655 & ~x656 & ~x671 & ~x684 & ~x689 & ~x693 & ~x702 & ~x704 & ~x755 & ~x783;
assign c5472 =  x411 &  x493 &  x497 &  x512 &  x528 & ~x6 & ~x60 & ~x92 & ~x142 & ~x185 & ~x648 & ~x651 & ~x762;
assign c5474 =  x211 & ~x11 & ~x26 & ~x57 & ~x90 & ~x118 & ~x138 & ~x148 & ~x149 & ~x216 & ~x226 & ~x233 & ~x309 & ~x587 & ~x717;
assign c5476 = ~x24 & ~x27 & ~x28 & ~x29 & ~x34 & ~x35 & ~x38 & ~x54 & ~x57 & ~x60 & ~x62 & ~x90 & ~x112 & ~x114 & ~x118 & ~x119 & ~x141 & ~x167 & ~x169 & ~x174 & ~x196 & ~x198 & ~x203 & ~x205 & ~x256 & ~x257 & ~x280 & ~x283 & ~x284 & ~x287 & ~x289 & ~x309 & ~x334 & ~x336 & ~x339 & ~x361 & ~x363 & ~x386 & ~x387 & ~x388 & ~x607 & ~x635 & ~x663 & ~x690 & ~x717 & ~x718 & ~x743 & ~x746 & ~x759 & ~x774;
assign c5478 = ~x1 & ~x3 & ~x4 & ~x5 & ~x6 & ~x8 & ~x11 & ~x14 & ~x32 & ~x33 & ~x35 & ~x36 & ~x37 & ~x38 & ~x55 & ~x56 & ~x61 & ~x62 & ~x63 & ~x65 & ~x85 & ~x90 & ~x91 & ~x93 & ~x110 & ~x111 & ~x112 & ~x115 & ~x118 & ~x121 & ~x139 & ~x141 & ~x145 & ~x146 & ~x150 & ~x169 & ~x172 & ~x173 & ~x174 & ~x176 & ~x195 & ~x198 & ~x199 & ~x202 & ~x203 & ~x231 & ~x252 & ~x254 & ~x257 & ~x259 & ~x261 & ~x284 & ~x309 & ~x310 & ~x334 & ~x364 & ~x365 & ~x449 & ~x476 & ~x477 & ~x479 & ~x504 & ~x505 & ~x506 & ~x606 & ~x607 & ~x633 & ~x635 & ~x688 & ~x716 & ~x719 & ~x728 & ~x743 & ~x772 & ~x781 & ~x782 & ~x783;
assign c5480 =  x483 &  x597 & ~x10 & ~x15 & ~x34 & ~x57 & ~x58 & ~x110 & ~x112 & ~x116 & ~x146 & ~x150 & ~x175 & ~x232 & ~x256 & ~x282 & ~x315 & ~x393 & ~x699 & ~x700 & ~x768;
assign c5482 =  x412 &  x481 &  x483 &  x490 &  x493 &  x499 & ~x7 & ~x10 & ~x11 & ~x14 & ~x22 & ~x33 & ~x45 & ~x48 & ~x51 & ~x55 & ~x64 & ~x66 & ~x71 & ~x81 & ~x82 & ~x88 & ~x90 & ~x91 & ~x92 & ~x93 & ~x98 & ~x104 & ~x105 & ~x115 & ~x120 & ~x125 & ~x138 & ~x140 & ~x148 & ~x149 & ~x161 & ~x163 & ~x165 & ~x171 & ~x179 & ~x180 & ~x183 & ~x195 & ~x199 & ~x204 & ~x205 & ~x206 & ~x212 & ~x224 & ~x228 & ~x242 & ~x243 & ~x258 & ~x259 & ~x288 & ~x339 & ~x363 & ~x559 & ~x560 & ~x575 & ~x578 & ~x589 & ~x591 & ~x592 & ~x595 & ~x600 & ~x614 & ~x627 & ~x631 & ~x642 & ~x646 & ~x650 & ~x654 & ~x656 & ~x659 & ~x662 & ~x664 & ~x667 & ~x671 & ~x688 & ~x693 & ~x707 & ~x712 & ~x716 & ~x726 & ~x749 & ~x751 & ~x753 & ~x756 & ~x758 & ~x783;
assign c5484 =  x273 &  x494 &  x522 &  x540 & ~x42 & ~x70 & ~x114 & ~x201 & ~x215 & ~x582 & ~x584 & ~x585 & ~x699 & ~x706;
assign c5486 =  x358 & ~x3 & ~x4 & ~x9 & ~x11 & ~x12 & ~x15 & ~x22 & ~x25 & ~x26 & ~x27 & ~x28 & ~x29 & ~x30 & ~x31 & ~x32 & ~x33 & ~x35 & ~x38 & ~x40 & ~x51 & ~x58 & ~x59 & ~x62 & ~x65 & ~x66 & ~x84 & ~x85 & ~x86 & ~x88 & ~x89 & ~x90 & ~x93 & ~x112 & ~x114 & ~x115 & ~x117 & ~x118 & ~x141 & ~x142 & ~x143 & ~x144 & ~x145 & ~x169 & ~x170 & ~x172 & ~x173 & ~x174 & ~x175 & ~x176 & ~x196 & ~x197 & ~x202 & ~x204 & ~x227 & ~x228 & ~x229 & ~x230 & ~x233 & ~x234 & ~x252 & ~x254 & ~x255 & ~x256 & ~x257 & ~x258 & ~x260 & ~x261 & ~x282 & ~x283 & ~x287 & ~x312 & ~x322 & ~x336 & ~x338 & ~x340 & ~x364 & ~x365 & ~x366 & ~x392 & ~x393 & ~x395 & ~x504 & ~x534 & ~x535 & ~x544 & ~x588 & ~x728 & ~x757;
assign c5488 =  x509 & ~x8 & ~x10 & ~x11 & ~x12 & ~x32 & ~x34 & ~x85 & ~x86 & ~x88 & ~x89 & ~x91 & ~x95 & ~x96 & ~x97 & ~x171 & ~x173 & ~x174 & ~x193 & ~x195 & ~x198 & ~x223 & ~x252 & ~x259 & ~x281 & ~x282 & ~x283 & ~x309 & ~x310 & ~x312 & ~x314 & ~x391 & ~x395 & ~x476 & ~x732 & ~x761 & ~x772 & ~x777;
assign c5490 =  x328 &  x355 & ~x12 & ~x28 & ~x43 & ~x64 & ~x174 & ~x206 & ~x232 & ~x233 & ~x257 & ~x281 & ~x365 & ~x407 & ~x672 & ~x759;
assign c5492 =  x397 & ~x8 & ~x16 & ~x24 & ~x29 & ~x43 & ~x62 & ~x72 & ~x73 & ~x82 & ~x83 & ~x89 & ~x97 & ~x100 & ~x102 & ~x137 & ~x179 & ~x205 & ~x206 & ~x223 & ~x235 & ~x241 & ~x257 & ~x335 & ~x336 & ~x363 & ~x420 & ~x587 & ~x614 & ~x615 & ~x646 & ~x661 & ~x692 & ~x714 & ~x735 & ~x754 & ~x756 & ~x759 & ~x769 & ~x770;
assign c5494 =  x105 & ~x2 & ~x3 & ~x9 & ~x55 & ~x56 & ~x63 & ~x82 & ~x89 & ~x90 & ~x110 & ~x111 & ~x114 & ~x116 & ~x146 & ~x169 & ~x170 & ~x171 & ~x172 & ~x195 & ~x196 & ~x198 & ~x201 & ~x202 & ~x203 & ~x229 & ~x256 & ~x284 & ~x311 & ~x314 & ~x337 & ~x341 & ~x342 & ~x343 & ~x366 & ~x368 & ~x370 & ~x419 & ~x420 & ~x448 & ~x615 & ~x616 & ~x643 & ~x671;
assign c5496 =  x584 & ~x4 & ~x6 & ~x19 & ~x23 & ~x30 & ~x38 & ~x39 & ~x63 & ~x91 & ~x92 & ~x110 & ~x112 & ~x115 & ~x140 & ~x168 & ~x200 & ~x224 & ~x227 & ~x229 & ~x233 & ~x253 & ~x260 & ~x308 & ~x476 & ~x478 & ~x590 & ~x745 & ~x748 & ~x756 & ~x776;
assign c5498 =  x397 &  x466 &  x480 &  x481 &  x489 &  x517 & ~x44 & ~x74 & ~x76 & ~x87 & ~x101 & ~x104 & ~x128 & ~x140 & ~x149 & ~x173 & ~x197 & ~x198 & ~x205 & ~x228 & ~x254 & ~x259 & ~x284 & ~x309 & ~x312 & ~x364 & ~x588 & ~x609 & ~x644 & ~x649 & ~x664 & ~x677 & ~x678 & ~x691 & ~x693 & ~x699 & ~x707 & ~x715 & ~x741 & ~x753 & ~x766;
assign c51 =  x206;
assign c53 =  x336;
assign c55 =  x351 &  x361 &  x378 &  x386 &  x387 &  x403 &  x404 &  x408 &  x414 &  x446 &  x471 &  x472 &  x474 & ~x0 & ~x4 & ~x25 & ~x29 & ~x44 & ~x57 & ~x68 & ~x74 & ~x84 & ~x90 & ~x94 & ~x98 & ~x105 & ~x106 & ~x113 & ~x118 & ~x131 & ~x156 & ~x164 & ~x171 & ~x181 & ~x195 & ~x206 & ~x208 & ~x223 & ~x261 & ~x282 & ~x312 & ~x588 & ~x651 & ~x652 & ~x671 & ~x678 & ~x679 & ~x685 & ~x692 & ~x703 & ~x712 & ~x715 & ~x719 & ~x722 & ~x724 & ~x735 & ~x737 & ~x742 & ~x747 & ~x748 & ~x768 & ~x773 & ~x775 & ~x776;
assign c57 = ~x130 & ~x246 & ~x275 & ~x330 & ~x451 & ~x529 & ~x726;
assign c59 =  x32;
assign c511 =  x258;
assign c513 =  x10;
assign c515 =  x380 &  x385 &  x387 &  x409 &  x417 &  x445 &  x471 & ~x2 & ~x3 & ~x24 & ~x34 & ~x35 & ~x37 & ~x50 & ~x60 & ~x61 & ~x63 & ~x81 & ~x82 & ~x96 & ~x103 & ~x110 & ~x111 & ~x113 & ~x115 & ~x125 & ~x132 & ~x133 & ~x136 & ~x141 & ~x144 & ~x162 & ~x173 & ~x192 & ~x228 & ~x260 & ~x280 & ~x311 & ~x313 & ~x314 & ~x338 & ~x342 & ~x363 & ~x364 & ~x365 & ~x367 & ~x369 & ~x393 & ~x588 & ~x591 & ~x617 & ~x621 & ~x624 & ~x626 & ~x642 & ~x648 & ~x659 & ~x660 & ~x673 & ~x679 & ~x686 & ~x696 & ~x699 & ~x700 & ~x713 & ~x722 & ~x736 & ~x751 & ~x753 & ~x760 & ~x763 & ~x773 & ~x774;
assign c517 = ~x300 & ~x385 & ~x440 & ~x557;
assign c519 =  x14;
assign c521 =  x310;
assign c523 =  x282;
assign c525 =  x372 &  x380 &  x417 &  x418 &  x424 & ~x6 & ~x31 & ~x45 & ~x70 & ~x82 & ~x92 & ~x103 & ~x108 & ~x111 & ~x112 & ~x133 & ~x139 & ~x146 & ~x182 & ~x193 & ~x196 & ~x210 & ~x211 & ~x217 & ~x219 & ~x222 & ~x245 & ~x273 & ~x336 & ~x337 & ~x341 & ~x562 & ~x594 & ~x604 & ~x613 & ~x640 & ~x650 & ~x688 & ~x691 & ~x706 & ~x709 & ~x710 & ~x721 & ~x725 & ~x728 & ~x756 & ~x777 & ~x778;
assign c527 = ~x276 & ~x361 & ~x389 & ~x397 & ~x417 & ~x474 & ~x529 & ~x645;
assign c529 =  x386 &  x410 &  x416 &  x417 &  x444 &  x445 &  x464 & ~x6 & ~x7 & ~x9 & ~x19 & ~x21 & ~x24 & ~x27 & ~x36 & ~x39 & ~x56 & ~x61 & ~x75 & ~x80 & ~x82 & ~x83 & ~x91 & ~x93 & ~x97 & ~x104 & ~x107 & ~x108 & ~x115 & ~x116 & ~x120 & ~x121 & ~x122 & ~x134 & ~x141 & ~x143 & ~x146 & ~x165 & ~x171 & ~x176 & ~x182 & ~x188 & ~x192 & ~x194 & ~x198 & ~x207 & ~x210 & ~x223 & ~x224 & ~x225 & ~x235 & ~x236 & ~x253 & ~x256 & ~x260 & ~x262 & ~x287 & ~x310 & ~x313 & ~x338 & ~x340 & ~x366 & ~x532 & ~x594 & ~x620 & ~x626 & ~x627 & ~x634 & ~x637 & ~x639 & ~x640 & ~x642 & ~x658 & ~x674 & ~x681 & ~x699 & ~x702 & ~x707 & ~x708 & ~x710 & ~x729 & ~x731 & ~x745 & ~x747 & ~x749 & ~x750 & ~x755 & ~x757 & ~x768 & ~x769 & ~x776;
assign c531 =  x345 &  x372 &  x373 &  x374 &  x423 &  x424 & ~x246 & ~x592;
assign c533 =  x272 &  x301 &  x302 &  x328 &  x351 &  x358 &  x386 &  x468 &  x520 &  x528 & ~x363 & ~x371;
assign c535 =  x661 & ~x362;
assign c537 = ~x3 & ~x6 & ~x9 & ~x11 & ~x15 & ~x27 & ~x47 & ~x55 & ~x56 & ~x64 & ~x76 & ~x77 & ~x78 & ~x87 & ~x90 & ~x94 & ~x100 & ~x107 & ~x112 & ~x114 & ~x127 & ~x130 & ~x136 & ~x137 & ~x140 & ~x141 & ~x143 & ~x148 & ~x152 & ~x153 & ~x171 & ~x180 & ~x181 & ~x195 & ~x198 & ~x203 & ~x208 & ~x222 & ~x238 & ~x251 & ~x254 & ~x290 & ~x291 & ~x310 & ~x316 & ~x318 & ~x335 & ~x341 & ~x365 & ~x370 & ~x396 & ~x399 & ~x425 & ~x426 & ~x428 & ~x448 & ~x588 & ~x617 & ~x618 & ~x620 & ~x644 & ~x647 & ~x653 & ~x654 & ~x655 & ~x658 & ~x663 & ~x668 & ~x674 & ~x677 & ~x681 & ~x683 & ~x685 & ~x686 & ~x688 & ~x696 & ~x699 & ~x700 & ~x713 & ~x723 & ~x725 & ~x730 & ~x736 & ~x740 & ~x745 & ~x751 & ~x757 & ~x770 & ~x771 & ~x773 & ~x783;
assign c539 =  x232;
assign c541 =  x145;
assign c543 =  x42;
assign c545 =  x305 &  x416 &  x427 & ~x231 & ~x236 & ~x300 & ~x562 & ~x563 & ~x585;
assign c547 =  x301 &  x358 &  x379 &  x384 &  x386 &  x415 &  x467 &  x517 &  x520 &  x528 & ~x8 & ~x178 & ~x234 & ~x318;
assign c549 =  x15;
assign c551 =  x269 &  x324 &  x330 &  x351 &  x386 &  x529 & ~x643 & ~x671 & ~x677;
assign c553 =  x91;
assign c555 =  x378 &  x405 &  x407 &  x411 &  x417 &  x434 &  x437 &  x445 & ~x13 & ~x17 & ~x64 & ~x88 & ~x104 & ~x107 & ~x154 & ~x164 & ~x166 & ~x175 & ~x342 & ~x369 & ~x420 & ~x592 & ~x625 & ~x630 & ~x631 & ~x637 & ~x648 & ~x697 & ~x711 & ~x734 & ~x757;
assign c557 =  x325 &  x351 &  x356 &  x357 &  x358 &  x360 &  x382 &  x416 &  x445 &  x467 &  x489 &  x496 &  x557 & ~x34 & ~x66 & ~x149 & ~x232 & ~x261;
assign c559 =  x229;
assign c561 = ~x48 & ~x136 & ~x197 & ~x217 & ~x248 & ~x274 & ~x275 & ~x302 & ~x342 & ~x368 & ~x453 & ~x557 & ~x558 & ~x613 & ~x640 & ~x752;
assign c563 =  x353 &  x375 &  x380 &  x381 &  x445 &  x469 & ~x43 & ~x52 & ~x78 & ~x105 & ~x369 & ~x393 & ~x628 & ~x670 & ~x721 & ~x724 & ~x743;
assign c565 =  x33;
assign c567 =  x319 &  x375 &  x401 &  x402 & ~x8 & ~x27 & ~x77 & ~x114 & ~x131 & ~x136 & ~x159 & ~x160 & ~x162 & ~x186 & ~x217 & ~x226 & ~x246 & ~x247 & ~x272 & ~x273 & ~x274 & ~x301 & ~x503 & ~x588 & ~x727 & ~x729 & ~x779;
assign c569 =  x296 &  x324 &  x352 &  x358 &  x378 &  x385 &  x386 &  x407 &  x408 &  x409 &  x434 &  x439 &  x441 &  x444 &  x467 &  x556 &  x573 &  x574 &  x576;
assign c571 =  x743;
assign c573 =  x147;
assign c575 =  x117;
assign c577 =  x32;
assign c579 =  x297 & ~x9 & ~x15 & ~x25 & ~x34 & ~x40 & ~x59 & ~x61 & ~x68 & ~x76 & ~x77 & ~x79 & ~x82 & ~x91 & ~x92 & ~x101 & ~x103 & ~x109 & ~x112 & ~x114 & ~x129 & ~x151 & ~x154 & ~x164 & ~x168 & ~x170 & ~x174 & ~x180 & ~x182 & ~x199 & ~x205 & ~x206 & ~x218 & ~x222 & ~x224 & ~x233 & ~x236 & ~x245 & ~x247 & ~x252 & ~x255 & ~x272 & ~x301 & ~x308 & ~x309 & ~x316 & ~x335 & ~x366 & ~x368 & ~x369 & ~x393 & ~x598 & ~x614 & ~x620 & ~x622 & ~x630 & ~x634 & ~x644 & ~x653 & ~x657 & ~x659 & ~x667 & ~x672 & ~x674 & ~x677 & ~x686 & ~x708 & ~x728 & ~x729 & ~x737 & ~x739 & ~x748 & ~x751 & ~x757 & ~x766;
assign c581 =  x322 &  x347 &  x354 &  x411 &  x415 &  x431 & ~x4 & ~x14 & ~x16 & ~x35 & ~x47 & ~x72 & ~x73 & ~x80 & ~x81 & ~x94 & ~x121 & ~x126 & ~x135 & ~x168 & ~x170 & ~x179 & ~x206 & ~x225 & ~x229 & ~x258 & ~x310 & ~x336 & ~x338 & ~x535 & ~x569 & ~x640 & ~x644 & ~x645 & ~x670 & ~x674 & ~x698 & ~x732 & ~x749 & ~x776;
assign c583 =  x426 &  x451 &  x453 &  x454 &  x455 &  x456 &  x485 & ~x6 & ~x33 & ~x60 & ~x93 & ~x111 & ~x118 & ~x131 & ~x160 & ~x165 & ~x221 & ~x225 & ~x237 & ~x248 & ~x261 & ~x282 & ~x335 & ~x715 & ~x757 & ~x777;
assign c585 =  x268 &  x319 &  x423 & ~x51 & ~x93 & ~x107 & ~x211 & ~x246 & ~x765;
assign c587 =  x297 &  x300 &  x330 &  x356 &  x358 &  x386 &  x467 &  x496 &  x500 &  x522 &  x527 & ~x56 & ~x60 & ~x112 & ~x261 & ~x370 & ~x371 & ~x421 & ~x760;
assign c589 = ~x33 & ~x108 & ~x136 & ~x246 & ~x278 & ~x328 & ~x426;
assign c591 =  x360 &  x408 &  x435 &  x465 &  x470 &  x551 & ~x0 & ~x4 & ~x5 & ~x18 & ~x27 & ~x31 & ~x42 & ~x57 & ~x58 & ~x80 & ~x103 & ~x104 & ~x105 & ~x108 & ~x110 & ~x126 & ~x152 & ~x160 & ~x164 & ~x165 & ~x170 & ~x177 & ~x205 & ~x226 & ~x233 & ~x255 & ~x262 & ~x308 & ~x311 & ~x315 & ~x335 & ~x660 & ~x671 & ~x687 & ~x696 & ~x752 & ~x768 & ~x773 & ~x779;
assign c593 =  x61;
assign c595 =  x309;
assign c597 =  x347 &  x375 &  x429 &  x488 &  x515 & ~x133 & ~x162 & ~x218 & ~x334;
assign c599 =  x757;
assign c5101 =  x373 &  x401 & ~x136 & ~x161 & ~x217 & ~x245 & ~x272 & ~x332 & ~x781;
assign c5103 =  x388 &  x445 & ~x13 & ~x23 & ~x27 & ~x42 & ~x58 & ~x86 & ~x103 & ~x104 & ~x110 & ~x123 & ~x144 & ~x147 & ~x161 & ~x185 & ~x192 & ~x193 & ~x195 & ~x205 & ~x212 & ~x234 & ~x239 & ~x247 & ~x264 & ~x265 & ~x273 & ~x274 & ~x289 & ~x301 & ~x336 & ~x338 & ~x560 & ~x598 & ~x621 & ~x622 & ~x667 & ~x670 & ~x675 & ~x720 & ~x748 & ~x779;
assign c5105 =  x303 &  x326 &  x351 &  x355 &  x360 &  x380 &  x382 &  x383 &  x384 &  x385 &  x410 &  x488 &  x493 & ~x3 & ~x6 & ~x20 & ~x24 & ~x26 & ~x27 & ~x54 & ~x59 & ~x62 & ~x65 & ~x114 & ~x150 & ~x167 & ~x174 & ~x199 & ~x201 & ~x205 & ~x233 & ~x257 & ~x280 & ~x286 & ~x315 & ~x336 & ~x369 & ~x370 & ~x395 & ~x398 & ~x420 & ~x448 & ~x717 & ~x728 & ~x730 & ~x731 & ~x759 & ~x760 & ~x761 & ~x763 & ~x774;
assign c5107 =  x281;
assign c5109 =  x35;
assign c5111 =  x783;
assign c5113 = ~x106 & ~x134 & ~x243 & ~x271 & ~x278 & ~x397 & ~x452 & ~x454 & ~x533;
assign c5115 =  x114;
assign c5117 =  x296 &  x351 &  x377 &  x389 &  x417 &  x441 & ~x27 & ~x29 & ~x53 & ~x64 & ~x95 & ~x105 & ~x106 & ~x129 & ~x146 & ~x148 & ~x154 & ~x165 & ~x192 & ~x193 & ~x217 & ~x235 & ~x258 & ~x263 & ~x367 & ~x392 & ~x593 & ~x598 & ~x600 & ~x603 & ~x606 & ~x618 & ~x640 & ~x649 & ~x653 & ~x677 & ~x680 & ~x696 & ~x710 & ~x723 & ~x749 & ~x757 & ~x763 & ~x768 & ~x770 & ~x774 & ~x780;
assign c5119 =  x202;
assign c5121 =  x89;
assign c5123 =  x174;
assign c5125 =  x353 &  x418 &  x473 & ~x47 & ~x68 & ~x143 & ~x199 & ~x217 & ~x220 & ~x304 & ~x563 & ~x721 & ~x751;
assign c5127 =  x35;
assign c5129 =  x203;
assign c5131 = ~x26 & ~x48 & ~x74 & ~x102 & ~x159 & ~x167 & ~x248 & ~x255 & ~x307 & ~x453 & ~x592 & ~x612 & ~x617 & ~x619 & ~x641 & ~x669 & ~x679 & ~x701 & ~x757 & ~x780;
assign c5133 =  x310;
assign c5135 =  x33;
assign c5137 =  x543 &  x635 & ~x306;
assign c5139 =  x85;
assign c5141 =  x633 & ~x362;
assign c5143 =  x418 & ~x2 & ~x11 & ~x29 & ~x34 & ~x38 & ~x40 & ~x41 & ~x56 & ~x59 & ~x61 & ~x65 & ~x70 & ~x75 & ~x77 & ~x78 & ~x103 & ~x108 & ~x111 & ~x129 & ~x135 & ~x145 & ~x149 & ~x154 & ~x159 & ~x166 & ~x171 & ~x186 & ~x211 & ~x217 & ~x219 & ~x222 & ~x235 & ~x247 & ~x251 & ~x252 & ~x255 & ~x260 & ~x274 & ~x280 & ~x283 & ~x285 & ~x301 & ~x315 & ~x331 & ~x366 & ~x562 & ~x563 & ~x590 & ~x591 & ~x608 & ~x609 & ~x616 & ~x628 & ~x637 & ~x646 & ~x662 & ~x666 & ~x673 & ~x675 & ~x684 & ~x687 & ~x696 & ~x699 & ~x707 & ~x713 & ~x715 & ~x729 & ~x734 & ~x745 & ~x748 & ~x752 & ~x756 & ~x760 & ~x761 & ~x769 & ~x782 & ~x783;
assign c5145 =  x268 &  x356 &  x380 &  x427 & ~x159 & ~x611;
assign c5147 =  x661;
assign c5149 = ~x27 & ~x79 & ~x220 & ~x274 & ~x425 & ~x453 & ~x557 & ~x612 & ~x613 & ~x645 & ~x704;
assign c5151 =  x175;
assign c5153 =  x145;
assign c5155 =  x213 &  x276 &  x297 &  x300 &  x324 &  x325 &  x330 &  x331 &  x352 &  x353 &  x381 &  x411 &  x489;
assign c5157 =  x378 &  x380 &  x389 &  x459 &  x488 & ~x0 & ~x3 & ~x10 & ~x20 & ~x25 & ~x26 & ~x40 & ~x46 & ~x51 & ~x77 & ~x78 & ~x81 & ~x89 & ~x117 & ~x123 & ~x146 & ~x158 & ~x172 & ~x189 & ~x204 & ~x207 & ~x260 & ~x280 & ~x314 & ~x336 & ~x343 & ~x392 & ~x394 & ~x560 & ~x588 & ~x618 & ~x623 & ~x647 & ~x654 & ~x656 & ~x658 & ~x671 & ~x673 & ~x682 & ~x686 & ~x694 & ~x702 & ~x704 & ~x705 & ~x708 & ~x717 & ~x720 & ~x721 & ~x724 & ~x726 & ~x729 & ~x751 & ~x752 & ~x757 & ~x768 & ~x775 & ~x780 & ~x782;
assign c5159 =  x243 &  x274 &  x275 &  x301 &  x303 &  x325 &  x330 &  x415 &  x467 &  x494 &  x518 &  x520 & ~x150;
assign c5161 =  x248 &  x300 &  x302 &  x326 &  x328 &  x352 &  x358 &  x378 &  x379 &  x382 &  x389 &  x408 &  x438 &  x487 &  x491 &  x493 & ~x94;
assign c5163 =  x353 &  x416 &  x444 &  x445 & ~x27 & ~x35 & ~x38 & ~x48 & ~x61 & ~x62 & ~x71 & ~x75 & ~x94 & ~x105 & ~x131 & ~x132 & ~x134 & ~x138 & ~x139 & ~x141 & ~x171 & ~x174 & ~x177 & ~x180 & ~x187 & ~x188 & ~x189 & ~x206 & ~x211 & ~x217 & ~x231 & ~x234 & ~x236 & ~x247 & ~x254 & ~x272 & ~x274 & ~x282 & ~x285 & ~x300 & ~x302 & ~x337 & ~x420 & ~x532 & ~x560 & ~x562 & ~x588 & ~x605 & ~x608 & ~x611 & ~x612 & ~x613 & ~x617 & ~x618 & ~x624 & ~x629 & ~x630 & ~x636 & ~x644 & ~x646 & ~x658 & ~x670 & ~x672 & ~x682 & ~x687 & ~x690 & ~x691 & ~x699 & ~x706 & ~x709 & ~x716 & ~x743 & ~x751 & ~x753 & ~x756 & ~x765 & ~x770 & ~x772 & ~x775 & ~x778 & ~x779 & ~x781;
assign c5165 =  x11;
assign c5167 = ~x75 & ~x130 & ~x158 & ~x304 & ~x369 & ~x370 & ~x424 & ~x426 & ~x561 & ~x649 & ~x755 & ~x780;
assign c5169 =  x205;
assign c5171 =  x11;
assign c5173 =  x59;
assign c5175 =  x30;
assign c5177 =  x202;
assign c5179 =  x268 &  x328 &  x330 &  x356 &  x357 &  x358 &  x381 &  x382 &  x414 &  x434 &  x543 & ~x453;
assign c5181 =  x297 &  x445 & ~x2 & ~x11 & ~x21 & ~x22 & ~x28 & ~x29 & ~x35 & ~x43 & ~x66 & ~x69 & ~x74 & ~x75 & ~x86 & ~x88 & ~x101 & ~x108 & ~x121 & ~x133 & ~x136 & ~x143 & ~x146 & ~x157 & ~x171 & ~x173 & ~x178 & ~x192 & ~x207 & ~x211 & ~x224 & ~x226 & ~x228 & ~x237 & ~x252 & ~x253 & ~x254 & ~x260 & ~x264 & ~x265 & ~x290 & ~x308 & ~x309 & ~x316 & ~x338 & ~x339 & ~x366 & ~x569 & ~x597 & ~x602 & ~x622 & ~x625 & ~x630 & ~x644 & ~x647 & ~x665 & ~x670 & ~x672 & ~x673 & ~x678 & ~x685 & ~x691 & ~x700 & ~x709 & ~x710 & ~x717 & ~x722 & ~x750 & ~x757 & ~x760 & ~x761 & ~x770 & ~x772;
assign c5183 =  x323 &  x349 &  x350 &  x356 &  x375 &  x379 &  x384 &  x457 &  x486 & ~x77 & ~x79 & ~x106 & ~x108 & ~x160 & ~x165 & ~x166 & ~x192 & ~x217 & ~x218 & ~x705;
assign c5185 =  x88;
assign c5187 =  x269 &  x351 &  x352 &  x357 &  x379 &  x408 &  x416 &  x467 &  x491 & ~x13 & ~x18 & ~x20 & ~x22 & ~x25 & ~x30 & ~x52 & ~x55 & ~x60 & ~x61 & ~x64 & ~x77 & ~x80 & ~x86 & ~x103 & ~x106 & ~x107 & ~x120 & ~x138 & ~x147 & ~x172 & ~x173 & ~x179 & ~x234 & ~x261 & ~x310 & ~x315 & ~x339 & ~x342 & ~x369 & ~x660 & ~x672 & ~x686 & ~x699 & ~x704 & ~x723 & ~x725 & ~x733 & ~x747 & ~x758 & ~x760 & ~x761 & ~x774 & ~x780 & ~x783;
assign c5189 = ~x1 & ~x8 & ~x13 & ~x14 & ~x18 & ~x23 & ~x24 & ~x27 & ~x29 & ~x35 & ~x36 & ~x47 & ~x48 & ~x49 & ~x51 & ~x53 & ~x55 & ~x56 & ~x57 & ~x59 & ~x60 & ~x61 & ~x64 & ~x66 & ~x67 & ~x69 & ~x77 & ~x80 & ~x81 & ~x83 & ~x89 & ~x92 & ~x99 & ~x105 & ~x106 & ~x107 & ~x114 & ~x117 & ~x119 & ~x124 & ~x130 & ~x131 & ~x132 & ~x136 & ~x142 & ~x145 & ~x149 & ~x151 & ~x161 & ~x162 & ~x163 & ~x164 & ~x166 & ~x167 & ~x176 & ~x177 & ~x178 & ~x181 & ~x182 & ~x184 & ~x191 & ~x192 & ~x197 & ~x218 & ~x219 & ~x220 & ~x221 & ~x222 & ~x223 & ~x224 & ~x230 & ~x233 & ~x235 & ~x238 & ~x239 & ~x252 & ~x254 & ~x257 & ~x258 & ~x263 & ~x265 & ~x286 & ~x290 & ~x291 & ~x293 & ~x307 & ~x309 & ~x313 & ~x335 & ~x339 & ~x341 & ~x344 & ~x363 & ~x365 & ~x366 & ~x369 & ~x392 & ~x420 & ~x531 & ~x587 & ~x588 & ~x616 & ~x620 & ~x639 & ~x640 & ~x643 & ~x656 & ~x673 & ~x674 & ~x675 & ~x690 & ~x698 & ~x701 & ~x704 & ~x710 & ~x711 & ~x713 & ~x715 & ~x719 & ~x735 & ~x742 & ~x745 & ~x749 & ~x754 & ~x755 & ~x756 & ~x760 & ~x761 & ~x762 & ~x763 & ~x770 & ~x777;
assign c5191 =  x337;
assign c5193 =  x150;
assign c5195 =  x203;
assign c5197 = ~x132 & ~x329 & ~x432 & ~x436 & ~x751;
assign c5199 =  x269 &  x350 &  x354 &  x417 &  x490 & ~x10 & ~x57 & ~x67 & ~x84 & ~x108 & ~x121 & ~x142 & ~x160 & ~x168 & ~x173 & ~x207 & ~x232 & ~x260 & ~x261 & ~x288 & ~x312 & ~x664 & ~x714 & ~x724 & ~x725 & ~x746 & ~x770;
assign c5201 =  x378 & ~x189 & ~x191;
assign c5203 =  x257;
assign c5205 =  x7;
assign c5207 =  x174;
assign c5209 =  x259;
assign c5211 =  x382 &  x390 &  x418 & ~x3 & ~x4 & ~x7 & ~x9 & ~x14 & ~x15 & ~x18 & ~x22 & ~x23 & ~x25 & ~x26 & ~x27 & ~x37 & ~x39 & ~x41 & ~x42 & ~x48 & ~x54 & ~x61 & ~x64 & ~x65 & ~x68 & ~x69 & ~x73 & ~x79 & ~x80 & ~x81 & ~x82 & ~x96 & ~x108 & ~x136 & ~x137 & ~x138 & ~x139 & ~x148 & ~x151 & ~x153 & ~x159 & ~x160 & ~x164 & ~x178 & ~x179 & ~x180 & ~x181 & ~x182 & ~x186 & ~x188 & ~x191 & ~x192 & ~x193 & ~x194 & ~x197 & ~x201 & ~x210 & ~x228 & ~x232 & ~x233 & ~x258 & ~x261 & ~x262 & ~x265 & ~x282 & ~x284 & ~x289 & ~x290 & ~x338 & ~x342 & ~x365 & ~x366 & ~x535 & ~x561 & ~x562 & ~x586 & ~x587 & ~x588 & ~x589 & ~x591 & ~x593 & ~x596 & ~x598 & ~x600 & ~x618 & ~x626 & ~x629 & ~x641 & ~x646 & ~x647 & ~x648 & ~x660 & ~x663 & ~x668 & ~x669 & ~x671 & ~x674 & ~x675 & ~x679 & ~x686 & ~x693 & ~x697 & ~x701 & ~x705 & ~x706 & ~x728 & ~x729 & ~x730 & ~x733 & ~x740 & ~x747 & ~x749 & ~x750 & ~x756 & ~x757 & ~x758 & ~x760 & ~x762 & ~x763 & ~x764 & ~x770 & ~x773 & ~x778 & ~x780 & ~x781 & ~x783;
assign c5213 =  x771;
assign c5215 =  x230;
assign c5217 =  x175;
assign c5219 =  x12;
assign c5221 =  x202;
assign c5223 =  x120;
assign c5225 =  x362 &  x411 &  x418 &  x436 &  x443 & ~x31 & ~x41 & ~x46 & ~x50 & ~x53 & ~x54 & ~x72 & ~x81 & ~x83 & ~x86 & ~x91 & ~x109 & ~x139 & ~x140 & ~x159 & ~x160 & ~x179 & ~x180 & ~x185 & ~x202 & ~x206 & ~x209 & ~x210 & ~x218 & ~x237 & ~x253 & ~x265 & ~x281 & ~x284 & ~x315 & ~x337 & ~x338 & ~x340 & ~x365 & ~x560 & ~x593 & ~x597 & ~x601 & ~x607 & ~x611 & ~x618 & ~x619 & ~x623 & ~x626 & ~x627 & ~x632 & ~x633 & ~x641 & ~x645 & ~x648 & ~x649 & ~x654 & ~x658 & ~x662 & ~x663 & ~x669 & ~x676 & ~x678 & ~x685 & ~x697 & ~x702 & ~x704 & ~x705 & ~x709 & ~x711 & ~x715 & ~x722 & ~x735 & ~x749 & ~x750 & ~x755 & ~x772 & ~x783;
assign c5229 =  x200;
assign c5231 =  x406 &  x440 &  x468 &  x469 &  x496 &  x547 &  x555 & ~x10 & ~x32 & ~x90 & ~x179 & ~x197 & ~x224 & ~x230 & ~x263 & ~x283 & ~x335 & ~x337 & ~x345 & ~x370 & ~x448 & ~x690 & ~x744 & ~x757;
assign c5233 =  x375 &  x378 &  x387 &  x410 &  x417 &  x429 &  x431 &  x464 & ~x4 & ~x36 & ~x40 & ~x55 & ~x133 & ~x171 & ~x177 & ~x261 & ~x311 & ~x312 & ~x369 & ~x393 & ~x628 & ~x642 & ~x654 & ~x701 & ~x704 & ~x715;
assign c5235 =  x58;
assign c5237 =  x9;
assign c5239 =  x172;
assign c5241 =  x174;
assign c5243 =  x117;
assign c5245 = ~x193 & ~x420 & ~x482 & ~x527 & ~x533 & ~x621 & ~x732 & ~x755 & ~x775 & ~x780;
assign c5247 =  x323 &  x356 &  x379 &  x384 &  x387 &  x408 &  x467 &  x470 &  x493 &  x495 &  x501 &  x517 &  x520 &  x528 &  x529 &  x545 & ~x31 & ~x91 & ~x113 & ~x118 & ~x140 & ~x175 & ~x176 & ~x203 & ~x231 & ~x233 & ~x261 & ~x775;
assign c5249 = ~x3 & ~x13 & ~x17 & ~x22 & ~x23 & ~x25 & ~x28 & ~x35 & ~x47 & ~x56 & ~x76 & ~x81 & ~x83 & ~x85 & ~x101 & ~x105 & ~x111 & ~x118 & ~x134 & ~x135 & ~x137 & ~x144 & ~x158 & ~x163 & ~x164 & ~x166 & ~x176 & ~x189 & ~x193 & ~x219 & ~x229 & ~x232 & ~x248 & ~x255 & ~x256 & ~x272 & ~x275 & ~x282 & ~x301 & ~x303 & ~x307 & ~x310 & ~x328 & ~x329 & ~x342 & ~x357 & ~x369 & ~x370 & ~x611 & ~x639 & ~x672 & ~x699 & ~x701 & ~x723 & ~x724 & ~x725 & ~x726 & ~x731 & ~x753 & ~x755 & ~x758 & ~x782;
assign c5251 =  x351 &  x381 &  x385 &  x388 &  x405 &  x415 &  x434 &  x439 &  x443 &  x444 &  x464 &  x465 & ~x10 & ~x11 & ~x22 & ~x28 & ~x39 & ~x50 & ~x60 & ~x68 & ~x79 & ~x81 & ~x95 & ~x102 & ~x109 & ~x112 & ~x115 & ~x149 & ~x151 & ~x154 & ~x161 & ~x171 & ~x172 & ~x174 & ~x175 & ~x201 & ~x209 & ~x210 & ~x217 & ~x221 & ~x225 & ~x229 & ~x234 & ~x253 & ~x287 & ~x309 & ~x310 & ~x336 & ~x392 & ~x560 & ~x591 & ~x614 & ~x617 & ~x619 & ~x627 & ~x631 & ~x638 & ~x644 & ~x645 & ~x650 & ~x651 & ~x655 & ~x662 & ~x670 & ~x685 & ~x702 & ~x706 & ~x724 & ~x726 & ~x733 & ~x745 & ~x750 & ~x768 & ~x771 & ~x774 & ~x781;
assign c5253 =  x14;
assign c5255 = ~x14 & ~x21 & ~x74 & ~x81 & ~x87 & ~x184 & ~x481 & ~x562 & ~x618 & ~x667 & ~x779;
assign c5257 = ~x7 & ~x80 & ~x81 & ~x104 & ~x107 & ~x110 & ~x114 & ~x134 & ~x160 & ~x193 & ~x242 & ~x243 & ~x271 & ~x327 & ~x342 & ~x343 & ~x365 & ~x369 & ~x494 & ~x612 & ~x613 & ~x673 & ~x674 & ~x675 & ~x695 & ~x730 & ~x752;
assign c5259 =  x388 &  x414 &  x439 &  x440 &  x441 &  x445 & ~x5 & ~x12 & ~x18 & ~x21 & ~x36 & ~x52 & ~x57 & ~x61 & ~x73 & ~x80 & ~x89 & ~x119 & ~x137 & ~x143 & ~x161 & ~x174 & ~x199 & ~x210 & ~x260 & ~x265 & ~x278 & ~x281 & ~x284 & ~x288 & ~x292 & ~x309 & ~x312 & ~x318 & ~x338 & ~x363 & ~x743 & ~x746;
assign c5261 = ~x1 & ~x5 & ~x48 & ~x81 & ~x105 & ~x142 & ~x167 & ~x224 & ~x273 & ~x279 & ~x303 & ~x330 & ~x369 & ~x371 & ~x448 & ~x531 & ~x532 & ~x559 & ~x638 & ~x639 & ~x640 & ~x666 & ~x673 & ~x697 & ~x699 & ~x703 & ~x724 & ~x733 & ~x758 & ~x761;
assign c5263 =  x298 &  x633;
assign c5265 =  x323 &  x361 &  x408 &  x466 &  x473 &  x491 &  x529 & ~x5 & ~x25 & ~x96 & ~x179 & ~x252 & ~x420 & ~x643 & ~x693 & ~x716 & ~x717;
assign c5267 =  x55;
assign c5269 =  x13;
assign c5271 =  x42;
assign c5273 =  x202;
assign c5275 =  x607 &  x671;
assign c5277 = ~x0 & ~x20 & ~x25 & ~x31 & ~x52 & ~x59 & ~x77 & ~x82 & ~x90 & ~x108 & ~x111 & ~x112 & ~x113 & ~x122 & ~x133 & ~x152 & ~x164 & ~x168 & ~x171 & ~x179 & ~x224 & ~x226 & ~x230 & ~x284 & ~x341 & ~x424 & ~x426 & ~x427 & ~x452 & ~x453 & ~x587 & ~x588 & ~x605 & ~x641 & ~x645 & ~x652 & ~x655 & ~x659 & ~x662 & ~x674 & ~x687 & ~x697 & ~x698 & ~x704 & ~x709 & ~x716 & ~x719 & ~x722 & ~x726 & ~x730 & ~x733 & ~x766 & ~x769 & ~x774 & ~x776 & ~x777;
assign c5279 = ~x165 & ~x192 & ~x453 & ~x528 & ~x549 & ~x610 & ~x731;
assign c5281 =  x716;
assign c5283 =  x330 &  x353 &  x383 &  x494 &  x498 &  x573 &  x575 &  x576 &  x581 &  x583 & ~x761;
assign c5285 =  x120;
assign c5287 =  x11;
assign c5289 =  x320 &  x373 &  x385 &  x390 & ~x85 & ~x245 & ~x256 & ~x301 & ~x585 & ~x613;
assign c5291 =  x56;
assign c5293 =  x560;
assign c5295 = ~x2 & ~x31 & ~x76 & ~x135 & ~x139 & ~x169 & ~x192 & ~x221 & ~x226 & ~x250 & ~x300 & ~x310 & ~x336 & ~x338 & ~x343 & ~x367 & ~x392 & ~x495 & ~x505 & ~x598 & ~x649 & ~x654 & ~x680 & ~x759;
assign c5297 = ~x453 & ~x485 & ~x542 & ~x549;
assign c5299 =  x346 &  x355 &  x372 & ~x107 & ~x134 & ~x136 & ~x162 & ~x245 & ~x251 & ~x274 & ~x302 & ~x584 & ~x585 & ~x618;
assign c5301 =  x113;
assign c5303 =  x43;
assign c5305 =  x167;
assign c5307 =  x771;
assign c5309 =  x22 &  x112;
assign c5311 =  x325 &  x358 &  x552 & ~x538;
assign c5313 =  x12;
assign c5315 =  x140;
assign c5317 =  x86;
assign c5321 =  x390 &  x408 &  x433 & ~x155 & ~x209 & ~x365 & ~x369 & ~x563 & ~x638 & ~x693 & ~x730 & ~x780;
assign c5323 =  x275 &  x297 &  x302 &  x606;
assign c5325 =  x12;
assign c5327 =  x282;
assign c5329 =  x146;
assign c5331 =  x441 &  x606 & ~x334 & ~x362 & ~x390;
assign c5333 = ~x301 & ~x530;
assign c5335 = ~x5 & ~x23 & ~x32 & ~x57 & ~x80 & ~x81 & ~x136 & ~x159 & ~x170 & ~x183 & ~x200 & ~x207 & ~x218 & ~x279 & ~x281 & ~x300 & ~x392 & ~x424 & ~x425 & ~x426 & ~x598 & ~x628 & ~x639 & ~x642 & ~x649 & ~x654 & ~x657 & ~x659 & ~x688 & ~x697 & ~x724 & ~x735 & ~x756 & ~x766;
assign c5337 =  x225;
assign c5339 =  x346 &  x349 &  x354 &  x372 &  x399 &  x422 &  x427 & ~x162 & ~x210 & ~x217 & ~x246;
assign c5341 =  x118;
assign c5343 =  x354 &  x356 &  x358 &  x385 &  x386 &  x406 &  x407 &  x409 &  x411 &  x413 &  x463 &  x489 &  x493 &  x518 &  x519 & ~x1 & ~x9 & ~x13 & ~x19 & ~x31 & ~x34 & ~x35 & ~x37 & ~x143 & ~x147 & ~x167 & ~x170 & ~x198 & ~x229 & ~x233 & ~x284 & ~x310 & ~x311 & ~x393 & ~x425 & ~x690 & ~x716 & ~x717 & ~x746 & ~x760;
assign c5345 =  x328 &  x331 &  x382 &  x470 &  x494 &  x517 & ~x42 & ~x112 & ~x123 & ~x149 & ~x234 & ~x251 & ~x372 & ~x397 & ~x400 & ~x451 & ~x453 & ~x749 & ~x763 & ~x767;
assign c5347 =  x204;
assign c5349 =  x213 &  x325 &  x326 &  x329 &  x351 &  x354 &  x355 &  x383 &  x384 &  x385 &  x386 &  x410 &  x439 &  x461 & ~x35 & ~x90 & ~x119 & ~x335 & ~x343 & ~x392;
assign c5351 =  x245 &  x301 &  x330 &  x352 &  x353 &  x357 &  x381 &  x387 &  x441 &  x489 &  x522 & ~x205 & ~x289 & ~x371 & ~x426;
assign c5353 =  x268 &  x297 &  x591;
assign c5355 =  x11 &  x63;
assign c5357 =  x302 &  x326 &  x329 &  x330 &  x331 &  x352 &  x357 &  x378 &  x380 &  x415 &  x489 &  x548 & ~x425;
assign c5359 =  x66;
assign c5361 =  x364;
assign c5363 =  x323 &  x324 &  x350 &  x353 &  x376 &  x377 &  x379 &  x380 &  x404 &  x410 &  x414 &  x416 &  x433 &  x435 &  x444 & ~x4 & ~x7 & ~x11 & ~x29 & ~x30 & ~x33 & ~x38 & ~x48 & ~x51 & ~x52 & ~x59 & ~x61 & ~x64 & ~x78 & ~x79 & ~x81 & ~x107 & ~x131 & ~x139 & ~x160 & ~x187 & ~x192 & ~x202 & ~x226 & ~x254 & ~x420 & ~x622 & ~x624 & ~x626 & ~x635 & ~x641 & ~x651 & ~x669 & ~x671 & ~x675 & ~x688 & ~x695 & ~x703 & ~x707 & ~x716 & ~x722 & ~x728 & ~x731 & ~x755 & ~x768 & ~x770 & ~x771;
assign c5365 =  x252;
assign c5367 =  x755;
assign c5369 =  x309;
assign c5371 =  x118;
assign c5373 =  x242 &  x298 &  x300 &  x328 &  x329 &  x330 &  x351 &  x356 &  x416 &  x492 &  x493 &  x518 & ~x27 & ~x92 & ~x93 & ~x138 & ~x167 & ~x198 & ~x230 & ~x260 & ~x284 & ~x288 & ~x316 & ~x344 & ~x368 & ~x369 & ~x370 & ~x689 & ~x690 & ~x691 & ~x744 & ~x745 & ~x758;
assign c5375 =  x303 &  x351 &  x381 &  x385 &  x387 &  x411 &  x462 &  x467 &  x493 &  x519 & ~x141 & ~x257 & ~x289 & ~x397 & ~x398 & ~x691 & ~x718;
assign c5377 =  x39 &  x280;
assign c5379 =  x11;
assign c5381 =  x58;
assign c5383 =  x226;
assign c5385 = ~x33 & ~x53 & ~x155 & ~x246 & ~x247 & ~x302 & ~x483 & ~x520 & ~x639 & ~x667 & ~x684 & ~x686;
assign c5387 =  x772;
assign c5389 =  x32;
assign c5391 =  x351 &  x352 &  x353 &  x354 &  x356 &  x360 &  x361 &  x380 &  x384 &  x385 &  x407 &  x408 &  x445 &  x489 &  x492 &  x514 &  x516 &  x520 &  x528 & ~x7 & ~x29 & ~x143 & ~x147 & ~x149 & ~x261 & ~x308 & ~x342 & ~x368 & ~x369 & ~x690 & ~x744;
assign c5393 =  x146;
assign c5395 =  x42 & ~x530;
assign c5397 =  x230;
assign c5399 =  x778;
assign c5401 =  x716;
assign c5403 =  x268 &  x275 &  x324 &  x331 &  x357 &  x360 &  x378 &  x435 &  x444 &  x488 &  x489 & ~x0 & ~x262;
assign c5405 = ~x25 & ~x50 & ~x184 & ~x206 & ~x236 & ~x250 & ~x255 & ~x275 & ~x302 & ~x315 & ~x317 & ~x338 & ~x478 & ~x603 & ~x613 & ~x633 & ~x646 & ~x672 & ~x676 & ~x679 & ~x708 & ~x739 & ~x768 & ~x774;
assign c5407 =  x196;
assign c5409 =  x273 &  x330 &  x358 &  x441 &  x544 & ~x402;
assign c5411 =  x329 &  x351 &  x355 &  x359 &  x378 &  x384 &  x405 &  x411 &  x414 &  x415 &  x438 &  x487 &  x488 &  x489 &  x493 & ~x0 & ~x12 & ~x26 & ~x65 & ~x66 & ~x87 & ~x140 & ~x143 & ~x144 & ~x145 & ~x199 & ~x206 & ~x228 & ~x233 & ~x259 & ~x280 & ~x281 & ~x315 & ~x343 & ~x369 & ~x504 & ~x689 & ~x690 & ~x772;
assign c5413 =  x297 &  x390 &  x418 &  x446 &  x472 & ~x11 & ~x12 & ~x21 & ~x26 & ~x48 & ~x55 & ~x66 & ~x86 & ~x102 & ~x106 & ~x109 & ~x110 & ~x112 & ~x121 & ~x177 & ~x185 & ~x211 & ~x238 & ~x254 & ~x309 & ~x314 & ~x335 & ~x342 & ~x366 & ~x560 & ~x600 & ~x606 & ~x607 & ~x612 & ~x624 & ~x638 & ~x640 & ~x649 & ~x654 & ~x657 & ~x660 & ~x667 & ~x697 & ~x698 & ~x708 & ~x721 & ~x729 & ~x743 & ~x747 & ~x757 & ~x779;
assign c5415 =  x272 &  x298 &  x302 &  x325 &  x331 &  x387 &  x407 &  x489 &  x546 &  x598 & ~x455;
assign c5417 =  x226;
assign c5419 =  x417 &  x445 & ~x6 & ~x11 & ~x54 & ~x61 & ~x64 & ~x71 & ~x78 & ~x82 & ~x90 & ~x91 & ~x101 & ~x102 & ~x112 & ~x119 & ~x131 & ~x134 & ~x138 & ~x140 & ~x141 & ~x149 & ~x150 & ~x151 & ~x155 & ~x160 & ~x163 & ~x165 & ~x173 & ~x191 & ~x198 & ~x223 & ~x227 & ~x235 & ~x244 & ~x246 & ~x254 & ~x265 & ~x285 & ~x286 & ~x300 & ~x301 & ~x316 & ~x342 & ~x365 & ~x392 & ~x393 & ~x394 & ~x532 & ~x533 & ~x561 & ~x600 & ~x614 & ~x638 & ~x648 & ~x650 & ~x651 & ~x653 & ~x657 & ~x663 & ~x681 & ~x695 & ~x700 & ~x721 & ~x723 & ~x732 & ~x736 & ~x737 & ~x744 & ~x758 & ~x771 & ~x775;
assign c5421 =  x320 &  x388 &  x403 &  x429 &  x432 &  x442 &  x443 & ~x2 & ~x53 & ~x71 & ~x161 & ~x174 & ~x201 & ~x209 & ~x251 & ~x596 & ~x598 & ~x649 & ~x667 & ~x694 & ~x746 & ~x782;
assign c5423 =  x690 & ~x473;
assign c5425 = ~x424 & ~x474 & ~x501 & ~x528;
assign c5427 =  x35;
assign c5429 =  x201;
assign c5431 =  x352 &  x378 &  x432 &  x437 &  x445 &  x462 &  x492 &  x493 & ~x7 & ~x15 & ~x21 & ~x25 & ~x26 & ~x32 & ~x40 & ~x70 & ~x82 & ~x96 & ~x104 & ~x171 & ~x173 & ~x194 & ~x195 & ~x201 & ~x224 & ~x234 & ~x364 & ~x369 & ~x392 & ~x664 & ~x713 & ~x725 & ~x728 & ~x732 & ~x735 & ~x736 & ~x755 & ~x756 & ~x765;
assign c5433 =  x304 &  x352 &  x411 &  x412 &  x415 &  x416 &  x439 &  x442 &  x465 & ~x6 & ~x24 & ~x36 & ~x57 & ~x87 & ~x114 & ~x232 & ~x254 & ~x259 & ~x335 & ~x343 & ~x369 & ~x393 & ~x420 & ~x717 & ~x779;
assign c5435 =  x354 &  x385 &  x464 &  x469 &  x494 &  x523 & ~x263 & ~x399 & ~x744;
assign c5437 =  x270 &  x271 &  x273 &  x328 &  x409 &  x414 &  x437 &  x466 &  x467 &  x495 &  x517 & ~x401;
assign c5439 =  x298 &  x323 &  x324 &  x332 &  x352 &  x354 &  x356 &  x358 &  x376 &  x379 &  x381 &  x384 &  x385 &  x387 &  x405 &  x410 &  x413 &  x417 &  x434 &  x437 &  x445 &  x460 &  x461 & ~x4 & ~x7 & ~x30 & ~x36 & ~x38 & ~x55 & ~x60 & ~x63 & ~x66 & ~x94 & ~x119 & ~x138 & ~x143 & ~x149 & ~x168 & ~x169 & ~x177 & ~x196 & ~x199 & ~x200 & ~x202 & ~x225 & ~x227 & ~x252 & ~x281 & ~x311 & ~x662 & ~x717;
assign c5441 =  x296 &  x353 &  x379 &  x406 &  x409 &  x433 &  x439 &  x462 &  x463 &  x464 &  x465 &  x486 &  x490 & ~x5 & ~x6 & ~x17 & ~x21 & ~x22 & ~x25 & ~x30 & ~x32 & ~x34 & ~x45 & ~x46 & ~x58 & ~x61 & ~x66 & ~x78 & ~x87 & ~x91 & ~x98 & ~x112 & ~x118 & ~x146 & ~x166 & ~x169 & ~x178 & ~x196 & ~x197 & ~x202 & ~x281 & ~x311 & ~x313 & ~x336 & ~x342 & ~x343 & ~x366 & ~x370 & ~x393 & ~x660 & ~x689 & ~x716 & ~x729 & ~x742 & ~x755 & ~x764 & ~x766 & ~x767 & ~x773 & ~x774 & ~x783;
assign c5443 =  x296 &  x297 &  x300 &  x330 &  x352 &  x379 &  x386 &  x405 &  x406 &  x434 &  x436 &  x461 &  x492 &  x493 &  x516 &  x517 &  x520 &  x521 & ~x36 & ~x150 & ~x230 & ~x289 & ~x312 & ~x369 & ~x370 & ~x371;
assign c5445 = ~x163 & ~x359 & ~x416 & ~x443 & ~x725;
assign c5447 =  x336;
assign c5449 =  x439 &  x462 & ~x4 & ~x14 & ~x25 & ~x26 & ~x30 & ~x44 & ~x55 & ~x58 & ~x62 & ~x69 & ~x93 & ~x94 & ~x147 & ~x149 & ~x150 & ~x154 & ~x161 & ~x162 & ~x169 & ~x171 & ~x205 & ~x212 & ~x230 & ~x238 & ~x239 & ~x251 & ~x257 & ~x259 & ~x264 & ~x265 & ~x266 & ~x311 & ~x316 & ~x337 & ~x370 & ~x392 & ~x394 & ~x643 & ~x646 & ~x703 & ~x716 & ~x722 & ~x730 & ~x731 & ~x759 & ~x764;
assign c5451 =  x325 &  x351 &  x417 &  x445 & ~x10 & ~x34 & ~x60 & ~x78 & ~x83 & ~x89 & ~x92 & ~x93 & ~x104 & ~x105 & ~x106 & ~x109 & ~x121 & ~x139 & ~x146 & ~x175 & ~x199 & ~x201 & ~x206 & ~x314 & ~x370 & ~x392 & ~x393 & ~x420 & ~x649 & ~x652 & ~x675 & ~x732 & ~x741 & ~x745 & ~x754 & ~x771 & ~x772;
assign c5453 =  x58;
assign c5455 =  x117;
assign c5457 =  x308;
assign c5459 =  x418 & ~x6 & ~x10 & ~x11 & ~x12 & ~x14 & ~x20 & ~x21 & ~x25 & ~x26 & ~x28 & ~x31 & ~x32 & ~x33 & ~x35 & ~x36 & ~x44 & ~x48 & ~x50 & ~x54 & ~x55 & ~x61 & ~x74 & ~x75 & ~x77 & ~x80 & ~x81 & ~x85 & ~x87 & ~x88 & ~x89 & ~x90 & ~x91 & ~x101 & ~x104 & ~x106 & ~x107 & ~x109 & ~x113 & ~x119 & ~x121 & ~x123 & ~x126 & ~x132 & ~x133 & ~x136 & ~x139 & ~x141 & ~x144 & ~x151 & ~x152 & ~x153 & ~x155 & ~x163 & ~x166 & ~x174 & ~x178 & ~x182 & ~x183 & ~x185 & ~x194 & ~x200 & ~x201 & ~x208 & ~x211 & ~x215 & ~x216 & ~x217 & ~x218 & ~x219 & ~x221 & ~x226 & ~x230 & ~x231 & ~x233 & ~x238 & ~x246 & ~x254 & ~x255 & ~x258 & ~x263 & ~x281 & ~x287 & ~x290 & ~x302 & ~x310 & ~x311 & ~x314 & ~x315 & ~x316 & ~x329 & ~x336 & ~x337 & ~x338 & ~x340 & ~x341 & ~x365 & ~x504 & ~x532 & ~x533 & ~x560 & ~x561 & ~x562 & ~x564 & ~x585 & ~x587 & ~x589 & ~x590 & ~x591 & ~x593 & ~x596 & ~x599 & ~x604 & ~x617 & ~x625 & ~x627 & ~x628 & ~x633 & ~x635 & ~x636 & ~x638 & ~x641 & ~x648 & ~x650 & ~x651 & ~x653 & ~x655 & ~x659 & ~x660 & ~x661 & ~x663 & ~x668 & ~x674 & ~x675 & ~x676 & ~x678 & ~x686 & ~x695 & ~x696 & ~x697 & ~x701 & ~x705 & ~x706 & ~x714 & ~x727 & ~x730 & ~x739 & ~x743 & ~x747 & ~x748 & ~x749 & ~x757 & ~x759 & ~x760 & ~x764 & ~x765 & ~x766 & ~x768 & ~x770 & ~x773 & ~x781;
assign c5461 =  x351 &  x352 &  x376 &  x410 &  x411 &  x437 &  x443 &  x444 &  x464 &  x472 &  x473 &  x486 &  x491 &  x494 & ~x2 & ~x10 & ~x14 & ~x34 & ~x84 & ~x113 & ~x177 & ~x195 & ~x227 & ~x228 & ~x230 & ~x289 & ~x314 & ~x317 & ~x342 & ~x344 & ~x367 & ~x368 & ~x369 & ~x370 & ~x420 & ~x760 & ~x769;
assign c5463 =  x227;
assign c5465 =  x257;
assign c5467 =  x325 &  x351 &  x352 &  x407 &  x411 &  x413 &  x414 &  x460 & ~x0 & ~x13 & ~x24 & ~x25 & ~x31 & ~x58 & ~x61 & ~x85 & ~x91 & ~x98 & ~x112 & ~x113 & ~x121 & ~x128 & ~x155 & ~x163 & ~x170 & ~x232 & ~x264 & ~x283 & ~x286 & ~x289 & ~x311 & ~x315 & ~x366 & ~x368 & ~x392 & ~x589 & ~x628 & ~x671 & ~x673 & ~x692 & ~x694 & ~x704 & ~x705 & ~x719 & ~x760 & ~x766 & ~x770 & ~x782;
assign c5469 =  x244 &  x245 &  x268 &  x275 &  x299 &  x300 &  x328 &  x414 &  x437 & ~x344 & ~x400;
assign c5471 = ~x219 & ~x485 & ~x494 & ~x543 & ~x677;
assign c5473 =  x380 &  x388 &  x466 &  x473 &  x493 &  x495 & ~x30 & ~x55 & ~x57 & ~x68 & ~x77 & ~x78 & ~x96 & ~x106 & ~x113 & ~x173 & ~x224 & ~x262 & ~x289 & ~x343 & ~x396 & ~x397 & ~x398 & ~x532 & ~x661 & ~x702 & ~x731 & ~x734 & ~x756;
assign c5475 =  x331 &  x332 &  x353 &  x359 &  x408 &  x445 &  x461 &  x496 & ~x178 & ~x452 & ~x453;
assign c5477 =  x230;
assign c5479 =  x351 &  x378 &  x379 &  x381 &  x383 &  x387 &  x411 &  x433 &  x441 &  x467 &  x473 &  x556 & ~x8 & ~x20 & ~x32 & ~x35 & ~x87 & ~x89 & ~x168 & ~x224 & ~x257 & ~x261 & ~x262 & ~x661 & ~x705 & ~x706 & ~x715 & ~x730 & ~x737 & ~x751 & ~x756;
assign c5481 =  x269 &  x351 &  x354 &  x376 &  x383 &  x384 &  x417 &  x486 &  x488 &  x493 &  x494 & ~x13 & ~x18 & ~x27 & ~x31 & ~x40 & ~x52 & ~x54 & ~x79 & ~x84 & ~x86 & ~x87 & ~x90 & ~x114 & ~x138 & ~x147 & ~x170 & ~x173 & ~x174 & ~x177 & ~x194 & ~x224 & ~x228 & ~x230 & ~x261 & ~x309 & ~x365 & ~x392 & ~x660 & ~x661 & ~x662 & ~x674 & ~x689 & ~x702 & ~x715 & ~x717 & ~x725 & ~x748 & ~x751 & ~x754 & ~x763 & ~x766 & ~x772 & ~x781;
assign c5483 =  x36;
assign c5485 =  x463 &  x489 &  x514 &  x579 & ~x107 & ~x163 & ~x192 & ~x278;
assign c5487 = ~x0 & ~x79 & ~x105 & ~x107 & ~x131 & ~x132 & ~x163 & ~x166 & ~x191 & ~x367 & ~x369 & ~x425 & ~x453 & ~x455 & ~x563 & ~x639 & ~x669 & ~x680 & ~x725 & ~x737 & ~x775;
assign c5489 =  x244 &  x245 &  x247 &  x303 &  x325 &  x328 &  x329 &  x356 &  x358 &  x381 &  x407 &  x415 &  x461 &  x517 &  x518 &  x520;
assign c5491 =  x364;
assign c5493 = ~x59 & ~x135 & ~x144 & ~x189 & ~x219 & ~x220 & ~x222 & ~x249 & ~x302 & ~x338 & ~x364 & ~x480 & ~x614 & ~x641 & ~x702 & ~x724 & ~x765;
assign c5495 =  x42;
assign c5497 =  x299 &  x330 &  x352 &  x355 &  x386 &  x410 &  x437 &  x468 &  x470 &  x472 &  x488 &  x495 &  x496 &  x518 &  x522 & ~x205 & ~x288 & ~x476 & ~x690 & ~x718 & ~x760 & ~x781;
assign c5499 = ~x219 & ~x243 & ~x317 & ~x421 & ~x500;
assign c60 =  x234 &  x266 &  x267 &  x323 &  x354 &  x438 &  x439 &  x457 &  x463 &  x543 &  x572 &  x596 &  x597 &  x603 &  x604 &  x633 &  x682 & ~x1 & ~x20 & ~x53 & ~x55 & ~x83 & ~x84 & ~x86 & ~x165 & ~x199 & ~x221 & ~x250 & ~x278 & ~x388 & ~x392 & ~x394 & ~x559 & ~x590 & ~x593 & ~x641 & ~x642 & ~x646 & ~x672 & ~x673 & ~x696 & ~x726 & ~x728 & ~x729 & ~x757 & ~x779;
assign c62 =  x75 &  x574 & ~x31 & ~x55 & ~x143 & ~x338 & ~x394 & ~x414 & ~x421 & ~x471 & ~x557 & ~x593 & ~x754 & ~x758 & ~x762 & ~x765 & ~x782;
assign c64 =  x339 & ~x3 & ~x169 & ~x279 & ~x760;
assign c66 =  x49 &  x525 & ~x762;
assign c68 =  x231 &  x301 &  x387 &  x413 & ~x20 & ~x28 & ~x30 & ~x56 & ~x57 & ~x82 & ~x83 & ~x85 & ~x113 & ~x115 & ~x137 & ~x138 & ~x166 & ~x167 & ~x193 & ~x194 & ~x221 & ~x222 & ~x223 & ~x225 & ~x250 & ~x279 & ~x281 & ~x306 & ~x307 & ~x308 & ~x309 & ~x334 & ~x335 & ~x420 & ~x448 & ~x449 & ~x476 & ~x615 & ~x728 & ~x729 & ~x757 & ~x763 & ~x764 & ~x779 & ~x783;
assign c610 = ~x2 & ~x17 & ~x45 & ~x46 & ~x279 & ~x307 & ~x447 & ~x467 & ~x674 & ~x757;
assign c612 =  x303 &  x315 &  x371 & ~x111 & ~x138 & ~x140 & ~x142 & ~x164 & ~x194 & ~x196 & ~x279 & ~x502 & ~x531 & ~x727 & ~x731 & ~x753 & ~x755 & ~x761 & ~x780 & ~x783;
assign c614 = ~x7 & ~x8 & ~x29 & ~x57 & ~x109 & ~x141 & ~x165 & ~x167 & ~x171 & ~x249 & ~x295 & ~x306 & ~x337 & ~x392 & ~x474 & ~x477 & ~x502 & ~x505 & ~x541 & ~x588 & ~x617 & ~x701 & ~x730 & ~x756;
assign c616 = ~x27 & ~x109 & ~x136 & ~x169 & ~x176 & ~x414 & ~x534 & ~x555 & ~x556 & ~x591 & ~x592 & ~x621 & ~x696;
assign c618 = ~x2 & ~x3 & ~x6 & ~x47 & ~x52 & ~x74 & ~x80 & ~x109 & ~x167 & ~x194 & ~x240 & ~x255 & ~x338 & ~x475 & ~x502 & ~x505 & ~x532 & ~x559 & ~x643 & ~x699 & ~x727 & ~x775 & ~x776 & ~x781;
assign c620 =  x339 & ~x167 & ~x223 & ~x308;
assign c622 =  x95 &  x241 &  x269 &  x320 &  x343 &  x346 &  x376 &  x377 &  x387 &  x414 &  x434 &  x437 &  x457 &  x490 &  x599 &  x604 &  x628 &  x632 &  x636 & ~x6 & ~x31 & ~x87 & ~x116 & ~x169 & ~x192 & ~x195 & ~x254 & ~x278 & ~x307 & ~x333 & ~x335 & ~x421 & ~x449 & ~x672;
assign c624 = ~x1 & ~x2 & ~x22 & ~x27 & ~x53 & ~x54 & ~x57 & ~x136 & ~x166 & ~x168 & ~x184 & ~x195 & ~x221 & ~x222 & ~x279 & ~x280 & ~x282 & ~x306 & ~x360 & ~x362 & ~x421 & ~x473 & ~x503 & ~x506 & ~x530 & ~x531 & ~x533 & ~x558 & ~x561 & ~x589 & ~x616 & ~x646 & ~x672 & ~x683 & ~x701 & ~x727 & ~x729 & ~x755;
assign c626 = ~x4 & ~x12 & ~x16 & ~x22 & ~x24 & ~x31 & ~x33 & ~x51 & ~x56 & ~x80 & ~x83 & ~x84 & ~x110 & ~x113 & ~x167 & ~x169 & ~x170 & ~x198 & ~x225 & ~x226 & ~x282 & ~x305 & ~x307 & ~x308 & ~x362 & ~x365 & ~x418 & ~x474 & ~x505 & ~x514 & ~x530 & ~x533 & ~x587 & ~x646 & ~x671 & ~x672 & ~x727 & ~x755;
assign c628 =  x345 &  x573 &  x652 & ~x3 & ~x7 & ~x20 & ~x21 & ~x22 & ~x24 & ~x28 & ~x29 & ~x31 & ~x52 & ~x60 & ~x88 & ~x110 & ~x144 & ~x169 & ~x172 & ~x198 & ~x223 & ~x225 & ~x248 & ~x337 & ~x338 & ~x363 & ~x365 & ~x387 & ~x394 & ~x417 & ~x425 & ~x448 & ~x451 & ~x452 & ~x454 & ~x472 & ~x480 & ~x502 & ~x504 & ~x528 & ~x529 & ~x531 & ~x534 & ~x555 & ~x558 & ~x562 & ~x584 & ~x588 & ~x610 & ~x638 & ~x646 & ~x667 & ~x674 & ~x676 & ~x697 & ~x698 & ~x702 & ~x705 & ~x728 & ~x730 & ~x733 & ~x751 & ~x760 & ~x761 & ~x781;
assign c630 =  x369 & ~x29 & ~x251 & ~x621 & ~x667 & ~x725;
assign c632 = ~x234 & ~x545 & ~x751;
assign c634 =  x287 &  x747 & ~x4 & ~x60 & ~x83 & ~x87 & ~x167 & ~x253 & ~x291 & ~x335 & ~x451 & ~x477 & ~x478 & ~x505 & ~x533 & ~x617 & ~x672 & ~x675 & ~x765;
assign c636 = ~x17 & ~x51 & ~x84 & ~x170 & ~x221 & ~x250 & ~x251 & ~x282 & ~x361 & ~x363 & ~x376 & ~x390 & ~x504 & ~x704 & ~x732 & ~x752 & ~x754;
assign c638 =  x36 &  x216 &  x317 &  x411 &  x427 & ~x2 & ~x15 & ~x24 & ~x28 & ~x59 & ~x110 & ~x136 & ~x141 & ~x142 & ~x170 & ~x193 & ~x195 & ~x196 & ~x225 & ~x308 & ~x336 & ~x363 & ~x364 & ~x365 & ~x391 & ~x475 & ~x756 & ~x757 & ~x782;
assign c640 =  x13 &  x15 &  x67 &  x104 &  x132 &  x178 &  x179 &  x203 &  x210 &  x212 &  x215 &  x242 &  x317 &  x495 &  x541 &  x599 &  x630 &  x632 &  x655 &  x657 & ~x18 & ~x20 & ~x86 & ~x108 & ~x166 & ~x227 & ~x254 & ~x278 & ~x309 & ~x419 & ~x474;
assign c642 =  x311 & ~x731;
assign c644 =  x35 &  x463 &  x482 & ~x83;
assign c646 = ~x11 & ~x27 & ~x83 & ~x169 & ~x238 & ~x350 & ~x378 & ~x532;
assign c648 =  x226;
assign c650 =  x268 &  x316 &  x437 &  x651 & ~x171 & ~x392 & ~x479 & ~x526 & ~x537 & ~x675 & ~x696 & ~x760;
assign c652 =  x15 &  x543 & ~x20 & ~x46 & ~x52 & ~x60 & ~x85 & ~x139 & ~x223 & ~x309 & ~x446 & ~x477 & ~x530 & ~x559 & ~x730 & ~x764;
assign c654 =  x260 &  x272 &  x686 &  x714 & ~x2 & ~x34 & ~x38 & ~x46 & ~x60 & ~x109 & ~x309 & ~x389 & ~x748 & ~x759;
assign c656 =  x146 &  x202 &  x742 & ~x5 & ~x10 & ~x20 & ~x21 & ~x22 & ~x32 & ~x33 & ~x36 & ~x37 & ~x51 & ~x61 & ~x88 & ~x112 & ~x143 & ~x144 & ~x167 & ~x198 & ~x252 & ~x279 & ~x307 & ~x335 & ~x337 & ~x361 & ~x365 & ~x422 & ~x448 & ~x450 & ~x531 & ~x532 & ~x586 & ~x757 & ~x776;
assign c658 = ~x17 & ~x122 & ~x248 & ~x392 & ~x411;
assign c660 =  x95 &  x263 &  x294 &  x318 &  x462 &  x518 & ~x27 & ~x59 & ~x79 & ~x86 & ~x108 & ~x109 & ~x111 & ~x146 & ~x173 & ~x202 & ~x249 & ~x250 & ~x253 & ~x255 & ~x278 & ~x307 & ~x333 & ~x366 & ~x391 & ~x478 & ~x504 & ~x561 & ~x587 & ~x615 & ~x618 & ~x619 & ~x670 & ~x729 & ~x756 & ~x782;
assign c662 =  x161 &  x746 & ~x9 & ~x17 & ~x27 & ~x35 & ~x37 & ~x46 & ~x82 & ~x86 & ~x136 & ~x168 & ~x224 & ~x473 & ~x533 & ~x588 & ~x757 & ~x758;
assign c664 =  x103 &  x129 &  x234 &  x297 &  x326 &  x327 &  x569 &  x624 &  x657 & ~x9 & ~x10 & ~x22 & ~x24 & ~x30 & ~x35 & ~x87 & ~x113 & ~x138 & ~x141 & ~x167 & ~x171 & ~x256 & ~x275 & ~x279 & ~x332 & ~x361 & ~x364 & ~x392 & ~x417 & ~x504 & ~x585 & ~x587 & ~x642 & ~x702 & ~x727;
assign c666 = ~x1 & ~x172 & ~x422 & ~x488 & ~x589 & ~x749;
assign c668 = ~x6 & ~x21 & ~x22 & ~x27 & ~x28 & ~x31 & ~x54 & ~x59 & ~x81 & ~x83 & ~x86 & ~x87 & ~x141 & ~x167 & ~x194 & ~x223 & ~x225 & ~x227 & ~x248 & ~x253 & ~x276 & ~x282 & ~x283 & ~x305 & ~x307 & ~x310 & ~x331 & ~x361 & ~x362 & ~x388 & ~x391 & ~x392 & ~x394 & ~x421 & ~x425 & ~x447 & ~x448 & ~x450 & ~x472 & ~x500 & ~x503 & ~x504 & ~x505 & ~x530 & ~x533 & ~x559 & ~x560 & ~x561 & ~x563 & ~x587 & ~x589 & ~x674 & ~x699 & ~x700 & ~x702 & ~x758 & ~x763 & ~x765 & ~x779;
assign c670 = ~x3 & ~x407 & ~x446 & ~x513;
assign c672 =  x40 &  x76 &  x237 &  x403 &  x576 &  x623 & ~x2 & ~x193 & ~x198 & ~x221 & ~x222 & ~x255 & ~x281 & ~x334 & ~x362 & ~x394 & ~x421 & ~x559 & ~x756 & ~x762 & ~x782;
assign c674 =  x177 &  x203 &  x210 &  x247 &  x260 &  x314 &  x352 & ~x24 & ~x25 & ~x27 & ~x83 & ~x138 & ~x140 & ~x166 & ~x196 & ~x448 & ~x476 & ~x756 & ~x760 & ~x762 & ~x763;
assign c676 =  x41 & ~x1 & ~x2 & ~x7 & ~x11 & ~x22 & ~x26 & ~x31 & ~x36 & ~x38 & ~x51 & ~x53 & ~x57 & ~x58 & ~x81 & ~x85 & ~x108 & ~x109 & ~x111 & ~x114 & ~x164 & ~x169 & ~x173 & ~x193 & ~x200 & ~x224 & ~x225 & ~x227 & ~x249 & ~x254 & ~x280 & ~x305 & ~x334 & ~x389 & ~x390 & ~x418 & ~x420 & ~x421 & ~x423 & ~x446 & ~x476 & ~x477 & ~x502 & ~x532 & ~x533 & ~x560 & ~x561 & ~x587 & ~x764 & ~x767 & ~x768 & ~x771 & ~x773 & ~x776;
assign c678 = ~x3 & ~x16 & ~x27 & ~x52 & ~x58 & ~x109 & ~x170 & ~x192 & ~x210 & ~x331 & ~x332 & ~x338 & ~x363 & ~x448 & ~x474 & ~x505 & ~x532 & ~x586;
assign c680 =  x706 &  x741 & ~x112 & ~x196 & ~x197 & ~x621 & ~x676 & ~x724 & ~x730;
assign c682 =  x67 &  x71 &  x96 &  x125 &  x129 &  x131 &  x157 &  x182 &  x185 &  x205 &  x233 &  x235 &  x513 &  x543 &  x607 &  x624 &  x627 &  x663 &  x712 &  x714 & ~x6 & ~x7 & ~x21 & ~x107 & ~x140 & ~x142 & ~x279 & ~x308 & ~x334 & ~x338 & ~x339 & ~x394 & ~x417 & ~x448 & ~x503 & ~x531 & ~x533 & ~x735 & ~x758 & ~x764;
assign c684 =  x14 &  x73 &  x92 &  x103 &  x126 &  x242 &  x298 &  x319 &  x325 &  x382 &  x401 &  x518 &  x572 &  x575 &  x625 &  x656 &  x657 &  x683 &  x714 & ~x0 & ~x9 & ~x29 & ~x31 & ~x55 & ~x80 & ~x107 & ~x135 & ~x143 & ~x193 & ~x197 & ~x199 & ~x249 & ~x254 & ~x307 & ~x308 & ~x339 & ~x363 & ~x393 & ~x422 & ~x501 & ~x531 & ~x562 & ~x587 & ~x618 & ~x726 & ~x727 & ~x781;
assign c686 =  x87;
assign c690 =  x272 &  x462 &  x550 &  x552 &  x679 &  x684 &  x707 &  x742 &  x743 & ~x393 & ~x532 & ~x563 & ~x583 & ~x587 & ~x639 & ~x699 & ~x752;
assign c692 = ~x5 & ~x6 & ~x16 & ~x20 & ~x25 & ~x27 & ~x28 & ~x33 & ~x51 & ~x52 & ~x53 & ~x55 & ~x57 & ~x60 & ~x81 & ~x111 & ~x112 & ~x113 & ~x139 & ~x140 & ~x143 & ~x165 & ~x170 & ~x197 & ~x198 & ~x221 & ~x224 & ~x252 & ~x334 & ~x365 & ~x419 & ~x430 & ~x449 & ~x474 & ~x476 & ~x478 & ~x503 & ~x505 & ~x531 & ~x588 & ~x589 & ~x643 & ~x644 & ~x645 & ~x669 & ~x671 & ~x701 & ~x702 & ~x726 & ~x727 & ~x728 & ~x729 & ~x730 & ~x758 & ~x759 & ~x778 & ~x780 & ~x781;
assign c694 =  x754;
assign c696 =  x13 &  x15 &  x65 &  x94 &  x104 &  x120 &  x409 &  x635 &  x657 & ~x4 & ~x18 & ~x21 & ~x136 & ~x170 & ~x449 & ~x532 & ~x534 & ~x561 & ~x586 & ~x644 & ~x729 & ~x776;
assign c698 =  x186 &  x214 &  x269 &  x270 &  x318 &  x320 &  x326 &  x327 &  x344 &  x345 &  x348 &  x435 &  x436 &  x455 &  x456 &  x467 &  x485 &  x487 &  x491 &  x495 &  x514 &  x516 &  x524 &  x541 &  x576 &  x596 &  x628 &  x661 & ~x0 & ~x13 & ~x55 & ~x111 & ~x420 & ~x476 & ~x647 & ~x697 & ~x725 & ~x758 & ~x760;
assign c6100 =  x63 &  x90 &  x203 &  x371 &  x399 &  x470 &  x564 &  x566 & ~x1 & ~x6 & ~x21 & ~x22 & ~x60 & ~x79 & ~x81 & ~x109 & ~x196 & ~x251 & ~x278 & ~x280 & ~x335 & ~x420 & ~x560 & ~x615 & ~x763;
assign c6102 =  x119 &  x124 &  x302 &  x689 & ~x17 & ~x38 & ~x53 & ~x79 & ~x81 & ~x109 & ~x163 & ~x167 & ~x306 & ~x391 & ~x474 & ~x476 & ~x477 & ~x504;
assign c6104 =  x88 & ~x40;
assign c6106 = ~x28 & ~x32 & ~x35 & ~x37 & ~x38 & ~x49 & ~x51 & ~x53 & ~x79 & ~x85 & ~x107 & ~x109 & ~x139 & ~x142 & ~x200 & ~x222 & ~x225 & ~x226 & ~x252 & ~x255 & ~x282 & ~x305 & ~x308 & ~x333 & ~x335 & ~x389 & ~x395 & ~x445 & ~x449 & ~x451 & ~x478 & ~x529 & ~x532 & ~x557 & ~x560 & ~x561 & ~x613 & ~x675 & ~x697 & ~x698 & ~x725 & ~x728 & ~x737 & ~x756 & ~x765 & ~x766 & ~x771;
assign c6108 =  x92 &  x119 &  x175 &  x203 &  x245 &  x272 &  x432 &  x487 &  x539 &  x573 &  x734 & ~x22 & ~x23 & ~x28 & ~x30 & ~x168 & ~x335 & ~x477 & ~x589 & ~x617 & ~x779;
assign c6110 = ~x46 & ~x214 & ~x264;
assign c6112 =  x747 &  x771 & ~x4 & ~x24 & ~x88 & ~x112 & ~x136 & ~x141 & ~x168 & ~x170 & ~x172 & ~x197 & ~x220 & ~x221 & ~x222 & ~x225 & ~x226 & ~x247 & ~x250 & ~x254 & ~x280 & ~x304 & ~x310 & ~x332 & ~x333 & ~x335 & ~x339 & ~x362 & ~x367 & ~x387 & ~x390 & ~x391 & ~x425 & ~x426 & ~x442 & ~x449 & ~x450 & ~x452 & ~x454 & ~x475 & ~x480 & ~x502 & ~x537 & ~x557 & ~x564 & ~x588 & ~x589 & ~x590 & ~x593 & ~x611 & ~x613 & ~x614 & ~x643 & ~x644 & ~x648 & ~x698 & ~x704 & ~x726 & ~x729 & ~x753 & ~x755 & ~x756 & ~x757 & ~x758 & ~x759;
assign c6114 =  x299 &  x495 &  x546 &  x574 &  x652 &  x658 &  x719 & ~x252 & ~x256 & ~x359 & ~x365 & ~x451 & ~x557 & ~x562 & ~x610 & ~x674 & ~x697 & ~x728;
assign c6116 =  x69 & ~x0 & ~x2 & ~x3 & ~x4 & ~x5 & ~x18 & ~x20 & ~x23 & ~x28 & ~x30 & ~x34 & ~x36 & ~x45 & ~x47 & ~x48 & ~x50 & ~x54 & ~x55 & ~x58 & ~x59 & ~x60 & ~x61 & ~x76 & ~x77 & ~x78 & ~x79 & ~x80 & ~x84 & ~x86 & ~x87 & ~x88 & ~x89 & ~x90 & ~x108 & ~x109 & ~x113 & ~x135 & ~x136 & ~x137 & ~x144 & ~x163 & ~x164 & ~x168 & ~x171 & ~x196 & ~x199 & ~x222 & ~x224 & ~x227 & ~x250 & ~x251 & ~x253 & ~x281 & ~x305 & ~x306 & ~x307 & ~x333 & ~x337 & ~x362 & ~x365 & ~x366 & ~x367 & ~x390 & ~x391 & ~x392 & ~x416 & ~x417 & ~x421 & ~x445 & ~x448 & ~x449 & ~x450 & ~x474 & ~x475 & ~x476 & ~x477 & ~x504 & ~x506 & ~x528 & ~x529 & ~x530 & ~x531 & ~x532 & ~x533 & ~x534 & ~x535 & ~x558 & ~x559 & ~x560 & ~x563 & ~x590 & ~x613 & ~x614 & ~x617 & ~x619 & ~x642 & ~x645 & ~x670 & ~x671 & ~x672 & ~x674 & ~x675 & ~x697 & ~x698 & ~x699 & ~x700 & ~x701 & ~x725 & ~x726 & ~x753 & ~x755 & ~x756 & ~x763 & ~x780 & ~x781;
assign c6118 =  x506;
assign c6120 =  x326 &  x439 &  x545 &  x578 & ~x2 & ~x54 & ~x81 & ~x82 & ~x138 & ~x140 & ~x169 & ~x171 & ~x172 & ~x193 & ~x395 & ~x426 & ~x443 & ~x447 & ~x448 & ~x555 & ~x562 & ~x584 & ~x585 & ~x611 & ~x697 & ~x759 & ~x777;
assign c6122 =  x137;
assign c6124 = ~x11 & ~x45 & ~x353 & ~x673;
assign c6126 =  x92 &  x122 &  x186 &  x269 &  x346 &  x349 &  x350 &  x375 &  x435 & ~x2 & ~x19 & ~x33 & ~x52 & ~x56 & ~x89 & ~x107 & ~x144 & ~x166 & ~x168 & ~x194 & ~x195 & ~x198 & ~x221 & ~x222 & ~x229 & ~x253 & ~x308 & ~x365 & ~x366 & ~x391 & ~x534 & ~x700;
assign c6128 =  x212 &  x383 &  x409 &  x428 &  x524 &  x602 &  x651 &  x690 &  x742 & ~x13 & ~x15 & ~x27 & ~x32 & ~x52 & ~x672 & ~x701;
assign c6130 =  x158 &  x262 &  x270 &  x271 &  x458 &  x459 &  x465 &  x599 &  x719 & ~x111 & ~x195 & ~x199 & ~x366 & ~x387 & ~x396 & ~x413 & ~x471 & ~x507 & ~x610 & ~x648 & ~x702 & ~x725 & ~x730 & ~x753;
assign c6132 =  x33;
assign c6134 =  x300 &  x742 & ~x2 & ~x24 & ~x59 & ~x86 & ~x139 & ~x141 & ~x167 & ~x220 & ~x221 & ~x222 & ~x225 & ~x252 & ~x278 & ~x337 & ~x338 & ~x363 & ~x365 & ~x366 & ~x478 & ~x562 & ~x587 & ~x699 & ~x728 & ~x735 & ~x758 & ~x763 & ~x766 & ~x775 & ~x776 & ~x777 & ~x782;
assign c6136 =  x36 &  x121 &  x182 &  x232 &  x234 &  x245 &  x246 &  x247 &  x263 &  x267 &  x290 &  x319 &  x429 &  x439 &  x513 &  x540 &  x552 &  x580 &  x600 &  x657 & ~x59 & ~x81 & ~x110 & ~x254 & ~x280 & ~x392;
assign c6138 = ~x131 & ~x169 & ~x214 & ~x304 & ~x319 & ~x466;
assign c6140 =  x15 &  x43 &  x73 &  x92 &  x98 &  x266 &  x712 & ~x1 & ~x10 & ~x19 & ~x21 & ~x46 & ~x51 & ~x85 & ~x106 & ~x108 & ~x113 & ~x136 & ~x138 & ~x142 & ~x144 & ~x169 & ~x170 & ~x193 & ~x390 & ~x393 & ~x421 & ~x423 & ~x445 & ~x446 & ~x447 & ~x475 & ~x476 & ~x478 & ~x558 & ~x561 & ~x562 & ~x614 & ~x615 & ~x641 & ~x697 & ~x698 & ~x727 & ~x729 & ~x757;
assign c6142 =  x63 &  x152 &  x180 &  x231 &  x286 &  x315 &  x345 &  x376 &  x513 &  x597 &  x624 &  x651 & ~x13 & ~x55 & ~x56 & ~x83 & ~x475 & ~x560 & ~x672;
assign c6144 =  x258 & ~x4 & ~x23 & ~x28 & ~x31 & ~x40 & ~x52 & ~x53 & ~x54 & ~x81 & ~x84 & ~x140 & ~x141 & ~x169 & ~x195 & ~x197 & ~x281 & ~x306 & ~x334 & ~x475 & ~x700 & ~x758 & ~x762 & ~x783;
assign c6146 = ~x158 & ~x235 & ~x505;
assign c6148 =  x132 &  x435 &  x624 & ~x6 & ~x47 & ~x111 & ~x112 & ~x140 & ~x162 & ~x167 & ~x190 & ~x361 & ~x392 & ~x444 & ~x447 & ~x451 & ~x532 & ~x588 & ~x590 & ~x618 & ~x670 & ~x726 & ~x727;
assign c6150 =  x231 & ~x18 & ~x22 & ~x26 & ~x28 & ~x44 & ~x55 & ~x84 & ~x140 & ~x142 & ~x193 & ~x196 & ~x224 & ~x250 & ~x251 & ~x252 & ~x278 & ~x306 & ~x336 & ~x363 & ~x391 & ~x392 & ~x616 & ~x644 & ~x671 & ~x672 & ~x756 & ~x757;
assign c6152 =  x65 &  x406 & ~x58 & ~x144 & ~x220 & ~x258 & ~x310 & ~x476 & ~x509 & ~x564 & ~x587 & ~x695 & ~x724;
assign c6154 =  x92 &  x123 &  x176 &  x242 &  x413 &  x442 &  x545 &  x688 & ~x10 & ~x17 & ~x28 & ~x47 & ~x111 & ~x140 & ~x311 & ~x335 & ~x393 & ~x449 & ~x475 & ~x476 & ~x478 & ~x729 & ~x783;
assign c6156 =  x133 &  x203 &  x232 &  x272 &  x429 &  x466 & ~x0 & ~x52 & ~x109 & ~x170 & ~x197 & ~x223 & ~x309 & ~x733 & ~x758 & ~x776;
assign c6158 =  x301 &  x636 &  x665 &  x693 & ~x4 & ~x5 & ~x27 & ~x28 & ~x53 & ~x57 & ~x81 & ~x86 & ~x167 & ~x169 & ~x170 & ~x194 & ~x196 & ~x336 & ~x363 & ~x394 & ~x419 & ~x449 & ~x476 & ~x503 & ~x504 & ~x531 & ~x727 & ~x762 & ~x765 & ~x772;
assign c6160 =  x156 &  x205 &  x411 &  x546 & ~x20 & ~x22 & ~x50 & ~x228 & ~x256 & ~x339 & ~x426 & ~x560 & ~x724 & ~x731 & ~x756;
assign c6162 =  x70 & ~x2 & ~x4 & ~x5 & ~x7 & ~x10 & ~x20 & ~x24 & ~x25 & ~x30 & ~x32 & ~x37 & ~x46 & ~x49 & ~x50 & ~x54 & ~x55 & ~x61 & ~x77 & ~x83 & ~x84 & ~x85 & ~x89 & ~x107 & ~x109 & ~x115 & ~x140 & ~x144 & ~x170 & ~x171 & ~x172 & ~x193 & ~x195 & ~x197 & ~x199 & ~x220 & ~x221 & ~x222 & ~x224 & ~x227 & ~x250 & ~x333 & ~x337 & ~x338 & ~x365 & ~x391 & ~x395 & ~x446 & ~x447 & ~x473 & ~x474 & ~x476 & ~x477 & ~x478 & ~x496 & ~x532 & ~x557 & ~x558 & ~x559 & ~x560 & ~x613 & ~x614 & ~x615 & ~x616 & ~x617 & ~x641 & ~x643 & ~x644 & ~x645 & ~x646 & ~x727 & ~x755 & ~x759 & ~x764;
assign c6164 =  x104 &  x185 &  x292 &  x320 &  x355 &  x456 &  x468 &  x713 &  x769 & ~x415 & ~x564;
assign c6166 =  x60;
assign c6168 = ~x295 & ~x383 & ~x776 & ~x778;
assign c6170 =  x282;
assign c6172 =  x59;
assign c6174 =  x369 &  x585 & ~x250 & ~x765;
assign c6176 = ~x3 & ~x11 & ~x21 & ~x83 & ~x88 & ~x110 & ~x112 & ~x136 & ~x166 & ~x197 & ~x236 & ~x390 & ~x450 & ~x477 & ~x506 & ~x557 & ~x587 & ~x590 & ~x641 & ~x671;
assign c6178 =  x33;
assign c6180 =  x585;
assign c6182 =  x48 &  x232 &  x457 &  x519 &  x580 &  x742 & ~x0 & ~x54 & ~x55 & ~x647 & ~x732 & ~x754 & ~x755 & ~x782;
assign c6184 = ~x4 & ~x20 & ~x30 & ~x57 & ~x58 & ~x88 & ~x111 & ~x114 & ~x136 & ~x449 & ~x474 & ~x479 & ~x502 & ~x507 & ~x528 & ~x562 & ~x615 & ~x643 & ~x648 & ~x656 & ~x674 & ~x699 & ~x704 & ~x728 & ~x758 & ~x777 & ~x778 & ~x783;
assign c6186 =  x101 &  x128 &  x158 &  x184 &  x270 &  x294 &  x317 &  x460 &  x496 &  x568 &  x569 &  x576 & ~x13 & ~x29 & ~x31 & ~x82 & ~x112 & ~x137 & ~x167 & ~x195 & ~x221 & ~x222 & ~x250 & ~x254 & ~x304 & ~x312 & ~x335 & ~x365 & ~x392 & ~x475;
assign c6188 =  x288 &  x712 & ~x7 & ~x28 & ~x32 & ~x46 & ~x49 & ~x54 & ~x55 & ~x76 & ~x88 & ~x89 & ~x115 & ~x141 & ~x169 & ~x196 & ~x223 & ~x225 & ~x226 & ~x307 & ~x309 & ~x361 & ~x364 & ~x530 & ~x532 & ~x558 & ~x588 & ~x613 & ~x673 & ~x776;
assign c6190 =  x609 & ~x646 & ~x647 & ~x701;
assign c6192 = ~x0 & ~x11 & ~x53 & ~x86 & ~x140 & ~x227 & ~x249 & ~x252 & ~x267 & ~x333 & ~x446 & ~x683 & ~x756 & ~x783;
assign c6194 =  x143;
assign c6196 =  x90 &  x612 & ~x171 & ~x308;
assign c6198 =  x200 &  x246 &  x287 &  x301 &  x408 &  x523 & ~x563 & ~x589 & ~x616 & ~x668 & ~x697 & ~x731 & ~x752;
assign c6200 =  x582 & ~x23 & ~x28 & ~x29 & ~x82 & ~x84 & ~x86 & ~x140 & ~x142 & ~x193 & ~x196 & ~x222 & ~x223 & ~x224 & ~x279 & ~x306 & ~x308 & ~x334 & ~x362 & ~x364 & ~x390 & ~x419 & ~x421 & ~x503 & ~x756 & ~x762;
assign c6202 =  x68 &  x96 &  x186 &  x209 &  x266 &  x326 &  x576 & ~x1 & ~x2 & ~x25 & ~x30 & ~x56 & ~x57 & ~x59 & ~x86 & ~x107 & ~x110 & ~x112 & ~x134 & ~x135 & ~x137 & ~x144 & ~x145 & ~x164 & ~x166 & ~x169 & ~x170 & ~x191 & ~x195 & ~x198 & ~x199 & ~x220 & ~x222 & ~x225 & ~x227 & ~x278 & ~x281 & ~x306 & ~x309 & ~x311 & ~x360 & ~x395 & ~x421 & ~x446 & ~x474 & ~x530 & ~x589 & ~x646 & ~x699 & ~x726 & ~x754 & ~x759 & ~x760 & ~x779;
assign c6204 =  x289 &  x401 &  x439 & ~x32 & ~x33 & ~x110 & ~x191 & ~x331 & ~x359 & ~x525 & ~x750;
assign c6206 =  x62 &  x188 &  x231 &  x236 &  x239 &  x376 &  x404 &  x456 &  x458 &  x462 &  x665 & ~x196 & ~x391 & ~x616 & ~x783;
assign c6208 =  x40 &  x43 &  x71 &  x133 &  x230 &  x231 &  x300 &  x328 &  x574 &  x607 &  x652 & ~x1 & ~x19 & ~x23 & ~x33 & ~x55 & ~x58 & ~x111 & ~x139 & ~x166 & ~x170 & ~x171 & ~x191 & ~x192 & ~x193 & ~x224 & ~x251 & ~x389 & ~x391 & ~x392 & ~x419 & ~x449 & ~x502 & ~x560 & ~x669 & ~x674 & ~x697 & ~x726 & ~x728 & ~x776;
assign c6210 =  x231 &  x357 &  x440 &  x491 &  x526 & ~x15 & ~x21 & ~x26 & ~x28 & ~x53 & ~x87 & ~x109 & ~x116 & ~x136 & ~x169 & ~x221 & ~x222 & ~x224 & ~x251 & ~x419 & ~x476 & ~x755 & ~x782;
assign c6212 =  x256 & ~x564 & ~x776 & ~x780;
assign c6214 =  x103 &  x131 &  x148 &  x158 &  x177 &  x208 &  x269 &  x272 &  x292 &  x326 &  x352 &  x384 &  x494 &  x495 &  x574 &  x627 &  x635 &  x655 &  x657 &  x694 & ~x5 & ~x54 & ~x81 & ~x138 & ~x167 & ~x193 & ~x194 & ~x219 & ~x309 & ~x332 & ~x367 & ~x589 & ~x672 & ~x728 & ~x756;
assign c6216 =  x69 & ~x10 & ~x19 & ~x21 & ~x36 & ~x45 & ~x47 & ~x51 & ~x53 & ~x63 & ~x79 & ~x83 & ~x84 & ~x85 & ~x88 & ~x111 & ~x117 & ~x139 & ~x143 & ~x166 & ~x171 & ~x192 & ~x252 & ~x254 & ~x307 & ~x311 & ~x339 & ~x389 & ~x420 & ~x421 & ~x423 & ~x444 & ~x448 & ~x474 & ~x475 & ~x534 & ~x563 & ~x587 & ~x642 & ~x672 & ~x701 & ~x756 & ~x759 & ~x764 & ~x775 & ~x783;
assign c6218 =  x289 &  x299 &  x460 & ~x172 & ~x539;
assign c6220 =  x92 &  x215 &  x326 &  x513 &  x572 &  x631 & ~x2 & ~x25 & ~x36 & ~x47 & ~x51 & ~x52 & ~x58 & ~x60 & ~x81 & ~x106 & ~x111 & ~x136 & ~x144 & ~x165 & ~x170 & ~x195 & ~x196 & ~x223 & ~x252 & ~x280 & ~x312 & ~x420 & ~x444 & ~x448 & ~x531 & ~x558 & ~x560 & ~x562 & ~x585 & ~x590 & ~x671 & ~x755 & ~x781;
assign c6222 =  x285 & ~x3 & ~x16 & ~x22 & ~x25 & ~x27 & ~x28 & ~x29 & ~x31 & ~x44 & ~x82 & ~x83 & ~x111 & ~x167 & ~x168 & ~x194 & ~x223 & ~x252 & ~x279 & ~x308 & ~x336 & ~x364 & ~x392 & ~x419 & ~x476 & ~x756 & ~x763;
assign c6224 =  x231 &  x397 &  x442 &  x480 &  x487 &  x526 & ~x1 & ~x6 & ~x14 & ~x25 & ~x29 & ~x51 & ~x56 & ~x57 & ~x58 & ~x82 & ~x108 & ~x110 & ~x114 & ~x137 & ~x141 & ~x143 & ~x193 & ~x196 & ~x225 & ~x251 & ~x279 & ~x281 & ~x335 & ~x336 & ~x337 & ~x392 & ~x758 & ~x780;
assign c6226 =  x118 &  x328 &  x743 & ~x2 & ~x3 & ~x6 & ~x8 & ~x26 & ~x30 & ~x54 & ~x55 & ~x56 & ~x57 & ~x59 & ~x60 & ~x87 & ~x109 & ~x111 & ~x113 & ~x115 & ~x116 & ~x136 & ~x137 & ~x138 & ~x139 & ~x143 & ~x165 & ~x167 & ~x194 & ~x250 & ~x251 & ~x252 & ~x308 & ~x336 & ~x362 & ~x366 & ~x393 & ~x420 & ~x446 & ~x449 & ~x477 & ~x503 & ~x505 & ~x587 & ~x671 & ~x702 & ~x726 & ~x728 & ~x729 & ~x756 & ~x758 & ~x783;
assign c6228 =  x59;
assign c6230 =  x213 &  x667 &  x752 & ~x136 & ~x141 & ~x759 & ~x763;
assign c6232 =  x137;
assign c6234 =  x119 &  x300 & ~x3 & ~x5 & ~x9 & ~x18 & ~x25 & ~x33 & ~x45 & ~x50 & ~x62 & ~x83 & ~x85 & ~x111 & ~x138 & ~x143 & ~x144 & ~x166 & ~x167 & ~x224 & ~x280 & ~x281 & ~x307 & ~x309 & ~x419 & ~x502 & ~x503 & ~x504 & ~x530 & ~x560 & ~x561 & ~x588 & ~x643 & ~x644 & ~x700 & ~x729 & ~x757 & ~x780;
assign c6236 =  x568 & ~x280 & ~x371 & ~x385 & ~x446 & ~x449 & ~x453 & ~x480 & ~x560 & ~x586 & ~x588 & ~x615 & ~x618 & ~x730 & ~x733 & ~x734 & ~x751 & ~x761 & ~x763;
assign c6238 = ~x3 & ~x25 & ~x28 & ~x32 & ~x58 & ~x76 & ~x84 & ~x86 & ~x87 & ~x88 & ~x110 & ~x111 & ~x137 & ~x141 & ~x168 & ~x193 & ~x197 & ~x224 & ~x250 & ~x251 & ~x254 & ~x269 & ~x280 & ~x306 & ~x307 & ~x309 & ~x334 & ~x336 & ~x337 & ~x338 & ~x362 & ~x363 & ~x391 & ~x392 & ~x418 & ~x422 & ~x474 & ~x475 & ~x502 & ~x514 & ~x560 & ~x587 & ~x615 & ~x700 & ~x701 & ~x759;
assign c6240 =  x36 &  x235 &  x412 &  x517 & ~x20 & ~x21 & ~x27 & ~x252 & ~x276 & ~x644;
assign c6242 =  x68 &  x73 &  x92 &  x101 &  x128 &  x129 &  x131 &  x156 &  x159 &  x178 &  x183 &  x209 &  x232 &  x236 &  x239 &  x267 &  x270 &  x289 &  x290 &  x297 &  x320 &  x323 &  x345 &  x373 &  x401 &  x435 &  x436 &  x457 &  x624 &  x630 &  x655 & ~x4 & ~x9 & ~x19 & ~x27 & ~x29 & ~x57 & ~x60 & ~x61 & ~x82 & ~x110 & ~x113 & ~x136 & ~x137 & ~x163 & ~x164 & ~x199 & ~x200 & ~x221 & ~x225 & ~x228 & ~x249 & ~x282 & ~x284 & ~x332 & ~x333 & ~x339 & ~x363 & ~x392 & ~x448 & ~x558 & ~x589 & ~x645 & ~x670;
assign c6244 =  x133 &  x202 &  x210 &  x407 &  x549 &  x718 & ~x25 & ~x222 & ~x727 & ~x736 & ~x765;
assign c6246 =  x60;
assign c6248 =  x203 &  x385 &  x413 &  x469 &  x472 & ~x0 & ~x2 & ~x21 & ~x22 & ~x24 & ~x25 & ~x55 & ~x81 & ~x108 & ~x109 & ~x110 & ~x138 & ~x170 & ~x171 & ~x194 & ~x195 & ~x198 & ~x221 & ~x223 & ~x224 & ~x226 & ~x252 & ~x254 & ~x280 & ~x306 & ~x310 & ~x335 & ~x338 & ~x362 & ~x364 & ~x391 & ~x447 & ~x503 & ~x644 & ~x671 & ~x673 & ~x763;
assign c6250 =  x103 &  x713 & ~x1 & ~x6 & ~x25 & ~x30 & ~x32 & ~x37 & ~x47 & ~x48 & ~x52 & ~x54 & ~x56 & ~x57 & ~x58 & ~x84 & ~x106 & ~x110 & ~x167 & ~x226 & ~x363 & ~x419 & ~x422 & ~x447 & ~x451 & ~x476 & ~x478 & ~x504 & ~x529 & ~x560 & ~x562 & ~x585 & ~x586 & ~x587 & ~x618 & ~x645 & ~x701 & ~x729 & ~x763 & ~x775;
assign c6252 =  x47 &  x185 &  x290 &  x295 &  x318 &  x373 &  x408 &  x430 &  x431 &  x522 &  x604 & ~x164 & ~x307 & ~x556 & ~x582 & ~x645 & ~x728;
assign c6254 =  x60;
assign c6256 =  x203 &  x484 & ~x0 & ~x2 & ~x3 & ~x6 & ~x14 & ~x15 & ~x21 & ~x24 & ~x28 & ~x30 & ~x51 & ~x53 & ~x55 & ~x57 & ~x82 & ~x84 & ~x85 & ~x87 & ~x108 & ~x109 & ~x110 & ~x112 & ~x113 & ~x114 & ~x137 & ~x138 & ~x142 & ~x143 & ~x165 & ~x166 & ~x167 & ~x169 & ~x170 & ~x196 & ~x197 & ~x221 & ~x222 & ~x223 & ~x225 & ~x226 & ~x250 & ~x251 & ~x279 & ~x281 & ~x391 & ~x422 & ~x447 & ~x449 & ~x474 & ~x476 & ~x477 & ~x478 & ~x502 & ~x531 & ~x559 & ~x586 & ~x588 & ~x589 & ~x616 & ~x617 & ~x645 & ~x646 & ~x670 & ~x672 & ~x673 & ~x698 & ~x699 & ~x700 & ~x728 & ~x731 & ~x751 & ~x752 & ~x755 & ~x757 & ~x761 & ~x778 & ~x779 & ~x782;
assign c6258 =  x46 &  x76 &  x204 &  x206 &  x261 &  x268 &  x270 &  x292 &  x295 &  x326 &  x434 &  x435 &  x457 &  x464 &  x466 &  x467 &  x516 &  x540 &  x549 &  x575 &  x605 & ~x27 & ~x29 & ~x87 & ~x107 & ~x165 & ~x166 & ~x170 & ~x363 & ~x393 & ~x558 & ~x560 & ~x562 & ~x672 & ~x697 & ~x783;
assign c6260 =  x326 &  x353 &  x436 &  x490 &  x602 & ~x29 & ~x32 & ~x49 & ~x85 & ~x191 & ~x225 & ~x279 & ~x335 & ~x360 & ~x417 & ~x526 & ~x528 & ~x558 & ~x610 & ~x613 & ~x672 & ~x676 & ~x698 & ~x700 & ~x724 & ~x730 & ~x782 & ~x783;
assign c6262 =  x41 &  x103 &  x681 & ~x2 & ~x4 & ~x21 & ~x25 & ~x34 & ~x37 & ~x46 & ~x47 & ~x59 & ~x61 & ~x77 & ~x83 & ~x106 & ~x108 & ~x111 & ~x136 & ~x167 & ~x279 & ~x362 & ~x391 & ~x393 & ~x474 & ~x475 & ~x529 & ~x531 & ~x559 & ~x618 & ~x643 & ~x671 & ~x674 & ~x754 & ~x755 & ~x765;
assign c6264 =  x203 &  x295 &  x322 &  x548 &  x666 &  x738 & ~x1 & ~x22 & ~x29 & ~x51 & ~x53 & ~x56 & ~x80 & ~x81 & ~x85 & ~x195 & ~x197 & ~x307 & ~x447 & ~x449 & ~x505 & ~x529 & ~x587 & ~x590 & ~x615 & ~x617;
assign c6266 =  x275 &  x385 & ~x57 & ~x109 & ~x668 & ~x698 & ~x701 & ~x728 & ~x732 & ~x759 & ~x779;
assign c6268 =  x266 &  x317 &  x349 &  x401 &  x432 &  x461 &  x545 & ~x32 & ~x52 & ~x53 & ~x138 & ~x139 & ~x140 & ~x170 & ~x192 & ~x196 & ~x220 & ~x221 & ~x222 & ~x250 & ~x280 & ~x281 & ~x283 & ~x303 & ~x308 & ~x309 & ~x333 & ~x342 & ~x358 & ~x367 & ~x394 & ~x414 & ~x421 & ~x453 & ~x469 & ~x475 & ~x477 & ~x531 & ~x536 & ~x556 & ~x564 & ~x585 & ~x588 & ~x639 & ~x729 & ~x732;
assign c6270 =  x273 &  x744 & ~x4 & ~x6 & ~x29 & ~x38 & ~x54 & ~x63 & ~x81 & ~x84 & ~x87 & ~x136 & ~x139 & ~x165 & ~x199 & ~x254 & ~x279 & ~x335 & ~x418 & ~x560 & ~x561 & ~x615 & ~x730 & ~x764 & ~x782;
assign c6272 =  x394;
assign c6274 =  x161 &  x267 &  x295 &  x371 &  x623 &  x658 & ~x82 & ~x83 & ~x335 & ~x475 & ~x736 & ~x748 & ~x756 & ~x774;
assign c6276 =  x35 &  x299 &  x301 &  x372 &  x408 &  x430 &  x468 &  x491 & ~x167 & ~x195;
assign c6278 =  x64 &  x148 &  x301 &  x353 &  x374 &  x538 &  x548 &  x608 &  x609 &  x611 & ~x80 & ~x113 & ~x227 & ~x366 & ~x447 & ~x478 & ~x589;
assign c6280 =  x64 &  x526 &  x612 &  x640 & ~x5 & ~x24 & ~x53 & ~x80 & ~x110 & ~x116 & ~x141 & ~x223 & ~x227 & ~x254 & ~x309 & ~x756;
assign c6282 =  x569 &  x742 & ~x22 & ~x30 & ~x278 & ~x421 & ~x422 & ~x530 & ~x587 & ~x736 & ~x748 & ~x756 & ~x764;
assign c6284 =  x359 &  x368 &  x480 & ~x11 & ~x14 & ~x197 & ~x277 & ~x278 & ~x309 & ~x336 & ~x756;
assign c6286 =  x93 &  x101 &  x401 &  x709 & ~x9 & ~x38 & ~x46 & ~x49 & ~x83 & ~x109 & ~x198 & ~x474 & ~x504 & ~x559 & ~x727 & ~x763;
assign c6288 =  x189 &  x216 & ~x5 & ~x19 & ~x21 & ~x23 & ~x32 & ~x33 & ~x58 & ~x59 & ~x83 & ~x107 & ~x110 & ~x111 & ~x163 & ~x165 & ~x166 & ~x167 & ~x168 & ~x170 & ~x171 & ~x193 & ~x194 & ~x199 & ~x220 & ~x225 & ~x249 & ~x253 & ~x309 & ~x335 & ~x338 & ~x392 & ~x395 & ~x417 & ~x422 & ~x446 & ~x504 & ~x531 & ~x532 & ~x559 & ~x561 & ~x587 & ~x588 & ~x618 & ~x674 & ~x701 & ~x749 & ~x764 & ~x777 & ~x782;
assign c6290 =  x64 &  x751 &  x752 & ~x446;
assign c6292 =  x563 & ~x22 & ~x139 & ~x140 & ~x142 & ~x195 & ~x198 & ~x221 & ~x418 & ~x760;
assign c6294 =  x282;
assign c6296 =  x92 &  x120 &  x237 &  x266 &  x299 &  x301 &  x350 &  x372 &  x401 &  x408 &  x520 &  x577 &  x609 &  x713 & ~x11 & ~x24 & ~x168 & ~x588 & ~x763;
assign c6298 =  x14 &  x91 &  x174 &  x300 &  x742 & ~x7 & ~x9 & ~x29 & ~x84 & ~x116 & ~x394 & ~x421 & ~x559 & ~x587 & ~x588 & ~x589 & ~x764 & ~x765;
assign c6300 =  x33;
assign c6302 =  x158 &  x326 &  x327 &  x383 &  x437 &  x541 &  x681 & ~x10 & ~x46 & ~x63 & ~x79 & ~x83 & ~x86 & ~x90 & ~x115 & ~x116 & ~x446 & ~x450 & ~x506 & ~x534 & ~x563 & ~x615 & ~x647 & ~x671 & ~x781;
assign c6304 =  x242 &  x289 &  x297 &  x298 &  x318 &  x348 &  x434 &  x439 &  x465 &  x492 &  x495 &  x571 &  x596 &  x597 &  x607 & ~x58 & ~x144 & ~x196 & ~x310 & ~x447 & ~x526 & ~x582 & ~x583 & ~x588 & ~x592 & ~x647 & ~x667 & ~x672 & ~x673 & ~x675 & ~x726 & ~x732 & ~x750 & ~x778 & ~x781;
assign c6306 =  x146 &  x741 & ~x0 & ~x22 & ~x27 & ~x31 & ~x46 & ~x47 & ~x49 & ~x52 & ~x53 & ~x54 & ~x107 & ~x141 & ~x193 & ~x226 & ~x306 & ~x310 & ~x335 & ~x362 & ~x421 & ~x615 & ~x727 & ~x729;
assign c6308 =  x60;
assign c6310 =  x637 &  x724 & ~x198 & ~x225 & ~x226 & ~x308 & ~x337 & ~x363 & ~x364 & ~x449 & ~x505 & ~x756 & ~x763;
assign c6312 = ~x18 & ~x36 & ~x47 & ~x80 & ~x112 & ~x170 & ~x390 & ~x411 & ~x448 & ~x476 & ~x644 & ~x754 & ~x781;
assign c6314 =  x105 &  x203 &  x272 &  x370 &  x371 &  x415 & ~x7 & ~x25 & ~x27 & ~x57 & ~x81 & ~x167 & ~x169 & ~x171 & ~x197 & ~x200 & ~x223 & ~x226 & ~x255 & ~x276 & ~x418 & ~x475 & ~x476 & ~x588 & ~x615 & ~x616 & ~x671 & ~x782 & ~x783;
assign c6316 = ~x1 & ~x2 & ~x4 & ~x5 & ~x21 & ~x23 & ~x25 & ~x26 & ~x27 & ~x28 & ~x29 & ~x30 & ~x32 & ~x33 & ~x49 & ~x51 & ~x56 & ~x57 & ~x58 & ~x59 & ~x79 & ~x82 & ~x83 & ~x84 & ~x85 & ~x86 & ~x108 & ~x110 & ~x111 & ~x112 & ~x114 & ~x115 & ~x136 & ~x137 & ~x138 & ~x139 & ~x140 & ~x141 & ~x144 & ~x165 & ~x166 & ~x170 & ~x192 & ~x195 & ~x196 & ~x197 & ~x221 & ~x223 & ~x224 & ~x225 & ~x227 & ~x248 & ~x249 & ~x250 & ~x251 & ~x252 & ~x277 & ~x279 & ~x282 & ~x306 & ~x333 & ~x334 & ~x336 & ~x339 & ~x362 & ~x364 & ~x365 & ~x367 & ~x389 & ~x390 & ~x391 & ~x392 & ~x393 & ~x394 & ~x417 & ~x418 & ~x420 & ~x446 & ~x449 & ~x450 & ~x473 & ~x474 & ~x475 & ~x476 & ~x478 & ~x502 & ~x506 & ~x529 & ~x531 & ~x542 & ~x558 & ~x560 & ~x561 & ~x587 & ~x589 & ~x613 & ~x617 & ~x618 & ~x643 & ~x644 & ~x671 & ~x698 & ~x699 & ~x700 & ~x701 & ~x727 & ~x728 & ~x756 & ~x757 & ~x777 & ~x780 & ~x781 & ~x782;
assign c6318 =  x92 &  x691 & ~x0 & ~x4 & ~x5 & ~x6 & ~x7 & ~x8 & ~x10 & ~x19 & ~x24 & ~x27 & ~x28 & ~x30 & ~x32 & ~x37 & ~x38 & ~x46 & ~x52 & ~x53 & ~x57 & ~x58 & ~x84 & ~x87 & ~x107 & ~x165 & ~x168 & ~x170 & ~x195 & ~x197 & ~x223 & ~x249 & ~x280 & ~x365 & ~x392 & ~x420 & ~x421 & ~x422 & ~x503 & ~x558 & ~x559 & ~x586 & ~x589 & ~x614 & ~x615 & ~x618 & ~x643 & ~x644 & ~x673 & ~x727 & ~x728 & ~x781 & ~x782;
assign c6320 =  x90 &  x91 &  x205 &  x286 &  x287 &  x300 &  x319 &  x341 &  x343 &  x345 &  x369 &  x376 &  x623 &  x654 & ~x110 & ~x248 & ~x278;
assign c6322 =  x93 &  x132 &  x211 &  x328 & ~x49 & ~x145 & ~x227 & ~x228 & ~x253 & ~x336 & ~x418 & ~x478 & ~x587 & ~x755 & ~x756 & ~x774;
assign c6324 =  x202 &  x343 & ~x0 & ~x27 & ~x58 & ~x85 & ~x448 & ~x565 & ~x620 & ~x676 & ~x697 & ~x732 & ~x754;
assign c6326 =  x123 &  x462 & ~x24 & ~x34 & ~x112 & ~x171 & ~x194 & ~x222 & ~x228 & ~x280 & ~x338 & ~x426 & ~x445 & ~x454 & ~x503 & ~x582 & ~x586 & ~x614 & ~x620 & ~x638 & ~x648 & ~x698 & ~x700 & ~x703;
assign c6328 =  x272 & ~x2 & ~x17 & ~x24 & ~x25 & ~x52 & ~x53 & ~x136 & ~x139 & ~x150 & ~x164 & ~x170 & ~x194 & ~x199 & ~x223 & ~x252 & ~x279 & ~x420 & ~x450 & ~x503 & ~x505 & ~x558 & ~x588 & ~x643 & ~x671 & ~x699 & ~x726 & ~x728 & ~x783;
assign c6330 =  x219 &  x287 &  x770 & ~x2 & ~x364 & ~x615;
assign c6332 =  x400 &  x658 &  x680 &  x707 & ~x21 & ~x26 & ~x60 & ~x109 & ~x136 & ~x137 & ~x168 & ~x170 & ~x220 & ~x390 & ~x391 & ~x395 & ~x448 & ~x450 & ~x506 & ~x535 & ~x554 & ~x558 & ~x563 & ~x582 & ~x587 & ~x589 & ~x590 & ~x618 & ~x642 & ~x698 & ~x727 & ~x754 & ~x756 & ~x757 & ~x783;
assign c6334 =  x231 & ~x53 & ~x111 & ~x112 & ~x263 & ~x280 & ~x308 & ~x758;
assign c6336 =  x342 & ~x1 & ~x13 & ~x23 & ~x25 & ~x28 & ~x41 & ~x53 & ~x56 & ~x57 & ~x81 & ~x84 & ~x85 & ~x111 & ~x112 & ~x114 & ~x142 & ~x167 & ~x169 & ~x195 & ~x197 & ~x222 & ~x307 & ~x363 & ~x448 & ~x503 & ~x756 & ~x782 & ~x783;
assign c6338 =  x230 &  x395 & ~x249;
assign c6340 =  x236 &  x316 &  x623 & ~x29 & ~x54 & ~x81 & ~x165 & ~x167 & ~x192 & ~x582 & ~x639 & ~x699 & ~x757 & ~x778;
assign c6342 = ~x38 & ~x167 & ~x280 & ~x281 & ~x456 & ~x530 & ~x586 & ~x766 & ~x776;
assign c6344 =  x43 &  x146 &  x328 &  x689 & ~x7 & ~x29 & ~x51 & ~x116 & ~x166 & ~x221 & ~x248 & ~x278 & ~x281 & ~x311 & ~x477 & ~x588 & ~x700 & ~x757 & ~x764 & ~x779;
assign c6346 =  x70 & ~x0 & ~x114 & ~x144 & ~x198 & ~x252 & ~x311 & ~x333 & ~x334 & ~x436 & ~x475 & ~x586 & ~x701 & ~x781 & ~x783;
assign c6348 = ~x149 & ~x319 & ~x429 & ~x494;
assign c6350 =  x97 &  x146 &  x316 &  x743 & ~x2 & ~x8 & ~x18 & ~x47 & ~x53 & ~x56 & ~x80 & ~x81 & ~x109 & ~x168 & ~x194 & ~x196 & ~x307 & ~x308 & ~x418 & ~x419 & ~x421 & ~x474 & ~x477 & ~x672 & ~x763;
assign c6352 =  x218 & ~x4 & ~x17 & ~x37 & ~x38 & ~x139 & ~x195 & ~x251 & ~x279 & ~x365 & ~x390 & ~x392 & ~x393 & ~x418 & ~x421 & ~x446 & ~x448 & ~x476 & ~x502 & ~x558 & ~x642 & ~x727 & ~x757 & ~x765;
assign c6354 =  x205 &  x569 &  x574 & ~x24 & ~x31 & ~x136 & ~x144 & ~x145 & ~x278 & ~x749 & ~x771;
assign c6356 =  x260 &  x462 &  x495 &  x680 & ~x23 & ~x51 & ~x53 & ~x55 & ~x80 & ~x81 & ~x193 & ~x198 & ~x224 & ~x303 & ~x304 & ~x335 & ~x342 & ~x416 & ~x417 & ~x445 & ~x479 & ~x480 & ~x504 & ~x557 & ~x563 & ~x584 & ~x699 & ~x730 & ~x752 & ~x757 & ~x780;
assign c6358 =  x40 &  x69 &  x97 &  x99 &  x119 &  x583 &  x714 & ~x37 & ~x47 & ~x83 & ~x170;
assign c6360 = ~x7 & ~x8 & ~x23 & ~x24 & ~x55 & ~x81 & ~x82 & ~x107 & ~x111 & ~x112 & ~x113 & ~x136 & ~x137 & ~x140 & ~x168 & ~x193 & ~x222 & ~x393 & ~x446 & ~x447 & ~x504 & ~x539 & ~x559 & ~x645 & ~x669 & ~x670 & ~x727 & ~x775;
assign c6362 =  x350 &  x495 & ~x60 & ~x164 & ~x199 & ~x503 & ~x532 & ~x561 & ~x694 & ~x766 & ~x778;
assign c6364 = ~x3 & ~x17 & ~x20 & ~x22 & ~x29 & ~x32 & ~x52 & ~x79 & ~x86 & ~x87 & ~x108 & ~x139 & ~x152 & ~x168 & ~x196 & ~x227 & ~x251 & ~x305 & ~x306 & ~x308 & ~x333 & ~x361 & ~x367 & ~x418 & ~x421 & ~x424 & ~x449 & ~x474 & ~x478 & ~x503 & ~x529 & ~x534 & ~x613 & ~x616 & ~x618 & ~x641 & ~x674 & ~x697 & ~x699 & ~x700 & ~x726 & ~x728 & ~x754 & ~x755 & ~x759 & ~x779;
assign c6366 =  x92 &  x608 &  x609 &  x752 & ~x110 & ~x194 & ~x309;
assign c6368 =  x451 & ~x29 & ~x53 & ~x86 & ~x198 & ~x363 & ~x587 & ~x760;
assign c6370 = ~x46 & ~x178 & ~x378 & ~x586;
assign c6372 =  x42 & ~x17 & ~x29 & ~x83 & ~x116 & ~x122 & ~x221 & ~x249 & ~x474 & ~x532 & ~x756;
assign c6374 =  x37 &  x76 &  x96 &  x185 &  x207 &  x238 &  x241 &  x244 &  x260 &  x295 &  x300 &  x321 &  x353 &  x354 &  x433 &  x462 &  x572 &  x636 &  x657 & ~x3 & ~x60 & ~x79 & ~x81 & ~x86 & ~x248 & ~x282 & ~x335 & ~x394 & ~x448;
assign c6376 =  x70 & ~x1 & ~x5 & ~x6 & ~x9 & ~x10 & ~x11 & ~x17 & ~x20 & ~x23 & ~x24 & ~x27 & ~x28 & ~x32 & ~x36 & ~x38 & ~x45 & ~x48 & ~x59 & ~x60 & ~x62 & ~x63 & ~x78 & ~x80 & ~x88 & ~x109 & ~x117 & ~x136 & ~x139 & ~x141 & ~x164 & ~x168 & ~x171 & ~x197 & ~x199 & ~x223 & ~x224 & ~x252 & ~x277 & ~x278 & ~x279 & ~x305 & ~x308 & ~x309 & ~x366 & ~x368 & ~x393 & ~x420 & ~x422 & ~x445 & ~x446 & ~x447 & ~x449 & ~x500 & ~x535 & ~x558 & ~x589 & ~x591 & ~x613 & ~x618 & ~x641 & ~x642 & ~x670 & ~x673 & ~x698 & ~x725 & ~x727 & ~x729 & ~x782;
assign c6378 =  x118 &  x294 &  x300 &  x371 &  x399 &  x492 &  x499 &  x604 & ~x20 & ~x22 & ~x30 & ~x138 & ~x166 & ~x171 & ~x193 & ~x221 & ~x228 & ~x252 & ~x277 & ~x279 & ~x280 & ~x337 & ~x422 & ~x504 & ~x700;
assign c6380 =  x41 & ~x1 & ~x2 & ~x22 & ~x27 & ~x34 & ~x53 & ~x54 & ~x55 & ~x60 & ~x87 & ~x108 & ~x116 & ~x141 & ~x143 & ~x167 & ~x169 & ~x193 & ~x222 & ~x255 & ~x308 & ~x333 & ~x334 & ~x420 & ~x421 & ~x449 & ~x474 & ~x502 & ~x503 & ~x505 & ~x587 & ~x599 & ~x615 & ~x617 & ~x645 & ~x757 & ~x764 & ~x777;
assign c6382 =  x15 &  x40 &  x73 &  x98 &  x103 &  x153 &  x161 &  x176 &  x373 &  x382 &  x514 &  x548 &  x656 &  x715 &  x716 & ~x2 & ~x18 & ~x36 & ~x49 & ~x82 & ~x83 & ~x108 & ~x112 & ~x142 & ~x197 & ~x249 & ~x253 & ~x279 & ~x280 & ~x335 & ~x364 & ~x422 & ~x644;
assign c6384 = ~x1 & ~x2 & ~x10 & ~x18 & ~x21 & ~x26 & ~x27 & ~x29 & ~x44 & ~x53 & ~x54 & ~x55 & ~x56 & ~x81 & ~x83 & ~x195 & ~x224 & ~x448 & ~x449 & ~x450 & ~x500 & ~x501 & ~x502 & ~x503 & ~x505 & ~x528 & ~x529 & ~x530 & ~x557 & ~x558 & ~x562 & ~x563 & ~x587 & ~x617 & ~x619 & ~x642 & ~x671 & ~x697 & ~x699 & ~x724 & ~x728 & ~x754 & ~x757 & ~x763 & ~x779;
assign c6386 =  x61 &  x329 &  x376 &  x651 & ~x756;
assign c6388 =  x441 &  x444 & ~x1 & ~x4 & ~x57 & ~x81 & ~x84 & ~x109 & ~x223 & ~x250 & ~x253 & ~x278 & ~x306 & ~x308 & ~x310 & ~x336 & ~x391 & ~x475 & ~x761 & ~x783;
assign c6390 =  x92 &  x128 &  x401 &  x425 &  x681 & ~x21 & ~x23 & ~x31 & ~x37 & ~x47 & ~x112 & ~x138 & ~x141 & ~x168 & ~x254 & ~x278 & ~x393 & ~x394 & ~x477;
assign c6392 =  x373 & ~x14 & ~x29 & ~x30 & ~x50 & ~x51 & ~x224 & ~x281 & ~x334 & ~x335 & ~x476 & ~x709;
assign c6394 =  x68 & ~x31 & ~x33 & ~x79 & ~x85 & ~x86 & ~x115 & ~x142 & ~x152 & ~x169 & ~x197 & ~x224 & ~x252 & ~x255 & ~x278 & ~x279 & ~x334 & ~x338 & ~x421 & ~x446 & ~x474 & ~x477 & ~x478 & ~x559 & ~x560 & ~x643 & ~x700 & ~x701 & ~x728 & ~x775;
assign c6396 =  x203 & ~x4 & ~x12 & ~x15 & ~x16 & ~x26 & ~x29 & ~x42 & ~x56 & ~x59 & ~x60 & ~x82 & ~x86 & ~x87 & ~x113 & ~x142 & ~x165 & ~x195 & ~x223 & ~x251 & ~x254 & ~x279 & ~x306 & ~x308 & ~x335 & ~x391 & ~x392 & ~x589 & ~x616 & ~x617 & ~x642 & ~x644 & ~x754 & ~x756 & ~x758;
assign c6398 =  x456 &  x545 &  x692 & ~x6 & ~x193 & ~x227 & ~x313 & ~x447 & ~x449 & ~x454 & ~x508 & ~x533 & ~x752;
assign c6400 =  x383 & ~x1 & ~x2 & ~x5 & ~x27 & ~x28 & ~x29 & ~x33 & ~x54 & ~x56 & ~x57 & ~x58 & ~x59 & ~x87 & ~x110 & ~x111 & ~x112 & ~x139 & ~x144 & ~x169 & ~x193 & ~x194 & ~x197 & ~x221 & ~x310 & ~x335 & ~x336 & ~x338 & ~x361 & ~x364 & ~x386 & ~x390 & ~x391 & ~x393 & ~x448 & ~x452 & ~x453 & ~x472 & ~x473 & ~x480 & ~x481 & ~x482 & ~x501 & ~x504 & ~x528 & ~x532 & ~x534 & ~x535 & ~x556 & ~x562 & ~x566 & ~x592 & ~x611 & ~x615 & ~x671 & ~x699 & ~x702 & ~x704 & ~x705 & ~x724 & ~x725 & ~x726 & ~x728 & ~x731 & ~x732 & ~x758 & ~x760 & ~x761 & ~x762;
assign c6402 =  x67 &  x92 &  x95 &  x119 &  x157 &  x206 &  x545 &  x580 &  x651 &  x657 & ~x2 & ~x111 & ~x135 & ~x141 & ~x194 & ~x251 & ~x277 & ~x363 & ~x367 & ~x447 & ~x473 & ~x755 & ~x757;
assign c6404 = ~x569 & ~x698;
assign c6406 = ~x504 & ~x675;
assign c6408 = ~x1 & ~x297 & ~x466 & ~x711;
assign c6410 = ~x26 & ~x30 & ~x55 & ~x81 & ~x109 & ~x111 & ~x112 & ~x114 & ~x117 & ~x144 & ~x145 & ~x172 & ~x191 & ~x197 & ~x221 & ~x249 & ~x252 & ~x277 & ~x304 & ~x310 & ~x333 & ~x338 & ~x390 & ~x392 & ~x418 & ~x421 & ~x446 & ~x448 & ~x477 & ~x671 & ~x679 & ~x698 & ~x726 & ~x728 & ~x730 & ~x740 & ~x755 & ~x761 & ~x782;
assign c6412 =  x64 &  x133 &  x161 &  x300 &  x315 &  x387 &  x596 & ~x1 & ~x108 & ~x138 & ~x144 & ~x194 & ~x223 & ~x280;
assign c6414 =  x716 & ~x18 & ~x30 & ~x37 & ~x57 & ~x60 & ~x84 & ~x392 & ~x588 & ~x608;
assign c6416 =  x118 &  x174 &  x175 &  x507 & ~x2 & ~x26 & ~x30 & ~x80 & ~x112 & ~x141 & ~x197 & ~x474 & ~x475 & ~x476 & ~x503 & ~x532 & ~x559 & ~x646 & ~x672 & ~x699 & ~x724 & ~x781;
assign c6418 =  x40 & ~x4 & ~x10 & ~x17 & ~x20 & ~x23 & ~x24 & ~x46 & ~x49 & ~x54 & ~x59 & ~x60 & ~x82 & ~x85 & ~x86 & ~x109 & ~x111 & ~x112 & ~x136 & ~x144 & ~x168 & ~x171 & ~x193 & ~x221 & ~x223 & ~x224 & ~x227 & ~x249 & ~x278 & ~x282 & ~x310 & ~x333 & ~x359 & ~x363 & ~x364 & ~x365 & ~x391 & ~x395 & ~x417 & ~x420 & ~x421 & ~x449 & ~x450 & ~x472 & ~x476 & ~x478 & ~x501 & ~x504 & ~x530 & ~x533 & ~x535 & ~x559 & ~x561 & ~x586 & ~x588 & ~x590 & ~x613 & ~x644 & ~x647 & ~x672 & ~x674 & ~x699 & ~x701 & ~x725 & ~x726 & ~x729 & ~x748 & ~x756 & ~x759 & ~x761 & ~x781;
assign c6420 =  x373 &  x409 &  x517 &  x579 & ~x49 & ~x87 & ~x138 & ~x140 & ~x166 & ~x171 & ~x334 & ~x337 & ~x338 & ~x361 & ~x391 & ~x417 & ~x446 & ~x447 & ~x504 & ~x643 & ~x721 & ~x748 & ~x749 & ~x760 & ~x762 & ~x780;
assign c6422 =  x329 &  x330 &  x459 & ~x24 & ~x53 & ~x195 & ~x563 & ~x587 & ~x611 & ~x669 & ~x674 & ~x761;
assign c6424 =  x231 &  x367 & ~x1 & ~x3 & ~x14 & ~x308;
assign c6426 =  x63 &  x552 &  x580 & ~x1 & ~x32 & ~x140 & ~x142 & ~x194 & ~x196 & ~x222 & ~x504 & ~x589 & ~x727 & ~x729 & ~x736 & ~x777;
assign c6428 =  x92 &  x713 & ~x23 & ~x26 & ~x31 & ~x37 & ~x38 & ~x83 & ~x310 & ~x367 & ~x417 & ~x447 & ~x474 & ~x502 & ~x697 & ~x728 & ~x753;
assign c6430 =  x47 & ~x0 & ~x12 & ~x14 & ~x25 & ~x30 & ~x138 & ~x168 & ~x170 & ~x199 & ~x223 & ~x250 & ~x281 & ~x336 & ~x366 & ~x425 & ~x450 & ~x588 & ~x612;
assign c6432 =  x119 & ~x1 & ~x4 & ~x26 & ~x31 & ~x42 & ~x81 & ~x82 & ~x83 & ~x87 & ~x111 & ~x222 & ~x223 & ~x251 & ~x252 & ~x307 & ~x475 & ~x756 & ~x757;
assign c6434 = ~x193 & ~x213 & ~x418 & ~x460 & ~x540 & ~x613;
assign c6436 =  x123 &  x177 &  x262 &  x271 &  x354 &  x401 &  x432 &  x435 &  x439 &  x519 &  x630 &  x709 & ~x6 & ~x59 & ~x107 & ~x136 & ~x137 & ~x193 & ~x252 & ~x335 & ~x339 & ~x361 & ~x416 & ~x419 & ~x422 & ~x470 & ~x482 & ~x647 & ~x668 & ~x670 & ~x674;
assign c6438 =  x310;
assign c6440 =  x300 & ~x23 & ~x27 & ~x28 & ~x53 & ~x55 & ~x57 & ~x59 & ~x81 & ~x85 & ~x86 & ~x101 & ~x110 & ~x167 & ~x168 & ~x223 & ~x251 & ~x279 & ~x308 & ~x391 & ~x447 & ~x503 & ~x613 & ~x642 & ~x643 & ~x645 & ~x701 & ~x726 & ~x728 & ~x729 & ~x730 & ~x756 & ~x758 & ~x761 & ~x763 & ~x781 & ~x782 & ~x783;
assign c6442 =  x12 &  x74 &  x91 &  x154 & ~x37 & ~x280 & ~x783;
assign c6444 =  x103 & ~x4 & ~x7 & ~x18 & ~x22 & ~x26 & ~x78 & ~x80 & ~x108 & ~x140 & ~x142 & ~x196 & ~x221 & ~x251 & ~x252 & ~x361 & ~x363 & ~x420 & ~x532 & ~x587 & ~x707 & ~x729 & ~x754 & ~x757 & ~x764 & ~x765 & ~x774 & ~x777 & ~x779 & ~x780 & ~x781 & ~x783;
assign c6446 =  x298 &  x574 & ~x140 & ~x166 & ~x249 & ~x285 & ~x553 & ~x557 & ~x581 & ~x583 & ~x591 & ~x638 & ~x640 & ~x755;
assign c6448 =  x632 & ~x83 & ~x98 & ~x221 & ~x392 & ~x648;
assign c6450 =  x244 &  x439 &  x546 &  x570 &  x580 & ~x0 & ~x1 & ~x3 & ~x5 & ~x23 & ~x54 & ~x84 & ~x108 & ~x113 & ~x114 & ~x115 & ~x137 & ~x141 & ~x164 & ~x196 & ~x224 & ~x502 & ~x534 & ~x582 & ~x590 & ~x615 & ~x616 & ~x618 & ~x645 & ~x647 & ~x668 & ~x728 & ~x732 & ~x752;
assign c6452 =  x43 &  x299 &  x326 &  x652 & ~x256 & ~x281 & ~x311 & ~x359 & ~x526 & ~x588 & ~x779;
assign c6454 =  x42 &  x43 &  x69 &  x769 & ~x6 & ~x7 & ~x21 & ~x24 & ~x27 & ~x28 & ~x34 & ~x49 & ~x52 & ~x53 & ~x54 & ~x56 & ~x59 & ~x85 & ~x88 & ~x108 & ~x111 & ~x112 & ~x113 & ~x115 & ~x135 & ~x136 & ~x139 & ~x164 & ~x165 & ~x166 & ~x167 & ~x168 & ~x171 & ~x192 & ~x194 & ~x196 & ~x197 & ~x223 & ~x250 & ~x255 & ~x333 & ~x336 & ~x337 & ~x361 & ~x362 & ~x366 & ~x394 & ~x419 & ~x421 & ~x422 & ~x475 & ~x501 & ~x503 & ~x506 & ~x530 & ~x532 & ~x533 & ~x534 & ~x558 & ~x614 & ~x615 & ~x642 & ~x643 & ~x644 & ~x670 & ~x699 & ~x701 & ~x728 & ~x754 & ~x755 & ~x758 & ~x759 & ~x781 & ~x782;
assign c6456 =  x79;
assign c6458 =  x74 &  x105 &  x238 &  x331 &  x556 &  x566 &  x582 & ~x4 & ~x25 & ~x83 & ~x136 & ~x194 & ~x283 & ~x334 & ~x420;
assign c6460 =  x261 &  x269 &  x439 &  x456 &  x652 &  x658 & ~x7 & ~x21 & ~x22 & ~x24 & ~x192 & ~x193 & ~x226 & ~x228 & ~x313 & ~x556 & ~x613 & ~x751 & ~x780;
assign c6462 = ~x0 & ~x28 & ~x81 & ~x112 & ~x197 & ~x199 & ~x227 & ~x248 & ~x254 & ~x275 & ~x276 & ~x278 & ~x304 & ~x310 & ~x333 & ~x339 & ~x363 & ~x365 & ~x391 & ~x421 & ~x422 & ~x445 & ~x474 & ~x476 & ~x562 & ~x614 & ~x643 & ~x672 & ~x699 & ~x705 & ~x710 & ~x727 & ~x780;
assign c6466 =  x259 &  x528 & ~x172 & ~x191 & ~x278 & ~x309 & ~x334 & ~x361;
assign c6468 =  x47 &  x259 &  x296 &  x303 &  x343 &  x399 &  x406 & ~x0 & ~x82;
assign c6470 =  x13 &  x104 &  x239 &  x241 &  x295 &  x403 &  x404 &  x583 &  x597 &  x604 &  x635 &  x715 & ~x19 & ~x364;
assign c6472 =  x142;
assign c6474 =  x35 & ~x3 & ~x4 & ~x12 & ~x14 & ~x16 & ~x24 & ~x27 & ~x31 & ~x57 & ~x59 & ~x81 & ~x83 & ~x86 & ~x110 & ~x113 & ~x114 & ~x138 & ~x169 & ~x308 & ~x335 & ~x336 & ~x423 & ~x477 & ~x506 & ~x560 & ~x589 & ~x646 & ~x672 & ~x673 & ~x729 & ~x755 & ~x756 & ~x780;
assign c6476 =  x147 &  x273 &  x382 &  x430 &  x458 &  x514 &  x602 &  x653 & ~x28 & ~x29 & ~x45 & ~x47 & ~x54 & ~x56 & ~x85 & ~x110 & ~x251 & ~x390 & ~x419 & ~x503 & ~x532 & ~x780;
assign c6478 =  x67 &  x95 &  x97 &  x104 &  x149 &  x160 &  x213 &  x215 &  x232 &  x269 &  x271 &  x297 &  x299 &  x347 &  x348 &  x350 &  x354 &  x374 &  x379 &  x382 &  x519 &  x521 &  x544 &  x596 &  x603 &  x625 &  x632 &  x657 &  x659 &  x681 &  x682 &  x770 & ~x6 & ~x34 & ~x52 & ~x83 & ~x140 & ~x171 & ~x194 & ~x251 & ~x254 & ~x278 & ~x309 & ~x360 & ~x420 & ~x588 & ~x589 & ~x700 & ~x757;
assign c6480 =  x43 &  x99 &  x119 &  x132 &  x386 & ~x19 & ~x31 & ~x37 & ~x46 & ~x55 & ~x79 & ~x195 & ~x221 & ~x222 & ~x339 & ~x422 & ~x589;
assign c6482 =  x34;
assign c6484 = ~x214 & ~x459;
assign c6486 =  x144 &  x301 & ~x779;
assign c6488 =  x40 & ~x4 & ~x5 & ~x17 & ~x33 & ~x36 & ~x37 & ~x38 & ~x46 & ~x48 & ~x49 & ~x55 & ~x57 & ~x64 & ~x76 & ~x83 & ~x86 & ~x87 & ~x88 & ~x107 & ~x110 & ~x111 & ~x138 & ~x166 & ~x168 & ~x169 & ~x193 & ~x194 & ~x197 & ~x222 & ~x250 & ~x279 & ~x280 & ~x305 & ~x334 & ~x361 & ~x364 & ~x365 & ~x388 & ~x390 & ~x393 & ~x417 & ~x418 & ~x421 & ~x449 & ~x477 & ~x502 & ~x503 & ~x504 & ~x558 & ~x560 & ~x587 & ~x675 & ~x698 & ~x699 & ~x725 & ~x727 & ~x729 & ~x748 & ~x753 & ~x757 & ~x758 & ~x775 & ~x776 & ~x781 & ~x782 & ~x783;
assign c6490 =  x344 &  x349 &  x351 &  x354 &  x484 &  x495 &  x664 &  x679 & ~x1 & ~x2 & ~x5 & ~x7 & ~x20 & ~x23 & ~x26 & ~x27 & ~x28 & ~x30 & ~x33 & ~x53 & ~x54 & ~x57 & ~x59 & ~x60 & ~x80 & ~x83 & ~x86 & ~x110 & ~x137 & ~x196 & ~x251 & ~x363 & ~x364 & ~x419 & ~x584 & ~x588 & ~x592 & ~x593 & ~x612 & ~x645 & ~x669 & ~x671 & ~x675 & ~x700 & ~x701 & ~x702 & ~x727 & ~x730 & ~x753 & ~x755 & ~x757 & ~x760 & ~x781 & ~x782;
assign c6492 =  x259 &  x372 & ~x6 & ~x19 & ~x23 & ~x26 & ~x29 & ~x37 & ~x45 & ~x53 & ~x56 & ~x57 & ~x82 & ~x83 & ~x84 & ~x112 & ~x114 & ~x136 & ~x137 & ~x169 & ~x250 & ~x308 & ~x335 & ~x336 & ~x392 & ~x619 & ~x643 & ~x673;
assign c6494 =  x119 &  x455 &  x684 & ~x4 & ~x10 & ~x32 & ~x46 & ~x83 & ~x167 & ~x195 & ~x196 & ~x504 & ~x532 & ~x534 & ~x557 & ~x559 & ~x588 & ~x590 & ~x618 & ~x641 & ~x647 & ~x669 & ~x671 & ~x673 & ~x726;
assign c6496 =  x104 &  x264 &  x538 & ~x114 & ~x219 & ~x474 & ~x477 & ~x765;
assign c6498 = ~x23 & ~x26 & ~x28 & ~x53 & ~x82 & ~x114 & ~x169 & ~x450 & ~x475 & ~x502 & ~x505 & ~x590 & ~x656 & ~x673 & ~x698 & ~x757 & ~x777;
assign c61 =  x38 &  x120 &  x121 &  x122 &  x131 &  x134 &  x149 &  x173 &  x256 &  x260 &  x273 &  x275 &  x577 & ~x31 & ~x51 & ~x83 & ~x114 & ~x140 & ~x170 & ~x194 & ~x253 & ~x362 & ~x418 & ~x476 & ~x502 & ~x503 & ~x531 & ~x561 & ~x643 & ~x645 & ~x671 & ~x730;
assign c63 =  x1;
assign c65 = ~x8 & ~x18 & ~x105 & ~x116 & ~x341 & ~x559 & ~x563 & ~x643 & ~x648 & ~x650 & ~x665 & ~x667 & ~x679 & ~x692 & ~x696 & ~x699 & ~x723;
assign c67 =  x121 &  x187 &  x375 &  x379 &  x431 &  x488 &  x515 &  x603 &  x629 &  x654 &  x660 &  x683 &  x687 &  x689 &  x711 &  x712 &  x713 &  x717 &  x741 & ~x8 & ~x22 & ~x23 & ~x26 & ~x32 & ~x51 & ~x54 & ~x111 & ~x141 & ~x193 & ~x251 & ~x282 & ~x333 & ~x334 & ~x364 & ~x389 & ~x394 & ~x423 & ~x472 & ~x478 & ~x479 & ~x532 & ~x561 & ~x563 & ~x587 & ~x588 & ~x613 & ~x619 & ~x620 & ~x668 & ~x694 & ~x698 & ~x700 & ~x705 & ~x706 & ~x721;
assign c69 =  x301 &  x329 &  x413 &  x469 &  x750 & ~x9 & ~x21 & ~x58 & ~x164 & ~x276 & ~x310 & ~x445 & ~x506 & ~x561 & ~x562 & ~x671 & ~x697 & ~x741 & ~x744 & ~x746 & ~x770;
assign c611 =  x420;
assign c613 =  x146 &  x229 &  x273 &  x287 &  x320 &  x341 &  x350 &  x353 &  x431 &  x437 &  x462 &  x463 &  x485 &  x486 &  x493 &  x526 &  x555 &  x583 &  x639 &  x649 &  x695 &  x705 & ~x9 & ~x19 & ~x25 & ~x26 & ~x54 & ~x85 & ~x115 & ~x167 & ~x253 & ~x308 & ~x310 & ~x337 & ~x505 & ~x534 & ~x585 & ~x614 & ~x617 & ~x702 & ~x727 & ~x730 & ~x753 & ~x758 & ~x769 & ~x771;
assign c615 =  x589;
assign c617 =  x39 &  x41 &  x43 &  x45 &  x232 &  x301 &  x346 &  x414 &  x431 &  x548 &  x572 &  x629 &  x635 &  x653 & ~x33 & ~x61 & ~x139 & ~x199 & ~x277 & ~x394 & ~x475 & ~x501 & ~x557 & ~x699 & ~x725 & ~x729 & ~x731 & ~x754;
assign c619 =  x197;
assign c621 =  x27;
assign c623 =  x504;
assign c625 =  x253;
assign c627 =  x726;
assign c629 =  x54;
assign c631 =  x42 &  x70 &  x72 &  x124 &  x126 &  x155 &  x157 &  x159 &  x176 &  x186 &  x205 &  x215 &  x216 &  x217 &  x237 &  x268 &  x273 &  x297 &  x352 &  x354 &  x409 &  x430 &  x487 &  x488 &  x494 &  x521 &  x548 &  x550 &  x568 &  x605 &  x627 &  x657 & ~x35 & ~x61 & ~x86 & ~x109 & ~x110 & ~x112 & ~x113 & ~x144 & ~x164 & ~x198 & ~x277 & ~x283 & ~x311 & ~x389 & ~x421 & ~x446 & ~x477 & ~x478 & ~x532 & ~x563 & ~x587 & ~x591 & ~x615 & ~x616 & ~x673 & ~x697 & ~x698 & ~x703 & ~x725 & ~x753 & ~x755 & ~x758 & ~x782;
assign c633 =  x783;
assign c635 =  x781;
assign c637 =  x228 &  x591;
assign c639 =  x571 &  x738 &  x740 & ~x0 & ~x28 & ~x220 & ~x221 & ~x306 & ~x307 & ~x414 & ~x425 & ~x442 & ~x443 & ~x446 & ~x448 & ~x451 & ~x452 & ~x472 & ~x478 & ~x481 & ~x527 & ~x530 & ~x537 & ~x556 & ~x593 & ~x611 & ~x616 & ~x617 & ~x619 & ~x621 & ~x638 & ~x639 & ~x641 & ~x645 & ~x647 & ~x651 & ~x666 & ~x668 & ~x670 & ~x679 & ~x693 & ~x707 & ~x722 & ~x723 & ~x732 & ~x759 & ~x777 & ~x779 & ~x782;
assign c641 =  x127 &  x153 &  x576 & ~x162 & ~x173 & ~x246 & ~x284 & ~x414 & ~x533 & ~x592 & ~x695;
assign c643 = ~x145 & ~x602 & ~x629 & ~x742;
assign c645 =  x126 &  x181 & ~x62 & ~x63 & ~x75 & ~x134 & ~x163 & ~x164 & ~x190 & ~x253 & ~x275 & ~x556;
assign c647 =  x736 & ~x356 & ~x412;
assign c649 =  x783;
assign c651 = ~x70 & ~x98 & ~x104 & ~x181;
assign c653 =  x467 &  x468 &  x497 &  x547 & ~x0 & ~x62 & ~x91;
assign c655 =  x30;
assign c657 =  x687 & ~x8 & ~x9 & ~x18 & ~x20 & ~x24 & ~x36 & ~x51 & ~x54 & ~x55 & ~x78 & ~x80 & ~x89 & ~x90 & ~x91 & ~x92 & ~x106 & ~x143 & ~x144 & ~x145 & ~x225 & ~x256 & ~x334 & ~x364 & ~x389 & ~x448 & ~x559 & ~x586 & ~x669 & ~x702 & ~x730;
assign c659 =  x728;
assign c661 =  x122 &  x129 &  x130 &  x147 &  x148 &  x217 &  x268 &  x274 &  x301 &  x313 &  x314 &  x317 &  x326 &  x355 &  x357 &  x358 &  x374 &  x398 &  x400 &  x429 &  x439 &  x442 &  x469 &  x510 &  x512 &  x525 &  x542 &  x546 &  x549 &  x568 & ~x20 & ~x24 & ~x81 & ~x109 & ~x112 & ~x166 & ~x192 & ~x221 & ~x248 & ~x250 & ~x255 & ~x394 & ~x417 & ~x422 & ~x505 & ~x529 & ~x530 & ~x562 & ~x644 & ~x646 & ~x727 & ~x730 & ~x753 & ~x755 & ~x759;
assign c663 =  x201 &  x257 &  x439 &  x648 &  x751 & ~x222 & ~x725;
assign c665 =  x448;
assign c667 =  x157 &  x380 &  x404 &  x436 &  x487 &  x492 &  x543 &  x603 &  x628 &  x655 &  x656 &  x657 & ~x4 & ~x9 & ~x18 & ~x75 & ~x76 & ~x87 & ~x107 & ~x137 & ~x195 & ~x227 & ~x304 & ~x305 & ~x364 & ~x392 & ~x419 & ~x476 & ~x477 & ~x503 & ~x506 & ~x532 & ~x559 & ~x562 & ~x616 & ~x671 & ~x757 & ~x763;
assign c669 =  x14 &  x16 &  x273 &  x568 &  x626 &  x680 & ~x24 & ~x31 & ~x110 & ~x279 & ~x306 & ~x362 & ~x476 & ~x503 & ~x558 & ~x617 & ~x727 & ~x759 & ~x781 & ~x782;
assign c671 =  x2;
assign c673 = ~x19 & ~x66 & ~x70 & ~x91 & ~x118 & ~x119 & ~x146;
assign c675 =  x1;
assign c677 =  x392;
assign c679 =  x252;
assign c681 =  x38 &  x98 & ~x416 & ~x528 & ~x563 & ~x580 & ~x669 & ~x673;
assign c683 =  x56;
assign c685 =  x755;
assign c687 =  x55;
assign c689 =  x27;
assign c691 =  x38 &  x123 &  x191 &  x243 &  x302 &  x625 & ~x393 & ~x447 & ~x529 & ~x730;
assign c693 =  x167;
assign c695 =  x27;
assign c697 =  x82;
assign c699 =  x84;
assign c6101 =  x252;
assign c6103 = ~x44 & ~x216 & ~x287 & ~x288 & ~x313;
assign c6105 =  x38 &  x39 &  x45 &  x147 &  x177 &  x325 &  x347 &  x435 &  x461 &  x522 &  x543 &  x576 &  x598 &  x627 &  x628 &  x654 &  x657 &  x690 & ~x3 & ~x25 & ~x59 & ~x107 & ~x109 & ~x110 & ~x113 & ~x136 & ~x137 & ~x144 & ~x165 & ~x168 & ~x169 & ~x223 & ~x277 & ~x279 & ~x280 & ~x305 & ~x308 & ~x334 & ~x363 & ~x419 & ~x422 & ~x449 & ~x473 & ~x476 & ~x501 & ~x502 & ~x505 & ~x507 & ~x533 & ~x534 & ~x535 & ~x559 & ~x563 & ~x588 & ~x618 & ~x642 & ~x699 & ~x703 & ~x725;
assign c6107 =  x39 &  x46 &  x70 &  x319 & ~x137 & ~x483 & ~x539;
assign c6109 =  x168;
assign c6111 =  x41 &  x76 &  x93 &  x101 &  x162 &  x174 &  x187 &  x229 &  x245 &  x246 &  x247 &  x258 &  x260 &  x402 &  x493 &  x523 &  x572 &  x634 & ~x8 & ~x23 & ~x113 & ~x138 & ~x141 & ~x280 & ~x446 & ~x532 & ~x558 & ~x559 & ~x783;
assign c6113 =  x757;
assign c6117 =  x190 &  x313 &  x356 &  x544 & ~x63 & ~x671 & ~x770;
assign c6119 = ~x67 & ~x97 & ~x147;
assign c6121 =  x57;
assign c6123 =  x192 & ~x694;
assign c6125 =  x420;
assign c6127 =  x42 &  x44 &  x214 &  x216 &  x288 &  x294 &  x319 &  x461 &  x463 &  x577 &  x634 &  x682 &  x688 & ~x3 & ~x7 & ~x25 & ~x35 & ~x110 & ~x113 & ~x138 & ~x222 & ~x249 & ~x277 & ~x279 & ~x333 & ~x334 & ~x335 & ~x389 & ~x391 & ~x392 & ~x417 & ~x423 & ~x450 & ~x451 & ~x474 & ~x530 & ~x532 & ~x564 & ~x617 & ~x619 & ~x642 & ~x644 & ~x675 & ~x696 & ~x698 & ~x704 & ~x780;
assign c6129 =  x383 &  x384 & ~x10 & ~x35 & ~x36 & ~x62 & ~x64 & ~x91 & ~x92;
assign c6131 =  x14 &  x94 &  x127 &  x426 &  x427 &  x430 &  x544 & ~x62 & ~x106 & ~x165 & ~x727;
assign c6133 =  x41 &  x63 &  x118 &  x121 &  x172 &  x173 &  x200 &  x256 &  x257 &  x568 &  x573 &  x597 & ~x365 & ~x366;
assign c6135 =  x54;
assign c6137 =  x318 &  x373 &  x517 &  x598 &  x607 &  x654 &  x708 &  x709 &  x710 &  x736 &  x737 &  x738 &  x764 &  x765 &  x766 &  x773 & ~x3 & ~x4 & ~x198 & ~x225 & ~x308 & ~x420 & ~x421 & ~x474 & ~x476 & ~x586 & ~x590 & ~x757;
assign c6139 = ~x201 & ~x244 & ~x261;
assign c6141 =  x71 &  x258 &  x709 &  x710 &  x711 &  x774 &  x775 & ~x80 & ~x558;
assign c6143 =  x392;
assign c6145 =  x476;
assign c6147 = ~x258 & ~x260 & ~x300 & ~x454;
assign c6149 =  x51 & ~x97;
assign c6151 =  x448;
assign c6153 =  x231 &  x324 &  x385 &  x498 &  x582 & ~x54 & ~x641 & ~x669 & ~x670 & ~x714 & ~x715 & ~x739 & ~x741 & ~x753;
assign c6155 =  x39 &  x45 &  x126 &  x129 &  x179 &  x238 &  x240 &  x259 &  x272 &  x273 &  x374 &  x408 &  x432 &  x437 &  x514 &  x521 &  x543 &  x578 &  x626 &  x627 &  x653 &  x662 & ~x0 & ~x3 & ~x28 & ~x59 & ~x89 & ~x107 & ~x167 & ~x172 & ~x255 & ~x311 & ~x416 & ~x445 & ~x475 & ~x529 & ~x531 & ~x532 & ~x589 & ~x590 & ~x618 & ~x647 & ~x669 & ~x673 & ~x725 & ~x758 & ~x780;
assign c6157 =  x252;
assign c6159 =  x28;
assign c6161 =  x128 &  x149 &  x152 &  x177 &  x229 &  x341 &  x386 &  x521 &  x626 &  x661 &  x691 & ~x32 & ~x86 & ~x139 & ~x143 & ~x227 & ~x445 & ~x534 & ~x557 & ~x613 & ~x769 & ~x772;
assign c6163 =  x11 &  x16 & ~x0 & ~x53 & ~x81 & ~x113 & ~x141 & ~x251 & ~x308 & ~x394 & ~x471 & ~x473 & ~x480 & ~x502 & ~x504 & ~x587 & ~x618 & ~x619 & ~x647 & ~x669 & ~x673 & ~x700 & ~x727 & ~x780;
assign c6165 =  x656 &  x740 & ~x89 & ~x201 & ~x230 & ~x231;
assign c6167 =  x486 &  x654 & ~x300;
assign c6169 =  x112;
assign c6171 = ~x42 & ~x89 & ~x174 & ~x177 & ~x204;
assign c6173 =  x83;
assign c6175 =  x341 &  x359 &  x368 &  x381 &  x458 &  x554 &  x582 &  x621 &  x733 & ~x136 & ~x194 & ~x699 & ~x753;
assign c6177 =  x224;
assign c6179 =  x251;
assign c6181 =  x392;
assign c6183 =  x71 &  x74 &  x103 &  x148 &  x320 &  x465 &  x598 &  x606 &  x634 &  x716 &  x744 & ~x115 & ~x420 & ~x506 & ~x536 & ~x587 & ~x612 & ~x616 & ~x671 & ~x693 & ~x695 & ~x721 & ~x761 & ~x778;
assign c6185 =  x26;
assign c6187 =  x140;
assign c6189 =  x82;
assign c6191 =  x759;
assign c6193 =  x22;
assign c6195 =  x476;
assign c6197 =  x111;
assign c6199 =  x392;
assign c6201 =  x259 &  x432 &  x464 &  x466 &  x485 &  x523 &  x540 &  x551 &  x568 &  x573 &  x576 &  x607 &  x628 &  x630 &  x659 &  x682 &  x684 &  x711 &  x714 &  x742 & ~x1 & ~x25 & ~x29 & ~x32 & ~x54 & ~x81 & ~x110 & ~x114 & ~x163 & ~x165 & ~x168 & ~x170 & ~x193 & ~x223 & ~x250 & ~x279 & ~x281 & ~x282 & ~x332 & ~x335 & ~x360 & ~x362 & ~x366 & ~x446 & ~x474 & ~x501 & ~x504 & ~x506 & ~x529 & ~x530 & ~x558 & ~x587 & ~x614 & ~x616 & ~x617 & ~x644 & ~x669 & ~x675 & ~x702 & ~x726 & ~x728;
assign c6203 =  x728;
assign c6205 =  x476;
assign c6207 =  x46 &  x74 &  x92 &  x94 &  x187 &  x319 &  x375 &  x410 &  x464 &  x492 &  x522 &  x625 &  x633 &  x634 & ~x26 & ~x52 & ~x53 & ~x55 & ~x58 & ~x114 & ~x138 & ~x143 & ~x223 & ~x305 & ~x361 & ~x391 & ~x418 & ~x422 & ~x450 & ~x504 & ~x557 & ~x585 & ~x587 & ~x590 & ~x613 & ~x616 & ~x645 & ~x673 & ~x701 & ~x725 & ~x757 & ~x770;
assign c6209 =  x180 &  x190 &  x208 &  x210 &  x215 &  x216 &  x218 &  x244 &  x262 &  x263 &  x268 &  x274 &  x287 &  x289 &  x294 &  x298 &  x318 &  x323 &  x326 &  x330 &  x385 &  x386 &  x397 &  x404 &  x405 &  x406 &  x430 &  x439 &  x453 &  x458 &  x459 &  x460 &  x467 &  x471 &  x491 &  x513 &  x516 &  x541 &  x543 &  x545 &  x549 &  x554 &  x555 &  x573 &  x605 & ~x1 & ~x5 & ~x28 & ~x30 & ~x54 & ~x60 & ~x61 & ~x110 & ~x111 & ~x167 & ~x615 & ~x617 & ~x673 & ~x674 & ~x702 & ~x753 & ~x767 & ~x770 & ~x771;
assign c6211 =  x159 &  x204 &  x232 &  x239 &  x241 &  x267 &  x272 &  x296 &  x321 &  x322 &  x377 &  x460 &  x489 &  x492 &  x493 &  x550 &  x575 &  x576 &  x686 &  x710 &  x713 &  x714 &  x741 & ~x22 & ~x60 & ~x84 & ~x138 & ~x139 & ~x196 & ~x198 & ~x250 & ~x282 & ~x338 & ~x417 & ~x475 & ~x507 & ~x530 & ~x622 & ~x640 & ~x648 & ~x668 & ~x696 & ~x701 & ~x702 & ~x722 & ~x727 & ~x733 & ~x734 & ~x752 & ~x757 & ~x759 & ~x760 & ~x761;
assign c6213 =  x39 &  x76 & ~x4 & ~x25 & ~x32 & ~x83 & ~x112 & ~x138 & ~x141 & ~x142 & ~x309 & ~x362 & ~x393 & ~x419 & ~x475 & ~x505 & ~x507 & ~x557 & ~x563 & ~x637 & ~x672 & ~x698 & ~x730 & ~x754;
assign c6215 =  x267 & ~x116 & ~x256 & ~x456 & ~x508;
assign c6217 =  x379 & ~x33 & ~x64 & ~x144 & ~x652 & ~x692 & ~x703;
assign c6219 =  x98 &  x99 &  x125 &  x153 &  x182 &  x236 &  x347 &  x576 &  x604 &  x684 & ~x31 & ~x49 & ~x62 & ~x106 & ~x146 & ~x173 & ~x194 & ~x256 & ~x332 & ~x366 & ~x418 & ~x421 & ~x477 & ~x478 & ~x616 & ~x726 & ~x729 & ~x756;
assign c6221 =  x14 &  x15 &  x16 &  x151 & ~x23 & ~x30 & ~x53 & ~x56 & ~x86 & ~x87 & ~x111 & ~x139 & ~x195 & ~x254 & ~x449 & ~x616 & ~x617 & ~x770 & ~x772;
assign c6223 =  x763;
assign c6225 =  x219 &  x528 &  x570 &  x625 & ~x671 & ~x772;
assign c6227 =  x587;
assign c6229 =  x308;
assign c6231 =  x94 &  x122 &  x127 &  x153 &  x187 &  x320 &  x380 &  x402 &  x433 &  x460 &  x465 &  x514 &  x548 &  x598 &  x599 &  x628 &  x632 &  x633 &  x655 &  x682 &  x688 &  x689 &  x711 &  x739 &  x745 & ~x0 & ~x35 & ~x54 & ~x56 & ~x80 & ~x82 & ~x83 & ~x110 & ~x111 & ~x140 & ~x167 & ~x169 & ~x195 & ~x222 & ~x224 & ~x225 & ~x278 & ~x311 & ~x337 & ~x339 & ~x362 & ~x364 & ~x367 & ~x388 & ~x390 & ~x419 & ~x445 & ~x447 & ~x472 & ~x474 & ~x476 & ~x480 & ~x501 & ~x502 & ~x507 & ~x585 & ~x586 & ~x589 & ~x614 & ~x615 & ~x616 & ~x619 & ~x645 & ~x676 & ~x698 & ~x729 & ~x730 & ~x733 & ~x734 & ~x750 & ~x752 & ~x755 & ~x759;
assign c6233 =  x44 &  x121 &  x124 &  x130 &  x154 &  x188 &  x207 &  x211 &  x212 &  x403 &  x459 &  x485 &  x542 &  x549 &  x550 &  x551 & ~x21 & ~x25 & ~x50 & ~x60 & ~x90 & ~x105 & ~x106 & ~x143 & ~x163 & ~x191 & ~x197 & ~x225 & ~x226 & ~x304 & ~x334 & ~x336 & ~x338 & ~x449 & ~x478 & ~x613 & ~x702 & ~x728;
assign c6235 =  x251;
assign c6237 =  x13 &  x482 &  x483 &  x511 &  x521 &  x566 &  x567 &  x580 & ~x106 & ~x277;
assign c6239 =  x252;
assign c6241 =  x174 &  x245 &  x259 &  x705 &  x722 &  x750 & ~x51 & ~x61 & ~x79 & ~x80 & ~x108 & ~x111 & ~x170 & ~x193 & ~x195 & ~x221 & ~x308 & ~x309 & ~x333 & ~x337 & ~x420 & ~x445 & ~x473 & ~x476 & ~x503 & ~x561 & ~x643 & ~x645 & ~x646 & ~x671 & ~x730 & ~x743 & ~x744 & ~x753 & ~x763 & ~x764 & ~x766 & ~x767 & ~x769;
assign c6243 =  x29;
assign c6245 =  x589;
assign c6247 =  x314 &  x315 &  x355 &  x408 &  x466 &  x468 &  x567 &  x568 &  x573 &  x657 & ~x62 & ~x76 & ~x140 & ~x199 & ~x558;
assign c6249 =  x196;
assign c6251 =  x448;
assign c6253 =  x67 &  x145 &  x201 &  x439 &  x521 &  x541 &  x631 & ~x29 & ~x86 & ~x449 & ~x553 & ~x728;
assign c6255 =  x126 &  x128 &  x184 &  x293 &  x351 &  x352 &  x377 &  x403 &  x408 &  x431 &  x489 &  x494 &  x521 &  x543 &  x548 &  x549 &  x661 &  x685 & ~x7 & ~x22 & ~x25 & ~x33 & ~x54 & ~x59 & ~x84 & ~x169 & ~x251 & ~x280 & ~x310 & ~x338 & ~x363 & ~x364 & ~x366 & ~x390 & ~x393 & ~x420 & ~x424 & ~x445 & ~x448 & ~x452 & ~x471 & ~x499 & ~x502 & ~x533 & ~x559 & ~x613 & ~x614 & ~x619 & ~x644 & ~x649 & ~x677 & ~x693 & ~x698 & ~x721 & ~x725 & ~x730 & ~x731 & ~x732 & ~x753 & ~x756;
assign c6257 =  x70 &  x94 &  x97 &  x130 &  x159 &  x204 &  x319 &  x374 &  x402 &  x435 &  x460 &  x542 &  x550 &  x711 &  x717 &  x718 & ~x2 & ~x24 & ~x25 & ~x80 & ~x84 & ~x196 & ~x391 & ~x393 & ~x395 & ~x416 & ~x424 & ~x447 & ~x471 & ~x527 & ~x530 & ~x585 & ~x610 & ~x617 & ~x641 & ~x645 & ~x650 & ~x704 & ~x730 & ~x734 & ~x758;
assign c6259 =  x392;
assign c6261 =  x16 & ~x386 & ~x538 & ~x622;
assign c6263 = ~x509 & ~x579 & ~x580 & ~x678;
assign c6265 =  x215 & ~x332 & ~x448 & ~x552 & ~x556 & ~x584 & ~x608 & ~x619 & ~x753;
assign c6267 =  x167;
assign c6269 =  x16 &  x38 &  x39 &  x42 &  x43 &  x45 &  x73 &  x94 &  x97 &  x124 &  x211 &  x234 &  x269 &  x654 &  x690 & ~x249 & ~x505 & ~x586;
assign c6271 =  x98 &  x275 &  x325 &  x527 &  x631 &  x705 & ~x137 & ~x559 & ~x730 & ~x769;
assign c6273 =  x41 &  x69 &  x70 & ~x110 & ~x193 & ~x195 & ~x364 & ~x385 & ~x390 & ~x392 & ~x395 & ~x424 & ~x455 & ~x469 & ~x483 & ~x506 & ~x525 & ~x527 & ~x530 & ~x553 & ~x554 & ~x558 & ~x581 & ~x619 & ~x637 & ~x670 & ~x673 & ~x674 & ~x726 & ~x754;
assign c6275 =  x220 &  x276;
assign c6277 =  x4;
assign c6279 =  x487 &  x543 &  x544 &  x628 &  x656 & ~x2 & ~x6 & ~x21 & ~x22 & ~x24 & ~x25 & ~x29 & ~x50 & ~x58 & ~x83 & ~x108 & ~x110 & ~x114 & ~x137 & ~x142 & ~x165 & ~x167 & ~x194 & ~x223 & ~x251 & ~x308 & ~x337 & ~x362 & ~x363 & ~x390 & ~x393 & ~x394 & ~x396 & ~x397 & ~x417 & ~x420 & ~x423 & ~x424 & ~x442 & ~x453 & ~x471 & ~x472 & ~x477 & ~x479 & ~x481 & ~x499 & ~x503 & ~x506 & ~x527 & ~x528 & ~x533 & ~x534 & ~x537 & ~x556 & ~x557 & ~x585 & ~x590 & ~x591 & ~x592 & ~x593 & ~x614 & ~x622 & ~x638 & ~x645 & ~x646 & ~x648 & ~x665 & ~x674 & ~x675 & ~x677 & ~x698 & ~x700 & ~x701 & ~x702 & ~x721 & ~x725 & ~x727 & ~x757 & ~x761 & ~x777 & ~x782;
assign c6281 =  x699;
assign c6283 =  x201 &  x410 &  x569 &  x625 &  x648 & ~x23 & ~x643;
assign c6285 =  x355 &  x438 &  x440 &  x464 &  x466 &  x469 &  x497 &  x539 &  x541 &  x543 &  x550 &  x554 &  x567 &  x581 &  x595 &  x596 &  x610 & ~x0 & ~x36 & ~x57 & ~x58 & ~x76 & ~x78 & ~x81 & ~x83 & ~x85 & ~x727 & ~x756;
assign c6287 =  x336;
assign c6289 =  x308;
assign c6291 =  x740 & ~x4 & ~x9 & ~x23 & ~x31 & ~x32 & ~x50 & ~x59 & ~x79 & ~x140 & ~x142 & ~x166 & ~x198 & ~x249 & ~x279 & ~x282 & ~x311 & ~x339 & ~x341 & ~x367 & ~x368 & ~x395 & ~x443 & ~x503 & ~x537 & ~x561 & ~x563 & ~x590 & ~x595 & ~x667 & ~x677 & ~x694 & ~x699 & ~x730 & ~x752 & ~x760 & ~x762 & ~x778;
assign c6293 =  x56;
assign c6295 =  x656 & ~x3 & ~x4 & ~x27 & ~x28 & ~x34 & ~x59 & ~x60 & ~x108 & ~x111 & ~x116 & ~x142 & ~x168 & ~x194 & ~x197 & ~x254 & ~x277 & ~x282 & ~x305 & ~x307 & ~x309 & ~x365 & ~x366 & ~x367 & ~x368 & ~x395 & ~x397 & ~x425 & ~x445 & ~x446 & ~x449 & ~x473 & ~x478 & ~x503 & ~x507 & ~x508 & ~x528 & ~x534 & ~x555 & ~x564 & ~x612 & ~x614 & ~x619 & ~x648 & ~x650 & ~x651 & ~x665 & ~x667 & ~x668 & ~x676 & ~x698 & ~x701 & ~x705 & ~x707 & ~x722 & ~x725 & ~x727 & ~x750 & ~x755 & ~x756;
assign c6297 =  x783;
assign c6299 = ~x3 & ~x5 & ~x19 & ~x21 & ~x22 & ~x33 & ~x35 & ~x47 & ~x56 & ~x75 & ~x76 & ~x78 & ~x80 & ~x82 & ~x85 & ~x86 & ~x88 & ~x90 & ~x91 & ~x103 & ~x104 & ~x106 & ~x112 & ~x118 & ~x133 & ~x140 & ~x141 & ~x161 & ~x162 & ~x163 & ~x171 & ~x172 & ~x173 & ~x190 & ~x225 & ~x388 & ~x391 & ~x395 & ~x479 & ~x507 & ~x562 & ~x615 & ~x617 & ~x642 & ~x643 & ~x668 & ~x674 & ~x703 & ~x724 & ~x726 & ~x752 & ~x753;
assign c6301 =  x76 &  x93 &  x101 &  x144 &  x626 &  x653 &  x708 &  x709 & ~x51 & ~x59 & ~x137 & ~x140 & ~x308 & ~x420 & ~x502 & ~x586 & ~x617;
assign c6303 =  x278;
assign c6305 =  x251;
assign c6307 =  x88;
assign c6309 = ~x18 & ~x71 & ~x90 & ~x92 & ~x125 & ~x127 & ~x132 & ~x752;
assign c6311 =  x41 &  x202 &  x767 &  x773;
assign c6313 =  x168;
assign c6315 =  x2;
assign c6317 =  x196;
assign c6319 =  x28;
assign c6321 =  x64 &  x77 &  x90 &  x95 &  x172 &  x174 &  x219 &  x573 &  x709 &  x741 & ~x364 & ~x730;
assign c6323 =  x38 &  x41 &  x42 &  x45 &  x70 &  x73 &  x95 &  x96 &  x97 &  x124 &  x125 &  x126 &  x127 &  x129 &  x130 &  x152 &  x154 &  x156 &  x158 &  x183 &  x262 &  x264 &  x266 &  x348 &  x374 &  x432 &  x435 &  x436 &  x437 &  x438 &  x459 &  x486 &  x515 &  x516 &  x541 &  x548 &  x549 &  x597 &  x598 &  x605 &  x660 &  x662 &  x682 &  x709 &  x710 &  x712 &  x716 & ~x24 & ~x28 & ~x58 & ~x60 & ~x84 & ~x114 & ~x142 & ~x167 & ~x198 & ~x224 & ~x225 & ~x279 & ~x305 & ~x310 & ~x336 & ~x338 & ~x364 & ~x366 & ~x367 & ~x418 & ~x423 & ~x446 & ~x450 & ~x451 & ~x477 & ~x502 & ~x507 & ~x529 & ~x557 & ~x586 & ~x646 & ~x671 & ~x698 & ~x702 & ~x703 & ~x727 & ~x753 & ~x754 & ~x780;
assign c6325 =  x758;
assign c6327 =  x475;
assign c6329 = ~x190 & ~x216 & ~x218 & ~x243 & ~x244;
assign c6331 =  x783;
assign c6333 =  x82;
assign c6335 = ~x0 & ~x1 & ~x4 & ~x5 & ~x9 & ~x11 & ~x29 & ~x35 & ~x56 & ~x65 & ~x90 & ~x92 & ~x93 & ~x111 & ~x115 & ~x118 & ~x119 & ~x138 & ~x145 & ~x169 & ~x170 & ~x201 & ~x227 & ~x228 & ~x229 & ~x254 & ~x366 & ~x392 & ~x393 & ~x475 & ~x476 & ~x504 & ~x559 & ~x758 & ~x775 & ~x782 & ~x783;
assign c6337 =  x590;
assign c6339 =  x14 &  x433 &  x455 &  x492 &  x541 &  x549 &  x550 &  x606 & ~x58 & ~x91 & ~x110 & ~x249 & ~x780;
assign c6341 =  x180 &  x235 & ~x7 & ~x22 & ~x36 & ~x60 & ~x85 & ~x192 & ~x197 & ~x199 & ~x221 & ~x250 & ~x255 & ~x282 & ~x309 & ~x361 & ~x393 & ~x394 & ~x422 & ~x478 & ~x506 & ~x557 & ~x590 & ~x636 & ~x699;
assign c6343 =  x190 &  x620 &  x732;
assign c6345 = ~x70 & ~x93;
assign c6347 =  x477;
assign c6349 =  x2;
assign c6351 =  x139;
assign c6353 =  x259 &  x722 &  x733 & ~x3 & ~x5 & ~x6 & ~x7 & ~x22 & ~x24 & ~x28 & ~x29 & ~x50 & ~x53 & ~x56 & ~x57 & ~x80 & ~x85 & ~x88 & ~x108 & ~x112 & ~x114 & ~x136 & ~x141 & ~x164 & ~x168 & ~x170 & ~x195 & ~x198 & ~x220 & ~x221 & ~x222 & ~x223 & ~x224 & ~x227 & ~x248 & ~x253 & ~x255 & ~x276 & ~x277 & ~x278 & ~x280 & ~x281 & ~x304 & ~x305 & ~x308 & ~x310 & ~x332 & ~x360 & ~x361 & ~x362 & ~x363 & ~x366 & ~x388 & ~x390 & ~x391 & ~x394 & ~x417 & ~x419 & ~x421 & ~x422 & ~x445 & ~x449 & ~x450 & ~x473 & ~x478 & ~x502 & ~x503 & ~x504 & ~x506 & ~x530 & ~x531 & ~x532 & ~x534 & ~x557 & ~x559 & ~x585 & ~x589 & ~x614 & ~x615 & ~x617 & ~x641 & ~x642 & ~x645 & ~x669 & ~x670 & ~x673 & ~x697 & ~x700 & ~x701 & ~x726 & ~x729 & ~x730 & ~x731 & ~x739 & ~x740 & ~x741 & ~x742 & ~x743 & ~x747 & ~x753 & ~x755 & ~x757 & ~x764 & ~x766 & ~x769 & ~x770 & ~x771 & ~x774 & ~x782 & ~x783;
assign c6355 =  x120 &  x150 &  x189 &  x217 &  x292 &  x324 &  x377 &  x410 &  x426 &  x429 &  x435 &  x459 &  x486 &  x538 &  x550 &  x566 & ~x4 & ~x19 & ~x56 & ~x60 & ~x61 & ~x137 & ~x138 & ~x165 & ~x223 & ~x224 & ~x281 & ~x305 & ~x337 & ~x339 & ~x449 & ~x450 & ~x560 & ~x590 & ~x702 & ~x730 & ~x741 & ~x776;
assign c6357 =  x82;
assign c6359 = ~x67 & ~x103 & ~x132 & ~x155 & ~x160;
assign c6361 =  x736 &  x766 &  x776;
assign c6363 =  x448;
assign c6365 =  x70 &  x99 &  x150 &  x156 &  x158 &  x177 &  x181 &  x210 &  x211 &  x233 &  x237 &  x272 &  x377 &  x404 &  x430 &  x436 &  x438 &  x462 &  x464 &  x465 &  x487 &  x519 &  x573 &  x603 & ~x9 & ~x18 & ~x58 & ~x64 & ~x78 & ~x81 & ~x85 & ~x86 & ~x87 & ~x135 & ~x163 & ~x166 & ~x196 & ~x226 & ~x254 & ~x255 & ~x308 & ~x334 & ~x335 & ~x419 & ~x422 & ~x560 & ~x673 & ~x726 & ~x727 & ~x783;
assign c6367 =  x83;
assign c6369 = ~x5 & ~x25 & ~x28 & ~x82 & ~x86 & ~x115 & ~x145 & ~x203 & ~x204 & ~x225 & ~x229 & ~x231 & ~x232 & ~x280 & ~x504 & ~x616 & ~x729;
assign c6371 =  x613;
assign c6373 =  x351 &  x491 &  x515 &  x519 &  x521 &  x544 &  x598 &  x605 &  x687 &  x711 &  x738 &  x744 &  x745 & ~x4 & ~x6 & ~x7 & ~x30 & ~x56 & ~x86 & ~x87 & ~x109 & ~x196 & ~x307 & ~x360 & ~x362 & ~x363 & ~x369 & ~x416 & ~x419 & ~x449 & ~x479 & ~x481 & ~x499 & ~x506 & ~x558 & ~x564 & ~x586 & ~x592 & ~x638 & ~x643 & ~x672 & ~x673 & ~x694 & ~x696 & ~x721 & ~x723 & ~x725 & ~x730 & ~x733;
assign c6375 =  x124 &  x127 &  x238 &  x244 &  x352 &  x354 &  x374 &  x435 &  x438 &  x510 &  x547 &  x550 &  x574 &  x576 & ~x9 & ~x88 & ~x114 & ~x137 & ~x167 & ~x277 & ~x308 & ~x338 & ~x360 & ~x451 & ~x472 & ~x506 & ~x640 & ~x668 & ~x670 & ~x675;
assign c6377 = ~x406 & ~x409;
assign c6379 =  x193;
assign c6381 =  x24;
assign c6383 =  x155 &  x370 &  x381 &  x438 &  x459 &  x463 &  x483 &  x520 &  x523 & ~x78 & ~x90 & ~x105 & ~x110 & ~x114 & ~x220 & ~x389;
assign c6385 =  x51 &  x756;
assign c6387 = ~x92 & ~x174 & ~x635 & ~x691 & ~x747;
assign c6389 =  x755;
assign c6391 =  x101 &  x119 &  x122 &  x131 &  x132 &  x134 &  x162 &  x173 &  x176 &  x189 &  x204 &  x219 &  x232 &  x264 &  x290 &  x409 &  x430 &  x432 &  x439 &  x518 &  x522 &  x545 &  x548 &  x550 &  x577 &  x602 &  x603 &  x625 &  x628 &  x655 &  x660 &  x663 &  x681 &  x691 & ~x6 & ~x8 & ~x55 & ~x85 & ~x86 & ~x112 & ~x137 & ~x196 & ~x222 & ~x225 & ~x282 & ~x305 & ~x504 & ~x559 & ~x586 & ~x588 & ~x589 & ~x642 & ~x670 & ~x671 & ~x730 & ~x754 & ~x756;
assign c6393 =  x40 &  x42 &  x70 &  x174 &  x201 &  x229 & ~x20 & ~x530 & ~x767;
assign c6395 =  x11 &  x16 &  x41 & ~x304 & ~x529 & ~x641 & ~x673 & ~x731 & ~x771 & ~x772;
assign c6397 =  x29;
assign c6399 =  x389;
assign c6401 = ~x18 & ~x19 & ~x28 & ~x30 & ~x34 & ~x51 & ~x81 & ~x83 & ~x107 & ~x112 & ~x135 & ~x199 & ~x251 & ~x366 & ~x588 & ~x645 & ~x673 & ~x686 & ~x687 & ~x697 & ~x703 & ~x712 & ~x713 & ~x724 & ~x725 & ~x728 & ~x742 & ~x744 & ~x768 & ~x770;
assign c6403 =  x93 &  x201 &  x481 &  x542 &  x733 & ~x447 & ~x557 & ~x670 & ~x737;
assign c6405 = ~x90 & ~x91 & ~x117 & ~x146 & ~x228 & ~x283 & ~x317;
assign c6407 =  x75 &  x76 &  x163 &  x173 &  x625 &  x681;
assign c6409 =  x13 &  x14 &  x122 &  x124 &  x125 &  x149 &  x150 &  x155 &  x156 &  x184 &  x240 & ~x0 & ~x24 & ~x26 & ~x29 & ~x34 & ~x50 & ~x79 & ~x90 & ~x105 & ~x109 & ~x135 & ~x199 & ~x224 & ~x255 & ~x334 & ~x389 & ~x503 & ~x617 & ~x729;
assign c6411 = ~x9 & ~x60 & ~x105 & ~x172 & ~x200 & ~x367 & ~x593 & ~x594 & ~x636 & ~x666 & ~x692 & ~x695 & ~x706 & ~x731 & ~x754;
assign c6413 =  x181 &  x401 &  x542 &  x575 &  x577 &  x625 &  x634 &  x663 &  x682 &  x687 &  x711 &  x712 &  x748 & ~x53 & ~x85 & ~x138 & ~x482 & ~x497 & ~x588 & ~x610;
assign c6415 =  x483 &  x599 & ~x29 & ~x33 & ~x47 & ~x90 & ~x104 & ~x105 & ~x106 & ~x107 & ~x110 & ~x117 & ~x135 & ~x225 & ~x280 & ~x615 & ~x781;
assign c6417 =  x401 &  x428 &  x439 &  x453 &  x568 &  x606 &  x625 &  x721 & ~x226 & ~x305 & ~x753;
assign c6419 =  x29;
assign c6423 =  x41 &  x43 &  x105 &  x228 &  x288 &  x402 &  x570 &  x712 & ~x33 & ~x142 & ~x198 & ~x337 & ~x417 & ~x449 & ~x502 & ~x504 & ~x645 & ~x698 & ~x757;
assign c6425 =  x39 &  x44 &  x69 &  x70 &  x96 &  x97 &  x98 &  x100 &  x102 &  x132 &  x147 &  x148 &  x149 &  x161 &  x177 &  x181 &  x184 &  x189 &  x190 &  x202 &  x205 &  x211 &  x212 &  x213 &  x241 &  x245 &  x257 &  x264 &  x272 &  x285 &  x287 &  x290 &  x319 &  x373 &  x376 &  x378 &  x381 &  x383 &  x405 &  x410 &  x411 &  x429 &  x431 &  x435 &  x437 &  x459 &  x460 &  x466 &  x488 &  x489 &  x516 &  x521 &  x543 &  x544 &  x548 &  x579 &  x597 &  x598 &  x602 &  x605 &  x606 &  x627 &  x629 &  x658 &  x662 & ~x1 & ~x3 & ~x6 & ~x27 & ~x51 & ~x57 & ~x59 & ~x110 & ~x137 & ~x193 & ~x195 & ~x249 & ~x251 & ~x282 & ~x306 & ~x335 & ~x338 & ~x389 & ~x392 & ~x417 & ~x420 & ~x445 & ~x446 & ~x478 & ~x557 & ~x559 & ~x561 & ~x585 & ~x588 & ~x613 & ~x615 & ~x616 & ~x641 & ~x644 & ~x669 & ~x671 & ~x697 & ~x699 & ~x702 & ~x730 & ~x754;
assign c6427 =  x243 &  x273 &  x343 &  x344 &  x381 &  x414 &  x427 &  x489 &  x512 &  x519 &  x520 &  x554 &  x567 &  x568 & ~x63 & ~x79 & ~x531;
assign c6429 =  x475;
assign c6433 =  x336;
assign c6435 =  x584 &  x640 &  x708;
assign c6437 =  x57;
assign c6439 =  x783;
assign c6441 =  x497 &  x511 & ~x24 & ~x63 & ~x77 & ~x106 & ~x738 & ~x740 & ~x744 & ~x759 & ~x768 & ~x770;
assign c6443 =  x195;
assign c6447 =  x660 &  x766 & ~x371;
assign c6449 = ~x91 & ~x98 & ~x147 & ~x181 & ~x205;
assign c6451 =  x420;
assign c6453 =  x462 &  x511 & ~x37 & ~x48 & ~x64 & ~x76 & ~x92;
assign c6455 =  x224;
assign c6457 =  x69 &  x120 &  x126 &  x151 &  x153 &  x156 &  x161 &  x175 &  x177 &  x180 &  x183 &  x184 &  x185 &  x188 &  x203 &  x209 &  x210 &  x216 &  x239 &  x263 &  x270 &  x301 &  x322 &  x346 &  x347 &  x351 &  x380 &  x385 &  x386 &  x403 &  x404 &  x425 &  x426 &  x427 &  x432 &  x461 &  x470 &  x494 &  x519 &  x526 &  x549 &  x638 & ~x28 & ~x31 & ~x51 & ~x53 & ~x54 & ~x88 & ~x113 & ~x114 & ~x136 & ~x137 & ~x138 & ~x170 & ~x171 & ~x192 & ~x193 & ~x194 & ~x222 & ~x223 & ~x249 & ~x308 & ~x361 & ~x393 & ~x418 & ~x419 & ~x445 & ~x476 & ~x477 & ~x504 & ~x505 & ~x506 & ~x531 & ~x534 & ~x557 & ~x558 & ~x560 & ~x589 & ~x615 & ~x618 & ~x641 & ~x642 & ~x669 & ~x672 & ~x725 & ~x758 & ~x764 & ~x765 & ~x766 & ~x767 & ~x768 & ~x769 & ~x772 & ~x776;
assign c6459 =  x56;
assign c6461 =  x427 &  x494 &  x511 &  x520 &  x525 &  x567 &  x581 & ~x55 & ~x91 & ~x118 & ~x532;
assign c6463 = ~x8 & ~x26 & ~x34 & ~x87 & ~x108 & ~x193 & ~x194 & ~x279 & ~x312 & ~x337 & ~x340 & ~x420 & ~x442 & ~x535 & ~x536 & ~x553 & ~x566 & ~x583 & ~x591 & ~x594 & ~x608 & ~x638 & ~x639 & ~x694 & ~x701 & ~x724 & ~x749 & ~x750 & ~x777 & ~x780;
assign c6465 =  x279;
assign c6467 =  x83;
assign c6469 =  x113;
assign c6471 = ~x15 & ~x35 & ~x90 & ~x176 & ~x201 & ~x205;
assign c6473 =  x39 &  x45 &  x231 &  x240 &  x431 &  x441 &  x442 &  x469 &  x497 &  x526 &  x547 &  x625 & ~x53 & ~x55 & ~x114 & ~x137 & ~x171 & ~x196 & ~x309 & ~x311 & ~x333 & ~x361 & ~x446 & ~x501 & ~x558 & ~x647 & ~x730;
assign c6475 =  x215 &  x316 & ~x64 & ~x733 & ~x734 & ~x762;
assign c6477 =  x504;
assign c6479 = ~x5 & ~x19 & ~x37 & ~x58 & ~x65 & ~x93 & ~x134 & ~x196 & ~x229 & ~x280 & ~x504 & ~x671 & ~x760;
assign c6481 =  x232 &  x259 &  x323 &  x402 &  x516 &  x548 &  x569 &  x579 &  x628 &  x634 &  x656 &  x658 &  x683 &  x685 &  x713 &  x736 &  x738 &  x743 & ~x59 & ~x138 & ~x222 & ~x253 & ~x364 & ~x394 & ~x421 & ~x449 & ~x501 & ~x502 & ~x585 & ~x614 & ~x647 & ~x649 & ~x667 & ~x678 & ~x697 & ~x703 & ~x723 & ~x779 & ~x781;
assign c6483 =  x39 &  x69 &  x71 &  x93 &  x119 &  x123 &  x124 &  x126 &  x127 &  x151 &  x154 &  x162 &  x219 &  x257 &  x378 &  x383 &  x485 &  x541 &  x547 &  x572 &  x628 &  x634 &  x654 &  x661 &  x662 &  x688 &  x709 &  x714 &  x719 & ~x7 & ~x20 & ~x55 & ~x111 & ~x113 & ~x140 & ~x166 & ~x167 & ~x222 & ~x252 & ~x253 & ~x279 & ~x280 & ~x337 & ~x419 & ~x448 & ~x504 & ~x505 & ~x558 & ~x586 & ~x614 & ~x617 & ~x670 & ~x700 & ~x757 & ~x759 & ~x783;
assign c6485 =  x308;
assign c6487 =  x55;
assign c6489 =  x39 &  x40 &  x150 &  x177 &  x259 &  x291 &  x377 &  x431 &  x520 &  x543 &  x576 &  x600 &  x716 &  x717 &  x737 &  x740 &  x743 & ~x8 & ~x24 & ~x27 & ~x28 & ~x80 & ~x81 & ~x168 & ~x282 & ~x361 & ~x393 & ~x472 & ~x557 & ~x587 & ~x645 & ~x734 & ~x762 & ~x778;
assign c6491 = ~x10 & ~x14 & ~x15 & ~x28 & ~x31 & ~x33 & ~x281 & ~x283 & ~x286 & ~x313 & ~x315 & ~x342 & ~x775;
assign c6493 =  x21;
assign c6495 =  x176 &  x287 &  x514 &  x522 &  x550 &  x578 &  x599 &  x627 &  x661 &  x662 &  x710 &  x716 & ~x30 & ~x32 & ~x50 & ~x58 & ~x168 & ~x193 & ~x335 & ~x337 & ~x363 & ~x390 & ~x393 & ~x417 & ~x444 & ~x449 & ~x472 & ~x479 & ~x535 & ~x561 & ~x563 & ~x587 & ~x612 & ~x614 & ~x668 & ~x670 & ~x675 & ~x698 & ~x700 & ~x705 & ~x706 & ~x721 & ~x726 & ~x734 & ~x762;
assign c6497 =  x515 & ~x75 & ~x104 & ~x118 & ~x119;
assign c70 =  x185 &  x324 &  x333 &  x429 & ~x0 & ~x7 & ~x9 & ~x10 & ~x23 & ~x40 & ~x48 & ~x52 & ~x55 & ~x65 & ~x88 & ~x89 & ~x110 & ~x111 & ~x115 & ~x134 & ~x137 & ~x139 & ~x172 & ~x177 & ~x256 & ~x281 & ~x282 & ~x283 & ~x288 & ~x337 & ~x531 & ~x705 & ~x723 & ~x730 & ~x748 & ~x749 & ~x761 & ~x762 & ~x764 & ~x776 & ~x780;
assign c72 =  x691;
assign c74 = ~x8 & ~x10 & ~x13 & ~x15 & ~x16 & ~x18 & ~x22 & ~x27 & ~x29 & ~x33 & ~x37 & ~x39 & ~x40 & ~x43 & ~x53 & ~x54 & ~x64 & ~x67 & ~x71 & ~x76 & ~x79 & ~x80 & ~x84 & ~x94 & ~x98 & ~x100 & ~x103 & ~x110 & ~x111 & ~x112 & ~x116 & ~x126 & ~x127 & ~x128 & ~x130 & ~x131 & ~x134 & ~x139 & ~x147 & ~x157 & ~x163 & ~x164 & ~x178 & ~x179 & ~x180 & ~x188 & ~x192 & ~x197 & ~x202 & ~x204 & ~x206 & ~x207 & ~x209 & ~x220 & ~x226 & ~x228 & ~x245 & ~x253 & ~x254 & ~x264 & ~x272 & ~x274 & ~x281 & ~x289 & ~x291 & ~x300 & ~x310 & ~x312 & ~x315 & ~x317 & ~x318 & ~x328 & ~x329 & ~x337 & ~x338 & ~x341 & ~x342 & ~x343 & ~x345 & ~x367 & ~x368 & ~x392 & ~x588 & ~x589 & ~x649 & ~x656 & ~x661 & ~x667 & ~x668 & ~x678 & ~x682 & ~x691 & ~x692 & ~x705 & ~x712 & ~x713 & ~x719 & ~x720 & ~x721 & ~x730 & ~x733 & ~x740 & ~x742 & ~x758 & ~x771 & ~x779 & ~x780;
assign c76 =  x276 & ~x0 & ~x4 & ~x9 & ~x12 & ~x13 & ~x14 & ~x15 & ~x16 & ~x21 & ~x23 & ~x28 & ~x37 & ~x38 & ~x42 & ~x47 & ~x57 & ~x60 & ~x61 & ~x62 & ~x80 & ~x85 & ~x90 & ~x108 & ~x119 & ~x138 & ~x139 & ~x141 & ~x149 & ~x150 & ~x151 & ~x171 & ~x174 & ~x178 & ~x196 & ~x199 & ~x202 & ~x206 & ~x209 & ~x230 & ~x231 & ~x252 & ~x284 & ~x309 & ~x314 & ~x315 & ~x339 & ~x476 & ~x558 & ~x584 & ~x585 & ~x608 & ~x611 & ~x612 & ~x613 & ~x616 & ~x640 & ~x641 & ~x643 & ~x644 & ~x664 & ~x688 & ~x693 & ~x694 & ~x697 & ~x700 & ~x714 & ~x715 & ~x727 & ~x746 & ~x754 & ~x760 & ~x764 & ~x767 & ~x773 & ~x775 & ~x778 & ~x780 & ~x783;
assign c78 =  x351 &  x445 & ~x7 & ~x9 & ~x10 & ~x13 & ~x16 & ~x17 & ~x22 & ~x23 & ~x31 & ~x32 & ~x35 & ~x36 & ~x41 & ~x43 & ~x44 & ~x48 & ~x52 & ~x58 & ~x67 & ~x70 & ~x73 & ~x74 & ~x75 & ~x76 & ~x77 & ~x79 & ~x85 & ~x86 & ~x91 & ~x96 & ~x97 & ~x99 & ~x104 & ~x106 & ~x109 & ~x111 & ~x112 & ~x128 & ~x129 & ~x137 & ~x138 & ~x139 & ~x140 & ~x141 & ~x143 & ~x147 & ~x150 & ~x151 & ~x167 & ~x172 & ~x174 & ~x179 & ~x191 & ~x193 & ~x201 & ~x205 & ~x217 & ~x220 & ~x225 & ~x227 & ~x229 & ~x230 & ~x249 & ~x255 & ~x256 & ~x284 & ~x285 & ~x286 & ~x311 & ~x315 & ~x339 & ~x342 & ~x365 & ~x391 & ~x393 & ~x397 & ~x419 & ~x588 & ~x646 & ~x674 & ~x676 & ~x677 & ~x684 & ~x692 & ~x698 & ~x702 & ~x707 & ~x714 & ~x718 & ~x727 & ~x729 & ~x737 & ~x739 & ~x747 & ~x755 & ~x758 & ~x763 & ~x765 & ~x768 & ~x772 & ~x777 & ~x779;
assign c710 =  x215 & ~x5 & ~x7 & ~x11 & ~x22 & ~x24 & ~x31 & ~x37 & ~x43 & ~x46 & ~x47 & ~x48 & ~x75 & ~x77 & ~x86 & ~x87 & ~x90 & ~x91 & ~x94 & ~x101 & ~x105 & ~x113 & ~x116 & ~x120 & ~x122 & ~x123 & ~x125 & ~x129 & ~x139 & ~x147 & ~x149 & ~x151 & ~x166 & ~x168 & ~x174 & ~x181 & ~x192 & ~x194 & ~x199 & ~x200 & ~x202 & ~x210 & ~x219 & ~x224 & ~x230 & ~x251 & ~x259 & ~x263 & ~x265 & ~x283 & ~x284 & ~x286 & ~x311 & ~x316 & ~x337 & ~x338 & ~x365 & ~x366 & ~x392 & ~x394 & ~x424 & ~x692 & ~x696 & ~x698 & ~x704 & ~x706 & ~x708 & ~x711 & ~x716 & ~x717 & ~x718 & ~x725 & ~x728 & ~x735 & ~x741 & ~x743 & ~x747 & ~x753 & ~x760 & ~x761 & ~x762 & ~x763 & ~x769 & ~x780;
assign c712 =  x324 &  x428 &  x457 &  x458 & ~x10 & ~x13 & ~x17 & ~x26 & ~x27 & ~x30 & ~x36 & ~x45 & ~x51 & ~x53 & ~x54 & ~x63 & ~x66 & ~x67 & ~x72 & ~x77 & ~x81 & ~x84 & ~x85 & ~x96 & ~x115 & ~x123 & ~x124 & ~x126 & ~x137 & ~x140 & ~x142 & ~x144 & ~x145 & ~x153 & ~x159 & ~x161 & ~x166 & ~x174 & ~x176 & ~x189 & ~x190 & ~x194 & ~x197 & ~x198 & ~x205 & ~x207 & ~x231 & ~x252 & ~x261 & ~x266 & ~x281 & ~x288 & ~x315 & ~x335 & ~x337 & ~x341 & ~x363 & ~x364 & ~x392 & ~x560 & ~x588 & ~x590 & ~x615 & ~x620 & ~x621 & ~x639 & ~x646 & ~x649 & ~x655 & ~x657 & ~x659 & ~x660 & ~x661 & ~x663 & ~x668 & ~x673 & ~x675 & ~x677 & ~x681 & ~x683 & ~x685 & ~x688 & ~x704 & ~x718 & ~x728 & ~x729 & ~x733 & ~x740 & ~x751 & ~x752 & ~x753 & ~x759 & ~x760 & ~x771 & ~x773 & ~x776 & ~x780;
assign c714 =  x423 &  x449 & ~x6 & ~x14 & ~x15 & ~x19 & ~x36 & ~x45 & ~x48 & ~x50 & ~x51 & ~x74 & ~x78 & ~x83 & ~x89 & ~x91 & ~x96 & ~x99 & ~x102 & ~x105 & ~x106 & ~x107 & ~x124 & ~x127 & ~x135 & ~x136 & ~x139 & ~x140 & ~x143 & ~x154 & ~x162 & ~x163 & ~x176 & ~x177 & ~x181 & ~x182 & ~x188 & ~x190 & ~x198 & ~x199 & ~x209 & ~x212 & ~x217 & ~x220 & ~x232 & ~x238 & ~x254 & ~x259 & ~x281 & ~x282 & ~x284 & ~x288 & ~x308 & ~x312 & ~x313 & ~x315 & ~x369 & ~x560 & ~x618 & ~x622 & ~x628 & ~x629 & ~x631 & ~x634 & ~x639 & ~x640 & ~x653 & ~x658 & ~x662 & ~x667 & ~x669 & ~x672 & ~x674 & ~x681 & ~x686 & ~x691 & ~x693 & ~x701 & ~x705 & ~x713 & ~x720 & ~x724 & ~x729 & ~x731 & ~x736 & ~x738 & ~x741 & ~x751 & ~x752 & ~x762 & ~x763 & ~x765 & ~x766;
assign c716 =  x355 &  x362 &  x409 &  x418 & ~x0 & ~x5 & ~x7 & ~x12 & ~x19 & ~x24 & ~x25 & ~x26 & ~x27 & ~x38 & ~x39 & ~x44 & ~x46 & ~x50 & ~x59 & ~x63 & ~x65 & ~x70 & ~x73 & ~x74 & ~x75 & ~x81 & ~x84 & ~x86 & ~x94 & ~x99 & ~x103 & ~x104 & ~x105 & ~x127 & ~x130 & ~x134 & ~x144 & ~x151 & ~x152 & ~x161 & ~x165 & ~x173 & ~x174 & ~x197 & ~x200 & ~x202 & ~x223 & ~x226 & ~x234 & ~x251 & ~x255 & ~x260 & ~x284 & ~x285 & ~x581 & ~x586 & ~x600 & ~x620 & ~x645 & ~x647 & ~x654 & ~x659 & ~x666 & ~x670 & ~x672 & ~x676 & ~x680 & ~x685 & ~x686 & ~x691 & ~x694 & ~x695 & ~x700 & ~x703 & ~x705 & ~x707 & ~x709 & ~x717 & ~x720 & ~x721 & ~x725 & ~x726 & ~x729 & ~x732 & ~x746 & ~x749 & ~x752 & ~x762 & ~x764 & ~x771 & ~x774 & ~x778;
assign c718 =  x359 &  x406 &  x407 &  x458 &  x467 &  x468 &  x471 &  x472 &  x511 &  x516 & ~x0 & ~x8 & ~x9 & ~x16 & ~x23 & ~x26 & ~x35 & ~x41 & ~x47 & ~x49 & ~x54 & ~x66 & ~x69 & ~x83 & ~x85 & ~x92 & ~x93 & ~x98 & ~x102 & ~x105 & ~x107 & ~x109 & ~x111 & ~x115 & ~x121 & ~x143 & ~x149 & ~x182 & ~x192 & ~x194 & ~x207 & ~x222 & ~x233 & ~x234 & ~x238 & ~x256 & ~x261 & ~x265 & ~x266 & ~x284 & ~x285 & ~x286 & ~x308 & ~x313 & ~x338 & ~x342 & ~x668 & ~x669 & ~x670 & ~x673 & ~x679 & ~x684 & ~x685 & ~x686 & ~x689 & ~x690 & ~x706 & ~x718 & ~x726 & ~x727 & ~x731 & ~x745 & ~x751 & ~x762 & ~x766 & ~x770 & ~x773 & ~x780;
assign c720 = ~x6 & ~x17 & ~x22 & ~x24 & ~x25 & ~x27 & ~x28 & ~x30 & ~x31 & ~x35 & ~x36 & ~x39 & ~x40 & ~x41 & ~x42 & ~x43 & ~x44 & ~x54 & ~x66 & ~x68 & ~x84 & ~x86 & ~x87 & ~x88 & ~x90 & ~x91 & ~x98 & ~x100 & ~x102 & ~x108 & ~x109 & ~x114 & ~x118 & ~x119 & ~x120 & ~x122 & ~x123 & ~x125 & ~x126 & ~x129 & ~x134 & ~x136 & ~x140 & ~x143 & ~x145 & ~x148 & ~x151 & ~x152 & ~x169 & ~x180 & ~x183 & ~x192 & ~x198 & ~x203 & ~x204 & ~x207 & ~x223 & ~x233 & ~x245 & ~x251 & ~x257 & ~x272 & ~x279 & ~x284 & ~x301 & ~x308 & ~x312 & ~x337 & ~x364 & ~x412 & ~x611 & ~x613 & ~x615 & ~x640 & ~x642 & ~x643 & ~x662 & ~x663 & ~x664 & ~x667 & ~x669 & ~x679 & ~x681 & ~x689 & ~x695 & ~x697 & ~x699 & ~x713 & ~x718 & ~x721 & ~x722 & ~x724 & ~x730 & ~x742 & ~x743 & ~x744 & ~x747 & ~x748 & ~x749 & ~x752 & ~x758 & ~x761 & ~x763 & ~x769 & ~x772 & ~x775 & ~x783;
assign c722 =  x460 &  x487 &  x489 &  x513 & ~x4 & ~x71 & ~x116 & ~x132 & ~x179 & ~x189 & ~x193 & ~x195 & ~x450 & ~x749 & ~x757;
assign c724 = ~x18 & ~x46 & ~x64 & ~x104 & ~x131 & ~x133 & ~x148 & ~x169 & ~x452 & ~x483 & ~x512 & ~x652 & ~x686 & ~x709 & ~x731 & ~x733 & ~x744 & ~x777;
assign c726 =  x362 &  x443 &  x471 &  x473 &  x484 & ~x10 & ~x22 & ~x44 & ~x48 & ~x92 & ~x204 & ~x206 & ~x232 & ~x314 & ~x477 & ~x700 & ~x756 & ~x765 & ~x766;
assign c728 =  x158 &  x472 & ~x24 & ~x36 & ~x42 & ~x43 & ~x63 & ~x113 & ~x116 & ~x120 & ~x139 & ~x146 & ~x150 & ~x169 & ~x336 & ~x338 & ~x393 & ~x724 & ~x746 & ~x752 & ~x766 & ~x772 & ~x778;
assign c730 =  x418 &  x449 & ~x2 & ~x5 & ~x6 & ~x7 & ~x9 & ~x40 & ~x42 & ~x55 & ~x60 & ~x79 & ~x85 & ~x97 & ~x100 & ~x118 & ~x124 & ~x127 & ~x135 & ~x136 & ~x142 & ~x151 & ~x162 & ~x164 & ~x165 & ~x169 & ~x175 & ~x176 & ~x181 & ~x183 & ~x195 & ~x201 & ~x204 & ~x244 & ~x251 & ~x254 & ~x300 & ~x336 & ~x595 & ~x598 & ~x609 & ~x610 & ~x613 & ~x627 & ~x634 & ~x637 & ~x651 & ~x654 & ~x661 & ~x666 & ~x667 & ~x676 & ~x679 & ~x680 & ~x683 & ~x686 & ~x688 & ~x691 & ~x704 & ~x705 & ~x708 & ~x711 & ~x713 & ~x718 & ~x719 & ~x742 & ~x750 & ~x772 & ~x783;
assign c732 =  x330 &  x524 &  x660 & ~x397 & ~x425;
assign c734 =  x215 & ~x3 & ~x5 & ~x6 & ~x11 & ~x17 & ~x28 & ~x29 & ~x30 & ~x32 & ~x33 & ~x36 & ~x38 & ~x49 & ~x52 & ~x59 & ~x70 & ~x80 & ~x81 & ~x83 & ~x89 & ~x101 & ~x124 & ~x128 & ~x132 & ~x149 & ~x155 & ~x178 & ~x179 & ~x230 & ~x237 & ~x256 & ~x260 & ~x261 & ~x282 & ~x283 & ~x310 & ~x336 & ~x339 & ~x340 & ~x365 & ~x369 & ~x395 & ~x419 & ~x425 & ~x449 & ~x450 & ~x644 & ~x661 & ~x667 & ~x680 & ~x691 & ~x714 & ~x715 & ~x717 & ~x721 & ~x729 & ~x730 & ~x736 & ~x742 & ~x745 & ~x748 & ~x753 & ~x757 & ~x763 & ~x774;
assign c736 =  x158 &  x185 &  x446 & ~x5 & ~x109;
assign c738 =  x457 &  x576 & ~x24 & ~x34 & ~x63 & ~x66 & ~x89 & ~x95 & ~x98 & ~x124 & ~x127 & ~x133 & ~x166 & ~x183 & ~x193 & ~x224 & ~x238 & ~x253 & ~x257 & ~x281 & ~x311 & ~x338 & ~x618 & ~x619 & ~x635 & ~x636 & ~x643 & ~x647 & ~x650 & ~x680 & ~x686 & ~x689 & ~x731 & ~x732 & ~x734 & ~x739 & ~x744 & ~x755;
assign c740 =  x489 & ~x17 & ~x23 & ~x100 & ~x106 & ~x119 & ~x122 & ~x143 & ~x179 & ~x196 & ~x203 & ~x223 & ~x290 & ~x291 & ~x295 & ~x337 & ~x365 & ~x371 & ~x736 & ~x755 & ~x776;
assign c742 =  x381 &  x558 &  x662 & ~x105 & ~x290 & ~x450 & ~x453;
assign c744 =  x389 & ~x9 & ~x10 & ~x14 & ~x17 & ~x18 & ~x19 & ~x20 & ~x26 & ~x35 & ~x37 & ~x38 & ~x40 & ~x41 & ~x55 & ~x57 & ~x59 & ~x60 & ~x66 & ~x69 & ~x83 & ~x89 & ~x90 & ~x106 & ~x112 & ~x137 & ~x146 & ~x147 & ~x160 & ~x169 & ~x170 & ~x178 & ~x198 & ~x200 & ~x202 & ~x208 & ~x209 & ~x210 & ~x223 & ~x234 & ~x257 & ~x282 & ~x313 & ~x501 & ~x645 & ~x662 & ~x667 & ~x670 & ~x686 & ~x691 & ~x693 & ~x696 & ~x704 & ~x708 & ~x712 & ~x714 & ~x736 & ~x743 & ~x750 & ~x755 & ~x771 & ~x772 & ~x778;
assign c746 =  x499 &  x632 & ~x40 & ~x150 & ~x205 & ~x279 & ~x336 & ~x752 & ~x776;
assign c748 =  x322 &  x418 &  x446 &  x526 &  x631 & ~x335 & ~x369;
assign c750 =  x277 &  x383 &  x446 & ~x4 & ~x5 & ~x6 & ~x7 & ~x11 & ~x12 & ~x14 & ~x18 & ~x19 & ~x20 & ~x22 & ~x24 & ~x25 & ~x28 & ~x31 & ~x32 & ~x36 & ~x38 & ~x47 & ~x53 & ~x54 & ~x57 & ~x58 & ~x62 & ~x82 & ~x89 & ~x90 & ~x91 & ~x93 & ~x94 & ~x114 & ~x121 & ~x122 & ~x143 & ~x144 & ~x148 & ~x149 & ~x167 & ~x172 & ~x177 & ~x178 & ~x196 & ~x201 & ~x205 & ~x206 & ~x207 & ~x226 & ~x228 & ~x229 & ~x230 & ~x232 & ~x234 & ~x235 & ~x252 & ~x254 & ~x255 & ~x256 & ~x257 & ~x258 & ~x259 & ~x260 & ~x261 & ~x262 & ~x279 & ~x281 & ~x282 & ~x283 & ~x286 & ~x287 & ~x309 & ~x311 & ~x312 & ~x339 & ~x364 & ~x365 & ~x585 & ~x586 & ~x610 & ~x611 & ~x612 & ~x613 & ~x614 & ~x637 & ~x641 & ~x643 & ~x667 & ~x668 & ~x670 & ~x671 & ~x690 & ~x694 & ~x695 & ~x696 & ~x697 & ~x699 & ~x700 & ~x714 & ~x727 & ~x757 & ~x760 & ~x761 & ~x771 & ~x773 & ~x776 & ~x781 & ~x782;
assign c752 =  x576 &  x579 & ~x16 & ~x19 & ~x29 & ~x30 & ~x32 & ~x33 & ~x37 & ~x39 & ~x43 & ~x45 & ~x48 & ~x49 & ~x51 & ~x64 & ~x77 & ~x90 & ~x91 & ~x92 & ~x100 & ~x101 & ~x104 & ~x106 & ~x112 & ~x113 & ~x123 & ~x125 & ~x131 & ~x134 & ~x137 & ~x145 & ~x150 & ~x165 & ~x166 & ~x167 & ~x168 & ~x170 & ~x172 & ~x175 & ~x178 & ~x197 & ~x201 & ~x204 & ~x225 & ~x226 & ~x231 & ~x232 & ~x255 & ~x257 & ~x290 & ~x310 & ~x342 & ~x365 & ~x593 & ~x613 & ~x617 & ~x627 & ~x631 & ~x633 & ~x636 & ~x643 & ~x649 & ~x668 & ~x685 & ~x705 & ~x710 & ~x713 & ~x715 & ~x718 & ~x721 & ~x722 & ~x728 & ~x731 & ~x735 & ~x736 & ~x741 & ~x742 & ~x743 & ~x744 & ~x751 & ~x752 & ~x755 & ~x756 & ~x766 & ~x770 & ~x771 & ~x778 & ~x782;
assign c754 =  x403 &  x411 &  x429 & ~x13 & ~x14 & ~x22 & ~x29 & ~x40 & ~x54 & ~x66 & ~x105 & ~x205 & ~x209 & ~x210 & ~x290 & ~x310 & ~x615 & ~x679 & ~x683 & ~x697 & ~x705 & ~x722 & ~x730 & ~x759 & ~x767;
assign c756 = ~x0 & ~x4 & ~x5 & ~x6 & ~x10 & ~x15 & ~x16 & ~x25 & ~x26 & ~x27 & ~x28 & ~x32 & ~x34 & ~x37 & ~x40 & ~x41 & ~x42 & ~x43 & ~x46 & ~x51 & ~x59 & ~x61 & ~x62 & ~x71 & ~x72 & ~x75 & ~x76 & ~x80 & ~x81 & ~x83 & ~x85 & ~x89 & ~x95 & ~x98 & ~x100 & ~x101 & ~x102 & ~x103 & ~x104 & ~x109 & ~x111 & ~x119 & ~x129 & ~x132 & ~x133 & ~x135 & ~x139 & ~x141 & ~x142 & ~x145 & ~x146 & ~x150 & ~x155 & ~x161 & ~x165 & ~x167 & ~x168 & ~x173 & ~x174 & ~x176 & ~x177 & ~x197 & ~x198 & ~x201 & ~x204 & ~x207 & ~x224 & ~x229 & ~x231 & ~x235 & ~x251 & ~x254 & ~x255 & ~x257 & ~x261 & ~x280 & ~x281 & ~x282 & ~x284 & ~x286 & ~x288 & ~x311 & ~x313 & ~x314 & ~x315 & ~x342 & ~x343 & ~x366 & ~x369 & ~x370 & ~x447 & ~x475 & ~x503 & ~x534 & ~x567 & ~x573 & ~x617 & ~x621 & ~x622 & ~x633 & ~x642 & ~x643 & ~x645 & ~x646 & ~x649 & ~x652 & ~x653 & ~x654 & ~x656 & ~x657 & ~x658 & ~x663 & ~x674 & ~x675 & ~x677 & ~x681 & ~x682 & ~x683 & ~x687 & ~x688 & ~x690 & ~x693 & ~x694 & ~x695 & ~x697 & ~x698 & ~x700 & ~x702 & ~x703 & ~x704 & ~x715 & ~x717 & ~x722 & ~x723 & ~x724 & ~x727 & ~x730 & ~x731 & ~x732 & ~x735 & ~x736 & ~x738 & ~x743 & ~x744 & ~x747 & ~x749 & ~x751 & ~x752 & ~x754 & ~x760 & ~x761 & ~x764 & ~x769 & ~x770 & ~x774 & ~x775 & ~x777 & ~x778 & ~x781 & ~x782;
assign c758 =  x333 &  x462 & ~x25 & ~x38 & ~x41 & ~x48 & ~x56 & ~x94 & ~x112 & ~x120 & ~x143 & ~x144 & ~x163 & ~x164 & ~x165 & ~x227 & ~x245 & ~x251 & ~x254 & ~x308 & ~x310 & ~x327 & ~x335 & ~x337 & ~x644 & ~x655 & ~x666 & ~x669 & ~x693 & ~x696 & ~x713 & ~x757 & ~x760;
assign c760 =  x451 & ~x438;
assign c762 =  x333 &  x362 &  x403 &  x435 &  x502 &  x550 &  x606 & ~x106 & ~x110 & ~x224 & ~x781;
assign c764 =  x330 &  x410 &  x412 & ~x52 & ~x55 & ~x64 & ~x68 & ~x70 & ~x71 & ~x77 & ~x105 & ~x114 & ~x120 & ~x129 & ~x136 & ~x167 & ~x169 & ~x194 & ~x221 & ~x233 & ~x235 & ~x259 & ~x261 & ~x262 & ~x280 & ~x313 & ~x336 & ~x391 & ~x420 & ~x452 & ~x672 & ~x675 & ~x711 & ~x715 & ~x724 & ~x737 & ~x747 & ~x749 & ~x750 & ~x759 & ~x769 & ~x771 & ~x777 & ~x783;
assign c766 =  x430 &  x606 &  x608 & ~x59 & ~x114 & ~x134 & ~x149 & ~x289 & ~x667;
assign c768 = ~x13 & ~x41 & ~x44 & ~x69 & ~x77 & ~x110 & ~x115 & ~x119 & ~x124 & ~x128 & ~x130 & ~x140 & ~x152 & ~x157 & ~x162 & ~x180 & ~x189 & ~x193 & ~x201 & ~x206 & ~x229 & ~x288 & ~x313 & ~x339 & ~x343 & ~x481 & ~x483 & ~x641 & ~x643 & ~x648 & ~x651 & ~x665 & ~x678 & ~x685 & ~x687 & ~x689 & ~x693 & ~x694 & ~x696 & ~x701 & ~x711 & ~x712 & ~x713 & ~x715 & ~x727 & ~x734 & ~x740 & ~x746 & ~x750 & ~x751 & ~x752 & ~x765 & ~x776;
assign c770 =  x578 &  x581 &  x582 &  x583 & ~x3 & ~x17 & ~x24 & ~x25 & ~x28 & ~x29 & ~x33 & ~x35 & ~x36 & ~x39 & ~x43 & ~x46 & ~x63 & ~x64 & ~x68 & ~x71 & ~x72 & ~x91 & ~x96 & ~x97 & ~x103 & ~x114 & ~x117 & ~x119 & ~x120 & ~x123 & ~x124 & ~x131 & ~x138 & ~x139 & ~x143 & ~x150 & ~x151 & ~x153 & ~x159 & ~x173 & ~x174 & ~x176 & ~x198 & ~x202 & ~x220 & ~x223 & ~x224 & ~x226 & ~x229 & ~x230 & ~x254 & ~x256 & ~x261 & ~x279 & ~x280 & ~x287 & ~x307 & ~x309 & ~x314 & ~x364 & ~x595 & ~x615 & ~x616 & ~x638 & ~x648 & ~x650 & ~x677 & ~x678 & ~x680 & ~x681 & ~x685 & ~x690 & ~x692 & ~x693 & ~x696 & ~x698 & ~x700 & ~x705 & ~x710 & ~x714 & ~x715 & ~x722 & ~x728 & ~x749 & ~x753 & ~x761 & ~x775;
assign c772 = ~x0 & ~x3 & ~x7 & ~x12 & ~x16 & ~x20 & ~x28 & ~x30 & ~x32 & ~x36 & ~x60 & ~x61 & ~x63 & ~x66 & ~x70 & ~x71 & ~x76 & ~x78 & ~x79 & ~x80 & ~x82 & ~x83 & ~x89 & ~x92 & ~x97 & ~x98 & ~x99 & ~x106 & ~x107 & ~x108 & ~x110 & ~x112 & ~x113 & ~x114 & ~x122 & ~x127 & ~x129 & ~x130 & ~x133 & ~x144 & ~x148 & ~x152 & ~x154 & ~x161 & ~x162 & ~x164 & ~x166 & ~x169 & ~x174 & ~x175 & ~x179 & ~x181 & ~x182 & ~x183 & ~x187 & ~x189 & ~x198 & ~x199 & ~x201 & ~x205 & ~x206 & ~x208 & ~x209 & ~x227 & ~x251 & ~x252 & ~x256 & ~x259 & ~x260 & ~x263 & ~x264 & ~x286 & ~x290 & ~x312 & ~x314 & ~x336 & ~x342 & ~x392 & ~x500 & ~x560 & ~x617 & ~x640 & ~x645 & ~x646 & ~x650 & ~x652 & ~x660 & ~x663 & ~x666 & ~x667 & ~x668 & ~x676 & ~x679 & ~x680 & ~x686 & ~x691 & ~x694 & ~x695 & ~x698 & ~x713 & ~x717 & ~x719 & ~x723 & ~x727 & ~x728 & ~x734 & ~x746 & ~x749 & ~x750 & ~x755 & ~x763 & ~x764 & ~x766 & ~x770 & ~x771 & ~x773 & ~x776 & ~x777;
assign c774 =  x359 &  x428 &  x436 & ~x18 & ~x36 & ~x38 & ~x43 & ~x73 & ~x84 & ~x94 & ~x101 & ~x144 & ~x149 & ~x171 & ~x207 & ~x234 & ~x340 & ~x450 & ~x616 & ~x693 & ~x728 & ~x753 & ~x782 & ~x783;
assign c776 =  x458 & ~x0 & ~x2 & ~x4 & ~x7 & ~x8 & ~x9 & ~x10 & ~x11 & ~x12 & ~x14 & ~x17 & ~x18 & ~x22 & ~x24 & ~x26 & ~x27 & ~x31 & ~x33 & ~x34 & ~x35 & ~x36 & ~x39 & ~x41 & ~x44 & ~x47 & ~x49 & ~x55 & ~x57 & ~x58 & ~x60 & ~x61 & ~x63 & ~x67 & ~x70 & ~x72 & ~x77 & ~x78 & ~x85 & ~x86 & ~x89 & ~x91 & ~x94 & ~x95 & ~x102 & ~x104 & ~x105 & ~x107 & ~x108 & ~x110 & ~x111 & ~x113 & ~x115 & ~x117 & ~x120 & ~x121 & ~x123 & ~x125 & ~x126 & ~x127 & ~x130 & ~x135 & ~x139 & ~x140 & ~x141 & ~x145 & ~x149 & ~x150 & ~x151 & ~x153 & ~x154 & ~x160 & ~x161 & ~x162 & ~x164 & ~x165 & ~x166 & ~x167 & ~x168 & ~x169 & ~x173 & ~x174 & ~x175 & ~x176 & ~x177 & ~x178 & ~x181 & ~x182 & ~x193 & ~x194 & ~x195 & ~x197 & ~x198 & ~x199 & ~x205 & ~x207 & ~x208 & ~x209 & ~x222 & ~x223 & ~x224 & ~x235 & ~x236 & ~x250 & ~x252 & ~x253 & ~x256 & ~x257 & ~x258 & ~x259 & ~x261 & ~x278 & ~x279 & ~x282 & ~x291 & ~x293 & ~x312 & ~x314 & ~x317 & ~x336 & ~x339 & ~x342 & ~x343 & ~x345 & ~x346 & ~x368 & ~x369 & ~x370 & ~x371 & ~x397 & ~x588 & ~x645 & ~x647 & ~x653 & ~x656 & ~x658 & ~x659 & ~x660 & ~x666 & ~x667 & ~x669 & ~x670 & ~x672 & ~x673 & ~x674 & ~x675 & ~x677 & ~x679 & ~x681 & ~x684 & ~x687 & ~x688 & ~x692 & ~x695 & ~x697 & ~x704 & ~x706 & ~x708 & ~x709 & ~x710 & ~x712 & ~x716 & ~x724 & ~x726 & ~x733 & ~x740 & ~x742 & ~x743 & ~x745 & ~x749 & ~x751 & ~x752 & ~x756 & ~x761 & ~x764 & ~x765 & ~x766 & ~x767 & ~x768 & ~x771 & ~x772 & ~x775 & ~x777 & ~x778 & ~x781;
assign c778 = ~x15 & ~x16 & ~x23 & ~x51 & ~x62 & ~x68 & ~x76 & ~x87 & ~x94 & ~x106 & ~x125 & ~x141 & ~x143 & ~x245 & ~x272 & ~x273 & ~x288 & ~x293 & ~x300 & ~x308 & ~x313 & ~x328 & ~x329 & ~x336 & ~x339 & ~x369 & ~x648 & ~x668 & ~x676 & ~x686 & ~x715 & ~x722 & ~x726 & ~x759 & ~x761;
assign c780 =  x369;
assign c782 = ~x8 & ~x11 & ~x15 & ~x23 & ~x44 & ~x58 & ~x67 & ~x76 & ~x85 & ~x101 & ~x108 & ~x129 & ~x130 & ~x140 & ~x142 & ~x163 & ~x164 & ~x178 & ~x181 & ~x182 & ~x199 & ~x208 & ~x231 & ~x232 & ~x233 & ~x257 & ~x310 & ~x339 & ~x397 & ~x428 & ~x533 & ~x596 & ~x599 & ~x612 & ~x650 & ~x653 & ~x688 & ~x689 & ~x690 & ~x706 & ~x724 & ~x726 & ~x729 & ~x739 & ~x742 & ~x758 & ~x759 & ~x766 & ~x771;
assign c784 =  x577 &  x578 & ~x1 & ~x2 & ~x10 & ~x12 & ~x17 & ~x18 & ~x22 & ~x24 & ~x33 & ~x38 & ~x45 & ~x51 & ~x53 & ~x54 & ~x58 & ~x66 & ~x68 & ~x78 & ~x82 & ~x84 & ~x92 & ~x102 & ~x103 & ~x120 & ~x124 & ~x125 & ~x145 & ~x151 & ~x159 & ~x165 & ~x169 & ~x175 & ~x187 & ~x188 & ~x200 & ~x205 & ~x209 & ~x218 & ~x225 & ~x226 & ~x250 & ~x253 & ~x278 & ~x280 & ~x281 & ~x307 & ~x310 & ~x311 & ~x338 & ~x339 & ~x364 & ~x392 & ~x629 & ~x644 & ~x660 & ~x669 & ~x672 & ~x679 & ~x681 & ~x683 & ~x684 & ~x694 & ~x697 & ~x700 & ~x702 & ~x704 & ~x705 & ~x707 & ~x710 & ~x721 & ~x722 & ~x732 & ~x742 & ~x746 & ~x750 & ~x758 & ~x768 & ~x771 & ~x775;
assign c786 =  x472 & ~x8 & ~x12 & ~x15 & ~x39 & ~x44 & ~x45 & ~x57 & ~x65 & ~x66 & ~x71 & ~x84 & ~x90 & ~x95 & ~x112 & ~x114 & ~x118 & ~x120 & ~x151 & ~x167 & ~x176 & ~x180 & ~x199 & ~x204 & ~x208 & ~x225 & ~x287 & ~x308 & ~x312 & ~x314 & ~x398 & ~x582 & ~x585 & ~x612 & ~x641 & ~x697 & ~x710 & ~x712 & ~x715 & ~x723 & ~x724 & ~x729 & ~x738 & ~x746 & ~x764 & ~x781;
assign c788 =  x293 &  x319 &  x344 &  x345 & ~x12 & ~x23 & ~x24 & ~x30 & ~x44 & ~x49 & ~x51 & ~x73 & ~x81 & ~x92 & ~x131 & ~x142 & ~x161 & ~x224 & ~x230 & ~x257 & ~x258 & ~x617 & ~x649 & ~x660 & ~x664 & ~x669 & ~x689 & ~x715 & ~x717 & ~x720 & ~x739 & ~x753 & ~x771;
assign c790 = ~x9 & ~x21 & ~x24 & ~x25 & ~x29 & ~x40 & ~x43 & ~x58 & ~x67 & ~x78 & ~x99 & ~x113 & ~x115 & ~x118 & ~x121 & ~x128 & ~x148 & ~x150 & ~x165 & ~x167 & ~x172 & ~x177 & ~x189 & ~x196 & ~x205 & ~x206 & ~x225 & ~x230 & ~x258 & ~x280 & ~x307 & ~x308 & ~x338 & ~x451 & ~x482 & ~x483 & ~x532 & ~x588 & ~x618 & ~x638 & ~x653 & ~x655 & ~x656 & ~x666 & ~x667 & ~x668 & ~x670 & ~x675 & ~x687 & ~x729 & ~x744 & ~x752 & ~x763 & ~x769;
assign c792 = ~x7 & ~x38 & ~x45 & ~x60 & ~x72 & ~x104 & ~x115 & ~x129 & ~x136 & ~x147 & ~x167 & ~x175 & ~x191 & ~x193 & ~x194 & ~x195 & ~x196 & ~x206 & ~x207 & ~x232 & ~x263 & ~x283 & ~x290 & ~x312 & ~x316 & ~x337 & ~x365 & ~x368 & ~x616 & ~x617 & ~x670 & ~x673 & ~x676 & ~x689 & ~x695 & ~x718 & ~x722 & ~x741 & ~x746 & ~x761 & ~x769 & ~x773 & ~x781 & ~x783;
assign c794 =  x334 &  x446 &  x458 &  x514 &  x524 &  x525 & ~x146 & ~x450;
assign c796 =  x334 & ~x17 & ~x18 & ~x19 & ~x21 & ~x28 & ~x33 & ~x59 & ~x61 & ~x111 & ~x113 & ~x114 & ~x117 & ~x119 & ~x142 & ~x147 & ~x172 & ~x197 & ~x233 & ~x235 & ~x254 & ~x261 & ~x509 & ~x532 & ~x598 & ~x780 & ~x781;
assign c798 =  x407 &  x417 & ~x6 & ~x17 & ~x19 & ~x24 & ~x46 & ~x97 & ~x101 & ~x104 & ~x105 & ~x110 & ~x111 & ~x131 & ~x134 & ~x136 & ~x148 & ~x162 & ~x175 & ~x188 & ~x197 & ~x218 & ~x231 & ~x247 & ~x256 & ~x278 & ~x283 & ~x369 & ~x393 & ~x615 & ~x638 & ~x667 & ~x668 & ~x672 & ~x686 & ~x703 & ~x704 & ~x712 & ~x716 & ~x720 & ~x722 & ~x723 & ~x733 & ~x739 & ~x741 & ~x744 & ~x746 & ~x747 & ~x751 & ~x754 & ~x756 & ~x760 & ~x762 & ~x765;
assign c7100 =  x390 & ~x0 & ~x2 & ~x15 & ~x19 & ~x25 & ~x28 & ~x42 & ~x51 & ~x54 & ~x55 & ~x56 & ~x58 & ~x63 & ~x66 & ~x71 & ~x73 & ~x86 & ~x88 & ~x89 & ~x93 & ~x97 & ~x125 & ~x136 & ~x141 & ~x143 & ~x145 & ~x152 & ~x154 & ~x170 & ~x171 & ~x172 & ~x173 & ~x174 & ~x175 & ~x176 & ~x179 & ~x182 & ~x189 & ~x190 & ~x194 & ~x200 & ~x201 & ~x205 & ~x211 & ~x220 & ~x226 & ~x232 & ~x234 & ~x235 & ~x258 & ~x259 & ~x262 & ~x272 & ~x282 & ~x285 & ~x288 & ~x300 & ~x301 & ~x311 & ~x314 & ~x596 & ~x603 & ~x611 & ~x614 & ~x626 & ~x629 & ~x636 & ~x638 & ~x645 & ~x650 & ~x652 & ~x655 & ~x661 & ~x665 & ~x668 & ~x674 & ~x676 & ~x678 & ~x679 & ~x682 & ~x684 & ~x694 & ~x698 & ~x708 & ~x709 & ~x712 & ~x713 & ~x715 & ~x718 & ~x721 & ~x722 & ~x723 & ~x724 & ~x728 & ~x729 & ~x734 & ~x739 & ~x740 & ~x742 & ~x747 & ~x749 & ~x758 & ~x766 & ~x768 & ~x769 & ~x770 & ~x771 & ~x773 & ~x774 & ~x775 & ~x777 & ~x781;
assign c7102 = ~x47 & ~x122 & ~x164 & ~x174 & ~x228 & ~x454 & ~x507 & ~x539 & ~x590 & ~x598 & ~x779 & ~x780;
assign c7104 =  x347 &  x350 &  x375 &  x401 &  x415 &  x427 &  x428 &  x433 &  x444 & ~x6 & ~x11 & ~x28 & ~x50 & ~x53 & ~x96 & ~x137 & ~x139 & ~x147 & ~x152 & ~x189 & ~x196 & ~x217 & ~x253 & ~x255 & ~x310 & ~x642 & ~x646 & ~x648 & ~x654 & ~x658 & ~x666 & ~x685 & ~x692 & ~x745 & ~x747 & ~x753 & ~x771;
assign c7106 = ~x8 & ~x14 & ~x22 & ~x44 & ~x46 & ~x49 & ~x55 & ~x85 & ~x100 & ~x105 & ~x113 & ~x115 & ~x136 & ~x140 & ~x144 & ~x149 & ~x150 & ~x153 & ~x173 & ~x176 & ~x177 & ~x281 & ~x336 & ~x337 & ~x346 & ~x368 & ~x372 & ~x397 & ~x399 & ~x426 & ~x452 & ~x564 & ~x687 & ~x705 & ~x713;
assign c7108 =  x323 &  x350 &  x386 &  x403 &  x417 &  x445 & ~x0 & ~x2 & ~x3 & ~x5 & ~x9 & ~x12 & ~x14 & ~x15 & ~x23 & ~x25 & ~x27 & ~x28 & ~x40 & ~x42 & ~x45 & ~x46 & ~x51 & ~x58 & ~x61 & ~x62 & ~x64 & ~x66 & ~x67 & ~x68 & ~x71 & ~x72 & ~x73 & ~x75 & ~x81 & ~x85 & ~x89 & ~x91 & ~x93 & ~x97 & ~x99 & ~x100 & ~x102 & ~x106 & ~x109 & ~x115 & ~x116 & ~x119 & ~x120 & ~x123 & ~x125 & ~x128 & ~x136 & ~x139 & ~x151 & ~x152 & ~x153 & ~x155 & ~x161 & ~x168 & ~x171 & ~x175 & ~x179 & ~x181 & ~x183 & ~x192 & ~x196 & ~x205 & ~x210 & ~x223 & ~x232 & ~x233 & ~x253 & ~x257 & ~x280 & ~x282 & ~x284 & ~x286 & ~x289 & ~x308 & ~x310 & ~x312 & ~x336 & ~x338 & ~x363 & ~x645 & ~x646 & ~x647 & ~x648 & ~x657 & ~x659 & ~x661 & ~x665 & ~x666 & ~x667 & ~x671 & ~x672 & ~x674 & ~x678 & ~x681 & ~x691 & ~x695 & ~x705 & ~x707 & ~x711 & ~x715 & ~x716 & ~x719 & ~x720 & ~x721 & ~x724 & ~x725 & ~x729 & ~x730 & ~x731 & ~x733 & ~x737 & ~x739 & ~x741 & ~x742 & ~x744 & ~x745 & ~x748 & ~x749 & ~x751 & ~x753 & ~x762 & ~x764 & ~x766 & ~x768 & ~x772 & ~x776 & ~x782;
assign c7110 = ~x7 & ~x13 & ~x56 & ~x62 & ~x107 & ~x110 & ~x127 & ~x141 & ~x151 & ~x162 & ~x170 & ~x173 & ~x177 & ~x206 & ~x226 & ~x231 & ~x280 & ~x290 & ~x335 & ~x393 & ~x452 & ~x453 & ~x454 & ~x455 & ~x596 & ~x599 & ~x628 & ~x687 & ~x696 & ~x701 & ~x751 & ~x753 & ~x769 & ~x773 & ~x777;
assign c7112 =  x390 & ~x11 & ~x51 & ~x203 & ~x272 & ~x300 & ~x301 & ~x581 & ~x584 & ~x585;
assign c7114 =  x361 &  x634 & ~x2 & ~x7 & ~x12 & ~x14 & ~x20 & ~x30 & ~x39 & ~x53 & ~x63 & ~x76 & ~x85 & ~x90 & ~x96 & ~x136 & ~x146 & ~x204 & ~x207 & ~x229 & ~x311 & ~x316 & ~x678 & ~x723 & ~x736 & ~x752;
assign c7116 =  x214 & ~x11 & ~x48 & ~x109 & ~x141 & ~x178 & ~x194 & ~x203 & ~x233 & ~x338 & ~x451 & ~x640 & ~x707 & ~x783;
assign c7118 =  x292 &  x318 & ~x5 & ~x11 & ~x13 & ~x16 & ~x20 & ~x27 & ~x29 & ~x38 & ~x41 & ~x43 & ~x46 & ~x50 & ~x53 & ~x55 & ~x56 & ~x61 & ~x66 & ~x71 & ~x73 & ~x79 & ~x82 & ~x88 & ~x91 & ~x92 & ~x98 & ~x99 & ~x105 & ~x108 & ~x110 & ~x111 & ~x113 & ~x115 & ~x124 & ~x131 & ~x135 & ~x136 & ~x140 & ~x145 & ~x149 & ~x150 & ~x159 & ~x161 & ~x168 & ~x169 & ~x171 & ~x172 & ~x173 & ~x174 & ~x177 & ~x191 & ~x195 & ~x196 & ~x198 & ~x200 & ~x202 & ~x203 & ~x204 & ~x224 & ~x225 & ~x227 & ~x228 & ~x230 & ~x231 & ~x232 & ~x251 & ~x260 & ~x286 & ~x336 & ~x419 & ~x590 & ~x606 & ~x616 & ~x618 & ~x620 & ~x622 & ~x645 & ~x646 & ~x649 & ~x650 & ~x651 & ~x661 & ~x663 & ~x668 & ~x669 & ~x675 & ~x676 & ~x678 & ~x679 & ~x683 & ~x689 & ~x691 & ~x695 & ~x697 & ~x699 & ~x702 & ~x704 & ~x705 & ~x707 & ~x710 & ~x712 & ~x713 & ~x715 & ~x717 & ~x721 & ~x723 & ~x724 & ~x729 & ~x730 & ~x744 & ~x746 & ~x747 & ~x756 & ~x761 & ~x762 & ~x772 & ~x774 & ~x776 & ~x777 & ~x779 & ~x782;
assign c7120 =  x213 &  x331 &  x514 & ~x9 & ~x12 & ~x19 & ~x65 & ~x76 & ~x94 & ~x116 & ~x119 & ~x120 & ~x137 & ~x164 & ~x166 & ~x175 & ~x194 & ~x198 & ~x204 & ~x206 & ~x221 & ~x222 & ~x235 & ~x258 & ~x259 & ~x262 & ~x280 & ~x283 & ~x286 & ~x307 & ~x308 & ~x309 & ~x314 & ~x338 & ~x747 & ~x766 & ~x783;
assign c7122 =  x371 &  x394 & ~x45 & ~x96 & ~x127 & ~x157 & ~x173 & ~x195 & ~x204 & ~x207 & ~x231 & ~x654 & ~x663 & ~x710 & ~x713 & ~x716 & ~x746;
assign c7124 =  x359 &  x409 &  x573 &  x574 &  x575 &  x576 &  x577 &  x578 & ~x3 & ~x4 & ~x6 & ~x14 & ~x15 & ~x20 & ~x29 & ~x31 & ~x46 & ~x51 & ~x52 & ~x53 & ~x55 & ~x57 & ~x61 & ~x65 & ~x69 & ~x71 & ~x73 & ~x75 & ~x76 & ~x77 & ~x83 & ~x89 & ~x92 & ~x96 & ~x104 & ~x105 & ~x106 & ~x108 & ~x121 & ~x133 & ~x134 & ~x135 & ~x141 & ~x144 & ~x146 & ~x147 & ~x151 & ~x152 & ~x163 & ~x164 & ~x169 & ~x174 & ~x177 & ~x196 & ~x199 & ~x205 & ~x208 & ~x235 & ~x254 & ~x258 & ~x260 & ~x262 & ~x281 & ~x283 & ~x285 & ~x286 & ~x287 & ~x288 & ~x309 & ~x310 & ~x311 & ~x312 & ~x315 & ~x391 & ~x613 & ~x627 & ~x636 & ~x676 & ~x700 & ~x714 & ~x717 & ~x718 & ~x722 & ~x726 & ~x731 & ~x735 & ~x738 & ~x740 & ~x743 & ~x745 & ~x749 & ~x756 & ~x775;
assign c7126 =  x462 &  x464 &  x542 & ~x0 & ~x7 & ~x14 & ~x17 & ~x38 & ~x39 & ~x42 & ~x50 & ~x52 & ~x58 & ~x62 & ~x65 & ~x72 & ~x73 & ~x74 & ~x76 & ~x108 & ~x111 & ~x117 & ~x120 & ~x140 & ~x146 & ~x151 & ~x167 & ~x168 & ~x174 & ~x203 & ~x205 & ~x234 & ~x254 & ~x261 & ~x279 & ~x281 & ~x340 & ~x342 & ~x343 & ~x367 & ~x448 & ~x585 & ~x616 & ~x635 & ~x641 & ~x662 & ~x675 & ~x694 & ~x696 & ~x704 & ~x714 & ~x723 & ~x726 & ~x727 & ~x736 & ~x738 & ~x739 & ~x740 & ~x751 & ~x753 & ~x754 & ~x764 & ~x765 & ~x778;
assign c7128 =  x297 &  x348 &  x374 & ~x3 & ~x4 & ~x14 & ~x29 & ~x33 & ~x65 & ~x66 & ~x85 & ~x88 & ~x111 & ~x115 & ~x120 & ~x121 & ~x123 & ~x125 & ~x134 & ~x151 & ~x171 & ~x192 & ~x193 & ~x194 & ~x260 & ~x274 & ~x314 & ~x619 & ~x642 & ~x656 & ~x670 & ~x672 & ~x674 & ~x693 & ~x729 & ~x730 & ~x738 & ~x751 & ~x766 & ~x768 & ~x772 & ~x776 & ~x781 & ~x782;
assign c7130 =  x446 & ~x5 & ~x10 & ~x13 & ~x15 & ~x17 & ~x25 & ~x30 & ~x32 & ~x36 & ~x37 & ~x40 & ~x52 & ~x54 & ~x61 & ~x65 & ~x67 & ~x81 & ~x82 & ~x87 & ~x106 & ~x108 & ~x109 & ~x110 & ~x117 & ~x119 & ~x125 & ~x146 & ~x165 & ~x168 & ~x173 & ~x179 & ~x193 & ~x196 & ~x205 & ~x225 & ~x231 & ~x255 & ~x281 & ~x285 & ~x308 & ~x338 & ~x341 & ~x365 & ~x367 & ~x395 & ~x398 & ~x424 & ~x504 & ~x613 & ~x616 & ~x644 & ~x661 & ~x664 & ~x667 & ~x672 & ~x677 & ~x679 & ~x680 & ~x684 & ~x694 & ~x695 & ~x700 & ~x705 & ~x706 & ~x708 & ~x711 & ~x713 & ~x714 & ~x717 & ~x720 & ~x722 & ~x729 & ~x732 & ~x739 & ~x741 & ~x747 & ~x759 & ~x760 & ~x763 & ~x774 & ~x775 & ~x778 & ~x780 & ~x783;
assign c7132 =  x130;
assign c7134 =  x554 & ~x8 & ~x16 & ~x20 & ~x24 & ~x26 & ~x35 & ~x47 & ~x52 & ~x54 & ~x80 & ~x90 & ~x102 & ~x106 & ~x107 & ~x112 & ~x123 & ~x163 & ~x164 & ~x201 & ~x222 & ~x231 & ~x249 & ~x286 & ~x309 & ~x314 & ~x339 & ~x421 & ~x424 & ~x451 & ~x675 & ~x703 & ~x706 & ~x707 & ~x723 & ~x727 & ~x728 & ~x735 & ~x743 & ~x749 & ~x771;
assign c7136 =  x361 &  x382 &  x444 &  x470 & ~x17 & ~x61 & ~x69 & ~x91 & ~x113 & ~x147 & ~x173 & ~x197 & ~x203 & ~x204 & ~x261 & ~x291 & ~x309 & ~x313 & ~x316 & ~x451 & ~x615 & ~x641 & ~x654 & ~x677 & ~x680 & ~x687 & ~x728 & ~x734 & ~x767;
assign c7138 =  x334 &  x362 &  x383 &  x419 & ~x114 & ~x137 & ~x167 & ~x338;
assign c7140 =  x541 &  x553 & ~x49 & ~x63 & ~x122 & ~x165 & ~x191 & ~x195 & ~x220 & ~x280 & ~x289 & ~x307 & ~x315 & ~x340 & ~x364 & ~x673 & ~x694 & ~x715 & ~x721 & ~x729 & ~x749 & ~x759 & ~x775 & ~x777 & ~x779;
assign c7142 =  x353 &  x417 &  x443 &  x444 & ~x4 & ~x5 & ~x6 & ~x18 & ~x26 & ~x45 & ~x76 & ~x81 & ~x84 & ~x97 & ~x100 & ~x103 & ~x113 & ~x119 & ~x146 & ~x150 & ~x151 & ~x154 & ~x166 & ~x176 & ~x177 & ~x190 & ~x203 & ~x226 & ~x228 & ~x230 & ~x251 & ~x253 & ~x257 & ~x258 & ~x259 & ~x261 & ~x313 & ~x315 & ~x342 & ~x366 & ~x369 & ~x392 & ~x585 & ~x615 & ~x616 & ~x654 & ~x668 & ~x675 & ~x684 & ~x696 & ~x698 & ~x704 & ~x709 & ~x724 & ~x727 & ~x735 & ~x741 & ~x752 & ~x756 & ~x759 & ~x769 & ~x774 & ~x783;
assign c7144 = ~x165 & ~x453;
assign c7146 =  x268 &  x379 &  x404 & ~x4 & ~x5 & ~x7 & ~x10 & ~x12 & ~x15 & ~x16 & ~x18 & ~x19 & ~x20 & ~x22 & ~x23 & ~x27 & ~x30 & ~x33 & ~x34 & ~x36 & ~x38 & ~x39 & ~x40 & ~x42 & ~x43 & ~x49 & ~x57 & ~x61 & ~x62 & ~x63 & ~x66 & ~x67 & ~x69 & ~x70 & ~x71 & ~x73 & ~x75 & ~x76 & ~x79 & ~x80 & ~x81 & ~x82 & ~x83 & ~x86 & ~x88 & ~x89 & ~x90 & ~x92 & ~x93 & ~x96 & ~x98 & ~x99 & ~x101 & ~x103 & ~x105 & ~x106 & ~x108 & ~x109 & ~x112 & ~x113 & ~x115 & ~x116 & ~x118 & ~x119 & ~x120 & ~x121 & ~x122 & ~x124 & ~x125 & ~x128 & ~x133 & ~x134 & ~x135 & ~x137 & ~x140 & ~x141 & ~x145 & ~x147 & ~x150 & ~x151 & ~x154 & ~x155 & ~x159 & ~x160 & ~x161 & ~x166 & ~x167 & ~x170 & ~x172 & ~x173 & ~x174 & ~x176 & ~x178 & ~x179 & ~x180 & ~x181 & ~x194 & ~x195 & ~x196 & ~x197 & ~x204 & ~x205 & ~x228 & ~x229 & ~x230 & ~x231 & ~x232 & ~x234 & ~x250 & ~x253 & ~x258 & ~x260 & ~x261 & ~x280 & ~x281 & ~x286 & ~x287 & ~x308 & ~x309 & ~x310 & ~x312 & ~x313 & ~x314 & ~x336 & ~x580 & ~x582 & ~x588 & ~x616 & ~x617 & ~x618 & ~x645 & ~x647 & ~x648 & ~x650 & ~x654 & ~x657 & ~x658 & ~x659 & ~x661 & ~x662 & ~x663 & ~x664 & ~x665 & ~x668 & ~x669 & ~x670 & ~x671 & ~x672 & ~x673 & ~x674 & ~x675 & ~x676 & ~x678 & ~x685 & ~x686 & ~x687 & ~x689 & ~x691 & ~x692 & ~x693 & ~x696 & ~x697 & ~x700 & ~x702 & ~x704 & ~x705 & ~x707 & ~x708 & ~x715 & ~x717 & ~x718 & ~x719 & ~x720 & ~x721 & ~x724 & ~x728 & ~x731 & ~x732 & ~x734 & ~x737 & ~x738 & ~x740 & ~x742 & ~x746 & ~x748 & ~x750 & ~x752 & ~x753 & ~x754 & ~x756 & ~x758 & ~x764 & ~x765 & ~x766 & ~x769 & ~x770 & ~x774 & ~x776 & ~x777 & ~x779 & ~x781 & ~x783;
assign c7148 = ~x7 & ~x52 & ~x65 & ~x78 & ~x80 & ~x84 & ~x88 & ~x92 & ~x101 & ~x112 & ~x120 & ~x124 & ~x133 & ~x134 & ~x137 & ~x138 & ~x148 & ~x164 & ~x172 & ~x179 & ~x189 & ~x200 & ~x205 & ~x223 & ~x232 & ~x234 & ~x288 & ~x309 & ~x315 & ~x339 & ~x342 & ~x344 & ~x369 & ~x370 & ~x527 & ~x534 & ~x560 & ~x561 & ~x623 & ~x629 & ~x640 & ~x641 & ~x645 & ~x653 & ~x715 & ~x717 & ~x720 & ~x745 & ~x746 & ~x754 & ~x759 & ~x777;
assign c7150 =  x372 &  x422 &  x423 &  x452 &  x483 &  x485 & ~x8 & ~x18 & ~x29 & ~x41 & ~x43 & ~x52 & ~x74 & ~x76 & ~x96 & ~x97 & ~x99 & ~x104 & ~x114 & ~x124 & ~x129 & ~x144 & ~x150 & ~x154 & ~x161 & ~x175 & ~x188 & ~x192 & ~x198 & ~x201 & ~x227 & ~x233 & ~x246 & ~x259 & ~x260 & ~x308 & ~x312 & ~x619 & ~x644 & ~x648 & ~x655 & ~x657 & ~x682 & ~x696 & ~x703 & ~x704 & ~x707 & ~x719 & ~x724 & ~x730 & ~x736 & ~x740 & ~x748 & ~x752 & ~x756 & ~x763 & ~x774 & ~x777;
assign c7152 =  x186 &  x214 &  x241 &  x243 &  x407 &  x429 & ~x12 & ~x35 & ~x54 & ~x59 & ~x81 & ~x118 & ~x615 & ~x667 & ~x712 & ~x716 & ~x745 & ~x747 & ~x769 & ~x781;
assign c7154 =  x214 &  x405 &  x429 &  x483 &  x488 &  x501 & ~x1 & ~x6 & ~x12 & ~x19 & ~x29 & ~x32 & ~x41 & ~x42 & ~x50 & ~x81 & ~x89 & ~x107 & ~x114 & ~x115 & ~x123 & ~x129 & ~x133 & ~x136 & ~x153 & ~x164 & ~x167 & ~x169 & ~x191 & ~x200 & ~x204 & ~x206 & ~x223 & ~x225 & ~x226 & ~x253 & ~x421 & ~x751 & ~x755 & ~x758 & ~x763 & ~x766 & ~x776 & ~x782;
assign c7156 =  x407 & ~x200 & ~x205 & ~x309 & ~x492 & ~x595 & ~x681;
assign c7158 = ~x8 & ~x14 & ~x19 & ~x26 & ~x27 & ~x31 & ~x41 & ~x45 & ~x48 & ~x50 & ~x61 & ~x64 & ~x66 & ~x69 & ~x70 & ~x83 & ~x88 & ~x89 & ~x92 & ~x93 & ~x98 & ~x105 & ~x107 & ~x110 & ~x111 & ~x113 & ~x117 & ~x122 & ~x123 & ~x125 & ~x131 & ~x132 & ~x140 & ~x141 & ~x147 & ~x162 & ~x166 & ~x168 & ~x171 & ~x173 & ~x176 & ~x181 & ~x182 & ~x189 & ~x200 & ~x201 & ~x202 & ~x206 & ~x209 & ~x230 & ~x231 & ~x250 & ~x253 & ~x254 & ~x255 & ~x257 & ~x258 & ~x279 & ~x285 & ~x307 & ~x308 & ~x309 & ~x313 & ~x314 & ~x337 & ~x339 & ~x340 & ~x342 & ~x453 & ~x454 & ~x455 & ~x622 & ~x624 & ~x642 & ~x666 & ~x669 & ~x672 & ~x679 & ~x680 & ~x681 & ~x688 & ~x689 & ~x693 & ~x696 & ~x702 & ~x706 & ~x708 & ~x712 & ~x717 & ~x719 & ~x722 & ~x728 & ~x738 & ~x739 & ~x741 & ~x742 & ~x743 & ~x747 & ~x748 & ~x754 & ~x756 & ~x760 & ~x762 & ~x766 & ~x767 & ~x769 & ~x773 & ~x783;
assign c7160 =  x350 &  x578 & ~x1 & ~x5 & ~x7 & ~x16 & ~x17 & ~x19 & ~x20 & ~x22 & ~x27 & ~x29 & ~x36 & ~x37 & ~x40 & ~x42 & ~x43 & ~x51 & ~x52 & ~x54 & ~x59 & ~x64 & ~x66 & ~x68 & ~x72 & ~x73 & ~x75 & ~x78 & ~x83 & ~x87 & ~x99 & ~x101 & ~x107 & ~x108 & ~x112 & ~x120 & ~x122 & ~x127 & ~x139 & ~x140 & ~x148 & ~x149 & ~x155 & ~x158 & ~x160 & ~x162 & ~x163 & ~x164 & ~x165 & ~x171 & ~x172 & ~x175 & ~x177 & ~x178 & ~x180 & ~x181 & ~x188 & ~x189 & ~x192 & ~x195 & ~x198 & ~x202 & ~x207 & ~x217 & ~x227 & ~x231 & ~x234 & ~x259 & ~x279 & ~x282 & ~x283 & ~x312 & ~x313 & ~x337 & ~x340 & ~x341 & ~x343 & ~x588 & ~x592 & ~x618 & ~x627 & ~x629 & ~x640 & ~x641 & ~x644 & ~x646 & ~x649 & ~x650 & ~x657 & ~x662 & ~x663 & ~x672 & ~x678 & ~x679 & ~x690 & ~x692 & ~x694 & ~x700 & ~x709 & ~x710 & ~x716 & ~x719 & ~x720 & ~x726 & ~x731 & ~x741 & ~x746 & ~x762 & ~x764 & ~x768 & ~x772 & ~x774 & ~x778 & ~x783;
assign c7162 =  x407 &  x461 & ~x3 & ~x6 & ~x7 & ~x23 & ~x26 & ~x30 & ~x34 & ~x35 & ~x39 & ~x41 & ~x43 & ~x50 & ~x55 & ~x58 & ~x61 & ~x73 & ~x79 & ~x89 & ~x90 & ~x94 & ~x98 & ~x101 & ~x111 & ~x130 & ~x132 & ~x136 & ~x137 & ~x139 & ~x145 & ~x147 & ~x149 & ~x153 & ~x161 & ~x166 & ~x167 & ~x174 & ~x182 & ~x198 & ~x203 & ~x225 & ~x230 & ~x285 & ~x287 & ~x308 & ~x317 & ~x342 & ~x343 & ~x370 & ~x393 & ~x447 & ~x560 & ~x586 & ~x599 & ~x600 & ~x644 & ~x646 & ~x651 & ~x652 & ~x656 & ~x662 & ~x664 & ~x672 & ~x678 & ~x684 & ~x685 & ~x690 & ~x691 & ~x695 & ~x696 & ~x704 & ~x706 & ~x708 & ~x718 & ~x720 & ~x721 & ~x726 & ~x730 & ~x736 & ~x742 & ~x757 & ~x772 & ~x778 & ~x779 & ~x781 & ~x782 & ~x783;
assign c7164 =  x269 &  x352 &  x382 &  x400 &  x406 &  x432 &  x458 &  x482 & ~x5 & ~x28 & ~x34 & ~x39 & ~x56 & ~x73 & ~x77 & ~x78 & ~x80 & ~x87 & ~x103 & ~x115 & ~x139 & ~x149 & ~x171 & ~x175 & ~x198 & ~x232 & ~x258 & ~x342 & ~x419 & ~x447 & ~x657 & ~x662 & ~x668 & ~x686 & ~x697 & ~x698 & ~x699 & ~x704 & ~x714 & ~x744 & ~x767;
assign c7166 =  x294 &  x319 &  x400 &  x401 & ~x2 & ~x3 & ~x7 & ~x9 & ~x13 & ~x14 & ~x18 & ~x19 & ~x20 & ~x22 & ~x23 & ~x32 & ~x41 & ~x42 & ~x52 & ~x61 & ~x70 & ~x72 & ~x74 & ~x75 & ~x78 & ~x79 & ~x81 & ~x97 & ~x99 & ~x101 & ~x102 & ~x104 & ~x105 & ~x109 & ~x120 & ~x125 & ~x126 & ~x131 & ~x132 & ~x137 & ~x142 & ~x143 & ~x145 & ~x146 & ~x149 & ~x164 & ~x173 & ~x178 & ~x199 & ~x200 & ~x201 & ~x221 & ~x245 & ~x587 & ~x588 & ~x618 & ~x639 & ~x641 & ~x661 & ~x662 & ~x664 & ~x667 & ~x670 & ~x671 & ~x673 & ~x678 & ~x682 & ~x683 & ~x695 & ~x697 & ~x702 & ~x706 & ~x708 & ~x711 & ~x715 & ~x716 & ~x717 & ~x719 & ~x721 & ~x724 & ~x729 & ~x741 & ~x743 & ~x747 & ~x750 & ~x751 & ~x766 & ~x772 & ~x775;
assign c7168 =  x269 &  x380 & ~x2 & ~x6 & ~x9 & ~x11 & ~x14 & ~x17 & ~x18 & ~x20 & ~x23 & ~x24 & ~x28 & ~x32 & ~x37 & ~x38 & ~x41 & ~x44 & ~x45 & ~x47 & ~x50 & ~x51 & ~x54 & ~x55 & ~x57 & ~x59 & ~x66 & ~x69 & ~x70 & ~x73 & ~x76 & ~x79 & ~x81 & ~x83 & ~x85 & ~x87 & ~x89 & ~x93 & ~x95 & ~x96 & ~x97 & ~x98 & ~x100 & ~x106 & ~x107 & ~x109 & ~x110 & ~x112 & ~x116 & ~x118 & ~x121 & ~x123 & ~x125 & ~x127 & ~x129 & ~x134 & ~x135 & ~x142 & ~x144 & ~x145 & ~x147 & ~x150 & ~x154 & ~x159 & ~x160 & ~x161 & ~x168 & ~x172 & ~x174 & ~x176 & ~x177 & ~x181 & ~x187 & ~x190 & ~x193 & ~x194 & ~x196 & ~x198 & ~x200 & ~x201 & ~x206 & ~x217 & ~x221 & ~x223 & ~x224 & ~x225 & ~x226 & ~x229 & ~x233 & ~x234 & ~x249 & ~x250 & ~x252 & ~x253 & ~x260 & ~x261 & ~x279 & ~x281 & ~x284 & ~x289 & ~x309 & ~x311 & ~x313 & ~x392 & ~x503 & ~x532 & ~x591 & ~x616 & ~x618 & ~x620 & ~x640 & ~x642 & ~x644 & ~x646 & ~x650 & ~x658 & ~x659 & ~x661 & ~x662 & ~x665 & ~x667 & ~x668 & ~x670 & ~x672 & ~x674 & ~x676 & ~x677 & ~x685 & ~x693 & ~x694 & ~x704 & ~x705 & ~x714 & ~x718 & ~x719 & ~x721 & ~x725 & ~x726 & ~x729 & ~x730 & ~x739 & ~x740 & ~x742 & ~x749 & ~x752 & ~x753 & ~x757 & ~x760 & ~x761 & ~x763 & ~x766 & ~x769 & ~x771 & ~x772 & ~x775 & ~x778 & ~x779 & ~x781 & ~x783;
assign c7170 =  x325 &  x355 &  x385 &  x430 &  x436 &  x458 &  x463 &  x545 &  x632 & ~x2 & ~x24 & ~x25 & ~x26 & ~x37 & ~x41 & ~x44 & ~x47 & ~x49 & ~x54 & ~x64 & ~x86 & ~x121 & ~x124 & ~x137 & ~x141 & ~x202 & ~x207 & ~x225 & ~x227 & ~x258 & ~x260 & ~x263 & ~x284 & ~x343 & ~x449 & ~x450 & ~x715 & ~x740 & ~x745 & ~x755 & ~x761;
assign c7172 =  x406 &  x484 &  x495 &  x499 &  x522 &  x523 & ~x0 & ~x7 & ~x15 & ~x26 & ~x36 & ~x39 & ~x44 & ~x50 & ~x53 & ~x66 & ~x70 & ~x75 & ~x76 & ~x78 & ~x81 & ~x82 & ~x90 & ~x95 & ~x97 & ~x98 & ~x107 & ~x114 & ~x117 & ~x123 & ~x131 & ~x154 & ~x160 & ~x172 & ~x197 & ~x200 & ~x205 & ~x209 & ~x221 & ~x222 & ~x229 & ~x233 & ~x253 & ~x256 & ~x258 & ~x281 & ~x314 & ~x339 & ~x393 & ~x425 & ~x642 & ~x648 & ~x660 & ~x669 & ~x698 & ~x706 & ~x719 & ~x721 & ~x727 & ~x732 & ~x753 & ~x754 & ~x766 & ~x778;
assign c7174 =  x606 & ~x9 & ~x18 & ~x45 & ~x63 & ~x71 & ~x154 & ~x160 & ~x197 & ~x199 & ~x206 & ~x254 & ~x262 & ~x283 & ~x290 & ~x397 & ~x636 & ~x660 & ~x667 & ~x672 & ~x674 & ~x691 & ~x692 & ~x765 & ~x775 & ~x779 & ~x782;
assign c7176 =  x130 &  x446 &  x551;
assign c7178 =  x389 &  x463 & ~x4 & ~x13 & ~x18 & ~x21 & ~x22 & ~x24 & ~x26 & ~x27 & ~x32 & ~x46 & ~x51 & ~x52 & ~x53 & ~x58 & ~x62 & ~x63 & ~x64 & ~x67 & ~x77 & ~x82 & ~x87 & ~x88 & ~x91 & ~x96 & ~x97 & ~x98 & ~x101 & ~x140 & ~x146 & ~x148 & ~x149 & ~x167 & ~x173 & ~x176 & ~x178 & ~x180 & ~x196 & ~x198 & ~x209 & ~x224 & ~x227 & ~x228 & ~x230 & ~x232 & ~x252 & ~x257 & ~x261 & ~x282 & ~x283 & ~x312 & ~x501 & ~x676 & ~x680 & ~x685 & ~x704 & ~x709 & ~x713 & ~x714 & ~x716 & ~x727 & ~x740 & ~x750 & ~x761 & ~x764 & ~x770 & ~x771 & ~x775 & ~x778 & ~x779;
assign c7180 =  x353 &  x374 & ~x3 & ~x12 & ~x17 & ~x26 & ~x27 & ~x28 & ~x29 & ~x32 & ~x38 & ~x39 & ~x42 & ~x43 & ~x46 & ~x52 & ~x56 & ~x61 & ~x63 & ~x66 & ~x68 & ~x69 & ~x71 & ~x73 & ~x74 & ~x79 & ~x80 & ~x81 & ~x83 & ~x85 & ~x89 & ~x91 & ~x95 & ~x97 & ~x98 & ~x99 & ~x100 & ~x101 & ~x102 & ~x103 & ~x104 & ~x105 & ~x107 & ~x108 & ~x112 & ~x124 & ~x125 & ~x139 & ~x144 & ~x146 & ~x149 & ~x154 & ~x159 & ~x166 & ~x168 & ~x170 & ~x175 & ~x176 & ~x178 & ~x180 & ~x198 & ~x200 & ~x202 & ~x203 & ~x205 & ~x216 & ~x226 & ~x227 & ~x228 & ~x231 & ~x257 & ~x280 & ~x312 & ~x526 & ~x590 & ~x641 & ~x644 & ~x650 & ~x651 & ~x657 & ~x659 & ~x663 & ~x664 & ~x665 & ~x666 & ~x669 & ~x677 & ~x681 & ~x686 & ~x687 & ~x689 & ~x692 & ~x694 & ~x695 & ~x696 & ~x698 & ~x700 & ~x706 & ~x713 & ~x714 & ~x715 & ~x717 & ~x720 & ~x724 & ~x726 & ~x729 & ~x740 & ~x742 & ~x747 & ~x751 & ~x752 & ~x756 & ~x758 & ~x760 & ~x763 & ~x764 & ~x768 & ~x770 & ~x772 & ~x776 & ~x778 & ~x779 & ~x783;
assign c7182 =  x631 & ~x78 & ~x82 & ~x141 & ~x163 & ~x175 & ~x180 & ~x192 & ~x393;
assign c7184 =  x359 &  x389 &  x415 &  x417 &  x439 &  x441 &  x445 &  x446 & ~x16 & ~x21 & ~x40 & ~x41 & ~x54 & ~x83 & ~x89 & ~x93 & ~x95 & ~x108 & ~x146 & ~x150 & ~x151 & ~x169 & ~x170 & ~x174 & ~x178 & ~x200 & ~x205 & ~x207 & ~x230 & ~x231 & ~x254 & ~x258 & ~x313 & ~x314 & ~x505 & ~x588 & ~x615 & ~x636 & ~x637 & ~x640 & ~x699 & ~x700 & ~x720 & ~x732 & ~x768 & ~x774 & ~x780;
assign c7186 =  x406 &  x407 &  x551 & ~x1 & ~x7 & ~x8 & ~x12 & ~x13 & ~x15 & ~x18 & ~x27 & ~x29 & ~x37 & ~x41 & ~x44 & ~x47 & ~x56 & ~x62 & ~x82 & ~x86 & ~x89 & ~x96 & ~x101 & ~x109 & ~x118 & ~x120 & ~x128 & ~x135 & ~x164 & ~x167 & ~x169 & ~x172 & ~x174 & ~x175 & ~x178 & ~x179 & ~x199 & ~x206 & ~x207 & ~x208 & ~x224 & ~x228 & ~x229 & ~x230 & ~x232 & ~x233 & ~x234 & ~x253 & ~x255 & ~x256 & ~x259 & ~x279 & ~x281 & ~x282 & ~x308 & ~x310 & ~x364 & ~x583 & ~x616 & ~x617 & ~x618 & ~x642 & ~x648 & ~x652 & ~x655 & ~x659 & ~x661 & ~x662 & ~x663 & ~x664 & ~x669 & ~x673 & ~x687 & ~x699 & ~x700 & ~x702 & ~x705 & ~x706 & ~x707 & ~x710 & ~x712 & ~x713 & ~x716 & ~x717 & ~x718 & ~x719 & ~x721 & ~x734 & ~x738 & ~x743 & ~x744 & ~x746 & ~x747 & ~x749 & ~x750 & ~x752 & ~x761 & ~x762 & ~x771 & ~x777 & ~x778;
assign c7188 =  x630 & ~x8 & ~x61 & ~x63 & ~x116 & ~x146 & ~x150 & ~x152 & ~x169 & ~x255 & ~x340 & ~x667 & ~x680 & ~x683 & ~x684 & ~x689 & ~x718 & ~x743 & ~x751 & ~x774;
assign c7190 =  x461 &  x606 & ~x9 & ~x15 & ~x20 & ~x23 & ~x32 & ~x108 & ~x112 & ~x135 & ~x171 & ~x174 & ~x181 & ~x197 & ~x199 & ~x203 & ~x232 & ~x234 & ~x259 & ~x307 & ~x309 & ~x312 & ~x342 & ~x365 & ~x368 & ~x589 & ~x642 & ~x651 & ~x667 & ~x670 & ~x677 & ~x703 & ~x704 & ~x710 & ~x718 & ~x719 & ~x726 & ~x735 & ~x761 & ~x767 & ~x774 & ~x781;
assign c7192 =  x292 &  x345 & ~x2 & ~x3 & ~x7 & ~x9 & ~x10 & ~x11 & ~x12 & ~x14 & ~x15 & ~x28 & ~x31 & ~x33 & ~x36 & ~x37 & ~x42 & ~x43 & ~x44 & ~x47 & ~x48 & ~x49 & ~x52 & ~x56 & ~x57 & ~x58 & ~x62 & ~x63 & ~x68 & ~x69 & ~x70 & ~x71 & ~x72 & ~x77 & ~x78 & ~x80 & ~x83 & ~x84 & ~x86 & ~x87 & ~x88 & ~x89 & ~x90 & ~x91 & ~x92 & ~x97 & ~x98 & ~x101 & ~x105 & ~x107 & ~x108 & ~x115 & ~x118 & ~x121 & ~x122 & ~x123 & ~x127 & ~x128 & ~x134 & ~x137 & ~x139 & ~x143 & ~x144 & ~x148 & ~x151 & ~x152 & ~x155 & ~x167 & ~x173 & ~x174 & ~x176 & ~x177 & ~x179 & ~x190 & ~x197 & ~x199 & ~x200 & ~x201 & ~x203 & ~x204 & ~x207 & ~x217 & ~x222 & ~x223 & ~x224 & ~x225 & ~x227 & ~x228 & ~x229 & ~x231 & ~x253 & ~x254 & ~x255 & ~x257 & ~x258 & ~x259 & ~x260 & ~x279 & ~x280 & ~x285 & ~x308 & ~x589 & ~x616 & ~x620 & ~x635 & ~x636 & ~x637 & ~x638 & ~x640 & ~x641 & ~x643 & ~x644 & ~x645 & ~x646 & ~x648 & ~x657 & ~x658 & ~x659 & ~x666 & ~x667 & ~x672 & ~x677 & ~x680 & ~x681 & ~x683 & ~x684 & ~x685 & ~x686 & ~x687 & ~x691 & ~x695 & ~x696 & ~x697 & ~x700 & ~x701 & ~x707 & ~x710 & ~x711 & ~x712 & ~x714 & ~x715 & ~x717 & ~x719 & ~x723 & ~x724 & ~x728 & ~x729 & ~x730 & ~x739 & ~x742 & ~x743 & ~x744 & ~x746 & ~x748 & ~x750 & ~x752 & ~x753 & ~x754 & ~x760 & ~x761 & ~x762 & ~x763 & ~x764 & ~x765 & ~x766 & ~x769 & ~x770 & ~x772 & ~x773 & ~x779 & ~x780 & ~x782 & ~x783;
assign c7194 =  x359 &  x411 &  x434 &  x437 &  x462 &  x491 & ~x0 & ~x1 & ~x7 & ~x11 & ~x15 & ~x27 & ~x37 & ~x41 & ~x42 & ~x46 & ~x49 & ~x52 & ~x54 & ~x60 & ~x61 & ~x62 & ~x66 & ~x69 & ~x70 & ~x74 & ~x75 & ~x76 & ~x81 & ~x83 & ~x85 & ~x86 & ~x87 & ~x93 & ~x97 & ~x104 & ~x105 & ~x111 & ~x117 & ~x118 & ~x119 & ~x125 & ~x128 & ~x130 & ~x131 & ~x133 & ~x135 & ~x138 & ~x139 & ~x143 & ~x144 & ~x146 & ~x147 & ~x148 & ~x149 & ~x152 & ~x155 & ~x159 & ~x164 & ~x166 & ~x168 & ~x176 & ~x178 & ~x179 & ~x180 & ~x181 & ~x182 & ~x190 & ~x193 & ~x194 & ~x195 & ~x198 & ~x201 & ~x203 & ~x211 & ~x218 & ~x220 & ~x221 & ~x224 & ~x227 & ~x231 & ~x232 & ~x252 & ~x253 & ~x255 & ~x257 & ~x259 & ~x260 & ~x262 & ~x279 & ~x280 & ~x281 & ~x282 & ~x286 & ~x307 & ~x315 & ~x317 & ~x335 & ~x338 & ~x339 & ~x341 & ~x343 & ~x344 & ~x365 & ~x393 & ~x420 & ~x643 & ~x644 & ~x651 & ~x655 & ~x660 & ~x662 & ~x664 & ~x666 & ~x668 & ~x669 & ~x673 & ~x676 & ~x679 & ~x680 & ~x681 & ~x683 & ~x684 & ~x696 & ~x697 & ~x700 & ~x711 & ~x718 & ~x721 & ~x722 & ~x723 & ~x731 & ~x733 & ~x735 & ~x736 & ~x740 & ~x743 & ~x744 & ~x747 & ~x748 & ~x749 & ~x757 & ~x758 & ~x763 & ~x764 & ~x765 & ~x767 & ~x769 & ~x770 & ~x774 & ~x777 & ~x779;
assign c7196 = ~x5 & ~x11 & ~x12 & ~x13 & ~x14 & ~x29 & ~x32 & ~x33 & ~x39 & ~x52 & ~x55 & ~x74 & ~x77 & ~x96 & ~x103 & ~x104 & ~x107 & ~x120 & ~x154 & ~x168 & ~x173 & ~x195 & ~x229 & ~x284 & ~x314 & ~x338 & ~x372 & ~x374 & ~x425 & ~x426 & ~x428 & ~x455 & ~x588 & ~x672 & ~x692 & ~x696 & ~x712 & ~x715 & ~x722 & ~x736 & ~x765 & ~x767 & ~x771;
assign c7198 = ~x35 & ~x70 & ~x96 & ~x129 & ~x131 & ~x151 & ~x182 & ~x300 & ~x311 & ~x351 & ~x430 & ~x682;
assign c7200 = ~x20 & ~x21 & ~x26 & ~x31 & ~x32 & ~x35 & ~x50 & ~x56 & ~x62 & ~x68 & ~x75 & ~x78 & ~x80 & ~x82 & ~x99 & ~x100 & ~x102 & ~x105 & ~x117 & ~x131 & ~x136 & ~x146 & ~x153 & ~x154 & ~x163 & ~x201 & ~x208 & ~x221 & ~x222 & ~x231 & ~x234 & ~x238 & ~x289 & ~x310 & ~x313 & ~x314 & ~x317 & ~x321 & ~x345 & ~x347 & ~x372 & ~x401 & ~x426 & ~x427 & ~x447 & ~x475 & ~x647 & ~x691 & ~x701 & ~x709 & ~x730 & ~x733 & ~x734 & ~x739 & ~x747 & ~x749 & ~x753 & ~x760 & ~x762 & ~x767 & ~x778;
assign c7202 = ~x2 & ~x13 & ~x14 & ~x17 & ~x18 & ~x22 & ~x24 & ~x26 & ~x33 & ~x34 & ~x35 & ~x40 & ~x48 & ~x53 & ~x58 & ~x59 & ~x61 & ~x65 & ~x68 & ~x69 & ~x72 & ~x74 & ~x77 & ~x104 & ~x105 & ~x106 & ~x126 & ~x127 & ~x140 & ~x141 & ~x147 & ~x148 & ~x149 & ~x155 & ~x157 & ~x159 & ~x160 & ~x163 & ~x164 & ~x166 & ~x175 & ~x176 & ~x177 & ~x181 & ~x196 & ~x198 & ~x220 & ~x226 & ~x227 & ~x228 & ~x229 & ~x246 & ~x255 & ~x261 & ~x280 & ~x281 & ~x285 & ~x286 & ~x303 & ~x314 & ~x337 & ~x392 & ~x425 & ~x426 & ~x620 & ~x621 & ~x629 & ~x646 & ~x649 & ~x650 & ~x657 & ~x659 & ~x665 & ~x669 & ~x675 & ~x676 & ~x688 & ~x689 & ~x690 & ~x692 & ~x695 & ~x697 & ~x698 & ~x707 & ~x708 & ~x712 & ~x713 & ~x718 & ~x720 & ~x730 & ~x740 & ~x741 & ~x744 & ~x747 & ~x753 & ~x760 & ~x772 & ~x776;
assign c7204 =  x617;
assign c7206 =  x241 &  x306 &  x607 & ~x83 & ~x169 & ~x319 & ~x452 & ~x753;
assign c7208 = ~x1 & ~x7 & ~x13 & ~x15 & ~x18 & ~x21 & ~x27 & ~x31 & ~x32 & ~x38 & ~x39 & ~x51 & ~x69 & ~x71 & ~x82 & ~x89 & ~x103 & ~x117 & ~x132 & ~x163 & ~x171 & ~x179 & ~x181 & ~x182 & ~x197 & ~x233 & ~x261 & ~x314 & ~x338 & ~x364 & ~x369 & ~x400 & ~x419 & ~x425 & ~x426 & ~x452 & ~x562 & ~x563 & ~x648 & ~x693 & ~x716 & ~x719 & ~x725 & ~x734 & ~x738 & ~x745 & ~x748 & ~x749 & ~x756 & ~x760 & ~x766 & ~x770 & ~x782;
assign c7210 = ~x3 & ~x4 & ~x6 & ~x14 & ~x16 & ~x17 & ~x19 & ~x25 & ~x33 & ~x37 & ~x39 & ~x42 & ~x43 & ~x45 & ~x49 & ~x52 & ~x60 & ~x65 & ~x66 & ~x73 & ~x86 & ~x92 & ~x102 & ~x107 & ~x110 & ~x111 & ~x116 & ~x117 & ~x124 & ~x133 & ~x137 & ~x138 & ~x141 & ~x142 & ~x143 & ~x148 & ~x150 & ~x169 & ~x177 & ~x183 & ~x184 & ~x185 & ~x193 & ~x195 & ~x198 & ~x203 & ~x216 & ~x223 & ~x225 & ~x243 & ~x244 & ~x245 & ~x247 & ~x251 & ~x253 & ~x272 & ~x279 & ~x300 & ~x308 & ~x392 & ~x511 & ~x512 & ~x561 & ~x589 & ~x594 & ~x605 & ~x611 & ~x615 & ~x653 & ~x668 & ~x670 & ~x671 & ~x676 & ~x711 & ~x728 & ~x736 & ~x738 & ~x739 & ~x740 & ~x747 & ~x749 & ~x770 & ~x773 & ~x774;
assign c7212 = ~x0 & ~x5 & ~x20 & ~x24 & ~x38 & ~x40 & ~x41 & ~x43 & ~x49 & ~x54 & ~x66 & ~x76 & ~x77 & ~x85 & ~x93 & ~x103 & ~x105 & ~x107 & ~x110 & ~x112 & ~x118 & ~x137 & ~x138 & ~x149 & ~x163 & ~x167 & ~x168 & ~x170 & ~x174 & ~x191 & ~x192 & ~x201 & ~x203 & ~x206 & ~x208 & ~x223 & ~x225 & ~x226 & ~x228 & ~x229 & ~x230 & ~x232 & ~x233 & ~x282 & ~x283 & ~x287 & ~x311 & ~x313 & ~x315 & ~x338 & ~x453 & ~x454 & ~x455 & ~x587 & ~x604 & ~x605 & ~x609 & ~x610 & ~x622 & ~x628 & ~x630 & ~x632 & ~x636 & ~x638 & ~x643 & ~x645 & ~x651 & ~x658 & ~x661 & ~x664 & ~x669 & ~x671 & ~x675 & ~x678 & ~x680 & ~x682 & ~x686 & ~x687 & ~x688 & ~x692 & ~x701 & ~x703 & ~x704 & ~x706 & ~x708 & ~x714 & ~x722 & ~x727 & ~x728 & ~x729 & ~x730 & ~x732 & ~x736 & ~x737 & ~x738 & ~x744 & ~x747 & ~x750 & ~x757 & ~x760 & ~x765 & ~x771 & ~x775 & ~x778 & ~x779 & ~x781;
assign c7214 =  x297 &  x321 &  x346 &  x350 &  x380 &  x381 & ~x1 & ~x3 & ~x4 & ~x5 & ~x6 & ~x8 & ~x10 & ~x11 & ~x13 & ~x16 & ~x17 & ~x19 & ~x21 & ~x22 & ~x24 & ~x25 & ~x27 & ~x31 & ~x34 & ~x35 & ~x38 & ~x39 & ~x40 & ~x41 & ~x42 & ~x44 & ~x45 & ~x46 & ~x48 & ~x49 & ~x52 & ~x54 & ~x55 & ~x56 & ~x57 & ~x58 & ~x59 & ~x60 & ~x61 & ~x63 & ~x66 & ~x68 & ~x70 & ~x71 & ~x72 & ~x75 & ~x76 & ~x77 & ~x79 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x87 & ~x88 & ~x90 & ~x92 & ~x93 & ~x94 & ~x96 & ~x97 & ~x100 & ~x101 & ~x102 & ~x105 & ~x106 & ~x107 & ~x109 & ~x110 & ~x113 & ~x114 & ~x118 & ~x120 & ~x121 & ~x122 & ~x125 & ~x126 & ~x128 & ~x129 & ~x133 & ~x134 & ~x139 & ~x143 & ~x145 & ~x147 & ~x148 & ~x149 & ~x150 & ~x151 & ~x152 & ~x156 & ~x160 & ~x165 & ~x168 & ~x170 & ~x171 & ~x174 & ~x175 & ~x176 & ~x177 & ~x179 & ~x180 & ~x195 & ~x197 & ~x198 & ~x200 & ~x202 & ~x203 & ~x204 & ~x205 & ~x208 & ~x224 & ~x226 & ~x228 & ~x231 & ~x233 & ~x234 & ~x235 & ~x252 & ~x253 & ~x255 & ~x256 & ~x258 & ~x259 & ~x260 & ~x261 & ~x280 & ~x281 & ~x283 & ~x285 & ~x286 & ~x288 & ~x308 & ~x309 & ~x311 & ~x312 & ~x560 & ~x588 & ~x589 & ~x616 & ~x617 & ~x618 & ~x640 & ~x641 & ~x642 & ~x643 & ~x648 & ~x650 & ~x651 & ~x654 & ~x655 & ~x656 & ~x660 & ~x661 & ~x665 & ~x666 & ~x668 & ~x669 & ~x670 & ~x673 & ~x674 & ~x675 & ~x676 & ~x678 & ~x685 & ~x687 & ~x688 & ~x691 & ~x692 & ~x698 & ~x700 & ~x703 & ~x705 & ~x706 & ~x707 & ~x708 & ~x710 & ~x714 & ~x716 & ~x719 & ~x720 & ~x721 & ~x726 & ~x728 & ~x730 & ~x732 & ~x735 & ~x736 & ~x737 & ~x738 & ~x739 & ~x743 & ~x744 & ~x745 & ~x748 & ~x749 & ~x750 & ~x751 & ~x752 & ~x753 & ~x754 & ~x755 & ~x756 & ~x757 & ~x758 & ~x764 & ~x765 & ~x766 & ~x768 & ~x769 & ~x771 & ~x772 & ~x775 & ~x776 & ~x778 & ~x779 & ~x780 & ~x781 & ~x782 & ~x783;
assign c7216 =  x362 &  x445 & ~x1 & ~x3 & ~x4 & ~x6 & ~x8 & ~x11 & ~x12 & ~x13 & ~x14 & ~x15 & ~x16 & ~x17 & ~x19 & ~x20 & ~x22 & ~x28 & ~x31 & ~x37 & ~x40 & ~x41 & ~x45 & ~x47 & ~x50 & ~x51 & ~x53 & ~x55 & ~x56 & ~x57 & ~x58 & ~x59 & ~x61 & ~x62 & ~x65 & ~x66 & ~x69 & ~x71 & ~x73 & ~x74 & ~x75 & ~x79 & ~x83 & ~x84 & ~x89 & ~x90 & ~x94 & ~x97 & ~x98 & ~x100 & ~x102 & ~x106 & ~x107 & ~x109 & ~x112 & ~x116 & ~x119 & ~x122 & ~x123 & ~x125 & ~x126 & ~x127 & ~x132 & ~x134 & ~x135 & ~x136 & ~x139 & ~x143 & ~x146 & ~x147 & ~x149 & ~x151 & ~x152 & ~x153 & ~x154 & ~x159 & ~x160 & ~x163 & ~x164 & ~x165 & ~x168 & ~x174 & ~x178 & ~x179 & ~x180 & ~x183 & ~x190 & ~x192 & ~x198 & ~x199 & ~x200 & ~x201 & ~x205 & ~x207 & ~x224 & ~x226 & ~x232 & ~x235 & ~x252 & ~x253 & ~x255 & ~x256 & ~x259 & ~x262 & ~x280 & ~x281 & ~x282 & ~x283 & ~x284 & ~x308 & ~x314 & ~x337 & ~x340 & ~x570 & ~x581 & ~x582 & ~x588 & ~x617 & ~x639 & ~x641 & ~x642 & ~x643 & ~x644 & ~x645 & ~x649 & ~x650 & ~x651 & ~x654 & ~x657 & ~x658 & ~x659 & ~x660 & ~x661 & ~x662 & ~x663 & ~x665 & ~x667 & ~x668 & ~x670 & ~x671 & ~x674 & ~x676 & ~x679 & ~x680 & ~x681 & ~x691 & ~x692 & ~x695 & ~x702 & ~x705 & ~x707 & ~x709 & ~x710 & ~x711 & ~x712 & ~x714 & ~x717 & ~x721 & ~x722 & ~x724 & ~x725 & ~x728 & ~x729 & ~x731 & ~x733 & ~x734 & ~x738 & ~x742 & ~x749 & ~x750 & ~x753 & ~x755 & ~x756 & ~x761 & ~x765 & ~x766 & ~x768 & ~x770 & ~x772 & ~x774 & ~x775 & ~x776 & ~x778 & ~x779;
assign c7218 =  x387 &  x388 &  x415 &  x416 &  x438 &  x445 & ~x2 & ~x3 & ~x4 & ~x5 & ~x9 & ~x10 & ~x12 & ~x13 & ~x14 & ~x16 & ~x17 & ~x19 & ~x22 & ~x24 & ~x25 & ~x26 & ~x28 & ~x30 & ~x31 & ~x32 & ~x35 & ~x38 & ~x39 & ~x40 & ~x41 & ~x44 & ~x45 & ~x46 & ~x47 & ~x48 & ~x49 & ~x50 & ~x51 & ~x59 & ~x64 & ~x67 & ~x71 & ~x73 & ~x75 & ~x77 & ~x78 & ~x81 & ~x83 & ~x84 & ~x91 & ~x93 & ~x96 & ~x98 & ~x99 & ~x100 & ~x101 & ~x102 & ~x104 & ~x105 & ~x106 & ~x109 & ~x110 & ~x115 & ~x117 & ~x122 & ~x123 & ~x124 & ~x125 & ~x127 & ~x129 & ~x130 & ~x136 & ~x137 & ~x138 & ~x139 & ~x141 & ~x145 & ~x146 & ~x148 & ~x150 & ~x152 & ~x160 & ~x165 & ~x167 & ~x169 & ~x170 & ~x172 & ~x177 & ~x178 & ~x181 & ~x191 & ~x192 & ~x193 & ~x194 & ~x195 & ~x201 & ~x202 & ~x203 & ~x217 & ~x223 & ~x225 & ~x226 & ~x227 & ~x228 & ~x245 & ~x250 & ~x251 & ~x252 & ~x253 & ~x254 & ~x273 & ~x282 & ~x309 & ~x338 & ~x366 & ~x392 & ~x560 & ~x589 & ~x615 & ~x618 & ~x619 & ~x621 & ~x622 & ~x629 & ~x632 & ~x633 & ~x634 & ~x635 & ~x636 & ~x640 & ~x641 & ~x649 & ~x652 & ~x655 & ~x656 & ~x657 & ~x658 & ~x659 & ~x663 & ~x664 & ~x665 & ~x667 & ~x669 & ~x672 & ~x675 & ~x676 & ~x678 & ~x680 & ~x681 & ~x682 & ~x683 & ~x686 & ~x689 & ~x690 & ~x691 & ~x696 & ~x698 & ~x699 & ~x700 & ~x703 & ~x705 & ~x706 & ~x707 & ~x713 & ~x715 & ~x721 & ~x722 & ~x723 & ~x724 & ~x729 & ~x730 & ~x731 & ~x735 & ~x738 & ~x739 & ~x740 & ~x742 & ~x746 & ~x748 & ~x751 & ~x753 & ~x754 & ~x755 & ~x758 & ~x759 & ~x762 & ~x763 & ~x764 & ~x769 & ~x771 & ~x773 & ~x774 & ~x777 & ~x782;
assign c7220 =  x293 &  x294 &  x319 &  x320 & ~x0 & ~x1 & ~x2 & ~x3 & ~x6 & ~x7 & ~x8 & ~x12 & ~x16 & ~x18 & ~x20 & ~x21 & ~x22 & ~x23 & ~x25 & ~x26 & ~x28 & ~x29 & ~x31 & ~x33 & ~x34 & ~x36 & ~x38 & ~x39 & ~x40 & ~x41 & ~x42 & ~x44 & ~x46 & ~x47 & ~x51 & ~x52 & ~x53 & ~x59 & ~x60 & ~x61 & ~x63 & ~x64 & ~x68 & ~x70 & ~x71 & ~x74 & ~x75 & ~x76 & ~x77 & ~x78 & ~x79 & ~x80 & ~x81 & ~x82 & ~x83 & ~x85 & ~x86 & ~x88 & ~x89 & ~x90 & ~x92 & ~x93 & ~x94 & ~x95 & ~x96 & ~x98 & ~x104 & ~x105 & ~x106 & ~x108 & ~x109 & ~x110 & ~x111 & ~x112 & ~x119 & ~x120 & ~x123 & ~x127 & ~x128 & ~x129 & ~x130 & ~x131 & ~x137 & ~x139 & ~x140 & ~x141 & ~x143 & ~x146 & ~x149 & ~x150 & ~x151 & ~x152 & ~x153 & ~x156 & ~x163 & ~x164 & ~x165 & ~x166 & ~x168 & ~x170 & ~x171 & ~x174 & ~x175 & ~x176 & ~x179 & ~x181 & ~x188 & ~x189 & ~x194 & ~x195 & ~x196 & ~x198 & ~x200 & ~x201 & ~x202 & ~x205 & ~x217 & ~x222 & ~x224 & ~x225 & ~x228 & ~x229 & ~x230 & ~x231 & ~x232 & ~x251 & ~x252 & ~x253 & ~x257 & ~x259 & ~x287 & ~x308 & ~x336 & ~x532 & ~x560 & ~x587 & ~x588 & ~x589 & ~x590 & ~x593 & ~x594 & ~x615 & ~x617 & ~x618 & ~x619 & ~x621 & ~x622 & ~x623 & ~x624 & ~x626 & ~x627 & ~x629 & ~x632 & ~x633 & ~x634 & ~x637 & ~x638 & ~x639 & ~x640 & ~x641 & ~x644 & ~x647 & ~x648 & ~x649 & ~x650 & ~x652 & ~x653 & ~x656 & ~x657 & ~x659 & ~x660 & ~x661 & ~x662 & ~x663 & ~x664 & ~x665 & ~x667 & ~x670 & ~x671 & ~x675 & ~x676 & ~x677 & ~x678 & ~x680 & ~x682 & ~x683 & ~x685 & ~x686 & ~x687 & ~x688 & ~x689 & ~x690 & ~x693 & ~x694 & ~x695 & ~x696 & ~x698 & ~x699 & ~x700 & ~x701 & ~x702 & ~x703 & ~x704 & ~x705 & ~x706 & ~x707 & ~x708 & ~x710 & ~x712 & ~x713 & ~x714 & ~x716 & ~x717 & ~x718 & ~x721 & ~x722 & ~x723 & ~x725 & ~x727 & ~x729 & ~x730 & ~x731 & ~x733 & ~x734 & ~x736 & ~x737 & ~x738 & ~x742 & ~x743 & ~x744 & ~x747 & ~x748 & ~x749 & ~x750 & ~x752 & ~x753 & ~x755 & ~x756 & ~x758 & ~x762 & ~x763 & ~x765 & ~x766 & ~x771 & ~x772 & ~x773 & ~x775 & ~x776 & ~x777 & ~x780 & ~x781;
assign c7222 =  x349 &  x374 &  x375 &  x401 &  x424 &  x426 &  x451 &  x478 & ~x5 & ~x9 & ~x35 & ~x58 & ~x62 & ~x72 & ~x83 & ~x96 & ~x131 & ~x144 & ~x170 & ~x173 & ~x179 & ~x222 & ~x231 & ~x252 & ~x253 & ~x255 & ~x259 & ~x286 & ~x308 & ~x617 & ~x619 & ~x650 & ~x654 & ~x660 & ~x661 & ~x665 & ~x666 & ~x668 & ~x677 & ~x678 & ~x681 & ~x682 & ~x691 & ~x698 & ~x705 & ~x712 & ~x720 & ~x726 & ~x727 & ~x728 & ~x732 & ~x743 & ~x745 & ~x748 & ~x750 & ~x756 & ~x761 & ~x762 & ~x779 & ~x780;
assign c7224 =  x439 &  x468 & ~x1 & ~x9 & ~x25 & ~x43 & ~x67 & ~x91 & ~x106 & ~x115 & ~x118 & ~x147 & ~x151 & ~x152 & ~x162 & ~x172 & ~x191 & ~x199 & ~x201 & ~x205 & ~x238 & ~x267 & ~x284 & ~x293 & ~x313 & ~x339 & ~x420 & ~x637 & ~x643 & ~x688 & ~x701 & ~x739 & ~x748;
assign c7226 =  x457 &  x606 & ~x25 & ~x210 & ~x668 & ~x693 & ~x773;
assign c7228 =  x463 & ~x14 & ~x26 & ~x29 & ~x35 & ~x37 & ~x39 & ~x45 & ~x52 & ~x54 & ~x62 & ~x63 & ~x64 & ~x71 & ~x72 & ~x73 & ~x74 & ~x84 & ~x88 & ~x90 & ~x106 & ~x108 & ~x110 & ~x111 & ~x113 & ~x114 & ~x115 & ~x116 & ~x119 & ~x124 & ~x139 & ~x141 & ~x152 & ~x155 & ~x156 & ~x167 & ~x170 & ~x178 & ~x180 & ~x202 & ~x228 & ~x230 & ~x233 & ~x235 & ~x259 & ~x261 & ~x262 & ~x282 & ~x307 & ~x310 & ~x311 & ~x312 & ~x313 & ~x315 & ~x316 & ~x337 & ~x397 & ~x420 & ~x555 & ~x614 & ~x616 & ~x621 & ~x630 & ~x646 & ~x649 & ~x650 & ~x651 & ~x666 & ~x669 & ~x673 & ~x684 & ~x685 & ~x689 & ~x690 & ~x694 & ~x696 & ~x698 & ~x707 & ~x708 & ~x712 & ~x714 & ~x715 & ~x718 & ~x721 & ~x722 & ~x728 & ~x732 & ~x741 & ~x743 & ~x746 & ~x753 & ~x756 & ~x757 & ~x764 & ~x766 & ~x771;
assign c7230 =  x305 &  x462 &  x660 & ~x374;
assign c7232 =  x348 &  x388 &  x400 &  x416 &  x445 & ~x5 & ~x9 & ~x16 & ~x30 & ~x32 & ~x35 & ~x44 & ~x46 & ~x47 & ~x49 & ~x53 & ~x62 & ~x65 & ~x68 & ~x74 & ~x76 & ~x78 & ~x82 & ~x89 & ~x99 & ~x101 & ~x102 & ~x103 & ~x113 & ~x116 & ~x119 & ~x125 & ~x127 & ~x129 & ~x131 & ~x135 & ~x140 & ~x144 & ~x149 & ~x151 & ~x161 & ~x167 & ~x173 & ~x183 & ~x189 & ~x190 & ~x195 & ~x198 & ~x199 & ~x203 & ~x216 & ~x222 & ~x224 & ~x228 & ~x231 & ~x246 & ~x254 & ~x281 & ~x283 & ~x588 & ~x615 & ~x618 & ~x620 & ~x623 & ~x629 & ~x631 & ~x634 & ~x636 & ~x637 & ~x641 & ~x649 & ~x654 & ~x665 & ~x667 & ~x671 & ~x672 & ~x675 & ~x681 & ~x689 & ~x690 & ~x691 & ~x699 & ~x700 & ~x706 & ~x707 & ~x709 & ~x710 & ~x711 & ~x718 & ~x720 & ~x723 & ~x725 & ~x728 & ~x730 & ~x737 & ~x740 & ~x744 & ~x754 & ~x772 & ~x782 & ~x783;
assign c7234 =  x323 &  x349 &  x353 &  x375 &  x384 &  x403 &  x451 &  x458 &  x460 &  x479 &  x483 &  x484 & ~x0 & ~x1 & ~x2 & ~x3 & ~x4 & ~x6 & ~x7 & ~x8 & ~x10 & ~x11 & ~x12 & ~x13 & ~x14 & ~x15 & ~x16 & ~x17 & ~x18 & ~x19 & ~x22 & ~x23 & ~x24 & ~x25 & ~x28 & ~x29 & ~x31 & ~x32 & ~x33 & ~x34 & ~x35 & ~x36 & ~x38 & ~x40 & ~x42 & ~x44 & ~x45 & ~x46 & ~x47 & ~x49 & ~x50 & ~x51 & ~x52 & ~x53 & ~x54 & ~x55 & ~x56 & ~x57 & ~x58 & ~x59 & ~x61 & ~x62 & ~x63 & ~x64 & ~x65 & ~x66 & ~x68 & ~x69 & ~x71 & ~x72 & ~x73 & ~x75 & ~x76 & ~x79 & ~x80 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x87 & ~x88 & ~x89 & ~x92 & ~x93 & ~x95 & ~x96 & ~x97 & ~x98 & ~x99 & ~x101 & ~x103 & ~x104 & ~x106 & ~x107 & ~x108 & ~x110 & ~x111 & ~x112 & ~x113 & ~x114 & ~x115 & ~x116 & ~x117 & ~x119 & ~x120 & ~x122 & ~x123 & ~x124 & ~x125 & ~x126 & ~x127 & ~x129 & ~x130 & ~x131 & ~x132 & ~x133 & ~x134 & ~x135 & ~x136 & ~x137 & ~x138 & ~x140 & ~x141 & ~x142 & ~x144 & ~x145 & ~x146 & ~x147 & ~x148 & ~x150 & ~x151 & ~x152 & ~x153 & ~x154 & ~x156 & ~x158 & ~x160 & ~x162 & ~x166 & ~x168 & ~x170 & ~x171 & ~x172 & ~x173 & ~x174 & ~x175 & ~x176 & ~x178 & ~x179 & ~x180 & ~x181 & ~x182 & ~x183 & ~x196 & ~x197 & ~x198 & ~x199 & ~x200 & ~x202 & ~x204 & ~x205 & ~x206 & ~x208 & ~x210 & ~x223 & ~x224 & ~x227 & ~x228 & ~x229 & ~x230 & ~x231 & ~x232 & ~x233 & ~x234 & ~x252 & ~x253 & ~x254 & ~x255 & ~x256 & ~x257 & ~x258 & ~x259 & ~x260 & ~x261 & ~x280 & ~x282 & ~x283 & ~x284 & ~x285 & ~x286 & ~x287 & ~x288 & ~x309 & ~x314 & ~x315 & ~x316 & ~x335 & ~x336 & ~x560 & ~x588 & ~x589 & ~x616 & ~x617 & ~x618 & ~x619 & ~x620 & ~x626 & ~x627 & ~x631 & ~x634 & ~x635 & ~x636 & ~x638 & ~x639 & ~x641 & ~x644 & ~x645 & ~x647 & ~x648 & ~x649 & ~x650 & ~x656 & ~x657 & ~x659 & ~x660 & ~x661 & ~x662 & ~x663 & ~x664 & ~x665 & ~x666 & ~x670 & ~x671 & ~x673 & ~x674 & ~x675 & ~x677 & ~x678 & ~x679 & ~x681 & ~x682 & ~x683 & ~x685 & ~x686 & ~x687 & ~x688 & ~x689 & ~x690 & ~x692 & ~x695 & ~x696 & ~x697 & ~x698 & ~x699 & ~x700 & ~x701 & ~x703 & ~x704 & ~x705 & ~x706 & ~x707 & ~x709 & ~x710 & ~x711 & ~x712 & ~x714 & ~x715 & ~x719 & ~x720 & ~x722 & ~x723 & ~x724 & ~x725 & ~x726 & ~x728 & ~x729 & ~x730 & ~x731 & ~x732 & ~x733 & ~x734 & ~x735 & ~x736 & ~x737 & ~x738 & ~x739 & ~x740 & ~x741 & ~x743 & ~x744 & ~x745 & ~x746 & ~x747 & ~x749 & ~x750 & ~x751 & ~x752 & ~x753 & ~x754 & ~x757 & ~x758 & ~x761 & ~x762 & ~x763 & ~x764 & ~x766 & ~x768 & ~x770 & ~x771 & ~x772 & ~x773 & ~x776 & ~x777 & ~x779 & ~x780 & ~x781 & ~x782 & ~x783;
assign c7236 = ~x28 & ~x70 & ~x116 & ~x149 & ~x171 & ~x222 & ~x225 & ~x260 & ~x313 & ~x392 & ~x454 & ~x481 & ~x482 & ~x483 & ~x588 & ~x589 & ~x686 & ~x694 & ~x707 & ~x725 & ~x729 & ~x754 & ~x768;
assign c7238 =  x347 &  x373 &  x441 &  x442 &  x469 &  x470 &  x471 &  x490 & ~x0 & ~x2 & ~x4 & ~x9 & ~x28 & ~x29 & ~x30 & ~x31 & ~x34 & ~x39 & ~x43 & ~x46 & ~x48 & ~x49 & ~x53 & ~x56 & ~x61 & ~x63 & ~x64 & ~x67 & ~x68 & ~x72 & ~x73 & ~x81 & ~x84 & ~x85 & ~x86 & ~x87 & ~x88 & ~x89 & ~x90 & ~x91 & ~x95 & ~x99 & ~x100 & ~x104 & ~x112 & ~x119 & ~x122 & ~x124 & ~x125 & ~x126 & ~x133 & ~x143 & ~x145 & ~x146 & ~x148 & ~x149 & ~x151 & ~x152 & ~x153 & ~x160 & ~x161 & ~x166 & ~x167 & ~x168 & ~x169 & ~x170 & ~x171 & ~x176 & ~x178 & ~x197 & ~x204 & ~x205 & ~x207 & ~x210 & ~x224 & ~x225 & ~x228 & ~x251 & ~x252 & ~x258 & ~x307 & ~x336 & ~x364 & ~x588 & ~x589 & ~x612 & ~x613 & ~x635 & ~x636 & ~x637 & ~x640 & ~x641 & ~x642 & ~x643 & ~x645 & ~x648 & ~x650 & ~x661 & ~x665 & ~x666 & ~x667 & ~x668 & ~x678 & ~x686 & ~x687 & ~x691 & ~x692 & ~x697 & ~x698 & ~x703 & ~x708 & ~x709 & ~x713 & ~x714 & ~x715 & ~x717 & ~x718 & ~x719 & ~x721 & ~x723 & ~x727 & ~x729 & ~x730 & ~x733 & ~x734 & ~x735 & ~x736 & ~x742 & ~x746 & ~x749 & ~x752 & ~x753 & ~x759 & ~x764 & ~x766 & ~x767 & ~x768 & ~x775 & ~x779 & ~x780 & ~x781 & ~x783;
assign c7240 =  x455 &  x456 &  x457 &  x483 &  x576 & ~x2 & ~x5 & ~x35 & ~x40 & ~x87 & ~x95 & ~x112 & ~x113 & ~x133 & ~x134 & ~x136 & ~x137 & ~x144 & ~x155 & ~x156 & ~x165 & ~x169 & ~x178 & ~x181 & ~x182 & ~x183 & ~x207 & ~x208 & ~x209 & ~x210 & ~x226 & ~x227 & ~x237 & ~x238 & ~x258 & ~x264 & ~x265 & ~x284 & ~x309 & ~x312 & ~x315 & ~x318 & ~x344 & ~x364 & ~x365 & ~x366 & ~x369 & ~x648 & ~x671 & ~x684 & ~x690 & ~x692 & ~x694 & ~x704 & ~x735 & ~x736 & ~x746 & ~x750 & ~x763 & ~x772 & ~x774;
assign c7242 =  x355 &  x378 &  x404 &  x433 & ~x0 & ~x1 & ~x4 & ~x5 & ~x9 & ~x10 & ~x11 & ~x13 & ~x17 & ~x20 & ~x21 & ~x22 & ~x24 & ~x27 & ~x29 & ~x32 & ~x34 & ~x35 & ~x36 & ~x41 & ~x43 & ~x45 & ~x47 & ~x48 & ~x49 & ~x50 & ~x54 & ~x56 & ~x57 & ~x59 & ~x61 & ~x62 & ~x64 & ~x65 & ~x66 & ~x69 & ~x71 & ~x72 & ~x73 & ~x75 & ~x77 & ~x80 & ~x84 & ~x85 & ~x88 & ~x89 & ~x92 & ~x95 & ~x96 & ~x97 & ~x101 & ~x104 & ~x105 & ~x106 & ~x107 & ~x109 & ~x110 & ~x114 & ~x115 & ~x117 & ~x119 & ~x120 & ~x122 & ~x123 & ~x124 & ~x126 & ~x127 & ~x129 & ~x131 & ~x133 & ~x135 & ~x136 & ~x137 & ~x138 & ~x140 & ~x141 & ~x142 & ~x143 & ~x145 & ~x147 & ~x148 & ~x149 & ~x152 & ~x153 & ~x160 & ~x161 & ~x163 & ~x164 & ~x167 & ~x171 & ~x173 & ~x176 & ~x177 & ~x178 & ~x180 & ~x181 & ~x182 & ~x189 & ~x190 & ~x196 & ~x197 & ~x198 & ~x199 & ~x201 & ~x202 & ~x206 & ~x208 & ~x223 & ~x224 & ~x226 & ~x227 & ~x228 & ~x229 & ~x231 & ~x232 & ~x235 & ~x236 & ~x251 & ~x252 & ~x253 & ~x256 & ~x259 & ~x260 & ~x283 & ~x284 & ~x285 & ~x286 & ~x288 & ~x289 & ~x309 & ~x310 & ~x311 & ~x312 & ~x313 & ~x314 & ~x315 & ~x337 & ~x339 & ~x340 & ~x343 & ~x364 & ~x392 & ~x420 & ~x447 & ~x496 & ~x588 & ~x616 & ~x617 & ~x618 & ~x619 & ~x644 & ~x645 & ~x646 & ~x647 & ~x648 & ~x650 & ~x651 & ~x654 & ~x655 & ~x658 & ~x659 & ~x662 & ~x663 & ~x664 & ~x665 & ~x666 & ~x668 & ~x671 & ~x673 & ~x676 & ~x677 & ~x680 & ~x681 & ~x683 & ~x684 & ~x686 & ~x694 & ~x695 & ~x696 & ~x697 & ~x698 & ~x699 & ~x700 & ~x701 & ~x702 & ~x703 & ~x704 & ~x706 & ~x707 & ~x710 & ~x711 & ~x713 & ~x714 & ~x716 & ~x717 & ~x718 & ~x719 & ~x722 & ~x723 & ~x725 & ~x726 & ~x727 & ~x729 & ~x730 & ~x731 & ~x732 & ~x733 & ~x734 & ~x735 & ~x736 & ~x737 & ~x740 & ~x741 & ~x744 & ~x745 & ~x747 & ~x748 & ~x749 & ~x750 & ~x751 & ~x753 & ~x754 & ~x756 & ~x758 & ~x759 & ~x760 & ~x761 & ~x762 & ~x764 & ~x767 & ~x769 & ~x770 & ~x771 & ~x772 & ~x774 & ~x776 & ~x778 & ~x780 & ~x781 & ~x782;
assign c7244 =  x296 &  x375 &  x418 & ~x13 & ~x143 & ~x235 & ~x283 & ~x285 & ~x286 & ~x479 & ~x532 & ~x783;
assign c7246 = ~x13 & ~x15 & ~x17 & ~x21 & ~x33 & ~x40 & ~x42 & ~x48 & ~x56 & ~x57 & ~x71 & ~x79 & ~x87 & ~x91 & ~x105 & ~x107 & ~x109 & ~x121 & ~x122 & ~x135 & ~x136 & ~x152 & ~x162 & ~x164 & ~x167 & ~x171 & ~x191 & ~x195 & ~x205 & ~x218 & ~x220 & ~x222 & ~x223 & ~x224 & ~x260 & ~x281 & ~x308 & ~x309 & ~x313 & ~x337 & ~x344 & ~x369 & ~x392 & ~x402 & ~x427 & ~x454 & ~x616 & ~x617 & ~x673 & ~x678 & ~x681 & ~x682 & ~x687 & ~x689 & ~x700 & ~x705 & ~x717 & ~x724 & ~x729 & ~x740 & ~x743 & ~x752 & ~x754 & ~x759 & ~x768 & ~x772;
assign c7248 = ~x0 & ~x1 & ~x6 & ~x29 & ~x33 & ~x34 & ~x38 & ~x41 & ~x43 & ~x62 & ~x64 & ~x67 & ~x71 & ~x77 & ~x78 & ~x83 & ~x84 & ~x87 & ~x90 & ~x91 & ~x98 & ~x99 & ~x100 & ~x101 & ~x111 & ~x114 & ~x119 & ~x120 & ~x122 & ~x125 & ~x126 & ~x128 & ~x129 & ~x131 & ~x138 & ~x152 & ~x154 & ~x168 & ~x174 & ~x175 & ~x176 & ~x178 & ~x193 & ~x196 & ~x198 & ~x205 & ~x207 & ~x225 & ~x235 & ~x253 & ~x254 & ~x261 & ~x262 & ~x263 & ~x280 & ~x286 & ~x287 & ~x289 & ~x290 & ~x307 & ~x316 & ~x338 & ~x341 & ~x344 & ~x370 & ~x396 & ~x398 & ~x399 & ~x560 & ~x588 & ~x645 & ~x646 & ~x652 & ~x654 & ~x663 & ~x673 & ~x675 & ~x676 & ~x677 & ~x685 & ~x686 & ~x687 & ~x690 & ~x693 & ~x694 & ~x699 & ~x700 & ~x701 & ~x707 & ~x709 & ~x710 & ~x714 & ~x718 & ~x720 & ~x721 & ~x723 & ~x728 & ~x738 & ~x740 & ~x745 & ~x748 & ~x756 & ~x761 & ~x765 & ~x771 & ~x778 & ~x780 & ~x783;
assign c7250 =  x634 & ~x4 & ~x21 & ~x27 & ~x28 & ~x55 & ~x64 & ~x146 & ~x148 & ~x150 & ~x163 & ~x165 & ~x170 & ~x177 & ~x194 & ~x195 & ~x202 & ~x235 & ~x255 & ~x285 & ~x314 & ~x315 & ~x338 & ~x342 & ~x369 & ~x393 & ~x398 & ~x424 & ~x699 & ~x722 & ~x752 & ~x758 & ~x768 & ~x775 & ~x783;
assign c7252 =  x215 &  x334 &  x353 &  x362 &  x457 &  x502 & ~x8 & ~x60 & ~x76 & ~x77 & ~x103 & ~x106 & ~x111 & ~x114 & ~x118 & ~x142 & ~x145 & ~x147 & ~x151 & ~x171 & ~x200 & ~x235 & ~x254 & ~x281 & ~x285 & ~x310 & ~x339 & ~x343 & ~x729 & ~x733 & ~x743 & ~x744 & ~x769 & ~x770;
assign c7254 =  x269 &  x351 &  x424 & ~x14 & ~x15 & ~x17 & ~x28 & ~x43 & ~x44 & ~x46 & ~x47 & ~x52 & ~x76 & ~x79 & ~x81 & ~x94 & ~x102 & ~x106 & ~x114 & ~x121 & ~x143 & ~x144 & ~x152 & ~x166 & ~x174 & ~x206 & ~x232 & ~x257 & ~x286 & ~x312 & ~x364 & ~x642 & ~x645 & ~x647 & ~x657 & ~x663 & ~x668 & ~x681 & ~x685 & ~x687 & ~x714 & ~x715 & ~x716 & ~x738 & ~x741 & ~x745 & ~x750 & ~x759 & ~x764 & ~x780;
assign c7256 =  x316;
assign c7258 =  x382 &  x606 &  x607 & ~x7 & ~x22 & ~x35 & ~x99 & ~x129 & ~x138 & ~x163 & ~x280 & ~x310 & ~x673 & ~x674 & ~x685 & ~x722 & ~x756 & ~x768 & ~x773;
assign c7260 =  x268 &  x294 &  x347 &  x373 &  x378 &  x381 &  x465 & ~x1 & ~x8 & ~x14 & ~x16 & ~x21 & ~x22 & ~x24 & ~x25 & ~x31 & ~x45 & ~x55 & ~x60 & ~x71 & ~x73 & ~x74 & ~x75 & ~x91 & ~x96 & ~x98 & ~x105 & ~x112 & ~x113 & ~x115 & ~x125 & ~x137 & ~x171 & ~x226 & ~x227 & ~x254 & ~x280 & ~x281 & ~x287 & ~x310 & ~x312 & ~x313 & ~x365 & ~x587 & ~x588 & ~x646 & ~x648 & ~x649 & ~x677 & ~x688 & ~x690 & ~x692 & ~x693 & ~x694 & ~x705 & ~x712 & ~x716 & ~x717 & ~x724 & ~x727 & ~x735 & ~x757 & ~x767 & ~x769 & ~x771 & ~x776;
assign c7262 =  x382 &  x457 &  x606 & ~x5 & ~x10 & ~x17 & ~x31 & ~x33 & ~x34 & ~x54 & ~x75 & ~x123 & ~x126 & ~x135 & ~x163 & ~x180 & ~x190 & ~x191 & ~x193 & ~x198 & ~x202 & ~x204 & ~x209 & ~x236 & ~x237 & ~x281 & ~x309 & ~x310 & ~x316 & ~x368 & ~x618 & ~x667 & ~x686 & ~x688 & ~x704 & ~x712 & ~x715 & ~x716 & ~x722 & ~x730 & ~x734 & ~x757 & ~x765 & ~x774;
assign c7264 =  x319 &  x382 & ~x60 & ~x128 & ~x130 & ~x199 & ~x503 & ~x551 & ~x554 & ~x710 & ~x717 & ~x730 & ~x752 & ~x769 & ~x782;
assign c7266 = ~x1 & ~x2 & ~x8 & ~x16 & ~x23 & ~x37 & ~x45 & ~x50 & ~x60 & ~x74 & ~x78 & ~x89 & ~x126 & ~x131 & ~x161 & ~x179 & ~x180 & ~x195 & ~x207 & ~x226 & ~x235 & ~x237 & ~x262 & ~x316 & ~x338 & ~x339 & ~x342 & ~x374 & ~x397 & ~x398 & ~x534 & ~x657 & ~x658 & ~x669 & ~x671 & ~x673 & ~x676 & ~x684 & ~x689 & ~x694 & ~x696 & ~x698 & ~x706 & ~x713 & ~x716 & ~x736 & ~x739 & ~x751 & ~x756 & ~x764;
assign c7268 =  x379 &  x402 &  x409 &  x415 &  x416 &  x444 &  x462 &  x483 & ~x0 & ~x7 & ~x17 & ~x34 & ~x35 & ~x43 & ~x52 & ~x64 & ~x65 & ~x67 & ~x85 & ~x88 & ~x105 & ~x112 & ~x117 & ~x118 & ~x120 & ~x124 & ~x133 & ~x142 & ~x145 & ~x149 & ~x168 & ~x169 & ~x174 & ~x182 & ~x189 & ~x190 & ~x202 & ~x203 & ~x205 & ~x209 & ~x225 & ~x226 & ~x227 & ~x255 & ~x280 & ~x308 & ~x310 & ~x313 & ~x339 & ~x364 & ~x366 & ~x369 & ~x370 & ~x394 & ~x475 & ~x618 & ~x645 & ~x646 & ~x659 & ~x660 & ~x669 & ~x678 & ~x679 & ~x685 & ~x687 & ~x688 & ~x690 & ~x695 & ~x696 & ~x697 & ~x701 & ~x705 & ~x707 & ~x708 & ~x709 & ~x713 & ~x720 & ~x722 & ~x723 & ~x728 & ~x729 & ~x733 & ~x734 & ~x735 & ~x742 & ~x747 & ~x750 & ~x751 & ~x752 & ~x753 & ~x755 & ~x762 & ~x764 & ~x768 & ~x770 & ~x779;
assign c7270 = ~x4 & ~x10 & ~x15 & ~x35 & ~x38 & ~x42 & ~x47 & ~x49 & ~x51 & ~x57 & ~x58 & ~x62 & ~x65 & ~x67 & ~x74 & ~x80 & ~x83 & ~x85 & ~x89 & ~x100 & ~x117 & ~x119 & ~x137 & ~x154 & ~x164 & ~x168 & ~x176 & ~x177 & ~x180 & ~x203 & ~x222 & ~x254 & ~x258 & ~x282 & ~x285 & ~x309 & ~x314 & ~x315 & ~x335 & ~x336 & ~x365 & ~x453 & ~x454 & ~x455 & ~x532 & ~x606 & ~x608 & ~x609 & ~x610 & ~x627 & ~x631 & ~x640 & ~x645 & ~x650 & ~x670 & ~x671 & ~x680 & ~x687 & ~x689 & ~x690 & ~x691 & ~x703 & ~x708 & ~x710 & ~x714 & ~x718 & ~x720 & ~x721 & ~x732 & ~x734 & ~x735 & ~x751 & ~x755 & ~x764 & ~x767;
assign c7272 =  x353 &  x417 &  x443 & ~x9 & ~x14 & ~x15 & ~x19 & ~x21 & ~x23 & ~x25 & ~x30 & ~x31 & ~x33 & ~x35 & ~x37 & ~x38 & ~x40 & ~x47 & ~x51 & ~x52 & ~x54 & ~x59 & ~x60 & ~x62 & ~x72 & ~x86 & ~x90 & ~x92 & ~x94 & ~x98 & ~x99 & ~x109 & ~x111 & ~x121 & ~x125 & ~x126 & ~x133 & ~x135 & ~x137 & ~x146 & ~x147 & ~x149 & ~x153 & ~x156 & ~x161 & ~x164 & ~x167 & ~x174 & ~x175 & ~x177 & ~x188 & ~x193 & ~x195 & ~x196 & ~x197 & ~x201 & ~x202 & ~x204 & ~x209 & ~x219 & ~x225 & ~x229 & ~x230 & ~x236 & ~x237 & ~x253 & ~x255 & ~x257 & ~x260 & ~x261 & ~x274 & ~x281 & ~x288 & ~x310 & ~x314 & ~x315 & ~x364 & ~x365 & ~x366 & ~x394 & ~x645 & ~x646 & ~x657 & ~x669 & ~x671 & ~x673 & ~x674 & ~x684 & ~x687 & ~x692 & ~x701 & ~x706 & ~x716 & ~x717 & ~x718 & ~x719 & ~x721 & ~x727 & ~x730 & ~x735 & ~x738 & ~x745 & ~x748 & ~x749 & ~x753 & ~x760 & ~x762 & ~x771 & ~x773 & ~x775 & ~x783;
assign c7274 =  x334 & ~x6 & ~x11 & ~x13 & ~x15 & ~x16 & ~x21 & ~x23 & ~x28 & ~x29 & ~x30 & ~x33 & ~x38 & ~x39 & ~x43 & ~x44 & ~x45 & ~x46 & ~x49 & ~x50 & ~x51 & ~x54 & ~x59 & ~x60 & ~x66 & ~x70 & ~x71 & ~x78 & ~x84 & ~x86 & ~x94 & ~x96 & ~x97 & ~x103 & ~x104 & ~x105 & ~x106 & ~x110 & ~x122 & ~x123 & ~x128 & ~x132 & ~x135 & ~x137 & ~x139 & ~x142 & ~x145 & ~x151 & ~x159 & ~x160 & ~x161 & ~x162 & ~x172 & ~x173 & ~x178 & ~x182 & ~x188 & ~x189 & ~x196 & ~x203 & ~x206 & ~x223 & ~x224 & ~x226 & ~x231 & ~x235 & ~x251 & ~x256 & ~x260 & ~x261 & ~x284 & ~x286 & ~x308 & ~x313 & ~x336 & ~x337 & ~x339 & ~x364 & ~x476 & ~x584 & ~x585 & ~x644 & ~x647 & ~x648 & ~x652 & ~x657 & ~x658 & ~x659 & ~x661 & ~x663 & ~x664 & ~x666 & ~x670 & ~x672 & ~x676 & ~x678 & ~x681 & ~x686 & ~x688 & ~x689 & ~x690 & ~x697 & ~x702 & ~x703 & ~x704 & ~x711 & ~x716 & ~x718 & ~x719 & ~x721 & ~x725 & ~x727 & ~x732 & ~x735 & ~x738 & ~x742 & ~x748 & ~x757 & ~x760 & ~x765 & ~x767 & ~x768 & ~x772 & ~x779 & ~x780 & ~x782 & ~x783;
assign c7276 = ~x23 & ~x34 & ~x39 & ~x40 & ~x41 & ~x42 & ~x44 & ~x59 & ~x69 & ~x84 & ~x91 & ~x99 & ~x114 & ~x115 & ~x123 & ~x135 & ~x149 & ~x163 & ~x177 & ~x183 & ~x195 & ~x197 & ~x201 & ~x204 & ~x209 & ~x224 & ~x232 & ~x233 & ~x251 & ~x253 & ~x254 & ~x255 & ~x261 & ~x263 & ~x284 & ~x285 & ~x286 & ~x309 & ~x311 & ~x313 & ~x344 & ~x453 & ~x557 & ~x619 & ~x648 & ~x651 & ~x662 & ~x663 & ~x682 & ~x691 & ~x700 & ~x740 & ~x741 & ~x742 & ~x755 & ~x767 & ~x771;
assign c7278 = ~x0 & ~x1 & ~x15 & ~x17 & ~x20 & ~x27 & ~x37 & ~x43 & ~x46 & ~x49 & ~x62 & ~x79 & ~x91 & ~x94 & ~x95 & ~x96 & ~x97 & ~x102 & ~x105 & ~x106 & ~x110 & ~x123 & ~x124 & ~x125 & ~x129 & ~x132 & ~x141 & ~x149 & ~x159 & ~x169 & ~x178 & ~x179 & ~x187 & ~x189 & ~x190 & ~x201 & ~x203 & ~x208 & ~x218 & ~x219 & ~x226 & ~x229 & ~x233 & ~x237 & ~x238 & ~x239 & ~x244 & ~x246 & ~x253 & ~x254 & ~x272 & ~x273 & ~x274 & ~x275 & ~x279 & ~x280 & ~x288 & ~x291 & ~x301 & ~x303 & ~x309 & ~x317 & ~x330 & ~x337 & ~x343 & ~x369 & ~x619 & ~x621 & ~x623 & ~x625 & ~x626 & ~x629 & ~x630 & ~x643 & ~x658 & ~x660 & ~x662 & ~x673 & ~x674 & ~x677 & ~x679 & ~x680 & ~x683 & ~x686 & ~x695 & ~x705 & ~x710 & ~x714 & ~x718 & ~x720 & ~x730 & ~x733 & ~x737 & ~x738 & ~x739 & ~x741 & ~x748 & ~x773 & ~x779 & ~x783;
assign c7280 =  x634 & ~x7 & ~x20 & ~x57 & ~x68 & ~x76 & ~x84 & ~x110 & ~x120 & ~x165 & ~x173 & ~x194 & ~x231 & ~x255 & ~x312 & ~x424 & ~x449 & ~x752 & ~x772;
assign c7282 =  x159 &  x187 &  x331 & ~x532;
assign c7284 =  x244 &  x328 &  x330 &  x468 & ~x6 & ~x10 & ~x13 & ~x16 & ~x28 & ~x37 & ~x47 & ~x49 & ~x167 & ~x168 & ~x174 & ~x197 & ~x206 & ~x234 & ~x293 & ~x371 & ~x450 & ~x680 & ~x783;
assign c7286 =  x450 &  x481 &  x513 & ~x4 & ~x9 & ~x17 & ~x22 & ~x30 & ~x42 & ~x43 & ~x45 & ~x47 & ~x51 & ~x55 & ~x57 & ~x64 & ~x66 & ~x71 & ~x72 & ~x78 & ~x82 & ~x84 & ~x85 & ~x90 & ~x91 & ~x96 & ~x100 & ~x101 & ~x109 & ~x122 & ~x125 & ~x126 & ~x129 & ~x132 & ~x137 & ~x141 & ~x144 & ~x145 & ~x151 & ~x152 & ~x154 & ~x158 & ~x161 & ~x173 & ~x175 & ~x178 & ~x194 & ~x197 & ~x199 & ~x204 & ~x224 & ~x225 & ~x226 & ~x227 & ~x228 & ~x229 & ~x280 & ~x309 & ~x313 & ~x314 & ~x556 & ~x557 & ~x589 & ~x619 & ~x641 & ~x643 & ~x644 & ~x646 & ~x647 & ~x652 & ~x654 & ~x655 & ~x659 & ~x660 & ~x663 & ~x664 & ~x665 & ~x668 & ~x669 & ~x670 & ~x672 & ~x673 & ~x680 & ~x682 & ~x685 & ~x687 & ~x688 & ~x689 & ~x691 & ~x694 & ~x698 & ~x711 & ~x716 & ~x731 & ~x736 & ~x743 & ~x753 & ~x767 & ~x768 & ~x783;
assign c7288 =  x476 & ~x239 & ~x265;
assign c7290 = ~x2 & ~x10 & ~x32 & ~x34 & ~x39 & ~x40 & ~x44 & ~x48 & ~x49 & ~x50 & ~x56 & ~x70 & ~x71 & ~x73 & ~x75 & ~x76 & ~x99 & ~x107 & ~x111 & ~x113 & ~x115 & ~x116 & ~x125 & ~x132 & ~x134 & ~x141 & ~x146 & ~x147 & ~x148 & ~x160 & ~x163 & ~x179 & ~x187 & ~x194 & ~x200 & ~x202 & ~x207 & ~x216 & ~x219 & ~x221 & ~x228 & ~x232 & ~x235 & ~x254 & ~x272 & ~x301 & ~x307 & ~x315 & ~x316 & ~x337 & ~x482 & ~x483 & ~x629 & ~x648 & ~x673 & ~x691 & ~x710 & ~x739 & ~x745 & ~x762 & ~x766 & ~x770 & ~x777 & ~x780;
assign c7292 =  x157 &  x185 & ~x50 & ~x146;
assign c7294 =  x418 & ~x3 & ~x5 & ~x6 & ~x8 & ~x9 & ~x12 & ~x13 & ~x14 & ~x18 & ~x20 & ~x22 & ~x23 & ~x24 & ~x25 & ~x26 & ~x28 & ~x30 & ~x31 & ~x32 & ~x36 & ~x37 & ~x38 & ~x43 & ~x44 & ~x47 & ~x48 & ~x49 & ~x50 & ~x51 & ~x54 & ~x57 & ~x58 & ~x60 & ~x61 & ~x62 & ~x67 & ~x68 & ~x70 & ~x71 & ~x73 & ~x74 & ~x75 & ~x77 & ~x79 & ~x80 & ~x81 & ~x82 & ~x84 & ~x85 & ~x88 & ~x90 & ~x92 & ~x93 & ~x94 & ~x95 & ~x96 & ~x101 & ~x102 & ~x103 & ~x106 & ~x108 & ~x110 & ~x111 & ~x114 & ~x116 & ~x117 & ~x118 & ~x119 & ~x120 & ~x121 & ~x122 & ~x123 & ~x125 & ~x126 & ~x129 & ~x130 & ~x131 & ~x133 & ~x134 & ~x136 & ~x137 & ~x138 & ~x140 & ~x144 & ~x146 & ~x147 & ~x148 & ~x149 & ~x152 & ~x153 & ~x156 & ~x158 & ~x159 & ~x160 & ~x161 & ~x163 & ~x165 & ~x169 & ~x170 & ~x171 & ~x172 & ~x173 & ~x176 & ~x178 & ~x180 & ~x181 & ~x182 & ~x183 & ~x185 & ~x186 & ~x187 & ~x188 & ~x189 & ~x191 & ~x194 & ~x197 & ~x198 & ~x199 & ~x200 & ~x201 & ~x202 & ~x203 & ~x210 & ~x212 & ~x214 & ~x215 & ~x221 & ~x225 & ~x227 & ~x228 & ~x230 & ~x244 & ~x246 & ~x248 & ~x251 & ~x255 & ~x257 & ~x259 & ~x273 & ~x274 & ~x283 & ~x284 & ~x301 & ~x308 & ~x336 & ~x365 & ~x561 & ~x563 & ~x588 & ~x589 & ~x590 & ~x592 & ~x593 & ~x594 & ~x596 & ~x597 & ~x598 & ~x601 & ~x603 & ~x604 & ~x605 & ~x607 & ~x608 & ~x609 & ~x610 & ~x611 & ~x615 & ~x618 & ~x620 & ~x621 & ~x622 & ~x623 & ~x627 & ~x629 & ~x630 & ~x631 & ~x634 & ~x636 & ~x637 & ~x638 & ~x639 & ~x640 & ~x641 & ~x643 & ~x644 & ~x645 & ~x646 & ~x647 & ~x648 & ~x649 & ~x650 & ~x651 & ~x652 & ~x653 & ~x654 & ~x655 & ~x656 & ~x657 & ~x659 & ~x662 & ~x664 & ~x665 & ~x667 & ~x668 & ~x669 & ~x670 & ~x671 & ~x673 & ~x674 & ~x675 & ~x677 & ~x678 & ~x679 & ~x681 & ~x682 & ~x684 & ~x686 & ~x687 & ~x688 & ~x689 & ~x691 & ~x692 & ~x693 & ~x695 & ~x698 & ~x699 & ~x700 & ~x705 & ~x706 & ~x707 & ~x708 & ~x709 & ~x710 & ~x711 & ~x712 & ~x713 & ~x714 & ~x715 & ~x716 & ~x719 & ~x721 & ~x723 & ~x725 & ~x726 & ~x727 & ~x729 & ~x730 & ~x731 & ~x732 & ~x733 & ~x734 & ~x736 & ~x737 & ~x738 & ~x740 & ~x743 & ~x744 & ~x746 & ~x747 & ~x749 & ~x753 & ~x754 & ~x757 & ~x758 & ~x759 & ~x760 & ~x761 & ~x763 & ~x765 & ~x769 & ~x770 & ~x776 & ~x777 & ~x780 & ~x781 & ~x783;
assign c7296 = ~x8 & ~x12 & ~x13 & ~x15 & ~x17 & ~x24 & ~x31 & ~x32 & ~x38 & ~x39 & ~x40 & ~x59 & ~x63 & ~x66 & ~x80 & ~x81 & ~x84 & ~x96 & ~x118 & ~x119 & ~x128 & ~x130 & ~x143 & ~x144 & ~x149 & ~x154 & ~x160 & ~x172 & ~x175 & ~x177 & ~x179 & ~x195 & ~x199 & ~x209 & ~x280 & ~x289 & ~x314 & ~x340 & ~x425 & ~x426 & ~x455 & ~x613 & ~x615 & ~x617 & ~x651 & ~x658 & ~x671 & ~x673 & ~x683 & ~x687 & ~x692 & ~x709 & ~x710 & ~x711 & ~x715 & ~x719 & ~x720 & ~x731 & ~x733 & ~x735 & ~x753 & ~x755 & ~x767 & ~x779;
assign c7298 =  x297 &  x429 &  x606 & ~x22 & ~x26 & ~x27 & ~x55 & ~x59 & ~x71 & ~x96 & ~x164 & ~x174 & ~x191 & ~x197 & ~x235 & ~x237 & ~x676 & ~x684 & ~x721 & ~x751 & ~x752 & ~x773 & ~x778;
assign c7300 =  x295 &  x321 &  x346 & ~x0 & ~x12 & ~x13 & ~x16 & ~x24 & ~x25 & ~x26 & ~x27 & ~x30 & ~x36 & ~x37 & ~x39 & ~x40 & ~x42 & ~x48 & ~x49 & ~x52 & ~x55 & ~x60 & ~x61 & ~x63 & ~x66 & ~x67 & ~x71 & ~x74 & ~x76 & ~x77 & ~x79 & ~x82 & ~x83 & ~x84 & ~x88 & ~x90 & ~x91 & ~x92 & ~x96 & ~x100 & ~x101 & ~x110 & ~x111 & ~x113 & ~x115 & ~x119 & ~x122 & ~x126 & ~x127 & ~x128 & ~x130 & ~x139 & ~x140 & ~x146 & ~x150 & ~x152 & ~x154 & ~x155 & ~x168 & ~x170 & ~x171 & ~x175 & ~x179 & ~x180 & ~x188 & ~x203 & ~x206 & ~x216 & ~x223 & ~x225 & ~x229 & ~x231 & ~x234 & ~x235 & ~x244 & ~x245 & ~x258 & ~x259 & ~x281 & ~x283 & ~x309 & ~x314 & ~x337 & ~x364 & ~x563 & ~x589 & ~x609 & ~x610 & ~x612 & ~x616 & ~x620 & ~x644 & ~x646 & ~x647 & ~x649 & ~x652 & ~x660 & ~x665 & ~x669 & ~x670 & ~x671 & ~x677 & ~x678 & ~x680 & ~x686 & ~x687 & ~x688 & ~x693 & ~x699 & ~x701 & ~x702 & ~x703 & ~x704 & ~x705 & ~x706 & ~x707 & ~x709 & ~x711 & ~x714 & ~x716 & ~x718 & ~x719 & ~x721 & ~x723 & ~x725 & ~x730 & ~x735 & ~x737 & ~x740 & ~x751 & ~x752 & ~x757 & ~x758 & ~x766 & ~x769 & ~x770 & ~x773;
assign c7302 =  x332 &  x334 &  x362 &  x414 &  x418 &  x440 &  x578 & ~x6 & ~x82 & ~x116 & ~x227 & ~x316 & ~x422 & ~x643;
assign c7304 =  x390 &  x632 & ~x32;
assign c7306 =  x394 & ~x25 & ~x26 & ~x44 & ~x51 & ~x53 & ~x82 & ~x87 & ~x103 & ~x124 & ~x128 & ~x144 & ~x152 & ~x178 & ~x200 & ~x206 & ~x227 & ~x230 & ~x232 & ~x252 & ~x257 & ~x258 & ~x287 & ~x567 & ~x585 & ~x662 & ~x680 & ~x710 & ~x713;
assign c7308 =  x660 & ~x165 & ~x424;
assign c7310 =  x242 &  x520 &  x526 & ~x1 & ~x6 & ~x8 & ~x13 & ~x16 & ~x28 & ~x39 & ~x46 & ~x55 & ~x56 & ~x59 & ~x78 & ~x96 & ~x108 & ~x140 & ~x173 & ~x174 & ~x191 & ~x198 & ~x223 & ~x254 & ~x288 & ~x289 & ~x310 & ~x344 & ~x399 & ~x452 & ~x697 & ~x713 & ~x775 & ~x777 & ~x782;
assign c7312 = ~x183 & ~x486 & ~x510 & ~x511 & ~x584;
assign c7314 =  x187 &  x333 & ~x0 & ~x7 & ~x22 & ~x46 & ~x69 & ~x110 & ~x288 & ~x669 & ~x695 & ~x706 & ~x714 & ~x718 & ~x764;
assign c7316 =  x577 &  x578 & ~x1 & ~x4 & ~x6 & ~x19 & ~x22 & ~x23 & ~x32 & ~x34 & ~x38 & ~x47 & ~x48 & ~x49 & ~x51 & ~x54 & ~x56 & ~x58 & ~x59 & ~x64 & ~x65 & ~x72 & ~x88 & ~x91 & ~x102 & ~x104 & ~x109 & ~x112 & ~x121 & ~x123 & ~x124 & ~x126 & ~x128 & ~x136 & ~x138 & ~x139 & ~x141 & ~x146 & ~x151 & ~x152 & ~x153 & ~x162 & ~x165 & ~x183 & ~x189 & ~x193 & ~x197 & ~x202 & ~x204 & ~x224 & ~x225 & ~x228 & ~x233 & ~x234 & ~x257 & ~x259 & ~x280 & ~x281 & ~x287 & ~x288 & ~x337 & ~x338 & ~x341 & ~x343 & ~x365 & ~x392 & ~x393 & ~x394 & ~x420 & ~x560 & ~x561 & ~x616 & ~x620 & ~x621 & ~x638 & ~x644 & ~x652 & ~x657 & ~x664 & ~x667 & ~x671 & ~x672 & ~x675 & ~x677 & ~x680 & ~x681 & ~x683 & ~x692 & ~x693 & ~x695 & ~x709 & ~x716 & ~x719 & ~x722 & ~x723 & ~x726 & ~x732 & ~x734 & ~x743 & ~x759 & ~x764 & ~x778 & ~x779;
assign c7318 =  x297 &  x349 &  x458 & ~x0 & ~x1 & ~x9 & ~x14 & ~x23 & ~x26 & ~x28 & ~x29 & ~x31 & ~x43 & ~x45 & ~x52 & ~x55 & ~x59 & ~x61 & ~x62 & ~x63 & ~x66 & ~x70 & ~x72 & ~x80 & ~x81 & ~x82 & ~x84 & ~x86 & ~x92 & ~x95 & ~x109 & ~x112 & ~x113 & ~x117 & ~x121 & ~x122 & ~x140 & ~x171 & ~x172 & ~x196 & ~x223 & ~x226 & ~x227 & ~x232 & ~x233 & ~x235 & ~x256 & ~x260 & ~x279 & ~x281 & ~x310 & ~x340 & ~x341 & ~x342 & ~x365 & ~x369 & ~x393 & ~x448 & ~x587 & ~x613 & ~x614 & ~x616 & ~x635 & ~x640 & ~x671 & ~x699 & ~x701 & ~x714 & ~x719 & ~x725 & ~x736 & ~x755 & ~x756 & ~x760 & ~x761 & ~x762 & ~x765 & ~x768 & ~x772 & ~x773 & ~x775 & ~x776 & ~x777 & ~x783;
assign c7320 =  x662;
assign c7322 =  x333 &  x462 & ~x1 & ~x2 & ~x3 & ~x4 & ~x5 & ~x7 & ~x9 & ~x10 & ~x11 & ~x12 & ~x14 & ~x15 & ~x16 & ~x19 & ~x23 & ~x24 & ~x25 & ~x27 & ~x28 & ~x30 & ~x31 & ~x32 & ~x33 & ~x34 & ~x35 & ~x36 & ~x38 & ~x39 & ~x41 & ~x42 & ~x43 & ~x45 & ~x48 & ~x50 & ~x51 & ~x52 & ~x53 & ~x55 & ~x56 & ~x62 & ~x63 & ~x64 & ~x65 & ~x68 & ~x71 & ~x72 & ~x73 & ~x74 & ~x76 & ~x77 & ~x78 & ~x79 & ~x80 & ~x81 & ~x84 & ~x87 & ~x89 & ~x90 & ~x91 & ~x92 & ~x93 & ~x94 & ~x95 & ~x96 & ~x97 & ~x103 & ~x104 & ~x105 & ~x106 & ~x108 & ~x109 & ~x111 & ~x113 & ~x114 & ~x115 & ~x116 & ~x117 & ~x132 & ~x134 & ~x135 & ~x136 & ~x137 & ~x138 & ~x142 & ~x144 & ~x146 & ~x147 & ~x148 & ~x150 & ~x151 & ~x152 & ~x153 & ~x169 & ~x171 & ~x173 & ~x174 & ~x175 & ~x176 & ~x178 & ~x195 & ~x198 & ~x199 & ~x200 & ~x201 & ~x202 & ~x203 & ~x205 & ~x207 & ~x223 & ~x224 & ~x225 & ~x226 & ~x227 & ~x228 & ~x229 & ~x230 & ~x234 & ~x236 & ~x252 & ~x253 & ~x254 & ~x255 & ~x256 & ~x257 & ~x261 & ~x279 & ~x281 & ~x283 & ~x284 & ~x285 & ~x286 & ~x288 & ~x308 & ~x309 & ~x310 & ~x311 & ~x312 & ~x314 & ~x315 & ~x335 & ~x337 & ~x339 & ~x341 & ~x364 & ~x365 & ~x367 & ~x392 & ~x537 & ~x616 & ~x618 & ~x644 & ~x647 & ~x669 & ~x670 & ~x671 & ~x673 & ~x674 & ~x675 & ~x677 & ~x678 & ~x681 & ~x682 & ~x684 & ~x688 & ~x691 & ~x692 & ~x697 & ~x698 & ~x699 & ~x700 & ~x701 & ~x704 & ~x705 & ~x706 & ~x707 & ~x708 & ~x709 & ~x710 & ~x712 & ~x713 & ~x714 & ~x715 & ~x716 & ~x720 & ~x722 & ~x723 & ~x724 & ~x725 & ~x726 & ~x727 & ~x729 & ~x730 & ~x731 & ~x732 & ~x735 & ~x736 & ~x737 & ~x738 & ~x740 & ~x742 & ~x743 & ~x744 & ~x746 & ~x747 & ~x748 & ~x749 & ~x750 & ~x751 & ~x752 & ~x753 & ~x754 & ~x755 & ~x759 & ~x763 & ~x764 & ~x765 & ~x766 & ~x767 & ~x768 & ~x769 & ~x772 & ~x773 & ~x776 & ~x778 & ~x779 & ~x780 & ~x782;
assign c7324 =  x382 &  x413 & ~x0 & ~x6 & ~x7 & ~x9 & ~x10 & ~x14 & ~x18 & ~x20 & ~x22 & ~x24 & ~x28 & ~x30 & ~x32 & ~x35 & ~x39 & ~x42 & ~x51 & ~x54 & ~x56 & ~x60 & ~x67 & ~x71 & ~x85 & ~x86 & ~x88 & ~x90 & ~x92 & ~x99 & ~x104 & ~x105 & ~x106 & ~x108 & ~x110 & ~x111 & ~x114 & ~x116 & ~x117 & ~x119 & ~x120 & ~x131 & ~x133 & ~x139 & ~x145 & ~x150 & ~x151 & ~x167 & ~x170 & ~x172 & ~x173 & ~x198 & ~x201 & ~x202 & ~x203 & ~x205 & ~x223 & ~x225 & ~x226 & ~x229 & ~x253 & ~x254 & ~x284 & ~x285 & ~x313 & ~x524 & ~x526 & ~x590 & ~x615 & ~x619 & ~x620 & ~x635 & ~x636 & ~x640 & ~x641 & ~x649 & ~x652 & ~x653 & ~x660 & ~x662 & ~x666 & ~x668 & ~x669 & ~x674 & ~x681 & ~x684 & ~x686 & ~x690 & ~x696 & ~x697 & ~x699 & ~x703 & ~x705 & ~x713 & ~x720 & ~x721 & ~x722 & ~x723 & ~x725 & ~x730 & ~x733 & ~x736 & ~x738 & ~x744 & ~x745 & ~x746 & ~x756 & ~x757 & ~x759 & ~x767 & ~x770 & ~x774 & ~x779 & ~x780;
assign c7326 = ~x1 & ~x4 & ~x12 & ~x14 & ~x16 & ~x17 & ~x19 & ~x23 & ~x27 & ~x29 & ~x33 & ~x37 & ~x38 & ~x46 & ~x53 & ~x55 & ~x56 & ~x69 & ~x70 & ~x72 & ~x73 & ~x75 & ~x76 & ~x78 & ~x80 & ~x81 & ~x82 & ~x83 & ~x84 & ~x86 & ~x92 & ~x96 & ~x98 & ~x100 & ~x104 & ~x110 & ~x112 & ~x115 & ~x117 & ~x120 & ~x121 & ~x125 & ~x129 & ~x132 & ~x135 & ~x136 & ~x137 & ~x138 & ~x139 & ~x147 & ~x153 & ~x155 & ~x166 & ~x167 & ~x169 & ~x171 & ~x173 & ~x176 & ~x180 & ~x181 & ~x191 & ~x195 & ~x196 & ~x197 & ~x200 & ~x206 & ~x207 & ~x209 & ~x224 & ~x226 & ~x228 & ~x229 & ~x230 & ~x252 & ~x253 & ~x254 & ~x256 & ~x258 & ~x261 & ~x262 & ~x280 & ~x282 & ~x289 & ~x290 & ~x291 & ~x313 & ~x316 & ~x336 & ~x338 & ~x339 & ~x340 & ~x341 & ~x344 & ~x346 & ~x347 & ~x364 & ~x367 & ~x368 & ~x370 & ~x371 & ~x373 & ~x396 & ~x397 & ~x399 & ~x425 & ~x426 & ~x534 & ~x618 & ~x643 & ~x644 & ~x647 & ~x652 & ~x661 & ~x662 & ~x664 & ~x669 & ~x670 & ~x673 & ~x674 & ~x679 & ~x681 & ~x683 & ~x684 & ~x685 & ~x687 & ~x692 & ~x693 & ~x694 & ~x696 & ~x697 & ~x699 & ~x704 & ~x706 & ~x708 & ~x709 & ~x710 & ~x712 & ~x714 & ~x715 & ~x719 & ~x722 & ~x724 & ~x727 & ~x737 & ~x738 & ~x741 & ~x742 & ~x745 & ~x747 & ~x751 & ~x758 & ~x759 & ~x761 & ~x763 & ~x767 & ~x769 & ~x770 & ~x771 & ~x772 & ~x774 & ~x780;
assign c7328 =  x750;
assign c7330 =  x634 & ~x17 & ~x20 & ~x56 & ~x61 & ~x67 & ~x70 & ~x85 & ~x137 & ~x143 & ~x154 & ~x162 & ~x181 & ~x191 & ~x199 & ~x200 & ~x232 & ~x261 & ~x286 & ~x339 & ~x368 & ~x743 & ~x744 & ~x758 & ~x765;
assign c7332 = ~x5 & ~x42 & ~x44 & ~x55 & ~x64 & ~x72 & ~x76 & ~x83 & ~x86 & ~x99 & ~x104 & ~x107 & ~x110 & ~x118 & ~x131 & ~x138 & ~x141 & ~x153 & ~x161 & ~x162 & ~x193 & ~x197 & ~x204 & ~x214 & ~x216 & ~x221 & ~x238 & ~x280 & ~x301 & ~x327 & ~x328 & ~x465 & ~x658 & ~x673 & ~x678 & ~x679 & ~x681 & ~x682 & ~x710 & ~x719 & ~x741 & ~x745 & ~x754 & ~x768 & ~x770;
assign c7334 =  x362 & ~x3 & ~x5 & ~x6 & ~x9 & ~x11 & ~x13 & ~x17 & ~x20 & ~x26 & ~x33 & ~x36 & ~x42 & ~x44 & ~x49 & ~x62 & ~x63 & ~x65 & ~x68 & ~x72 & ~x73 & ~x74 & ~x75 & ~x78 & ~x84 & ~x85 & ~x87 & ~x96 & ~x97 & ~x104 & ~x105 & ~x109 & ~x117 & ~x118 & ~x123 & ~x126 & ~x127 & ~x131 & ~x139 & ~x143 & ~x145 & ~x146 & ~x148 & ~x149 & ~x155 & ~x165 & ~x172 & ~x175 & ~x176 & ~x177 & ~x181 & ~x183 & ~x198 & ~x201 & ~x203 & ~x204 & ~x205 & ~x206 & ~x208 & ~x224 & ~x225 & ~x226 & ~x229 & ~x230 & ~x232 & ~x235 & ~x251 & ~x252 & ~x254 & ~x256 & ~x258 & ~x284 & ~x286 & ~x307 & ~x364 & ~x505 & ~x534 & ~x561 & ~x590 & ~x591 & ~x592 & ~x595 & ~x601 & ~x602 & ~x629 & ~x632 & ~x639 & ~x641 & ~x642 & ~x643 & ~x651 & ~x655 & ~x658 & ~x662 & ~x665 & ~x666 & ~x668 & ~x670 & ~x682 & ~x685 & ~x687 & ~x689 & ~x696 & ~x701 & ~x704 & ~x705 & ~x714 & ~x716 & ~x719 & ~x720 & ~x723 & ~x726 & ~x727 & ~x729 & ~x730 & ~x731 & ~x735 & ~x736 & ~x738 & ~x739 & ~x744 & ~x745 & ~x746 & ~x747 & ~x749 & ~x751 & ~x757 & ~x758 & ~x759 & ~x765 & ~x766 & ~x767 & ~x768 & ~x773 & ~x774 & ~x776 & ~x780;
assign c7336 = ~x16 & ~x18 & ~x20 & ~x32 & ~x49 & ~x50 & ~x52 & ~x58 & ~x62 & ~x67 & ~x68 & ~x78 & ~x82 & ~x83 & ~x92 & ~x94 & ~x111 & ~x131 & ~x141 & ~x142 & ~x143 & ~x145 & ~x150 & ~x151 & ~x153 & ~x160 & ~x162 & ~x166 & ~x167 & ~x171 & ~x176 & ~x178 & ~x179 & ~x187 & ~x190 & ~x191 & ~x197 & ~x198 & ~x206 & ~x210 & ~x219 & ~x220 & ~x221 & ~x223 & ~x226 & ~x229 & ~x245 & ~x252 & ~x260 & ~x263 & ~x272 & ~x274 & ~x280 & ~x285 & ~x287 & ~x291 & ~x300 & ~x312 & ~x328 & ~x337 & ~x364 & ~x367 & ~x369 & ~x397 & ~x645 & ~x646 & ~x649 & ~x659 & ~x664 & ~x681 & ~x687 & ~x701 & ~x706 & ~x707 & ~x716 & ~x724 & ~x730 & ~x736 & ~x738 & ~x745 & ~x750 & ~x753 & ~x754 & ~x755 & ~x761 & ~x765 & ~x769 & ~x775 & ~x781;
assign c7338 =  x350 &  x351 &  x375 &  x376 &  x401 &  x445 & ~x4 & ~x10 & ~x15 & ~x16 & ~x19 & ~x27 & ~x35 & ~x36 & ~x37 & ~x38 & ~x39 & ~x41 & ~x47 & ~x50 & ~x54 & ~x56 & ~x60 & ~x61 & ~x65 & ~x67 & ~x71 & ~x73 & ~x76 & ~x83 & ~x85 & ~x87 & ~x89 & ~x90 & ~x92 & ~x96 & ~x99 & ~x101 & ~x106 & ~x108 & ~x121 & ~x122 & ~x124 & ~x125 & ~x131 & ~x132 & ~x136 & ~x140 & ~x142 & ~x149 & ~x150 & ~x151 & ~x154 & ~x161 & ~x168 & ~x169 & ~x170 & ~x171 & ~x172 & ~x175 & ~x186 & ~x189 & ~x200 & ~x202 & ~x203 & ~x204 & ~x223 & ~x228 & ~x230 & ~x233 & ~x244 & ~x254 & ~x256 & ~x259 & ~x260 & ~x261 & ~x280 & ~x288 & ~x289 & ~x308 & ~x364 & ~x561 & ~x588 & ~x591 & ~x593 & ~x617 & ~x618 & ~x621 & ~x623 & ~x646 & ~x648 & ~x651 & ~x652 & ~x653 & ~x656 & ~x659 & ~x660 & ~x661 & ~x663 & ~x664 & ~x665 & ~x667 & ~x668 & ~x676 & ~x684 & ~x685 & ~x687 & ~x688 & ~x691 & ~x698 & ~x702 & ~x705 & ~x710 & ~x711 & ~x712 & ~x713 & ~x716 & ~x719 & ~x720 & ~x724 & ~x725 & ~x727 & ~x729 & ~x732 & ~x738 & ~x744 & ~x747 & ~x750 & ~x769 & ~x770 & ~x771 & ~x772 & ~x774 & ~x777 & ~x778 & ~x780;
assign c7340 =  x418 & ~x2 & ~x7 & ~x8 & ~x13 & ~x14 & ~x16 & ~x36 & ~x41 & ~x51 & ~x57 & ~x61 & ~x62 & ~x63 & ~x67 & ~x84 & ~x94 & ~x95 & ~x104 & ~x107 & ~x108 & ~x111 & ~x119 & ~x123 & ~x126 & ~x127 & ~x131 & ~x132 & ~x133 & ~x141 & ~x142 & ~x145 & ~x151 & ~x156 & ~x159 & ~x161 & ~x165 & ~x166 & ~x172 & ~x177 & ~x188 & ~x193 & ~x194 & ~x200 & ~x202 & ~x218 & ~x219 & ~x221 & ~x246 & ~x259 & ~x274 & ~x276 & ~x280 & ~x281 & ~x302 & ~x308 & ~x309 & ~x310 & ~x337 & ~x364 & ~x392 & ~x621 & ~x645 & ~x653 & ~x664 & ~x675 & ~x677 & ~x678 & ~x696 & ~x722 & ~x730 & ~x731 & ~x744 & ~x754 & ~x762 & ~x772 & ~x774 & ~x777 & ~x779;
assign c7342 =  x319 &  x321 &  x345 &  x357 & ~x0 & ~x3 & ~x5 & ~x8 & ~x9 & ~x15 & ~x18 & ~x19 & ~x20 & ~x25 & ~x26 & ~x29 & ~x30 & ~x31 & ~x34 & ~x35 & ~x36 & ~x41 & ~x46 & ~x49 & ~x51 & ~x53 & ~x54 & ~x58 & ~x60 & ~x61 & ~x63 & ~x66 & ~x68 & ~x69 & ~x71 & ~x76 & ~x78 & ~x79 & ~x82 & ~x84 & ~x95 & ~x97 & ~x99 & ~x101 & ~x104 & ~x107 & ~x110 & ~x115 & ~x117 & ~x119 & ~x120 & ~x123 & ~x127 & ~x128 & ~x132 & ~x133 & ~x134 & ~x135 & ~x139 & ~x141 & ~x142 & ~x146 & ~x149 & ~x152 & ~x154 & ~x155 & ~x161 & ~x167 & ~x168 & ~x170 & ~x171 & ~x173 & ~x175 & ~x176 & ~x181 & ~x197 & ~x199 & ~x200 & ~x204 & ~x206 & ~x225 & ~x226 & ~x229 & ~x230 & ~x231 & ~x234 & ~x252 & ~x254 & ~x257 & ~x258 & ~x259 & ~x281 & ~x285 & ~x313 & ~x336 & ~x337 & ~x364 & ~x588 & ~x589 & ~x616 & ~x639 & ~x643 & ~x644 & ~x645 & ~x647 & ~x648 & ~x652 & ~x656 & ~x659 & ~x664 & ~x665 & ~x666 & ~x670 & ~x676 & ~x678 & ~x679 & ~x681 & ~x683 & ~x684 & ~x686 & ~x687 & ~x688 & ~x690 & ~x693 & ~x700 & ~x702 & ~x705 & ~x709 & ~x713 & ~x719 & ~x720 & ~x722 & ~x725 & ~x726 & ~x728 & ~x730 & ~x731 & ~x732 & ~x739 & ~x742 & ~x743 & ~x744 & ~x746 & ~x747 & ~x749 & ~x750 & ~x751 & ~x752 & ~x755 & ~x757 & ~x761 & ~x763 & ~x766 & ~x771 & ~x775 & ~x781 & ~x783;
assign c7344 = ~x5 & ~x27 & ~x40 & ~x49 & ~x53 & ~x67 & ~x69 & ~x73 & ~x106 & ~x125 & ~x126 & ~x128 & ~x134 & ~x146 & ~x163 & ~x189 & ~x195 & ~x205 & ~x228 & ~x245 & ~x246 & ~x252 & ~x279 & ~x300 & ~x359 & ~x365 & ~x637 & ~x662 & ~x665 & ~x675 & ~x679 & ~x687 & ~x695 & ~x701 & ~x707 & ~x715 & ~x738 & ~x753;
assign c7346 =  x242 &  x271 &  x326 &  x354 & ~x2 & ~x3 & ~x6 & ~x12 & ~x16 & ~x21 & ~x22 & ~x27 & ~x31 & ~x35 & ~x42 & ~x48 & ~x50 & ~x57 & ~x60 & ~x83 & ~x86 & ~x91 & ~x94 & ~x99 & ~x103 & ~x107 & ~x125 & ~x137 & ~x143 & ~x146 & ~x170 & ~x172 & ~x174 & ~x189 & ~x190 & ~x218 & ~x227 & ~x234 & ~x235 & ~x236 & ~x248 & ~x291 & ~x308 & ~x310 & ~x311 & ~x314 & ~x316 & ~x317 & ~x339 & ~x343 & ~x676 & ~x678 & ~x693 & ~x694 & ~x703 & ~x706 & ~x707 & ~x708 & ~x713 & ~x715 & ~x716 & ~x720 & ~x725 & ~x732 & ~x735 & ~x738 & ~x752 & ~x760 & ~x761 & ~x765 & ~x768 & ~x776 & ~x779;
assign c7348 =  x297 &  x348 &  x381 & ~x1 & ~x4 & ~x8 & ~x9 & ~x13 & ~x18 & ~x19 & ~x20 & ~x23 & ~x24 & ~x25 & ~x26 & ~x30 & ~x32 & ~x35 & ~x36 & ~x40 & ~x44 & ~x48 & ~x52 & ~x55 & ~x59 & ~x61 & ~x65 & ~x68 & ~x70 & ~x73 & ~x75 & ~x76 & ~x78 & ~x79 & ~x80 & ~x81 & ~x82 & ~x83 & ~x91 & ~x94 & ~x100 & ~x102 & ~x108 & ~x111 & ~x113 & ~x119 & ~x120 & ~x126 & ~x127 & ~x128 & ~x130 & ~x136 & ~x142 & ~x151 & ~x152 & ~x153 & ~x154 & ~x157 & ~x158 & ~x160 & ~x163 & ~x165 & ~x173 & ~x174 & ~x175 & ~x176 & ~x180 & ~x182 & ~x184 & ~x195 & ~x201 & ~x205 & ~x206 & ~x209 & ~x224 & ~x226 & ~x230 & ~x253 & ~x255 & ~x274 & ~x280 & ~x283 & ~x286 & ~x287 & ~x313 & ~x616 & ~x645 & ~x646 & ~x648 & ~x653 & ~x666 & ~x667 & ~x670 & ~x678 & ~x680 & ~x681 & ~x685 & ~x686 & ~x688 & ~x689 & ~x691 & ~x694 & ~x698 & ~x699 & ~x701 & ~x702 & ~x704 & ~x710 & ~x712 & ~x722 & ~x726 & ~x740 & ~x744 & ~x755 & ~x757 & ~x759 & ~x761 & ~x766 & ~x771 & ~x775 & ~x776 & ~x777 & ~x778 & ~x782;
assign c7350 =  x320 &  x396 &  x398 & ~x4 & ~x8 & ~x29 & ~x35 & ~x48 & ~x53 & ~x63 & ~x71 & ~x78 & ~x86 & ~x87 & ~x113 & ~x116 & ~x119 & ~x127 & ~x131 & ~x133 & ~x135 & ~x136 & ~x138 & ~x153 & ~x165 & ~x169 & ~x204 & ~x209 & ~x218 & ~x227 & ~x233 & ~x244 & ~x245 & ~x252 & ~x254 & ~x259 & ~x335 & ~x619 & ~x621 & ~x644 & ~x647 & ~x655 & ~x656 & ~x675 & ~x682 & ~x689 & ~x699 & ~x709 & ~x710 & ~x715 & ~x742 & ~x755 & ~x762 & ~x764 & ~x772 & ~x782;
assign c7352 =  x645;
assign c7354 =  x605 &  x606 & ~x641 & ~x642 & ~x757;
assign c7356 =  x68;
assign c7358 =  x417 &  x444 &  x445 & ~x0 & ~x1 & ~x2 & ~x4 & ~x5 & ~x6 & ~x9 & ~x15 & ~x17 & ~x19 & ~x22 & ~x26 & ~x28 & ~x29 & ~x30 & ~x31 & ~x34 & ~x35 & ~x36 & ~x41 & ~x44 & ~x50 & ~x52 & ~x54 & ~x56 & ~x62 & ~x63 & ~x64 & ~x65 & ~x67 & ~x69 & ~x70 & ~x73 & ~x74 & ~x76 & ~x79 & ~x81 & ~x87 & ~x89 & ~x92 & ~x94 & ~x95 & ~x98 & ~x100 & ~x103 & ~x107 & ~x110 & ~x111 & ~x112 & ~x118 & ~x119 & ~x123 & ~x128 & ~x130 & ~x132 & ~x134 & ~x135 & ~x136 & ~x137 & ~x141 & ~x143 & ~x149 & ~x151 & ~x154 & ~x159 & ~x163 & ~x165 & ~x173 & ~x175 & ~x177 & ~x179 & ~x180 & ~x181 & ~x187 & ~x189 & ~x192 & ~x193 & ~x194 & ~x195 & ~x196 & ~x200 & ~x202 & ~x204 & ~x217 & ~x218 & ~x220 & ~x227 & ~x229 & ~x245 & ~x246 & ~x247 & ~x252 & ~x254 & ~x255 & ~x256 & ~x259 & ~x273 & ~x274 & ~x281 & ~x282 & ~x284 & ~x301 & ~x307 & ~x309 & ~x312 & ~x337 & ~x364 & ~x365 & ~x392 & ~x617 & ~x618 & ~x619 & ~x643 & ~x648 & ~x650 & ~x651 & ~x653 & ~x658 & ~x659 & ~x665 & ~x675 & ~x681 & ~x684 & ~x685 & ~x686 & ~x687 & ~x690 & ~x691 & ~x693 & ~x694 & ~x695 & ~x699 & ~x701 & ~x703 & ~x708 & ~x709 & ~x710 & ~x711 & ~x712 & ~x713 & ~x714 & ~x715 & ~x716 & ~x717 & ~x719 & ~x720 & ~x726 & ~x728 & ~x730 & ~x732 & ~x737 & ~x741 & ~x742 & ~x743 & ~x745 & ~x746 & ~x747 & ~x749 & ~x752 & ~x754 & ~x757 & ~x758 & ~x759 & ~x760 & ~x764 & ~x767 & ~x773 & ~x774 & ~x779 & ~x781;
assign c7360 =  x444 &  x470 & ~x6 & ~x7 & ~x9 & ~x18 & ~x20 & ~x21 & ~x27 & ~x29 & ~x30 & ~x31 & ~x33 & ~x44 & ~x45 & ~x46 & ~x47 & ~x49 & ~x50 & ~x51 & ~x52 & ~x53 & ~x55 & ~x57 & ~x60 & ~x62 & ~x68 & ~x69 & ~x70 & ~x71 & ~x75 & ~x78 & ~x79 & ~x80 & ~x81 & ~x87 & ~x89 & ~x92 & ~x93 & ~x94 & ~x96 & ~x97 & ~x101 & ~x107 & ~x108 & ~x113 & ~x116 & ~x122 & ~x123 & ~x135 & ~x136 & ~x140 & ~x142 & ~x143 & ~x144 & ~x145 & ~x150 & ~x153 & ~x158 & ~x160 & ~x162 & ~x164 & ~x165 & ~x171 & ~x176 & ~x177 & ~x178 & ~x180 & ~x181 & ~x189 & ~x190 & ~x192 & ~x193 & ~x194 & ~x197 & ~x199 & ~x202 & ~x204 & ~x205 & ~x218 & ~x219 & ~x220 & ~x223 & ~x225 & ~x226 & ~x229 & ~x232 & ~x249 & ~x251 & ~x259 & ~x272 & ~x281 & ~x300 & ~x301 & ~x308 & ~x336 & ~x392 & ~x560 & ~x585 & ~x587 & ~x593 & ~x595 & ~x597 & ~x598 & ~x600 & ~x601 & ~x606 & ~x609 & ~x610 & ~x612 & ~x618 & ~x626 & ~x630 & ~x636 & ~x644 & ~x646 & ~x647 & ~x648 & ~x649 & ~x653 & ~x661 & ~x662 & ~x664 & ~x667 & ~x672 & ~x673 & ~x674 & ~x677 & ~x678 & ~x682 & ~x683 & ~x686 & ~x689 & ~x690 & ~x691 & ~x695 & ~x696 & ~x697 & ~x698 & ~x699 & ~x701 & ~x702 & ~x708 & ~x709 & ~x710 & ~x716 & ~x719 & ~x720 & ~x722 & ~x723 & ~x724 & ~x726 & ~x727 & ~x729 & ~x730 & ~x731 & ~x732 & ~x734 & ~x737 & ~x738 & ~x743 & ~x754 & ~x755 & ~x756 & ~x759 & ~x760 & ~x764 & ~x770 & ~x774 & ~x783;
assign c7362 =  x406 &  x492 &  x494 &  x521 & ~x0 & ~x2 & ~x5 & ~x12 & ~x15 & ~x21 & ~x25 & ~x30 & ~x34 & ~x36 & ~x37 & ~x40 & ~x41 & ~x42 & ~x43 & ~x49 & ~x50 & ~x57 & ~x64 & ~x76 & ~x77 & ~x89 & ~x96 & ~x99 & ~x103 & ~x104 & ~x106 & ~x107 & ~x111 & ~x114 & ~x115 & ~x139 & ~x140 & ~x142 & ~x145 & ~x146 & ~x148 & ~x170 & ~x174 & ~x175 & ~x200 & ~x202 & ~x205 & ~x206 & ~x226 & ~x227 & ~x228 & ~x230 & ~x253 & ~x257 & ~x308 & ~x314 & ~x556 & ~x557 & ~x588 & ~x613 & ~x615 & ~x635 & ~x636 & ~x639 & ~x640 & ~x643 & ~x644 & ~x662 & ~x666 & ~x668 & ~x672 & ~x678 & ~x690 & ~x691 & ~x693 & ~x694 & ~x696 & ~x700 & ~x704 & ~x708 & ~x711 & ~x716 & ~x717 & ~x718 & ~x720 & ~x722 & ~x723 & ~x726 & ~x731 & ~x733 & ~x735 & ~x739 & ~x740 & ~x741 & ~x744 & ~x757 & ~x758 & ~x760 & ~x761 & ~x764 & ~x766 & ~x768 & ~x769 & ~x773 & ~x774 & ~x775 & ~x777 & ~x778;
assign c7364 = ~x1 & ~x5 & ~x15 & ~x18 & ~x24 & ~x38 & ~x66 & ~x68 & ~x69 & ~x74 & ~x76 & ~x94 & ~x99 & ~x111 & ~x115 & ~x120 & ~x122 & ~x147 & ~x149 & ~x150 & ~x179 & ~x204 & ~x219 & ~x221 & ~x226 & ~x231 & ~x234 & ~x252 & ~x253 & ~x254 & ~x259 & ~x261 & ~x280 & ~x289 & ~x291 & ~x344 & ~x365 & ~x370 & ~x393 & ~x395 & ~x398 & ~x399 & ~x425 & ~x451 & ~x655 & ~x663 & ~x665 & ~x666 & ~x689 & ~x702 & ~x715 & ~x725 & ~x729 & ~x741 & ~x744 & ~x760 & ~x773 & ~x783;
assign c7366 =  x388 &  x444 &  x461 & ~x0 & ~x7 & ~x8 & ~x11 & ~x16 & ~x18 & ~x24 & ~x26 & ~x27 & ~x29 & ~x34 & ~x36 & ~x37 & ~x42 & ~x53 & ~x54 & ~x56 & ~x58 & ~x62 & ~x66 & ~x69 & ~x71 & ~x75 & ~x82 & ~x84 & ~x90 & ~x93 & ~x95 & ~x101 & ~x108 & ~x109 & ~x110 & ~x111 & ~x114 & ~x117 & ~x120 & ~x134 & ~x138 & ~x140 & ~x141 & ~x149 & ~x151 & ~x175 & ~x177 & ~x179 & ~x183 & ~x197 & ~x207 & ~x227 & ~x230 & ~x231 & ~x252 & ~x254 & ~x255 & ~x283 & ~x285 & ~x311 & ~x314 & ~x315 & ~x364 & ~x526 & ~x617 & ~x644 & ~x649 & ~x650 & ~x667 & ~x668 & ~x670 & ~x679 & ~x680 & ~x686 & ~x691 & ~x693 & ~x697 & ~x706 & ~x707 & ~x708 & ~x709 & ~x715 & ~x717 & ~x718 & ~x720 & ~x721 & ~x726 & ~x728 & ~x729 & ~x738 & ~x739 & ~x754 & ~x759 & ~x761 & ~x764 & ~x767 & ~x781;
assign c7368 =  x186 &  x353 &  x417 &  x472 & ~x20 & ~x47 & ~x106 & ~x116 & ~x167 & ~x194 & ~x224 & ~x532 & ~x560;
assign c7370 =  x590 &  x606 & ~x643;
assign c7372 =  x298 & ~x9 & ~x21 & ~x33 & ~x42 & ~x48 & ~x52 & ~x64 & ~x73 & ~x82 & ~x99 & ~x101 & ~x104 & ~x108 & ~x137 & ~x150 & ~x154 & ~x161 & ~x172 & ~x175 & ~x181 & ~x184 & ~x194 & ~x195 & ~x219 & ~x221 & ~x229 & ~x232 & ~x235 & ~x267 & ~x282 & ~x284 & ~x287 & ~x289 & ~x290 & ~x308 & ~x314 & ~x315 & ~x316 & ~x342 & ~x364 & ~x369 & ~x370 & ~x647 & ~x648 & ~x672 & ~x685 & ~x695 & ~x700 & ~x703 & ~x707 & ~x708 & ~x719 & ~x726 & ~x734 & ~x736 & ~x737 & ~x742 & ~x754 & ~x758 & ~x760 & ~x766 & ~x773 & ~x777;
assign c7374 =  x633 & ~x43 & ~x45 & ~x47 & ~x66 & ~x106 & ~x109 & ~x163 & ~x165 & ~x207 & ~x229 & ~x254 & ~x476 & ~x745 & ~x777;
assign c7376 =  x277 &  x390 &  x526 & ~x22 & ~x30 & ~x46 & ~x60 & ~x84 & ~x88 & ~x281 & ~x310 & ~x505;
assign c7378 = ~x5 & ~x8 & ~x21 & ~x22 & ~x24 & ~x43 & ~x54 & ~x74 & ~x75 & ~x76 & ~x77 & ~x83 & ~x85 & ~x92 & ~x93 & ~x96 & ~x138 & ~x154 & ~x172 & ~x195 & ~x197 & ~x198 & ~x206 & ~x207 & ~x230 & ~x232 & ~x236 & ~x238 & ~x252 & ~x253 & ~x261 & ~x264 & ~x281 & ~x291 & ~x293 & ~x314 & ~x316 & ~x318 & ~x322 & ~x347 & ~x365 & ~x372 & ~x373 & ~x398 & ~x424 & ~x643 & ~x695 & ~x708 & ~x724 & ~x726 & ~x736 & ~x743 & ~x746 & ~x747 & ~x750 & ~x752;
assign c7380 =  x382 &  x435 &  x443 & ~x9 & ~x11 & ~x13 & ~x38 & ~x57 & ~x58 & ~x60 & ~x62 & ~x70 & ~x78 & ~x109 & ~x117 & ~x123 & ~x140 & ~x152 & ~x169 & ~x181 & ~x207 & ~x219 & ~x227 & ~x228 & ~x238 & ~x256 & ~x259 & ~x284 & ~x285 & ~x293 & ~x370 & ~x394 & ~x420 & ~x475 & ~x709 & ~x716 & ~x732 & ~x747 & ~x752 & ~x783;
assign c7382 =  x104;
assign c7384 =  x130;
assign c7386 =  x319 &  x320 &  x345 &  x372 & ~x8 & ~x19 & ~x35 & ~x49 & ~x52 & ~x58 & ~x60 & ~x66 & ~x85 & ~x109 & ~x117 & ~x137 & ~x150 & ~x172 & ~x174 & ~x188 & ~x189 & ~x196 & ~x216 & ~x273 & ~x307 & ~x626 & ~x640 & ~x648 & ~x652 & ~x657 & ~x660 & ~x678 & ~x688 & ~x694 & ~x703 & ~x709 & ~x717 & ~x725 & ~x730 & ~x740 & ~x757;
assign c7388 =  x319 &  x320 &  x346 & ~x15 & ~x18 & ~x20 & ~x21 & ~x22 & ~x24 & ~x25 & ~x26 & ~x30 & ~x31 & ~x40 & ~x54 & ~x55 & ~x56 & ~x57 & ~x58 & ~x61 & ~x67 & ~x70 & ~x81 & ~x85 & ~x86 & ~x88 & ~x91 & ~x93 & ~x94 & ~x96 & ~x101 & ~x105 & ~x107 & ~x114 & ~x120 & ~x121 & ~x122 & ~x123 & ~x124 & ~x125 & ~x126 & ~x127 & ~x129 & ~x133 & ~x135 & ~x138 & ~x141 & ~x142 & ~x146 & ~x150 & ~x151 & ~x164 & ~x166 & ~x173 & ~x174 & ~x175 & ~x176 & ~x177 & ~x179 & ~x181 & ~x189 & ~x194 & ~x195 & ~x196 & ~x201 & ~x202 & ~x205 & ~x224 & ~x226 & ~x227 & ~x231 & ~x251 & ~x252 & ~x254 & ~x255 & ~x256 & ~x259 & ~x273 & ~x284 & ~x310 & ~x336 & ~x364 & ~x609 & ~x613 & ~x616 & ~x618 & ~x619 & ~x640 & ~x643 & ~x646 & ~x649 & ~x652 & ~x654 & ~x655 & ~x657 & ~x659 & ~x662 & ~x663 & ~x669 & ~x678 & ~x684 & ~x687 & ~x688 & ~x689 & ~x693 & ~x696 & ~x700 & ~x701 & ~x702 & ~x705 & ~x706 & ~x708 & ~x709 & ~x711 & ~x713 & ~x717 & ~x719 & ~x723 & ~x724 & ~x730 & ~x731 & ~x735 & ~x740 & ~x741 & ~x743 & ~x744 & ~x746 & ~x747 & ~x749 & ~x751 & ~x756 & ~x760 & ~x761 & ~x765 & ~x771 & ~x775 & ~x782;
assign c7390 = ~x14 & ~x21 & ~x22 & ~x34 & ~x45 & ~x46 & ~x66 & ~x67 & ~x106 & ~x112 & ~x124 & ~x125 & ~x126 & ~x127 & ~x137 & ~x142 & ~x150 & ~x151 & ~x193 & ~x202 & ~x205 & ~x227 & ~x254 & ~x259 & ~x281 & ~x283 & ~x288 & ~x308 & ~x311 & ~x312 & ~x315 & ~x426 & ~x481 & ~x482 & ~x588 & ~x647 & ~x679 & ~x683 & ~x690 & ~x694 & ~x702 & ~x706 & ~x725 & ~x732 & ~x736 & ~x740 & ~x741 & ~x745 & ~x757 & ~x764 & ~x767 & ~x771 & ~x782;
assign c7392 =  x270 & ~x5 & ~x13 & ~x36 & ~x39 & ~x41 & ~x73 & ~x79 & ~x86 & ~x92 & ~x104 & ~x112 & ~x142 & ~x146 & ~x149 & ~x152 & ~x167 & ~x180 & ~x195 & ~x197 & ~x229 & ~x230 & ~x246 & ~x257 & ~x263 & ~x274 & ~x281 & ~x309 & ~x364 & ~x597 & ~x600 & ~x601 & ~x602 & ~x646 & ~x710 & ~x717 & ~x732 & ~x739 & ~x743 & ~x747 & ~x749 & ~x756 & ~x781;
assign c7394 =  x359 &  x386 &  x387 &  x416 &  x430 &  x455 &  x468 & ~x1 & ~x4 & ~x9 & ~x15 & ~x21 & ~x24 & ~x41 & ~x46 & ~x50 & ~x53 & ~x54 & ~x58 & ~x69 & ~x72 & ~x78 & ~x83 & ~x98 & ~x107 & ~x116 & ~x118 & ~x143 & ~x152 & ~x168 & ~x172 & ~x173 & ~x208 & ~x225 & ~x233 & ~x258 & ~x280 & ~x281 & ~x286 & ~x288 & ~x308 & ~x309 & ~x312 & ~x315 & ~x335 & ~x337 & ~x338 & ~x339 & ~x340 & ~x341 & ~x364 & ~x367 & ~x368 & ~x370 & ~x394 & ~x395 & ~x420 & ~x588 & ~x615 & ~x638 & ~x643 & ~x645 & ~x647 & ~x650 & ~x657 & ~x660 & ~x661 & ~x662 & ~x667 & ~x676 & ~x705 & ~x708 & ~x709 & ~x710 & ~x712 & ~x721 & ~x724 & ~x725 & ~x732 & ~x738 & ~x743 & ~x749 & ~x757 & ~x758 & ~x763 & ~x765 & ~x768 & ~x775;
assign c7396 = ~x71 & ~x183 & ~x500 & ~x501 & ~x516 & ~x521 & ~x534 & ~x566 & ~x628 & ~x773;
assign c7398 =  x484 &  x485 &  x515 & ~x0 & ~x2 & ~x17 & ~x21 & ~x27 & ~x32 & ~x37 & ~x43 & ~x47 & ~x48 & ~x49 & ~x55 & ~x56 & ~x66 & ~x78 & ~x86 & ~x87 & ~x92 & ~x95 & ~x109 & ~x110 & ~x118 & ~x119 & ~x120 & ~x137 & ~x168 & ~x178 & ~x203 & ~x233 & ~x234 & ~x235 & ~x257 & ~x260 & ~x287 & ~x310 & ~x368 & ~x396 & ~x397 & ~x421 & ~x422 & ~x476 & ~x608 & ~x609 & ~x624 & ~x643 & ~x698 & ~x699 & ~x700 & ~x706 & ~x707 & ~x721 & ~x728 & ~x739 & ~x741 & ~x744 & ~x746 & ~x761 & ~x765 & ~x773 & ~x775 & ~x776 & ~x778 & ~x782;
assign c7400 =  x378 &  x445 &  x574 &  x577 & ~x17 & ~x23 & ~x26 & ~x28 & ~x40 & ~x44 & ~x46 & ~x49 & ~x55 & ~x63 & ~x70 & ~x71 & ~x76 & ~x82 & ~x95 & ~x96 & ~x101 & ~x102 & ~x106 & ~x117 & ~x120 & ~x121 & ~x122 & ~x123 & ~x138 & ~x142 & ~x150 & ~x152 & ~x158 & ~x171 & ~x174 & ~x191 & ~x194 & ~x198 & ~x201 & ~x206 & ~x221 & ~x222 & ~x223 & ~x226 & ~x258 & ~x282 & ~x588 & ~x618 & ~x643 & ~x645 & ~x647 & ~x648 & ~x649 & ~x651 & ~x663 & ~x664 & ~x665 & ~x671 & ~x672 & ~x678 & ~x688 & ~x694 & ~x701 & ~x704 & ~x711 & ~x712 & ~x732 & ~x739 & ~x742 & ~x745 & ~x751 & ~x764 & ~x772 & ~x777;
assign c7402 =  x214 & ~x0 & ~x10 & ~x18 & ~x21 & ~x23 & ~x48 & ~x58 & ~x64 & ~x71 & ~x82 & ~x90 & ~x124 & ~x125 & ~x169 & ~x173 & ~x196 & ~x199 & ~x203 & ~x206 & ~x209 & ~x210 & ~x228 & ~x234 & ~x253 & ~x257 & ~x266 & ~x285 & ~x309 & ~x367 & ~x450 & ~x643 & ~x675 & ~x676 & ~x679 & ~x681 & ~x746 & ~x751 & ~x752 & ~x757 & ~x770 & ~x771 & ~x774;
assign c7404 = ~x4 & ~x14 & ~x17 & ~x21 & ~x35 & ~x37 & ~x44 & ~x47 & ~x48 & ~x55 & ~x57 & ~x60 & ~x64 & ~x65 & ~x70 & ~x83 & ~x88 & ~x91 & ~x94 & ~x110 & ~x120 & ~x141 & ~x147 & ~x150 & ~x151 & ~x152 & ~x167 & ~x177 & ~x180 & ~x200 & ~x203 & ~x208 & ~x226 & ~x230 & ~x231 & ~x235 & ~x283 & ~x342 & ~x364 & ~x425 & ~x483 & ~x532 & ~x627 & ~x638 & ~x679 & ~x695 & ~x697 & ~x717 & ~x719 & ~x722 & ~x730 & ~x736 & ~x737 & ~x743 & ~x747 & ~x749 & ~x754 & ~x765 & ~x772 & ~x777 & ~x783;
assign c7406 =  x270 & ~x4 & ~x7 & ~x9 & ~x14 & ~x15 & ~x16 & ~x23 & ~x24 & ~x25 & ~x28 & ~x31 & ~x35 & ~x39 & ~x41 & ~x42 & ~x49 & ~x50 & ~x53 & ~x58 & ~x59 & ~x62 & ~x64 & ~x66 & ~x67 & ~x68 & ~x69 & ~x71 & ~x73 & ~x89 & ~x98 & ~x100 & ~x103 & ~x110 & ~x111 & ~x113 & ~x116 & ~x121 & ~x122 & ~x124 & ~x129 & ~x132 & ~x133 & ~x136 & ~x138 & ~x140 & ~x141 & ~x142 & ~x147 & ~x148 & ~x151 & ~x152 & ~x153 & ~x154 & ~x162 & ~x163 & ~x166 & ~x173 & ~x175 & ~x180 & ~x182 & ~x196 & ~x200 & ~x201 & ~x204 & ~x224 & ~x227 & ~x231 & ~x233 & ~x253 & ~x255 & ~x259 & ~x285 & ~x287 & ~x288 & ~x308 & ~x310 & ~x312 & ~x337 & ~x369 & ~x396 & ~x420 & ~x570 & ~x572 & ~x616 & ~x619 & ~x644 & ~x647 & ~x652 & ~x653 & ~x657 & ~x660 & ~x664 & ~x669 & ~x670 & ~x672 & ~x673 & ~x676 & ~x677 & ~x678 & ~x679 & ~x680 & ~x686 & ~x687 & ~x696 & ~x698 & ~x701 & ~x703 & ~x705 & ~x707 & ~x712 & ~x717 & ~x729 & ~x734 & ~x738 & ~x739 & ~x740 & ~x744 & ~x752 & ~x763 & ~x764 & ~x765 & ~x769 & ~x777 & ~x778 & ~x782 & ~x783;
assign c7408 =  x188 &  x270 &  x301 &  x418 &  x446 &  x470 &  x502 & ~x13 & ~x36 & ~x116 & ~x338 & ~x420 & ~x733 & ~x735;
assign c7410 =  x305 & ~x11 & ~x16 & ~x17 & ~x22 & ~x31 & ~x32 & ~x35 & ~x38 & ~x39 & ~x55 & ~x58 & ~x59 & ~x63 & ~x67 & ~x72 & ~x79 & ~x84 & ~x85 & ~x100 & ~x106 & ~x117 & ~x118 & ~x122 & ~x126 & ~x135 & ~x147 & ~x154 & ~x170 & ~x175 & ~x176 & ~x180 & ~x201 & ~x203 & ~x204 & ~x222 & ~x224 & ~x229 & ~x232 & ~x256 & ~x257 & ~x259 & ~x544 & ~x545 & ~x622 & ~x635 & ~x636 & ~x639 & ~x640 & ~x641 & ~x654 & ~x655 & ~x663 & ~x666 & ~x670 & ~x678 & ~x685 & ~x686 & ~x687 & ~x697 & ~x700 & ~x708 & ~x710 & ~x712 & ~x718 & ~x724 & ~x726 & ~x734 & ~x738 & ~x741 & ~x742 & ~x746 & ~x747 & ~x749 & ~x751 & ~x752 & ~x757 & ~x762 & ~x769 & ~x770 & ~x776 & ~x779 & ~x781;
assign c7412 =  x660 &  x661 &  x669;
assign c7414 =  x489 & ~x1 & ~x3 & ~x5 & ~x6 & ~x8 & ~x13 & ~x20 & ~x21 & ~x22 & ~x28 & ~x36 & ~x37 & ~x40 & ~x48 & ~x54 & ~x57 & ~x58 & ~x66 & ~x75 & ~x82 & ~x91 & ~x92 & ~x101 & ~x105 & ~x108 & ~x109 & ~x113 & ~x117 & ~x119 & ~x124 & ~x125 & ~x129 & ~x134 & ~x135 & ~x140 & ~x143 & ~x144 & ~x145 & ~x148 & ~x149 & ~x150 & ~x154 & ~x162 & ~x163 & ~x164 & ~x165 & ~x173 & ~x175 & ~x177 & ~x194 & ~x196 & ~x198 & ~x204 & ~x206 & ~x217 & ~x218 & ~x220 & ~x227 & ~x230 & ~x237 & ~x249 & ~x250 & ~x262 & ~x285 & ~x288 & ~x289 & ~x307 & ~x313 & ~x314 & ~x315 & ~x319 & ~x341 & ~x342 & ~x365 & ~x366 & ~x367 & ~x368 & ~x370 & ~x371 & ~x397 & ~x615 & ~x622 & ~x623 & ~x628 & ~x636 & ~x648 & ~x649 & ~x650 & ~x660 & ~x664 & ~x674 & ~x680 & ~x687 & ~x689 & ~x691 & ~x696 & ~x703 & ~x705 & ~x707 & ~x708 & ~x712 & ~x716 & ~x720 & ~x730 & ~x731 & ~x733 & ~x741 & ~x744 & ~x746 & ~x754 & ~x755 & ~x765 & ~x770 & ~x774 & ~x781 & ~x782;
assign c7416 =  x187 & ~x19 & ~x79 & ~x138 & ~x177 & ~x200 & ~x394 & ~x664 & ~x776;
assign c7418 = ~x11 & ~x94 & ~x204 & ~x454 & ~x509 & ~x533 & ~x567 & ~x779;
assign c7420 = ~x3 & ~x6 & ~x8 & ~x9 & ~x10 & ~x12 & ~x16 & ~x18 & ~x22 & ~x36 & ~x47 & ~x49 & ~x52 & ~x53 & ~x56 & ~x59 & ~x60 & ~x63 & ~x65 & ~x66 & ~x67 & ~x71 & ~x73 & ~x74 & ~x75 & ~x83 & ~x84 & ~x86 & ~x88 & ~x92 & ~x93 & ~x95 & ~x100 & ~x103 & ~x104 & ~x107 & ~x111 & ~x112 & ~x114 & ~x115 & ~x119 & ~x122 & ~x123 & ~x124 & ~x125 & ~x131 & ~x136 & ~x137 & ~x145 & ~x149 & ~x150 & ~x152 & ~x153 & ~x155 & ~x156 & ~x163 & ~x169 & ~x171 & ~x174 & ~x180 & ~x181 & ~x197 & ~x198 & ~x202 & ~x203 & ~x224 & ~x225 & ~x226 & ~x230 & ~x232 & ~x233 & ~x252 & ~x253 & ~x255 & ~x257 & ~x258 & ~x260 & ~x261 & ~x262 & ~x284 & ~x288 & ~x289 & ~x290 & ~x291 & ~x308 & ~x309 & ~x339 & ~x344 & ~x364 & ~x371 & ~x392 & ~x396 & ~x397 & ~x398 & ~x422 & ~x537 & ~x588 & ~x618 & ~x643 & ~x645 & ~x652 & ~x655 & ~x660 & ~x662 & ~x664 & ~x675 & ~x679 & ~x681 & ~x682 & ~x685 & ~x690 & ~x693 & ~x694 & ~x695 & ~x697 & ~x699 & ~x700 & ~x704 & ~x705 & ~x706 & ~x708 & ~x710 & ~x711 & ~x714 & ~x718 & ~x719 & ~x720 & ~x728 & ~x729 & ~x731 & ~x735 & ~x737 & ~x738 & ~x741 & ~x742 & ~x745 & ~x751 & ~x753 & ~x759 & ~x760 & ~x762 & ~x767 & ~x768 & ~x769 & ~x776 & ~x777 & ~x782;
assign c7422 =  x321 &  x346 &  x378 &  x379 &  x429 &  x488 &  x489 &  x493 & ~x12 & ~x19 & ~x21 & ~x25 & ~x30 & ~x34 & ~x40 & ~x43 & ~x48 & ~x69 & ~x74 & ~x90 & ~x98 & ~x100 & ~x103 & ~x111 & ~x116 & ~x129 & ~x131 & ~x132 & ~x145 & ~x148 & ~x150 & ~x162 & ~x165 & ~x174 & ~x199 & ~x203 & ~x229 & ~x252 & ~x257 & ~x258 & ~x308 & ~x336 & ~x649 & ~x655 & ~x657 & ~x659 & ~x664 & ~x669 & ~x676 & ~x686 & ~x687 & ~x688 & ~x695 & ~x696 & ~x698 & ~x702 & ~x705 & ~x713 & ~x720 & ~x747 & ~x749 & ~x751 & ~x755 & ~x760 & ~x762 & ~x768 & ~x774;
assign c7424 =  x554 &  x633 & ~x27 & ~x126 & ~x138 & ~x319 & ~x365 & ~x700 & ~x771;
assign c7426 =  x362 &  x419 & ~x9 & ~x17 & ~x20 & ~x51 & ~x85 & ~x87 & ~x198 & ~x225 & ~x254 & ~x279 & ~x286 & ~x308 & ~x587 & ~x759;
assign c7428 =  x158 &  x446 & ~x35 & ~x45 & ~x228 & ~x232 & ~x339 & ~x694;
assign c7430 =  x361 &  x463 & ~x7 & ~x8 & ~x9 & ~x10 & ~x12 & ~x18 & ~x19 & ~x28 & ~x30 & ~x31 & ~x34 & ~x37 & ~x38 & ~x40 & ~x41 & ~x42 & ~x48 & ~x49 & ~x50 & ~x51 & ~x54 & ~x55 & ~x58 & ~x64 & ~x65 & ~x66 & ~x72 & ~x76 & ~x77 & ~x80 & ~x81 & ~x82 & ~x83 & ~x84 & ~x88 & ~x90 & ~x91 & ~x93 & ~x94 & ~x95 & ~x99 & ~x100 & ~x106 & ~x107 & ~x108 & ~x111 & ~x118 & ~x120 & ~x121 & ~x123 & ~x135 & ~x145 & ~x148 & ~x152 & ~x167 & ~x172 & ~x174 & ~x176 & ~x178 & ~x200 & ~x201 & ~x205 & ~x206 & ~x207 & ~x208 & ~x227 & ~x228 & ~x229 & ~x230 & ~x231 & ~x234 & ~x252 & ~x256 & ~x257 & ~x258 & ~x259 & ~x260 & ~x261 & ~x279 & ~x287 & ~x288 & ~x308 & ~x309 & ~x312 & ~x314 & ~x316 & ~x337 & ~x340 & ~x342 & ~x531 & ~x556 & ~x557 & ~x588 & ~x610 & ~x635 & ~x637 & ~x638 & ~x639 & ~x640 & ~x642 & ~x650 & ~x662 & ~x666 & ~x668 & ~x670 & ~x675 & ~x677 & ~x682 & ~x687 & ~x688 & ~x690 & ~x693 & ~x695 & ~x698 & ~x699 & ~x702 & ~x703 & ~x705 & ~x708 & ~x710 & ~x711 & ~x717 & ~x719 & ~x724 & ~x727 & ~x737 & ~x743 & ~x746 & ~x749 & ~x750 & ~x751 & ~x754 & ~x758 & ~x760 & ~x761 & ~x763 & ~x765 & ~x770 & ~x771 & ~x781 & ~x782;
assign c7432 =  x355 & ~x4 & ~x5 & ~x18 & ~x19 & ~x27 & ~x33 & ~x39 & ~x55 & ~x59 & ~x61 & ~x74 & ~x99 & ~x100 & ~x106 & ~x113 & ~x143 & ~x145 & ~x149 & ~x152 & ~x169 & ~x173 & ~x177 & ~x198 & ~x200 & ~x208 & ~x226 & ~x231 & ~x234 & ~x281 & ~x283 & ~x285 & ~x289 & ~x313 & ~x342 & ~x497 & ~x612 & ~x613 & ~x638 & ~x646 & ~x665 & ~x666 & ~x702 & ~x717 & ~x719 & ~x722 & ~x737 & ~x761 & ~x764 & ~x765 & ~x772;
assign c7434 =  x269 & ~x39 & ~x81 & ~x92 & ~x95 & ~x122 & ~x137 & ~x138 & ~x147 & ~x158 & ~x161 & ~x163 & ~x170 & ~x171 & ~x174 & ~x190 & ~x191 & ~x257 & ~x272 & ~x273 & ~x274 & ~x286 & ~x300 & ~x301 & ~x313 & ~x314 & ~x604 & ~x605 & ~x610 & ~x666 & ~x701 & ~x707 & ~x709 & ~x766 & ~x774;
assign c7436 =  x385 &  x410 &  x460 & ~x5 & ~x13 & ~x16 & ~x32 & ~x52 & ~x58 & ~x72 & ~x99 & ~x122 & ~x145 & ~x149 & ~x165 & ~x173 & ~x197 & ~x204 & ~x223 & ~x227 & ~x281 & ~x289 & ~x316 & ~x340 & ~x366 & ~x538 & ~x681 & ~x699 & ~x702 & ~x732 & ~x767;
assign c7438 =  x390 & ~x42 & ~x44 & ~x72 & ~x102 & ~x106 & ~x118 & ~x122 & ~x165 & ~x188 & ~x193 & ~x300 & ~x309 & ~x339 & ~x533 & ~x566 & ~x584 & ~x591 & ~x619 & ~x629 & ~x656 & ~x658 & ~x680 & ~x684 & ~x696 & ~x703 & ~x736;
assign c7440 =  x704;
assign c7442 = ~x7 & ~x37 & ~x39 & ~x40 & ~x45 & ~x73 & ~x74 & ~x76 & ~x77 & ~x80 & ~x83 & ~x93 & ~x95 & ~x106 & ~x116 & ~x128 & ~x131 & ~x133 & ~x134 & ~x153 & ~x154 & ~x159 & ~x162 & ~x170 & ~x173 & ~x176 & ~x181 & ~x189 & ~x195 & ~x203 & ~x218 & ~x222 & ~x228 & ~x229 & ~x231 & ~x256 & ~x309 & ~x441 & ~x536 & ~x589 & ~x590 & ~x594 & ~x629 & ~x631 & ~x643 & ~x645 & ~x653 & ~x657 & ~x658 & ~x660 & ~x662 & ~x670 & ~x673 & ~x680 & ~x684 & ~x685 & ~x687 & ~x691 & ~x696 & ~x710 & ~x711 & ~x717 & ~x730 & ~x731 & ~x733 & ~x736 & ~x737 & ~x738 & ~x739 & ~x741 & ~x745 & ~x752 & ~x755 & ~x767 & ~x769 & ~x770 & ~x771 & ~x773 & ~x774 & ~x776 & ~x780 & ~x782;
assign c7444 = ~x0 & ~x2 & ~x7 & ~x21 & ~x29 & ~x31 & ~x35 & ~x40 & ~x46 & ~x52 & ~x53 & ~x57 & ~x67 & ~x71 & ~x72 & ~x73 & ~x79 & ~x86 & ~x92 & ~x97 & ~x99 & ~x103 & ~x104 & ~x107 & ~x118 & ~x119 & ~x121 & ~x130 & ~x131 & ~x133 & ~x140 & ~x148 & ~x157 & ~x161 & ~x167 & ~x168 & ~x171 & ~x177 & ~x180 & ~x182 & ~x190 & ~x204 & ~x207 & ~x252 & ~x254 & ~x256 & ~x259 & ~x313 & ~x316 & ~x338 & ~x363 & ~x365 & ~x370 & ~x392 & ~x393 & ~x396 & ~x399 & ~x419 & ~x503 & ~x581 & ~x588 & ~x617 & ~x647 & ~x649 & ~x656 & ~x665 & ~x668 & ~x678 & ~x680 & ~x693 & ~x694 & ~x696 & ~x701 & ~x704 & ~x709 & ~x719 & ~x722 & ~x732 & ~x739 & ~x746 & ~x747 & ~x748 & ~x758 & ~x760 & ~x771 & ~x775 & ~x776 & ~x778 & ~x783;
assign c7446 =  x463 & ~x68 & ~x76 & ~x82 & ~x100 & ~x181 & ~x350 & ~x426 & ~x691 & ~x693 & ~x694 & ~x740 & ~x750 & ~x778;
assign c7448 =  x385 &  x446 & ~x1 & ~x3 & ~x5 & ~x10 & ~x12 & ~x13 & ~x14 & ~x15 & ~x17 & ~x18 & ~x19 & ~x20 & ~x24 & ~x26 & ~x31 & ~x33 & ~x37 & ~x39 & ~x49 & ~x53 & ~x67 & ~x69 & ~x70 & ~x77 & ~x83 & ~x89 & ~x93 & ~x95 & ~x98 & ~x100 & ~x102 & ~x105 & ~x106 & ~x107 & ~x110 & ~x112 & ~x116 & ~x118 & ~x120 & ~x122 & ~x126 & ~x127 & ~x131 & ~x132 & ~x136 & ~x139 & ~x140 & ~x141 & ~x143 & ~x144 & ~x146 & ~x147 & ~x148 & ~x152 & ~x153 & ~x162 & ~x164 & ~x165 & ~x180 & ~x181 & ~x192 & ~x197 & ~x200 & ~x201 & ~x203 & ~x204 & ~x206 & ~x210 & ~x221 & ~x222 & ~x224 & ~x229 & ~x230 & ~x231 & ~x236 & ~x239 & ~x251 & ~x257 & ~x260 & ~x262 & ~x263 & ~x265 & ~x282 & ~x287 & ~x290 & ~x308 & ~x309 & ~x310 & ~x311 & ~x312 & ~x314 & ~x336 & ~x338 & ~x340 & ~x394 & ~x589 & ~x644 & ~x660 & ~x662 & ~x664 & ~x668 & ~x678 & ~x683 & ~x688 & ~x691 & ~x694 & ~x699 & ~x702 & ~x703 & ~x709 & ~x711 & ~x712 & ~x713 & ~x714 & ~x716 & ~x720 & ~x721 & ~x722 & ~x724 & ~x726 & ~x733 & ~x734 & ~x735 & ~x736 & ~x737 & ~x740 & ~x742 & ~x747 & ~x748 & ~x751 & ~x755 & ~x756 & ~x757 & ~x762 & ~x769 & ~x770 & ~x772 & ~x773 & ~x778 & ~x779 & ~x780 & ~x781 & ~x783;
assign c7450 =  x506 & ~x0 & ~x1 & ~x4 & ~x9 & ~x16 & ~x18 & ~x20 & ~x21 & ~x27 & ~x34 & ~x37 & ~x39 & ~x41 & ~x48 & ~x50 & ~x60 & ~x62 & ~x63 & ~x64 & ~x65 & ~x66 & ~x67 & ~x68 & ~x72 & ~x80 & ~x84 & ~x87 & ~x93 & ~x96 & ~x102 & ~x104 & ~x106 & ~x107 & ~x108 & ~x109 & ~x113 & ~x115 & ~x121 & ~x125 & ~x128 & ~x132 & ~x146 & ~x147 & ~x149 & ~x152 & ~x158 & ~x163 & ~x167 & ~x176 & ~x179 & ~x181 & ~x192 & ~x193 & ~x200 & ~x201 & ~x203 & ~x207 & ~x208 & ~x210 & ~x220 & ~x225 & ~x228 & ~x231 & ~x245 & ~x246 & ~x251 & ~x253 & ~x259 & ~x272 & ~x273 & ~x282 & ~x300 & ~x301 & ~x308 & ~x309 & ~x364 & ~x365 & ~x618 & ~x620 & ~x644 & ~x649 & ~x651 & ~x656 & ~x658 & ~x663 & ~x667 & ~x669 & ~x677 & ~x686 & ~x688 & ~x689 & ~x690 & ~x699 & ~x700 & ~x701 & ~x702 & ~x706 & ~x711 & ~x720 & ~x721 & ~x722 & ~x733 & ~x738 & ~x743 & ~x747 & ~x748 & ~x752 & ~x758 & ~x771 & ~x772 & ~x775 & ~x777 & ~x781;
assign c7452 =  x405 &  x429 &  x430 &  x488 &  x492 &  x532 & ~x4 & ~x27 & ~x46 & ~x60 & ~x67 & ~x75 & ~x87 & ~x93 & ~x98 & ~x103 & ~x104 & ~x115 & ~x119 & ~x129 & ~x151 & ~x153 & ~x160 & ~x173 & ~x175 & ~x203 & ~x204 & ~x223 & ~x307 & ~x312 & ~x392 & ~x475 & ~x660 & ~x667 & ~x693 & ~x703 & ~x711 & ~x722 & ~x723 & ~x732 & ~x741;
assign c7454 =  x605 & ~x40 & ~x81 & ~x120 & ~x169 & ~x196 & ~x203 & ~x234 & ~x235 & ~x255 & ~x262 & ~x337 & ~x637 & ~x641 & ~x689 & ~x696 & ~x713 & ~x727 & ~x752;
assign c7456 = ~x3 & ~x14 & ~x24 & ~x31 & ~x41 & ~x88 & ~x94 & ~x101 & ~x121 & ~x132 & ~x134 & ~x138 & ~x144 & ~x160 & ~x166 & ~x169 & ~x194 & ~x201 & ~x204 & ~x220 & ~x259 & ~x282 & ~x284 & ~x288 & ~x337 & ~x369 & ~x397 & ~x503 & ~x547 & ~x635 & ~x656 & ~x658 & ~x659 & ~x665 & ~x679 & ~x683 & ~x686 & ~x694 & ~x699 & ~x701 & ~x703 & ~x705 & ~x717 & ~x723 & ~x727 & ~x736 & ~x748 & ~x754 & ~x756 & ~x761 & ~x766 & ~x771 & ~x780;
assign c7458 =  x412 &  x578 & ~x5 & ~x16 & ~x25 & ~x28 & ~x32 & ~x38 & ~x44 & ~x45 & ~x49 & ~x52 & ~x55 & ~x58 & ~x73 & ~x88 & ~x90 & ~x92 & ~x99 & ~x100 & ~x102 & ~x106 & ~x111 & ~x124 & ~x141 & ~x147 & ~x151 & ~x171 & ~x172 & ~x173 & ~x174 & ~x198 & ~x206 & ~x238 & ~x254 & ~x255 & ~x258 & ~x264 & ~x290 & ~x310 & ~x311 & ~x313 & ~x366 & ~x392 & ~x607 & ~x609 & ~x610 & ~x633 & ~x635 & ~x676 & ~x686 & ~x695 & ~x703 & ~x707 & ~x712 & ~x721 & ~x723 & ~x726 & ~x734 & ~x737 & ~x742 & ~x757 & ~x758 & ~x768 & ~x770 & ~x779 & ~x780;
assign c7460 = ~x41 & ~x71 & ~x91 & ~x99 & ~x103 & ~x165 & ~x176 & ~x193 & ~x198 & ~x228 & ~x229 & ~x230 & ~x246 & ~x301 & ~x439 & ~x662 & ~x756;
assign c7462 =  x297 &  x351 &  x352 &  x377 &  x380 &  x382 &  x403 &  x404 &  x429 & ~x1 & ~x2 & ~x4 & ~x5 & ~x6 & ~x7 & ~x8 & ~x9 & ~x11 & ~x13 & ~x15 & ~x16 & ~x18 & ~x19 & ~x21 & ~x22 & ~x23 & ~x24 & ~x25 & ~x26 & ~x27 & ~x28 & ~x29 & ~x30 & ~x31 & ~x32 & ~x33 & ~x34 & ~x35 & ~x37 & ~x38 & ~x39 & ~x40 & ~x41 & ~x42 & ~x43 & ~x44 & ~x45 & ~x46 & ~x48 & ~x49 & ~x50 & ~x51 & ~x52 & ~x55 & ~x56 & ~x57 & ~x58 & ~x59 & ~x61 & ~x63 & ~x64 & ~x65 & ~x66 & ~x67 & ~x68 & ~x69 & ~x70 & ~x71 & ~x72 & ~x73 & ~x74 & ~x75 & ~x76 & ~x77 & ~x78 & ~x79 & ~x80 & ~x81 & ~x82 & ~x83 & ~x84 & ~x85 & ~x86 & ~x87 & ~x88 & ~x89 & ~x90 & ~x91 & ~x92 & ~x94 & ~x95 & ~x96 & ~x98 & ~x99 & ~x101 & ~x102 & ~x103 & ~x104 & ~x105 & ~x106 & ~x107 & ~x109 & ~x110 & ~x111 & ~x112 & ~x113 & ~x114 & ~x116 & ~x117 & ~x118 & ~x119 & ~x125 & ~x126 & ~x127 & ~x129 & ~x132 & ~x133 & ~x134 & ~x135 & ~x136 & ~x137 & ~x138 & ~x141 & ~x142 & ~x143 & ~x144 & ~x145 & ~x146 & ~x147 & ~x148 & ~x149 & ~x150 & ~x151 & ~x152 & ~x153 & ~x154 & ~x155 & ~x158 & ~x159 & ~x160 & ~x161 & ~x162 & ~x164 & ~x165 & ~x166 & ~x167 & ~x168 & ~x170 & ~x171 & ~x172 & ~x173 & ~x174 & ~x175 & ~x176 & ~x177 & ~x178 & ~x179 & ~x180 & ~x189 & ~x194 & ~x196 & ~x197 & ~x199 & ~x201 & ~x202 & ~x203 & ~x204 & ~x205 & ~x206 & ~x207 & ~x208 & ~x223 & ~x224 & ~x226 & ~x227 & ~x228 & ~x229 & ~x232 & ~x233 & ~x234 & ~x235 & ~x251 & ~x252 & ~x253 & ~x255 & ~x256 & ~x257 & ~x258 & ~x260 & ~x261 & ~x262 & ~x279 & ~x280 & ~x281 & ~x282 & ~x283 & ~x284 & ~x286 & ~x287 & ~x288 & ~x307 & ~x308 & ~x310 & ~x312 & ~x313 & ~x314 & ~x315 & ~x316 & ~x335 & ~x336 & ~x338 & ~x342 & ~x343 & ~x364 & ~x392 & ~x560 & ~x588 & ~x589 & ~x615 & ~x616 & ~x617 & ~x618 & ~x619 & ~x620 & ~x621 & ~x622 & ~x624 & ~x627 & ~x629 & ~x630 & ~x632 & ~x633 & ~x634 & ~x635 & ~x636 & ~x637 & ~x638 & ~x639 & ~x640 & ~x641 & ~x642 & ~x643 & ~x644 & ~x646 & ~x647 & ~x648 & ~x649 & ~x650 & ~x651 & ~x653 & ~x654 & ~x655 & ~x656 & ~x657 & ~x658 & ~x659 & ~x662 & ~x663 & ~x664 & ~x665 & ~x666 & ~x667 & ~x668 & ~x669 & ~x670 & ~x671 & ~x672 & ~x673 & ~x675 & ~x676 & ~x677 & ~x680 & ~x681 & ~x682 & ~x683 & ~x684 & ~x685 & ~x687 & ~x688 & ~x689 & ~x690 & ~x692 & ~x693 & ~x694 & ~x695 & ~x696 & ~x697 & ~x698 & ~x699 & ~x701 & ~x702 & ~x703 & ~x704 & ~x705 & ~x706 & ~x707 & ~x708 & ~x709 & ~x711 & ~x712 & ~x713 & ~x715 & ~x716 & ~x718 & ~x719 & ~x720 & ~x721 & ~x723 & ~x724 & ~x726 & ~x727 & ~x728 & ~x729 & ~x730 & ~x731 & ~x732 & ~x733 & ~x734 & ~x735 & ~x737 & ~x738 & ~x740 & ~x741 & ~x742 & ~x743 & ~x744 & ~x745 & ~x746 & ~x747 & ~x748 & ~x749 & ~x750 & ~x751 & ~x755 & ~x756 & ~x757 & ~x758 & ~x759 & ~x761 & ~x763 & ~x764 & ~x765 & ~x766 & ~x767 & ~x768 & ~x769 & ~x771 & ~x772 & ~x773 & ~x774 & ~x775 & ~x776 & ~x777 & ~x778 & ~x779 & ~x780 & ~x781 & ~x782 & ~x783;
assign c7464 = ~x4 & ~x10 & ~x14 & ~x18 & ~x22 & ~x28 & ~x30 & ~x34 & ~x42 & ~x46 & ~x47 & ~x49 & ~x53 & ~x54 & ~x58 & ~x67 & ~x69 & ~x73 & ~x74 & ~x79 & ~x82 & ~x83 & ~x84 & ~x89 & ~x92 & ~x94 & ~x96 & ~x97 & ~x100 & ~x101 & ~x104 & ~x109 & ~x110 & ~x113 & ~x114 & ~x115 & ~x116 & ~x119 & ~x122 & ~x127 & ~x139 & ~x144 & ~x145 & ~x154 & ~x158 & ~x161 & ~x162 & ~x164 & ~x168 & ~x170 & ~x180 & ~x181 & ~x182 & ~x188 & ~x190 & ~x191 & ~x196 & ~x200 & ~x203 & ~x209 & ~x225 & ~x226 & ~x227 & ~x228 & ~x230 & ~x232 & ~x236 & ~x238 & ~x256 & ~x258 & ~x261 & ~x280 & ~x291 & ~x313 & ~x315 & ~x335 & ~x337 & ~x344 & ~x364 & ~x368 & ~x369 & ~x370 & ~x397 & ~x535 & ~x536 & ~x561 & ~x589 & ~x615 & ~x617 & ~x620 & ~x621 & ~x622 & ~x624 & ~x632 & ~x634 & ~x638 & ~x643 & ~x648 & ~x653 & ~x654 & ~x655 & ~x660 & ~x663 & ~x666 & ~x668 & ~x669 & ~x672 & ~x675 & ~x677 & ~x678 & ~x680 & ~x689 & ~x693 & ~x700 & ~x701 & ~x704 & ~x705 & ~x707 & ~x714 & ~x722 & ~x726 & ~x728 & ~x729 & ~x734 & ~x738 & ~x743 & ~x744 & ~x745 & ~x747 & ~x748 & ~x750 & ~x754 & ~x756 & ~x761 & ~x762 & ~x763 & ~x766 & ~x767 & ~x769 & ~x775 & ~x781;
assign c7466 =  x665 & ~x346;
assign c7468 =  x326 &  x417 &  x440 &  x472 & ~x0 & ~x1 & ~x7 & ~x8 & ~x14 & ~x18 & ~x20 & ~x25 & ~x31 & ~x33 & ~x41 & ~x42 & ~x51 & ~x55 & ~x58 & ~x63 & ~x64 & ~x72 & ~x73 & ~x75 & ~x78 & ~x82 & ~x87 & ~x101 & ~x107 & ~x109 & ~x123 & ~x126 & ~x133 & ~x135 & ~x139 & ~x143 & ~x146 & ~x151 & ~x155 & ~x160 & ~x166 & ~x167 & ~x174 & ~x176 & ~x177 & ~x189 & ~x191 & ~x192 & ~x194 & ~x195 & ~x201 & ~x203 & ~x204 & ~x220 & ~x224 & ~x235 & ~x236 & ~x256 & ~x264 & ~x267 & ~x284 & ~x287 & ~x290 & ~x365 & ~x366 & ~x368 & ~x395 & ~x421 & ~x645 & ~x663 & ~x664 & ~x671 & ~x672 & ~x675 & ~x683 & ~x696 & ~x700 & ~x708 & ~x718 & ~x726 & ~x735 & ~x740 & ~x754 & ~x755 & ~x764 & ~x778;
assign c7470 = ~x10 & ~x11 & ~x26 & ~x42 & ~x43 & ~x45 & ~x51 & ~x56 & ~x65 & ~x76 & ~x82 & ~x97 & ~x102 & ~x106 & ~x129 & ~x133 & ~x153 & ~x159 & ~x162 & ~x193 & ~x204 & ~x210 & ~x227 & ~x229 & ~x244 & ~x271 & ~x273 & ~x301 & ~x316 & ~x336 & ~x356 & ~x572 & ~x616 & ~x679 & ~x681 & ~x732 & ~x735 & ~x745 & ~x753 & ~x755 & ~x762 & ~x772 & ~x777;
assign c7472 =  x605 & ~x11 & ~x13 & ~x34 & ~x42 & ~x48 & ~x62 & ~x67 & ~x80 & ~x97 & ~x112 & ~x118 & ~x119 & ~x148 & ~x154 & ~x163 & ~x167 & ~x168 & ~x179 & ~x181 & ~x283 & ~x284 & ~x588 & ~x589 & ~x615 & ~x637 & ~x640 & ~x642 & ~x650 & ~x665 & ~x672 & ~x678 & ~x684 & ~x688 & ~x691 & ~x708 & ~x713 & ~x721 & ~x733 & ~x744 & ~x764 & ~x769 & ~x782;
assign c7474 =  x633 &  x634 &  x639 & ~x290 & ~x312;
assign c7476 =  x185 & ~x5 & ~x175 & ~x634 & ~x636 & ~x657 & ~x668 & ~x758;
assign c7478 = ~x7 & ~x20 & ~x21 & ~x63 & ~x71 & ~x81 & ~x85 & ~x109 & ~x145 & ~x150 & ~x170 & ~x197 & ~x254 & ~x283 & ~x313 & ~x316 & ~x342 & ~x449 & ~x481 & ~x483 & ~x532 & ~x638 & ~x695 & ~x696 & ~x712 & ~x717 & ~x718 & ~x729 & ~x735 & ~x753 & ~x755 & ~x765 & ~x772 & ~x773;
assign c7480 = ~x3 & ~x8 & ~x9 & ~x15 & ~x18 & ~x19 & ~x21 & ~x27 & ~x28 & ~x32 & ~x34 & ~x37 & ~x41 & ~x46 & ~x51 & ~x55 & ~x58 & ~x65 & ~x66 & ~x69 & ~x83 & ~x85 & ~x86 & ~x87 & ~x88 & ~x93 & ~x98 & ~x100 & ~x101 & ~x102 & ~x105 & ~x106 & ~x108 & ~x118 & ~x122 & ~x128 & ~x130 & ~x133 & ~x140 & ~x141 & ~x151 & ~x152 & ~x154 & ~x161 & ~x165 & ~x170 & ~x175 & ~x178 & ~x182 & ~x190 & ~x201 & ~x203 & ~x208 & ~x210 & ~x220 & ~x221 & ~x222 & ~x224 & ~x231 & ~x251 & ~x253 & ~x255 & ~x273 & ~x282 & ~x284 & ~x307 & ~x309 & ~x310 & ~x312 & ~x313 & ~x395 & ~x426 & ~x428 & ~x588 & ~x608 & ~x622 & ~x646 & ~x647 & ~x651 & ~x657 & ~x658 & ~x661 & ~x667 & ~x671 & ~x672 & ~x676 & ~x679 & ~x688 & ~x691 & ~x692 & ~x696 & ~x698 & ~x701 & ~x704 & ~x713 & ~x717 & ~x720 & ~x733 & ~x735 & ~x745 & ~x748 & ~x751 & ~x752 & ~x755 & ~x760 & ~x761 & ~x762 & ~x764 & ~x770 & ~x773 & ~x780;
assign c7482 =  x186 &  x415 & ~x3 & ~x8 & ~x9 & ~x15 & ~x40 & ~x50 & ~x63 & ~x84 & ~x101 & ~x116 & ~x143 & ~x163 & ~x167 & ~x197 & ~x223 & ~x227 & ~x255 & ~x284 & ~x311 & ~x312 & ~x649 & ~x669 & ~x710 & ~x712 & ~x728 & ~x739 & ~x749 & ~x750 & ~x752 & ~x770;
assign c7484 =  x350 &  x353 &  x382 &  x402 &  x462 & ~x0 & ~x11 & ~x25 & ~x28 & ~x34 & ~x38 & ~x42 & ~x51 & ~x57 & ~x65 & ~x79 & ~x83 & ~x85 & ~x88 & ~x111 & ~x117 & ~x131 & ~x133 & ~x142 & ~x149 & ~x164 & ~x169 & ~x175 & ~x176 & ~x182 & ~x188 & ~x193 & ~x199 & ~x206 & ~x210 & ~x211 & ~x224 & ~x237 & ~x255 & ~x310 & ~x342 & ~x343 & ~x367 & ~x368 & ~x394 & ~x617 & ~x649 & ~x652 & ~x655 & ~x657 & ~x663 & ~x665 & ~x674 & ~x684 & ~x693 & ~x695 & ~x698 & ~x707 & ~x711 & ~x714 & ~x724 & ~x735 & ~x739 & ~x744 & ~x763 & ~x765 & ~x773 & ~x776 & ~x778;
assign c7486 =  x75;
assign c7488 = ~x1 & ~x3 & ~x5 & ~x10 & ~x15 & ~x22 & ~x23 & ~x24 & ~x29 & ~x31 & ~x37 & ~x40 & ~x42 & ~x43 & ~x45 & ~x49 & ~x55 & ~x56 & ~x58 & ~x60 & ~x61 & ~x67 & ~x68 & ~x69 & ~x71 & ~x72 & ~x74 & ~x76 & ~x78 & ~x80 & ~x82 & ~x84 & ~x92 & ~x95 & ~x96 & ~x99 & ~x101 & ~x104 & ~x107 & ~x108 & ~x115 & ~x117 & ~x118 & ~x121 & ~x127 & ~x129 & ~x131 & ~x135 & ~x136 & ~x137 & ~x138 & ~x140 & ~x141 & ~x146 & ~x148 & ~x151 & ~x152 & ~x154 & ~x155 & ~x156 & ~x159 & ~x160 & ~x162 & ~x163 & ~x165 & ~x166 & ~x167 & ~x169 & ~x170 & ~x171 & ~x172 & ~x176 & ~x177 & ~x178 & ~x183 & ~x187 & ~x188 & ~x192 & ~x193 & ~x194 & ~x197 & ~x198 & ~x199 & ~x200 & ~x201 & ~x203 & ~x204 & ~x205 & ~x207 & ~x208 & ~x210 & ~x213 & ~x217 & ~x222 & ~x223 & ~x224 & ~x226 & ~x227 & ~x229 & ~x231 & ~x237 & ~x238 & ~x245 & ~x253 & ~x255 & ~x258 & ~x261 & ~x262 & ~x279 & ~x280 & ~x281 & ~x284 & ~x285 & ~x287 & ~x312 & ~x314 & ~x315 & ~x316 & ~x336 & ~x342 & ~x343 & ~x364 & ~x392 & ~x526 & ~x528 & ~x529 & ~x588 & ~x622 & ~x636 & ~x637 & ~x647 & ~x649 & ~x650 & ~x651 & ~x652 & ~x658 & ~x663 & ~x668 & ~x670 & ~x671 & ~x672 & ~x674 & ~x676 & ~x679 & ~x687 & ~x689 & ~x691 & ~x693 & ~x694 & ~x700 & ~x703 & ~x705 & ~x707 & ~x709 & ~x710 & ~x713 & ~x714 & ~x717 & ~x719 & ~x726 & ~x733 & ~x738 & ~x739 & ~x740 & ~x742 & ~x743 & ~x744 & ~x746 & ~x750 & ~x752 & ~x757 & ~x758 & ~x761 & ~x763 & ~x764 & ~x765 & ~x767 & ~x769 & ~x770 & ~x781;
assign c7490 = ~x15 & ~x24 & ~x28 & ~x45 & ~x46 & ~x52 & ~x59 & ~x62 & ~x71 & ~x73 & ~x77 & ~x84 & ~x104 & ~x133 & ~x146 & ~x160 & ~x173 & ~x182 & ~x195 & ~x203 & ~x206 & ~x209 & ~x210 & ~x229 & ~x230 & ~x253 & ~x257 & ~x259 & ~x261 & ~x285 & ~x288 & ~x289 & ~x309 & ~x312 & ~x392 & ~x424 & ~x453 & ~x454 & ~x455 & ~x597 & ~x702 & ~x727 & ~x733 & ~x738 & ~x746 & ~x753 & ~x763 & ~x770 & ~x772 & ~x782;
assign c7492 =  x474 &  x606 & ~x0 & ~x1 & ~x37 & ~x42 & ~x79 & ~x86 & ~x106 & ~x112 & ~x117 & ~x120 & ~x142 & ~x146 & ~x165 & ~x197 & ~x282 & ~x283 & ~x284 & ~x287 & ~x344 & ~x364 & ~x371 & ~x397 & ~x398 & ~x451 & ~x768 & ~x782;
assign c7494 =  x577 & ~x0 & ~x8 & ~x11 & ~x16 & ~x22 & ~x26 & ~x30 & ~x31 & ~x34 & ~x37 & ~x41 & ~x48 & ~x49 & ~x50 & ~x52 & ~x53 & ~x57 & ~x59 & ~x63 & ~x66 & ~x67 & ~x70 & ~x74 & ~x76 & ~x77 & ~x81 & ~x86 & ~x91 & ~x92 & ~x94 & ~x96 & ~x97 & ~x100 & ~x104 & ~x106 & ~x111 & ~x115 & ~x118 & ~x120 & ~x124 & ~x126 & ~x131 & ~x132 & ~x136 & ~x139 & ~x142 & ~x143 & ~x144 & ~x145 & ~x148 & ~x151 & ~x154 & ~x160 & ~x165 & ~x166 & ~x167 & ~x176 & ~x177 & ~x178 & ~x181 & ~x189 & ~x195 & ~x196 & ~x197 & ~x199 & ~x200 & ~x218 & ~x220 & ~x221 & ~x222 & ~x226 & ~x235 & ~x236 & ~x255 & ~x257 & ~x259 & ~x260 & ~x262 & ~x263 & ~x278 & ~x280 & ~x283 & ~x288 & ~x309 & ~x313 & ~x315 & ~x340 & ~x365 & ~x367 & ~x368 & ~x649 & ~x660 & ~x668 & ~x669 & ~x678 & ~x687 & ~x691 & ~x693 & ~x702 & ~x705 & ~x707 & ~x708 & ~x709 & ~x710 & ~x713 & ~x721 & ~x722 & ~x727 & ~x730 & ~x734 & ~x740 & ~x741 & ~x744 & ~x748 & ~x751 & ~x752 & ~x756 & ~x757 & ~x759 & ~x760 & ~x765 & ~x770 & ~x772 & ~x779 & ~x781;
assign c7496 =  x322 &  x347 &  x371 &  x423 & ~x33 & ~x73 & ~x75 & ~x78 & ~x91 & ~x94 & ~x168 & ~x177 & ~x179 & ~x228 & ~x258 & ~x259 & ~x313 & ~x602 & ~x614 & ~x615 & ~x624 & ~x649 & ~x657 & ~x676 & ~x689 & ~x692 & ~x693 & ~x708 & ~x723 & ~x772 & ~x782 & ~x783;
assign c7498 =  x269 &  x347 &  x349 &  x353 &  x373 & ~x3 & ~x9 & ~x10 & ~x11 & ~x12 & ~x15 & ~x16 & ~x18 & ~x24 & ~x25 & ~x30 & ~x33 & ~x37 & ~x42 & ~x45 & ~x53 & ~x54 & ~x65 & ~x66 & ~x69 & ~x70 & ~x72 & ~x75 & ~x80 & ~x82 & ~x86 & ~x87 & ~x105 & ~x109 & ~x111 & ~x113 & ~x114 & ~x115 & ~x117 & ~x118 & ~x120 & ~x122 & ~x136 & ~x137 & ~x141 & ~x142 & ~x144 & ~x145 & ~x146 & ~x149 & ~x150 & ~x151 & ~x154 & ~x160 & ~x162 & ~x169 & ~x170 & ~x176 & ~x177 & ~x178 & ~x180 & ~x200 & ~x202 & ~x204 & ~x208 & ~x223 & ~x227 & ~x233 & ~x234 & ~x235 & ~x258 & ~x259 & ~x260 & ~x279 & ~x280 & ~x286 & ~x309 & ~x310 & ~x312 & ~x336 & ~x588 & ~x589 & ~x615 & ~x616 & ~x617 & ~x626 & ~x641 & ~x655 & ~x657 & ~x663 & ~x666 & ~x675 & ~x677 & ~x678 & ~x679 & ~x682 & ~x683 & ~x688 & ~x689 & ~x690 & ~x693 & ~x696 & ~x697 & ~x700 & ~x702 & ~x706 & ~x710 & ~x713 & ~x717 & ~x722 & ~x723 & ~x728 & ~x741 & ~x753 & ~x757 & ~x762 & ~x764 & ~x765 & ~x766 & ~x774 & ~x776 & ~x778 & ~x781 & ~x782;
assign c71 =  x240 &  x295 &  x296 &  x299 &  x303 &  x304 &  x381 &  x415 &  x441 &  x490 &  x506 &  x516 &  x518 &  x522 &  x530 &  x534 &  x540 &  x543 &  x545 &  x547 &  x557 &  x564 &  x567 &  x570 &  x573 &  x599 & ~x26 & ~x35 & ~x43 & ~x60 & ~x67 & ~x101 & ~x105 & ~x110 & ~x120 & ~x123 & ~x134 & ~x153 & ~x173 & ~x225 & ~x235 & ~x256 & ~x259 & ~x309 & ~x343 & ~x371 & ~x662 & ~x688 & ~x689 & ~x706 & ~x771;
assign c73 =  x207;
assign c75 =  x357 & ~x270 & ~x417 & ~x418 & ~x421;
assign c77 =  x143;
assign c79 =  x439 &  x473 &  x563 & ~x63 & ~x80 & ~x124 & ~x401 & ~x632 & ~x710;
assign c711 =  x648 &  x651;
assign c713 =  x629 &  x667 & ~x689;
assign c715 =  x613 &  x669;
assign c717 =  x70;
assign c721 =  x261;
assign c723 =  x601 &  x611 &  x620 &  x628 &  x652 &  x653;
assign c725 =  x89 &  x144;
assign c727 =  x387 & ~x393 & ~x404 & ~x450 & ~x461;
assign c729 = ~x249 & ~x278 & ~x419 & ~x444;
assign c731 =  x573 &  x613 & ~x98 & ~x162 & ~x631 & ~x754 & ~x764;
assign c733 =  x437 & ~x333 & ~x334 & ~x387 & ~x390;
assign c735 =  x466 & ~x270 & ~x271 & ~x362 & ~x389;
assign c737 =  x44;
assign c739 =  x695;
assign c741 =  x641 & ~x661;
assign c743 =  x602 &  x626 & ~x634;
assign c745 =  x175;
assign c747 =  x18;
assign c749 = ~x436 & ~x463;
assign c751 =  x201;
assign c753 =  x194;
assign c755 =  x203;
assign c757 = ~x242 & ~x390 & ~x394 & ~x416 & ~x418 & ~x574 & ~x581;
assign c759 =  x301 &  x557 & ~x2 & ~x5 & ~x17 & ~x20 & ~x21 & ~x26 & ~x29 & ~x31 & ~x32 & ~x33 & ~x40 & ~x41 & ~x47 & ~x48 & ~x57 & ~x62 & ~x65 & ~x66 & ~x71 & ~x78 & ~x84 & ~x89 & ~x97 & ~x107 & ~x111 & ~x112 & ~x113 & ~x115 & ~x126 & ~x127 & ~x129 & ~x132 & ~x136 & ~x138 & ~x142 & ~x145 & ~x147 & ~x151 & ~x154 & ~x155 & ~x156 & ~x157 & ~x159 & ~x163 & ~x166 & ~x167 & ~x178 & ~x198 & ~x200 & ~x201 & ~x227 & ~x232 & ~x256 & ~x257 & ~x260 & ~x263 & ~x279 & ~x290 & ~x308 & ~x367 & ~x370 & ~x392 & ~x393 & ~x394 & ~x531 & ~x559 & ~x618 & ~x634 & ~x646 & ~x648 & ~x656 & ~x661 & ~x673 & ~x677 & ~x685 & ~x696 & ~x702 & ~x711 & ~x712 & ~x718 & ~x721 & ~x725 & ~x733 & ~x738 & ~x739 & ~x742 & ~x748 & ~x751 & ~x758 & ~x760 & ~x769 & ~x775 & ~x782;
assign c761 =  x207;
assign c763 =  x82;
assign c765 =  x511 & ~x378 & ~x407 & ~x420;
assign c767 =  x47;
assign c769 =  x191 &  x585;
assign c771 = ~x417 & ~x418 & ~x577 & ~x582 & ~x585;
assign c773 =  x72;
assign c775 = ~x4 & ~x25 & ~x29 & ~x130 & ~x131 & ~x231 & ~x280 & ~x376 & ~x393 & ~x394 & ~x421 & ~x433 & ~x448 & ~x729 & ~x734;
assign c777 =  x135;
assign c779 =  x337;
assign c781 =  x258 &  x308;
assign c783 =  x308;
assign c785 =  x93;
assign c787 =  x54;
assign c789 =  x168;
assign c791 =  x295 &  x296 &  x473 &  x534 &  x555 & ~x52 & ~x428 & ~x662 & ~x702 & ~x708;
assign c793 =  x314;
assign c795 = ~x416 & ~x417 & ~x418 & ~x565 & ~x584 & ~x704;
assign c797 =  x710;
assign c799 = ~x248 & ~x418 & ~x421 & ~x444 & ~x614;
assign c7101 =  x224;
assign c7103 =  x37;
assign c7105 =  x454 & ~x101 & ~x107 & ~x119 & ~x155 & ~x158 & ~x228 & ~x236 & ~x242 & ~x244 & ~x258 & ~x261 & ~x262 & ~x268 & ~x269 & ~x287 & ~x309 & ~x339 & ~x651 & ~x682 & ~x699 & ~x770 & ~x783;
assign c7107 =  x21;
assign c7109 =  x512 &  x526 & ~x242 & ~x634;
assign c7111 =  x595 &  x613 &  x614 &  x644;
assign c7113 =  x13;
assign c7115 =  x315;
assign c7117 =  x268 &  x300 &  x304 &  x489 &  x495 &  x508 &  x513 &  x538 &  x553 & ~x20 & ~x30 & ~x69 & ~x70 & ~x76 & ~x85 & ~x91 & ~x126 & ~x138 & ~x279 & ~x289 & ~x312 & ~x606 & ~x607 & ~x619 & ~x629 & ~x632 & ~x675 & ~x711 & ~x714 & ~x722 & ~x730;
assign c7119 =  x425 &  x453 & ~x241 & ~x306 & ~x311;
assign c7121 =  x473 &  x509 &  x556 &  x565 &  x569 &  x584 &  x613 & ~x423 & ~x477;
assign c7125 =  x56;
assign c7127 =  x439 & ~x333 & ~x353;
assign c7129 =  x202;
assign c7131 =  x246 &  x248 &  x298 &  x506 &  x534 &  x601 &  x611 & ~x476;
assign c7133 =  x227;
assign c7135 = ~x319 & ~x406 & ~x407 & ~x435 & ~x449 & ~x615 & ~x744;
assign c7137 = ~x351 & ~x577;
assign c7139 =  x221 &  x556 &  x557 &  x570 &  x612 & ~x74 & ~x101 & ~x729;
assign c7141 =  x481 &  x495 & ~x418 & ~x445;
assign c7143 =  x257;
assign c7145 =  x670;
assign c7147 =  x269 &  x295 &  x296 &  x298 &  x303 &  x305 &  x325 &  x327 &  x333 &  x351 &  x357 &  x359 &  x361 &  x408 &  x413 &  x433 &  x462 &  x467 &  x493 &  x508 &  x515 &  x553 &  x557 &  x582 & ~x5 & ~x12 & ~x49 & ~x68 & ~x70 & ~x82 & ~x87 & ~x93 & ~x102 & ~x103 & ~x108 & ~x109 & ~x120 & ~x123 & ~x140 & ~x147 & ~x171 & ~x179 & ~x206 & ~x225 & ~x233 & ~x255 & ~x307 & ~x314 & ~x315 & ~x363 & ~x366 & ~x371 & ~x374 & ~x391 & ~x393 & ~x659 & ~x680 & ~x687 & ~x708 & ~x725 & ~x751 & ~x764 & ~x772;
assign c7149 =  x219 &  x490 &  x574 &  x612 & ~x143 & ~x280 & ~x391 & ~x689;
assign c7151 =  x364;
assign c7153 =  x572 &  x573 &  x614 & ~x633 & ~x661;
assign c7155 =  x537 & ~x4 & ~x8 & ~x21 & ~x36 & ~x39 & ~x62 & ~x66 & ~x77 & ~x88 & ~x93 & ~x99 & ~x112 & ~x122 & ~x132 & ~x134 & ~x140 & ~x145 & ~x146 & ~x149 & ~x156 & ~x168 & ~x185 & ~x199 & ~x200 & ~x201 & ~x206 & ~x225 & ~x226 & ~x251 & ~x262 & ~x281 & ~x315 & ~x337 & ~x341 & ~x345 & ~x346 & ~x364 & ~x375 & ~x421 & ~x423 & ~x616 & ~x620 & ~x633 & ~x643 & ~x646 & ~x654 & ~x656 & ~x686 & ~x692 & ~x696 & ~x707 & ~x712 & ~x734 & ~x748 & ~x751 & ~x755 & ~x757 & ~x758 & ~x759 & ~x760 & ~x761 & ~x763 & ~x768 & ~x774;
assign c7157 =  x277 &  x470 &  x501 &  x534 & ~x58 & ~x187 & ~x401 & ~x424 & ~x426 & ~x634 & ~x688 & ~x743;
assign c7159 = ~x313 & ~x371 & ~x477;
assign c7161 =  x336;
assign c7163 =  x719;
assign c7165 =  x762;
assign c7167 =  x510 & ~x86 & ~x126 & ~x181 & ~x184 & ~x185 & ~x478 & ~x643 & ~x672;
assign c7169 =  x168;
assign c7171 =  x771;
assign c7173 =  x710;
assign c7177 =  x171;
assign c7179 =  x198 &  x756;
assign c7181 =  x225;
assign c7183 =  x218 &  x557 & ~x306;
assign c7185 =  x191 &  x613;
assign c7187 =  x296 &  x327 &  x329 &  x330 &  x382 &  x439 &  x466 &  x481 &  x497 &  x502 &  x510 &  x511 &  x514 &  x524 & ~x2 & ~x32 & ~x36 & ~x45 & ~x46 & ~x47 & ~x52 & ~x56 & ~x60 & ~x61 & ~x75 & ~x80 & ~x81 & ~x84 & ~x85 & ~x92 & ~x96 & ~x103 & ~x105 & ~x109 & ~x111 & ~x116 & ~x119 & ~x122 & ~x125 & ~x127 & ~x129 & ~x131 & ~x137 & ~x144 & ~x151 & ~x154 & ~x157 & ~x161 & ~x164 & ~x168 & ~x173 & ~x179 & ~x189 & ~x204 & ~x220 & ~x231 & ~x259 & ~x291 & ~x337 & ~x364 & ~x588 & ~x590 & ~x603 & ~x606 & ~x623 & ~x624 & ~x641 & ~x653 & ~x654 & ~x655 & ~x657 & ~x658 & ~x666 & ~x668 & ~x671 & ~x678 & ~x686 & ~x690 & ~x699 & ~x716 & ~x720 & ~x721 & ~x723 & ~x729 & ~x740 & ~x741 & ~x748 & ~x749 & ~x753 & ~x766 & ~x767 & ~x769 & ~x770 & ~x771 & ~x776 & ~x781;
assign c7189 =  x312;
assign c7191 = ~x334 & ~x389 & ~x395 & ~x549 & ~x583;
assign c7193 =  x537 &  x538 &  x552 &  x553 & ~x61 & ~x79 & ~x132 & ~x138 & ~x147 & ~x202 & ~x259 & ~x288 & ~x320 & ~x345 & ~x606 & ~x616 & ~x618 & ~x623 & ~x630 & ~x632 & ~x662 & ~x676 & ~x697 & ~x714 & ~x726;
assign c7195 =  x62;
assign c7197 =  x258;
assign c7199 =  x118;
assign c7201 =  x667;
assign c7203 =  x616;
assign c7205 =  x573 &  x609 &  x611 & ~x9 & ~x449 & ~x634 & ~x659 & ~x660 & ~x661 & ~x704;
assign c7207 =  x242 &  x247 &  x248 &  x267 &  x270 &  x276 &  x325 &  x414 &  x433 &  x462 &  x490 &  x515 &  x535 &  x583 & ~x57 & ~x76 & ~x88 & ~x120 & ~x251 & ~x310 & ~x317 & ~x344 & ~x660 & ~x702 & ~x721 & ~x739 & ~x745 & ~x759;
assign c7209 =  x585 &  x649;
assign c7211 =  x780;
assign c7213 =  x114;
assign c7215 = ~x4 & ~x8 & ~x22 & ~x25 & ~x28 & ~x45 & ~x50 & ~x53 & ~x59 & ~x63 & ~x85 & ~x91 & ~x99 & ~x102 & ~x104 & ~x122 & ~x124 & ~x142 & ~x143 & ~x156 & ~x158 & ~x160 & ~x172 & ~x179 & ~x185 & ~x198 & ~x232 & ~x255 & ~x258 & ~x259 & ~x262 & ~x282 & ~x284 & ~x287 & ~x289 & ~x290 & ~x308 & ~x318 & ~x394 & ~x395 & ~x422 & ~x450 & ~x451 & ~x476 & ~x477 & ~x478 & ~x560 & ~x644 & ~x645 & ~x646 & ~x660 & ~x661 & ~x671 & ~x673 & ~x675 & ~x676 & ~x702 & ~x717 & ~x722 & ~x728 & ~x738 & ~x741 & ~x746 & ~x770 & ~x777 & ~x782;
assign c7217 =  x697;
assign c7219 =  x757;
assign c7221 =  x212 &  x557 &  x570 &  x573 &  x597 &  x611 &  x640 &  x641 & ~x79 & ~x315 & ~x690 & ~x719 & ~x766 & ~x771;
assign c7223 =  x283 &  x761;
assign c7225 =  x19;
assign c7227 =  x41;
assign c7229 =  x193 &  x611;
assign c7233 =  x100;
assign c7235 =  x235;
assign c7237 = ~x0 & ~x1 & ~x2 & ~x3 & ~x6 & ~x9 & ~x10 & ~x12 & ~x14 & ~x16 & ~x17 & ~x18 & ~x19 & ~x21 & ~x24 & ~x25 & ~x27 & ~x29 & ~x31 & ~x32 & ~x33 & ~x36 & ~x37 & ~x40 & ~x41 & ~x42 & ~x43 & ~x44 & ~x46 & ~x47 & ~x50 & ~x53 & ~x55 & ~x58 & ~x59 & ~x60 & ~x64 & ~x65 & ~x66 & ~x68 & ~x72 & ~x74 & ~x75 & ~x80 & ~x81 & ~x82 & ~x83 & ~x87 & ~x89 & ~x90 & ~x92 & ~x93 & ~x94 & ~x95 & ~x99 & ~x100 & ~x101 & ~x102 & ~x103 & ~x106 & ~x107 & ~x109 & ~x110 & ~x111 & ~x114 & ~x115 & ~x117 & ~x118 & ~x120 & ~x122 & ~x124 & ~x130 & ~x131 & ~x132 & ~x134 & ~x135 & ~x136 & ~x137 & ~x138 & ~x140 & ~x141 & ~x142 & ~x143 & ~x144 & ~x146 & ~x147 & ~x150 & ~x151 & ~x152 & ~x153 & ~x154 & ~x155 & ~x157 & ~x159 & ~x161 & ~x162 & ~x165 & ~x166 & ~x167 & ~x168 & ~x173 & ~x174 & ~x175 & ~x178 & ~x180 & ~x181 & ~x184 & ~x185 & ~x187 & ~x190 & ~x192 & ~x193 & ~x194 & ~x195 & ~x198 & ~x204 & ~x206 & ~x212 & ~x213 & ~x214 & ~x216 & ~x217 & ~x222 & ~x223 & ~x224 & ~x225 & ~x226 & ~x228 & ~x229 & ~x230 & ~x231 & ~x234 & ~x241 & ~x250 & ~x252 & ~x255 & ~x258 & ~x259 & ~x263 & ~x280 & ~x285 & ~x286 & ~x287 & ~x288 & ~x308 & ~x310 & ~x336 & ~x339 & ~x340 & ~x363 & ~x364 & ~x365 & ~x366 & ~x367 & ~x392 & ~x393 & ~x394 & ~x395 & ~x550 & ~x559 & ~x560 & ~x561 & ~x562 & ~x564 & ~x565 & ~x577 & ~x578 & ~x579 & ~x582 & ~x583 & ~x584 & ~x589 & ~x592 & ~x594 & ~x595 & ~x596 & ~x597 & ~x599 & ~x601 & ~x603 & ~x605 & ~x606 & ~x607 & ~x608 & ~x610 & ~x611 & ~x612 & ~x614 & ~x615 & ~x616 & ~x623 & ~x625 & ~x626 & ~x630 & ~x634 & ~x636 & ~x637 & ~x638 & ~x639 & ~x640 & ~x642 & ~x644 & ~x647 & ~x648 & ~x649 & ~x651 & ~x652 & ~x654 & ~x656 & ~x657 & ~x658 & ~x660 & ~x663 & ~x664 & ~x666 & ~x667 & ~x668 & ~x670 & ~x672 & ~x674 & ~x678 & ~x680 & ~x681 & ~x682 & ~x684 & ~x685 & ~x686 & ~x687 & ~x688 & ~x692 & ~x693 & ~x694 & ~x696 & ~x702 & ~x703 & ~x707 & ~x708 & ~x709 & ~x711 & ~x712 & ~x713 & ~x715 & ~x717 & ~x718 & ~x719 & ~x720 & ~x721 & ~x723 & ~x725 & ~x726 & ~x730 & ~x732 & ~x734 & ~x736 & ~x739 & ~x743 & ~x746 & ~x749 & ~x750 & ~x753 & ~x756 & ~x758 & ~x760 & ~x761 & ~x762 & ~x766 & ~x767 & ~x768 & ~x769 & ~x770 & ~x771 & ~x775 & ~x776 & ~x778 & ~x779 & ~x780 & ~x781;
assign c7239 =  x257;
assign c7241 =  x439 &  x456 & ~x295 & ~x296;
assign c7243 = ~x386 & ~x388;
assign c7245 =  x276 &  x299 &  x302 &  x408 &  x557 &  x567 &  x568 &  x571 &  x572 &  x584 & ~x13 & ~x15 & ~x33 & ~x55 & ~x86 & ~x115 & ~x119 & ~x138 & ~x145 & ~x316 & ~x339 & ~x559 & ~x633 & ~x646 & ~x659 & ~x661 & ~x674 & ~x690 & ~x753 & ~x774 & ~x780;
assign c7247 =  x358 & ~x417 & ~x418;
assign c7249 =  x20;
assign c7251 = ~x349 & ~x393 & ~x578;
assign c7253 =  x329 &  x330 &  x332 &  x497 & ~x18 & ~x88 & ~x89 & ~x91 & ~x123 & ~x131 & ~x137 & ~x168 & ~x180 & ~x185 & ~x186 & ~x218 & ~x229 & ~x231 & ~x242 & ~x640 & ~x683 & ~x706 & ~x734 & ~x743 & ~x770;
assign c7255 =  x55;
assign c7257 =  x695;
assign c7259 =  x669;
assign c7261 =  x336;
assign c7263 =  x256;
assign c7265 =  x229;
assign c7267 =  x136;
assign c7269 =  x68;
assign c7271 =  x482 & ~x4 & ~x83 & ~x105 & ~x118 & ~x124 & ~x151 & ~x164 & ~x173 & ~x182 & ~x214 & ~x215 & ~x216 & ~x217 & ~x345 & ~x366 & ~x578 & ~x614 & ~x632 & ~x668 & ~x776;
assign c7273 = ~x444;
assign c7275 =  x178;
assign c7277 =  x547 &  x585 & ~x2 & ~x4 & ~x16 & ~x24 & ~x28 & ~x35 & ~x36 & ~x44 & ~x46 & ~x47 & ~x56 & ~x60 & ~x63 & ~x64 & ~x81 & ~x84 & ~x85 & ~x89 & ~x96 & ~x97 & ~x99 & ~x107 & ~x115 & ~x119 & ~x137 & ~x142 & ~x169 & ~x173 & ~x176 & ~x179 & ~x201 & ~x208 & ~x228 & ~x230 & ~x252 & ~x254 & ~x284 & ~x308 & ~x316 & ~x338 & ~x341 & ~x346 & ~x398 & ~x399 & ~x420 & ~x589 & ~x606 & ~x619 & ~x620 & ~x632 & ~x634 & ~x635 & ~x647 & ~x662 & ~x676 & ~x677 & ~x686 & ~x692 & ~x698 & ~x708 & ~x715 & ~x719 & ~x730 & ~x738 & ~x741 & ~x743 & ~x748 & ~x749 & ~x763 & ~x766 & ~x771 & ~x774 & ~x775 & ~x779 & ~x781 & ~x783;
assign c7279 =  x244 & ~x418;
assign c7281 =  x276 &  x297 &  x303 &  x305 &  x328 &  x329 &  x354 &  x360 &  x381 &  x417 &  x418 &  x436 &  x438 &  x461 &  x464 &  x473 &  x485 &  x489 &  x491 &  x507 &  x509 &  x524 &  x540 &  x541 &  x553 &  x567 &  x581 &  x582 & ~x0 & ~x3 & ~x7 & ~x13 & ~x16 & ~x20 & ~x42 & ~x51 & ~x60 & ~x62 & ~x69 & ~x77 & ~x90 & ~x91 & ~x115 & ~x118 & ~x137 & ~x139 & ~x142 & ~x145 & ~x147 & ~x148 & ~x195 & ~x207 & ~x225 & ~x229 & ~x259 & ~x261 & ~x281 & ~x287 & ~x288 & ~x289 & ~x339 & ~x346 & ~x363 & ~x372 & ~x391 & ~x392 & ~x399 & ~x658 & ~x660 & ~x661 & ~x681 & ~x687 & ~x690 & ~x701 & ~x706 & ~x708 & ~x721 & ~x727 & ~x730 & ~x731 & ~x733 & ~x736 & ~x742 & ~x746 & ~x757 & ~x768 & ~x778 & ~x780;
assign c7283 =  x332 &  x356 &  x358 &  x412 & ~x2 & ~x5 & ~x7 & ~x10 & ~x13 & ~x14 & ~x23 & ~x34 & ~x35 & ~x38 & ~x61 & ~x69 & ~x80 & ~x87 & ~x88 & ~x90 & ~x99 & ~x126 & ~x133 & ~x135 & ~x137 & ~x152 & ~x155 & ~x157 & ~x165 & ~x167 & ~x170 & ~x172 & ~x181 & ~x184 & ~x200 & ~x212 & ~x218 & ~x219 & ~x259 & ~x282 & ~x307 & ~x309 & ~x316 & ~x319 & ~x419 & ~x607 & ~x617 & ~x625 & ~x626 & ~x636 & ~x640 & ~x646 & ~x652 & ~x671 & ~x678 & ~x687 & ~x692 & ~x697 & ~x723 & ~x727 & ~x728 & ~x736 & ~x737 & ~x738 & ~x745 & ~x749 & ~x767 & ~x772 & ~x776 & ~x777 & ~x779 & ~x780 & ~x782;
assign c7285 =  x379 &  x453 & ~x240 & ~x263 & ~x268 & ~x269 & ~x334;
assign c7287 =  x682;
assign c7291 = ~x72 & ~x129 & ~x347 & ~x423 & ~x432 & ~x450 & ~x634 & ~x654;
assign c7293 =  x465 & ~x334 & ~x361 & ~x362 & ~x389 & ~x390 & ~x395;
assign c7297 =  x512 & ~x379 & ~x407 & ~x421;
assign c7299 =  x111;
assign c7301 =  x123;
assign c7303 =  x511 & ~x186 & ~x348 & ~x451;
assign c7305 =  x71;
assign c7307 =  x275 &  x277 &  x295 &  x296 &  x322 &  x324 &  x353 &  x357 &  x380 &  x384 &  x385 &  x389 &  x413 &  x414 &  x433 &  x442 &  x443 &  x444 &  x463 &  x464 &  x471 &  x514 &  x523 &  x541 &  x543 &  x548 &  x569 &  x570 & ~x3 & ~x10 & ~x11 & ~x26 & ~x33 & ~x34 & ~x37 & ~x43 & ~x44 & ~x47 & ~x54 & ~x57 & ~x60 & ~x63 & ~x77 & ~x104 & ~x128 & ~x130 & ~x141 & ~x146 & ~x150 & ~x152 & ~x155 & ~x172 & ~x176 & ~x208 & ~x228 & ~x230 & ~x253 & ~x261 & ~x279 & ~x284 & ~x307 & ~x309 & ~x311 & ~x318 & ~x341 & ~x363 & ~x368 & ~x393 & ~x661 & ~x672 & ~x673 & ~x674 & ~x687 & ~x689 & ~x700 & ~x715 & ~x740 & ~x744 & ~x746 & ~x748 & ~x753 & ~x754 & ~x760 & ~x768;
assign c7309 =  x247 &  x379 &  x465 &  x473 &  x529 &  x572 &  x573 &  x584 &  x585 &  x613 & ~x0 & ~x11 & ~x64 & ~x72 & ~x75 & ~x101 & ~x145 & ~x148 & ~x231 & ~x251 & ~x281 & ~x284 & ~x343 & ~x391 & ~x420 & ~x660 & ~x685 & ~x688 & ~x701 & ~x716 & ~x718 & ~x737 & ~x746 & ~x753 & ~x773;
assign c7311 =  x248 &  x537 &  x554 &  x555 &  x570 &  x582 &  x583 & ~x17 & ~x20 & ~x29 & ~x32 & ~x44 & ~x49 & ~x54 & ~x65 & ~x67 & ~x73 & ~x93 & ~x95 & ~x106 & ~x124 & ~x127 & ~x130 & ~x133 & ~x163 & ~x169 & ~x199 & ~x200 & ~x255 & ~x262 & ~x280 & ~x283 & ~x308 & ~x338 & ~x340 & ~x364 & ~x397 & ~x448 & ~x616 & ~x619 & ~x634 & ~x650 & ~x652 & ~x659 & ~x662 & ~x666 & ~x671 & ~x672 & ~x689 & ~x706 & ~x713 & ~x720 & ~x734 & ~x742 & ~x748 & ~x751 & ~x760 & ~x774;
assign c7313 =  x249 &  x533 & ~x428 & ~x633;
assign c7315 =  x682;
assign c7317 = ~x418 & ~x423;
assign c7319 =  x681;
assign c7321 =  x330 &  x333 &  x356 &  x357 &  x495 & ~x8 & ~x15 & ~x22 & ~x25 & ~x28 & ~x29 & ~x35 & ~x48 & ~x49 & ~x63 & ~x64 & ~x70 & ~x81 & ~x92 & ~x96 & ~x101 & ~x115 & ~x120 & ~x129 & ~x134 & ~x140 & ~x141 & ~x164 & ~x169 & ~x181 & ~x185 & ~x193 & ~x194 & ~x203 & ~x212 & ~x213 & ~x220 & ~x226 & ~x242 & ~x243 & ~x245 & ~x311 & ~x392 & ~x621 & ~x668 & ~x695 & ~x707 & ~x708 & ~x727 & ~x732 & ~x738 & ~x745 & ~x746 & ~x749 & ~x751 & ~x752 & ~x753 & ~x773 & ~x775 & ~x783;
assign c7323 =  x38 &  x92;
assign c7325 =  x442 &  x534 &  x582 &  x596 &  x610 &  x638;
assign c7327 =  x198;
assign c7329 =  x454 & ~x45 & ~x418;
assign c7333 =  x149;
assign c7335 =  x253;
assign c7337 =  x369 & ~x394;
assign c7343 =  x5;
assign c7345 =  x425 & ~x394 & ~x423;
assign c7347 =  x453 & ~x101 & ~x241 & ~x242 & ~x250 & ~x252 & ~x287 & ~x421 & ~x423 & ~x629 & ~x769;
assign c7349 =  x300 & ~x4 & ~x7 & ~x13 & ~x17 & ~x20 & ~x28 & ~x30 & ~x42 & ~x43 & ~x50 & ~x51 & ~x52 & ~x53 & ~x59 & ~x64 & ~x68 & ~x70 & ~x71 & ~x72 & ~x90 & ~x94 & ~x96 & ~x105 & ~x108 & ~x110 & ~x114 & ~x115 & ~x116 & ~x121 & ~x122 & ~x125 & ~x129 & ~x135 & ~x140 & ~x141 & ~x142 & ~x143 & ~x146 & ~x149 & ~x156 & ~x157 & ~x158 & ~x169 & ~x170 & ~x179 & ~x183 & ~x184 & ~x187 & ~x190 & ~x194 & ~x202 & ~x208 & ~x209 & ~x214 & ~x215 & ~x230 & ~x234 & ~x251 & ~x256 & ~x261 & ~x285 & ~x287 & ~x290 & ~x291 & ~x311 & ~x313 & ~x315 & ~x318 & ~x336 & ~x338 & ~x339 & ~x340 & ~x392 & ~x393 & ~x612 & ~x614 & ~x617 & ~x620 & ~x630 & ~x632 & ~x643 & ~x647 & ~x651 & ~x652 & ~x654 & ~x655 & ~x660 & ~x664 & ~x665 & ~x667 & ~x668 & ~x669 & ~x670 & ~x674 & ~x685 & ~x689 & ~x692 & ~x695 & ~x697 & ~x702 & ~x703 & ~x711 & ~x713 & ~x721 & ~x726 & ~x728 & ~x731 & ~x732 & ~x735 & ~x736 & ~x741 & ~x748 & ~x755 & ~x756 & ~x763 & ~x768 & ~x770 & ~x775 & ~x778 & ~x782 & ~x783;
assign c7351 =  x714;
assign c7353 =  x220 &  x221 &  x247 &  x573 &  x583 &  x611 & ~x16 & ~x197 & ~x198 & ~x715 & ~x739;
assign c7355 =  x285;
assign c7359 =  x540 &  x564 &  x583 &  x584 & ~x605 & ~x659 & ~x695;
assign c7361 = ~x372 & ~x384 & ~x478 & ~x578;
assign c7363 =  x548 &  x553 &  x554 &  x555 &  x569 &  x582 & ~x2 & ~x11 & ~x16 & ~x17 & ~x20 & ~x28 & ~x30 & ~x32 & ~x37 & ~x40 & ~x53 & ~x55 & ~x56 & ~x58 & ~x63 & ~x70 & ~x72 & ~x73 & ~x75 & ~x79 & ~x85 & ~x87 & ~x90 & ~x94 & ~x97 & ~x101 & ~x104 & ~x105 & ~x112 & ~x113 & ~x115 & ~x117 & ~x128 & ~x130 & ~x131 & ~x141 & ~x151 & ~x153 & ~x157 & ~x165 & ~x167 & ~x168 & ~x174 & ~x180 & ~x181 & ~x200 & ~x225 & ~x231 & ~x254 & ~x260 & ~x262 & ~x263 & ~x280 & ~x289 & ~x291 & ~x308 & ~x309 & ~x316 & ~x318 & ~x319 & ~x342 & ~x391 & ~x420 & ~x588 & ~x606 & ~x617 & ~x620 & ~x631 & ~x632 & ~x634 & ~x648 & ~x652 & ~x653 & ~x654 & ~x656 & ~x659 & ~x661 & ~x669 & ~x670 & ~x680 & ~x685 & ~x689 & ~x696 & ~x712 & ~x715 & ~x721 & ~x723 & ~x727 & ~x730 & ~x739 & ~x740 & ~x743 & ~x747 & ~x756 & ~x762 & ~x778 & ~x781 & ~x782;
assign c7365 = ~x353 & ~x398 & ~x477;
assign c7367 = ~x26 & ~x120 & ~x278 & ~x306 & ~x333 & ~x339 & ~x361 & ~x577 & ~x581;
assign c7369 =  x276 &  x301 &  x534 &  x546 &  x547 &  x554 &  x555 &  x556 & ~x60 & ~x65 & ~x74 & ~x89 & ~x94 & ~x101 & ~x153 & ~x252 & ~x290 & ~x317 & ~x346 & ~x373 & ~x391 & ~x397 & ~x399 & ~x423 & ~x476 & ~x634 & ~x646 & ~x660 & ~x671 & ~x688 & ~x689 & ~x704 & ~x716 & ~x771;
assign c7371 =  x572 &  x583 & ~x12 & ~x19 & ~x402 & ~x633 & ~x661 & ~x673 & ~x698;
assign c7373 =  x191;
assign c7375 =  x501 &  x613 &  x628 &  x641 & ~x690;
assign c7377 =  x154 &  x217 &  x573 &  x583 &  x584 &  x611 &  x612;
assign c7379 =  x761;
assign c7383 = ~x241 & ~x263 & ~x268 & ~x269 & ~x339 & ~x390 & ~x555 & ~x570 & ~x582 & ~x584;
assign c7385 =  x398 &  x481 & ~x241 & ~x269 & ~x368;
assign c7387 = ~x82 & ~x349 & ~x434;
assign c7389 =  x178;
assign c7391 =  x249 &  x534 &  x583 &  x584 &  x610 & ~x132 & ~x345 & ~x400 & ~x662 & ~x688 & ~x755;
assign c7393 = ~x10 & ~x278 & ~x336 & ~x394 & ~x395 & ~x417 & ~x418 & ~x419 & ~x579 & ~x608;
assign c7395 =  x12;
assign c7397 =  x136;
assign c7399 =  x426 &  x482 &  x512 &  x514 &  x526 & ~x8 & ~x16 & ~x27 & ~x39 & ~x70 & ~x124 & ~x129 & ~x134 & ~x146 & ~x169 & ~x243 & ~x341 & ~x643 & ~x646 & ~x678 & ~x727 & ~x732 & ~x736 & ~x739 & ~x757 & ~x781;
assign c7401 =  x315;
assign c7403 = ~x187 & ~x269 & ~x270 & ~x388 & ~x390 & ~x607 & ~x617 & ~x633;
assign c7405 =  x628 & ~x429 & ~x690 & ~x717;
assign c7407 =  x711;
assign c7409 =  x285;
assign c7411 =  x557 & ~x457;
assign c7413 =  x777;
assign c7415 =  x220 &  x246 &  x507 &  x549 &  x584 &  x593 &  x611;
assign c7417 =  x286;
assign c7419 =  x203;
assign c7421 =  x485 & ~x416 & ~x443;
assign c7423 =  x246 &  x248 &  x268 &  x269 &  x270 &  x272 &  x275 &  x323 &  x329 &  x385 &  x388 &  x406 &  x413 &  x437 &  x470 &  x471 &  x490 &  x492 &  x495 &  x498 &  x499 &  x515 &  x525 &  x528 &  x548 &  x549 &  x556 &  x570 &  x571 &  x572 & ~x7 & ~x24 & ~x27 & ~x30 & ~x32 & ~x34 & ~x53 & ~x60 & ~x62 & ~x77 & ~x90 & ~x94 & ~x99 & ~x102 & ~x107 & ~x175 & ~x176 & ~x224 & ~x226 & ~x227 & ~x228 & ~x235 & ~x284 & ~x319 & ~x337 & ~x338 & ~x339 & ~x346 & ~x370 & ~x391 & ~x399 & ~x423 & ~x426 & ~x427 & ~x447 & ~x676 & ~x707 & ~x708 & ~x741 & ~x743 & ~x757 & ~x775 & ~x776 & ~x783;
assign c7425 =  x203;
assign c7427 =  x9;
assign c7429 =  x772;
assign c7431 = ~x241 & ~x366 & ~x417 & ~x418 & ~x564 & ~x577 & ~x704;
assign c7433 =  x207;
assign c7435 = ~x214 & ~x320 & ~x405 & ~x449 & ~x462;
assign c7437 =  x482 & ~x444 & ~x446;
assign c7439 =  x261;
assign c7441 = ~x13 & ~x368 & ~x434 & ~x449 & ~x634 & ~x661 & ~x689 & ~x749;
assign c7443 =  x199;
assign c7445 =  x539 &  x557 & ~x384 & ~x401 & ~x477 & ~x479;
assign c7447 =  x309;
assign c7449 =  x60;
assign c7451 =  x712;
assign c7453 =  x240 &  x245 &  x247 &  x270 &  x296 &  x534 &  x549 &  x556 &  x566 &  x570 & ~x88 & ~x97 & ~x143 & ~x161 & ~x254 & ~x291 & ~x401 & ~x646 & ~x674;
assign c7455 =  x410 &  x439 &  x444 & ~x61 & ~x90 & ~x142 & ~x306 & ~x334 & ~x337 & ~x363 & ~x373 & ~x374 & ~x402 & ~x504 & ~x689;
assign c7457 =  x572 &  x600 &  x652 & ~x429;
assign c7459 =  x269 &  x276 &  x297 &  x301 &  x303 &  x329 &  x332 &  x357 &  x463 &  x515 &  x520 &  x528 &  x534 &  x549 &  x564 &  x568 &  x569 &  x571 & ~x0 & ~x30 & ~x32 & ~x44 & ~x58 & ~x75 & ~x78 & ~x81 & ~x92 & ~x94 & ~x98 & ~x104 & ~x114 & ~x129 & ~x130 & ~x133 & ~x150 & ~x153 & ~x155 & ~x228 & ~x229 & ~x260 & ~x279 & ~x282 & ~x292 & ~x345 & ~x347 & ~x396 & ~x399 & ~x660 & ~x661 & ~x688 & ~x689 & ~x701 & ~x706 & ~x708 & ~x717 & ~x733 & ~x743 & ~x750 & ~x768;
assign c7461 =  x45;
assign c7463 =  x93;
assign c7465 =  x653 &  x656;
assign c7467 =  x47;
assign c7469 =  x18;
assign c7471 =  x282;
assign c7473 =  x249 &  x268 &  x277 &  x302 &  x354 &  x379 &  x384 &  x385 &  x412 &  x434 &  x438 &  x461 &  x462 &  x493 &  x500 &  x501 &  x507 &  x521 &  x522 &  x529 &  x543 &  x545 & ~x4 & ~x6 & ~x18 & ~x20 & ~x23 & ~x30 & ~x35 & ~x37 & ~x53 & ~x56 & ~x59 & ~x65 & ~x69 & ~x70 & ~x71 & ~x72 & ~x80 & ~x96 & ~x113 & ~x122 & ~x131 & ~x133 & ~x159 & ~x173 & ~x174 & ~x199 & ~x201 & ~x251 & ~x282 & ~x283 & ~x286 & ~x290 & ~x309 & ~x313 & ~x373 & ~x399 & ~x400 & ~x421 & ~x645 & ~x656 & ~x659 & ~x660 & ~x662 & ~x663 & ~x670 & ~x672 & ~x689 & ~x691 & ~x728 & ~x732 & ~x736 & ~x752 & ~x770 & ~x777;
assign c7475 =  x529 & ~x423 & ~x450 & ~x458;
assign c7477 =  x191 &  x611;
assign c7479 =  x773;
assign c7481 =  x239 &  x491 &  x537 &  x597 &  x611 & ~x153 & ~x399;
assign c7483 =  x717;
assign c7487 =  x195;
assign c7489 = ~x380 & ~x381;
assign c7491 =  x425 & ~x350 & ~x394;
assign c7493 =  x528 &  x556 &  x557 & ~x1 & ~x31 & ~x38 & ~x48 & ~x88 & ~x92 & ~x234 & ~x379 & ~x559 & ~x716;
assign c7495 =  x499 & ~x5 & ~x22 & ~x36 & ~x57 & ~x60 & ~x90 & ~x96 & ~x102 & ~x116 & ~x121 & ~x124 & ~x150 & ~x156 & ~x157 & ~x182 & ~x200 & ~x214 & ~x220 & ~x224 & ~x226 & ~x229 & ~x230 & ~x231 & ~x254 & ~x259 & ~x311 & ~x316 & ~x335 & ~x366 & ~x394 & ~x395 & ~x421 & ~x578 & ~x591 & ~x600 & ~x606 & ~x607 & ~x625 & ~x630 & ~x644 & ~x655 & ~x667 & ~x669 & ~x676 & ~x680 & ~x682 & ~x696 & ~x711 & ~x746 & ~x749 & ~x778;
assign c7497 =  x105;
assign c7499 = ~x333 & ~x386 & ~x394;
assign c80 =  x427 &  x537 &  x567 & ~x17 & ~x47 & ~x50 & ~x60 & ~x70 & ~x77 & ~x139 & ~x195;
assign c82 =  x578 &  x579 & ~x43 & ~x59 & ~x62 & ~x66 & ~x72 & ~x85 & ~x89 & ~x101 & ~x532 & ~x689 & ~x715 & ~x745;
assign c84 =  x97 &  x163 &  x499 & ~x646 & ~x754;
assign c86 =  x571 & ~x11 & ~x94 & ~x217 & ~x294 & ~x301 & ~x316 & ~x322 & ~x330 & ~x331 & ~x445 & ~x530;
assign c88 = ~x488 & ~x514 & ~x543 & ~x571;
assign c810 =  x290 &  x295 &  x317 &  x322 &  x327 &  x353 &  x355 &  x372 &  x374 &  x377 &  x402 &  x411 & ~x7 & ~x34 & ~x35 & ~x52 & ~x56 & ~x84 & ~x86 & ~x137 & ~x199 & ~x225 & ~x252 & ~x309 & ~x391 & ~x448 & ~x508 & ~x536 & ~x564 & ~x728 & ~x754 & ~x757 & ~x761 & ~x763 & ~x780;
assign c812 =  x213 & ~x652 & ~x653 & ~x654 & ~x666 & ~x681 & ~x684 & ~x695;
assign c814 =  x41 &  x719 & ~x9 & ~x10 & ~x11 & ~x12 & ~x19 & ~x144 & ~x227 & ~x228 & ~x256;
assign c816 =  x372 &  x387 &  x428 &  x488 &  x499 &  x523 &  x527 &  x555 &  x583 &  x628 &  x631 &  x639 &  x662 &  x665 &  x666 &  x686 &  x687 &  x693 &  x714 & ~x0 & ~x773 & ~x775 & ~x778 & ~x780;
assign c818 =  x306 & ~x656 & ~x691 & ~x741;
assign c820 =  x631 &  x632 & ~x10 & ~x35 & ~x49 & ~x53 & ~x64 & ~x77 & ~x80 & ~x90 & ~x132 & ~x145 & ~x171 & ~x217 & ~x220 & ~x231 & ~x778;
assign c822 =  x438 & ~x11 & ~x28 & ~x53 & ~x98 & ~x103 & ~x194 & ~x418 & ~x557;
assign c824 =  x142;
assign c826 = ~x122 & ~x371 & ~x399 & ~x407 & ~x410 & ~x442;
assign c828 =  x109;
assign c830 =  x252;
assign c832 =  x167;
assign c834 =  x356 & ~x9 & ~x11 & ~x63 & ~x78 & ~x104 & ~x107 & ~x126 & ~x154 & ~x161 & ~x189 & ~x201 & ~x212 & ~x218 & ~x220 & ~x240;
assign c836 =  x538 &  x595 & ~x11 & ~x53 & ~x63 & ~x90 & ~x128 & ~x135 & ~x167 & ~x224 & ~x363;
assign c838 =  x474 & ~x450 & ~x779;
assign c840 =  x186 & ~x442 & ~x485 & ~x486;
assign c842 =  x281;
assign c844 =  x458 & ~x36 & ~x37 & ~x48 & ~x60 & ~x62 & ~x77 & ~x89 & ~x92 & ~x105 & ~x124 & ~x134 & ~x162 & ~x173 & ~x184 & ~x185 & ~x193 & ~x420;
assign c846 =  x260 &  x441 &  x454 &  x483 & ~x12 & ~x27 & ~x35 & ~x281 & ~x751 & ~x753 & ~x754 & ~x768 & ~x769 & ~x770;
assign c848 =  x326 & ~x10 & ~x44 & ~x50 & ~x78 & ~x612 & ~x637 & ~x724;
assign c850 =  x602 &  x603 &  x604 & ~x12 & ~x135 & ~x151 & ~x273;
assign c852 =  x589 & ~x17 & ~x642 & ~x729;
assign c854 =  x620 & ~x2 & ~x9 & ~x64 & ~x70 & ~x78 & ~x79 & ~x81 & ~x92 & ~x755;
assign c856 =  x421 &  x505;
assign c858 =  x606 &  x635 & ~x12 & ~x26 & ~x35 & ~x39 & ~x47 & ~x50 & ~x76 & ~x93 & ~x250 & ~x307 & ~x504 & ~x562 & ~x644 & ~x759;
assign c860 =  x585 & ~x395;
assign c862 =  x306 &  x334 & ~x107 & ~x651;
assign c864 =  x364;
assign c866 =  x316 &  x426 &  x676 &  x705 &  x708 &  x713 &  x716 &  x720 &  x734 &  x738 &  x739 &  x742 &  x744;
assign c868 = ~x17 & ~x78 & ~x515 & ~x540 & ~x627 & ~x735;
assign c870 =  x538 & ~x19 & ~x47 & ~x103 & ~x106 & ~x246 & ~x259 & ~x303 & ~x358;
assign c872 =  x538 & ~x133 & ~x270;
assign c874 =  x232 &  x378 &  x499 &  x668 &  x735 & ~x673;
assign c876 =  x344 &  x401 &  x438 &  x439 &  x442 &  x484 &  x499 &  x518 &  x523 &  x525 &  x545 &  x547 &  x552 &  x595 &  x599 &  x610 &  x611 &  x625 &  x630 &  x637 &  x657 &  x664 &  x665 &  x667 &  x687 &  x695 &  x710 &  x721 &  x722 &  x736 & ~x4 & ~x31 & ~x59 & ~x114 & ~x197 & ~x699 & ~x727 & ~x728 & ~x756;
assign c878 =  x281;
assign c880 =  x14 & ~x70 & ~x98 & ~x118 & ~x531 & ~x561;
assign c882 =  x366 &  x619;
assign c884 =  x354 & ~x45 & ~x46 & ~x224 & ~x416;
assign c886 = ~x11 & ~x16 & ~x105 & ~x218 & ~x294 & ~x316 & ~x349 & ~x350 & ~x357 & ~x445 & ~x528;
assign c888 =  x262 & ~x579 & ~x580 & ~x626 & ~x627 & ~x682;
assign c890 =  x95 &  x146 &  x148 &  x151 &  x201 &  x202 &  x229 &  x230 &  x244 &  x323 &  x371 &  x427 &  x510 &  x525 &  x565 &  x566 &  x602 &  x637 &  x649 &  x706 &  x707 &  x712 &  x713 & ~x253 & ~x699 & ~x754;
assign c892 =  x591 & ~x11 & ~x36 & ~x47 & ~x71 & ~x106 & ~x224 & ~x672;
assign c894 =  x439 &  x460 &  x466 &  x485 &  x495 &  x513 &  x514 &  x521 &  x522 &  x541 &  x542 &  x547 &  x548 & ~x1 & ~x7 & ~x9 & ~x10 & ~x20 & ~x30 & ~x31 & ~x33 & ~x51 & ~x56 & ~x58 & ~x59 & ~x60 & ~x77 & ~x78 & ~x109 & ~x110 & ~x111 & ~x112 & ~x118 & ~x135 & ~x137 & ~x141 & ~x164 & ~x168 & ~x169 & ~x172 & ~x200 & ~x223 & ~x226 & ~x248 & ~x254 & ~x280 & ~x307 & ~x309 & ~x394 & ~x395 & ~x419 & ~x422 & ~x423 & ~x424 & ~x506 & ~x643 & ~x671 & ~x700 & ~x705 & ~x727 & ~x755 & ~x762 & ~x779 & ~x780 & ~x782 & ~x783;
assign c896 = ~x9 & ~x10 & ~x11 & ~x12 & ~x16 & ~x17 & ~x18 & ~x19 & ~x37 & ~x86 & ~x87 & ~x557 & ~x576 & ~x582 & ~x728 & ~x754 & ~x768 & ~x769;
assign c898 =  x532;
assign c8100 =  x547 &  x658 & ~x18 & ~x79 & ~x220 & ~x238 & ~x304;
assign c8102 =  x317 &  x327 &  x522 & ~x698 & ~x711 & ~x712 & ~x719 & ~x751 & ~x783;
assign c8104 =  x395 &  x566 & ~x46 & ~x47 & ~x60 & ~x88;
assign c8106 =  x421 &  x578;
assign c8108 =  x357 &  x372 &  x412 &  x433 &  x488 &  x512 &  x539 &  x543 &  x548 &  x571 &  x572 &  x628 &  x630 &  x631 &  x683 &  x708 &  x714 &  x720 & ~x6 & ~x60 & ~x84 & ~x143 & ~x194 & ~x306 & ~x307 & ~x448;
assign c8110 =  x308;
assign c8112 =  x232 & ~x17 & ~x531 & ~x712 & ~x722 & ~x751 & ~x752 & ~x754 & ~x764 & ~x776 & ~x779;
assign c8114 =  x3;
assign c8116 =  x310 & ~x735 & ~x745;
assign c8118 =  x224;
assign c8122 =  x764 & ~x463;
assign c8124 =  x417 &  x500 & ~x36 & ~x46 & ~x104 & ~x121 & ~x164 & ~x653 & ~x657;
assign c8126 = ~x95 & ~x134 & ~x371 & ~x655 & ~x656 & ~x657 & ~x661 & ~x685 & ~x697;
assign c8128 =  x550 & ~x38 & ~x295;
assign c8130 =  x49 &  x565 &  x705 &  x707;
assign c8132 =  x569 &  x579 &  x596 &  x624 &  x635 &  x660 &  x684 &  x690 &  x713 &  x714 &  x715 &  x718 & ~x1 & ~x6 & ~x7 & ~x20 & ~x25 & ~x30 & ~x36 & ~x60 & ~x63 & ~x64 & ~x91 & ~x135 & ~x137 & ~x144 & ~x165 & ~x220 & ~x281 & ~x306 & ~x309 & ~x390 & ~x728;
assign c8134 =  x381 & ~x39 & ~x73 & ~x130 & ~x240 & ~x425;
assign c8136 =  x454 &  x463 &  x594 & ~x750 & ~x769;
assign c8138 =  x372 &  x398 &  x523 & ~x2 & ~x22 & ~x48 & ~x53 & ~x64 & ~x68 & ~x111 & ~x254 & ~x532;
assign c8140 =  x625 &  x649 & ~x30 & ~x139 & ~x336 & ~x749 & ~x751 & ~x753 & ~x759 & ~x769 & ~x770 & ~x772 & ~x773 & ~x779;
assign c8142 =  x572 & ~x94 & ~x101 & ~x111 & ~x129 & ~x215 & ~x218;
assign c8144 =  x400 &  x544 &  x682 &  x684 & ~x19 & ~x88 & ~x339 & ~x564;
assign c8146 =  x425 &  x676 &  x718 &  x719 &  x734 & ~x589;
assign c8148 =  x138 & ~x106;
assign c8150 =  x63 &  x147 &  x150 &  x180 &  x454 &  x482 &  x593;
assign c8152 =  x745 & ~x210 & ~x229 & ~x289;
assign c8154 =  x559;
assign c8156 =  x13 &  x682 & ~x69;
assign c8158 =  x348 &  x372 &  x544 &  x579 &  x582 &  x609 & ~x38 & ~x48 & ~x49 & ~x57 & ~x62 & ~x63 & ~x66 & ~x78 & ~x504 & ~x560 & ~x755 & ~x756 & ~x780 & ~x782;
assign c8160 =  x397 & ~x23 & ~x62 & ~x88 & ~x98 & ~x99 & ~x108 & ~x588 & ~x755 & ~x778;
assign c8162 =  x569 &  x605 &  x606 &  x607 &  x631 &  x661 &  x662 &  x663 & ~x3 & ~x19 & ~x22 & ~x45 & ~x46 & ~x61 & ~x76 & ~x79 & ~x89 & ~x108 & ~x134 & ~x197 & ~x250 & ~x274 & ~x281 & ~x307 & ~x365;
assign c8164 =  x575 &  x628 & ~x182 & ~x216;
assign c8166 =  x599 &  x634 & ~x122 & ~x134 & ~x160 & ~x177;
assign c8168 =  x514 &  x516 &  x522 &  x550 & ~x6 & ~x18 & ~x24 & ~x30 & ~x35 & ~x52 & ~x59 & ~x63 & ~x113 & ~x114 & ~x130 & ~x154 & ~x168 & ~x192 & ~x193 & ~x392 & ~x448 & ~x449 & ~x476 & ~x504;
assign c8170 =  x365;
assign c8172 =  x277 &  x329 &  x528 &  x583 & ~x753;
assign c8174 =  x418 &  x554;
assign c8176 =  x266 & ~x449 & ~x477 & ~x664 & ~x684 & ~x686 & ~x719 & ~x734 & ~x742;
assign c8178 =  x340 & ~x36 & ~x64 & ~x90 & ~x126 & ~x173 & ~x420;
assign c8180 =  x41 &  x50;
assign c8182 =  x14 & ~x69 & ~x104;
assign c8184 =  x192 &  x220 &  x631 &  x638 &  x694 & ~x774 & ~x781;
assign c8186 = ~x127 & ~x369 & ~x634 & ~x651 & ~x656 & ~x685 & ~x739;
assign c8188 =  x429 &  x494 &  x495 &  x518 &  x522 &  x542 &  x546 &  x547 &  x550 &  x551 &  x635 &  x691 & ~x5 & ~x32 & ~x36 & ~x49 & ~x63 & ~x90 & ~x106 & ~x107 & ~x114 & ~x134 & ~x168 & ~x193 & ~x220 & ~x307 & ~x420 & ~x474 & ~x531 & ~x589 & ~x779;
assign c8190 =  x317 &  x319 &  x327 &  x328 &  x330 &  x389 &  x442 &  x443 &  x471 &  x496 &  x497 &  x526 &  x554 & ~x8 & ~x9 & ~x10 & ~x111 & ~x727 & ~x753 & ~x754 & ~x783;
assign c8192 = ~x246 & ~x273 & ~x316 & ~x349 & ~x416 & ~x443;
assign c8194 =  x500 & ~x44 & ~x143;
assign c8196 =  x300 &  x304 &  x352 &  x372 &  x385 &  x458 &  x469 &  x470 &  x499 &  x526 &  x527 & ~x699 & ~x752 & ~x776 & ~x778;
assign c8198 =  x684 &  x688 & ~x16 & ~x247 & ~x288 & ~x289 & ~x304;
assign c8200 =  x489 & ~x2 & ~x10 & ~x17 & ~x21 & ~x28 & ~x32 & ~x36 & ~x37 & ~x48 & ~x66 & ~x82 & ~x90 & ~x104 & ~x107 & ~x111 & ~x114 & ~x118 & ~x148 & ~x168 & ~x196 & ~x254 & ~x424 & ~x621 & ~x700 & ~x731 & ~x756 & ~x757 & ~x778 & ~x779;
assign c8202 =  x448;
assign c8204 =  x247 &  x276 &  x334 &  x499 &  x524 &  x526 &  x527 &  x553 &  x555;
assign c8206 =  x476;
assign c8208 = ~x4 & ~x10 & ~x11 & ~x47 & ~x77 & ~x132 & ~x145 & ~x146 & ~x164 & ~x176 & ~x184 & ~x190 & ~x192 & ~x218 & ~x265 & ~x266 & ~x269 & ~x273 & ~x307 & ~x644 & ~x781;
assign c8210 =  x336;
assign c8212 =  x470 &  x473 & ~x77 & ~x449 & ~x682 & ~x737;
assign c8214 =  x336;
assign c8216 =  x223;
assign c8218 =  x411 &  x435 &  x439 & ~x24 & ~x35 & ~x90 & ~x141 & ~x174 & ~x204 & ~x248;
assign c8220 =  x589 & ~x38 & ~x108;
assign c8222 = ~x7 & ~x8 & ~x9 & ~x10 & ~x18 & ~x23 & ~x41 & ~x42 & ~x50 & ~x53 & ~x60 & ~x65 & ~x68 & ~x69 & ~x70 & ~x80 & ~x81 & ~x333 & ~x505 & ~x532 & ~x559 & ~x615 & ~x644;
assign c8224 =  x177 &  x399 &  x439 &  x640 &  x694 &  x695 &  x707 & ~x615 & ~x698;
assign c8226 =  x56;
assign c8228 =  x409 &  x463 &  x470 &  x527 &  x574 &  x583 &  x628 &  x639 &  x667 &  x688 &  x690 &  x692 &  x694 &  x707 & ~x31 & ~x778 & ~x779;
assign c8230 =  x610 & ~x106 & ~x210 & ~x306;
assign c8232 =  x25;
assign c8234 =  x346 &  x353 & ~x47 & ~x80 & ~x394 & ~x658 & ~x685;
assign c8236 =  x358 &  x526 & ~x11 & ~x79 & ~x116 & ~x118 & ~x156;
assign c8238 =  x109;
assign c8240 = ~x106 & ~x331 & ~x343 & ~x434 & ~x441 & ~x498 & ~x512;
assign c8242 =  x506 &  x649 & ~x37 & ~x48 & ~x111 & ~x728;
assign c8244 = ~x10 & ~x11 & ~x18 & ~x78 & ~x92 & ~x164 & ~x175 & ~x187 & ~x209 & ~x210 & ~x220 & ~x238 & ~x245 & ~x248 & ~x306 & ~x473;
assign c8246 =  x513 &  x548 & ~x10 & ~x11 & ~x20 & ~x53 & ~x68 & ~x150 & ~x185 & ~x204 & ~x218 & ~x249;
assign c8248 =  x718 & ~x321;
assign c8250 =  x372 &  x377 &  x383 &  x400 &  x402 &  x521 & ~x6 & ~x10 & ~x18 & ~x19 & ~x22 & ~x54 & ~x83 & ~x87 & ~x92 & ~x107 & ~x112 & ~x168 & ~x254 & ~x394 & ~x477 & ~x505 & ~x778;
assign c8252 = ~x18 & ~x538 & ~x539 & ~x541 & ~x567 & ~x570 & ~x597 & ~x708 & ~x711;
assign c8254 =  x4;
assign c8256 =  x14 &  x622 &  x715 &  x736;
assign c8258 = ~x413 & ~x429 & ~x434 & ~x437 & ~x511;
assign c8260 = ~x45 & ~x62 & ~x64 & ~x67 & ~x74 & ~x91 & ~x92 & ~x103 & ~x132 & ~x218 & ~x652 & ~x657 & ~x664 & ~x681 & ~x684 & ~x685 & ~x707 & ~x709 & ~x712 & ~x734 & ~x739;
assign c8262 =  x309;
assign c8264 = ~x12 & ~x17 & ~x93 & ~x120 & ~x126 & ~x132 & ~x134 & ~x230 & ~x293 & ~x316 & ~x322 & ~x474 & ~x528 & ~x669;
assign c8266 = ~x16 & ~x67 & ~x76 & ~x79 & ~x85 & ~x120 & ~x159 & ~x164 & ~x176 & ~x202 & ~x204 & ~x259 & ~x274 & ~x302 & ~x303 & ~x332 & ~x390 & ~x417 & ~x421 & ~x445 & ~x449 & ~x477 & ~x499 & ~x529 & ~x561 & ~x585;
assign c8268 =  x90 &  x229 &  x357 &  x410 &  x463 &  x598 &  x705 &  x707 &  x712 & ~x83 & ~x197 & ~x419 & ~x643;
assign c8270 = ~x10 & ~x42 & ~x46 & ~x54 & ~x399 & ~x540 & ~x557 & ~x582 & ~x585 & ~x755 & ~x779;
assign c8272 =  x684 &  x717 & ~x201 & ~x212 & ~x221;
assign c8274 =  x31 &  x140;
assign c8276 =  x280;
assign c8278 =  x308;
assign c8280 = ~x16 & ~x161 & ~x162 & ~x458 & ~x467 & ~x485 & ~x496;
assign c8282 =  x224;
assign c8284 =  x542 &  x577 & ~x266 & ~x274;
assign c8286 =  x706 &  x707 &  x711 &  x718 &  x735 &  x737 & ~x144 & ~x164 & ~x200 & ~x646;
assign c8288 =  x532 &  x705;
assign c8290 =  x351 & ~x137 & ~x196 & ~x238 & ~x244 & ~x588;
assign c8292 =  x290 &  x327 & ~x23 & ~x394 & ~x654;
assign c8294 =  x570 &  x571 &  x577 &  x599 &  x601 &  x602 &  x604 &  x607 & ~x1 & ~x29 & ~x35 & ~x50 & ~x78 & ~x106 & ~x108 & ~x221 & ~x238 & ~x246 & ~x301 & ~x306 & ~x757 & ~x758 & ~x782;
assign c8296 =  x356 & ~x493 & ~x548;
assign c8298 = ~x6 & ~x10 & ~x11 & ~x18 & ~x32 & ~x35 & ~x38 & ~x39 & ~x46 & ~x49 & ~x64 & ~x65 & ~x66 & ~x75 & ~x81 & ~x103 & ~x104 & ~x108 & ~x117 & ~x119 & ~x121 & ~x177 & ~x203 & ~x204 & ~x246 & ~x247 & ~x265 & ~x272 & ~x273 & ~x293 & ~x305;
assign c8300 =  x452 &  x509 &  x537 &  x538 &  x614 &  x621 & ~x76;
assign c8304 =  x400 &  x411 &  x548 & ~x36 & ~x75 & ~x107 & ~x119 & ~x121 & ~x134 & ~x193 & ~x221 & ~x223 & ~x504 & ~x757 & ~x777;
assign c8306 =  x308;
assign c8308 =  x364;
assign c8310 =  x314 & ~x20 & ~x44 & ~x48 & ~x57 & ~x73 & ~x615 & ~x702 & ~x715 & ~x721 & ~x723 & ~x728 & ~x729 & ~x731 & ~x733 & ~x739 & ~x740 & ~x753 & ~x768 & ~x780;
assign c8312 =  x714 & ~x11 & ~x19 & ~x62 & ~x77 & ~x86 & ~x107 & ~x108 & ~x145 & ~x182 & ~x222 & ~x229;
assign c8314 =  x220 &  x317 &  x359 & ~x169 & ~x309 & ~x392 & ~x753 & ~x773 & ~x774 & ~x778;
assign c8316 = ~x9 & ~x11 & ~x18 & ~x50 & ~x107 & ~x273 & ~x297 & ~x298 & ~x301 & ~x302 & ~x316 & ~x357 & ~x440 & ~x529;
assign c8318 = ~x3 & ~x12 & ~x50 & ~x56 & ~x59 & ~x63 & ~x65 & ~x67 & ~x74 & ~x103 & ~x114 & ~x165 & ~x177 & ~x188 & ~x189 & ~x194 & ~x204 & ~x258 & ~x259 & ~x302 & ~x305 & ~x333 & ~x335 & ~x337 & ~x362 & ~x472 & ~x474 & ~x700 & ~x757 & ~x758 & ~x783;
assign c8320 =  x570 & ~x162 & ~x345 & ~x349;
assign c8322 =  x558 &  x578 & ~x75 & ~x535;
assign c8324 =  x599 &  x605 &  x636 & ~x1 & ~x5 & ~x8 & ~x19 & ~x37 & ~x64 & ~x78 & ~x88 & ~x92 & ~x106 & ~x108 & ~x115 & ~x118 & ~x146 & ~x147 & ~x165 & ~x170 & ~x193 & ~x199 & ~x279 & ~x307;
assign c8326 =  x51;
assign c8328 =  x695 &  x735 &  x737 & ~x672 & ~x771 & ~x772 & ~x773 & ~x779;
assign c8330 =  x555 & ~x89 & ~x108 & ~x128 & ~x533 & ~x588;
assign c8332 =  x475;
assign c8334 = ~x24 & ~x31 & ~x41 & ~x48 & ~x49 & ~x52 & ~x60 & ~x63 & ~x65 & ~x77 & ~x98 & ~x100 & ~x126 & ~x129 & ~x132 & ~x140 & ~x170;
assign c8336 =  x325 &  x326 &  x327 &  x356 &  x411 &  x412 & ~x7 & ~x31 & ~x43 & ~x51 & ~x54 & ~x64 & ~x225 & ~x534 & ~x560 & ~x673 & ~x749 & ~x754 & ~x757 & ~x781;
assign c8338 =  x400 &  x439 &  x569 &  x624 &  x631 & ~x3 & ~x8 & ~x9 & ~x136 & ~x141 & ~x162 & ~x169 & ~x200 & ~x279 & ~x282 & ~x362 & ~x391 & ~x416 & ~x418 & ~x421 & ~x422 & ~x504 & ~x532 & ~x536 & ~x562 & ~x587 & ~x615 & ~x645 & ~x648 & ~x667 & ~x757;
assign c8340 = ~x70 & ~x267 & ~x291 & ~x321 & ~x327 & ~x385 & ~x444;
assign c8342 =  x300 &  x301 &  x351 &  x375 &  x377 &  x378 &  x380 &  x381 &  x467 &  x490 &  x495 & ~x25 & ~x28 & ~x81 & ~x84 & ~x143 & ~x166 & ~x199 & ~x618 & ~x699 & ~x733;
assign c8344 =  x523 &  x524 &  x580 & ~x47 & ~x48 & ~x62 & ~x106 & ~x218 & ~x220 & ~x266;
assign c8346 =  x456 &  x510 &  x576 &  x666 &  x712 &  x734 &  x735 &  x737 & ~x754 & ~x775 & ~x776 & ~x778 & ~x780;
assign c8348 =  x766 & ~x17 & ~x265;
assign c8350 = ~x39 & ~x92 & ~x101 & ~x107 & ~x129 & ~x372 & ~x377 & ~x595;
assign c8352 =  x427 &  x493 &  x496 &  x550 & ~x35 & ~x37 & ~x40 & ~x64 & ~x78 & ~x168 & ~x200 & ~x253 & ~x281 & ~x364 & ~x508 & ~x755 & ~x783;
assign c8354 =  x512 &  x637 & ~x10 & ~x19 & ~x64 & ~x80 & ~x88 & ~x112 & ~x119 & ~x249 & ~x250 & ~x361;
assign c8356 =  x663 & ~x11 & ~x47 & ~x134 & ~x163 & ~x185;
assign c8358 =  x252;
assign c8360 =  x402 &  x543 &  x579 &  x580 &  x666 &  x708 & ~x6 & ~x12 & ~x20 & ~x21 & ~x24 & ~x35 & ~x36 & ~x59 & ~x138 & ~x199;
assign c8362 =  x234 &  x286 &  x427 &  x511 &  x704 &  x708 &  x717 &  x721;
assign c8364 =  x344 &  x702 &  x706 & ~x725;
assign c8366 =  x415 & ~x11 & ~x17 & ~x20 & ~x45 & ~x48 & ~x51 & ~x61 & ~x62 & ~x63 & ~x64 & ~x77 & ~x78 & ~x107 & ~x158 & ~x534 & ~x779;
assign c8368 = ~x9 & ~x36 & ~x46 & ~x70 & ~x106 & ~x154 & ~x238 & ~x244 & ~x273 & ~x294 & ~x295 & ~x305 & ~x442;
assign c8370 =  x349 &  x372 &  x375 &  x380 &  x405 &  x439 &  x493 &  x519 &  x521 &  x523 &  x553 & ~x32 & ~x58 & ~x86 & ~x111 & ~x139 & ~x252 & ~x643 & ~x644 & ~x697 & ~x698 & ~x750 & ~x751 & ~x755 & ~x772 & ~x773 & ~x775 & ~x776 & ~x780 & ~x782;
assign c8372 =  x375 &  x552 &  x649 & ~x36 & ~x39 & ~x65;
assign c8374 = ~x12 & ~x58 & ~x79 & ~x93 & ~x115 & ~x118 & ~x162 & ~x200 & ~x201 & ~x238 & ~x244 & ~x266 & ~x335 & ~x448 & ~x534;
assign c8376 =  x482 &  x529 &  x539 &  x566 &  x574 &  x622 &  x634 &  x649 &  x659;
assign c8378 =  x195;
assign c8380 =  x707 & ~x36 & ~x64 & ~x70 & ~x107 & ~x198;
assign c8382 =  x459 &  x469 & ~x35 & ~x108 & ~x182 & ~x560;
assign c8384 =  x309 & ~x218 & ~x679;
assign c8386 =  x513 &  x548 & ~x37 & ~x39 & ~x60 & ~x78 & ~x94 & ~x118 & ~x136 & ~x215 & ~x243 & ~x477 & ~x778;
assign c8388 =  x145 &  x151 &  x205 &  x453 &  x481;
assign c8390 =  x291 &  x297 &  x345 &  x357 &  x402 &  x416 &  x483 &  x495 &  x498 &  x569 &  x610 &  x626 &  x637 &  x638 &  x677 &  x679 & ~x25 & ~x727 & ~x781;
assign c8392 =  x649 & ~x17 & ~x60 & ~x62 & ~x88 & ~x107 & ~x114 & ~x696;
assign c8394 =  x141;
assign c8396 =  x276 &  x498 &  x527 & ~x614;
assign c8398 =  x705 & ~x135 & ~x275;
assign c8400 =  x234 & ~x3 & ~x6 & ~x11 & ~x39 & ~x43 & ~x46 & ~x47 & ~x48 & ~x51 & ~x52 & ~x77 & ~x113 & ~x691 & ~x703 & ~x710 & ~x712 & ~x738 & ~x743 & ~x750 & ~x752 & ~x753 & ~x768 & ~x773;
assign c8402 =  x276 &  x289 &  x290 &  x301 &  x302 &  x303 &  x304 &  x317 &  x332 &  x345 &  x360 &  x379 &  x415 & ~x140 & ~x167 & ~x279 & ~x393 & ~x560 & ~x672 & ~x780;
assign c8404 =  x559;
assign c8406 =  x291 &  x356 &  x380 &  x383 &  x403 &  x409 &  x412 &  x466 & ~x19 & ~x47 & ~x53 & ~x75 & ~x84 & ~x226 & ~x560 & ~x668 & ~x696 & ~x730 & ~x749 & ~x779 & ~x781;
assign c8408 =  x602 &  x633 & ~x105 & ~x149 & ~x726;
assign c8410 =  x651 & ~x36 & ~x46 & ~x75 & ~x132 & ~x133 & ~x163 & ~x164 & ~x238 & ~x250;
assign c8412 =  x176 &  x343 &  x370 &  x400 &  x401 &  x427 &  x469 &  x484 &  x495 & ~x24 & ~x58 & ~x753 & ~x771 & ~x773 & ~x778 & ~x783;
assign c8414 =  x303 &  x343 &  x417 &  x677 &  x694;
assign c8416 =  x85;
assign c8418 =  x547 &  x602 &  x604 &  x607 &  x658 & ~x18 & ~x35 & ~x105 & ~x162 & ~x274 & ~x361;
assign c8420 =  x262 & ~x568 & ~x597 & ~x680 & ~x707 & ~x711;
assign c8422 = ~x42 & ~x50 & ~x62 & ~x67 & ~x71 & ~x78 & ~x80 & ~x99 & ~x132 & ~x268 & ~x531 & ~x654 & ~x657 & ~x660 & ~x661 & ~x665 & ~x681 & ~x682 & ~x685 & ~x688 & ~x692 & ~x711 & ~x714 & ~x721 & ~x722 & ~x737;
assign c8424 =  x500 & ~x164 & ~x772;
assign c8426 =  x263 &  x270 &  x271 & ~x601 & ~x724;
assign c8428 =  x271 &  x276 &  x301 &  x304 &  x319 &  x322 &  x469 &  x526 &  x527 &  x528 &  x551 &  x554 & ~x746 & ~x748 & ~x750 & ~x779;
assign c8430 = ~x372 & ~x508 & ~x511 & ~x597 & ~x627 & ~x675;
assign c8432 = ~x1 & ~x10 & ~x11 & ~x29 & ~x34 & ~x37 & ~x38 & ~x46 & ~x47 & ~x50 & ~x54 & ~x61 & ~x62 & ~x64 & ~x76 & ~x78 & ~x89 & ~x90 & ~x91 & ~x103 & ~x104 & ~x105 & ~x106 & ~x107 & ~x111 & ~x114 & ~x115 & ~x120 & ~x134 & ~x138 & ~x140 & ~x161 & ~x162 & ~x163 & ~x164 & ~x165 & ~x169 & ~x170 & ~x175 & ~x176 & ~x182 & ~x190 & ~x201 & ~x211 & ~x217 & ~x218 & ~x219 & ~x220 & ~x249 & ~x251 & ~x258 & ~x337 & ~x363;
assign c8434 =  x448;
assign c8436 =  x395 &  x650 &  x653 &  x677 &  x680 &  x681 &  x707 &  x713 & ~x252 & ~x337 & ~x754;
assign c8440 = ~x10 & ~x12 & ~x38 & ~x47 & ~x65 & ~x73 & ~x74 & ~x191 & ~x259 & ~x271 & ~x272 & ~x299 & ~x405 & ~x442 & ~x530;
assign c8442 = ~x69 & ~x154 & ~x164 & ~x174 & ~x187 & ~x240 & ~x268 & ~x294 & ~x501;
assign c8444 =  x343 &  x344 &  x356 &  x519 &  x524 &  x546 & ~x38 & ~x53 & ~x57 & ~x63 & ~x77 & ~x85 & ~x171 & ~x729 & ~x731 & ~x762;
assign c8446 = ~x0 & ~x8 & ~x9 & ~x10 & ~x12 & ~x16 & ~x17 & ~x26 & ~x36 & ~x45 & ~x47 & ~x48 & ~x51 & ~x62 & ~x75 & ~x93 & ~x102 & ~x105 & ~x107 & ~x115 & ~x120 & ~x132 & ~x136 & ~x140 & ~x158 & ~x161 & ~x173 & ~x176 & ~x187 & ~x188 & ~x193 & ~x196 & ~x203 & ~x220 & ~x366 & ~x394 & ~x425 & ~x450 & ~x476 & ~x477 & ~x481 & ~x612 & ~x672 & ~x724 & ~x729 & ~x758;
assign c8448 =  x523 &  x547 &  x569 & ~x126 & ~x160 & ~x190 & ~x448;
assign c8450 =  x447;
assign c8452 =  x314 &  x327 & ~x2 & ~x20 & ~x28 & ~x32 & ~x36 & ~x42 & ~x50 & ~x60 & ~x702 & ~x732 & ~x761;
assign c8454 =  x292 & ~x399 & ~x623 & ~x654 & ~x684;
assign c8456 = ~x625 & ~x653;
assign c8458 = ~x554 & ~x627 & ~x697 & ~x721 & ~x737;
assign c8460 =  x339 &  x592 & ~x36 & ~x78;
assign c8462 =  x14 & ~x51 & ~x70 & ~x77 & ~x168 & ~x198 & ~x282;
assign c8464 = ~x10 & ~x17 & ~x18 & ~x77 & ~x79 & ~x89 & ~x104 & ~x106 & ~x116 & ~x132 & ~x133 & ~x246 & ~x272 & ~x274 & ~x293 & ~x301 & ~x321 & ~x325 & ~x330 & ~x343;
assign c8466 =  x487 &  x523 &  x546 & ~x2 & ~x59 & ~x78 & ~x80 & ~x138 & ~x274 & ~x276 & ~x592 & ~x777 & ~x783;
assign c8468 = ~x9 & ~x10 & ~x12 & ~x16 & ~x32 & ~x39 & ~x45 & ~x93 & ~x94 & ~x102 & ~x161 & ~x162 & ~x176 & ~x200 & ~x755;
assign c8470 = ~x12 & ~x20 & ~x73 & ~x107 & ~x130 & ~x176 & ~x187 & ~x199 & ~x215 & ~x230 & ~x231 & ~x232 & ~x233 & ~x243 & ~x247 & ~x259 & ~x260 & ~x273 & ~x287 & ~x300 & ~x329 & ~x331 & ~x583;
assign c8472 =  x348 & ~x10 & ~x88 & ~x422 & ~x567 & ~x569 & ~x596 & ~x627;
assign c8474 =  x222 &  x389 & ~x71 & ~x105;
assign c8476 =  x686 &  x692 & ~x65 & ~x227 & ~x771;
assign c8478 =  x560;
assign c8480 =  x693 &  x763 & ~x31;
assign c8482 = ~x77 & ~x106 & ~x442 & ~x456 & ~x485 & ~x486 & ~x514;
assign c8484 = ~x246 & ~x293 & ~x299 & ~x301 & ~x343 & ~x455;
assign c8486 =  x660 &  x744 & ~x11 & ~x38 & ~x65 & ~x131 & ~x216;
assign c8488 =  x664 &  x675 & ~x772;
assign c8490 =  x460 &  x469 &  x522 &  x549 &  x551 &  x580 &  x581 &  x659 &  x680 &  x693 & ~x115 & ~x167 & ~x170 & ~x336 & ~x529 & ~x589 & ~x700 & ~x758 & ~x778;
assign c8492 =  x14 & ~x69;
assign c8494 =  x682 & ~x57 & ~x61 & ~x98 & ~x117 & ~x182 & ~x306 & ~x781;
assign c8496 =  x401 &  x428 &  x542 &  x551 &  x553 &  x554 &  x598 &  x637 &  x712 &  x734 &  x737 &  x738 &  x740 & ~x56 & ~x141 & ~x142 & ~x167 & ~x336 & ~x530 & ~x780;
assign c8498 =  x561 & ~x217;
assign c81 =  x119 & ~x3 & ~x33 & ~x50 & ~x59 & ~x79 & ~x84 & ~x107 & ~x109 & ~x111 & ~x115 & ~x136 & ~x137 & ~x143 & ~x191 & ~x193 & ~x198 & ~x220 & ~x222 & ~x226 & ~x249 & ~x250 & ~x277 & ~x306 & ~x309 & ~x477 & ~x531 & ~x533 & ~x558 & ~x643 & ~x755;
assign c83 =  x747 & ~x2 & ~x4 & ~x5 & ~x22 & ~x23 & ~x24 & ~x25 & ~x26 & ~x28 & ~x29 & ~x30 & ~x31 & ~x32 & ~x51 & ~x53 & ~x54 & ~x56 & ~x57 & ~x58 & ~x81 & ~x82 & ~x84 & ~x85 & ~x87 & ~x109 & ~x110 & ~x111 & ~x113 & ~x114 & ~x137 & ~x138 & ~x141 & ~x166 & ~x167 & ~x169 & ~x195 & ~x196 & ~x222 & ~x223 & ~x224 & ~x252 & ~x279 & ~x307 & ~x308 & ~x362 & ~x363 & ~x364 & ~x391 & ~x392 & ~x419 & ~x447 & ~x453 & ~x475 & ~x497 & ~x503 & ~x555 & ~x559 & ~x561 & ~x562 & ~x563 & ~x564 & ~x565 & ~x584 & ~x585 & ~x586 & ~x587 & ~x590 & ~x591 & ~x592 & ~x611 & ~x613 & ~x614 & ~x618 & ~x620 & ~x638 & ~x639 & ~x640 & ~x641 & ~x642 & ~x643 & ~x644 & ~x645 & ~x646 & ~x647 & ~x648 & ~x649 & ~x667 & ~x668 & ~x669 & ~x670 & ~x671 & ~x672 & ~x673 & ~x674 & ~x675 & ~x676 & ~x695 & ~x696 & ~x697 & ~x698 & ~x699 & ~x700 & ~x701 & ~x702 & ~x703 & ~x704 & ~x705 & ~x724 & ~x725 & ~x726 & ~x727 & ~x729 & ~x731 & ~x732 & ~x733 & ~x752 & ~x753 & ~x755 & ~x756 & ~x757 & ~x758 & ~x759 & ~x760 & ~x761 & ~x779 & ~x780 & ~x781 & ~x783;
assign c85 =  x62 & ~x50 & ~x51 & ~x53 & ~x251 & ~x446 & ~x504 & ~x614;
assign c87 = ~x81 & ~x83 & ~x147 & ~x243 & ~x271 & ~x677;
assign c89 =  x163 &  x416 &  x529 & ~x223 & ~x280;
assign c811 = ~x208 & ~x282 & ~x312 & ~x630 & ~x674;
assign c813 =  x294 & ~x68 & ~x72 & ~x173 & ~x282 & ~x286 & ~x310 & ~x312;
assign c815 =  x77 &  x135 &  x192 &  x200 & ~x29;
assign c817 =  x120 &  x173 &  x213 &  x228 &  x275 & ~x52 & ~x81 & ~x108 & ~x166 & ~x194 & ~x559;
assign c819 =  x315 &  x594 & ~x1 & ~x28 & ~x50 & ~x115 & ~x138 & ~x143 & ~x194 & ~x224 & ~x249 & ~x277 & ~x389 & ~x392 & ~x446 & ~x478 & ~x502 & ~x505 & ~x533 & ~x587 & ~x764;
assign c821 =  x201 &  x339 &  x367 &  x368 & ~x80 & ~x197 & ~x222 & ~x335;
assign c823 = ~x167 & ~x310 & ~x314 & ~x363 & ~x390 & ~x620 & ~x649 & ~x667 & ~x770;
assign c825 =  x481 &  x509 & ~x33 & ~x111 & ~x165 & ~x171 & ~x248 & ~x389 & ~x725 & ~x726 & ~x764;
assign c827 = ~x6 & ~x20 & ~x22 & ~x28 & ~x52 & ~x57 & ~x82 & ~x95 & ~x99 & ~x100 & ~x101 & ~x109 & ~x137 & ~x139 & ~x195 & ~x250 & ~x281 & ~x334 & ~x364 & ~x419 & ~x475 & ~x510 & ~x532 & ~x560 & ~x757 & ~x758 & ~x760 & ~x761 & ~x762;
assign c829 =  x360 &  x585 & ~x289;
assign c831 =  x44 &  x510 & ~x0 & ~x1 & ~x23 & ~x26 & ~x27 & ~x28 & ~x29 & ~x31 & ~x48 & ~x51 & ~x58 & ~x60 & ~x86 & ~x87 & ~x88 & ~x112 & ~x136 & ~x138 & ~x192 & ~x195 & ~x196 & ~x251 & ~x253 & ~x282 & ~x305 & ~x306 & ~x307 & ~x333 & ~x334 & ~x362 & ~x363 & ~x365 & ~x367 & ~x394 & ~x417 & ~x445 & ~x450 & ~x477 & ~x504 & ~x532 & ~x560 & ~x561 & ~x646 & ~x669 & ~x670 & ~x697 & ~x701 & ~x725 & ~x727 & ~x755 & ~x781;
assign c833 = ~x14 & ~x121 & ~x312 & ~x314 & ~x717;
assign c835 = ~x86 & ~x198 & ~x310 & ~x338 & ~x340 & ~x423 & ~x449 & ~x505 & ~x517 & ~x729;
assign c837 =  x442 & ~x14 & ~x198 & ~x227 & ~x281 & ~x310 & ~x337 & ~x746;
assign c839 =  x218 & ~x260 & ~x281;
assign c841 =  x178 &  x265 &  x347 &  x349 &  x377 &  x431 &  x660 & ~x34 & ~x57 & ~x111 & ~x133 & ~x161 & ~x251 & ~x640;
assign c843 = ~x14 & ~x96 & ~x125 & ~x143 & ~x340 & ~x341 & ~x367 & ~x420 & ~x454 & ~x506;
assign c845 =  x538 & ~x4 & ~x19 & ~x25 & ~x51 & ~x86 & ~x137 & ~x143 & ~x227 & ~x363 & ~x419 & ~x475 & ~x589 & ~x735;
assign c847 =  x184 &  x187 &  x536 & ~x51 & ~x255 & ~x276 & ~x333 & ~x391;
assign c849 = ~x8 & ~x31 & ~x52 & ~x222 & ~x280 & ~x306 & ~x336 & ~x337 & ~x339 & ~x399 & ~x412 & ~x413 & ~x448 & ~x455 & ~x511 & ~x525 & ~x528 & ~x529 & ~x537 & ~x538 & ~x555 & ~x559 & ~x566 & ~x590 & ~x593 & ~x615 & ~x617 & ~x622 & ~x645 & ~x646 & ~x667 & ~x672 & ~x675 & ~x676 & ~x695 & ~x696 & ~x705 & ~x726 & ~x760 & ~x778;
assign c851 =  x454 & ~x630;
assign c853 = ~x72 & ~x289 & ~x314 & ~x315 & ~x340 & ~x365 & ~x717;
assign c855 =  x590 &  x618 &  x641;
assign c857 =  x407 &  x486 &  x493 &  x570 &  x598 & ~x25 & ~x29 & ~x30 & ~x57 & ~x58 & ~x81 & ~x82 & ~x279 & ~x363 & ~x441 & ~x502 & ~x526 & ~x557 & ~x561 & ~x588 & ~x592 & ~x593 & ~x616 & ~x669 & ~x781;
assign c859 = ~x166 & ~x186 & ~x241 & ~x534 & ~x577 & ~x669 & ~x764;
assign c861 =  x36 &  x256 &  x550 & ~x23 & ~x51 & ~x54 & ~x109 & ~x197 & ~x334 & ~x335 & ~x363;
assign c863 =  x426 &  x482 & ~x225 & ~x227 & ~x255 & ~x283 & ~x589 & ~x618 & ~x767 & ~x771;
assign c865 =  x622 & ~x370 & ~x426;
assign c867 =  x12 &  x41 &  x42 & ~x0 & ~x6 & ~x34 & ~x51 & ~x57 & ~x79 & ~x110 & ~x114 & ~x116 & ~x166 & ~x223 & ~x224 & ~x277 & ~x311 & ~x419 & ~x421 & ~x422 & ~x474 & ~x478 & ~x501 & ~x505 & ~x530 & ~x558 & ~x559 & ~x617 & ~x643 & ~x763;
assign c869 =  x409 & ~x40 & ~x41 & ~x174 & ~x191 & ~x275;
assign c871 =  x498 & ~x224 & ~x276 & ~x308 & ~x336 & ~x393 & ~x748 & ~x756 & ~x763;
assign c873 =  x47 &  x118 & ~x5 & ~x24 & ~x31 & ~x51 & ~x54 & ~x59 & ~x84 & ~x86 & ~x109 & ~x166 & ~x224 & ~x226 & ~x250 & ~x279 & ~x280 & ~x334 & ~x337 & ~x364 & ~x391 & ~x392 & ~x475 & ~x476 & ~x477 & ~x531 & ~x560 & ~x588 & ~x616 & ~x755 & ~x781;
assign c875 =  x220 &  x540 & ~x555;
assign c877 =  x117 & ~x505 & ~x533 & ~x584 & ~x586 & ~x587 & ~x592 & ~x611 & ~x615 & ~x620 & ~x643 & ~x755;
assign c879 = ~x236 & ~x310 & ~x340 & ~x367 & ~x766;
assign c881 =  x304 &  x332 &  x389 &  x596 & ~x14 & ~x25 & ~x337;
assign c883 =  x40 &  x41 &  x42 &  x43 &  x358 & ~x29 & ~x33 & ~x34 & ~x52 & ~x79 & ~x83 & ~x84 & ~x108 & ~x109 & ~x110 & ~x137 & ~x142 & ~x169 & ~x193 & ~x252 & ~x253 & ~x278 & ~x281 & ~x306 & ~x362 & ~x363 & ~x364 & ~x390 & ~x391 & ~x394 & ~x418 & ~x421 & ~x422 & ~x446 & ~x448 & ~x449 & ~x477 & ~x505 & ~x559 & ~x561 & ~x588 & ~x589 & ~x617 & ~x758;
assign c885 =  x300 & ~x289 & ~x310 & ~x337 & ~x776;
assign c887 =  x187 &  x316 &  x467 &  x706 & ~x82 & ~x83 & ~x168 & ~x363 & ~x448 & ~x507 & ~x529 & ~x534 & ~x556 & ~x560 & ~x562 & ~x584 & ~x590 & ~x619 & ~x671 & ~x672 & ~x674 & ~x675 & ~x703 & ~x727 & ~x754;
assign c889 =  x171 &  x255 & ~x166;
assign c891 =  x570 &  x597 &  x598 &  x634 & ~x3 & ~x4 & ~x24 & ~x25 & ~x26 & ~x27 & ~x28 & ~x29 & ~x30 & ~x51 & ~x52 & ~x54 & ~x55 & ~x82 & ~x83 & ~x86 & ~x112 & ~x140 & ~x142 & ~x166 & ~x168 & ~x169 & ~x194 & ~x195 & ~x196 & ~x197 & ~x222 & ~x252 & ~x391 & ~x475 & ~x504 & ~x537 & ~x582 & ~x592 & ~x593 & ~x610 & ~x611 & ~x615 & ~x617 & ~x620 & ~x621 & ~x639 & ~x649 & ~x667 & ~x668 & ~x670 & ~x677 & ~x695 & ~x696 & ~x704 & ~x705 & ~x733 & ~x752 & ~x757 & ~x761 & ~x781;
assign c893 =  x185 &  x330 &  x500 &  x508 &  x535 & ~x193;
assign c895 =  x174 &  x208 &  x387 &  x536 &  x556 &  x606 & ~x53 & ~x81 & ~x109 & ~x142 & ~x166 & ~x169 & ~x198 & ~x226 & ~x254 & ~x334;
assign c897 =  x442 & ~x1 & ~x141 & ~x252 & ~x262 & ~x281 & ~x309 & ~x336 & ~x339 & ~x744 & ~x770;
assign c899 = ~x1 & ~x8 & ~x32 & ~x56 & ~x75 & ~x79 & ~x80 & ~x136 & ~x138 & ~x143 & ~x223 & ~x226 & ~x277 & ~x279 & ~x307 & ~x309 & ~x334 & ~x389 & ~x391 & ~x422 & ~x446 & ~x450 & ~x478 & ~x502 & ~x505 & ~x558 & ~x562 & ~x586 & ~x614 & ~x615 & ~x617 & ~x645 & ~x672 & ~x673 & ~x701 & ~x735 & ~x763 & ~x773 & ~x781 & ~x783;
assign c8101 =  x748 & ~x57 & ~x497 & ~x621;
assign c8103 =  x426 &  x481 & ~x169 & ~x200 & ~x227 & ~x253 & ~x255 & ~x256 & ~x668 & ~x671;
assign c8105 =  x320 &  x515 &  x516 & ~x72 & ~x561 & ~x593;
assign c8107 = ~x2 & ~x5 & ~x141 & ~x143 & ~x163 & ~x194 & ~x197 & ~x225 & ~x236 & ~x253 & ~x278 & ~x306 & ~x334 & ~x365 & ~x505 & ~x511 & ~x533 & ~x617 & ~x699 & ~x728 & ~x759 & ~x761 & ~x762;
assign c8109 =  x632 & ~x13 & ~x22 & ~x25 & ~x29 & ~x32 & ~x41 & ~x51 & ~x55 & ~x84 & ~x138 & ~x167 & ~x168 & ~x195 & ~x279 & ~x363 & ~x419 & ~x447 & ~x476 & ~x531 & ~x559 & ~x589 & ~x644 & ~x647 & ~x667 & ~x669 & ~x675 & ~x727 & ~x728 & ~x729 & ~x731 & ~x757 & ~x782;
assign c8111 =  x129 &  x259 &  x470 & ~x116 & ~x135 & ~x139 & ~x191 & ~x276 & ~x305;
assign c8113 =  x160 &  x388 & ~x79;
assign c8115 =  x739 & ~x6 & ~x14 & ~x251 & ~x469 & ~x554 & ~x555 & ~x621 & ~x667;
assign c8117 =  x750 & ~x505 & ~x748;
assign c8119 =  x751 & ~x736;
assign c8121 =  x207 & ~x79 & ~x189 & ~x313 & ~x330 & ~x342 & ~x366 & ~x388 & ~x529 & ~x557 & ~x583 & ~x783;
assign c8123 =  x287 &  x694 & ~x110 & ~x112 & ~x141 & ~x196 & ~x276 & ~x277 & ~x283 & ~x305 & ~x307 & ~x336 & ~x450 & ~x501 & ~x505 & ~x534 & ~x559 & ~x562 & ~x701 & ~x702 & ~x727 & ~x754;
assign c8125 =  x349 &  x375 & ~x84 & ~x280 & ~x298 & ~x727;
assign c8127 =  x488 &  x630 &  x655 & ~x3 & ~x13 & ~x28 & ~x39 & ~x42 & ~x43 & ~x57 & ~x109 & ~x114 & ~x139 & ~x140 & ~x250 & ~x251 & ~x335 & ~x363 & ~x587 & ~x668 & ~x760;
assign c8129 =  x105 &  x737 & ~x0 & ~x3 & ~x4 & ~x14 & ~x24 & ~x166;
assign c8131 =  x204 &  x317 &  x481 &  x509 &  x604 &  x662 & ~x59 & ~x82 & ~x87 & ~x137 & ~x140 & ~x170 & ~x198 & ~x224 & ~x226 & ~x248 & ~x249 & ~x250 & ~x277 & ~x307 & ~x309 & ~x334 & ~x335 & ~x362 & ~x475 & ~x674 & ~x697 & ~x701 & ~x755;
assign c8133 =  x456 & ~x223 & ~x257 & ~x282 & ~x634 & ~x650;
assign c8135 =  x69 &  x442 &  x537 &  x681 & ~x5 & ~x50 & ~x81 & ~x361 & ~x418 & ~x449;
assign c8137 =  x425 & ~x579;
assign c8139 =  x443 & ~x229 & ~x232 & ~x288 & ~x309 & ~x314 & ~x339;
assign c8141 =  x200 & ~x592 & ~x593 & ~x611 & ~x620 & ~x641 & ~x648 & ~x675 & ~x695 & ~x697 & ~x704 & ~x757 & ~x783;
assign c8143 =  x571 & ~x5 & ~x23 & ~x32 & ~x56 & ~x110 & ~x141 & ~x250 & ~x276 & ~x280 & ~x281 & ~x305 & ~x309 & ~x364 & ~x391 & ~x476 & ~x507 & ~x529 & ~x530 & ~x532 & ~x535 & ~x557 & ~x558 & ~x585 & ~x590 & ~x591 & ~x613 & ~x614 & ~x647 & ~x670 & ~x675 & ~x759 & ~x764 & ~x773 & ~x783;
assign c8145 = ~x334 & ~x548 & ~x561 & ~x591;
assign c8147 = ~x57 & ~x90 & ~x143 & ~x202 & ~x234 & ~x288 & ~x310 & ~x317 & ~x344 & ~x368 & ~x393 & ~x395 & ~x419 & ~x422;
assign c8149 =  x399 & ~x262 & ~x661;
assign c8151 =  x535 &  x536 &  x556 & ~x253 & ~x762 & ~x763;
assign c8153 =  x515 &  x655 & ~x496 & ~x696 & ~x731;
assign c8155 = ~x170 & ~x202 & ~x261 & ~x292 & ~x309 & ~x367 & ~x368 & ~x369 & ~x422;
assign c8157 =  x481 & ~x313;
assign c8159 =  x160 &  x444 &  x619;
assign c8161 =  x655 &  x656 & ~x0 & ~x1 & ~x2 & ~x13 & ~x24 & ~x28 & ~x29 & ~x32 & ~x57 & ~x68 & ~x83 & ~x85 & ~x111 & ~x224 & ~x337 & ~x365 & ~x366 & ~x368 & ~x369 & ~x394 & ~x395 & ~x397 & ~x421 & ~x449 & ~x450 & ~x451 & ~x478 & ~x671 & ~x699 & ~x730;
assign c8163 = ~x362 & ~x374 & ~x402 & ~x486;
assign c8165 = ~x171 & ~x283 & ~x287 & ~x310 & ~x770;
assign c8167 =  x129 &  x479 &  x480 &  x585 & ~x137;
assign c8169 = ~x115 & ~x205 & ~x255 & ~x262 & ~x263 & ~x282 & ~x337 & ~x365;
assign c8171 =  x564 & ~x193 & ~x222 & ~x225 & ~x254 & ~x278 & ~x280 & ~x447 & ~x474 & ~x671 & ~x764 & ~x766;
assign c8173 = ~x402 & ~x502 & ~x538;
assign c8175 =  x360 & ~x315 & ~x340;
assign c8177 = ~x150 & ~x234 & ~x254 & ~x282 & ~x283 & ~x289 & ~x314 & ~x336 & ~x337 & ~x745 & ~x746;
assign c8179 = ~x142 & ~x340 & ~x393 & ~x439 & ~x473 & ~x589 & ~x608;
assign c8181 =  x39 &  x42 &  x43 & ~x7 & ~x48 & ~x49 & ~x51 & ~x79 & ~x115 & ~x196 & ~x281 & ~x306 & ~x365 & ~x389 & ~x390 & ~x445 & ~x450 & ~x533 & ~x614 & ~x643 & ~x669 & ~x783;
assign c8183 =  x232 &  x243 &  x266 &  x288 &  x470 &  x493 & ~x135 & ~x143 & ~x163 & ~x192 & ~x198 & ~x252 & ~x276 & ~x337 & ~x420;
assign c8185 =  x452 &  x454 & ~x309 & ~x595;
assign c8187 =  x93 &  x94 &  x201 &  x368 & ~x61 & ~x136 & ~x477;
assign c8189 = ~x14 & ~x42 & ~x255 & ~x258 & ~x282 & ~x340 & ~x367 & ~x420 & ~x729 & ~x756;
assign c8191 =  x102 &  x129 &  x228 &  x284 &  x292 &  x549 & ~x137 & ~x252;
assign c8193 =  x736 & ~x25 & ~x28 & ~x55 & ~x59 & ~x87 & ~x138 & ~x309 & ~x340 & ~x369 & ~x452 & ~x454 & ~x474 & ~x476 & ~x480 & ~x530 & ~x535 & ~x560 & ~x587 & ~x671 & ~x756 & ~x758 & ~x783;
assign c8195 =  x463 &  x661 & ~x13 & ~x14 & ~x564 & ~x584 & ~x590 & ~x641;
assign c8197 =  x15 &  x40 &  x42 & ~x51 & ~x58 & ~x108 & ~x140 & ~x170 & ~x335 & ~x365 & ~x448 & ~x587 & ~x616;
assign c8199 =  x174 &  x201 &  x228 &  x247 &  x303 &  x456 &  x569 &  x663 & ~x137;
assign c8201 =  x214 &  x244 &  x272 &  x436 &  x568 &  x601 &  x653;
assign c8203 =  x214 &  x266 &  x576 &  x579 & ~x33 & ~x50 & ~x51 & ~x57 & ~x78 & ~x79 & ~x80 & ~x90 & ~x107 & ~x135 & ~x140 & ~x168 & ~x192 & ~x194 & ~x196 & ~x248 & ~x391 & ~x392 & ~x394 & ~x445 & ~x447 & ~x448 & ~x449 & ~x473 & ~x474 & ~x477 & ~x502 & ~x504 & ~x587 & ~x669 & ~x730 & ~x734 & ~x758 & ~x781;
assign c8205 = ~x206 & ~x235 & ~x285 & ~x340;
assign c8207 =  x130 &  x724;
assign c8209 = ~x0 & ~x3 & ~x5 & ~x23 & ~x25 & ~x28 & ~x32 & ~x35 & ~x49 & ~x53 & ~x55 & ~x56 & ~x58 & ~x59 & ~x61 & ~x78 & ~x79 & ~x82 & ~x83 & ~x87 & ~x113 & ~x138 & ~x139 & ~x166 & ~x169 & ~x252 & ~x279 & ~x335 & ~x477 & ~x478 & ~x479 & ~x502 & ~x527 & ~x528 & ~x529 & ~x535 & ~x557 & ~x558 & ~x559 & ~x561 & ~x562 & ~x563 & ~x587 & ~x589 & ~x590 & ~x591 & ~x613 & ~x617 & ~x618 & ~x619 & ~x642 & ~x644 & ~x646 & ~x647 & ~x669 & ~x674 & ~x675 & ~x698 & ~x699 & ~x701 & ~x702 & ~x703 & ~x725 & ~x726 & ~x730 & ~x754 & ~x756 & ~x757 & ~x763 & ~x765 & ~x766 & ~x773 & ~x776;
assign c8211 =  x259 &  x442 & ~x5 & ~x167 & ~x198 & ~x220 & ~x222 & ~x227 & ~x249 & ~x276 & ~x277 & ~x280 & ~x305 & ~x306 & ~x307 & ~x333 & ~x335 & ~x337 & ~x447 & ~x731 & ~x764;
assign c8213 =  x345 & ~x30 & ~x151 & ~x166 & ~x536 & ~x649;
assign c8215 =  x175 &  x526 & ~x145 & ~x163 & ~x198 & ~x220 & ~x255 & ~x361;
assign c8217 = ~x55 & ~x72 & ~x338 & ~x344 & ~x771;
assign c8219 =  x65 &  x91 &  x120 & ~x108 & ~x250 & ~x252 & ~x531;
assign c8221 =  x471 & ~x289 & ~x311;
assign c8223 = ~x1 & ~x28 & ~x55 & ~x164 & ~x278 & ~x339 & ~x551 & ~x617 & ~x641 & ~x726 & ~x729 & ~x736;
assign c8225 =  x454 & ~x227 & ~x773;
assign c8227 =  x248 &  x625 & ~x14 & ~x476;
assign c8229 = ~x179 & ~x208 & ~x228 & ~x335 & ~x340 & ~x687 & ~x755 & ~x773;
assign c8231 = ~x0 & ~x2 & ~x5 & ~x6 & ~x21 & ~x22 & ~x24 & ~x27 & ~x52 & ~x53 & ~x54 & ~x56 & ~x57 & ~x59 & ~x81 & ~x82 & ~x83 & ~x84 & ~x86 & ~x109 & ~x112 & ~x114 & ~x139 & ~x141 & ~x142 & ~x163 & ~x165 & ~x166 & ~x194 & ~x196 & ~x197 & ~x198 & ~x202 & ~x222 & ~x223 & ~x224 & ~x225 & ~x228 & ~x247 & ~x251 & ~x258 & ~x279 & ~x286 & ~x301 & ~x314 & ~x329 & ~x332 & ~x333 & ~x337 & ~x338 & ~x342 & ~x357 & ~x362 & ~x363 & ~x364 & ~x365 & ~x366 & ~x367 & ~x369 & ~x386 & ~x393 & ~x394 & ~x395 & ~x398 & ~x413 & ~x414 & ~x416 & ~x417 & ~x418 & ~x419 & ~x420 & ~x421 & ~x422 & ~x423 & ~x424 & ~x425 & ~x441 & ~x443 & ~x444 & ~x447 & ~x451 & ~x452 & ~x454 & ~x470 & ~x471 & ~x472 & ~x474 & ~x475 & ~x480 & ~x498 & ~x499 & ~x500 & ~x501 & ~x502 & ~x503 & ~x505 & ~x506 & ~x507 & ~x508 & ~x509 & ~x510 & ~x526 & ~x527 & ~x529 & ~x530 & ~x535 & ~x538 & ~x555 & ~x558 & ~x561 & ~x562 & ~x563 & ~x582 & ~x583 & ~x585 & ~x587 & ~x588 & ~x591 & ~x592 & ~x611 & ~x613 & ~x614 & ~x616 & ~x618 & ~x619 & ~x621 & ~x638 & ~x641 & ~x646 & ~x647 & ~x648 & ~x667 & ~x670 & ~x672 & ~x673 & ~x675 & ~x676 & ~x696 & ~x697 & ~x698 & ~x700 & ~x702 & ~x704 & ~x705 & ~x724 & ~x725 & ~x728 & ~x730 & ~x732 & ~x751 & ~x753 & ~x755 & ~x757 & ~x758 & ~x759 & ~x782;
assign c8233 = ~x0 & ~x1 & ~x2 & ~x17 & ~x21 & ~x25 & ~x26 & ~x27 & ~x32 & ~x33 & ~x35 & ~x48 & ~x50 & ~x51 & ~x53 & ~x59 & ~x60 & ~x61 & ~x63 & ~x76 & ~x78 & ~x79 & ~x85 & ~x88 & ~x107 & ~x112 & ~x113 & ~x114 & ~x116 & ~x135 & ~x137 & ~x139 & ~x141 & ~x143 & ~x166 & ~x171 & ~x192 & ~x194 & ~x195 & ~x196 & ~x223 & ~x225 & ~x227 & ~x249 & ~x251 & ~x253 & ~x275 & ~x278 & ~x279 & ~x280 & ~x305 & ~x306 & ~x308 & ~x310 & ~x334 & ~x338 & ~x362 & ~x363 & ~x365 & ~x366 & ~x367 & ~x389 & ~x392 & ~x395 & ~x417 & ~x445 & ~x446 & ~x475 & ~x476 & ~x503 & ~x505 & ~x506 & ~x530 & ~x531 & ~x533 & ~x534 & ~x560 & ~x585 & ~x588 & ~x617 & ~x645 & ~x646 & ~x669 & ~x671 & ~x673 & ~x692 & ~x698 & ~x700 & ~x703 & ~x725 & ~x728 & ~x753 & ~x759 & ~x776 & ~x781 & ~x783;
assign c8235 =  x333 & ~x119 & ~x255 & ~x316 & ~x364;
assign c8237 = ~x15 & ~x43 & ~x121 & ~x229 & ~x254 & ~x261 & ~x311 & ~x369 & ~x372 & ~x425;
assign c8239 =  x426 & ~x117 & ~x589 & ~x679 & ~x703;
assign c8241 =  x42 &  x43 & ~x28 & ~x38 & ~x52 & ~x110 & ~x142 & ~x167 & ~x169 & ~x223 & ~x309 & ~x419 & ~x502 & ~x507 & ~x529 & ~x558 & ~x587 & ~x591 & ~x619 & ~x620 & ~x640 & ~x643 & ~x648 & ~x671 & ~x731 & ~x757 & ~x779;
assign c8243 =  x44 &  x71 & ~x75 & ~x532 & ~x533;
assign c8245 = ~x355;
assign c8247 =  x486 & ~x399 & ~x452 & ~x468 & ~x479;
assign c8249 =  x66 &  x485 &  x513 &  x541 & ~x0 & ~x1 & ~x56 & ~x169 & ~x197 & ~x363 & ~x482 & ~x640 & ~x667 & ~x668;
assign c8251 =  x243 &  x267 &  x271 &  x288 &  x325 &  x347 &  x466 &  x488 &  x491 &  x600 &  x651 & ~x0 & ~x22 & ~x25 & ~x26 & ~x28 & ~x111 & ~x139 & ~x140 & ~x336 & ~x391 & ~x395 & ~x419 & ~x421 & ~x424 & ~x444 & ~x447 & ~x448 & ~x449 & ~x450 & ~x472 & ~x474 & ~x475 & ~x477 & ~x479 & ~x480 & ~x500 & ~x501 & ~x502 & ~x503 & ~x504 & ~x507 & ~x528 & ~x529 & ~x535 & ~x560 & ~x562 & ~x563 & ~x584 & ~x586 & ~x591 & ~x592 & ~x613 & ~x614 & ~x615 & ~x617 & ~x618 & ~x640 & ~x641 & ~x642 & ~x644 & ~x645 & ~x646 & ~x647 & ~x668 & ~x669 & ~x671 & ~x674 & ~x675 & ~x697 & ~x698 & ~x702 & ~x703 & ~x724 & ~x725 & ~x730 & ~x731 & ~x752 & ~x756 & ~x760 & ~x781 & ~x782;
assign c8253 =  x46 &  x736 &  x772 & ~x33 & ~x51 & ~x475;
assign c8255 = ~x310 & ~x372 & ~x400;
assign c8257 = ~x122 & ~x367 & ~x490 & ~x577;
assign c8259 =  x187 &  x414 &  x526 &  x579 &  x635 &  x653 &  x660 & ~x50 & ~x80 & ~x192 & ~x226 & ~x249 & ~x310 & ~x333 & ~x334 & ~x389 & ~x393 & ~x503;
assign c8261 = ~x96 & ~x113 & ~x151 & ~x236 & ~x310 & ~x659;
assign c8263 =  x126 & ~x34 & ~x54 & ~x121 & ~x140 & ~x141 & ~x170 & ~x198 & ~x279 & ~x308 & ~x309 & ~x394 & ~x448 & ~x452 & ~x559;
assign c8265 =  x397 & ~x250 & ~x590;
assign c8267 =  x434 &  x582 & ~x50 & ~x144 & ~x191 & ~x198 & ~x219 & ~x227 & ~x247 & ~x248 & ~x276 & ~x280 & ~x389 & ~x418 & ~x419 & ~x503 & ~x531 & ~x669 & ~x698 & ~x699 & ~x702 & ~x726 & ~x730 & ~x781;
assign c8269 = ~x142 & ~x144 & ~x145 & ~x151 & ~x152 & ~x253 & ~x256 & ~x532 & ~x563 & ~x675 & ~x724 & ~x777 & ~x780;
assign c8271 =  x40 &  x41 &  x42 &  x43 & ~x8 & ~x19 & ~x23 & ~x31 & ~x33 & ~x35 & ~x48 & ~x53 & ~x55 & ~x80 & ~x81 & ~x87 & ~x107 & ~x111 & ~x139 & ~x194 & ~x199 & ~x222 & ~x224 & ~x254 & ~x333 & ~x336 & ~x365 & ~x366 & ~x389 & ~x448 & ~x477 & ~x503 & ~x505 & ~x615 & ~x617 & ~x645 & ~x672 & ~x674 & ~x727 & ~x730 & ~x753 & ~x755 & ~x759 & ~x781;
assign c8273 =  x641 &  x703 &  x725;
assign c8275 = ~x59 & ~x143 & ~x166 & ~x168 & ~x170 & ~x226 & ~x253 & ~x306 & ~x384 & ~x392 & ~x419 & ~x477 & ~x504 & ~x526 & ~x527 & ~x530 & ~x537 & ~x555 & ~x561 & ~x564 & ~x583 & ~x584 & ~x610 & ~x617 & ~x622 & ~x666 & ~x697 & ~x704 & ~x734 & ~x777 & ~x779 & ~x781;
assign c8277 =  x538 &  x733 & ~x34 & ~x365 & ~x389 & ~x502 & ~x562 & ~x674 & ~x764;
assign c8279 =  x12 &  x42 & ~x50 & ~x166 & ~x420 & ~x588;
assign c8281 =  x9;
assign c8283 =  x485 &  x603 &  x694 & ~x28 & ~x31 & ~x50 & ~x51 & ~x52 & ~x53 & ~x85 & ~x107 & ~x109 & ~x111 & ~x113 & ~x164 & ~x195 & ~x197 & ~x219 & ~x248 & ~x250 & ~x276 & ~x279 & ~x304 & ~x305 & ~x362 & ~x367 & ~x392 & ~x420 & ~x451 & ~x475 & ~x477 & ~x478 & ~x529 & ~x534 & ~x669 & ~x702 & ~x726 & ~x753 & ~x754 & ~x755 & ~x757;
assign c8285 = ~x311 & ~x340 & ~x411 & ~x530;
assign c8287 = ~x2 & ~x6 & ~x13 & ~x14 & ~x42 & ~x55 & ~x57 & ~x170 & ~x173 & ~x194 & ~x251 & ~x253 & ~x285 & ~x309 & ~x338 & ~x341 & ~x368 & ~x370 & ~x392 & ~x399 & ~x424 & ~x427 & ~x533;
assign c8289 =  x41 &  x42 &  x43 &  x70 & ~x0 & ~x4 & ~x56 & ~x59 & ~x64 & ~x168 & ~x223 & ~x253 & ~x308 & ~x333 & ~x420 & ~x421 & ~x448 & ~x449 & ~x450 & ~x475 & ~x478 & ~x729 & ~x756 & ~x782;
assign c8291 =  x508 &  x511 & ~x142 & ~x199 & ~x254 & ~x281 & ~x282 & ~x283 & ~x310 & ~x338 & ~x645 & ~x710 & ~x782;
assign c8293 = ~x28 & ~x31 & ~x55 & ~x141 & ~x147 & ~x168 & ~x259 & ~x287 & ~x329 & ~x340 & ~x369 & ~x371 & ~x394 & ~x397 & ~x422 & ~x425 & ~x426 & ~x450 & ~x452 & ~x453 & ~x477 & ~x478 & ~x480 & ~x481 & ~x499 & ~x500 & ~x502 & ~x506 & ~x507 & ~x509 & ~x510 & ~x527 & ~x533 & ~x535 & ~x556 & ~x562 & ~x563 & ~x565 & ~x582 & ~x610 & ~x640 & ~x760;
assign c8295 =  x315 &  x665 & ~x13 & ~x15 & ~x53 & ~x476 & ~x583 & ~x591 & ~x647 & ~x668 & ~x670 & ~x702;
assign c8297 = ~x20 & ~x55 & ~x59 & ~x63 & ~x138 & ~x169 & ~x170 & ~x197 & ~x227 & ~x252 & ~x332 & ~x335 & ~x360 & ~x366 & ~x390 & ~x394 & ~x395 & ~x445 & ~x446 & ~x473 & ~x474 & ~x479 & ~x535 & ~x559 & ~x585 & ~x613 & ~x614 & ~x616 & ~x617 & ~x664 & ~x669 & ~x670 & ~x673 & ~x692 & ~x702 & ~x730 & ~x755 & ~x759 & ~x763 & ~x775 & ~x776 & ~x777;
assign c8299 =  x593 & ~x24 & ~x30 & ~x50 & ~x57 & ~x79 & ~x169 & ~x365 & ~x395 & ~x422 & ~x616 & ~x701 & ~x765;
assign c8301 =  x40 &  x41 &  x43 & ~x26 & ~x36 & ~x37 & ~x48 & ~x58 & ~x61 & ~x78 & ~x79 & ~x111 & ~x196 & ~x221 & ~x362 & ~x365 & ~x391 & ~x420 & ~x560 & ~x755;
assign c8303 =  x173 &  x661 & ~x733;
assign c8305 =  x40 &  x69 & ~x64 & ~x77;
assign c8307 = ~x64 & ~x143 & ~x178 & ~x204 & ~x252 & ~x281 & ~x314 & ~x339 & ~x340 & ~x713 & ~x744 & ~x745;
assign c8309 = ~x269 & ~x278 & ~x563 & ~x625 & ~x706;
assign c8311 = ~x232 & ~x478 & ~x517;
assign c8313 =  x374 & ~x25 & ~x58 & ~x113 & ~x133 & ~x166 & ~x192 & ~x194 & ~x224 & ~x252 & ~x253 & ~x335 & ~x475 & ~x533 & ~x587 & ~x613 & ~x615 & ~x618 & ~x753 & ~x754 & ~x766;
assign c8315 =  x160 &  x585 & ~x365;
assign c8317 =  x70 &  x537 &  x564 & ~x50 & ~x277 & ~x305 & ~x337 & ~x361;
assign c8319 =  x266 &  x288 &  x656 & ~x2 & ~x26 & ~x53 & ~x83 & ~x85 & ~x110 & ~x139 & ~x307 & ~x421 & ~x445 & ~x448 & ~x451 & ~x452 & ~x471 & ~x473 & ~x479 & ~x500 & ~x528 & ~x529 & ~x533 & ~x556 & ~x558 & ~x559 & ~x562 & ~x563 & ~x585 & ~x586 & ~x589 & ~x591 & ~x642 & ~x644 & ~x668 & ~x669 & ~x674 & ~x675 & ~x698 & ~x699 & ~x724 & ~x725 & ~x726 & ~x728 & ~x755 & ~x759 & ~x779 & ~x780;
assign c8321 =  x44 &  x70 &  x469 &  x510 & ~x50 & ~x138 & ~x250 & ~x279 & ~x334 & ~x365 & ~x645;
assign c8323 =  x405 &  x627 &  x655 &  x683 &  x715 & ~x3 & ~x11 & ~x23 & ~x24 & ~x28 & ~x29 & ~x57 & ~x82 & ~x112 & ~x138 & ~x140 & ~x196 & ~x224 & ~x251 & ~x307 & ~x364 & ~x390 & ~x394 & ~x395 & ~x415 & ~x421 & ~x443 & ~x445 & ~x448 & ~x449 & ~x453 & ~x454 & ~x471 & ~x474 & ~x475 & ~x477 & ~x479 & ~x498 & ~x501 & ~x502 & ~x504 & ~x509 & ~x531 & ~x532 & ~x535 & ~x536 & ~x557 & ~x559 & ~x560 & ~x565 & ~x584 & ~x585 & ~x592 & ~x611 & ~x612 & ~x613 & ~x614 & ~x615 & ~x639 & ~x641 & ~x645 & ~x668 & ~x669 & ~x673 & ~x674 & ~x695 & ~x698 & ~x704 & ~x723 & ~x724 & ~x756 & ~x758 & ~x760 & ~x780;
assign c8325 = ~x255 & ~x309 & ~x338 & ~x392 & ~x633;
assign c8327 = ~x283 & ~x311 & ~x312;
assign c8329 =  x179 &  x264 & ~x161 & ~x174 & ~x223 & ~x475 & ~x508 & ~x536 & ~x555 & ~x583 & ~x584 & ~x619 & ~x675 & ~x754 & ~x782;
assign c8331 =  x324 &  x436 &  x492 &  x604 &  x626 & ~x11 & ~x31 & ~x57 & ~x58 & ~x83 & ~x86 & ~x114 & ~x117 & ~x145 & ~x164 & ~x192 & ~x195 & ~x220 & ~x223 & ~x249 & ~x250 & ~x252 & ~x255 & ~x276 & ~x278 & ~x279 & ~x304 & ~x309 & ~x339 & ~x389 & ~x451 & ~x477 & ~x588 & ~x590 & ~x614 & ~x617 & ~x618 & ~x642 & ~x646 & ~x669 & ~x673 & ~x701 & ~x725 & ~x726 & ~x755 & ~x756 & ~x764;
assign c8333 =  x17 &  x44 & ~x50;
assign c8335 =  x40 &  x41 &  x42 & ~x0 & ~x2 & ~x6 & ~x21 & ~x24 & ~x25 & ~x27 & ~x29 & ~x30 & ~x32 & ~x34 & ~x35 & ~x36 & ~x49 & ~x50 & ~x51 & ~x52 & ~x54 & ~x55 & ~x56 & ~x57 & ~x58 & ~x60 & ~x77 & ~x79 & ~x81 & ~x82 & ~x83 & ~x85 & ~x86 & ~x87 & ~x107 & ~x109 & ~x111 & ~x112 & ~x114 & ~x117 & ~x138 & ~x141 & ~x143 & ~x163 & ~x165 & ~x167 & ~x168 & ~x170 & ~x193 & ~x194 & ~x195 & ~x219 & ~x224 & ~x249 & ~x250 & ~x255 & ~x277 & ~x278 & ~x304 & ~x309 & ~x310 & ~x332 & ~x333 & ~x334 & ~x335 & ~x338 & ~x360 & ~x361 & ~x362 & ~x363 & ~x365 & ~x366 & ~x392 & ~x393 & ~x395 & ~x416 & ~x418 & ~x419 & ~x422 & ~x423 & ~x444 & ~x445 & ~x446 & ~x448 & ~x449 & ~x450 & ~x451 & ~x473 & ~x474 & ~x475 & ~x476 & ~x478 & ~x479 & ~x501 & ~x502 & ~x503 & ~x530 & ~x531 & ~x532 & ~x559 & ~x561 & ~x586 & ~x590 & ~x613 & ~x614 & ~x615 & ~x616 & ~x643 & ~x646 & ~x675 & ~x700 & ~x725 & ~x726 & ~x754 & ~x758 & ~x781;
assign c8337 = ~x14 & ~x204 & ~x229 & ~x281 & ~x288 & ~x769 & ~x770;
assign c8339 =  x556 & ~x339 & ~x365;
assign c8341 =  x749 & ~x26 & ~x363 & ~x643 & ~x649 & ~x668 & ~x724 & ~x751 & ~x752;
assign c8343 = ~x141 & ~x143 & ~x179 & ~x253 & ~x255 & ~x281 & ~x326 & ~x365 & ~x392 & ~x394 & ~x765;
assign c8345 =  x398 & ~x605 & ~x661;
assign c8347 =  x540 & ~x26 & ~x34 & ~x50 & ~x55 & ~x58 & ~x59 & ~x81 & ~x111 & ~x143 & ~x171 & ~x200 & ~x225 & ~x226 & ~x228 & ~x229 & ~x255 & ~x281 & ~x282 & ~x283 & ~x285 & ~x286 & ~x287 & ~x308 & ~x309 & ~x312 & ~x314 & ~x336 & ~x337 & ~x339 & ~x343 & ~x364 & ~x365 & ~x392 & ~x395 & ~x700 & ~x729 & ~x733 & ~x755 & ~x757 & ~x759 & ~x760 & ~x762;
assign c8349 = ~x2 & ~x5 & ~x13 & ~x14 & ~x15 & ~x31 & ~x42 & ~x86 & ~x112 & ~x169 & ~x252 & ~x253 & ~x280 & ~x338 & ~x342 & ~x364 & ~x366 & ~x368 & ~x392 & ~x394 & ~x395 & ~x396 & ~x420 & ~x424 & ~x425 & ~x448 & ~x449 & ~x450 & ~x451 & ~x452 & ~x453 & ~x477 & ~x478 & ~x480 & ~x587 & ~x756 & ~x781;
assign c8351 =  x406 &  x462 & ~x141 & ~x201 & ~x224 & ~x315;
assign c8353 = ~x2 & ~x13 & ~x14 & ~x26 & ~x32 & ~x140 & ~x422 & ~x424 & ~x478 & ~x501 & ~x505 & ~x507 & ~x533 & ~x583 & ~x586 & ~x590 & ~x592 & ~x593 & ~x612 & ~x615 & ~x616 & ~x619 & ~x639 & ~x648 & ~x668 & ~x697 & ~x700 & ~x702 & ~x729;
assign c8355 =  x599 &  x684 & ~x14 & ~x41 & ~x42 & ~x449 & ~x451 & ~x700 & ~x728;
assign c8357 = ~x227 & ~x281 & ~x312 & ~x374 & ~x765 & ~x766 & ~x768;
assign c8359 =  x267 & ~x72 & ~x232;
assign c8361 = ~x262 & ~x281 & ~x578;
assign c8363 =  x395 &  x423 &  x424 &  x443 & ~x621 & ~x762;
assign c8365 = ~x373;
assign c8367 = ~x143 & ~x151 & ~x178 & ~x179 & ~x403 & ~x743;
assign c8369 =  x533 &  x534;
assign c8371 = ~x179 & ~x208 & ~x423;
assign c8373 =  x361 & ~x316;
assign c8375 =  x47 &  x77 &  x116 &  x133 &  x173 & ~x82 & ~x85;
assign c8377 =  x737 & ~x2 & ~x5 & ~x14 & ~x27 & ~x33 & ~x115 & ~x167 & ~x195 & ~x255 & ~x308 & ~x336 & ~x337 & ~x370 & ~x422 & ~x454 & ~x479 & ~x671 & ~x756 & ~x760;
assign c8379 =  x593 & ~x14 & ~x280 & ~x310 & ~x341 & ~x365 & ~x366 & ~x367 & ~x394 & ~x420 & ~x423 & ~x450 & ~x559 & ~x756;
assign c8381 =  x499 &  x564 &  x612 &  x696 &  x724 & ~x109 & ~x365;
assign c8383 =  x69 &  x71 &  x72 &  x768 & ~x3 & ~x33 & ~x49 & ~x52 & ~x140 & ~x194 & ~x224 & ~x365 & ~x389 & ~x391 & ~x504 & ~x643;
assign c8385 =  x295 &  x434 & ~x5 & ~x8 & ~x24 & ~x25 & ~x26 & ~x27 & ~x50 & ~x52 & ~x56 & ~x82 & ~x83 & ~x85 & ~x86 & ~x88 & ~x90 & ~x111 & ~x112 & ~x113 & ~x116 & ~x118 & ~x138 & ~x145 & ~x146 & ~x161 & ~x169 & ~x171 & ~x172 & ~x173 & ~x174 & ~x191 & ~x192 & ~x193 & ~x197 & ~x198 & ~x200 & ~x201 & ~x218 & ~x219 & ~x225 & ~x226 & ~x228 & ~x247 & ~x254 & ~x255 & ~x256 & ~x280 & ~x281 & ~x283 & ~x308 & ~x309 & ~x335 & ~x336 & ~x338 & ~x364 & ~x533 & ~x562 & ~x588 & ~x641 & ~x642 & ~x644 & ~x669 & ~x672 & ~x674 & ~x675 & ~x697 & ~x698 & ~x701 & ~x725 & ~x753 & ~x754 & ~x759 & ~x760;
assign c8387 = ~x29 & ~x34 & ~x59 & ~x157 & ~x166 & ~x197 & ~x198 & ~x248 & ~x254 & ~x255 & ~x282 & ~x361 & ~x589 & ~x705 & ~x766 & ~x776;
assign c8389 =  x385 & ~x378 & ~x768;
assign c8391 =  x13 &  x15 &  x41 & ~x49 & ~x51;
assign c8393 =  x229 &  x444 &  x516 &  x572 & ~x169 & ~x193 & ~x306 & ~x334;
assign c8395 =  x344 & ~x224 & ~x308 & ~x389 & ~x390 & ~x418 & ~x423 & ~x547;
assign c8397 = ~x0 & ~x3 & ~x11 & ~x13 & ~x14 & ~x15 & ~x23 & ~x25 & ~x41 & ~x54 & ~x57 & ~x84 & ~x167 & ~x252 & ~x280 & ~x284 & ~x313 & ~x340 & ~x368 & ~x369 & ~x392 & ~x396 & ~x425 & ~x450 & ~x452 & ~x453 & ~x481 & ~x507 & ~x536 & ~x756;
assign c8399 =  x47 & ~x0 & ~x3 & ~x13 & ~x23 & ~x33 & ~x82 & ~x109 & ~x111 & ~x250 & ~x728 & ~x763;
assign c8401 = ~x319;
assign c8403 = ~x213 & ~x281 & ~x365 & ~x605 & ~x619 & ~x768;
assign c8405 =  x453 & ~x654;
assign c8407 = ~x286 & ~x562 & ~x578 & ~x593;
assign c8409 =  x360 &  x653 & ~x667;
assign c8411 = ~x282 & ~x283 & ~x309 & ~x313 & ~x617 & ~x660 & ~x739;
assign c8413 =  x174 & ~x20 & ~x83 & ~x225 & ~x263;
assign c8415 = ~x291 & ~x336 & ~x338 & ~x367 & ~x647;
assign c8417 =  x206 &  x374 &  x515 &  x632 & ~x14 & ~x71 & ~x112 & ~x167 & ~x393;
assign c8419 =  x123 &  x465 & ~x48 & ~x50 & ~x483 & ~x724;
assign c8421 =  x40 &  x41 &  x69 &  x516 & ~x48 & ~x333 & ~x337 & ~x392 & ~x450 & ~x558;
assign c8423 = ~x231 & ~x235 & ~x281 & ~x284 & ~x310 & ~x312 & ~x374 & ~x771;
assign c8425 = ~x16 & ~x46 & ~x60 & ~x70 & ~x110 & ~x112 & ~x125 & ~x140 & ~x149 & ~x151 & ~x171 & ~x172 & ~x198 & ~x207 & ~x230 & ~x254 & ~x258 & ~x262 & ~x281 & ~x310 & ~x311 & ~x312 & ~x338 & ~x705 & ~x714 & ~x726 & ~x745 & ~x748 & ~x751 & ~x755 & ~x757 & ~x767 & ~x768 & ~x770 & ~x771;
assign c8427 =  x134 &  x679 & ~x5 & ~x14 & ~x28 & ~x29 & ~x336 & ~x364 & ~x419 & ~x475 & ~x560 & ~x587 & ~x760 & ~x761 & ~x780;
assign c8429 =  x406 &  x462 &  x517 &  x545 &  x601 &  x711 & ~x1 & ~x27 & ~x32 & ~x139 & ~x196 & ~x222 & ~x303 & ~x330 & ~x341 & ~x397 & ~x415 & ~x505 & ~x560 & ~x564 & ~x612 & ~x641 & ~x647 & ~x672 & ~x701 & ~x725 & ~x783;
assign c8431 =  x101 &  x154 &  x536 &  x556 & ~x137 & ~x165 & ~x193 & ~x364;
assign c8433 = ~x78 & ~x110 & ~x198 & ~x309 & ~x551 & ~x557 & ~x590 & ~x649 & ~x701 & ~x703 & ~x734;
assign c8435 =  x344 & ~x354 & ~x391 & ~x417 & ~x447 & ~x644 & ~x701 & ~x775;
assign c8437 =  x70 & ~x85 & ~x141 & ~x169 & ~x504 & ~x699;
assign c8439 =  x41 &  x42 & ~x0 & ~x22 & ~x38 & ~x58 & ~x81 & ~x84 & ~x171 & ~x191 & ~x308 & ~x474 & ~x477 & ~x506 & ~x507 & ~x531 & ~x560 & ~x669 & ~x673 & ~x701 & ~x726;
assign c8441 = ~x261 & ~x523;
assign c8443 =  x98;
assign c8445 = ~x234 & ~x366 & ~x689;
assign c8447 =  x499 &  x526 & ~x1 & ~x28 & ~x29 & ~x138 & ~x139 & ~x141 & ~x253 & ~x280 & ~x309 & ~x310 & ~x335 & ~x337 & ~x419 & ~x447 & ~x587 & ~x700 & ~x748 & ~x766;
assign c8449 =  x445 & ~x143 & ~x310 & ~x740;
assign c8451 =  x569 & ~x112 & ~x393 & ~x421 & ~x450 & ~x478 & ~x617 & ~x701 & ~x702 & ~x745 & ~x765;
assign c8453 =  x510 & ~x139 & ~x198 & ~x200 & ~x224 & ~x254 & ~x256 & ~x282 & ~x310 & ~x311 & ~x312 & ~x313 & ~x336 & ~x337 & ~x338 & ~x340 & ~x662;
assign c8455 =  x67 &  x70 & ~x6 & ~x20 & ~x25 & ~x31 & ~x48 & ~x49 & ~x53 & ~x54 & ~x56 & ~x85 & ~x108 & ~x110 & ~x116 & ~x138 & ~x141 & ~x167 & ~x170 & ~x172 & ~x304 & ~x307 & ~x390 & ~x395 & ~x418 & ~x419 & ~x503 & ~x674 & ~x697 & ~x727 & ~x753 & ~x782;
assign c8457 =  x415 & ~x178 & ~x262 & ~x311 & ~x336 & ~x580;
assign c8459 = ~x208 & ~x550 & ~x607;
assign c8461 = ~x403 & ~x563 & ~x583 & ~x714;
assign c8463 =  x646;
assign c8465 =  x276 & ~x421 & ~x453;
assign c8467 =  x121 &  x129 &  x130 &  x159 &  x179 &  x186 &  x201 &  x275 &  x284 &  x287 &  x606 &  x635 &  x663 &  x691 & ~x80 & ~x137 & ~x140 & ~x194 & ~x250 & ~x363 & ~x531;
assign c8469 = ~x230 & ~x253 & ~x262 & ~x289 & ~x773;
assign c8471 =  x11 & ~x50 & ~x254;
assign c8473 = ~x121 & ~x148 & ~x262 & ~x311 & ~x317 & ~x318 & ~x396;
assign c8475 =  x436 &  x637 &  x653 &  x688 & ~x649 & ~x724;
assign c8477 =  x70 & ~x36 & ~x75 & ~x532;
assign c8479 = ~x84 & ~x151 & ~x248 & ~x253 & ~x255 & ~x311 & ~x689;
assign c8481 =  x259 &  x318 &  x538 &  x653 & ~x24 & ~x32 & ~x82 & ~x108 & ~x163 & ~x166 & ~x198 & ~x220 & ~x254 & ~x276 & ~x282 & ~x311 & ~x333 & ~x334 & ~x338 & ~x389 & ~x390 & ~x421 & ~x450 & ~x674 & ~x776;
assign c8483 =  x66 &  x288 &  x457 &  x541 &  x597 &  x625 &  x652 & ~x0 & ~x1 & ~x3 & ~x22 & ~x54 & ~x56 & ~x57 & ~x84 & ~x195 & ~x280 & ~x588 & ~x590 & ~x614 & ~x615 & ~x617 & ~x619 & ~x641 & ~x644 & ~x646 & ~x647 & ~x668 & ~x669 & ~x671 & ~x674 & ~x675 & ~x696 & ~x697 & ~x699 & ~x703 & ~x731 & ~x752 & ~x754 & ~x758 & ~x781 & ~x782 & ~x783;
assign c8485 =  x410 &  x415 &  x444 &  x466 &  x493 &  x494 &  x507 &  x508 &  x520 &  x546 & ~x52 & ~x56 & ~x58 & ~x137 & ~x139 & ~x166 & ~x222 & ~x251 & ~x252 & ~x253 & ~x337;
assign c8487 =  x172 &  x201 &  x219 &  x684 & ~x52 & ~x53;
assign c8489 =  x183 & ~x11 & ~x54 & ~x57 & ~x146 & ~x174 & ~x224 & ~x418 & ~x478 & ~x500 & ~x505 & ~x528 & ~x561 & ~x614 & ~x647 & ~x672;
assign c8491 =  x231 & ~x58 & ~x79 & ~x80 & ~x85 & ~x109 & ~x170 & ~x198 & ~x252 & ~x278 & ~x338 & ~x390 & ~x446 & ~x475 & ~x476 & ~x748;
assign c8493 = ~x230 & ~x309 & ~x340 & ~x715;
assign c8495 =  x374 &  x604 &  x605 &  x710 &  x739 & ~x52 & ~x336 & ~x413 & ~x424 & ~x502 & ~x506 & ~x531 & ~x564 & ~x616 & ~x619 & ~x646 & ~x675;
assign c8497 =  x107 &  x135 & ~x13 & ~x14 & ~x26 & ~x365 & ~x393;
assign c8499 =  x37 & ~x0 & ~x3 & ~x5 & ~x6 & ~x23 & ~x24 & ~x28 & ~x31 & ~x32 & ~x50 & ~x52 & ~x53 & ~x54 & ~x55 & ~x59 & ~x80 & ~x81 & ~x85 & ~x108 & ~x109 & ~x111 & ~x112 & ~x113 & ~x114 & ~x137 & ~x140 & ~x141 & ~x165 & ~x166 & ~x168 & ~x169 & ~x194 & ~x195 & ~x196 & ~x226 & ~x250 & ~x253 & ~x334 & ~x335 & ~x336 & ~x337 & ~x363 & ~x393 & ~x394 & ~x418 & ~x419 & ~x421 & ~x448 & ~x450 & ~x474 & ~x475 & ~x476 & ~x502 & ~x506 & ~x532 & ~x561 & ~x587 & ~x589 & ~x615 & ~x644 & ~x669 & ~x699 & ~x700 & ~x701 & ~x726 & ~x727 & ~x728 & ~x729 & ~x756 & ~x757 & ~x782;
assign c90 =  x237 &  x242 &  x351 &  x378 &  x381 &  x384 &  x407 &  x409 &  x412 &  x435 &  x437 &  x462 &  x491 &  x545 &  x573 & ~x6 & ~x30 & ~x59 & ~x61 & ~x63 & ~x115 & ~x117 & ~x140 & ~x141 & ~x149 & ~x176 & ~x199 & ~x225 & ~x226 & ~x228 & ~x258 & ~x285 & ~x288 & ~x309 & ~x316 & ~x336 & ~x344 & ~x393 & ~x398 & ~x425 & ~x426 & ~x700 & ~x729 & ~x730 & ~x771 & ~x773 & ~x774;
assign c92 =  x302 &  x330 &  x356 &  x359 &  x387 & ~x28 & ~x54 & ~x56 & ~x58 & ~x62 & ~x64 & ~x83 & ~x114 & ~x116 & ~x117 & ~x141 & ~x145 & ~x167 & ~x169 & ~x176 & ~x224 & ~x228 & ~x229 & ~x281 & ~x284 & ~x306 & ~x312 & ~x335 & ~x337 & ~x342 & ~x363 & ~x366 & ~x369 & ~x370 & ~x394 & ~x395 & ~x399 & ~x419 & ~x420 & ~x454 & ~x482 & ~x484 & ~x531 & ~x757;
assign c94 =  x387 &  x543 & ~x1 & ~x11 & ~x20 & ~x34 & ~x40 & ~x45 & ~x62 & ~x67 & ~x68 & ~x83 & ~x84 & ~x88 & ~x92 & ~x94 & ~x109 & ~x110 & ~x131 & ~x132 & ~x135 & ~x147 & ~x163 & ~x165 & ~x167 & ~x171 & ~x174 & ~x179 & ~x180 & ~x182 & ~x196 & ~x209 & ~x233 & ~x234 & ~x235 & ~x251 & ~x260 & ~x287 & ~x288 & ~x291 & ~x308 & ~x313 & ~x316 & ~x317 & ~x318 & ~x340 & ~x346 & ~x590 & ~x604 & ~x605 & ~x617 & ~x620 & ~x623 & ~x648 & ~x660 & ~x677 & ~x694 & ~x703 & ~x712 & ~x727 & ~x730 & ~x735 & ~x737 & ~x745 & ~x751 & ~x760 & ~x774 & ~x783;
assign c96 =  x276 &  x354 &  x524 & ~x55 & ~x77 & ~x94 & ~x176 & ~x216 & ~x287 & ~x576 & ~x660 & ~x720 & ~x721 & ~x750 & ~x780;
assign c98 =  x545 &  x557 &  x571 & ~x22 & ~x26 & ~x33 & ~x35 & ~x38 & ~x125 & ~x169 & ~x225 & ~x258 & ~x262 & ~x338 & ~x341 & ~x399 & ~x426 & ~x429 & ~x454 & ~x455 & ~x456 & ~x688 & ~x729 & ~x741 & ~x754 & ~x764 & ~x774 & ~x776 & ~x782;
assign c910 = ~x48 & ~x52 & ~x142 & ~x171 & ~x179 & ~x196 & ~x307 & ~x315 & ~x319 & ~x419 & ~x456 & ~x482 & ~x483 & ~x515 & ~x538 & ~x541 & ~x758;
assign c912 =  x534 & ~x14 & ~x29 & ~x54 & ~x74 & ~x78 & ~x100 & ~x106 & ~x107 & ~x108 & ~x131 & ~x142 & ~x144 & ~x145 & ~x179 & ~x200 & ~x208 & ~x224 & ~x230 & ~x235 & ~x280 & ~x284 & ~x336 & ~x339 & ~x340 & ~x343 & ~x368 & ~x370 & ~x393 & ~x398 & ~x420 & ~x427 & ~x428 & ~x687 & ~x689 & ~x704 & ~x707 & ~x712 & ~x715 & ~x732 & ~x740 & ~x747 & ~x752 & ~x754 & ~x769 & ~x774;
assign c914 =  x527 & ~x1 & ~x9 & ~x12 & ~x16 & ~x24 & ~x54 & ~x57 & ~x58 & ~x68 & ~x69 & ~x72 & ~x85 & ~x86 & ~x88 & ~x90 & ~x95 & ~x96 & ~x97 & ~x112 & ~x116 & ~x117 & ~x119 & ~x122 & ~x125 & ~x140 & ~x143 & ~x151 & ~x170 & ~x171 & ~x201 & ~x205 & ~x253 & ~x257 & ~x259 & ~x261 & ~x263 & ~x280 & ~x281 & ~x283 & ~x286 & ~x289 & ~x308 & ~x311 & ~x315 & ~x335 & ~x338 & ~x341 & ~x369 & ~x391 & ~x392 & ~x393 & ~x426 & ~x427 & ~x428 & ~x481 & ~x511 & ~x512 & ~x757 & ~x758;
assign c916 =  x298 & ~x52 & ~x53 & ~x77 & ~x185 & ~x364 & ~x577 & ~x606 & ~x684;
assign c918 =  x534 &  x551 &  x569 &  x572 & ~x5 & ~x18 & ~x29 & ~x68 & ~x81 & ~x113 & ~x226 & ~x233 & ~x284 & ~x335 & ~x337 & ~x371 & ~x400 & ~x428 & ~x644 & ~x659 & ~x660 & ~x677 & ~x705 & ~x727 & ~x737 & ~x748 & ~x771;
assign c920 =  x265 &  x293 &  x322 &  x348 &  x375 &  x409 &  x412 &  x431 &  x435 &  x437 &  x459 &  x460 &  x546 & ~x1 & ~x26 & ~x33 & ~x56 & ~x64 & ~x196 & ~x225 & ~x230 & ~x258 & ~x283 & ~x286 & ~x312 & ~x689 & ~x690 & ~x692 & ~x729 & ~x746 & ~x760 & ~x761 & ~x771 & ~x775 & ~x778;
assign c922 =  x327 &  x329 &  x352 &  x438 &  x493 &  x599 & ~x30 & ~x39 & ~x45 & ~x47 & ~x48 & ~x57 & ~x68 & ~x72 & ~x74 & ~x76 & ~x79 & ~x87 & ~x91 & ~x98 & ~x102 & ~x116 & ~x150 & ~x199 & ~x260 & ~x312 & ~x343 & ~x345 & ~x369 & ~x397 & ~x399 & ~x428 & ~x702 & ~x730 & ~x739;
assign c924 =  x110;
assign c926 =  x19;
assign c928 =  x539 & ~x16 & ~x344 & ~x578 & ~x654 & ~x780;
assign c930 =  x299 &  x328 &  x415 &  x435 &  x449 &  x468 &  x469 &  x490 &  x541 & ~x3 & ~x10 & ~x14 & ~x27 & ~x72 & ~x88 & ~x144 & ~x197 & ~x208 & ~x289 & ~x560 & ~x618 & ~x653 & ~x689 & ~x701 & ~x714 & ~x745 & ~x754 & ~x755 & ~x760;
assign c932 =  x665 & ~x13 & ~x29 & ~x43 & ~x75 & ~x78 & ~x80 & ~x83 & ~x99 & ~x108 & ~x113 & ~x125 & ~x141 & ~x171 & ~x205 & ~x255 & ~x280 & ~x337 & ~x363 & ~x449 & ~x748 & ~x779;
assign c934 =  x277 &  x417 & ~x154 & ~x155 & ~x566;
assign c936 = ~x22 & ~x195 & ~x287 & ~x318 & ~x334 & ~x374 & ~x428 & ~x566 & ~x596 & ~x597 & ~x598 & ~x729 & ~x773;
assign c938 =  x479 &  x507 &  x573 & ~x227 & ~x398;
assign c940 =  x218 &  x273 &  x300 &  x325 &  x329 &  x351 &  x352 &  x356 &  x358 &  x378 &  x379 &  x381 &  x383 &  x385 &  x406 &  x407 &  x410 &  x435 &  x436 &  x438 &  x439 &  x463 &  x490 &  x491 &  x492 &  x494 &  x546 &  x573 &  x599 &  x600 & ~x8 & ~x9 & ~x28 & ~x29 & ~x32 & ~x33 & ~x56 & ~x59 & ~x60 & ~x62 & ~x86 & ~x87 & ~x90 & ~x91 & ~x113 & ~x118 & ~x120 & ~x139 & ~x145 & ~x147 & ~x148 & ~x168 & ~x170 & ~x172 & ~x196 & ~x198 & ~x228 & ~x252 & ~x256 & ~x260 & ~x280 & ~x281 & ~x283 & ~x286 & ~x311 & ~x336 & ~x341 & ~x342 & ~x365 & ~x367 & ~x369 & ~x371 & ~x393 & ~x394 & ~x397 & ~x398 & ~x427 & ~x448 & ~x453 & ~x454 & ~x756 & ~x758 & ~x759;
assign c942 =  x190 &  x218 &  x240 &  x243 &  x244 &  x245 &  x268 &  x271 &  x272 &  x273 &  x295 &  x296 &  x300 &  x323 &  x324 &  x325 &  x326 &  x327 &  x328 &  x329 &  x351 &  x352 &  x356 &  x359 &  x379 &  x380 &  x384 &  x385 &  x409 &  x411 &  x412 &  x463 &  x489 &  x492 &  x545 & ~x0 & ~x2 & ~x3 & ~x4 & ~x6 & ~x10 & ~x29 & ~x30 & ~x31 & ~x32 & ~x34 & ~x36 & ~x38 & ~x55 & ~x56 & ~x57 & ~x58 & ~x61 & ~x62 & ~x63 & ~x64 & ~x84 & ~x85 & ~x88 & ~x113 & ~x114 & ~x115 & ~x116 & ~x120 & ~x139 & ~x140 & ~x141 & ~x142 & ~x144 & ~x169 & ~x171 & ~x174 & ~x197 & ~x198 & ~x199 & ~x224 & ~x225 & ~x227 & ~x252 & ~x254 & ~x256 & ~x257 & ~x280 & ~x282 & ~x283 & ~x308 & ~x309 & ~x314 & ~x336 & ~x337 & ~x339 & ~x364 & ~x365 & ~x366 & ~x368 & ~x393 & ~x394 & ~x395 & ~x397 & ~x426 & ~x448 & ~x452 & ~x532 & ~x728 & ~x759 & ~x783;
assign c944 =  x380 &  x382 &  x445 & ~x11 & ~x16 & ~x22 & ~x23 & ~x25 & ~x121 & ~x123 & ~x127 & ~x158 & ~x257 & ~x287 & ~x364 & ~x700 & ~x749 & ~x752;
assign c946 =  x540 & ~x3 & ~x9 & ~x67 & ~x93 & ~x98 & ~x156 & ~x164 & ~x257 & ~x281 & ~x338 & ~x630 & ~x685 & ~x689 & ~x740 & ~x741 & ~x745 & ~x753 & ~x775;
assign c948 =  x382 &  x415 &  x451 & ~x63 & ~x65 & ~x100 & ~x156 & ~x157 & ~x194 & ~x563 & ~x622 & ~x664 & ~x719 & ~x751 & ~x779 & ~x783;
assign c950 =  x604 &  x630 &  x648 &  x656 &  x658 & ~x1 & ~x2 & ~x3 & ~x4 & ~x6 & ~x7 & ~x8 & ~x9 & ~x10 & ~x13 & ~x24 & ~x26 & ~x27 & ~x28 & ~x29 & ~x30 & ~x31 & ~x32 & ~x33 & ~x34 & ~x35 & ~x36 & ~x38 & ~x52 & ~x53 & ~x54 & ~x55 & ~x57 & ~x58 & ~x59 & ~x60 & ~x61 & ~x62 & ~x63 & ~x64 & ~x83 & ~x84 & ~x85 & ~x87 & ~x89 & ~x90 & ~x92 & ~x111 & ~x112 & ~x113 & ~x114 & ~x116 & ~x117 & ~x118 & ~x121 & ~x140 & ~x141 & ~x142 & ~x143 & ~x144 & ~x145 & ~x168 & ~x169 & ~x170 & ~x171 & ~x175 & ~x196 & ~x197 & ~x198 & ~x199 & ~x200 & ~x225 & ~x226 & ~x227 & ~x228 & ~x229 & ~x231 & ~x232 & ~x252 & ~x253 & ~x254 & ~x256 & ~x257 & ~x258 & ~x260 & ~x261 & ~x281 & ~x283 & ~x284 & ~x285 & ~x286 & ~x287 & ~x308 & ~x309 & ~x313 & ~x314 & ~x315 & ~x337 & ~x341 & ~x342 & ~x343 & ~x344 & ~x364 & ~x365 & ~x366 & ~x367 & ~x368 & ~x369 & ~x370 & ~x371 & ~x372 & ~x392 & ~x393 & ~x394 & ~x395 & ~x397 & ~x399 & ~x400 & ~x420 & ~x423 & ~x424 & ~x425 & ~x426 & ~x427 & ~x428 & ~x448 & ~x449 & ~x450 & ~x452 & ~x476 & ~x504 & ~x700 & ~x701 & ~x727 & ~x729 & ~x758 & ~x759 & ~x761 & ~x772 & ~x773 & ~x774;
assign c952 =  x129 &  x157 &  x185 &  x186 &  x245 &  x324 &  x352 &  x379 &  x380 &  x384 &  x385 &  x409 &  x410 &  x413 &  x441 &  x466 &  x491 &  x494 & ~x4 & ~x5 & ~x6 & ~x7 & ~x25 & ~x27 & ~x29 & ~x30 & ~x32 & ~x33 & ~x37 & ~x56 & ~x58 & ~x61 & ~x65 & ~x86 & ~x87 & ~x91 & ~x114 & ~x117 & ~x118 & ~x140 & ~x141 & ~x142 & ~x144 & ~x168 & ~x170 & ~x176 & ~x195 & ~x196 & ~x197 & ~x198 & ~x225 & ~x228 & ~x252 & ~x254 & ~x256 & ~x282 & ~x283 & ~x286 & ~x308 & ~x310 & ~x336 & ~x337 & ~x340 & ~x341 & ~x364 & ~x365 & ~x392 & ~x393 & ~x396 & ~x397 & ~x398 & ~x476 & ~x728 & ~x729 & ~x756 & ~x757 & ~x758 & ~x773 & ~x776;
assign c954 =  x219 &  x244 &  x247 &  x272 &  x275 &  x276 &  x329 &  x331 &  x332 &  x388 &  x485 &  x487 &  x489 &  x546 & ~x2 & ~x3 & ~x36 & ~x54 & ~x65 & ~x88 & ~x118 & ~x145 & ~x201 & ~x226 & ~x230 & ~x252 & ~x253 & ~x257 & ~x312 & ~x313 & ~x340 & ~x758 & ~x759 & ~x778 & ~x782;
assign c956 =  x494 &  x614 & ~x8 & ~x20 & ~x80 & ~x113 & ~x144 & ~x200 & ~x230 & ~x316 & ~x399 & ~x560 & ~x659 & ~x733 & ~x738 & ~x767;
assign c958 =  x354 &  x379 &  x492 &  x561 &  x640 & ~x1 & ~x4 & ~x7 & ~x29 & ~x47 & ~x60 & ~x67 & ~x77 & ~x82 & ~x84 & ~x86 & ~x87 & ~x94 & ~x110 & ~x114 & ~x141 & ~x176 & ~x200 & ~x228 & ~x233 & ~x257 & ~x260 & ~x285 & ~x313 & ~x314 & ~x337 & ~x342 & ~x369 & ~x672 & ~x674 & ~x734 & ~x737 & ~x738 & ~x742 & ~x745 & ~x752 & ~x761 & ~x766 & ~x772 & ~x780 & ~x782;
assign c960 =  x578 &  x580 &  x614 &  x642 & ~x1 & ~x5 & ~x6 & ~x16 & ~x20 & ~x21 & ~x58 & ~x63 & ~x67 & ~x69 & ~x83 & ~x94 & ~x114 & ~x143 & ~x199 & ~x204 & ~x223 & ~x229 & ~x230 & ~x236 & ~x290 & ~x291 & ~x292 & ~x317 & ~x319 & ~x335 & ~x343 & ~x363 & ~x370 & ~x372 & ~x394 & ~x448 & ~x476 & ~x644 & ~x758 & ~x759;
assign c962 =  x298 & ~x0 & ~x1 & ~x5 & ~x7 & ~x11 & ~x23 & ~x24 & ~x26 & ~x27 & ~x29 & ~x32 & ~x33 & ~x34 & ~x35 & ~x38 & ~x39 & ~x55 & ~x57 & ~x58 & ~x59 & ~x61 & ~x62 & ~x63 & ~x64 & ~x66 & ~x88 & ~x89 & ~x113 & ~x116 & ~x118 & ~x120 & ~x122 & ~x123 & ~x140 & ~x141 & ~x142 & ~x143 & ~x144 & ~x148 & ~x151 & ~x169 & ~x170 & ~x171 & ~x173 & ~x174 & ~x178 & ~x179 & ~x195 & ~x196 & ~x197 & ~x198 & ~x200 & ~x201 & ~x225 & ~x228 & ~x231 & ~x232 & ~x252 & ~x255 & ~x258 & ~x259 & ~x261 & ~x262 & ~x263 & ~x281 & ~x282 & ~x283 & ~x288 & ~x291 & ~x312 & ~x314 & ~x316 & ~x318 & ~x335 & ~x337 & ~x341 & ~x342 & ~x346 & ~x368 & ~x369 & ~x370 & ~x372 & ~x373 & ~x398 & ~x399 & ~x400 & ~x421 & ~x423 & ~x424 & ~x426 & ~x427 & ~x428 & ~x448 & ~x455 & ~x476 & ~x511 & ~x512 & ~x644 & ~x700 & ~x718 & ~x728 & ~x745 & ~x755 & ~x757 & ~x758 & ~x760 & ~x774 & ~x781 & ~x783;
assign c964 =  x138;
assign c966 =  x218 &  x220 &  x246 &  x271 &  x303 &  x304 &  x331 &  x352 &  x436 &  x493 & ~x1 & ~x3 & ~x4 & ~x54 & ~x172 & ~x254 & ~x280 & ~x281 & ~x314 & ~x367 & ~x448 & ~x693 & ~x729 & ~x758 & ~x764 & ~x779;
assign c968 =  x581 &  x614 & ~x7 & ~x92 & ~x177 & ~x260 & ~x289 & ~x312 & ~x662 & ~x671 & ~x731;
assign c970 =  x277 &  x301 &  x388 &  x413 &  x628 &  x629 &  x641 & ~x9 & ~x25 & ~x26 & ~x29 & ~x31 & ~x33 & ~x34 & ~x36 & ~x41 & ~x42 & ~x57 & ~x85 & ~x92 & ~x93 & ~x95 & ~x112 & ~x118 & ~x121 & ~x144 & ~x169 & ~x175 & ~x199 & ~x200 & ~x227 & ~x229 & ~x252 & ~x253 & ~x255 & ~x282 & ~x284 & ~x286 & ~x309 & ~x311 & ~x313 & ~x316 & ~x317 & ~x336 & ~x337 & ~x340 & ~x367 & ~x369 & ~x449 & ~x700 & ~x701 & ~x702 & ~x729 & ~x730 & ~x732 & ~x733 & ~x756 & ~x765 & ~x778 & ~x782 & ~x783;
assign c972 =  x354 &  x378 &  x381 &  x414 &  x438 &  x440 &  x463 &  x464 &  x545 &  x547 &  x573 &  x601 &  x683 &  x684 & ~x0 & ~x2 & ~x3 & ~x7 & ~x29 & ~x30 & ~x31 & ~x34 & ~x35 & ~x57 & ~x58 & ~x61 & ~x62 & ~x84 & ~x85 & ~x87 & ~x93 & ~x118 & ~x120 & ~x141 & ~x142 & ~x146 & ~x149 & ~x170 & ~x172 & ~x173 & ~x174 & ~x176 & ~x199 & ~x200 & ~x205 & ~x225 & ~x231 & ~x258 & ~x280 & ~x281 & ~x284 & ~x288 & ~x308 & ~x309 & ~x310 & ~x339 & ~x344 & ~x365 & ~x367 & ~x368 & ~x369 & ~x426 & ~x428 & ~x449 & ~x476 & ~x479 & ~x504 & ~x509 & ~x728 & ~x757 & ~x759 & ~x782 & ~x783;
assign c974 = ~x2 & ~x3 & ~x6 & ~x7 & ~x9 & ~x10 & ~x11 & ~x25 & ~x27 & ~x29 & ~x30 & ~x34 & ~x36 & ~x37 & ~x53 & ~x57 & ~x60 & ~x64 & ~x66 & ~x84 & ~x85 & ~x86 & ~x87 & ~x88 & ~x89 & ~x90 & ~x93 & ~x94 & ~x111 & ~x112 & ~x114 & ~x116 & ~x117 & ~x118 & ~x141 & ~x142 & ~x143 & ~x145 & ~x146 & ~x147 & ~x148 & ~x149 & ~x150 & ~x168 & ~x169 & ~x170 & ~x173 & ~x174 & ~x177 & ~x180 & ~x199 & ~x200 & ~x201 & ~x203 & ~x207 & ~x229 & ~x233 & ~x234 & ~x251 & ~x254 & ~x255 & ~x256 & ~x257 & ~x263 & ~x279 & ~x285 & ~x289 & ~x291 & ~x306 & ~x307 & ~x308 & ~x309 & ~x311 & ~x313 & ~x314 & ~x316 & ~x317 & ~x318 & ~x319 & ~x334 & ~x335 & ~x338 & ~x339 & ~x342 & ~x345 & ~x346 & ~x363 & ~x364 & ~x367 & ~x370 & ~x371 & ~x372 & ~x373 & ~x374 & ~x392 & ~x393 & ~x394 & ~x395 & ~x396 & ~x397 & ~x398 & ~x399 & ~x400 & ~x401 & ~x402 & ~x419 & ~x422 & ~x423 & ~x424 & ~x425 & ~x426 & ~x448 & ~x449 & ~x452 & ~x453 & ~x457 & ~x475 & ~x476 & ~x478 & ~x479 & ~x481 & ~x482 & ~x483 & ~x484 & ~x539 & ~x728 & ~x730 & ~x745 & ~x756 & ~x757 & ~x758 & ~x760 & ~x771 & ~x772 & ~x773 & ~x783;
assign c976 =  x222 &  x250 &  x324 &  x356 &  x358 &  x379 &  x385 &  x409 &  x434 & ~x5 & ~x15 & ~x42 & ~x64 & ~x117 & ~x139 & ~x147 & ~x259 & ~x261 & ~x367;
assign c978 = ~x39 & ~x107 & ~x141 & ~x374 & ~x439;
assign c980 =  x413 &  x469 &  x493 &  x496 & ~x1 & ~x32 & ~x57 & ~x59 & ~x64 & ~x84 & ~x85 & ~x111 & ~x167 & ~x226 & ~x253 & ~x256 & ~x307 & ~x315 & ~x335 & ~x342 & ~x344 & ~x363 & ~x367 & ~x398 & ~x426 & ~x427 & ~x428 & ~x455 & ~x565 & ~x701 & ~x746 & ~x747 & ~x758;
assign c982 =  x358 &  x445 &  x564 & ~x5 & ~x7 & ~x8 & ~x30 & ~x38 & ~x50 & ~x53 & ~x73 & ~x80 & ~x92 & ~x102 & ~x113 & ~x146 & ~x168 & ~x203 & ~x229 & ~x260 & ~x308 & ~x310 & ~x342 & ~x366 & ~x370 & ~x422 & ~x428 & ~x750 & ~x756 & ~x757;
assign c984 =  x269 &  x299 &  x324 &  x325 &  x327 &  x354 &  x358 &  x409 &  x414 &  x465 &  x545 &  x575 &  x599 &  x602 &  x626 & ~x0 & ~x7 & ~x9 & ~x26 & ~x31 & ~x32 & ~x38 & ~x58 & ~x60 & ~x62 & ~x85 & ~x87 & ~x93 & ~x112 & ~x118 & ~x119 & ~x143 & ~x144 & ~x147 & ~x169 & ~x173 & ~x196 & ~x197 & ~x198 & ~x200 & ~x201 & ~x224 & ~x226 & ~x227 & ~x230 & ~x232 & ~x254 & ~x255 & ~x256 & ~x261 & ~x281 & ~x310 & ~x316 & ~x317 & ~x336 & ~x367 & ~x370 & ~x372 & ~x396 & ~x397 & ~x419 & ~x421 & ~x447 & ~x531 & ~x560 & ~x671 & ~x728 & ~x758 & ~x773;
assign c986 =  x212 &  x268 &  x324 &  x353 &  x498 &  x499 &  x542 & ~x0 & ~x8 & ~x12 & ~x23 & ~x33 & ~x41 & ~x62 & ~x176 & ~x177 & ~x225 & ~x226 & ~x341 & ~x362 & ~x367 & ~x368 & ~x393 & ~x690 & ~x731 & ~x740 & ~x776;
assign c988 =  x329 &  x357 &  x383 &  x385 &  x413 & ~x2 & ~x5 & ~x8 & ~x25 & ~x29 & ~x30 & ~x34 & ~x52 & ~x64 & ~x69 & ~x92 & ~x106 & ~x146 & ~x148 & ~x174 & ~x203 & ~x313 & ~x314 & ~x365 & ~x455 & ~x663 & ~x700 & ~x709 & ~x776;
assign c990 =  x382 &  x423 &  x491 & ~x11 & ~x77 & ~x121 & ~x134 & ~x135 & ~x136 & ~x257 & ~x261 & ~x671 & ~x729 & ~x759 & ~x771;
assign c992 =  x249 &  x277 & ~x11 & ~x17 & ~x49 & ~x68 & ~x83 & ~x106 & ~x115 & ~x140 & ~x142 & ~x206 & ~x253 & ~x289 & ~x392 & ~x482 & ~x692 & ~x693;
assign c994 =  x506 &  x562 &  x592 &  x593 &  x602 &  x612 & ~x10 & ~x15 & ~x18 & ~x55 & ~x60 & ~x69 & ~x76 & ~x116 & ~x124 & ~x126 & ~x147 & ~x168 & ~x172 & ~x203 & ~x616 & ~x701 & ~x709 & ~x728 & ~x748 & ~x749 & ~x751 & ~x758;
assign c996 =  x327 &  x575 &  x598 & ~x11 & ~x16 & ~x38 & ~x42 & ~x47 & ~x48 & ~x52 & ~x78 & ~x95 & ~x97 & ~x110 & ~x117 & ~x121 & ~x130 & ~x133 & ~x169 & ~x174 & ~x199 & ~x204 & ~x254 & ~x282 & ~x292 & ~x315 & ~x342 & ~x393 & ~x421 & ~x427 & ~x662 & ~x671 & ~x694 & ~x709 & ~x717 & ~x727 & ~x740 & ~x744 & ~x745 & ~x759;
assign c998 =  x293 &  x300 &  x301 &  x349 &  x351 &  x360 &  x377 &  x378 &  x384 &  x388 &  x404 &  x411 &  x416 &  x463 & ~x11 & ~x25 & ~x51 & ~x58 & ~x99 & ~x119 & ~x201 & ~x202 & ~x226 & ~x227 & ~x228 & ~x285 & ~x308 & ~x340 & ~x365 & ~x678 & ~x683 & ~x689 & ~x699 & ~x763 & ~x772 & ~x775;
assign c9100 =  x295 &  x328 &  x378 &  x386 &  x414 &  x435 &  x463 &  x467 &  x496 &  x547 &  x576 &  x582 &  x599 &  x603 & ~x35 & ~x37 & ~x59 & ~x64 & ~x65 & ~x86 & ~x87 & ~x88 & ~x118 & ~x142 & ~x167 & ~x169 & ~x170 & ~x200 & ~x205 & ~x222 & ~x252 & ~x254 & ~x279 & ~x282 & ~x284 & ~x286 & ~x307 & ~x316 & ~x337 & ~x366 & ~x371 & ~x392 & ~x394 & ~x397 & ~x476 & ~x504 & ~x532 & ~x700 & ~x760 & ~x761 & ~x783;
assign c9102 =  x516 & ~x44 & ~x85 & ~x115 & ~x178 & ~x180 & ~x225 & ~x374 & ~x589 & ~x605 & ~x624 & ~x765 & ~x779;
assign c9104 =  x580 & ~x3 & ~x29 & ~x41 & ~x49 & ~x120 & ~x122 & ~x129 & ~x139 & ~x170 & ~x253 & ~x280 & ~x286 & ~x290 & ~x316 & ~x424 & ~x426 & ~x429 & ~x450 & ~x457;
assign c9106 =  x213 &  x270 &  x296 &  x298 &  x299 &  x327 &  x355 &  x380 &  x381 &  x385 &  x463 &  x519 &  x548 &  x573 & ~x1 & ~x2 & ~x8 & ~x9 & ~x27 & ~x28 & ~x31 & ~x33 & ~x36 & ~x55 & ~x60 & ~x63 & ~x64 & ~x84 & ~x89 & ~x90 & ~x92 & ~x116 & ~x117 & ~x120 & ~x140 & ~x142 & ~x144 & ~x147 & ~x167 & ~x171 & ~x196 & ~x198 & ~x200 & ~x203 & ~x205 & ~x227 & ~x228 & ~x230 & ~x252 & ~x253 & ~x254 & ~x255 & ~x259 & ~x281 & ~x282 & ~x284 & ~x287 & ~x288 & ~x307 & ~x309 & ~x313 & ~x314 & ~x339 & ~x342 & ~x364 & ~x365 & ~x366 & ~x367 & ~x368 & ~x369 & ~x370 & ~x371 & ~x372 & ~x373 & ~x396 & ~x398 & ~x399 & ~x421 & ~x425 & ~x426 & ~x447 & ~x448 & ~x451 & ~x456 & ~x478 & ~x479 & ~x728 & ~x758 & ~x760 & ~x781 & ~x782;
assign c9108 = ~x182 & ~x207 & ~x263 & ~x335 & ~x406 & ~x481 & ~x511 & ~x541 & ~x744;
assign c9110 =  x161 &  x162 &  x164 &  x187 &  x190 &  x192 &  x212 &  x213 &  x214 &  x217 &  x218 &  x270 &  x273 &  x327 &  x328 &  x357 &  x385 &  x386 &  x410 &  x411 &  x548 &  x549 &  x572 & ~x28 & ~x30 & ~x31 & ~x32 & ~x38 & ~x55 & ~x58 & ~x59 & ~x62 & ~x63 & ~x84 & ~x86 & ~x89 & ~x90 & ~x91 & ~x115 & ~x116 & ~x118 & ~x142 & ~x143 & ~x145 & ~x148 & ~x149 & ~x224 & ~x225 & ~x228 & ~x229 & ~x230 & ~x254 & ~x279 & ~x311 & ~x314 & ~x315 & ~x336 & ~x341 & ~x343 & ~x364 & ~x367 & ~x368 & ~x371 & ~x425 & ~x452 & ~x728 & ~x757;
assign c9112 =  x194;
assign c9114 =  x299 &  x324 &  x361 &  x434 &  x466 & ~x13 & ~x42 & ~x74 & ~x92 & ~x100 & ~x141 & ~x172 & ~x186 & ~x203 & ~x226 & ~x315 & ~x559 & ~x605 & ~x622 & ~x688 & ~x689 & ~x697 & ~x737 & ~x743 & ~x774;
assign c9116 =  x267 &  x275 &  x324 &  x325 &  x349 &  x416 &  x471 &  x473 &  x486 &  x512 &  x555 & ~x11 & ~x36 & ~x76 & ~x94 & ~x169 & ~x284 & ~x289 & ~x366 & ~x722;
assign c9118 =  x181 &  x237 &  x245 &  x349 &  x351 &  x383 &  x384 &  x434 &  x490 &  x518 &  x599 & ~x3 & ~x5 & ~x6 & ~x10 & ~x29 & ~x82 & ~x116 & ~x117 & ~x168 & ~x171 & ~x226 & ~x336 & ~x340 & ~x364 & ~x393 & ~x394 & ~x729 & ~x761 & ~x772;
assign c9120 =  x103 &  x156 &  x159 &  x160 &  x186 &  x188 &  x211 &  x213 &  x301 &  x328 &  x330 &  x354 &  x378 &  x603 &  x648;
assign c9122 =  x274 &  x415 &  x597 &  x613 & ~x11 & ~x31 & ~x32 & ~x65 & ~x86 & ~x87 & ~x117 & ~x139 & ~x225 & ~x227 & ~x280 & ~x316 & ~x339 & ~x633 & ~x659 & ~x701 & ~x744 & ~x776;
assign c9124 =  x408 &  x413 &  x519 & ~x60 & ~x87 & ~x91 & ~x141 & ~x217 & ~x258 & ~x288 & ~x314 & ~x559 & ~x560 & ~x564;
assign c9126 =  x605 & ~x3 & ~x4 & ~x6 & ~x13 & ~x30 & ~x35 & ~x36 & ~x56 & ~x57 & ~x58 & ~x59 & ~x60 & ~x62 & ~x64 & ~x66 & ~x87 & ~x112 & ~x122 & ~x140 & ~x142 & ~x143 & ~x144 & ~x145 & ~x149 & ~x150 & ~x171 & ~x174 & ~x178 & ~x179 & ~x196 & ~x198 & ~x203 & ~x204 & ~x224 & ~x225 & ~x226 & ~x227 & ~x291 & ~x307 & ~x308 & ~x311 & ~x312 & ~x314 & ~x315 & ~x335 & ~x339 & ~x365 & ~x402 & ~x421 & ~x422 & ~x423 & ~x429 & ~x456 & ~x457 & ~x476 & ~x482 & ~x483 & ~x484 & ~x720 & ~x730 & ~x744 & ~x746 & ~x757 & ~x758 & ~x760 & ~x763 & ~x764 & ~x772 & ~x773 & ~x774 & ~x775;
assign c9128 =  x351 & ~x83 & ~x88 & ~x139 & ~x176 & ~x195 & ~x214 & ~x313 & ~x399 & ~x681;
assign c9130 =  x409 &  x489 &  x491 &  x501 &  x520 &  x527 &  x535 &  x544 & ~x8 & ~x46 & ~x79 & ~x229 & ~x285 & ~x337 & ~x371 & ~x448 & ~x606 & ~x711;
assign c9132 = ~x14 & ~x63 & ~x64 & ~x66 & ~x76 & ~x80 & ~x89 & ~x118 & ~x142 & ~x169 & ~x171 & ~x178 & ~x258 & ~x263 & ~x284 & ~x344 & ~x368 & ~x396 & ~x400 & ~x424 & ~x447 & ~x448 & ~x453 & ~x454 & ~x458 & ~x594;
assign c9134 =  x376 &  x409 &  x411 &  x434 &  x490 &  x627 & ~x2 & ~x6 & ~x7 & ~x19 & ~x25 & ~x38 & ~x53 & ~x56 & ~x57 & ~x58 & ~x87 & ~x92 & ~x116 & ~x120 & ~x142 & ~x143 & ~x175 & ~x176 & ~x178 & ~x225 & ~x226 & ~x228 & ~x229 & ~x231 & ~x254 & ~x285 & ~x287 & ~x315 & ~x316 & ~x336 & ~x342 & ~x393 & ~x397 & ~x662 & ~x701 & ~x702 & ~x730 & ~x742 & ~x746 & ~x762 & ~x771 & ~x782;
assign c9136 =  x354 &  x356 &  x358 &  x384 &  x387 &  x467 &  x496 & ~x8 & ~x11 & ~x26 & ~x30 & ~x31 & ~x36 & ~x57 & ~x63 & ~x65 & ~x86 & ~x112 & ~x143 & ~x147 & ~x167 & ~x169 & ~x223 & ~x224 & ~x225 & ~x229 & ~x251 & ~x255 & ~x307 & ~x308 & ~x311 & ~x335 & ~x343 & ~x369 & ~x373 & ~x395 & ~x397 & ~x475 & ~x509 & ~x728 & ~x762 & ~x772 & ~x783;
assign c9138 =  x298 & ~x0 & ~x22 & ~x59 & ~x87 & ~x94 & ~x112 & ~x126 & ~x144 & ~x168 & ~x199 & ~x200 & ~x207 & ~x208 & ~x232 & ~x234 & ~x235 & ~x257 & ~x289 & ~x291 & ~x307 & ~x337 & ~x343 & ~x363 & ~x369 & ~x373 & ~x391 & ~x393 & ~x396 & ~x397 & ~x399 & ~x401 & ~x425 & ~x426 & ~x448 & ~x455 & ~x456 & ~x457 & ~x479 & ~x481 & ~x482 & ~x483 & ~x760 & ~x773;
assign c9140 =  x245 &  x269 &  x295 &  x351 &  x354 &  x358 &  x409 &  x486 &  x501 &  x570 & ~x30 & ~x66 & ~x91 & ~x119 & ~x228 & ~x232 & ~x286 & ~x287 & ~x336 & ~x337 & ~x340 & ~x342 & ~x369 & ~x616 & ~x671 & ~x720 & ~x744 & ~x745 & ~x776;
assign c9142 =  x461 &  x462 &  x549 &  x562 &  x571 &  x583 & ~x10 & ~x16 & ~x39 & ~x74 & ~x78 & ~x91 & ~x119 & ~x143 & ~x167 & ~x171 & ~x177 & ~x283 & ~x335 & ~x392 & ~x394 & ~x396 & ~x476 & ~x739 & ~x749 & ~x758 & ~x781;
assign c9144 =  x250 &  x278 &  x409 &  x410 &  x614 & ~x117 & ~x147 & ~x308 & ~x338;
assign c9146 =  x212 &  x243 &  x299 &  x324 &  x355 &  x468 &  x522 &  x528 & ~x16 & ~x38 & ~x42 & ~x59 & ~x78 & ~x81 & ~x94 & ~x101 & ~x109 & ~x119 & ~x146 & ~x147 & ~x168 & ~x368 & ~x369 & ~x392 & ~x687 & ~x688 & ~x732 & ~x737 & ~x739 & ~x744 & ~x755 & ~x760 & ~x774;
assign c9148 = ~x0 & ~x48 & ~x54 & ~x146 & ~x172 & ~x259 & ~x453 & ~x455 & ~x456 & ~x482 & ~x483 & ~x485 & ~x486 & ~x513 & ~x594;
assign c9150 =  x299 &  x354 &  x355 &  x376 &  x378 &  x434 &  x490 &  x494 &  x497 & ~x20 & ~x23 & ~x39 & ~x44 & ~x45 & ~x60 & ~x70 & ~x98 & ~x107 & ~x132 & ~x152 & ~x156 & ~x199 & ~x255 & ~x260 & ~x262 & ~x311 & ~x342 & ~x343 & ~x344 & ~x587 & ~x588 & ~x595 & ~x619 & ~x643 & ~x651 & ~x663 & ~x670 & ~x672 & ~x687 & ~x691 & ~x697 & ~x698 & ~x702 & ~x704 & ~x728 & ~x733 & ~x745 & ~x776 & ~x779 & ~x782;
assign c9152 =  x240 &  x270 &  x323 &  x350 &  x378 &  x379 &  x386 &  x407 &  x409 &  x414 &  x438 &  x440 &  x462 &  x489 &  x490 &  x492 &  x545 &  x546 &  x652 &  x653 &  x655 & ~x7 & ~x25 & ~x62 & ~x63 & ~x84 & ~x85 & ~x118 & ~x120 & ~x140 & ~x141 & ~x149 & ~x230 & ~x231 & ~x252 & ~x255 & ~x282 & ~x284 & ~x287 & ~x311 & ~x363 & ~x369 & ~x371 & ~x420 & ~x422 & ~x425 & ~x426 & ~x476 & ~x728 & ~x757 & ~x761;
assign c9154 =  x688 &  x715 &  x735 &  x737 &  x740 & ~x482 & ~x484 & ~x509 & ~x510;
assign c9156 = ~x13 & ~x69 & ~x96 & ~x104 & ~x140 & ~x182 & ~x210 & ~x289 & ~x317 & ~x429 & ~x509 & ~x510 & ~x512 & ~x747;
assign c9158 = ~x3 & ~x5 & ~x6 & ~x7 & ~x8 & ~x11 & ~x27 & ~x29 & ~x32 & ~x36 & ~x86 & ~x89 & ~x114 & ~x119 & ~x140 & ~x141 & ~x142 & ~x144 & ~x146 & ~x147 & ~x167 & ~x168 & ~x171 & ~x198 & ~x228 & ~x229 & ~x231 & ~x232 & ~x234 & ~x253 & ~x254 & ~x283 & ~x285 & ~x287 & ~x291 & ~x311 & ~x315 & ~x318 & ~x334 & ~x339 & ~x344 & ~x362 & ~x363 & ~x367 & ~x371 & ~x393 & ~x398 & ~x401 & ~x419 & ~x426 & ~x454 & ~x478 & ~x483 & ~x484 & ~x507 & ~x508 & ~x509 & ~x510 & ~x512 & ~x531 & ~x534 & ~x538 & ~x539 & ~x747 & ~x759 & ~x760 & ~x774 & ~x783;
assign c9160 =  x294 & ~x11 & ~x160 & ~x169 & ~x173 & ~x196 & ~x604 & ~x723 & ~x760 & ~x778;
assign c9162 =  x300 &  x381 &  x385 &  x444 &  x494 &  x553 &  x582 & ~x45 & ~x50 & ~x56 & ~x102 & ~x186 & ~x369 & ~x777;
assign c9164 =  x304 &  x388 &  x501 & ~x241 & ~x345 & ~x745;
assign c9166 =  x246 &  x450 &  x518 & ~x29 & ~x199;
assign c9168 =  x614 & ~x242;
assign c9170 =  x506 &  x585 & ~x619 & ~x634 & ~x655 & ~x717 & ~x774;
assign c9172 = ~x87 & ~x92 & ~x168 & ~x193 & ~x206 & ~x292 & ~x403 & ~x515 & ~x538 & ~x540;
assign c9174 =  x379 &  x452 & ~x9 & ~x13 & ~x596 & ~x669 & ~x680 & ~x752;
assign c9176 =  x302 &  x507 &  x517 &  x608 &  x609 & ~x17 & ~x29 & ~x62 & ~x68 & ~x96 & ~x106 & ~x124 & ~x198 & ~x251 & ~x260 & ~x337 & ~x685 & ~x687 & ~x724 & ~x744 & ~x751 & ~x780;
assign c9178 =  x270 &  x351 &  x378 &  x379 &  x408 &  x409 &  x413 &  x414 &  x438 &  x492 &  x522 &  x547 &  x572 &  x600 &  x601 &  x648 &  x683 & ~x10 & ~x30 & ~x36 & ~x62 & ~x65 & ~x113 & ~x120 & ~x140 & ~x146 & ~x148 & ~x149 & ~x173 & ~x198 & ~x203 & ~x225 & ~x228 & ~x233 & ~x284 & ~x287 & ~x308 & ~x311 & ~x316 & ~x336 & ~x365 & ~x393 & ~x395 & ~x423 & ~x424 & ~x425 & ~x449 & ~x454 & ~x783;
assign c9180 = ~x443 & ~x444 & ~x455 & ~x515 & ~x539;
assign c9182 =  x277 &  x493 & ~x82 & ~x129 & ~x186 & ~x315 & ~x372 & ~x577;
assign c9184 =  x526 &  x609 &  x610 &  x613 & ~x4 & ~x8 & ~x66 & ~x70 & ~x141 & ~x208 & ~x425 & ~x447 & ~x726 & ~x731 & ~x767;
assign c9186 =  x580 & ~x0 & ~x1 & ~x2 & ~x9 & ~x10 & ~x30 & ~x34 & ~x36 & ~x38 & ~x42 & ~x57 & ~x58 & ~x63 & ~x64 & ~x84 & ~x92 & ~x94 & ~x111 & ~x114 & ~x117 & ~x118 & ~x124 & ~x140 & ~x149 & ~x176 & ~x179 & ~x180 & ~x200 & ~x203 & ~x205 & ~x227 & ~x229 & ~x232 & ~x233 & ~x234 & ~x252 & ~x254 & ~x259 & ~x262 & ~x279 & ~x282 & ~x286 & ~x289 & ~x291 & ~x309 & ~x335 & ~x337 & ~x340 & ~x342 & ~x343 & ~x363 & ~x365 & ~x368 & ~x372 & ~x373 & ~x374 & ~x393 & ~x397 & ~x420 & ~x422 & ~x424 & ~x426 & ~x448 & ~x455 & ~x484 & ~x485 & ~x772 & ~x783;
assign c9188 =  x350 &  x416 &  x488 &  x545 &  x591 & ~x8 & ~x36 & ~x64 & ~x65 & ~x66 & ~x92 & ~x94 & ~x113 & ~x117 & ~x139 & ~x149 & ~x169 & ~x173 & ~x176 & ~x200 & ~x203 & ~x227 & ~x252 & ~x258 & ~x287 & ~x339 & ~x393 & ~x397 & ~x660 & ~x700 & ~x717 & ~x742 & ~x772 & ~x773;
assign c9190 =  x405 &  x458 &  x521 &  x534 &  x561 & ~x4 & ~x11 & ~x17 & ~x30 & ~x38 & ~x67 & ~x86 & ~x144 & ~x146 & ~x171 & ~x177 & ~x201 & ~x280 & ~x371 & ~x693 & ~x717 & ~x744 & ~x755 & ~x757 & ~x762;
assign c9192 =  x249 &  x332 &  x410 &  x470 &  x494 & ~x60 & ~x62 & ~x146 & ~x399 & ~x633 & ~x741 & ~x749 & ~x760;
assign c9194 =  x271 &  x327 &  x354 & ~x3 & ~x7 & ~x9 & ~x10 & ~x11 & ~x12 & ~x23 & ~x24 & ~x25 & ~x26 & ~x27 & ~x28 & ~x29 & ~x30 & ~x34 & ~x35 & ~x49 & ~x53 & ~x55 & ~x57 & ~x61 & ~x62 & ~x63 & ~x80 & ~x84 & ~x85 & ~x90 & ~x91 & ~x93 & ~x114 & ~x118 & ~x120 & ~x123 & ~x143 & ~x149 & ~x169 & ~x172 & ~x173 & ~x176 & ~x179 & ~x198 & ~x200 & ~x205 & ~x206 & ~x207 & ~x223 & ~x225 & ~x226 & ~x227 & ~x228 & ~x229 & ~x231 & ~x233 & ~x253 & ~x256 & ~x258 & ~x261 & ~x264 & ~x280 & ~x283 & ~x285 & ~x288 & ~x289 & ~x291 & ~x308 & ~x314 & ~x315 & ~x317 & ~x337 & ~x339 & ~x341 & ~x346 & ~x363 & ~x367 & ~x369 & ~x372 & ~x374 & ~x392 & ~x395 & ~x398 & ~x401 & ~x420 & ~x421 & ~x422 & ~x423 & ~x424 & ~x428 & ~x429 & ~x448 & ~x453 & ~x454 & ~x455 & ~x456 & ~x699 & ~x727 & ~x729 & ~x757 & ~x760 & ~x775 & ~x776 & ~x783;
assign c9196 =  x560 &  x576;
assign c9198 = ~x12 & ~x28 & ~x29 & ~x33 & ~x36 & ~x44 & ~x48 & ~x65 & ~x66 & ~x69 & ~x77 & ~x82 & ~x110 & ~x117 & ~x122 & ~x138 & ~x142 & ~x143 & ~x144 & ~x179 & ~x180 & ~x196 & ~x202 & ~x203 & ~x208 & ~x223 & ~x225 & ~x232 & ~x259 & ~x261 & ~x263 & ~x281 & ~x283 & ~x284 & ~x285 & ~x289 & ~x309 & ~x312 & ~x313 & ~x314 & ~x317 & ~x318 & ~x339 & ~x343 & ~x346 & ~x369 & ~x397 & ~x398 & ~x400 & ~x401 & ~x402 & ~x419 & ~x423 & ~x425 & ~x426 & ~x427 & ~x451 & ~x453 & ~x454 & ~x455 & ~x456 & ~x457 & ~x482 & ~x483 & ~x484 & ~x537 & ~x587 & ~x759;
assign c9200 =  x160 &  x184 &  x211 &  x212 &  x267 &  x323 &  x324 &  x351 &  x352 &  x354 &  x358 &  x378 &  x379 &  x381 &  x382 &  x384 &  x385 &  x408 &  x410 &  x438 &  x441 &  x489 &  x490 &  x491 &  x494 &  x520 &  x599 &  x600 & ~x60 & ~x62 & ~x83 & ~x113 & ~x171 & ~x224 & ~x227 & ~x230 & ~x280 & ~x308 & ~x339 & ~x363 & ~x366 & ~x368 & ~x425 & ~x426 & ~x759 & ~x782 & ~x783;
assign c9202 =  x218 &  x220 &  x352 &  x358 &  x416 &  x548 &  x572 &  x573 & ~x2 & ~x7 & ~x8 & ~x9 & ~x10 & ~x13 & ~x14 & ~x16 & ~x17 & ~x21 & ~x22 & ~x25 & ~x26 & ~x31 & ~x34 & ~x37 & ~x38 & ~x40 & ~x41 & ~x50 & ~x53 & ~x54 & ~x56 & ~x59 & ~x60 & ~x61 & ~x62 & ~x66 & ~x67 & ~x83 & ~x86 & ~x87 & ~x88 & ~x90 & ~x91 & ~x112 & ~x114 & ~x115 & ~x117 & ~x118 & ~x119 & ~x120 & ~x122 & ~x139 & ~x142 & ~x143 & ~x144 & ~x145 & ~x149 & ~x167 & ~x198 & ~x199 & ~x200 & ~x202 & ~x224 & ~x225 & ~x226 & ~x227 & ~x228 & ~x230 & ~x252 & ~x255 & ~x281 & ~x284 & ~x308 & ~x310 & ~x313 & ~x336 & ~x338 & ~x340 & ~x364 & ~x366 & ~x367 & ~x393 & ~x448 & ~x476 & ~x701 & ~x729 & ~x732 & ~x733 & ~x755 & ~x756 & ~x757 & ~x761 & ~x763 & ~x764 & ~x773 & ~x774 & ~x776 & ~x779 & ~x782;
assign c9204 =  x248 &  x249 &  x376 &  x377 &  x520 &  x527 &  x545 & ~x65 & ~x130 & ~x168 & ~x341 & ~x392 & ~x644;
assign c9206 =  x248 &  x268 &  x325 &  x555 & ~x0 & ~x1 & ~x16 & ~x56 & ~x83 & ~x89 & ~x121 & ~x173 & ~x227 & ~x231 & ~x253 & ~x264 & ~x312 & ~x336 & ~x341 & ~x343 & ~x476 & ~x671 & ~x721 & ~x745 & ~x749 & ~x764;
assign c9208 =  x276 &  x350 &  x403 &  x405 &  x492 &  x541 &  x544 &  x545 & ~x229 & ~x233 & ~x255 & ~x426 & ~x606 & ~x746 & ~x759;
assign c9210 =  x444 &  x460 &  x473 &  x543 & ~x95 & ~x191 & ~x213 & ~x400;
assign c9212 =  x351 &  x356 &  x441 &  x469 &  x522 &  x527 & ~x28 & ~x36 & ~x37 & ~x54 & ~x62 & ~x65 & ~x92 & ~x226 & ~x234 & ~x262 & ~x335 & ~x342 & ~x344 & ~x365 & ~x368 & ~x393 & ~x394 & ~x401 & ~x426 & ~x428 & ~x635 & ~x691 & ~x720 & ~x745 & ~x771;
assign c9214 =  x435 &  x556 & ~x7 & ~x35 & ~x70 & ~x73 & ~x94 & ~x102 & ~x107 & ~x116 & ~x136 & ~x171 & ~x176 & ~x205 & ~x225 & ~x234 & ~x339 & ~x340 & ~x341 & ~x370 & ~x398 & ~x606 & ~x673 & ~x693 & ~x698 & ~x720 & ~x748;
assign c9216 =  x276 &  x328 &  x414 &  x435 &  x468 &  x493 &  x494 &  x495 &  x518 &  x655 & ~x0 & ~x4 & ~x5 & ~x11 & ~x17 & ~x24 & ~x26 & ~x28 & ~x31 & ~x35 & ~x37 & ~x56 & ~x57 & ~x60 & ~x63 & ~x65 & ~x67 & ~x88 & ~x91 & ~x92 & ~x112 & ~x115 & ~x139 & ~x141 & ~x144 & ~x145 & ~x146 & ~x150 & ~x168 & ~x196 & ~x198 & ~x200 & ~x224 & ~x225 & ~x226 & ~x228 & ~x229 & ~x233 & ~x252 & ~x254 & ~x258 & ~x259 & ~x281 & ~x282 & ~x284 & ~x288 & ~x310 & ~x312 & ~x313 & ~x316 & ~x317 & ~x335 & ~x336 & ~x343 & ~x364 & ~x365 & ~x367 & ~x392 & ~x394 & ~x420 & ~x448 & ~x476 & ~x729 & ~x746 & ~x758 & ~x760 & ~x770 & ~x771;
assign c9218 =  x472 &  x556 &  x571 & ~x28 & ~x44 & ~x54 & ~x56 & ~x59 & ~x94 & ~x100 & ~x140 & ~x150 & ~x151 & ~x159 & ~x186 & ~x235 & ~x262 & ~x395 & ~x399 & ~x674 & ~x699 & ~x783;
assign c9220 =  x463 &  x533 &  x538 &  x540 &  x565 & ~x39 & ~x279 & ~x621 & ~x632 & ~x726;
assign c9222 = ~x0 & ~x1 & ~x3 & ~x5 & ~x11 & ~x28 & ~x35 & ~x36 & ~x60 & ~x62 & ~x63 & ~x86 & ~x87 & ~x88 & ~x89 & ~x117 & ~x118 & ~x140 & ~x143 & ~x146 & ~x149 & ~x170 & ~x200 & ~x223 & ~x224 & ~x228 & ~x251 & ~x256 & ~x257 & ~x281 & ~x286 & ~x288 & ~x308 & ~x310 & ~x338 & ~x340 & ~x343 & ~x344 & ~x368 & ~x370 & ~x476 & ~x500 & ~x507 & ~x508 & ~x509 & ~x510 & ~x511 & ~x672 & ~x690 & ~x745 & ~x747 & ~x748 & ~x772 & ~x773 & ~x775;
assign c9224 = ~x319 & ~x377 & ~x453 & ~x455 & ~x485 & ~x513 & ~x515 & ~x538;
assign c9226 =  x324 &  x351 &  x354 &  x355 &  x379 &  x409 &  x436 &  x437 &  x466 &  x494 &  x522 &  x687 & ~x1 & ~x27 & ~x28 & ~x31 & ~x57 & ~x60 & ~x63 & ~x114 & ~x145 & ~x168 & ~x251 & ~x288 & ~x307 & ~x316 & ~x344 & ~x369 & ~x397 & ~x422 & ~x425 & ~x728 & ~x757 & ~x759 & ~x772;
assign c9228 =  x298 &  x377 &  x446 &  x467 & ~x574 & ~x595 & ~x675 & ~x773 & ~x775;
assign c9230 =  x277 &  x333 &  x468 &  x527 &  x558 & ~x1 & ~x6 & ~x369 & ~x605 & ~x682;
assign c9232 = ~x129 & ~x412;
assign c9234 = ~x41 & ~x45 & ~x47 & ~x72 & ~x74 & ~x75 & ~x88 & ~x100 & ~x110 & ~x135 & ~x141 & ~x145 & ~x167 & ~x176 & ~x183 & ~x199 & ~x260 & ~x290 & ~x319 & ~x343 & ~x372 & ~x373 & ~x399 & ~x421 & ~x448 & ~x452 & ~x455 & ~x672 & ~x708 & ~x714 & ~x718 & ~x747 & ~x750 & ~x753 & ~x754 & ~x781;
assign c9236 =  x472 &  x548 &  x583 & ~x1 & ~x4 & ~x6 & ~x7 & ~x8 & ~x28 & ~x29 & ~x34 & ~x61 & ~x64 & ~x84 & ~x86 & ~x96 & ~x140 & ~x141 & ~x176 & ~x204 & ~x232 & ~x256 & ~x257 & ~x279 & ~x281 & ~x285 & ~x288 & ~x292 & ~x314 & ~x319 & ~x335 & ~x337 & ~x339 & ~x340 & ~x373 & ~x374 & ~x396 & ~x398 & ~x422 & ~x426 & ~x449 & ~x455 & ~x456 & ~x717 & ~x749 & ~x751 & ~x758 & ~x767 & ~x774 & ~x775 & ~x780 & ~x781;
assign c9238 =  x266 &  x267 &  x325 &  x327 &  x331 &  x353 &  x360 &  x389 &  x431 &  x482 &  x490 & ~x12 & ~x21 & ~x27 & ~x40 & ~x66 & ~x87 & ~x111 & ~x115 & ~x169 & ~x258 & ~x314 & ~x365 & ~x730 & ~x757 & ~x765;
assign c9240 =  x403 &  x444 &  x462 & ~x184 & ~x281 & ~x345 & ~x534;
assign c9242 =  x74 &  x75 &  x185 &  x212 &  x213 &  x296 &  x324 &  x357 &  x381 &  x408 &  x409 &  x410 &  x436 &  x463 &  x469 &  x491 &  x494 &  x520 & ~x148 & ~x198 & ~x199 & ~x339 & ~x344 & ~x420 & ~x428;
assign c9244 =  x586 & ~x25 & ~x55 & ~x57 & ~x83 & ~x179 & ~x187 & ~x283 & ~x309 & ~x340 & ~x560 & ~x699 & ~x720 & ~x721;
assign c9246 = ~x8 & ~x28 & ~x44 & ~x46 & ~x56 & ~x68 & ~x69 & ~x70 & ~x86 & ~x87 & ~x114 & ~x117 & ~x122 & ~x124 & ~x129 & ~x142 & ~x146 & ~x168 & ~x171 & ~x177 & ~x200 & ~x207 & ~x234 & ~x283 & ~x290 & ~x307 & ~x337 & ~x339 & ~x363 & ~x391 & ~x394 & ~x399 & ~x403 & ~x425 & ~x537 & ~x538 & ~x539 & ~x700 & ~x701 & ~x732 & ~x733 & ~x744 & ~x771 & ~x778;
assign c9248 =  x276 &  x451 & ~x228 & ~x314 & ~x318 & ~x661 & ~x691;
assign c9250 =  x154 &  x240 &  x266 &  x269 &  x298 &  x321 &  x327 &  x354 &  x378 &  x381 &  x408 &  x411 &  x414 &  x432 &  x434 &  x462 &  x465 &  x490 & ~x11 & ~x30 & ~x90 & ~x91 & ~x112 & ~x118 & ~x141 & ~x197 & ~x339 & ~x700;
assign c9252 =  x300 &  x381 &  x443 &  x500 & ~x5 & ~x93 & ~x203 & ~x214 & ~x318 & ~x606;
assign c9254 =  x221 &  x462 &  x506 &  x544 & ~x45 & ~x92 & ~x117 & ~x143 & ~x199 & ~x705 & ~x713 & ~x722 & ~x765;
assign c9256 =  x132 &  x158 &  x159 &  x160 &  x182 &  x185 &  x214 &  x215 &  x326 &  x351 &  x414 &  x441 &  x545 &  x547 &  x548 &  x573 &  x601 & ~x366 & ~x367 & ~x393 & ~x453 & ~x454 & ~x455 & ~x476 & ~x482 & ~x757;
assign c9258 =  x190 &  x191 &  x269 &  x273 &  x301 &  x302 &  x331 &  x354 &  x357 &  x359 &  x409 &  x411 &  x412 &  x413 &  x415 &  x521 &  x572 &  x574 & ~x0 & ~x3 & ~x5 & ~x7 & ~x11 & ~x27 & ~x28 & ~x30 & ~x33 & ~x35 & ~x37 & ~x62 & ~x63 & ~x86 & ~x88 & ~x91 & ~x119 & ~x142 & ~x143 & ~x145 & ~x169 & ~x170 & ~x205 & ~x225 & ~x228 & ~x232 & ~x281 & ~x310 & ~x365 & ~x367 & ~x368 & ~x393 & ~x395 & ~x396 & ~x421 & ~x424 & ~x426 & ~x476 & ~x701 & ~x728 & ~x755 & ~x756 & ~x773;
assign c9260 =  x126 &  x155 &  x158 &  x211 &  x213 &  x215 &  x242 &  x244 &  x271 &  x324 &  x378 &  x381 &  x408 &  x463 &  x469 &  x677 &  x681;
assign c9262 = ~x3 & ~x6 & ~x9 & ~x16 & ~x18 & ~x27 & ~x30 & ~x34 & ~x42 & ~x44 & ~x56 & ~x62 & ~x65 & ~x88 & ~x118 & ~x122 & ~x124 & ~x141 & ~x143 & ~x151 & ~x153 & ~x169 & ~x177 & ~x225 & ~x227 & ~x229 & ~x232 & ~x254 & ~x258 & ~x260 & ~x261 & ~x263 & ~x279 & ~x281 & ~x284 & ~x285 & ~x291 & ~x308 & ~x313 & ~x318 & ~x335 & ~x337 & ~x341 & ~x349 & ~x363 & ~x394 & ~x395 & ~x427 & ~x429 & ~x454 & ~x455 & ~x484 & ~x509 & ~x510 & ~x746 & ~x756 & ~x771 & ~x774 & ~x777;
assign c9264 =  x321 &  x351 &  x358 &  x405 &  x432 &  x489 &  x491 &  x518 & ~x36 & ~x86 & ~x115 & ~x198 & ~x224 & ~x228 & ~x255 & ~x283 & ~x364 & ~x369 & ~x370 & ~x371 & ~x421 & ~x423 & ~x425 & ~x580 & ~x643 & ~x671 & ~x721 & ~x772;
assign c9266 =  x222 &  x383 &  x386 &  x411 &  x466 & ~x4 & ~x12 & ~x31 & ~x37 & ~x63 & ~x89 & ~x92 & ~x119 & ~x145 & ~x197 & ~x229 & ~x231 & ~x233 & ~x261 & ~x732 & ~x778 & ~x783;
assign c9268 =  x247 &  x248 &  x359 &  x414 &  x461 &  x520 &  x546 &  x571 &  x601 &  x602 &  x613 &  x626 & ~x0 & ~x2 & ~x4 & ~x7 & ~x9 & ~x11 & ~x24 & ~x26 & ~x28 & ~x34 & ~x35 & ~x37 & ~x38 & ~x58 & ~x59 & ~x60 & ~x64 & ~x83 & ~x85 & ~x89 & ~x91 & ~x92 & ~x93 & ~x94 & ~x115 & ~x116 & ~x117 & ~x119 & ~x120 & ~x148 & ~x150 & ~x168 & ~x170 & ~x205 & ~x226 & ~x227 & ~x229 & ~x254 & ~x257 & ~x279 & ~x280 & ~x282 & ~x308 & ~x311 & ~x314 & ~x336 & ~x337 & ~x338 & ~x339 & ~x343 & ~x365 & ~x366 & ~x367 & ~x369 & ~x392 & ~x394 & ~x425 & ~x427 & ~x758 & ~x759;
assign c9270 =  x351 &  x478 &  x491 &  x492 &  x539 & ~x111 & ~x142 & ~x182 & ~x215 & ~x340 & ~x371 & ~x392 & ~x677 & ~x736 & ~x772 & ~x776;
assign c9272 =  x215 &  x410 &  x492 &  x547 &  x548 &  x605 &  x631 &  x659 &  x678 &  x682 & ~x1 & ~x7 & ~x27 & ~x29 & ~x30 & ~x32 & ~x35 & ~x57 & ~x61 & ~x85 & ~x92 & ~x119 & ~x139 & ~x144 & ~x148 & ~x171 & ~x172 & ~x177 & ~x199 & ~x224 & ~x227 & ~x228 & ~x230 & ~x232 & ~x281 & ~x316 & ~x335 & ~x338 & ~x340 & ~x344 & ~x363 & ~x370 & ~x392 & ~x394 & ~x420 & ~x427 & ~x428 & ~x450 & ~x451 & ~x455 & ~x482 & ~x532 & ~x728 & ~x757 & ~x783;
assign c9274 =  x379 &  x576 &  x577 &  x583 &  x584 &  x601 &  x610 &  x612 & ~x5 & ~x10 & ~x37 & ~x65 & ~x83 & ~x90 & ~x92 & ~x111 & ~x119 & ~x121 & ~x123 & ~x124 & ~x147 & ~x173 & ~x208 & ~x224 & ~x225 & ~x230 & ~x233 & ~x255 & ~x307 & ~x308 & ~x367 & ~x394 & ~x430 & ~x447 & ~x449 & ~x476 & ~x771 & ~x774;
assign c9276 =  x133 &  x218 &  x243 &  x269 &  x296 &  x324 &  x351 &  x353 &  x358 &  x381 &  x386 &  x409 &  x434 &  x493 &  x573 &  x600 &  x601 & ~x5 & ~x9 & ~x10 & ~x11 & ~x32 & ~x34 & ~x35 & ~x36 & ~x55 & ~x60 & ~x112 & ~x115 & ~x140 & ~x141 & ~x143 & ~x149 & ~x224 & ~x225 & ~x252 & ~x255 & ~x310 & ~x340 & ~x364 & ~x366 & ~x367 & ~x371 & ~x393 & ~x395 & ~x421 & ~x447 & ~x448 & ~x700 & ~x727 & ~x774;
assign c9278 =  x351 &  x487 &  x507 &  x526 &  x535 & ~x56 & ~x125 & ~x178 & ~x234 & ~x283 & ~x371 & ~x393 & ~x559 & ~x620 & ~x633 & ~x699 & ~x707 & ~x711 & ~x728;
assign c9280 =  x462 &  x590 & ~x78 & ~x81 & ~x84 & ~x115 & ~x167 & ~x255 & ~x256 & ~x310 & ~x316 & ~x366 & ~x397 & ~x424 & ~x455 & ~x693 & ~x738 & ~x749 & ~x783;
assign c9282 =  x477 &  x543 & ~x124 & ~x399 & ~x760;
assign c9284 =  x299 &  x327 &  x356 & ~x26 & ~x28 & ~x29 & ~x34 & ~x48 & ~x50 & ~x62 & ~x74 & ~x92 & ~x100 & ~x114 & ~x151 & ~x179 & ~x201 & ~x230 & ~x252 & ~x254 & ~x256 & ~x510 & ~x674 & ~x675 & ~x713 & ~x726 & ~x757 & ~x761 & ~x770 & ~x773 & ~x774 & ~x780;
assign c9286 =  x461 &  x534 &  x547 &  x552 & ~x40 & ~x62 & ~x79 & ~x148 & ~x154 & ~x226 & ~x227 & ~x283 & ~x313 & ~x315 & ~x342 & ~x365 & ~x604 & ~x648 & ~x701 & ~x717 & ~x770;
assign c9288 =  x354 &  x384 & ~x23 & ~x33 & ~x36 & ~x93 & ~x118 & ~x119 & ~x125 & ~x176 & ~x318 & ~x369 & ~x447 & ~x454 & ~x455 & ~x671 & ~x726 & ~x727 & ~x748 & ~x781;
assign c9290 =  x381 &  x414 &  x439 &  x440 &  x462 &  x544 & ~x11 & ~x48 & ~x51 & ~x78 & ~x86 & ~x94 & ~x116 & ~x141 & ~x145 & ~x170 & ~x182 & ~x202 & ~x226 & ~x228 & ~x230 & ~x236 & ~x253 & ~x367 & ~x395 & ~x397 & ~x399 & ~x400 & ~x589 & ~x631 & ~x648 & ~x665 & ~x678 & ~x685 & ~x691 & ~x696 & ~x698 & ~x703 & ~x718 & ~x730 & ~x735 & ~x741 & ~x756 & ~x757 & ~x771 & ~x777 & ~x779;
assign c9292 =  x156 &  x211 &  x212 &  x218 &  x239 &  x240 &  x243 &  x244 &  x269 &  x272 &  x325 &  x329 &  x332 &  x380 &  x381 &  x383 &  x385 &  x407 &  x409 &  x410 &  x435 &  x437 &  x441 &  x463 &  x469 &  x489 &  x491 &  x547 &  x599;
assign c9294 =  x243 &  x271 &  x298 &  x299 &  x410 & ~x9 & ~x28 & ~x29 & ~x60 & ~x61 & ~x84 & ~x90 & ~x257 & ~x309 & ~x311 & ~x336 & ~x339 & ~x340 & ~x364 & ~x367 & ~x369 & ~x426 & ~x478 & ~x505 & ~x507 & ~x508 & ~x509 & ~x511 & ~x512 & ~x535 & ~x539 & ~x540 & ~x745 & ~x746 & ~x758 & ~x759;
assign c9296 =  x435 &  x436 &  x562 &  x619 &  x623 &  x625 &  x628 &  x629 & ~x2 & ~x9 & ~x10 & ~x13 & ~x29 & ~x41 & ~x57 & ~x59 & ~x60 & ~x64 & ~x143 & ~x168 & ~x199 & ~x205 & ~x224 & ~x225 & ~x226 & ~x227 & ~x229 & ~x253 & ~x258 & ~x337 & ~x340 & ~x341 & ~x368 & ~x370 & ~x392 & ~x426 & ~x476 & ~x700 & ~x734 & ~x767;
assign c9298 =  x461 &  x517 &  x563 &  x564 &  x593 &  x613 & ~x37 & ~x62 & ~x65 & ~x106 & ~x114 & ~x119 & ~x141 & ~x149 & ~x172 & ~x178 & ~x254 & ~x260 & ~x707 & ~x723 & ~x732 & ~x742 & ~x745 & ~x753;
assign c9300 =  x383 &  x543 &  x546 &  x553 &  x565 &  x570 & ~x24 & ~x119 & ~x142 & ~x173 & ~x200 & ~x204 & ~x205 & ~x234 & ~x283 & ~x339 & ~x362 & ~x755 & ~x756 & ~x778;
assign c9302 =  x274 &  x301 &  x331 &  x351 &  x357 &  x381 &  x386 &  x414 &  x494 &  x665 & ~x8 & ~x28 & ~x32 & ~x34 & ~x35 & ~x37 & ~x56 & ~x89 & ~x93 & ~x119 & ~x145 & ~x149 & ~x170 & ~x173 & ~x174 & ~x201 & ~x202 & ~x203 & ~x205 & ~x224 & ~x225 & ~x227 & ~x232 & ~x233 & ~x252 & ~x254 & ~x287 & ~x288 & ~x308 & ~x336 & ~x366 & ~x757 & ~x758 & ~x759;
assign c9304 =  x352 &  x411 &  x436 &  x437 &  x438 &  x478 &  x483 &  x501 & ~x7 & ~x70 & ~x80 & ~x99 & ~x101 & ~x102 & ~x119 & ~x120 & ~x135 & ~x139 & ~x178 & ~x208 & ~x265 & ~x279 & ~x307 & ~x372 & ~x623 & ~x645 & ~x727;
assign c9306 =  x387 &  x507 &  x599 &  x612 & ~x14 & ~x25 & ~x90 & ~x142 & ~x343 & ~x768 & ~x769;
assign c9308 =  x608 &  x612 & ~x3 & ~x20 & ~x83 & ~x121 & ~x122 & ~x141 & ~x153 & ~x174 & ~x228 & ~x262 & ~x363 & ~x392 & ~x419 & ~x648 & ~x690 & ~x731;
assign c9310 =  x221 &  x351 &  x353 &  x354 &  x356 &  x434 &  x445 & ~x0 & ~x2 & ~x14 & ~x36 & ~x37 & ~x49 & ~x51 & ~x61 & ~x85 & ~x89 & ~x91 & ~x98 & ~x110 & ~x121 & ~x122 & ~x143 & ~x148 & ~x149 & ~x168 & ~x170 & ~x172 & ~x197 & ~x198 & ~x202 & ~x223 & ~x227 & ~x229 & ~x310 & ~x315 & ~x338 & ~x340 & ~x343 & ~x364 & ~x369 & ~x701 & ~x722 & ~x730 & ~x748 & ~x750 & ~x762 & ~x778 & ~x780 & ~x783;
assign c9312 =  x265 &  x359 &  x375 &  x376 &  x405 &  x434 &  x460 &  x490 &  x491 &  x543 &  x570 & ~x31 & ~x56 & ~x143 & ~x308 & ~x315 & ~x344 & ~x364 & ~x718 & ~x747;
assign c9314 =  x351 &  x378 &  x379 &  x380 &  x381 &  x382 &  x407 &  x409 &  x461 &  x546 &  x573 &  x599 &  x600 &  x601 &  x626 &  x676 &  x677 &  x681 & ~x1 & ~x29 & ~x32 & ~x33 & ~x59 & ~x113 & ~x197 & ~x228 & ~x230 & ~x284 & ~x288 & ~x311 & ~x335 & ~x367 & ~x368 & ~x392 & ~x422 & ~x426 & ~x504 & ~x757 & ~x761;
assign c9316 = ~x6 & ~x10 & ~x70 & ~x91 & ~x170 & ~x173 & ~x174 & ~x179 & ~x197 & ~x198 & ~x238 & ~x335 & ~x372 & ~x392 & ~x395 & ~x398 & ~x419 & ~x479 & ~x487 & ~x511 & ~x538 & ~x539 & ~x773;
assign c9318 =  x694 & ~x29 & ~x64 & ~x170 & ~x231 & ~x258 & ~x363 & ~x371 & ~x391 & ~x425 & ~x540 & ~x566 & ~x567;
assign c9320 = ~x17 & ~x32 & ~x37 & ~x39 & ~x41 & ~x43 & ~x52 & ~x53 & ~x59 & ~x67 & ~x76 & ~x91 & ~x92 & ~x99 & ~x109 & ~x122 & ~x131 & ~x138 & ~x142 & ~x151 & ~x156 & ~x162 & ~x164 & ~x168 & ~x169 & ~x176 & ~x183 & ~x187 & ~x206 & ~x234 & ~x264 & ~x286 & ~x290 & ~x292 & ~x308 & ~x316 & ~x335 & ~x337 & ~x338 & ~x371 & ~x391 & ~x401 & ~x420 & ~x425 & ~x428 & ~x646 & ~x674 & ~x686 & ~x688 & ~x693 & ~x716 & ~x717 & ~x718 & ~x739 & ~x747 & ~x748 & ~x762 & ~x774 & ~x777 & ~x783;
assign c9322 = ~x20 & ~x29 & ~x33 & ~x36 & ~x40 & ~x46 & ~x48 & ~x55 & ~x59 & ~x71 & ~x72 & ~x76 & ~x80 & ~x84 & ~x96 & ~x116 & ~x145 & ~x146 & ~x180 & ~x197 & ~x206 & ~x253 & ~x257 & ~x282 & ~x283 & ~x287 & ~x307 & ~x310 & ~x311 & ~x335 & ~x363 & ~x391 & ~x396 & ~x420 & ~x421 & ~x480 & ~x481 & ~x487 & ~x511 & ~x732 & ~x743 & ~x782;
assign c9324 =  x212 &  x240 &  x352 &  x414 &  x438 & ~x1 & ~x27 & ~x34 & ~x56 & ~x59 & ~x64 & ~x86 & ~x142 & ~x144 & ~x149 & ~x176 & ~x203 & ~x205 & ~x224 & ~x229 & ~x251 & ~x254 & ~x256 & ~x260 & ~x283 & ~x285 & ~x288 & ~x334 & ~x338 & ~x344 & ~x367 & ~x368 & ~x371 & ~x395 & ~x396 & ~x400 & ~x448 & ~x587 & ~x756 & ~x760 & ~x774 & ~x775;
assign c9326 =  x468 &  x501 & ~x25 & ~x168 & ~x261 & ~x314 & ~x316 & ~x550 & ~x610 & ~x634 & ~x690 & ~x699 & ~x719 & ~x773;
assign c9328 =  x298 &  x302 &  x358 &  x437 & ~x39 & ~x174 & ~x180 & ~x213 & ~x215 & ~x284 & ~x338 & ~x604 & ~x631;
assign c9330 =  x218 &  x219 &  x247 &  x304 &  x351 &  x353 &  x379 &  x381 &  x382 &  x388 &  x409 &  x412 &  x445 &  x461 &  x462 &  x492 & ~x2 & ~x3 & ~x6 & ~x7 & ~x26 & ~x28 & ~x31 & ~x37 & ~x55 & ~x65 & ~x82 & ~x84 & ~x92 & ~x93 & ~x113 & ~x118 & ~x122 & ~x138 & ~x139 & ~x144 & ~x170 & ~x196 & ~x199 & ~x200 & ~x201 & ~x202 & ~x224 & ~x229 & ~x230 & ~x261 & ~x287 & ~x310 & ~x311 & ~x337 & ~x338 & ~x344 & ~x366 & ~x420 & ~x448 & ~x476 & ~x728 & ~x767 & ~x772 & ~x773 & ~x775 & ~x776;
assign c9332 =  x380 &  x585 & ~x15 & ~x83 & ~x180 & ~x202 & ~x606 & ~x688;
assign c9334 =  x273 &  x329 &  x405 &  x408 &  x440 &  x490 & ~x175 & ~x181 & ~x253 & ~x260 & ~x559 & ~x630 & ~x650 & ~x656 & ~x696 & ~x707 & ~x783;
assign c9336 =  x219 &  x406 &  x435 &  x490 &  x521 &  x546 &  x547 &  x574 &  x584 &  x598 & ~x5 & ~x6 & ~x8 & ~x21 & ~x25 & ~x27 & ~x29 & ~x32 & ~x36 & ~x47 & ~x49 & ~x57 & ~x65 & ~x87 & ~x90 & ~x91 & ~x93 & ~x94 & ~x106 & ~x117 & ~x139 & ~x140 & ~x141 & ~x144 & ~x145 & ~x148 & ~x168 & ~x169 & ~x172 & ~x175 & ~x177 & ~x202 & ~x225 & ~x226 & ~x228 & ~x254 & ~x255 & ~x256 & ~x281 & ~x282 & ~x285 & ~x309 & ~x310 & ~x311 & ~x312 & ~x336 & ~x338 & ~x368 & ~x720 & ~x721 & ~x731 & ~x738 & ~x744 & ~x745 & ~x747 & ~x756 & ~x763 & ~x764 & ~x775 & ~x778;
assign c9338 =  x636 & ~x3 & ~x9 & ~x26 & ~x28 & ~x29 & ~x30 & ~x37 & ~x38 & ~x57 & ~x63 & ~x65 & ~x83 & ~x89 & ~x91 & ~x95 & ~x122 & ~x142 & ~x145 & ~x147 & ~x151 & ~x170 & ~x171 & ~x172 & ~x178 & ~x179 & ~x203 & ~x205 & ~x228 & ~x230 & ~x234 & ~x255 & ~x256 & ~x258 & ~x260 & ~x261 & ~x263 & ~x281 & ~x282 & ~x285 & ~x287 & ~x288 & ~x289 & ~x291 & ~x307 & ~x308 & ~x309 & ~x313 & ~x314 & ~x319 & ~x335 & ~x341 & ~x343 & ~x345 & ~x363 & ~x364 & ~x367 & ~x370 & ~x371 & ~x372 & ~x374 & ~x391 & ~x395 & ~x396 & ~x399 & ~x402 & ~x419 & ~x421 & ~x423 & ~x424 & ~x425 & ~x453 & ~x454 & ~x455 & ~x456 & ~x457 & ~x479 & ~x480 & ~x481 & ~x483 & ~x729;
assign c9340 =  x301 &  x303 &  x357 & ~x281;
assign c9342 =  x245 &  x267 &  x331 &  x348 &  x375 &  x501 &  x518 & ~x8 & ~x337 & ~x643 & ~x711;
assign c9344 =  x211 &  x238 &  x275 &  x321 &  x330 &  x349 &  x350 &  x358 &  x416 &  x444 &  x445 &  x471 &  x518 &  x527 &  x529 &  x583 & ~x6 & ~x14 & ~x26 & ~x27 & ~x29 & ~x31 & ~x60 & ~x84 & ~x87 & ~x91 & ~x111 & ~x112 & ~x117 & ~x119 & ~x148 & ~x172 & ~x174 & ~x230 & ~x252 & ~x258 & ~x311 & ~x314 & ~x366 & ~x368 & ~x755 & ~x756 & ~x783;
assign c9346 =  x694 & ~x0 & ~x2 & ~x3 & ~x8 & ~x28 & ~x31 & ~x32 & ~x33 & ~x35 & ~x36 & ~x37 & ~x55 & ~x56 & ~x57 & ~x61 & ~x62 & ~x86 & ~x87 & ~x88 & ~x89 & ~x90 & ~x91 & ~x92 & ~x93 & ~x111 & ~x114 & ~x116 & ~x117 & ~x118 & ~x119 & ~x120 & ~x121 & ~x140 & ~x141 & ~x171 & ~x199 & ~x232 & ~x233 & ~x253 & ~x255 & ~x256 & ~x257 & ~x258 & ~x259 & ~x260 & ~x280 & ~x281 & ~x282 & ~x283 & ~x284 & ~x286 & ~x288 & ~x307 & ~x308 & ~x309 & ~x315 & ~x316 & ~x334 & ~x336 & ~x342 & ~x343 & ~x344 & ~x362 & ~x363 & ~x368 & ~x372 & ~x390 & ~x392 & ~x393 & ~x396 & ~x419 & ~x421 & ~x422 & ~x424 & ~x425 & ~x426 & ~x427 & ~x447 & ~x448 & ~x452 & ~x456 & ~x475 & ~x476 & ~x478 & ~x481 & ~x503 & ~x511 & ~x531 & ~x559 & ~x759;
assign c9348 =  x184 &  x212 &  x242 &  x243 &  x247 &  x269 &  x301 &  x407 &  x413 &  x435 &  x436 &  x441 &  x464 &  x467 &  x492 &  x497 &  x520 &  x522 &  x637 & ~x2 & ~x8 & ~x11 & ~x26 & ~x27 & ~x29 & ~x34 & ~x62 & ~x65 & ~x85 & ~x86 & ~x94 & ~x111 & ~x115 & ~x144 & ~x146 & ~x149 & ~x173 & ~x175 & ~x176 & ~x196 & ~x200 & ~x224 & ~x226 & ~x229 & ~x232 & ~x254 & ~x255 & ~x308 & ~x313 & ~x392 & ~x420 & ~x422 & ~x756 & ~x759 & ~x783;
assign c9350 =  x386 &  x466 &  x552 & ~x8 & ~x35 & ~x114 & ~x231 & ~x233 & ~x252 & ~x287 & ~x308 & ~x315 & ~x342 & ~x369 & ~x400 & ~x401 & ~x606 & ~x731 & ~x762;
assign c9352 =  x159 &  x160 &  x186 &  x241 &  x270 &  x272 &  x296 &  x324 &  x325 &  x328 &  x359 &  x379 &  x381 &  x384 &  x385 &  x387 &  x410 &  x469 &  x599 &  x600 & ~x7 & ~x55 & ~x60 & ~x91 & ~x111 & ~x113 & ~x115 & ~x116 & ~x145 & ~x167 & ~x170 & ~x224 & ~x257 & ~x281 & ~x285 & ~x311 & ~x312 & ~x313 & ~x337 & ~x338 & ~x340 & ~x342 & ~x368 & ~x369 & ~x397 & ~x398;
assign c9354 =  x328 &  x353 &  x358 &  x376 &  x489 &  x494 &  x626 & ~x32 & ~x59 & ~x256 & ~x338;
assign c9356 =  x215 &  x245 &  x295 &  x416 &  x516 &  x543 &  x545 &  x602 &  x603 &  x625 & ~x6 & ~x8 & ~x10 & ~x27 & ~x29 & ~x34 & ~x57 & ~x61 & ~x85 & ~x87 & ~x112 & ~x114 & ~x115 & ~x117 & ~x118 & ~x119 & ~x120 & ~x168 & ~x196 & ~x197 & ~x199 & ~x223 & ~x224 & ~x225 & ~x226 & ~x227 & ~x232 & ~x253 & ~x282 & ~x286 & ~x309 & ~x310 & ~x311 & ~x316 & ~x336 & ~x337 & ~x340 & ~x341 & ~x364 & ~x372 & ~x393 & ~x394 & ~x397 & ~x420 & ~x447 & ~x475 & ~x476 & ~x755 & ~x756 & ~x757 & ~x758 & ~x760 & ~x776 & ~x783;
assign c9358 = ~x2 & ~x31 & ~x33 & ~x42 & ~x56 & ~x84 & ~x93 & ~x94 & ~x101 & ~x107 & ~x115 & ~x136 & ~x141 & ~x158 & ~x163 & ~x263 & ~x309 & ~x340 & ~x455 & ~x457 & ~x744 & ~x783;
assign c9360 =  x463 &  x543 &  x612 & ~x2 & ~x8 & ~x19 & ~x28 & ~x35 & ~x49 & ~x53 & ~x56 & ~x58 & ~x60 & ~x61 & ~x63 & ~x65 & ~x66 & ~x74 & ~x111 & ~x114 & ~x117 & ~x146 & ~x150 & ~x178 & ~x255 & ~x256 & ~x283 & ~x308 & ~x371 & ~x476 & ~x644 & ~x685 & ~x687 & ~x692 & ~x701 & ~x715 & ~x726 & ~x733 & ~x734 & ~x737 & ~x751 & ~x756 & ~x761 & ~x764 & ~x772;
assign c9362 =  x326 & ~x6 & ~x28 & ~x31 & ~x40 & ~x52 & ~x57 & ~x58 & ~x64 & ~x86 & ~x95 & ~x115 & ~x118 & ~x119 & ~x151 & ~x169 & ~x170 & ~x174 & ~x175 & ~x176 & ~x203 & ~x206 & ~x226 & ~x228 & ~x234 & ~x257 & ~x308 & ~x313 & ~x315 & ~x336 & ~x340 & ~x395 & ~x420 & ~x505 & ~x506 & ~x507 & ~x564 & ~x566 & ~x567 & ~x596 & ~x643 & ~x672 & ~x744 & ~x745 & ~x760 & ~x775 & ~x776;
assign c9364 = ~x4 & ~x26 & ~x37 & ~x44 & ~x52 & ~x55 & ~x59 & ~x67 & ~x79 & ~x84 & ~x94 & ~x95 & ~x97 & ~x114 & ~x124 & ~x132 & ~x140 & ~x164 & ~x199 & ~x201 & ~x205 & ~x207 & ~x210 & ~x225 & ~x226 & ~x232 & ~x258 & ~x285 & ~x289 & ~x291 & ~x292 & ~x307 & ~x366 & ~x374 & ~x419 & ~x422 & ~x429 & ~x448 & ~x700 & ~x756 & ~x770;
assign c9366 =  x409 &  x538 & ~x13 & ~x19 & ~x85 & ~x86 & ~x122 & ~x138 & ~x179 & ~x187 & ~x203 & ~x287 & ~x290 & ~x367 & ~x400 & ~x697 & ~x712 & ~x730 & ~x771 & ~x778;
assign c9368 =  x328 &  x377 &  x472 &  x583 & ~x49 & ~x68 & ~x127 & ~x173 & ~x253 & ~x724;
assign c9370 =  x238 &  x275 &  x330 &  x386 &  x518 &  x519 &  x546 &  x552 &  x583 &  x585 & ~x2 & ~x8 & ~x10 & ~x19 & ~x27 & ~x58 & ~x59 & ~x61 & ~x89 & ~x91 & ~x113 & ~x115 & ~x119 & ~x120 & ~x123 & ~x140 & ~x168 & ~x171 & ~x177 & ~x206 & ~x225 & ~x254 & ~x257 & ~x336 & ~x339 & ~x342 & ~x368 & ~x369 & ~x747 & ~x772;
assign c9372 =  x103 &  x128 &  x155 &  x159 &  x183 &  x184 &  x212 &  x213 &  x240 &  x268 &  x269 &  x296 &  x297 &  x325 &  x357 &  x407 &  x408 &  x435 &  x463 &  x464 &  x497 &  x520 & ~x33 & ~x62 & ~x84 & ~x91 & ~x92 & ~x117 & ~x233 & ~x257 & ~x259 & ~x309 & ~x316 & ~x342 & ~x364 & ~x759;
assign c9374 =  x321 &  x467 &  x520 & ~x10 & ~x23 & ~x28 & ~x35 & ~x44 & ~x168 & ~x181 & ~x186 & ~x198 & ~x204 & ~x228 & ~x234 & ~x252 & ~x285 & ~x368 & ~x398 & ~x671 & ~x691 & ~x699 & ~x728 & ~x741 & ~x753 & ~x778;
assign c9376 = ~x17 & ~x28 & ~x86 & ~x114 & ~x136 & ~x178 & ~x180 & ~x182 & ~x225 & ~x309 & ~x338 & ~x358 & ~x360 & ~x426 & ~x776;
assign c9378 =  x249 &  x414 &  x586 &  x604 &  x614 &  x641 &  x642 &  x656 & ~x6 & ~x8 & ~x12 & ~x84 & ~x87 & ~x119 & ~x206 & ~x229 & ~x286 & ~x308 & ~x420 & ~x426 & ~x427 & ~x728 & ~x757 & ~x758;
assign c9380 = ~x0 & ~x1 & ~x5 & ~x8 & ~x11 & ~x14 & ~x24 & ~x26 & ~x27 & ~x30 & ~x35 & ~x36 & ~x37 & ~x42 & ~x53 & ~x54 & ~x56 & ~x59 & ~x60 & ~x61 & ~x63 & ~x64 & ~x70 & ~x76 & ~x82 & ~x86 & ~x87 & ~x93 & ~x94 & ~x96 & ~x97 & ~x111 & ~x112 & ~x114 & ~x121 & ~x143 & ~x148 & ~x150 & ~x152 & ~x172 & ~x173 & ~x176 & ~x178 & ~x179 & ~x180 & ~x196 & ~x197 & ~x199 & ~x201 & ~x204 & ~x205 & ~x207 & ~x225 & ~x229 & ~x231 & ~x233 & ~x235 & ~x236 & ~x251 & ~x254 & ~x257 & ~x259 & ~x260 & ~x261 & ~x280 & ~x283 & ~x285 & ~x291 & ~x314 & ~x319 & ~x335 & ~x336 & ~x337 & ~x343 & ~x344 & ~x345 & ~x363 & ~x365 & ~x366 & ~x367 & ~x391 & ~x392 & ~x396 & ~x400 & ~x401 & ~x420 & ~x422 & ~x426 & ~x428 & ~x448 & ~x449 & ~x455 & ~x482 & ~x483 & ~x484 & ~x531 & ~x644 & ~x746 & ~x758 & ~x770 & ~x773 & ~x775;
assign c9382 =  x273 &  x274 &  x275 &  x293 &  x333 &  x360 &  x413 &  x432 &  x433 &  x445 & ~x24 & ~x116 & ~x141 & ~x176 & ~x203 & ~x260 & ~x285 & ~x369 & ~x608;
assign c9384 =  x604 & ~x4 & ~x6 & ~x7 & ~x10 & ~x16 & ~x32 & ~x35 & ~x52 & ~x54 & ~x64 & ~x68 & ~x69 & ~x73 & ~x74 & ~x75 & ~x83 & ~x85 & ~x90 & ~x102 & ~x104 & ~x115 & ~x140 & ~x146 & ~x147 & ~x152 & ~x153 & ~x179 & ~x180 & ~x225 & ~x228 & ~x254 & ~x261 & ~x280 & ~x291 & ~x312 & ~x336 & ~x368 & ~x479 & ~x510 & ~x512 & ~x702 & ~x728 & ~x742 & ~x747 & ~x768 & ~x772 & ~x773 & ~x774;
assign c9386 =  x294 &  x302 &  x349 &  x350 &  x379 &  x389 &  x426 &  x488 & ~x47 & ~x49 & ~x77 & ~x115 & ~x252 & ~x258 & ~x279 & ~x289 & ~x728 & ~x748 & ~x773;
assign c9388 =  x299 &  x301 &  x302 &  x327 &  x329 &  x332 &  x384 &  x386 &  x407 &  x408 &  x411 &  x413 &  x434 &  x437 &  x466 &  x467 &  x493 &  x494 &  x519 &  x520 &  x653 &  x654 & ~x1 & ~x2 & ~x4 & ~x6 & ~x8 & ~x29 & ~x31 & ~x55 & ~x60 & ~x61 & ~x64 & ~x85 & ~x86 & ~x88 & ~x92 & ~x112 & ~x117 & ~x118 & ~x121 & ~x141 & ~x142 & ~x143 & ~x144 & ~x145 & ~x168 & ~x199 & ~x224 & ~x225 & ~x227 & ~x229 & ~x251 & ~x253 & ~x254 & ~x255 & ~x256 & ~x288 & ~x310 & ~x313 & ~x314 & ~x315 & ~x316 & ~x336 & ~x338 & ~x364 & ~x370 & ~x371 & ~x393 & ~x397 & ~x398 & ~x421 & ~x427 & ~x729 & ~x756;
assign c9390 =  x303 &  x409 &  x436 &  x440 &  x460 &  x473 & ~x16 & ~x76 & ~x97 & ~x110 & ~x116 & ~x145 & ~x154 & ~x176 & ~x178 & ~x205 & ~x262 & ~x341 & ~x420 & ~x602 & ~x603 & ~x604 & ~x605 & ~x635 & ~x640 & ~x651 & ~x657 & ~x666 & ~x679 & ~x681 & ~x683 & ~x700 & ~x712 & ~x760 & ~x768;
assign c9392 =  x638 & ~x2 & ~x37 & ~x61 & ~x95 & ~x105 & ~x116 & ~x121 & ~x133 & ~x229 & ~x279 & ~x307 & ~x309 & ~x310 & ~x316 & ~x336 & ~x338 & ~x346 & ~x362 & ~x391 & ~x394 & ~x419 & ~x424 & ~x451 & ~x730 & ~x767 & ~x771;
assign c9394 =  x421 &  x443 & ~x161 & ~x686;
assign c9396 = ~x26 & ~x29 & ~x34 & ~x37 & ~x44 & ~x52 & ~x58 & ~x66 & ~x94 & ~x96 & ~x98 & ~x99 & ~x105 & ~x107 & ~x112 & ~x139 & ~x145 & ~x148 & ~x149 & ~x162 & ~x164 & ~x165 & ~x176 & ~x180 & ~x190 & ~x195 & ~x196 & ~x197 & ~x225 & ~x234 & ~x254 & ~x307 & ~x319 & ~x335 & ~x336 & ~x341 & ~x359 & ~x363 & ~x393 & ~x398 & ~x399 & ~x424 & ~x744 & ~x746 & ~x756 & ~x776;
assign c9398 = ~x54 & ~x68 & ~x180 & ~x291 & ~x319 & ~x401 & ~x419 & ~x425 & ~x460 & ~x482 & ~x510 & ~x511 & ~x512 & ~x690 & ~x745 & ~x770;
assign c9400 =  x580 &  x582 & ~x31 & ~x32 & ~x40 & ~x42 & ~x73 & ~x105 & ~x125 & ~x136 & ~x178 & ~x179 & ~x200 & ~x202 & ~x206 & ~x225 & ~x226 & ~x285 & ~x370 & ~x428 & ~x631 & ~x646 & ~x681 & ~x683 & ~x690 & ~x693 & ~x721 & ~x727 & ~x728 & ~x731 & ~x733 & ~x773 & ~x776 & ~x779;
assign c9402 =  x705 & ~x334 & ~x446 & ~x511;
assign c9404 = ~x3 & ~x4 & ~x5 & ~x8 & ~x10 & ~x11 & ~x12 & ~x16 & ~x27 & ~x29 & ~x30 & ~x32 & ~x33 & ~x34 & ~x35 & ~x36 & ~x38 & ~x40 & ~x42 & ~x48 & ~x49 & ~x50 & ~x54 & ~x57 & ~x59 & ~x60 & ~x62 & ~x63 & ~x65 & ~x66 & ~x67 & ~x68 & ~x69 & ~x83 & ~x89 & ~x91 & ~x93 & ~x94 & ~x95 & ~x110 & ~x111 & ~x112 & ~x115 & ~x118 & ~x121 & ~x122 & ~x123 & ~x124 & ~x140 & ~x142 & ~x143 & ~x145 & ~x150 & ~x151 & ~x153 & ~x168 & ~x169 & ~x170 & ~x171 & ~x173 & ~x176 & ~x177 & ~x179 & ~x195 & ~x196 & ~x197 & ~x198 & ~x199 & ~x201 & ~x202 & ~x203 & ~x205 & ~x206 & ~x208 & ~x230 & ~x231 & ~x233 & ~x236 & ~x251 & ~x252 & ~x253 & ~x255 & ~x260 & ~x262 & ~x263 & ~x283 & ~x286 & ~x287 & ~x289 & ~x291 & ~x307 & ~x309 & ~x312 & ~x313 & ~x314 & ~x315 & ~x319 & ~x335 & ~x337 & ~x339 & ~x343 & ~x344 & ~x363 & ~x364 & ~x365 & ~x368 & ~x370 & ~x373 & ~x374 & ~x391 & ~x392 & ~x393 & ~x395 & ~x397 & ~x399 & ~x400 & ~x420 & ~x421 & ~x423 & ~x427 & ~x428 & ~x429 & ~x448 & ~x449 & ~x451 & ~x454 & ~x455 & ~x457 & ~x477 & ~x478 & ~x482 & ~x483 & ~x484 & ~x727 & ~x729 & ~x746 & ~x747 & ~x756 & ~x757 & ~x758 & ~x759 & ~x763 & ~x773 & ~x775;
assign c9406 =  x212 &  x245 &  x248 &  x269 &  x472 & ~x64 & ~x67 & ~x139 & ~x146 & ~x339 & ~x393 & ~x617 & ~x654;
assign c9408 =  x306 &  x331 &  x547 &  x571 & ~x20 & ~x43 & ~x140 & ~x204 & ~x279 & ~x341 & ~x365 & ~x713 & ~x726 & ~x765 & ~x766;
assign c9410 =  x266 &  x268 &  x301 &  x303 &  x406 &  x459 &  x489 & ~x23 & ~x138 & ~x142 & ~x148 & ~x168 & ~x312 & ~x314 & ~x336 & ~x691 & ~x766;
assign c9412 =  x272 &  x681 & ~x458;
assign c9414 =  x580 & ~x0 & ~x1 & ~x2 & ~x3 & ~x4 & ~x5 & ~x8 & ~x10 & ~x23 & ~x24 & ~x27 & ~x28 & ~x29 & ~x31 & ~x32 & ~x36 & ~x37 & ~x38 & ~x39 & ~x53 & ~x55 & ~x59 & ~x60 & ~x61 & ~x62 & ~x64 & ~x65 & ~x85 & ~x86 & ~x87 & ~x89 & ~x92 & ~x93 & ~x94 & ~x96 & ~x112 & ~x113 & ~x114 & ~x117 & ~x119 & ~x121 & ~x123 & ~x143 & ~x145 & ~x147 & ~x149 & ~x170 & ~x171 & ~x172 & ~x174 & ~x175 & ~x177 & ~x178 & ~x179 & ~x195 & ~x196 & ~x197 & ~x198 & ~x199 & ~x200 & ~x202 & ~x223 & ~x224 & ~x225 & ~x227 & ~x229 & ~x230 & ~x232 & ~x234 & ~x253 & ~x254 & ~x255 & ~x256 & ~x258 & ~x261 & ~x262 & ~x263 & ~x280 & ~x281 & ~x286 & ~x287 & ~x289 & ~x290 & ~x291 & ~x308 & ~x310 & ~x311 & ~x315 & ~x316 & ~x319 & ~x336 & ~x339 & ~x344 & ~x346 & ~x364 & ~x365 & ~x368 & ~x369 & ~x372 & ~x374 & ~x392 & ~x395 & ~x396 & ~x397 & ~x398 & ~x401 & ~x419 & ~x420 & ~x421 & ~x422 & ~x423 & ~x424 & ~x425 & ~x426 & ~x427 & ~x428 & ~x429 & ~x447 & ~x448 & ~x455 & ~x484 & ~x727 & ~x729 & ~x756 & ~x757 & ~x758 & ~x759;
assign c9416 =  x187 &  x215 &  x216 &  x243 &  x354 &  x410 &  x438 &  x601 & ~x0 & ~x4 & ~x5 & ~x9 & ~x31 & ~x34 & ~x35 & ~x59 & ~x60 & ~x61 & ~x64 & ~x85 & ~x88 & ~x111 & ~x112 & ~x114 & ~x116 & ~x118 & ~x143 & ~x149 & ~x197 & ~x198 & ~x251 & ~x252 & ~x253 & ~x256 & ~x259 & ~x279 & ~x308 & ~x311 & ~x336 & ~x338 & ~x340 & ~x342 & ~x364 & ~x365 & ~x366 & ~x370 & ~x372 & ~x394 & ~x395 & ~x399 & ~x400 & ~x425 & ~x426 & ~x427 & ~x428 & ~x453 & ~x454 & ~x455 & ~x456 & ~x477 & ~x478 & ~x480 & ~x481 & ~x482 & ~x483 & ~x505 & ~x509 & ~x510 & ~x511 & ~x538 & ~x539 & ~x757 & ~x759 & ~x772 & ~x773;
assign c9418 =  x249 &  x270 &  x295 &  x356 &  x493 &  x518 & ~x36 & ~x42 & ~x113 & ~x120 & ~x223 & ~x225 & ~x226 & ~x258 & ~x338 & ~x341 & ~x365 & ~x659 & ~x663 & ~x699 & ~x731 & ~x736 & ~x758 & ~x761 & ~x764 & ~x783;
assign c9420 =  x183 &  x211 &  x212 &  x241 &  x242 &  x273 &  x276 &  x295 &  x301 &  x302 &  x328 &  x330 &  x332 &  x382 &  x387 &  x520 &  x527 & ~x7 & ~x27 & ~x28 & ~x33 & ~x61 & ~x62 & ~x83 & ~x114 & ~x116 & ~x117 & ~x118 & ~x140 & ~x141 & ~x145 & ~x168 & ~x169 & ~x197 & ~x198 & ~x224 & ~x228 & ~x252 & ~x255 & ~x256 & ~x257 & ~x281 & ~x314 & ~x336 & ~x364 & ~x365 & ~x366 & ~x367 & ~x419 & ~x757 & ~x760 & ~x783;
assign c9422 = ~x0 & ~x5 & ~x7 & ~x8 & ~x10 & ~x24 & ~x27 & ~x29 & ~x30 & ~x37 & ~x38 & ~x39 & ~x57 & ~x60 & ~x62 & ~x65 & ~x66 & ~x84 & ~x88 & ~x90 & ~x95 & ~x113 & ~x114 & ~x115 & ~x116 & ~x135 & ~x140 & ~x141 & ~x147 & ~x150 & ~x170 & ~x225 & ~x229 & ~x256 & ~x258 & ~x281 & ~x284 & ~x290 & ~x311 & ~x317 & ~x344 & ~x345 & ~x362 & ~x365 & ~x373 & ~x374 & ~x390 & ~x393 & ~x395 & ~x396 & ~x397 & ~x398 & ~x419 & ~x421 & ~x424 & ~x448 & ~x504 & ~x587 & ~x729 & ~x745 & ~x758 & ~x759;
assign c9424 =  x238 &  x376 &  x480 & ~x77 & ~x122 & ~x226;
assign c9426 =  x554 & ~x9 & ~x370 & ~x562 & ~x578 & ~x603 & ~x623 & ~x624 & ~x666 & ~x712;
assign c9428 =  x221 &  x488 &  x516 & ~x9 & ~x27 & ~x34 & ~x46 & ~x77 & ~x99 & ~x100 & ~x117 & ~x175 & ~x308 & ~x672 & ~x673 & ~x690 & ~x701 & ~x714 & ~x745;
assign c9430 =  x418 &  x538 &  x540 & ~x7 & ~x33 & ~x345 & ~x364 & ~x392 & ~x578 & ~x653;
assign c9432 =  x715 &  x735 &  x742;
assign c9434 =  x386 &  x387 &  x388 &  x473 &  x553 & ~x13 & ~x49 & ~x309 & ~x372 & ~x603 & ~x655;
assign c9436 =  x266 &  x302 &  x305 &  x356 &  x437 &  x463 &  x466 & ~x19 & ~x108 & ~x145 & ~x146 & ~x173 & ~x175 & ~x233 & ~x782;
assign c9438 = ~x31 & ~x37 & ~x83 & ~x117 & ~x118 & ~x121 & ~x142 & ~x169 & ~x253 & ~x265 & ~x394 & ~x400 & ~x424 & ~x426 & ~x429 & ~x454 & ~x455 & ~x457 & ~x475 & ~x482 & ~x483 & ~x484 & ~x487 & ~x509 & ~x510 & ~x537 & ~x538 & ~x539 & ~x587;
assign c9440 =  x127 &  x155 &  x156 &  x158 &  x184 &  x185 &  x211 &  x212 &  x213 &  x239 &  x242 &  x243 &  x269 &  x270 &  x351 &  x379 &  x381 &  x407 &  x410 &  x435 &  x465 &  x469 &  x493 &  x545 &  x574 &  x656 &  x683 & ~x2 & ~x9 & ~x27 & ~x34 & ~x139 & ~x144 & ~x223 & ~x283 & ~x288 & ~x316 & ~x339 & ~x368 & ~x394 & ~x397 & ~x399 & ~x423 & ~x453 & ~x756;
assign c9442 = ~x2 & ~x5 & ~x15 & ~x36 & ~x39 & ~x41 & ~x42 & ~x67 & ~x73 & ~x88 & ~x91 & ~x124 & ~x151 & ~x179 & ~x180 & ~x200 & ~x206 & ~x208 & ~x223 & ~x225 & ~x232 & ~x239 & ~x262 & ~x280 & ~x290 & ~x316 & ~x317 & ~x344 & ~x345 & ~x363 & ~x368 & ~x369 & ~x372 & ~x391 & ~x420 & ~x422 & ~x423 & ~x428 & ~x560 & ~x731 & ~x732 & ~x733 & ~x742 & ~x745 & ~x748 & ~x750 & ~x760 & ~x782;
assign c9444 =  x192 &  x217 &  x218 &  x246 &  x247 &  x248 &  x270 &  x274 &  x275 &  x304 &  x330 &  x357 &  x358 &  x386 &  x408 &  x409 &  x411 &  x435 &  x438 &  x490 &  x491 &  x492 &  x493 & ~x0 & ~x5 & ~x7 & ~x9 & ~x12 & ~x26 & ~x30 & ~x31 & ~x32 & ~x33 & ~x34 & ~x56 & ~x57 & ~x58 & ~x60 & ~x62 & ~x63 & ~x65 & ~x66 & ~x67 & ~x87 & ~x89 & ~x93 & ~x113 & ~x115 & ~x119 & ~x141 & ~x143 & ~x146 & ~x169 & ~x170 & ~x172 & ~x197 & ~x198 & ~x199 & ~x227 & ~x230 & ~x252 & ~x253 & ~x254 & ~x256 & ~x258 & ~x259 & ~x282 & ~x288 & ~x314 & ~x315 & ~x336 & ~x338 & ~x339 & ~x340 & ~x365 & ~x366 & ~x367 & ~x393 & ~x396 & ~x398 & ~x399 & ~x421 & ~x448 & ~x728 & ~x756 & ~x757 & ~x759 & ~x783;
assign c9446 =  x239 &  x348 &  x350 &  x375 &  x572 & ~x2 & ~x3 & ~x7 & ~x15 & ~x25 & ~x26 & ~x28 & ~x34 & ~x36 & ~x37 & ~x60 & ~x85 & ~x87 & ~x90 & ~x110 & ~x111 & ~x115 & ~x139 & ~x148 & ~x149 & ~x169 & ~x175 & ~x200 & ~x205 & ~x226 & ~x227 & ~x229 & ~x252 & ~x253 & ~x257 & ~x258 & ~x261 & ~x285 & ~x286 & ~x288 & ~x308 & ~x309 & ~x312 & ~x336 & ~x338 & ~x341 & ~x366 & ~x396 & ~x397 & ~x398 & ~x421 & ~x587 & ~x663 & ~x699 & ~x718 & ~x720 & ~x756 & ~x757 & ~x759 & ~x774;
assign c9448 =  x464 &  x520 &  x529 &  x547 & ~x68 & ~x180 & ~x185 & ~x197 & ~x346 & ~x374 & ~x701;
assign c9450 = ~x1 & ~x33 & ~x41 & ~x46 & ~x49 & ~x55 & ~x69 & ~x70 & ~x73 & ~x79 & ~x84 & ~x102 & ~x108 & ~x120 & ~x123 & ~x133 & ~x140 & ~x144 & ~x148 & ~x150 & ~x178 & ~x182 & ~x195 & ~x197 & ~x198 & ~x226 & ~x234 & ~x236 & ~x254 & ~x263 & ~x286 & ~x287 & ~x291 & ~x309 & ~x337 & ~x338 & ~x366 & ~x367 & ~x368 & ~x393 & ~x395 & ~x420 & ~x422 & ~x482 & ~x483 & ~x484 & ~x675 & ~x731 & ~x755 & ~x761 & ~x762;
assign c9452 =  x156 &  x161 &  x185 &  x188 &  x189 &  x190 &  x211 &  x218 &  x246 &  x272 &  x296 &  x301 &  x303 &  x351 &  x413 &  x415 &  x440 &  x441 & ~x3 & ~x5 & ~x9 & ~x27 & ~x32 & ~x59 & ~x89 & ~x146 & ~x229 & ~x256 & ~x286 & ~x316 & ~x392 & ~x420 & ~x729;
assign c9454 = ~x4 & ~x71 & ~x86 & ~x94 & ~x96 & ~x152 & ~x180 & ~x231 & ~x266 & ~x279 & ~x286 & ~x307 & ~x310 & ~x318 & ~x335 & ~x369 & ~x431 & ~x482 & ~x487 & ~x513 & ~x537 & ~x538;
assign c9456 =  x591 &  x603 &  x622 &  x623 &  x626 & ~x2 & ~x37 & ~x56 & ~x57 & ~x60 & ~x65 & ~x66 & ~x67 & ~x86 & ~x87 & ~x91 & ~x95 & ~x145 & ~x149 & ~x169 & ~x170 & ~x171 & ~x172 & ~x174 & ~x175 & ~x176 & ~x197 & ~x224 & ~x228 & ~x254 & ~x280 & ~x313 & ~x316 & ~x336 & ~x342 & ~x343 & ~x344 & ~x345 & ~x363 & ~x365 & ~x369 & ~x370 & ~x373 & ~x394 & ~x398 & ~x420 & ~x423 & ~x425 & ~x426 & ~x428 & ~x448 & ~x454 & ~x455 & ~x456 & ~x478 & ~x482 & ~x483 & ~x700 & ~x756 & ~x758 & ~x760;
assign c9458 =  x497 &  x524 &  x528 & ~x104 & ~x176 & ~x204 & ~x214 & ~x246 & ~x603 & ~x632 & ~x648 & ~x653 & ~x741 & ~x778;
assign c9460 =  x377 &  x517 & ~x29 & ~x162 & ~x163 & ~x363 & ~x364 & ~x372 & ~x531 & ~x621 & ~x661;
assign c9462 =  x555 &  x580 &  x583 &  x598 & ~x36 & ~x44 & ~x54 & ~x68 & ~x87 & ~x95 & ~x109 & ~x392 & ~x633 & ~x751;
assign c9464 = ~x4 & ~x11 & ~x17 & ~x18 & ~x19 & ~x22 & ~x25 & ~x27 & ~x32 & ~x34 & ~x39 & ~x41 & ~x66 & ~x69 & ~x70 & ~x76 & ~x78 & ~x96 & ~x112 & ~x113 & ~x120 & ~x176 & ~x178 & ~x206 & ~x208 & ~x232 & ~x253 & ~x263 & ~x285 & ~x288 & ~x289 & ~x309 & ~x317 & ~x335 & ~x391 & ~x392 & ~x395 & ~x419 & ~x421 & ~x423 & ~x426 & ~x448 & ~x453 & ~x457 & ~x482 & ~x483 & ~x671 & ~x736 & ~x745 & ~x747 & ~x751 & ~x770 & ~x773 & ~x776 & ~x780;
assign c9466 =  x464 &  x467 &  x491 &  x497 &  x507 &  x549 & ~x1 & ~x41 & ~x51 & ~x54 & ~x77 & ~x92 & ~x159 & ~x182 & ~x197 & ~x204 & ~x232 & ~x312 & ~x317 & ~x320 & ~x399 & ~x744 & ~x749 & ~x775;
assign c9468 =  x299 &  x300 &  x303 &  x356 &  x386 &  x414 &  x525 &  x527 &  x583 & ~x5 & ~x8 & ~x10 & ~x15 & ~x37 & ~x39 & ~x60 & ~x64 & ~x92 & ~x114 & ~x115 & ~x117 & ~x147 & ~x174 & ~x230 & ~x231 & ~x232 & ~x252 & ~x281 & ~x283 & ~x284 & ~x290 & ~x340 & ~x344 & ~x368 & ~x397 & ~x430 & ~x448 & ~x758;
assign c9470 =  x300 &  x379 & ~x16 & ~x45 & ~x120 & ~x149 & ~x152 & ~x176 & ~x186 & ~x252 & ~x310 & ~x562 & ~x577 & ~x634 & ~x636 & ~x697;
assign c9472 =  x303 &  x304 &  x499 &  x534 & ~x16 & ~x39 & ~x41 & ~x51 & ~x66 & ~x94 & ~x102 & ~x120 & ~x124 & ~x128 & ~x142 & ~x148 & ~x153 & ~x231 & ~x401 & ~x423 & ~x631 & ~x644 & ~x678 & ~x695 & ~x717 & ~x765 & ~x782;
assign c9474 =  x294 &  x449 &  x472 & ~x21 & ~x31 & ~x34 & ~x39 & ~x87 & ~x96 & ~x153 & ~x171 & ~x195 & ~x228 & ~x253 & ~x261 & ~x672 & ~x695 & ~x759 & ~x770;
assign c9476 =  x299 &  x423 & ~x476;
assign c9478 =  x471 & ~x13 & ~x133 & ~x185 & ~x289 & ~x373 & ~x591 & ~x730;
assign c9480 =  x21;
assign c9482 =  x185 &  x188 &  x192 &  x246 &  x247 &  x248 &  x296 &  x304 &  x305 &  x386 &  x388 &  x435 & ~x6 & ~x29 & ~x33 & ~x35 & ~x59 & ~x60 & ~x63 & ~x67 & ~x92 & ~x116 & ~x121 & ~x140 & ~x141 & ~x145 & ~x177 & ~x196 & ~x199 & ~x225 & ~x228 & ~x256 & ~x258 & ~x280 & ~x281 & ~x282 & ~x283 & ~x284 & ~x286 & ~x309 & ~x313 & ~x337 & ~x366 & ~x368 & ~x398 & ~x420 & ~x759 & ~x760 & ~x762 & ~x783;
assign c9484 = ~x22 & ~x25 & ~x40 & ~x42 & ~x111 & ~x207 & ~x230 & ~x231 & ~x232 & ~x288 & ~x307 & ~x335 & ~x373 & ~x400 & ~x401 & ~x425 & ~x451 & ~x478 & ~x511 & ~x512 & ~x515 & ~x539 & ~x746 & ~x760;
assign c9486 =  x220 &  x245 &  x246 &  x247 &  x248 &  x269 &  x270 &  x273 &  x298 &  x300 &  x301 &  x327 &  x329 &  x354 &  x358 &  x435 &  x436 &  x513 & ~x4 & ~x27 & ~x35 & ~x37 & ~x55 & ~x58 & ~x64 & ~x67 & ~x84 & ~x85 & ~x90 & ~x94 & ~x197 & ~x198 & ~x204 & ~x254 & ~x258 & ~x287 & ~x340 & ~x367 & ~x368 & ~x690 & ~x691 & ~x755 & ~x756 & ~x757 & ~x770 & ~x771 & ~x781 & ~x782;
assign c9488 =  x409 &  x604 &  x605 &  x626 &  x647 &  x648 &  x658 &  x681 & ~x60 & ~x63 & ~x85 & ~x89 & ~x112 & ~x171 & ~x230 & ~x310 & ~x335 & ~x393 & ~x396 & ~x397 & ~x420 & ~x447 & ~x476 & ~x478 & ~x532 & ~x755 & ~x758 & ~x760;
assign c9490 =  x272 &  x273 &  x274 &  x297 &  x298 &  x324 &  x325 &  x356 &  x357 &  x358 &  x381 &  x385 &  x410 &  x464 &  x465 &  x467 &  x469 & ~x2 & ~x4 & ~x9 & ~x28 & ~x31 & ~x35 & ~x36 & ~x39 & ~x56 & ~x62 & ~x65 & ~x66 & ~x67 & ~x84 & ~x86 & ~x87 & ~x89 & ~x93 & ~x113 & ~x114 & ~x116 & ~x118 & ~x119 & ~x146 & ~x149 & ~x168 & ~x171 & ~x174 & ~x175 & ~x176 & ~x177 & ~x178 & ~x196 & ~x197 & ~x199 & ~x200 & ~x203 & ~x224 & ~x226 & ~x229 & ~x232 & ~x233 & ~x234 & ~x256 & ~x258 & ~x280 & ~x282 & ~x283 & ~x287 & ~x288 & ~x291 & ~x308 & ~x310 & ~x313 & ~x315 & ~x335 & ~x337 & ~x339 & ~x341 & ~x344 & ~x346 & ~x364 & ~x365 & ~x370 & ~x371 & ~x392 & ~x393 & ~x395 & ~x396 & ~x397 & ~x400 & ~x420 & ~x429 & ~x453 & ~x454 & ~x615 & ~x699 & ~x727 & ~x755 & ~x756 & ~x758;
assign c9492 =  x183 &  x405 &  x496 &  x514 & ~x3 & ~x36 & ~x54 & ~x59 & ~x60 & ~x90 & ~x117 & ~x119 & ~x146 & ~x171 & ~x173 & ~x204 & ~x205 & ~x226 & ~x313 & ~x314 & ~x338 & ~x339 & ~x395 & ~x420 & ~x447 & ~x448 & ~x746 & ~x748 & ~x749 & ~x756 & ~x770 & ~x773;
assign c9494 =  x358 &  x479 &  x537 & ~x73 & ~x117 & ~x605 & ~x657 & ~x715;
assign c9496 =  x271 &  x715;
assign c9498 = ~x1 & ~x23 & ~x38 & ~x59 & ~x89 & ~x99 & ~x173 & ~x223 & ~x311 & ~x336 & ~x396 & ~x514 & ~x538 & ~x567 & ~x746;
assign c91 =  x318 & ~x244;
assign c93 =  x269 &  x270 &  x271 &  x272 &  x275 &  x298 &  x301 &  x303 &  x332 &  x359 &  x383 &  x385 &  x387 &  x409 &  x410 &  x412 &  x413 &  x415 &  x432 &  x441 &  x444 &  x462 &  x463 &  x465 &  x467 &  x469 &  x470 &  x474 &  x491 &  x492 &  x496 &  x497 &  x514 &  x524 & ~x6 & ~x8 & ~x15 & ~x17 & ~x27 & ~x28 & ~x32 & ~x34 & ~x44 & ~x45 & ~x46 & ~x49 & ~x57 & ~x66 & ~x70 & ~x72 & ~x74 & ~x75 & ~x78 & ~x84 & ~x85 & ~x88 & ~x89 & ~x92 & ~x96 & ~x97 & ~x109 & ~x111 & ~x114 & ~x124 & ~x127 & ~x134 & ~x139 & ~x140 & ~x142 & ~x145 & ~x154 & ~x155 & ~x161 & ~x165 & ~x167 & ~x170 & ~x176 & ~x193 & ~x195 & ~x199 & ~x201 & ~x204 & ~x223 & ~x224 & ~x233 & ~x234 & ~x236 & ~x254 & ~x256 & ~x279 & ~x280 & ~x289 & ~x308 & ~x314 & ~x319 & ~x339 & ~x341 & ~x342 & ~x364 & ~x369 & ~x370 & ~x397 & ~x398 & ~x419 & ~x422 & ~x448 & ~x615 & ~x623 & ~x627 & ~x628 & ~x629 & ~x631 & ~x633 & ~x634 & ~x635 & ~x636 & ~x639 & ~x642 & ~x645 & ~x648 & ~x650 & ~x655 & ~x660 & ~x667 & ~x670 & ~x672 & ~x676 & ~x677 & ~x687 & ~x690 & ~x697 & ~x698 & ~x707 & ~x709 & ~x713 & ~x721 & ~x722 & ~x723 & ~x727 & ~x737 & ~x748 & ~x750 & ~x751 & ~x757 & ~x760 & ~x771 & ~x775 & ~x782;
assign c95 = ~x303 & ~x329;
assign c97 =  x305 &  x352 &  x383 &  x386 &  x466 &  x471 &  x512 &  x522 &  x527 &  x529 &  x570 &  x578 & ~x20 & ~x24 & ~x28 & ~x33 & ~x35 & ~x40 & ~x42 & ~x45 & ~x65 & ~x79 & ~x89 & ~x101 & ~x115 & ~x117 & ~x123 & ~x131 & ~x138 & ~x143 & ~x146 & ~x148 & ~x149 & ~x159 & ~x163 & ~x181 & ~x183 & ~x200 & ~x209 & ~x219 & ~x235 & ~x251 & ~x252 & ~x254 & ~x256 & ~x264 & ~x283 & ~x284 & ~x312 & ~x313 & ~x319 & ~x335 & ~x368 & ~x588 & ~x615 & ~x634 & ~x636 & ~x640 & ~x642 & ~x652 & ~x666 & ~x669 & ~x684 & ~x687 & ~x693 & ~x698 & ~x709 & ~x711 & ~x713 & ~x718 & ~x720 & ~x723 & ~x733 & ~x735 & ~x736 & ~x738 & ~x745 & ~x751 & ~x759 & ~x762 & ~x777;
assign c99 = ~x301 & ~x531 & ~x670 & ~x698;
assign c911 =  x120;
assign c913 =  x59;
assign c915 =  x145;
assign c917 =  x203;
assign c919 =  x8;
assign c921 = ~x459 & ~x634;
assign c925 =  x232;
assign c927 = ~x36 & ~x53 & ~x105 & ~x110 & ~x209 & ~x340 & ~x346 & ~x395 & ~x398 & ~x422 & ~x478 & ~x504 & ~x560 & ~x598 & ~x601 & ~x602 & ~x604 & ~x608 & ~x609 & ~x626 & ~x628 & ~x629 & ~x635 & ~x637 & ~x638 & ~x642 & ~x671 & ~x684 & ~x687 & ~x730 & ~x741 & ~x751 & ~x762 & ~x763 & ~x765;
assign c929 =  x367;
assign c931 =  x91;
assign c933 =  x773;
assign c935 =  x241 &  x324 &  x333 &  x350 &  x380 &  x381 &  x384 &  x407 &  x409 &  x412 &  x415 &  x416 &  x436 &  x445 &  x463 &  x473 &  x485 &  x490 &  x511 & ~x0 & ~x3 & ~x4 & ~x11 & ~x12 & ~x14 & ~x21 & ~x22 & ~x31 & ~x37 & ~x38 & ~x39 & ~x42 & ~x47 & ~x52 & ~x53 & ~x54 & ~x59 & ~x66 & ~x70 & ~x71 & ~x74 & ~x78 & ~x79 & ~x91 & ~x93 & ~x100 & ~x101 & ~x108 & ~x111 & ~x113 & ~x114 & ~x117 & ~x119 & ~x122 & ~x123 & ~x124 & ~x131 & ~x132 & ~x133 & ~x139 & ~x153 & ~x154 & ~x165 & ~x167 & ~x168 & ~x170 & ~x173 & ~x177 & ~x178 & ~x180 & ~x181 & ~x183 & ~x194 & ~x195 & ~x196 & ~x198 & ~x201 & ~x204 & ~x217 & ~x222 & ~x223 & ~x227 & ~x231 & ~x232 & ~x249 & ~x253 & ~x256 & ~x282 & ~x284 & ~x287 & ~x308 & ~x311 & ~x314 & ~x316 & ~x317 & ~x367 & ~x420 & ~x588 & ~x593 & ~x619 & ~x626 & ~x627 & ~x631 & ~x642 & ~x646 & ~x650 & ~x654 & ~x665 & ~x668 & ~x670 & ~x676 & ~x682 & ~x684 & ~x693 & ~x700 & ~x701 & ~x706 & ~x713 & ~x715 & ~x719 & ~x720 & ~x726 & ~x730 & ~x731 & ~x734 & ~x738 & ~x746 & ~x747 & ~x754 & ~x755 & ~x756 & ~x761 & ~x763 & ~x767 & ~x769 & ~x771 & ~x773 & ~x775 & ~x778 & ~x781;
assign c937 =  x117;
assign c939 =  x397 & ~x273;
assign c941 =  x297 & ~x1 & ~x20 & ~x22 & ~x33 & ~x34 & ~x45 & ~x63 & ~x88 & ~x96 & ~x104 & ~x116 & ~x121 & ~x129 & ~x153 & ~x154 & ~x179 & ~x232 & ~x235 & ~x253 & ~x254 & ~x277 & ~x320 & ~x364 & ~x394 & ~x448 & ~x692 & ~x722 & ~x749 & ~x752 & ~x770 & ~x779;
assign c943 =  x443 & ~x463 & ~x561;
assign c945 =  x3 &  x149 &  x420;
assign c947 = ~x361 & ~x610;
assign c949 =  x283;
assign c951 = ~x492 & ~x607;
assign c953 =  x289;
assign c955 =  x270 &  x440 &  x466 &  x482 &  x483 &  x512 & ~x33 & ~x45 & ~x54 & ~x83 & ~x85 & ~x124 & ~x141 & ~x166 & ~x230 & ~x313 & ~x314 & ~x368 & ~x503 & ~x506 & ~x643 & ~x671 & ~x718 & ~x768;
assign c957 =  x87;
assign c959 =  x226;
assign c961 =  x88;
assign c963 =  x342;
assign c965 =  x119;
assign c967 =  x242 &  x352 &  x355 &  x359 &  x388 &  x414 &  x440 &  x441 &  x459 &  x460 &  x471 &  x473 &  x482 &  x516 &  x556 &  x557 &  x604 &  x605 & ~x3 & ~x31 & ~x36 & ~x47 & ~x55 & ~x85 & ~x103 & ~x113 & ~x114 & ~x134 & ~x141 & ~x145 & ~x147 & ~x148 & ~x151 & ~x154 & ~x176 & ~x182 & ~x237 & ~x263 & ~x288 & ~x307 & ~x315 & ~x337 & ~x363 & ~x371 & ~x421 & ~x588 & ~x648 & ~x659 & ~x663 & ~x666 & ~x674 & ~x679 & ~x698 & ~x712 & ~x739 & ~x740 & ~x741 & ~x761 & ~x767 & ~x768 & ~x777;
assign c969 =  x368;
assign c971 =  x35;
assign c973 =  x118;
assign c975 =  x455 & ~x348 & ~x423 & ~x424 & ~x450 & ~x690;
assign c977 =  x341 &  x392;
assign c979 = ~x115 & ~x120 & ~x503 & ~x545 & ~x606 & ~x634;
assign c981 =  x332 &  x405 &  x442 &  x446 &  x513 & ~x1 & ~x3 & ~x10 & ~x22 & ~x23 & ~x41 & ~x99 & ~x225 & ~x257 & ~x321 & ~x336 & ~x394 & ~x397 & ~x422 & ~x447 & ~x450 & ~x588 & ~x662 & ~x667 & ~x705 & ~x717 & ~x747 & ~x772;
assign c983 =  x54;
assign c985 =  x36;
assign c987 =  x273 &  x512 & ~x1 & ~x5 & ~x8 & ~x9 & ~x10 & ~x15 & ~x21 & ~x22 & ~x27 & ~x35 & ~x38 & ~x41 & ~x53 & ~x64 & ~x70 & ~x72 & ~x80 & ~x90 & ~x91 & ~x105 & ~x109 & ~x113 & ~x123 & ~x126 & ~x137 & ~x138 & ~x139 & ~x143 & ~x144 & ~x148 & ~x165 & ~x166 & ~x169 & ~x175 & ~x199 & ~x206 & ~x209 & ~x223 & ~x235 & ~x254 & ~x258 & ~x260 & ~x261 & ~x281 & ~x287 & ~x289 & ~x310 & ~x316 & ~x319 & ~x336 & ~x339 & ~x344 & ~x368 & ~x392 & ~x393 & ~x396 & ~x422 & ~x424 & ~x448 & ~x449 & ~x478 & ~x479 & ~x644 & ~x671 & ~x672 & ~x674 & ~x689 & ~x691 & ~x710 & ~x712 & ~x713 & ~x714 & ~x715 & ~x724 & ~x725 & ~x731 & ~x732 & ~x736 & ~x744 & ~x753 & ~x760 & ~x764 & ~x768 & ~x769 & ~x771 & ~x780;
assign c989 = ~x461;
assign c991 =  x60;
assign c993 =  x359 & ~x1 & ~x4 & ~x7 & ~x8 & ~x14 & ~x25 & ~x29 & ~x30 & ~x31 & ~x33 & ~x35 & ~x43 & ~x44 & ~x45 & ~x49 & ~x51 & ~x53 & ~x57 & ~x59 & ~x61 & ~x65 & ~x68 & ~x71 & ~x77 & ~x81 & ~x84 & ~x88 & ~x90 & ~x94 & ~x95 & ~x106 & ~x110 & ~x115 & ~x119 & ~x121 & ~x122 & ~x124 & ~x127 & ~x129 & ~x130 & ~x134 & ~x139 & ~x145 & ~x147 & ~x148 & ~x149 & ~x151 & ~x155 & ~x157 & ~x159 & ~x160 & ~x161 & ~x164 & ~x170 & ~x173 & ~x174 & ~x175 & ~x176 & ~x183 & ~x189 & ~x190 & ~x197 & ~x198 & ~x200 & ~x205 & ~x208 & ~x220 & ~x221 & ~x222 & ~x224 & ~x229 & ~x235 & ~x236 & ~x237 & ~x247 & ~x248 & ~x249 & ~x250 & ~x253 & ~x254 & ~x256 & ~x280 & ~x282 & ~x283 & ~x287 & ~x307 & ~x312 & ~x315 & ~x316 & ~x342 & ~x365 & ~x391 & ~x394 & ~x419 & ~x447 & ~x475 & ~x560 & ~x589 & ~x620 & ~x624 & ~x627 & ~x629 & ~x632 & ~x636 & ~x639 & ~x640 & ~x642 & ~x645 & ~x646 & ~x649 & ~x651 & ~x654 & ~x658 & ~x660 & ~x663 & ~x664 & ~x666 & ~x672 & ~x675 & ~x676 & ~x682 & ~x683 & ~x686 & ~x694 & ~x695 & ~x697 & ~x699 & ~x701 & ~x702 & ~x703 & ~x704 & ~x708 & ~x709 & ~x711 & ~x714 & ~x719 & ~x727 & ~x731 & ~x733 & ~x734 & ~x737 & ~x740 & ~x741 & ~x752 & ~x753 & ~x757 & ~x759 & ~x760 & ~x761 & ~x762 & ~x764 & ~x769 & ~x772 & ~x773 & ~x775 & ~x776 & ~x777 & ~x779 & ~x783;
assign c995 = ~x351 & ~x383;
assign c997 =  x746;
assign c999 =  x280;
assign c9101 =  x8;
assign c9103 =  x745;
assign c9105 =  x233;
assign c9107 =  x56;
assign c9109 =  x120;
assign c9111 =  x141;
assign c9113 =  x772;
assign c9115 =  x370;
assign c9117 =  x6 &  x771;
assign c9119 =  x415 & ~x0 & ~x2 & ~x9 & ~x10 & ~x14 & ~x18 & ~x34 & ~x37 & ~x38 & ~x43 & ~x62 & ~x63 & ~x68 & ~x69 & ~x91 & ~x96 & ~x142 & ~x145 & ~x150 & ~x166 & ~x176 & ~x224 & ~x229 & ~x281 & ~x282 & ~x311 & ~x364 & ~x393 & ~x395 & ~x396 & ~x397 & ~x398 & ~x421 & ~x476 & ~x506 & ~x590 & ~x633 & ~x636 & ~x643 & ~x698 & ~x715 & ~x717 & ~x719 & ~x720 & ~x729 & ~x732 & ~x742 & ~x758 & ~x759 & ~x762 & ~x764 & ~x769 & ~x773 & ~x777;
assign c9121 =  x115;
assign c9123 =  x12;
assign c9125 =  x149;
assign c9127 = ~x323 & ~x517 & ~x631;
assign c9129 =  x214 &  x242 &  x359 &  x386 &  x388 &  x414 &  x418 &  x446 &  x458 &  x462 &  x500 &  x513 &  x542 &  x550 &  x551 &  x552 & ~x3 & ~x19 & ~x20 & ~x52 & ~x60 & ~x65 & ~x82 & ~x84 & ~x87 & ~x109 & ~x136 & ~x162 & ~x166 & ~x174 & ~x181 & ~x195 & ~x200 & ~x292 & ~x310 & ~x339 & ~x343 & ~x395 & ~x398 & ~x399 & ~x420 & ~x422 & ~x450 & ~x476 & ~x588 & ~x649 & ~x682 & ~x683 & ~x706 & ~x714 & ~x734 & ~x736 & ~x738 & ~x752 & ~x754 & ~x778;
assign c9131 =  x326 &  x468 &  x510 &  x549 & ~x41 & ~x42 & ~x209 & ~x221 & ~x394 & ~x395 & ~x475 & ~x613 & ~x631 & ~x638 & ~x640 & ~x648 & ~x651 & ~x661 & ~x694 & ~x721 & ~x725;
assign c9133 = ~x379;
assign c9135 =  x269 & ~x90 & ~x93 & ~x96 & ~x109 & ~x121 & ~x140 & ~x147 & ~x211 & ~x320 & ~x366 & ~x422 & ~x536 & ~x633 & ~x671 & ~x698 & ~x722 & ~x741 & ~x775 & ~x777 & ~x779;
assign c9137 =  x325 &  x347 & ~x273 & ~x589 & ~x590 & ~x617 & ~x620;
assign c9139 = ~x323 & ~x353;
assign c9141 =  x368;
assign c9143 =  x120;
assign c9145 =  x268 &  x400 &  x468 &  x482 & ~x10 & ~x20 & ~x43 & ~x65 & ~x66 & ~x75 & ~x76 & ~x120 & ~x122 & ~x124 & ~x134 & ~x143 & ~x147 & ~x150 & ~x163 & ~x167 & ~x172 & ~x187 & ~x194 & ~x223 & ~x245 & ~x252 & ~x338 & ~x419 & ~x532 & ~x615 & ~x655 & ~x664 & ~x666 & ~x702 & ~x705 & ~x734 & ~x737 & ~x750 & ~x773 & ~x780;
assign c9147 =  x417 & ~x20 & ~x50 & ~x249 & ~x349 & ~x718;
assign c9149 = ~x407;
assign c9151 =  x368;
assign c9153 =  x242 &  x528 &  x529 & ~x28 & ~x56 & ~x173 & ~x282 & ~x293 & ~x392 & ~x506 & ~x670 & ~x777;
assign c9155 =  x412 &  x442 & ~x16 & ~x321 & ~x376 & ~x636;
assign c9159 =  x370;
assign c9161 =  x312;
assign c9163 =  x399 &  x514 &  x537 & ~x159 & ~x210 & ~x245 & ~x307;
assign c9167 =  x261;
assign c9169 =  x372;
assign c9171 =  x758;
assign c9173 =  x439 &  x467 &  x508 & ~x9 & ~x12 & ~x13 & ~x15 & ~x17 & ~x18 & ~x19 & ~x21 & ~x26 & ~x30 & ~x33 & ~x34 & ~x35 & ~x38 & ~x42 & ~x44 & ~x45 & ~x51 & ~x54 & ~x66 & ~x74 & ~x77 & ~x83 & ~x85 & ~x88 & ~x91 & ~x102 & ~x105 & ~x113 & ~x125 & ~x133 & ~x135 & ~x137 & ~x138 & ~x141 & ~x146 & ~x166 & ~x170 & ~x173 & ~x175 & ~x179 & ~x193 & ~x195 & ~x222 & ~x223 & ~x229 & ~x251 & ~x283 & ~x289 & ~x290 & ~x308 & ~x310 & ~x311 & ~x342 & ~x364 & ~x366 & ~x421 & ~x422 & ~x423 & ~x585 & ~x608 & ~x609 & ~x644 & ~x645 & ~x652 & ~x661 & ~x663 & ~x665 & ~x673 & ~x674 & ~x675 & ~x677 & ~x683 & ~x686 & ~x691 & ~x693 & ~x707 & ~x709 & ~x712 & ~x723 & ~x726 & ~x729 & ~x730 & ~x732 & ~x733 & ~x735 & ~x738 & ~x739 & ~x749 & ~x754 & ~x758 & ~x760 & ~x779 & ~x782;
assign c9175 =  x373 &  x375 &  x384 &  x494 &  x516 & ~x6 & ~x68 & ~x71 & ~x72 & ~x93 & ~x96 & ~x97 & ~x98 & ~x105 & ~x108 & ~x118 & ~x121 & ~x201 & ~x250 & ~x365 & ~x420 & ~x587 & ~x593 & ~x635 & ~x636 & ~x652 & ~x673 & ~x695 & ~x710 & ~x723 & ~x734 & ~x737 & ~x742 & ~x781 & ~x782;
assign c9177 =  x91;
assign c9179 =  x399 & ~x394;
assign c9181 =  x343;
assign c9183 =  x66;
assign c9185 =  x270 &  x271 &  x361 &  x383 &  x384 &  x385 &  x389 &  x414 &  x417 &  x418 &  x442 &  x446 &  x482 &  x483 &  x487 &  x493 &  x495 &  x498 &  x500 &  x501 &  x521 &  x525 &  x526 &  x528 & ~x0 & ~x1 & ~x11 & ~x24 & ~x35 & ~x36 & ~x37 & ~x40 & ~x41 & ~x57 & ~x65 & ~x69 & ~x72 & ~x84 & ~x91 & ~x93 & ~x94 & ~x96 & ~x100 & ~x106 & ~x107 & ~x112 & ~x114 & ~x118 & ~x124 & ~x125 & ~x128 & ~x129 & ~x130 & ~x138 & ~x141 & ~x154 & ~x155 & ~x160 & ~x161 & ~x166 & ~x171 & ~x173 & ~x179 & ~x190 & ~x194 & ~x198 & ~x222 & ~x225 & ~x233 & ~x234 & ~x254 & ~x257 & ~x258 & ~x262 & ~x263 & ~x280 & ~x284 & ~x307 & ~x312 & ~x315 & ~x319 & ~x335 & ~x338 & ~x366 & ~x367 & ~x391 & ~x392 & ~x419 & ~x422 & ~x503 & ~x615 & ~x632 & ~x642 & ~x644 & ~x646 & ~x653 & ~x657 & ~x660 & ~x661 & ~x662 & ~x663 & ~x669 & ~x673 & ~x679 & ~x687 & ~x697 & ~x705 & ~x706 & ~x710 & ~x713 & ~x716 & ~x718 & ~x720 & ~x722 & ~x724 & ~x743 & ~x744 & ~x752 & ~x755 & ~x757 & ~x761 & ~x764 & ~x769 & ~x771 & ~x772 & ~x777 & ~x780 & ~x781;
assign c9187 =  x717;
assign c9189 =  x337;
assign c9191 = ~x397 & ~x545 & ~x562 & ~x589 & ~x601 & ~x618 & ~x634;
assign c9193 = ~x54 & ~x113 & ~x146 & ~x197 & ~x222 & ~x223 & ~x259 & ~x339 & ~x525 & ~x580 & ~x589 & ~x590 & ~x608 & ~x750 & ~x777;
assign c9195 = ~x6 & ~x17 & ~x18 & ~x22 & ~x27 & ~x52 & ~x64 & ~x81 & ~x96 & ~x105 & ~x114 & ~x115 & ~x141 & ~x191 & ~x201 & ~x203 & ~x232 & ~x233 & ~x249 & ~x250 & ~x283 & ~x364 & ~x420 & ~x447 & ~x584 & ~x586 & ~x610 & ~x644 & ~x650 & ~x652 & ~x667 & ~x696 & ~x698 & ~x724 & ~x739 & ~x750 & ~x767 & ~x779 & ~x781;
assign c9197 =  x306 & ~x324 & ~x348 & ~x375;
assign c9201 =  x4;
assign c9203 =  x8;
assign c9205 =  x371;
assign c9207 =  x36;
assign c9209 =  x367;
assign c9211 =  x343;
assign c9213 =  x259 &  x315;
assign c9215 =  x369;
assign c9217 =  x214 &  x299 &  x301 &  x325 &  x327 &  x328 &  x351 &  x378 &  x381 &  x386 &  x388 &  x405 &  x415 &  x416 &  x431 &  x434 &  x436 &  x437 &  x439 &  x442 &  x457 &  x459 &  x462 &  x463 &  x470 &  x471 &  x486 &  x493 &  x496 &  x497 &  x508 &  x509 &  x511 &  x512 &  x514 &  x518 &  x520 &  x523 &  x526 &  x528 & ~x10 & ~x13 & ~x15 & ~x17 & ~x26 & ~x27 & ~x30 & ~x31 & ~x33 & ~x40 & ~x43 & ~x45 & ~x46 & ~x47 & ~x49 & ~x51 & ~x57 & ~x58 & ~x61 & ~x62 & ~x63 & ~x65 & ~x73 & ~x76 & ~x78 & ~x81 & ~x82 & ~x85 & ~x92 & ~x95 & ~x96 & ~x100 & ~x104 & ~x106 & ~x112 & ~x115 & ~x124 & ~x125 & ~x130 & ~x132 & ~x135 & ~x136 & ~x137 & ~x139 & ~x141 & ~x145 & ~x148 & ~x150 & ~x160 & ~x164 & ~x166 & ~x171 & ~x172 & ~x175 & ~x176 & ~x179 & ~x189 & ~x191 & ~x193 & ~x195 & ~x197 & ~x203 & ~x207 & ~x208 & ~x209 & ~x224 & ~x227 & ~x229 & ~x231 & ~x233 & ~x236 & ~x252 & ~x255 & ~x256 & ~x259 & ~x263 & ~x281 & ~x282 & ~x291 & ~x307 & ~x310 & ~x311 & ~x312 & ~x336 & ~x363 & ~x365 & ~x371 & ~x372 & ~x391 & ~x423 & ~x424 & ~x449 & ~x588 & ~x616 & ~x619 & ~x644 & ~x652 & ~x659 & ~x662 & ~x665 & ~x669 & ~x672 & ~x673 & ~x675 & ~x677 & ~x678 & ~x683 & ~x688 & ~x689 & ~x693 & ~x697 & ~x702 & ~x704 & ~x706 & ~x709 & ~x711 & ~x712 & ~x713 & ~x715 & ~x716 & ~x718 & ~x719 & ~x729 & ~x737 & ~x739 & ~x741 & ~x743 & ~x746 & ~x753 & ~x754 & ~x762 & ~x763 & ~x764 & ~x765 & ~x770 & ~x773 & ~x778 & ~x780;
assign c9219 =  x142;
assign c9221 = ~x517 & ~x579;
assign c9223 =  x149;
assign c9225 = ~x525 & ~x543 & ~x580 & ~x666;
assign c9227 =  x445 &  x471 &  x499 & ~x9 & ~x12 & ~x29 & ~x41 & ~x42 & ~x57 & ~x98 & ~x109 & ~x148 & ~x150 & ~x176 & ~x184 & ~x200 & ~x289 & ~x312 & ~x315 & ~x318 & ~x343 & ~x367 & ~x395 & ~x396 & ~x420 & ~x507 & ~x636 & ~x643 & ~x660 & ~x661 & ~x662 & ~x663 & ~x690 & ~x692 & ~x719 & ~x771;
assign c9229 =  x481 & ~x131 & ~x222 & ~x278 & ~x503 & ~x609 & ~x631 & ~x634 & ~x635 & ~x642 & ~x665 & ~x688 & ~x694;
assign c9231 =  x393;
assign c9233 =  x176;
assign c9235 = ~x489 & ~x586;
assign c9237 = ~x489 & ~x610;
assign c9239 =  x142;
assign c9241 =  x286 &  x288;
assign c9243 =  x60;
assign c9245 =  x65;
assign c9247 =  x312;
assign c9249 =  x62;
assign c9251 =  x420;
assign c9253 =  x229;
assign c9255 =  x341;
assign c9257 =  x11;
assign c9261 =  x399 & ~x245;
assign c9263 =  x168;
assign c9265 =  x365;
assign c9267 =  x448 & ~x273;
assign c9269 =  x145;
assign c9271 =  x215 &  x538 & ~x9 & ~x13 & ~x24 & ~x27 & ~x28 & ~x29 & ~x37 & ~x60 & ~x116 & ~x140 & ~x166 & ~x203 & ~x222 & ~x228 & ~x230 & ~x280 & ~x284 & ~x294 & ~x336 & ~x422 & ~x450 & ~x675 & ~x724 & ~x725 & ~x727 & ~x760 & ~x767 & ~x782;
assign c9273 =  x62;
assign c9275 =  x62;
assign c9277 =  x470 &  x498 &  x510 & ~x155 & ~x195 & ~x422 & ~x479 & ~x643;
assign c9279 =  x556 & ~x492;
assign c9281 =  x175;
assign c9283 =  x32;
assign c9285 =  x399 & ~x245 & ~x273;
assign c9287 =  x93 &  x772;
assign c9289 =  x400 &  x509 &  x549 & ~x32 & ~x109 & ~x151 & ~x160 & ~x189 & ~x206 & ~x219 & ~x222 & ~x223 & ~x229 & ~x610 & ~x622 & ~x639 & ~x642 & ~x648 & ~x654;
assign c9291 =  x365;
assign c9293 = ~x0 & ~x11 & ~x16 & ~x22 & ~x25 & ~x28 & ~x29 & ~x31 & ~x32 & ~x35 & ~x36 & ~x43 & ~x46 & ~x51 & ~x52 & ~x53 & ~x67 & ~x71 & ~x73 & ~x77 & ~x90 & ~x91 & ~x96 & ~x98 & ~x113 & ~x115 & ~x120 & ~x125 & ~x130 & ~x137 & ~x138 & ~x141 & ~x145 & ~x151 & ~x156 & ~x157 & ~x166 & ~x173 & ~x174 & ~x193 & ~x194 & ~x197 & ~x198 & ~x202 & ~x207 & ~x225 & ~x229 & ~x232 & ~x239 & ~x253 & ~x257 & ~x263 & ~x280 & ~x282 & ~x289 & ~x293 & ~x336 & ~x343 & ~x366 & ~x368 & ~x394 & ~x395 & ~x396 & ~x420 & ~x423 & ~x560 & ~x573 & ~x594 & ~x603 & ~x616 & ~x621 & ~x625 & ~x633 & ~x644 & ~x645 & ~x646 & ~x648 & ~x656 & ~x657 & ~x664 & ~x667 & ~x669 & ~x676 & ~x677 & ~x678 & ~x680 & ~x683 & ~x684 & ~x685 & ~x686 & ~x691 & ~x693 & ~x694 & ~x695 & ~x705 & ~x721 & ~x725 & ~x726 & ~x728 & ~x729 & ~x732 & ~x734 & ~x739 & ~x750 & ~x752 & ~x753 & ~x756 & ~x757 & ~x758 & ~x771 & ~x772 & ~x776 & ~x783;
assign c9295 =  x452 & ~x247 & ~x555;
assign c9297 =  x313;
assign c9299 =  x325 &  x414 &  x466 &  x502 & ~x3 & ~x4 & ~x8 & ~x25 & ~x35 & ~x48 & ~x51 & ~x52 & ~x53 & ~x62 & ~x63 & ~x79 & ~x89 & ~x96 & ~x106 & ~x111 & ~x117 & ~x126 & ~x135 & ~x139 & ~x140 & ~x160 & ~x165 & ~x171 & ~x179 & ~x183 & ~x222 & ~x224 & ~x228 & ~x235 & ~x261 & ~x264 & ~x284 & ~x312 & ~x338 & ~x593 & ~x600 & ~x612 & ~x614 & ~x617 & ~x620 & ~x636 & ~x642 & ~x666 & ~x673 & ~x675 & ~x677 & ~x691 & ~x698 & ~x708 & ~x710 & ~x714 & ~x736 & ~x741 & ~x749 & ~x763 & ~x765 & ~x768 & ~x769;
assign c9301 =  x120;
assign c9303 =  x418 &  x445 & ~x409;
assign c9305 =  x539 & ~x406 & ~x407;
assign c9307 =  x372 & ~x586 & ~x614;
assign c9309 =  x392;
assign c9311 =  x198;
assign c9313 = ~x553 & ~x580 & ~x583 & ~x585 & ~x610 & ~x611 & ~x636 & ~x653 & ~x666;
assign c9315 =  x297 &  x325 &  x326 &  x477 & ~x187 & ~x668;
assign c9317 =  x771;
assign c9319 =  x28;
assign c9321 = ~x15 & ~x81 & ~x149 & ~x161 & ~x177 & ~x249 & ~x250 & ~x275 & ~x309 & ~x367 & ~x531 & ~x532 & ~x560 & ~x612 & ~x706 & ~x720 & ~x722 & ~x726 & ~x750;
assign c9323 = ~x489 & ~x551 & ~x579 & ~x606;
assign c9325 =  x242 &  x243 &  x297 &  x333 &  x353 &  x355 &  x381 &  x414 &  x416 &  x445 &  x458 &  x513 &  x514 &  x525 &  x526 &  x555 &  x605 & ~x12 & ~x14 & ~x18 & ~x47 & ~x54 & ~x61 & ~x67 & ~x72 & ~x73 & ~x74 & ~x79 & ~x84 & ~x104 & ~x108 & ~x113 & ~x125 & ~x139 & ~x144 & ~x148 & ~x163 & ~x173 & ~x178 & ~x197 & ~x199 & ~x226 & ~x252 & ~x289 & ~x309 & ~x310 & ~x338 & ~x339 & ~x365 & ~x423 & ~x451 & ~x698 & ~x714 & ~x716 & ~x723 & ~x730 & ~x733 & ~x734 & ~x736 & ~x738 & ~x743 & ~x744 & ~x770 & ~x773 & ~x781 & ~x783;
assign c9327 =  x60;
assign c9329 =  x242 &  x270 &  x356 &  x360 &  x380 &  x382 &  x384 &  x387 &  x388 &  x406 &  x407 &  x409 &  x441 &  x442 &  x456 &  x461 &  x464 &  x465 &  x474 &  x492 &  x493 &  x495 &  x498 &  x508 & ~x3 & ~x4 & ~x8 & ~x9 & ~x12 & ~x13 & ~x17 & ~x20 & ~x23 & ~x25 & ~x26 & ~x29 & ~x31 & ~x34 & ~x37 & ~x41 & ~x42 & ~x46 & ~x49 & ~x51 & ~x55 & ~x59 & ~x61 & ~x65 & ~x70 & ~x75 & ~x80 & ~x83 & ~x84 & ~x85 & ~x87 & ~x93 & ~x94 & ~x100 & ~x104 & ~x106 & ~x109 & ~x110 & ~x113 & ~x117 & ~x118 & ~x121 & ~x125 & ~x132 & ~x136 & ~x148 & ~x160 & ~x161 & ~x164 & ~x166 & ~x167 & ~x172 & ~x176 & ~x182 & ~x183 & ~x191 & ~x192 & ~x193 & ~x195 & ~x196 & ~x198 & ~x200 & ~x201 & ~x202 & ~x210 & ~x224 & ~x225 & ~x231 & ~x235 & ~x252 & ~x254 & ~x257 & ~x261 & ~x264 & ~x280 & ~x285 & ~x286 & ~x288 & ~x289 & ~x308 & ~x310 & ~x316 & ~x317 & ~x339 & ~x341 & ~x343 & ~x345 & ~x364 & ~x366 & ~x371 & ~x392 & ~x397 & ~x399 & ~x422 & ~x423 & ~x424 & ~x425 & ~x448 & ~x615 & ~x617 & ~x633 & ~x636 & ~x637 & ~x638 & ~x642 & ~x643 & ~x644 & ~x646 & ~x648 & ~x652 & ~x653 & ~x662 & ~x663 & ~x664 & ~x665 & ~x667 & ~x668 & ~x670 & ~x681 & ~x685 & ~x688 & ~x692 & ~x694 & ~x695 & ~x698 & ~x701 & ~x703 & ~x709 & ~x714 & ~x724 & ~x727 & ~x737 & ~x738 & ~x739 & ~x742 & ~x743 & ~x746 & ~x748 & ~x754 & ~x755 & ~x758 & ~x759 & ~x763 & ~x764 & ~x770 & ~x771 & ~x777;
assign c9331 =  x85;
assign c9333 =  x387 &  x415 & ~x8 & ~x11 & ~x17 & ~x18 & ~x19 & ~x51 & ~x78 & ~x89 & ~x103 & ~x111 & ~x174 & ~x179 & ~x180 & ~x194 & ~x198 & ~x223 & ~x232 & ~x247 & ~x248 & ~x276 & ~x315 & ~x448 & ~x532 & ~x561 & ~x775;
assign c9335 =  x117;
assign c9337 =  x745;
assign c9339 =  x757;
assign c9341 =  x358 & ~x354 & ~x586;
assign c9343 =  x253;
assign c9345 = ~x273 & ~x527;
assign c9347 =  x311;
assign c9349 =  x417 &  x499 & ~x407 & ~x604;
assign c9351 =  x479 & ~x273 & ~x602 & ~x613;
assign c9353 =  x596 & ~x0 & ~x49 & ~x53 & ~x102 & ~x141 & ~x177 & ~x194 & ~x200 & ~x205 & ~x206 & ~x227 & ~x262 & ~x317 & ~x321 & ~x368 & ~x615 & ~x636 & ~x692;
assign c9355 =  x282;
assign c9357 =  x400 & ~x272 & ~x613;
assign c9359 =  x362 & ~x461;
assign c9361 = ~x305 & ~x489;
assign c9363 =  x309;
assign c9365 =  x29;
assign c9367 =  x242 & ~x1 & ~x9 & ~x20 & ~x22 & ~x24 & ~x29 & ~x32 & ~x34 & ~x37 & ~x51 & ~x55 & ~x60 & ~x78 & ~x79 & ~x80 & ~x87 & ~x100 & ~x105 & ~x118 & ~x129 & ~x130 & ~x136 & ~x142 & ~x178 & ~x183 & ~x193 & ~x194 & ~x208 & ~x223 & ~x237 & ~x256 & ~x309 & ~x312 & ~x340 & ~x364 & ~x365 & ~x370 & ~x392 & ~x393 & ~x394 & ~x449 & ~x450 & ~x504 & ~x604 & ~x607 & ~x608 & ~x634 & ~x646 & ~x657 & ~x661 & ~x664 & ~x665 & ~x681 & ~x690 & ~x694 & ~x697 & ~x698 & ~x702 & ~x707 & ~x713 & ~x715 & ~x720 & ~x725 & ~x729 & ~x731 & ~x754 & ~x757 & ~x764 & ~x773 & ~x780 & ~x782;
assign c9369 =  x339;
assign c9371 =  x147;
assign c9373 =  x30;
assign c9375 =  x26;
assign c9377 =  x271 &  x272 &  x297 &  x352 &  x358 &  x381 &  x384 &  x413 &  x430 &  x432 &  x438 &  x456 &  x460 &  x474 &  x494 &  x512 &  x553 &  x604 & ~x28 & ~x42 & ~x45 & ~x48 & ~x50 & ~x84 & ~x115 & ~x140 & ~x143 & ~x182 & ~x201 & ~x206 & ~x229 & ~x253 & ~x261 & ~x285 & ~x291 & ~x368 & ~x392 & ~x394 & ~x396 & ~x651 & ~x662 & ~x663 & ~x707 & ~x723 & ~x726 & ~x738 & ~x742 & ~x745 & ~x757 & ~x758 & ~x769 & ~x774 & ~x776;
assign c9379 =  x324 & ~x292 & ~x543 & ~x601 & ~x608;
assign c9381 = ~x379;
assign c9383 =  x205;
assign c9385 = ~x4 & ~x5 & ~x6 & ~x10 & ~x11 & ~x16 & ~x17 & ~x18 & ~x22 & ~x25 & ~x26 & ~x33 & ~x35 & ~x36 & ~x50 & ~x52 & ~x53 & ~x56 & ~x57 & ~x60 & ~x68 & ~x77 & ~x78 & ~x79 & ~x81 & ~x83 & ~x85 & ~x86 & ~x101 & ~x103 & ~x104 & ~x108 & ~x109 & ~x110 & ~x115 & ~x116 & ~x117 & ~x120 & ~x122 & ~x124 & ~x129 & ~x133 & ~x134 & ~x137 & ~x148 & ~x150 & ~x158 & ~x160 & ~x163 & ~x169 & ~x170 & ~x177 & ~x179 & ~x181 & ~x182 & ~x189 & ~x193 & ~x195 & ~x196 & ~x205 & ~x207 & ~x208 & ~x226 & ~x229 & ~x251 & ~x252 & ~x253 & ~x254 & ~x259 & ~x260 & ~x262 & ~x263 & ~x280 & ~x281 & ~x286 & ~x315 & ~x316 & ~x336 & ~x344 & ~x364 & ~x365 & ~x367 & ~x392 & ~x393 & ~x395 & ~x422 & ~x423 & ~x476 & ~x535 & ~x616 & ~x617 & ~x620 & ~x621 & ~x622 & ~x625 & ~x632 & ~x633 & ~x639 & ~x642 & ~x643 & ~x644 & ~x645 & ~x647 & ~x649 & ~x650 & ~x651 & ~x657 & ~x664 & ~x668 & ~x669 & ~x671 & ~x673 & ~x674 & ~x675 & ~x677 & ~x691 & ~x693 & ~x694 & ~x695 & ~x696 & ~x699 & ~x701 & ~x702 & ~x703 & ~x705 & ~x718 & ~x722 & ~x723 & ~x734 & ~x735 & ~x736 & ~x741 & ~x742 & ~x745 & ~x746 & ~x749 & ~x751 & ~x752 & ~x753 & ~x754 & ~x756 & ~x757 & ~x758 & ~x763 & ~x765 & ~x766 & ~x767 & ~x772 & ~x773 & ~x774 & ~x775 & ~x780 & ~x781;
assign c9387 =  x92;
assign c9389 =  x566 & ~x350;
assign c9391 = ~x13 & ~x36 & ~x51 & ~x53 & ~x81 & ~x115 & ~x136 & ~x252 & ~x320 & ~x363 & ~x422 & ~x423 & ~x579 & ~x580 & ~x631 & ~x632 & ~x691 & ~x754 & ~x762 & ~x763 & ~x773;
assign c9393 =  x443 & ~x494;
assign c9395 =  x167;
assign c9397 =  x757;
assign c9399 =  x390 &  x446 & ~x321;
assign c9401 =  x362 & ~x280 & ~x348 & ~x506 & ~x615 & ~x643;
assign c9403 =  x215 &  x243 &  x324 &  x387 &  x416 &  x469 &  x471 &  x488 &  x497 &  x511 & ~x10 & ~x12 & ~x16 & ~x17 & ~x19 & ~x23 & ~x40 & ~x43 & ~x45 & ~x58 & ~x61 & ~x65 & ~x68 & ~x71 & ~x72 & ~x73 & ~x85 & ~x86 & ~x87 & ~x88 & ~x93 & ~x96 & ~x98 & ~x104 & ~x117 & ~x129 & ~x135 & ~x138 & ~x141 & ~x148 & ~x164 & ~x182 & ~x191 & ~x192 & ~x193 & ~x199 & ~x200 & ~x203 & ~x207 & ~x208 & ~x209 & ~x254 & ~x258 & ~x279 & ~x319 & ~x347 & ~x365 & ~x397 & ~x420 & ~x422 & ~x425 & ~x452 & ~x476 & ~x645 & ~x672 & ~x674 & ~x678 & ~x689 & ~x691 & ~x699 & ~x713 & ~x714 & ~x718 & ~x723 & ~x728 & ~x742 & ~x743 & ~x745 & ~x749 & ~x758 & ~x762 & ~x770 & ~x774 & ~x782;
assign c9405 =  x6;
assign c9407 =  x744;
assign c9409 =  x487 &  x492 & ~x3 & ~x12 & ~x14 & ~x26 & ~x28 & ~x32 & ~x54 & ~x111 & ~x140 & ~x149 & ~x173 & ~x174 & ~x199 & ~x200 & ~x219 & ~x251 & ~x256 & ~x341 & ~x393 & ~x556 & ~x582 & ~x589 & ~x609 & ~x611 & ~x612 & ~x615 & ~x666 & ~x668 & ~x676 & ~x727 & ~x762 & ~x763 & ~x782;
assign c9411 =  x140;
assign c9413 =  x30;
assign c9415 = ~x350 & ~x353;
assign c9417 =  x287;
assign c9419 =  x229;
assign c9421 =  x280;
assign c9423 =  x93;
assign c9425 =  x318;
assign c9427 =  x284;
assign c9429 =  x224;
assign c9431 =  x756;
assign c9433 = ~x407;
assign c9435 =  x56;
assign c9437 =  x389 &  x390 &  x415 & ~x277 & ~x421;
assign c9439 =  x324 & ~x71 & ~x106 & ~x121 & ~x132 & ~x153 & ~x225 & ~x227 & ~x261 & ~x264 & ~x346 & ~x370 & ~x396 & ~x450 & ~x451 & ~x634 & ~x635 & ~x683 & ~x698 & ~x716 & ~x733 & ~x737;
assign c9441 =  x116;
assign c9443 = ~x279 & ~x289 & ~x305 & ~x579 & ~x635 & ~x636 & ~x781 & ~x782;
assign c9445 =  x298 &  x326 &  x351 &  x381 &  x400 &  x418 &  x427 &  x428 &  x487 & ~x0 & ~x1 & ~x4 & ~x13 & ~x17 & ~x18 & ~x21 & ~x23 & ~x27 & ~x41 & ~x45 & ~x54 & ~x57 & ~x63 & ~x64 & ~x68 & ~x73 & ~x85 & ~x89 & ~x95 & ~x97 & ~x100 & ~x101 & ~x105 & ~x109 & ~x113 & ~x131 & ~x137 & ~x148 & ~x152 & ~x159 & ~x160 & ~x163 & ~x167 & ~x168 & ~x181 & ~x184 & ~x189 & ~x190 & ~x194 & ~x195 & ~x202 & ~x226 & ~x257 & ~x262 & ~x279 & ~x281 & ~x283 & ~x284 & ~x289 & ~x290 & ~x307 & ~x309 & ~x310 & ~x314 & ~x337 & ~x365 & ~x394 & ~x395 & ~x421 & ~x448 & ~x648 & ~x650 & ~x655 & ~x658 & ~x662 & ~x664 & ~x691 & ~x692 & ~x695 & ~x716 & ~x724 & ~x725 & ~x726 & ~x731 & ~x735 & ~x741 & ~x748 & ~x751 & ~x769 & ~x770 & ~x780;
assign c9447 = ~x6 & ~x8 & ~x19 & ~x25 & ~x28 & ~x30 & ~x31 & ~x35 & ~x48 & ~x51 & ~x65 & ~x81 & ~x88 & ~x90 & ~x115 & ~x116 & ~x141 & ~x146 & ~x147 & ~x173 & ~x174 & ~x195 & ~x198 & ~x204 & ~x227 & ~x234 & ~x255 & ~x258 & ~x280 & ~x309 & ~x314 & ~x315 & ~x340 & ~x368 & ~x398 & ~x422 & ~x423 & ~x450 & ~x560 & ~x579 & ~x580 & ~x608 & ~x651 & ~x664 & ~x666 & ~x721 & ~x726 & ~x728 & ~x729 & ~x730 & ~x734 & ~x735 & ~x749 & ~x750 & ~x758 & ~x763 & ~x771 & ~x777;
assign c9449 = ~x1 & ~x3 & ~x25 & ~x50 & ~x58 & ~x60 & ~x67 & ~x83 & ~x128 & ~x142 & ~x151 & ~x195 & ~x223 & ~x235 & ~x267 & ~x294 & ~x295 & ~x314 & ~x371 & ~x394 & ~x449 & ~x616 & ~x662 & ~x665 & ~x698 & ~x720 & ~x776;
assign c9451 =  x30;
assign c9453 =  x281;
assign c9455 =  x67 &  x745;
assign c9457 = ~x591 & ~x609 & ~x612 & ~x648 & ~x722;
assign c9459 =  x316;
assign c9461 =  x400 &  x511 &  x548 & ~x15 & ~x17 & ~x58 & ~x73 & ~x111 & ~x121 & ~x172 & ~x201 & ~x223 & ~x586 & ~x731 & ~x735 & ~x782;
assign c9463 =  x280;
assign c9465 = ~x324 & ~x325;
assign c9467 =  x177 &  x316;
assign c9469 =  x84;
assign c9471 =  x286;
assign c9473 =  x57;
assign c9475 =  x399 & ~x246;
assign c9477 =  x144;
assign c9479 =  x12 &  x253;
assign c9481 =  x145;
assign c9483 =  x332 &  x333 &  x384 &  x387 &  x409 &  x416 &  x440 &  x444 &  x471 &  x546 &  x550 & ~x0 & ~x2 & ~x8 & ~x14 & ~x17 & ~x28 & ~x29 & ~x34 & ~x38 & ~x48 & ~x50 & ~x54 & ~x55 & ~x57 & ~x66 & ~x67 & ~x69 & ~x74 & ~x77 & ~x78 & ~x79 & ~x81 & ~x94 & ~x103 & ~x115 & ~x118 & ~x126 & ~x127 & ~x130 & ~x132 & ~x134 & ~x135 & ~x139 & ~x146 & ~x147 & ~x152 & ~x162 & ~x165 & ~x170 & ~x175 & ~x176 & ~x179 & ~x188 & ~x194 & ~x199 & ~x202 & ~x207 & ~x218 & ~x221 & ~x227 & ~x234 & ~x247 & ~x251 & ~x256 & ~x257 & ~x258 & ~x259 & ~x262 & ~x263 & ~x286 & ~x311 & ~x312 & ~x313 & ~x335 & ~x364 & ~x367 & ~x391 & ~x592 & ~x593 & ~x632 & ~x643 & ~x646 & ~x647 & ~x649 & ~x651 & ~x653 & ~x661 & ~x665 & ~x671 & ~x677 & ~x682 & ~x685 & ~x686 & ~x687 & ~x689 & ~x692 & ~x697 & ~x704 & ~x707 & ~x712 & ~x714 & ~x717 & ~x723 & ~x725 & ~x730 & ~x735 & ~x738 & ~x740 & ~x749 & ~x752 & ~x756 & ~x759 & ~x765 & ~x768 & ~x780;
assign c9485 =  x255;
assign c9487 =  x120;
assign c9489 = ~x215 & ~x361;
assign c9491 =  x230;
assign c9493 =  x147;
assign c9495 =  x372 & ~x642;
assign c9497 = ~x323 & ~x581;
assign c9499 =  x63;

endmodule